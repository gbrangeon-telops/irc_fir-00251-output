

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LQ2vJKYKktoZrCpK4juRqJANqbtQy3/ocOY3ZqWcaeltVJ85vibXAMA5tlVvS0pp5GAf58wutyGk
pEVV5Zv68g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oMuoQxHU8xamO4YIRqVhC5y86VVKXTIB4hGEIvLUCrdkutaN+fgAx1w1DFW4AV5UF4/dcrqjOzkY
K71n5sVp1APv9EcDNy4SK12rfM6JNEmec1W0js2v54algVfB410d4rZG0ryxf2jOEEtG3y1R1uZT
docKTvmf8ciwTam2vyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RwKTb0xAeUUC/Zlh40ZbRUmoUjB02ejSjmyrw31uw3LFcwmpLfrEGeQFx9W8nBY5yWIBOz4idUaq
fc3pMxhJHFC7jCdnh3Y8hC14pp9rspO1hZLfCOxHKu7GOhZZlRDfFJE9YTYvNMQlQ719mBEfy5DV
yB6StZ3JnfaWR9muuKfjZivHmkGfCe6IBabrX2L7+LYnKKp4Bj89EkuYxLdjSsxwwHL5yBSzQWsD
f3NymUlojWqzg7COUuAovEX4Cr2S0yo+Zr9C4jJ43pknI50nQ+b7CaiUKqbCSj+K5CzuK/dZ/FYE
aO9kMeHqHP3vuIYIBhuz7gnYm8SB2OlUmalvFg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yN6ERKfUqtxcEaZPhTWcKmh6+v/ubkhs44a1yogYIxw8eK2NURIBs5ApjPyj6y69SFt7ufKFYnlE
zs+yxTyZOIDjE0iu1eOyuLmYVN1yfs8OFxlynJLngPXQyLVxs9254patixjWMGwWk4PkkE6mKJuY
ZOkdptcpF67u2/mYpXY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t5IcFW6UoqOUfYz1GOxoQECi+9Dv8vBS33YPIONcGWTXCbnB+Rky6dyYF4Y8M27ZqAdkRtAsKEP1
XbHsYeeN9tcVjnhsAEW+ZxZyVmGkxa8lAjUHEo6bSWwd4akFKgw3xIpbktgKgaV0fLwj4wfHvTcJ
XEKHWYqSYc/CYMdUUlUPXn3ng5DzustWIyUHmy7pVesXYKHPGiFba8n7HX/7Kf+2y3k3y0XUfQRM
e1vWugHsLB14SmtA740nmVJ5TRRb/gYA8FobWc86Rp4qtvRHvVvYBe1XopHUWeY1WEaPGutqYtgU
FjBA3NC9aJ03W8dZxVcVFZhyW8E1aSZwJp996w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1517888)
`protect data_block
4jCYyQvZR2ysdb7IowijAXyYHO1u+o3TaA7ShyAsosVyPc46/pOhbIK98D9TBrx4z8oxMeO3MYry
2kJmzAii5Ow13Oc5dL8RoLIrXLY8YsC+XkGXtq1sAF6X7m6gwxZUr+XXI3O6c+EavXQEltE8l8xg
GElQrHL3eyctEWV0DBO+OQkJCl7tgP2Ol+Nnp4O+MbRU3B6mit44m0S/luXtRw1oa6ix1NtXdx/+
PKymx6FeGO08QnSuRXdq8L3no/d+Oas8QwvBNpyiDSZuYtINZlPHG8iVzcSEIr7olatQKywuLTBk
zMODrw98IPiglsaKMIYxJBCfzgtAxXIPQtEhDRD4cEYXE+xP5eMSa1InsTs19rsrx3DhneIZfR2u
VSfImvGPPIZjOz4AoRoREoP5BczPM9R8GqN6cUyhwdfaP/LmCihyEuSPFfSIo29bdA1D3/nDX350
6nJe70ue8wKjuOWu1wmjp/+e79wdQtDolcKryj1jagiPFO4eAGnCZ5+843YN7IfMofXslXeq3l8B
58+TLCb86PAZ6aJQQ4KiFUtLN4JmGHuibrwQ5Cgo+/aA+t9azZ7I6EpuB+kpbQStxJPoSDyGRgZd
cMoI5DZZv7By6TDorIvqgNVdatRxZ6d9h05lqFx6MxRGk+2lROzoKR1h1F64n0xV4jJ9gJkCktpi
HW0sMLREwJCq1zu2gGZe2u0puXCinH3QyTLcFncb39RrdeeonvFcNzlgbCuaZFXzrZvBATW4ZKqA
mBalczyOL1xBSXp+JrfrZVP706VbD/eMpN4/8zXGf1Q6m1WTsrTAQbEW/F+Wn6qfEmJmLzZt+Ba+
T6wHfudICNl0BGgj6ZK17h2+V89n3eEv8nCXUYOLxIL7dLumhleRmiFwFPQtmuyZtsYVlLGXJGkD
0qoUFMDiW6+qrTKCLlBI1tFTYt9u5iVsuMGbZpUK6gWTS+v1wmAArgPYc7aMFsStwn1xyGRBDerx
nrDFBk4Wayp50fFTUTGpuwpk1e5Ub6/LK6+OEel1oVyxhQhqoZxRlFDWbcJzxi/1wENHmCaeQIHF
Zm2RbwRCbom8agNJ5I82xtx62EotD2OazS30t5AeO3rb8jYxYuiDPWRXZRTejYzdm7PJbtMcu+p7
5p9jI7tbncym8Bp62aUDiKvH0VVMtCsw5yAi92XDn+Gu/tcOQZXd3vqwkxwgQ668yVHdUXdnY2MJ
1vs3KQlDtkyQWCv/dQd/mhPEBnAYXLF9AyZN9RyFQKgOBLxJWsRz15BXqdV4FNfgmwWc/1Q9eIpX
CF4SZMTxKvn3q4raYbldI5h1QZdaruA2gJ5PXRZHXcbu1J6BkacmDpYg2gXS8rN/fSwgRtse3Ey9
si13oOglXnvnPQssc3TYKBL9byzV8YiVplqA3ZM4vBktktoXfYGNLvXZJpKd7q4C+FgcgbYxrx17
qcvva4a8Klp5pOE0YTbH1OnWZLr7Fzh5whean4JqzphPGuYx4nEKuXDkkc0usiVC8MXiJgiweydB
HzOKCxsltICU9oPQjlZP4ryn4PIgE8sYpg99Pyyg1v/FvFWSgME7PQe0peWiJBXDo9ovXWcrJ81Q
q0yjN/spC/1VOpdcSqeqDpmSSeSziyjE/ETl4x4H1K2VCpvdsidn7rXV1Nl9/Cvws5qk1WTkj1a9
xzZ8IYs8XHZuwCa35pwyh3UU9pWodPbkByiEBE6WxHfmNcg6WyZIwTtf2qtfjuvojFb0SJobJWfF
0djg2igCKZ9B3FCJgTq22KQQV3Q3OP3GF2Mvudn+N14+Y8w4BB/MvcLLVddEBoZMgYg4tJHfNbTH
k5AvDDAWbGnARfC58hyqm1qQhjgPFm5U6md13tIefZ+j3lSAKT7jDvto9wE7XuOuKFrO3ingcNxR
6jzbLtzvUMJK9G62tiK6OBt+NYpSuce0bqIgZyKBR6LAatQ1zPn2UpbGwFw3eEj0c7YfGe3vxsf8
+VnaEhveSkl+EJHDIGLgHI3BIt6+o+vy/u83wdDpRAUPWtys6oAUCkqQTrK6HrslJty8S+HM5cju
UneuwjffB1eeulBwHK+UZNDihnNbDPvCrgvTN4TEApQmv74N1YEY9pB2iCa3mHGk3+vKUs1BBqt1
0Pje9es15pPGwgZzdS6u4qv9IHBNz/hvydyWAS/BExrqevERJQ9U2uIx9hIdVAambSi8ePTVv1FG
lsL2LdQKc2rG2lpz97ggUblIiuWkQ5R+OSVnYcXJPtAVCXnnk3LdJJqyFeZNLnAY70Mz9Yj/QvTs
x7WVU7ZLzTNxzCnl/IYmHE/fLz4iLdyyatn7/Lrio0BHi1r0rFuXCHFK8qhS13QxGUkFdJvcN+uJ
LlDYpP6CthUUwlVieFUQEAXg9ZWvFdeZJrB2cFKmo4iWzbwaFQa3CQWdHEQDIMlQ9E5efXBE9UNv
AMMUEprcFwqaALiWRcWT6HkBGZwpZVpAY+Kyy+aRtmBPVWF7cTK1XEvoJRyxisuV6IFJE0L85AzA
NfEdc/mi6HIB47esGVLAoiuavvOTug7k4lf2mGwrjBpb27k2vgNOmnL/39oWEaQmMRh/FJY46Puq
m2/JA/zMiAJwkOKDNB2RdDF5I/d3BRLwp9NM+mIFaLfXzveXF56RT9pT1TywbU1Zezvp78blro6x
ulofpuqrQvTTYWEy9lnimRTWTmx+aOaXxh2hPC5OQTaRukW5pkf33wYQ8iyC8h/ZMuTH4Vuh40hW
3Gy0ki9gbVR3hwo2YkA1wLoeS1BMuyQLNrfetxSXNjjMxDc5J/HWfzcsoIfV9PcseyMVyHigIR1Z
Mnl9poT7q8jOWpirdRStyS7xK9LyRD7XVkJR7vPLRUd/4ULACND6gBrHntZRm2kiVfHEGUbXLzGY
FUkf7hQ6qFEFW2/vmAp4oaicI3w+sHTqbcZ14x3cGcLqKpqrnlYegS8T138WjVzsd1q9mVs6kvPg
9TndHXdVOmyrkQErU/RjbX1svDrzis5SfJL8y4q0Di7uoBvPuSPOGiKa1ccgF1r8MmzODkTo1jS3
lJV21K4OIknNQfNXNKzaM+wwEROLFZm6vlWKm5UlNjbIZlDQcGu90MpzitQAXDRAznQYusPbcmSe
mgFDdm92cJULjhts3EywDjnTXms6URStJD+YDZY1t7QiWtakEHecPUhgbeU2bPBjSyJ7z+0Sm/z1
zntBj46EV2aToP26mAvnCvEtmTsRLGv0Z8C+LIl51SpXEX/aY52PtJN7ClxuToV7Pd2fS5JKYkcN
WzJvrV/c4/JklipnBRT+/pDeLMVOKYMqtRPIepiYtwGk2aDPDz4HsFxUEDpa5vSb71o7aqr0n01X
4HmZleVd3h3dlVqq23pMBTFQySAGY7MWVDaKFj4t/YDNmJxHm4YneeY3f/j/qmWR2UHB9Znmkq6y
tYvERAc0MH6LgFFTQ1oRIUQQlf8Xf/8cmjDUHrBzZxaLvwhDeJWssk6QVp6uKPSVPmV1p81a7Ish
93EyAhLTLOkEKtq54WaE14nGLPrYWvhdEdSrK2edtMpEl/HkiXau4oJA0diSdKkhK8eQzN5RmWor
3BRA4VCQicnPJ739A7GntbRvamxQ8t/MInTuOMIzijk5NC8cfbypjlipwOYeeh3j8SSHruDUgujj
/Eo/r8e1HyytVLGf53oZpJ47YsP1wN/X6XMlpTAIw2ArzVcx7vq+h15rFLUbDJtYZyUkBZxK7qR4
AWt9A8tgjDLRHhD/bq5l5C7VXwQFnQSreyVMrMbdfhEVR7GTfzTTHqgsl91gswFxwRfGc9I8j/Gt
/49+ZlBRhdhzDxz+FNf2IfTehRYPVPCOMZYsr1IO5gGE7LD/Lt3SHeuz1lin2KTxfjACFMOvBElD
tGIky9mKOkeezf14VzKhZgorxuMMnLNX07krb1TuMzRhXf77F3htzcM+u8ZDsu+stnRO3kFbY4aP
gKIfuW2CINkDk+9wRxluiv8/Qu0S06NyJy5vgD8wi2LMQXVH+SjIyR8CX2EAcR8Wo3KqgVG4kThQ
uQ8vbVbH1rBMGYbLvbkk2G8lwKKB6muSSqvxpky2DlxZ0ZC9BidpB2v9DGfXIj47nC/TQkkHxMdj
UXhu7yu2JajecbzTckdFepeZJSOmNiGuZ4ZZKq1gV9joEeUFUvBnGpbHveL8FFruDcZGMgbOJWbP
syiETw3jrwBHHOPuDjIXfJm2yZaGHu4gjR5pplEWkAnUFwE7wEgPSa0yHBbmWZ/Vhh2EiEpGSM/O
YQhG+nBoznjrpnBgTJdyhnUIhh0bh9gVMkg2vLFw7q8xwxHWZRLgO7pCc91spieGWokhy5rsnXCd
nlMQ+CoqwPJ8MW8Zv3aLFdhwmA3m6yppqGCcKnA+geXcxARuJravDUrD76vdW3h4WbhOXeo3yTnq
dxygHQ8tmslTYsePXEG1sqvLxXwDRG9Xmny7K0yYS3yMImGqZlyxX8fOQtGNEp7rKcqC2VRFwf8s
QX9o8CkikRgNbJPbFmjw/zS9IKEDvTx2byozFgLm8Kq/NOv5pgb5KMrnTw3vgUqGUerqnhAlCbZ2
35o9Hj0lvjE9Ozs8KqYl94YblVBZvpzGsXbkzKQ97Veu7XHlNb2BsYR/ZK6ZR0/71dXRiCNhcOTP
TWl9Ta5UUniQMQN3BWtMkoLpXlcZWD1RQFkimcU6JtIzdLABRwPdCjWMogAZSMibvFo3jMu9qliR
Orrt03MaU4B3kbFwlLiCLq/BWD9PIU4tk11K5ywvvG/mdp2S4JKYfdqYpdYigccv+RQnWs3LKiv0
3oaf3u6iMLZbfa0XwlNZjNtOKHZGS+MUY9UIxv64FEKF/C9xTD3ewGTGhZi8us3OVz9nwdRJP02W
TMMSrt5TopvD94o2bplGcZBPrV1b2CdjwPs4NW5KEFP7MD2xgLjU07FNtrIHn9QJaKM2TfqamaMK
Nq/3Cd9iH5sD/Stj3Z6jYXQptDFEunh1PlvcmDypPL0KkFsf4GUk/118HNX9oUkpOqMiZQUFFjE1
ioE17ENiOBcAYhaL+jS3h9qsXfpIf6I0XoyUWV5AloW6svEZYZiNEYEDBnI6A/WuBkqBuCDOgcfJ
eFEOurnxzvTJe3D0f9faIoh5ey3mBogcnrLX6W+DZ2HdkCpmfoVaM9/ZiDZOmFCGohWHJ4lbOS1I
v4TUdDq3UrNWnbGbSXzstVLVFr/7Gvm5CRGIyXCGo5YzTdpEt4DtagBHoybKwdgOuD2kxl2MsSmZ
p3mb8XwEqgfsnTOPfEHQu9XOcK5cOwtK730GOz1Rr1Ok9kovt82CBKbViwtPH9nlR6WqsveJf2Up
TtWyOsFtEhSa+E222VP892iLO7quy4ceuU9GEkI9dCj9Zulf7RRT+SulKPjjGFsCP9nzExUb8J3H
jxvv9uVSL8GTYqqlNa+EQCYUEd+g6LAwSCQLg1bTy3DaoCpUJ/cuD0zF87s1ztk2IeXKyHymbeuo
XPSaQHEseOoRCc+sUBagpGsxGGfIFvjYqsjw9NKjTtCSzsW6JHjv2+2mgnByM8z03ZoT2c7BuHP1
4VJWd0kWclIPYBda9gVgT2L1tDGw+fCkGB77WsNUOccyCOeYQcKLzlxsjsCTBBwrWFD9+eO/iOOH
n5Uhtd/SEXF1e2RDBR58nr2tzqxXd9OLqtOjNBLRtQT90Tfc6+WbM0GlD5nP2xy8fpzCt7pzlUFD
G+kCSIiPN+PycKDIjyrYo6Pn3iV3F1GerfJ5dJS6oFv6q84fOHRfqdjoTFTau5+sTPVFAsVGF8qJ
SToIMdb/NIEMk7DLSpIxjZTtDJuQrwtRjyfuzkqypbiRswAuTktOxywFB5YjqIZqS2tV9Qm5dih9
RFe2F0Hm9J24MNq04XmATml9fC19we/Ms96dRe+gZxRfWkLyv44n/CdD7Co024Qm+dMpPhCy4ExC
84FV/40+6gzLy793lm8b5Fzm0pN4DBLEpy6IoPaZ0jRZk4f+3+I+CbM5eIFLHcgpAxk2MeifPhH4
ADP5VuDU9oTedpThGL0wth6uWQv36Di9mvf9uuGc7OJyQZv07Lhr0Q4pNldtm/XJxXsGHwBYy+Oz
LVbjc7yp2tGIP7V5XmoTrpnIvElNwKerZU6QRoGI8lOo9Um6aHJPRgENDalbeFTs8gftlGzHMdGR
RfSGlJm10L/KNm67fPWkGM4RQZthkv50SI+t5QhJTpmUHVtLomQTc5olbfBOLT7tosWXyiFlLIYP
RfyLv2FOXk8hVd1nmcmUmE4q9Pg8/89ddHcRwOkF+gi6iGjz5a5VcmOV8eVepmR9y7U7v5cIq3PH
WrqfXu8C08WjP0l4urHjG6GrtOZa5D+9bHTx21DcUYOxA+sFu0nE8WQT5a9FDMhKoABDiqewWPOa
eELQTpmzMO/5uMq9+VEajW6Zb2eHvs08zX28eozMsDPeXBwkLICbCtisqtUbez/ScMyAOooKYV3t
72uNeIKYKROcwP2fNOf6GJs9if1zjH00s1ZqxmJW97c6JP76Sd/mxMOSvdA35XihWpfwiiTVguQk
ECqMJINg4Y2zziYxDJMGw8nn+lm1JyNIw/yNwMMcr7q/W2N01ppn+WOiwofdcMzfpxwI2m7yq5ZF
IQtMo663hrUsSacX6KorgonkZXI6o6mXF02YZRbaA59JZIa/gYHaysbmHBj04nqwSo5DmO3nDGmO
qMvA19LvxVfktu1xDVpGw6OlsJDfhOGx1iraFMDwqW3RWSPCGUGWHcAwFQTwXjD8ciNG4T4yoWlY
1Kfh8l4DviikOIZwTgPFKk3Jc5BKvBpplKEIUsSvvfXsEWCeFJN7uxiHt0DW/PO5YR6h2Pn4tife
4fdP9GGvmw9Vy51K1TuD3cCEAly3mxkprdvUQ/G2hIVIKoQRhZalCsE7GAaazO9P0YxzDXxFpgA9
X8RZe6Cxl/7hqwjsGv7bq3nX4fcK/vjYWtdamIERU9aNw7uZRhnZ3+tFegPZ7p4YMfCFksIOXNGb
7d2I/WU/jqb5J8ytsGkl7+GAdhlqOIa1mpQ5fDgYLz5iB+lcVtxPX7ACtRpR1eftl1zwIfTa6HnA
+NkmD4O1LHGmLlpLLZ9GKRmfTYO8ZY7Kk4aI7+2U/dxWsGn7UbOYC4c3RSW1v0uKzZ2bEgEkbKmB
+qVyhb/9yQZfuDoERE0B7NhbnIiEToh/qu9wm9fy7w8CV3K+WBD2H63Yjgbq5h4WxxHWXdTDmmhb
h0aunBsd/e3lDFHrC3vl9zR8ShJgolkR0ZcdAt0XMxw8AfSABXlFxQvQIbIAXeaLvfkk4bfjLWzF
CG6t+2SgvBZMwiQg2WcOvfnGg2hgYbn01GxsEovMlnUHtp2JSPuf9HmUsRjSK1i8a6NQkPhcxCsT
UaTBfttfyHgcm022PfvJ/7iWne8o6Iv0utrwePbxh2vgEPPdEeSmQHnipUFw4jN5hGrLUwLA3h0C
90F8SzSh6pZ/Bi0AYDGbU31GoTf4mbzm9kLyZJ685L5wGu3VUq6Oa8PqTIU4eIYKpwa9598g+e1L
Ax2tYnGrPzb8O9Xsw4O6lbkQlqAAAUOmz9vEQPHBCy4qMTVhUnJHEl29cSGjd5dOwIDb3rUBf409
cV39M3yhc99/cme98O5GWltnSl/rkkA2KIRX7yWQRdiw15sjwWKM7Hzt0YVxT9j8/jSPESwFxwMs
opwi4zWrl7NP89g64RPrf00hIX4piZUB0FhWZDgaR7lUUco8tLRjzLSkeu/+ckzWsuabX3v/Uutl
bxviirHkSiUcwmEfX9Qdeobk+KrmWFVmSBcPwT+iYIsx6j6PvDGw2gk1XOM3cRFw/TDh7Ns3gJJM
ljm6QPyO01FnM2IBennXiz0RgtUzlGBSQuuvkd0LxuQjdksjIDO2ziLSDdBYsaBEwDpHtYyhz1XX
zW5gAQuIvi77KjQ3vd28qqunWuMkFdY4Niy/UKDZ7JepfY5a6poRieATe/aoSvuzoTHpwt6f4Byz
G9zt28k/o6B3X8Dfp1KcP/bbNu6qLk08ksgf6NiYko7f1ssEdLOGWYukzoybhxiLB/dWCLhAsHDz
tRx724sFuVjo5GP4xT2/efj9rcXc+VQcMl57DlkcJkqVfd/rjn6TS9TyO9jRyqupqtVLOj1JwiPL
E9X0XWzOpJ2Rnk1SCUxn4Ls+vr4aI3BQkxu3++RKIYeLGe6dS8c2+znIgWj/ttT1s+86Y3pDilmL
g5D3ymMPZmJzGktUpvYO2OsYZnIVWNonQIuIzsdG5ItAPgeTQviqPNPLMvt11CO5ub9xbMrdc2YY
5Es0swTi0kir65Jc8TV3vgvZxRSfBFEDiWI784m0UYicclLaYvU3SBJ/B+J+CKttTzl2wJGX9Z4B
yQTqf7c3cPNUOcoBSAPoBHBEsbGPmCnj+8GEnczCBR8fdX5oZgl5hLs4gZ/6Y592OeFnvp2Zzl8e
4bzMnEaL2RyW2xjJbOqKsxAhSX+KcRO6pKNb289fSCSq7dIsXiIFTU7RvxheD/qtjXq/agjJntRN
tZbv/z1vN1ANkG25ViZ8uA/O00viWi1rlemMelvV48H+OIQ/VcYxieK1p2J3/xeQKg6Uwh8ZS7jK
K75I1gw8gQ8CIHacY779A/deVBCLcUTJDbPLfkiPUqhhe2s4lCQZF5defNFlPOu9BDgJOuRHPoGy
pURq6cV+3P1tUOEt+t+dPlE/dGatkCl0Gl2p2e/OQJ7U+KAlYJMfPtTxPJfbaOtRQAS5bDUhpEkz
1JTK95QkhIEqi+ndRpD0AQ8lr89CVQ64vZDrEi9rBSetmaFFF/fECwsOkC12vVZdpUW2JAv7/Q/N
UvelJdq6hDGcUq3m7PPg3Cr1iTCQcG30slD6zkkt+4eTJhKSyeQKbU55tcDe5rxKSK1m3PRUgoFh
WmYAEJslupUiKkekYO4eNZ2i9bN5WkJlvgLgJjCvoLoBF9RDz505XcMgxUZ46c/r3BFbcvp2Zf7T
jxDg6FNbm+Qmcjm2g89Y8Ar6xv/L5xldNvT5ZHsdcsQG2ZtUqn0Zy41p4JJ0v2QnLD1MJfKeBXo8
ffBiwCXg9hqkXgb100rCXzkok0VGwVmlTAfdYpbrVhUE6w9V2jijYtC6HU3rhmtRAdqAfH0H4Qxk
Fv3mpS0BiZyfv2pYREK2NAUZyBTDnawmTAGLe+fqeRuTRnSeUH8Qvk+QpgIEvLGgz2y0oQDKbvwU
ICeuLJiianajNaf1e56AUI1tWuNJFnwu9XboNTpRYE53TLyifnUMtxGk8MoBfohVuzg15FwLBrGO
LyE5kYYBp2AdKnRVvdFa4fmupccTsUGPSdFzOYLym28ow8Hr455EHl+bRLaHIssyJmp+HdhNqyWs
VTgAU2gN6GXdTPfcNtjjtgDdhj2kflflHkn1K6r9PH5o1RK3zZfjuh2euj3bTBoyvNKP9QwK21pk
KWNDxJBx9Orn6v4RS1ZxcSUItknnEtkKwQF8D3bUp3B+4cCmQzdpT3NlRc5W9PcZPeSBCKZm2YaG
jqCDOhdZlIAuZs+qKmRjzMiB4q/v/OS4q2TcC3Iogw3rCyNPqAODXZyeg07qm40ZKPX5nDcrmTSb
w0OUVkXwUhJzB2Vn4EmzNg7vKHk9mQIyCM+iL/Ltnr/M4SYrjBimunL4eEa0XM6HvoDuKS7CUW7M
ZDHM/kMcaMOA6uXfwW5G9L4kg1kf2Uig3gzfZFYw8vore1sP/h/98M+TXQgM1pr6SeHCTM/uAJyu
wcXp0Ln7KKOM0EgwgpxR+bQFW69lGWniGj0+D87hGi1a5ik2OyXcs8ot/X/Oqgp7g+ryXKIG6mGB
fLVEbolqmxdZaAoG2t8ZEJ07AGw2HpST9pZLKd7n+6srv30EORKr3b8iFzq03m6P63iYVBtPLYs5
21NDJv3G83P7+R4TOkrZbc67RN3dFu0Mxk2LsUskVHBHza5dbah93LaSi+6xpIpB6c/xbETUPOOo
OIDi4RWlm3jLuoZLsvH+K3T7ZJC7tW+uZb3CC97PKjJuJ1LUPyqs1D5KX3kdaE/3T5ea3fsl2wVX
9COjj8zraUiCJ5YYhVu7dXTDpkZEsFT/lOndxOrVz3bJ4WoJ3y6tCapTMZv6pbhPdKT1RlPpm0JF
jNJ/twFjWDca9SoC1PQHrJC4Z+LDtq6GzjT/f42/nCBr4hhcNAmgHi3BPAvxikuX0wHYuYNkghYG
v5OwXCOLuFEfPAulcoHF9QASIMk0Pd2FE33Dzbn6SX5v14kb4JsvwokLW1uMdnuvCd8pfawI8Bel
vu6scR/LV5fVQvsyE0TQ1PF3YC/edSRwbnUTsY9mfjrUCuhSZjbe1dwLAutnH5Z80o4kJ0Uw0xWk
ZlRViXPQIsxORmaSwO/QAo2k61THuvdq+al3EVd81V8N6+pn0umh9GhNMC503/FWknC0jCiDmgyN
vyigdJfWtyowG+nmplrXNk1G340bcVd4IE5BPhbOTJ0Gen7XNG6J8ghzc2JCRTEvm5UWsUd9z24z
Hpcadom9s7Lub2yyhfkzpcZBFDItNouylFx0AC5T080vOQa3z9ySCouW6IlZTtPYSWfrpvU06ZRz
4NWPMOC1yeZaDWk2RcmIfN9DfSiKQ47Aix7TH+L6mWV3QLw0jOWvLckd0GuHKrKyGGlPSuw5UhS/
Id2HzPuYty68CNYyuinKme2psKwqHGqYzN0y5Yl0jDfWGSFY3k31dZS/RvHTFjxYI3Lu8jQhgWmZ
/IUl7Vkz/jWN/8hmobza2c/jQh702iP8zT0c7DpHqb63ZAti0AuzOGuZ+EV2aladzc3KFctOADBp
xlO+mXfhuCPsU9+JU2lzY52t3hKrVY6gA9IDNvgPuUJD9wDHbj33wM/orQZ6e7F9qu34+XQVxlfh
Cod6lGSbHLqWuFo37Z6TdC6vOWxeYe+xIFDVbHYkkFoY1v+uOqFLMQh3gjiJyy3j19HlRm+GKhqo
vyehHVnH4J/UdOUN58Be/p+6RcfxHxDy8drlWRl6CipW6vdauQqf0A9bpijCyVXYTrZYn8VVzPP5
3ZKRotOGRS9734xnfwEKso7D/bnlBFh38wjuRmjbtNtbifmotBWt1owimMg3HSi38/EEieuI8wzZ
X9gwWhJpKpsiUqCE8rn3tkABeqWh9JZOBAyDWbmfVrUIW2Lb5Dr7/kU2WkCnMWEUIdbkNWmj/03G
tQN8jhTEdJWe5gngDupn/xRgxw9yMXnlXFSFv/rfKMm89mgLugOrnoOYy/9k0C0SVQRxaHRtbFVX
MIHiHvGhlvwUROKnazCWXpGMVlEOc/AGexORXEX8PszVK5OGkC0WQjrTfhfH+PBEaNtP74EeMXow
Jn5hg7mLYrfC+zyz5XGNEs5eXzCzcpqgAeu6zm5kwO1fidrlWIK6hk3mHoqFkQ/ySfJ1XuUaKpxd
J/F5eqvxlULlsuJedNL3PkBBa5xwMIPDAh6G+MALk2FISDTsMqHWKZR33NBpBbRxFMRIgjaCa+k8
QJSUyd9o6MnY02MtfboPe62PjEYGLncJ4cYX+H1EGAZH1F09OiRDoUiyh2ojnj2907oYT5pel1pJ
vCeUFEblEyBD7lXVYMuRC5hGnFuaAKsU+9qIW4k0QVuAiG0mcpTprpGrM2XOLgF39YuYfjfmoyMk
7Z40HTAMUqfdAcpjACNBem/Gp+cccxOEtvbiKzgHfar71PvisHYgmpoh/y4vtqtVNK52QEuGOwJI
dOj89QIr8jEvOIAegLiFiEkpqVSlOvCaFRQzUbAKkvuWFdabdS7RWGj7i4L0p4ZaZNdHtoqxl6IU
rlkOfciDgIOw1kFWPFmEYLPAE/oM5ACoVL+JR/riOwgDp5nU5kSLND3SjHbdly5Ie6Eit2Ek9IqR
ueYl1bERkwulLzgv8b1158mZJcatHEWU9xBci59GR3QZ5wwfA2H8Ofr/HMH4emWEMloLqbZdv+bW
BfnW+/NvowiGZh87mWPxhDwavFb606Ohep/lQJdl0MC3BU0SX6p6u5rrRn522bxLvGPh81vdk7kN
btq96+yZGfaV5tXWWS7Wl7pQVeAkfBoSsZk8KEXglWLDb8q7W0UBUBkofmUXpDQrceID2jCs5fOj
MO/hjxHtmlYjOoGCZ7GV+jxD/UPdG0TX6q+jeRArj0ma4nt+pl0ZPtMpkf3LU0Q8fXij3qn7JdQx
VJ4XCpfYsP2S3LID9edhnwRU5StdUXwYVUcLv633KWnbLiZlcd5/tH9Io51AIn3LJPUpJ7xMF9wV
J4Y4Sx/DULPUQPQF5w2EbG2cNRXOd0dWJpGba7SMdzodlVuzWDf2v124liT2Xq7fFCcTGCdVcP1s
fgTxc5QReiRKCppoHjELQWml+APKHHd8B842ibNVJfbL8EbcKidPTuCl9EaAUZ+G2QSxdtHPS2x+
ee1MUYhM5jGeoDGBq2zAqHBfh0SqlnPqBQByGyvEPTiev/qdTXvLgmTSGWj/l0ZrsNMde+jf1Fks
xixIi3KcM01D7fdV9prTevcJQtHK2Y3cVktz4j5Cc4L+pAqxCkcYUPHPZJVdwAdb+UgnY6pZts+v
RJpxeLgtA6yh4EctKNttsCMJ9dAI+jrBn9ZOI4UU5ul7i3/Z0T8PDhhgvS20JdvH27TDEsl3TJCO
VwZnDuJDQpIk4foxlX15gx1kpOi/9nZnN416zfy2hw/9vAdCweCyhWQGZmsghP4oeydBZVLdxyZj
7I6I2JUkeld7vjkMbrNe1hdhlmDaOazIKQVSqb+fXJGylZOTcnQY+HZZaR+kcsW4c8C3pZLC20Pz
i/NHttfJbVPEdWMsiFy1szwZPW/Jbud2LrNLryAIJpT4WJ9HX3QMCMFHi86CRo3KxGwdzWAETZjk
yMk9m8MAB3scuK7DLmvRBnas6AcqpOAbnNBItWPnKrx1+lO6gYKElHeL5TD9elQWHmsCTDO58DuS
Th+jtzoPqQ+ujO4fpGgNX7KPkfH7dZBumndlZj6vRE8Zv800yFtvIlpHBWvcLBqQdoOHEid+0/A5
47caWPpEHICzHm5jO2kwQgKZNp9Qy7mSO+91nbl98RIoRqSF7wNijHQVmNjVLEnTUmgODzz/5R0f
bjIVFX/tKsGdWgDNrBLC4pBvIqh3tWSRO3e+TmqTmnKYzH/8f887YbI7t8l6sK4j7kB5CvnP0td0
QR34o6A1gCPLRoS+oYWCzApfaSnyhfjTcxPgTwNVeoC7HhV407vMoJCVCHMyDAfUtDmCRMMqtQdL
p6IHWaWPS9SXgxctRTqCXxGBdSaO1mGsbyOhb2u8c6MxVsIV26kx1XquOmt4QtOZY5fHZLxJWRRz
FEf76JNN+s+/SbRBXTDJsNmCnpkafWFGWY9Ls9/g5WVWr7xW8aD08Mumf1ajHtifmZHdyE9i8JfG
BRoH4e8sL3lneFDpF8AgVS29+x3c7Dm/YeAv4ombmPhzuMtHjUO28AlyOnz4hx/XOahmMCUoL4ct
0F1H+ifhDMdDGrmn/JWvGFBHWk2ktJOOrgMxhgnDeXL+bnBFreS3E3CPT038RAMDaBYMZlamKO2R
SH4Jx3fgIdni2P2n9gHpvg+MzlefbB87uVoRqkFr9I3FjH3fVlbfmuiORYDp/at3pBLb1VG1yArT
oDvd+xwjtRXMVO5IsmWXf/De6RVQbosJf80hCC0Vs7BAdeEvm4I23HClAp5EkUWPVmUsbVimhdBW
3yWN9BE0VutA2PN6GQPddRuh7E8qXct5/zTnuA4lIgSgFlztFbCze+9+ve/Lwh0HD6E9a2fl/wgO
aqZ6agoJQ6R55yc+2M8o/B7vbK8IkBWV6RbKN9SNkEKxSgn9xoZmMnO9UhQPmQWjO0iwKdyQTubs
fw9AwDEvmd1FzIw0HekSBZYhuA2YOC5QLoIK3Ung5bmJXWre/DTsSG9vFryeIqoTS0F5N7ZsSHEl
Cgxs6b/7jQ2Zikz4nOE7JBct43d6TG0qTVh0ycsVU9n8shkl6euqsKgx/v3enw3HfOvJMSEHJ2Qw
s/no5IJ+uueOuLAzgNlHHTm11FSl0vI36KMt63Rdyjl9E+QlQKblEGbMILJ+JUMMSwtQcTXZgUVa
TT2QgpGYlwa9YAE2uWyEd4+Zc0nHtOzpC3IJz9p7azZTfqIcK3XtNxKpL1+ibxehhLKyF0lGB98q
DdTX1T1ekoltmGDwUeZAqaeTO//J1kKOXCHRXOF8S1t9xHuqyzZKAaE1wqn35gbT7Q/dXkgDKKkS
50ogCtlysOysDOrzoILz6yfxktZR9Tcbq0wdNT7toMP0u1zHdKgwKnCZLsYghh3fLQOFTKV/haYh
yfJG2TBzzOzR0G/wWq9drOX2nyOGfTQ5wo9KxUTanOkCLuLxuOkh9Ko/H2LLdZiGZmXak5Qgtilp
ceTyQS3FXeYdLw5sFHRL49/9mMg1dnhru0EVyBJNVGrymWr+9DuX41AzsdF5i4SFbJgrj818HEUx
OpTIuzLFcdnMQVTpoeLJsA63pDiOGqYp3DNuOtUkLbeXRHMa7xmNNxIVzL+0pDrXQOXC8X2EmGvT
msqkU9+epESSrjGbYzSTwtkTDL14O9HUqYfOlngoxfQB0rVYih5yvuJcKa9FZ54DWTmBLZ8uNPTh
5SXUI87qGpCWW8f+kaftWzKnBUU338q+zWKaYg/V/xq5NHaK8BLQl7Dqdl5sf7Xc9vQGZ36NoWS9
oH4547hrzL9hT0bqWOLApvxURapyAE52HacDfSEdjb8eSMlXKIvVoCx1bnp0dznZMVyCkOItmxES
LB+v0TP8P3joSnuWgPbVSulPVD8LAuGLZYC24FN3+5slez4GKpJHZ6kiS+lpZ4NImtBKI2Rx0hmg
Q8aA8kX7bpgKk/nh+bzibDYm5VwAnmTbrplH/a+UA83/SZx0nY4SIyKtcIKwsCZM2/2fdrEbaPzk
XKgD04UrK2B4HPlm+Dlb8yGb94tLbqX0Tc2/Zb5eziE5PUfqqnhhlas+AtDAs6EgX9o+Qr57GqTw
UJ793UBsjY7uyWzEVgd8ANSq877KRz6wmtFR1S7EazJA6bCHDTTf/3sK8Co6i01bUYR5Pf2iPOW0
kqqhKER7ZwuiIXz/LKjqkjpNLVLQrf3hkS0+f7uSe9vZVtfMUuuG07b2OU1stOvFmNQ+FpuoqskE
t2aa8hvSvg2wCpvwErif5j0lpsueD7WsRKjAy+9oNJNdAwqNzfPgnQKVeT1MXVPElZKAi7A1Pw/E
55z/QdY7vAdGh/lmo7JwFiipot8+rrGn/gGikfE5qQQOKOppeIKSaT1nAcdeSgpye236BgBEnpt3
V9Txrj7prhVe9o46JvZLIl9NIGV/IzzplvDxqYvPFV9oTVyjT/rMCD5A0zdtm2ZHyfdJWj7IE9xf
FOlwikgHNWogcoR7GEHdQxfqhkhh3iOqMKXZ3XszviGIFZcuh8waONsjMPo+ksjmkbjtZyreCFmS
4xw2Kk6MFRduSzv2RsdbiXLao/j6MQNxZwDSkUcLofJu4xr2aTluz5Datd4mCcOIJ8JZI3b1iUOu
er6t5H8U6af5VnlmsouFYhq8FFxtu6lqhFJ2pLLEFGAGcurSA4L7yWAsHnpshfr+te1GpPzRo+bW
4+3wRjEiWkGCqETJ7SoXV8AQpU+N93OZUZlfeAVO+VaxFg7VoPKIJLSS240/hnEKhNEDNOMn3xi1
zB+E6/F1r7jzh4msqz3P/8zh+rqRNwJZVWWaGlOkZXzhJRA3QTstNcviK9GAuK287tC/QG09EQyq
SNY9go44dYHXz/gtU6ZN7CxnDXRoT0BkZWIVNwb41u3ltWsjmnjPxI/NKY9AJtcOJCRXwgLCS0A7
7QE+8CePGCiUI38w6hlZF2+3PH1uFeyLaAbwbUaWs22QyK8ZAYxv2ImE00OIaPS09jEDQoeVAjT1
usCDRDLmhVz8jIU1VAybu0EJN3dBl4zYMbaxLfs6UaelX8+4oNTsVwG3q8nwyOgIDu2vtvu+i47/
8MYKCzAkaXVx8jdzQP7tc+ZUhE0riK4h2ALSwvHmv3wprj83OV57FFUUQPoLrn/Kkzj1rGM7sRTz
L49KH8UfhMWsUxVMWmtDFmdmPgpFBCC90mehWAXOxMnmx137DpaQDwdVmzK1679cLMKjG5eCJbrF
kwgpvO/pjmpR3i7JpYBx9fNEeyYNUHV91HxuYlp0s3UqPOz+XNI/nLois8pGKuj5W7UGtNv3HGu4
PmEQXyNgj6ydUH9yNiUjt4rkcXQK0+KA+hlYxWaxzs7R3NtOSRvBq/zQEigOKu88PMjs8KzNQOJo
EEygb4/Tg+LMxOtDhMihx3GrVaQvVSqjmuSWX9nl2RyD+/sgtibbjGV8QIyTSs2p1QzEwXS8Jvo2
focMCisjQOLPAaVFEAZVr6Ss/tgnhB5mZFmbnrS4hGnv75+ZmNI8vHVbIZ47Dnttth3/yalzQsT3
fpHOcL97goYHOqREtGBj1po2hP/SYietZWg27cZuVhE4NSsr0FJEg7ElvOl2vuLEMYewMTM0GBBZ
tjGApbYWTjNVVGs5qAXj4GzOSNN+Rf4GpSMSmuqOvMdFqz881gI+UlsNKXEEheTFhMwjdJHq7YCz
iKumJNA6yL8w9cvDCLtRZ9laOOVwkSs6ReUh4ksFuuXu/+O7jz9XyYZny7bBnkTf941NmfVd4YrX
MpkEaPSvDbM4cPj+/uJ6KN9TkjJQZi5r9Lz6awyXwLUc/F67XlGc1tyjmd+3F6rCrCN9fdMtF6Ss
LI42QUCenAz2ORk9mqy6/TgH/tGp5u+qTUHKYo6+WgefE7JC8Hkt5+SVYZRIqXKcScdqXPlSAn9p
QiLNtdTArDcYmds3U7gunkrf0Y3EjLZrZrwI1KPBnr7w+7OJVqrrYjaczkyGyA/+cW+U3RWwvq1T
CxN8tSOR4ilWjXTWHseD+aINLw8g7xuTV3omT6P0vWwo+XMp9Qs7aA/Ch/Eksy6bIg5R1F1Qqkxd
fTKanmPpyZFSujm1MSo9DqhoZAd99I7BuAR7b1trg9yq0PKP95Wpx6Zst7Yk1VQPGcr7FYAM0x3J
77BSL4f0k9UwYBBXM2+cNgDFdVy5zn+oLXttVe3IIVoD9S9e1iv8Dvo1T3a9Ul+Ptbv7NU8GTSAL
u1cHCKcWWe4E0apPhMIFAUFEYSlmsy492lkc8vEazfQiUa1Pm8TWHkm0l9Okp/5YIebC3xIrcJr6
8PX9WW7fQIk75LFs77d31g/nOLx239d+ffbOWPujQrrhO1M5kjYrfhlRzcewioHY4hPUhIaDsa3l
s+VjQtuDDomLBzP1MAXvkHhO7MApfbcpsgjxJUvZkxrJPXoisAX9a4LZbB2QVcacaVOV4CwFTru8
nZ9JpL2almi71julLTnqlsWNrSDwveWOtVD2CxT4hCyGEarksU8Jv2TbJ66uKqhWLpO/bTNrT7qk
GCYm3GKBNc/k67uWn3oPYI3mKl8ik+NinSHy71YZzzzMUVIk3du1tHWzggK/V96NHT2yUqZ1022x
/R/t1lW/gjde2LaJQ05ppv+fmUAKETZVRMZHrfSdaUVsmf66jt80b7mW92GqD1Ws0OF8H0ZwFasn
XpWXStWa3/pi82wb/mMixeNXcTL5QhuNqDtLtjAjspc51qBqbLkutSMgzykGYm1sKNFzUodKUqgV
vhXQblKMWiRiIXbPW8CCsqoelMsCt/HRF1LysnuHjpBr3OUfVBLFPYbhHn6jB2V4bLNNeaZ23jsY
nNokAIv54+diEQp4QFMFbrdMOO2/LiC+k1j/BRb3xkThlNnIPfp6lI1BoZtTb4q2G0hqZMb8+ATb
n3lT9KdK6g/qv8A5UKxrRaujI71PlGlxYnYND/uRx3INPjILBajkPRL36Hu/Y+4+pAFwYZFH8v+w
ccx4LasXd7wlOGmk4E38UuNOD3jfM28hKRNKQuSDR+jUqzztmtrKoX1hsHqyn33pUzNbUfHpmgLh
4WPmBOHp4fCp6yfah59JZmuRClJ9THYn5N7oiOJmPTh7c6lobkDiRIlD1uJpGBPWcWiVb21tdunl
wTi4LJ1ZipeL3B2A/ZiXYMV6SgvbnIYtEzp478i8BjYzWgKG4XehPOY2OuYdKFqriZmUVRGtBgHB
DCqAL6j5s/r4FL2OofGMB79FiMI4PE2zIahSV+yzD9QHl23skfQdH1+hllOd3IA444x4CoTOCRH8
sDStB+UCnSmXZpppRgKuFr6GsOPVpJYkLeDe2zI0xCwq79ZfLBShX5OHub3LmHxsK1WneoKPa07N
B7jec8lx4lo4HxIT+qpdOW46aVG0k3z1BaN47mvi6o3/XkOrAxyc2CMocBtGDq9LpXr4XAN4fucq
8F7lF9F1PZh4PMF0X0FHGcc5Duns48joFOnsqKQSpWJ30xwQMIKGFyY28LcKr1oL40vIC8dddLSm
rie2UsH5dD2NdMMhlIyL9CYmpJ/b6VFtsive0A5zQ6tP6McP0bDXRXJAXwdRBQT9K1fYeGjU89jl
DtiDlWmnY4fiabXhXy/kWLvmXPvngOOd8VoWu0pN+qma7o+sYeni9h4cnNKBWAH42MlNK41p2Pdd
uPetHM3OsFSzDUrI7+r3wnYCy4XhObBBY2RnTQskPLtkltezIqcv3yrFkqi6gYixabjnkfNHr6oc
3SaQS9kuSFN0KX1HtWiSGT4gNEsVlpokSQE5K+zvdB1GtdWj9Gz0R3Gd+MotZiKpwlffsqQnOG1b
MpQGo8GJTanxlRxo7mOEk9joO49I9+Fb9w8LJmFMK6AyVz3J17SNBQHfDYdU4pvFtJzHsNiVkETJ
/LLx7af/tcVrLE0dbRp/l2Sjo1g40n6Ojuj58gekyntImZEiTlXa8z/S+ew8qSZj3/ibTAFcAWE5
UI7Pp/fmB3rzVKajf7zqaBOUcdjvE/6tKenDCVZTGeTeE3WSXHUbeIfN3ZvzQvIjBFPbGFu1SrJu
i3QtxyhiWCbEqkcf3UJveI5iH32QNpf2Ybc1JQ1uJoiGBdOHjKUl6puo0byQ4wYFtoVmz0E3o7X5
KSyTXm0dBBsDB5KiVm7CFgr723f2mbPKkY+dww6z5PhnnAY252tWx0hmtnLNW8yO7/ygBDuQziQ+
ZULt/seOnybIAr0+ZasW4nm+Xbadil9WUW5i3QrXTa9ABulngRMyjwVrmTzxWVK+ga9k2sc4paIb
9WicIvPwu0jWMRF51CMVFkT0lPLlb1oGMM2ROA3kpKNmOzMv4jkMUwz4Sq7q0kuxlLqqwdXP0xva
y3vd8FJOmSIDwa8M9dPc+v/YXLm/oNeaNfJuAGD3wlX10i6xqHTdMxiYa70lBWPoK6y8ad+nrHDx
ySEdlAQp0/6uxqOEt6ZVPpPcHCgCevzV1yWjYo1OB8BaIXlWWL+S7JM9NLjX5/3XUgfrP2pgtSgA
Lq/smIzjM15VZfrIjJGveUjG2ovV4Ow7wXP/+siSgkaGE8G2UOyrt0C+tGi/96GTDGPi754F3gSL
GHIWjfG/o7LAd6737sErlrPVFuHa9bNtYGIIVvuOjUxPb4f3PQVJGM8v9KMFm464hV2Ugp/5TF4u
XR3qA/9yUbTdDf/z0DUXHIFTTbahX+cXeXKNawpdbZ534XVzMbxNh3+t6C2XKqy6akJTsbjEvCFf
pa7qZ0d7GXYU7pxGAA0KyCbHmeX5/UwgWAdv10gB6r7c0Ax3hgkNvQl6qDDdT3Og1l1pxMEh9UCz
anrjp5HPeZToS1Lium844+0UpuMctO2keOuXSm6TxI02qsE+ocQBgmbcV1kxv4VB/LbFhkWHRBOg
QK/YOEw8x6hdvQ9ZUnuQxo6SY9leweqiAZEKNm2KwYQEKxcCq+GzA/VRnuW6wCNh813MJ4R0r6Bx
rqAeHbGdYyF8jEzr/k+qUxS3vtXQ6t1aRvZcr8WbMqif4+z1vRf2kVhALVpkV3cZzKdF4COxOG1b
dQ0olK34Qpqkq0Hv+hlLVAkepg5vYcRDvL2pHjHCjKJ4pSdMxNpuWxMt9JPOA73w8jfgYH65k97R
GWjyIrd//BrxBHZ9jsqtVs7agXWInyOX92oEteAKzedr3uAxSktblCpzU9QOoSrF0dxtu8GaOjmz
+G9rwzcUESw8jAgZUuU4biagb3wVaUDb82YuzQcqkOXBuZOqNk3FFqLvLl8gJEibJ9Lu0OzApld2
VQ5CNGPM+wR6wV4PmT/JdnsqBGmUIxKJvr4CZB+qLQTM0ZuKv8iBbxrSdRlaRCu9QB+O9oV8Zc+/
UPnunS1K+3Xg5IhynrDGKpHqhalXaoL5urzg+RVCUwQHMfWStu02o/1uMw7xrQN+a6+oqf0C7vpX
w+XA8s40FRx502/WN3O1II03QP7+rkyVq9lSSJPCkhy3JRgkYW42Boby2iYg8sXNHYNhkzb+WopQ
xcBorzVEy6uO3kBkGgbR98DTolZvtXjQrl4L8RhEkAqZ6xgMR7RpKwsYPmQxyx//3Z148JhQDuLn
ywvFkF9gWCvNizqkTZImIj+nWqgc6eMbQM4s+EYnLUTXqT7i1xDTsgQCs8JCW7Fh0KwsAeTFEB1K
LG9chFT8P6Dm94ZjWCJT2OMW8uLN/b/yX5zqG7s6c0deJY0YudILd+2tPyTI2M5xaS7GdPdaf/Xg
HZQFn/7pY8t+VVNJanVoFgxHtA6efPlx23eH4YBdZnj/OAv9tajp2tQRoFwmJmHCKCYpd4phhz6S
fYlpdVcCo29UpCe1ysJ5YEu7mRicyclOxTLi96f6vK7KFwUdb62pMnGepeLq3gd1ifZyN0SyjGzR
c3iiHMVEIBr8nJszMQxZg3XwtFjvR7aieT34xH7W3CJzB7v+tgIutCqUCUte4rH3bHeMwj8yK6cp
9SYtsJQLZsDGXLJOBUUHCChu8KYdvRkd75wC6jLOv9J2pQ36qM8QWcQ6CpjCR2pY1AfCkseS9PGq
X1C2bO3r6gWVEGSmjrF2U9AAK4N1tylwiMTWYRucbq47gqGEEEA9R2OCeApsxkB+S+lgtK/fG5gW
a8aH746diPXV/N0RaWXziOIxfeKSqWq7cmqRlMLMRveIfq3AEdH7xjMtRdiu7uByYrh9Gv9VDn2Y
XKlqmx7X06ysDEGtG2/FH2gxcJsmN4VOKo5OFVqfOa0kj/JD5pDobasJqGE2EllPZJjXHuKreyQ0
Z9M3KwwI8z1+pjJxe8fdJWZI8k/RWvy8nAz4RI/yL0CW7gNL3BMUr2DjyjSsyDoMEE/mhuLpHkxt
RKVNQiNoZ5B4HT4Ad3X2Df7D/9UaKWGO4eHz4+cSz24aF5NZO5PTQAYj0psvivhf+aN3gcEaTwoH
+f5wYRLHZMemfaRnCAbnbcIRfDqwbYm2cRK5Cq10ZTAU6MfyfiKBcsa6/XF2UDjzU4bBi7+aEwVG
vgn5UuikYzDxsYjszUDL9+fgYIf8pn50S/bOtz6Ri8vy3BTxSpF3wIZnrSAgfYPeS/SeJh0BtvAL
ePinjQAOZCh3HHfPW8ahM1CC7plqlKaBTbFXSfnNpoX6BtIn1u07bmhOQKC6MI2yBfkWJ+aREv6X
jjmI9vS21REH1oTEqeafjXjemUZNo/OczeTlFuy+ixZIGe7OYInnmhLGdT7B46aVu6YWTvUi6y4s
cWpI/KYB6a18HilvCwO1Ls09rMyFfEwW6eD1vP8oNFF5L7vuvetzpn2fihhLhYjpdA0EqSAn+Lf9
8genZGvZeIn7g1q5a3bzSMDkWXcwQ/kqsioauqhg0431/FqWcRUIcqa5lrjahF1N7zQFcTyWqKA0
57Qs75k33a8/l5Bv1dlN5hinrrtACPU4CFH8Nhg1+NUvfI9lKsinms3bnHN1IJcOKNJAh16a2Jev
zCtKtD4KYEMGBFB+D8n9WAbf8T+wezCNsSFx9TMs60VQZr8duU3Q5ki7++NFg5coIjru8TC2c/JT
ng1sWph9g8O1S+wtz0jXPPpexd8xWOTtatcnWOvp1OZL3n19VJQMgUFMEliQ9epZdLfnWBc0TOWu
cThUiJkbKaDUi1rwXOj5EvIZ6EdRfOiwXsCZuyza9Ujr3HDpL3tYgBOwHGL0ae04fq9XC83SB73c
nw/mGZKOMOVx24O09h5iUsYVKkp3TdBE2ywssWjsbPZ1dLO9DE6w61rC1XP74EWCfM4YdbAkQVbI
AtmjRMVUl6kNrs8hY8hV5AgqVSm+YSpRDor1BzQqfMXbCqxcKzZfdL/9LNf/FaEkwLsS4BXkANVA
40YIbQ58NA1+h2EuZ+fozTzYH04ysQAZHDlq61thIluIvMMCQPtc2jzWlJoa4X4sMchlbuVcwWME
hIL0+W6tZzRw6ST6Nl86X4nwgwFnEgfIKrO9fMJ1nYnZdc9YXCDPdFp3wSGIR3T45DAXDoYm93iQ
TL39xnKbfryenqjNwCuenh11q5r1Hzh+w0OfceACsILnpz7pVtImbli6Ij1B435y+AzOYlfTRNT2
dF7Zj5E4XZh1ovlRrAck2vdmxWzWIjF1ltMaOuzPf3dYCqzW5ODUZUg6+PIYSc+zwmfvrHdr9B0O
3kFWprvglCAL5sf5HKEpPQuGNfod69ejKfXXdJQd6U5VIjiSFNC2K3jzalc2e9n1fgAYM4B3NrTy
sxuKQ3ESBm6ry2UCHTXQhCQyTT0Ej5oKWOJnyuDQS9+kat70tjPss9ksUsZyFK4ApTzBwmtFa1J1
6Kgmttt8GX8DqFUBNgzTNVHfXO1xlUnnsXasQ8xlgjeiTfeakrnBkNc72EhqApsJcplG+Wxhpfuv
IdoddZrKckjJNZke2XN5r2wkpNJkQ3FxLHGTVHfyoIoJ95j26n9ATjxlqQtHs0bQ8Tt5Nys8B7MR
iEbDUCC1CH9Oiq6DsYf71h77847fmFFaxcbvsKom4y55DvAVHuFpfA+8ebwlrIb8JUaxd0d5w7nP
zSbzUwtZ3RFPSeZ9qbkYKgzhtWEIip42W+e8vGy/BvMA2GX6FN2vxTFm8tx5g+F0VZm2299zdENm
32AR0iJo/WFMRGFTze6z3xUPEpQ5ToWgmyzJVp2uNx07A0ruz4kQVVgognMP+Rn5BLn78Jg363Kz
2+75BRs15WCs6SXPZI2y9Y8SvYf3I2uuETK46vgZXNARVlXy3KHJFbPTcPmscmF0JP0s2Al/7ngF
W8OMYhv4q8h+3HVGIOSz5vGIjFtGGI4GphdQKs4m0l4uZU00irN4heW6Uam1/RABL/xSrqeKmsFo
Dn/OqQ/lZwjh30CC8kkTE8kkmTq9IuuCKLytZAm34NquYupPAN93RKQHgMTsNT6ov4qft1u7ZOUd
sQErb+VbWCbm35yH9RzAtpyZuArXcwJ6RqKA2l0aMO14pATA4Ma8VY9247U/Xw9qF2AUGyvhcLao
xLVER7fSS2FwMrYTUGxdi9AYd8NFZTvXnwfgg3wIwseNOOjpYPEAblVyj5/hhh1/cD2HZSxt1c7+
8f7o8cGJ+yRySQMOEDJf7ichH0lQQve9FiHOVlWyQMddxbmuRplUlo0YUjKojbUY58fVwR0zZZMp
0/yHgZ/1quQYSMJUfOoATjS2Fmg0EcdNZg0U/s4vs5Yw9GUnpnSmJJmihGMFUnza65kcyr1pdBuk
X2FvUr2TfNvPWM0c9JlScgD2bHQd686OfkDvCkU0cTvbpZQx0vZRNU4fOTHfxj99/ytSTi/tHGOa
aGzp2PVZY/+BjuZnZ0LTJxmzI1Xh3/qVwduKyv9uLwJ1aKaIoMShMAYgWJQcyd7kbq1DBo5uAefT
YcY8PsC5SWOGuHSAtPsZm5Kbd1fJ+XzMMO63/CBL6a42uoaTadUjsGUn4v1tLqhntxlI6lAC2iw4
bDxwRw+IsxpG2w9rXOQeO/h/gWfOoyuTScB7hyxOi2SolSZ1Mdd/b5/7JnEL5e9zYdp7DNl4BDam
+VzUdjbelw3CAIsomUL+kxv3UgBajIYYFOxvIv+q3ap6IokIbSYFPn8aN/tRoERgadmCdupoUVgU
3OTc0Q8gRGMoGZMUjzvF5Bq24dY3cy5XBdiEVGnO7+lFrxpGMko/qohf4mMaxTV8Mg8SBLJ7b4Yn
s850Fn/LdBvXeJBh82qluql7hsjKt70/jnyVFukalkNjLpyjPPztFf8T8Q7Kf6F2eLu7XTdAIBOL
I/qXLaXcgjlhhMTU8naZofnJ3MnR//wvg8L6ogBPk83CoKrpasgXa7BtIabbSXHWC9s9B0Bf2lRt
8edIsrO3/Op8BSDltFWXInt3gGG8wmBC72GGQATpm3uRDIX/pgF1cyrA2jIYMIMWjjfWeHFyjZrk
mXuQXdMjoBBpHaS2LjDU94nEoRFR0Ro6LAoLf8xu7mxCMS23IQJ91X5MQ3oYJQBe394jBPux1wMn
6ficLsV5hwiJQFctzhuHPqCwZmaiGpiYupSzXL+5WSgOFm7ylnBHom7GiOVQ9JHEQxNXRUYmyMdU
jRyWOt/B0EYf9DE63T7mxXi/jwg+EjymKz4nDPdMVLDqfH8fsfCR1+ixebTA0ZJa/awLZTjDt5La
sis2wQyHIcQUml968L5saDrtmT+C3kWUNV/78WYoiFdDqhn4Iwa5uB6LEcUpKPt4chYcrwIsJLWJ
rvX9n406BktiiLXUkig2l5kqHNLqWTkBLxJM2qQAOblUIqP+3JQUOghFqNsSbEGFW4RirKhEVxUX
8c//HvdBOBok9AL2BI+FZ3/SOTZDO5w6L2JadSpGr199Hs1xc9aEB+C+8gM+lJpHe2Y52YJ6tC2D
WDEBRen2Z5l3ENwFn6dOpSN6wK1VS79wIkDKiZt5Nj9PcPksM5NtlgDGrH8GxjrSfOBjybzKAEef
VJaYzxcC2i3cD7/84E9Yih4WYZC8W5enTRtycSg/zmlBiSmcHrBMLjrb03WsU5jAfqv6/SjRfwHQ
KJgLpWzYh0tfr7KqsFMDJiKCbCGskPAcXMUOU4if/sKjSlk6sADBmwTbszJGjct3aFt0cp4mb49Z
vLv0YPWOiJhTgcuL7MIJ98iu/EXR6O8IWpFemUFCz5muvsf/SwXKvPOc6aFFg27vS6LJB8rPqKTF
tvEvTMMv0mCCsab1H16YFT8EEn1zS/mW3VQcfKffHHd6qf8UaXLl+dpNIoSsiM0zHZfjosgyDcwr
q0TDQsiiXw47jUE7IAred92E5xt9QtEytPKBgM+VUgiU5IODHA1ybowbDhPrMgHYFAGBaoT+XaVp
IucLCvAsMxs+J6ex0ylhJRdggiHiRq2+VIThm/VoKu1j1W/HkSAkZTVeLodOuJOfsGuz+qUmjHQN
QhpTCOv+n6iV8zFbzKVUwqqW/cw3AvI1UWaAdOwS31gzypCuqmlQgMgJSMMh3wVZmM2OxBEvJEW3
7vjCYdxIgC6MEIMElyh7WOCObG6hVQW4EEukkvyD+bUgbJ42vGWzY/QsJngRizRbZ+EWxURUTWKA
JSLHUyB5LKVNRG0fUDgdtoSA+1DExzN1E8fgwRVk4d+3iP+umw7Q47wqxovYfmYIXlr2Qcl14Gy9
GmHggfbzc8WzGc3GZdAbGExroDzg3Uv0SEjBZ2osSQbotWeIEp2HGnNMOErc7xbuUl6xcmHhgygu
1bw6zbqBPIqCfJT61psbLn9PwG87LZQd3qA2fuh3G40kb49WU9bepxPyGCvregNETiLuP4OhHEyy
Ut73cYLrRMb2gOHWJRqs1zis1iam92sUcEw9xG21hyqz8x+SzIKA4Tq261vZA2zV+071bu9ZORoH
OzdAVeZLUL3/tEoqbnblngFcFAes8X051G3YaoDjiBNP/Rj6NdKHTmLzd/DWsK02jlkp3brmESi7
F3hzzaI+o7wjjrtEpbOL+thEX+SiExoGzlTM0HGLLJ2h3BCnwQbjaK4BdAuRPZRon+rn0vBxQirY
irZAZV+sp3eLXXnDBCxxSxamcwNY2ELsIh8USdQfmenRH5PqtdyBe7YmNrrHIF9qGLDWUyLxuoqF
eohPyQ4JW5ADtg0crDA2cqRrqMwEyNvNtkIBtLBMoSMVW8qb0b3uw/aAmnVgTSPxpAgo7JTgYJKc
uDba+tIGrXJasHlXzqJg99ey4nz2DldLgfpSE30qWavGP5dqkEuKB3ECEsUjphOOWFIK9nEBtRLr
VK5VaGTxbTJ20y5Wu1+GQTpHx98l4q/95G8yr9+w3TRTXz0uo2pC7ZjqeNQTx62w17/NMl6GwKfG
M7jv4XNxko9jYimN3sWlkk7zjjQUtlUeVtyJAGIy4qTSSlo6Psd4qIHsIlJSghuhgX7HfTvzxjrV
7i+Awo/3D8rhU9iWXLHT3UuPcZL1V6CKkEe/EI8MTTxdZdzocQTEg9+i6bX3hdSAGll/QC+dmczm
y/kFsc2x/agfgQO3FVf3v7bpr5ZxM8WCo0aTCKNVZs+6gCHUpQLGCn3orX9huai+ndr2KDuUhcMC
dJzqeCPL5hvzpR5LYJWT0EEejr2T2nbbB8PijiwIiBcotWftCuBuiBsgpLZGiaHICp9tnHP9kiAW
eLsm0+CRINg99BkixUs2VmD34VSSdeFc+4mXOH3hAhsTZUK/Q02QcfCEJLvvY9HAc87TdkSAFl8F
oDyqL1N2qR91On2kmADMloJRADsG9UGHs4neliF6C5y11yW1ziKURP3KjwfnGHCpcyoAscK8uyhP
xhI6I0HLlB79w+rLNLD45hThmcrtOF3QzRCexMBSBkpvqEHLWcYmmRzko0EJFew6dSCsuo5ZGVX1
45J+NgLzxJVjPy1KNJhF/nLEj6OPlnkdw8dIqwe3WBanAzMyCHpTrPgqw6zQrxf9wZFQy7OWsDcA
CqOHVAAUsT9pAhL7ubFvRQrYmLt2gyn1gnFqQCLfzFj9QJiGC50cQa1dDECgmEi/Tn1fODo4X4tg
bTc/I36WJ4DXRGLphZDMpRDMp1Hh8HALkZ0yVe2k9+yjFsJeyhrEHl3FKTPnGX6v6nRsOJESj/L0
wdPjGki7QrmgTue/cv+qELnZMNNcRnDt6ZirJVDZoigNk7dz/12mvkjvw+WVqoyButbGgYVzDEIr
uvWfhuO9kkAfoT86GM0MPU2bPC1M17v5fVT3Cfogwd6g/5QSLUFBXL829CCEOtjNI6Jq1wIObpZZ
v3cLS9rSgmDlpeYXr3cVWyn3MbjSFi/jUsfw7pcL1EmDxxJ37kFBgwE4ApPTeszye6CkEF/kd02S
2tEL4l1umVeAoArG0ukdeyaugQ+YAcvuNJ/ke//+JSOOZqNVYUM4Yr6TFaCJaP2iIlfbsRcedlK+
pH9/y39yAcncgKbcjfDs+keJEXVpPfTi++zHme3ikQ6y+qUpDDlndXBPgweYYrr0jybojVTYqyhi
W4GKbGtQIe09cBv13NUIU5ItsN0RMtnmbVTBwcfn0XpNcag+LqMccSre0ngrVMH9IArcKIJDUKD2
9G/OXAD2AFDvZoWBJ0Phj8uiNwOJvN/Ezr46jsl8uOtTlIUT26nWtTqsvFX5y8WMF6SXsn92t6xC
ymzlbticDpqWz6CoxUNpwc9WOuU/lGLmFVZJSuo8SkuVUTQBnTIdJSdlJjUxF2e3FRh3HSqpUGVD
FTDZkQSpE9uYjvfrndVkWCALFr3hErJDnbVe9h8FZ1ly/YNUzWFTaOfzLV69HHVL0eQS0d3C3J1w
i8wJUhWhT9XLPgy+eM341vC8hojObW0/sIcLyoL/Ai9jj8EbGvNIHi/iJycnMt7eH9WJw3w7mX6M
tUpRroNE8cunFVEL/DlGIYBoeJc9PPIG6lomV4kk7J7ibsGdpCL897CghREBjaQRn0dsXM1zyBma
fPCgGbyN7tuhAidO/9Xl2/S+AtCPfzsZ332OwccmNAU5/FS1YyHRB9pSU30ct1TFe8YwP2CbI5ge
pn8zxmrUe4c41wmM17X2A0OeZuJ422wetNLm2LyzU/LMkJFSg9iMnLNeCO9NtUlY7qw7VGlbYcV/
pDYznQyajf+KAKg7jrK2wWuSVsxhvIJfpV9iq+OU0qwBxFun/jfKchuCEzgesY4L3unkpgI7nNFz
S18MwTMp95IJTMTRYqUgV0JHmLoVzGMzpT9Ai1/Klf756s7xAje4xT1azBJnd+t7xxstGpzqisvY
MqqcuPsI9Y+HWM0Q/S9tyWhzdEWb511Jpk6Z8ZiWoo5TYsxrTERgJBI3GG6Jpq2bUgZEUCU7FyeP
obDfzdbkZ21Q+KLzpH4As93FV3K9QKelKxVY+/MS6yjjJ83tp1VgkwID+vPcinkitzinoTQxazGs
jBJ78S5oqPKKQRP3P1mAGOVpoJTUpqRrAzai169hU57sEg3ahsT4sKPKAzGDTgAVIGxpPvS99IS1
8KMSuhFxAapoJ0Yf5Uk5zFWau/E/Xsj1Qqmzl+7NFdlC7y2HGEU7HqxkLkzJdZGzpQI37/7IDxFB
dt6tHh8gcrjUkF5GvdaNNl77O32ba/CXOwOcWa7fHk+8dPAudpe0AEm6omgAttUJvH9v/ciIOhBI
nrHzV+YBpifC2P1Y6ORG4RS3z3UsXBjHH/1Fe4c8B4s9mbs01mIKocAmhOKVuJOWshnNrZFCt31I
/5SREE4hPwKwYiwuvfu0QBiWw863CZCWkYwgDgHgSzKNm6Y27c4qyFyZyEKe5zDYFzHkXIfbqrpw
8cuAZEonFbi4wlnWFsGnYCitnPEf0ux2dCz0zmXHlqjettqSNqrUezfs1csfSKECoF+XjPu/Y2f5
FSMjXcVOZi8lA4dUNXa7pthaYKhQRwq32DWaUqhtDyZ/OUHcvaTd0cKJgbRqRRNOiIhZf203ZwO/
sUQfcOzzY10begvwip7GBqFlRcVpe78QPbFVVWEVsdl9jjozp9ZALd8HqZnKLDlaM8Pimiy4lJAQ
HKhIH6RylQ44xGfCQQT3WUthZinxRa8KjKbPKC07NIFws/Q7H/EUK/BUO1V0xJOrDViS2n3oo+km
FaeE7YrZEWrIp/8EL7fKGGDN26mUa7E9HXGg6bgnnfh1khgKDvYr+xNi74Gzoruf/Ce31NGpncBT
qmi+5JUmp7D5JWp4c8Lh82aygV6lz/PjySUPtCQJARo+OasIshYw39hy+i7wgdREKpuPDke5ysv0
3aMx9DlRCmyNV8hiL4/fm/74ONJPQcAjv5Z4iN+2AQW/7GZ5Q4X56b5y7mKTQikQKh9NJSO+Cl4j
ePZocmZ5YkYt6fY9zgVe060nsjjM0d2bDcDjPcBojAjjLD/1AGRgmisKy5VZY6wAZvyGmQyyEh3i
3KHvNK555aiHoGzg1G49JOm6r+SUhdMHYizOrbua+3rt0h9jRT0anywg7xRWD3CYgJXusF0u4O5O
WEQh5wVvNQ87q8JYBuq1uq7zEbXKOed3jQHMmi+sOAqkeh2PUyXE7EzGsPSliS4hWsyblDWWg+Xs
Mzs+7DXskkMw+gSEZzbZqsH3pR09KRoOw1JLcoO7y0LzHb0tYNMBLV0tIbyEsMiajVbISP7dIoSW
mKtyP/yYsxvEQvjXjfpe7HKfYzH0YKVK3snpdJ3Q7R6q697FPF5cOtm7oYnBlSlp72AcMLybZDWx
o2Bz0p/gBQA3hcRsJ2jjfkNxv1iJOPeboQcFp/Wx01JwLBFEO0tkT+l5SVTt9zZOlp1UW7Om5WGu
kY1jg/4wIyeF0F4GkBPy6XxOnKM40MiSpDAuAt5eisRcWwgbN0X8n/ezJJNgDw3t10OPANUIWxIZ
hURB+Jtc0gEqstVIiF7+3RfCGvz4+sSFUNUbEOTzLwPnzy1iWGSDG8oSpJWyIKTXQrjZFYSAT2vp
y3tGum8LoO90RYui36IPlUSWzr+82o7niMLMiiZw7dys6rtluSYJ7doDZrZ6M1ubFzrXrJyWJc2u
LERHWaK70vDFsxwJCOT+6R4+qVhfJKNfQPJ3YI0m2J4dxjbixwZmND13ILjsH0ZRAM1LHmBieo05
kQ+AN/WJss27JPnaZYGXg7vUb60qIunYkXoKlPCKQ/8YowLUaRvYNvYQ03wyEpz/DEwUZCOhW7w/
OlPEwzjF58OMOeedpsavk5dPo3dXZP1/hEYQy8IPRBsH30h+XkB4PEoymdenoJxb8+5R617lQtrB
ZptuheVGE2hDjG5H+zxxgSf9k2IAxFV7bytgaagDwN5VxC5naAT1r4dAuxm+AuOMsTQvmbt7ONYv
yf1ubIEHCSlh2o/9l/chI4co+7NUHEgpI1L7uzjsvTj8c1zgGP+5Vn7uuMeCBIBYQ8zVm+ZFxaTy
FUoCYH7Iy7UE2QjFxSahJiJHLwHRehdgQClgAKnKlsAmyLQF5c70mYEdwA3x+02C/tI5/M66ZgYS
9bTvqGnII0OtkJmns++efNn2SrTahqZoT27ph1JAZ29WpC9YfJbNRmTrVIBYb6pGx5GS/E/Sf0vY
hM80xhd0/XXUSqDxACBXjBwAtEtOguiX7RgLnbnRmQNPi0El/nGRQ/IKHovQD4LC7P8m6Wb8Trem
3WuyERy4oGp16CO0mQZyx/Hd4+MTO+fb3pd2oDJOjAI/Z7wW4CpHFFfjzpOWRH7OOjywJCa5G04v
OpBaB2nGN+cnYZtislx3L3g7o4tHhQHZOAo0awkQjL96SDZ9BOelaevmW1Qyn+pWzp4u70u81OXU
1Wo/kgzUe0bywJHp8o3669kPVS3R5U2hGFoBZlml1jAB988YDqd51NvWfPwS1Z+A98cxkMJFvLvp
Ds/ZLh6GHDOd1Ac/x119SKyfpyX6cPYH3tNzDYkndfLG78QFNlYpO27HkNw5OMa9z/2E3ZyCQdcU
3x60nt8pYSoLcLOq4A6mjZS6By0UD0X+G2Iof79CDwrA38zsuKgUrwITxeQkAeH3uJSntihe7U0M
hH1qp4CY7cIbAiFR6lnk0pNF2KPkNlzTAyD40/VjfVNNfcnvsA1JQ7GtEClr0QdvKyLKPHgf+E4G
W7rwmcCrlzQVNZ1VIkE45yc6pLwuPHw9Co96txhWijMO9P3BUYDLGDpU81vtJvuG8ff1VnD/8/J5
byeM0kPUrFQpJd5JUK2ItzaMLBnGT390ypJ1WKHMfVKe8pbCwh0I+AcxHyMkS1AYfOU3M1u6X/N1
CxEUJfGevTgIH/wzK03+FqdOPvqqe8lY0LtY2rR9lz3R9psCnYZV1UhTfx4eFevwswzICQgbnEyG
jFk4Qgk4CRmVEgtJanJ+ibkM0YGImtqUtjIrK/FN5QRpw7hKUnb+SjTsSB17/j+FtLvnTlr605FE
rHWuJImJEpr5ZgEtmSmtQA8YVHbtcJeExxMK2NTDC+X2VMYmKoMvdTJ5SxqpvAXgkIFSzm5EuyXi
glWV6soku3gysTEstWRR6z5vGK7SwuFs3MaFVgax0PydIoQlPAiyB2j7KRTSwtsTCI4ct+S3YcCl
2Bgfqk+NQKBH9zmNlTW4Qs/yDAyF/1GpaXIi8HCeFHXD34DNC58Nfr/11aiavDhB8datkMVgrOti
BeRE5msij4ipHZFRrDqXqN1pJe3E8mw8/dtcCVnjwnuhs26qMbfSwBKqOrhErKxGT8MGZUvxihrJ
CxE5NcSVMnzPsCKUI0GQ/CkEMny0PCm6/IUT6niT/vse5qoaJO9NosmqK81iCtuPgwm0mCnsqkir
RITkYjXxUtJcKd2TpsWPkSWxkGhPg4+daqv0P5bO2O082HvdzXh75cr1EY4JipUE0c9JWKcNRdaM
eBuhut0bQvnqI8oV34sVGB+s7HkKDUCGyBRPaGhm2HnPdgzFReWTranB4mgO9s/BlyaZn8bPHdRA
T7L+PWCBQDY2jiNYSmU7EpLOxcThjWAX4ihWcowruQrUL4GTBKBMjIucqe7zxa56MXhCYpzwtVyW
4zMW+tZTiJGxME8fX/hE1rzEDkPk0+kZ27Ib7p1d3X0rbPcyxgWi8WYmyCFl4pbWb8LBYtksWxQu
AkoaD5D74Lsto/eELiWeN8f7JmQfNwhRe1/ZRV1TE2Bc6Hz36xTIYboivgjNKa/taeJhzTQq16H4
J4yNew2plQtoqYq9c5SmlYM2A9CU5wazYC29DWR6p2zqKvX08HRzWokiNNktOdvelUEQWNyDSrHF
xZXfuCKihM/uf8UNbMTeSQPE8a0aG6fj6zgK+wpErMo79uRDZgxBvQh/9Y6//wOjZcYH13jzprxM
v1x8jgUyT5GB1YFoeA/XOUIbq2fnLS+DXlzYoxSOyEIQDa7czCMqWNO3Ry9lUdZKZ0cyaMIG8jSK
nQj4t0vwErxdut0W4xfGAQRmGJ0sDitceNYSIXtk5O3A2BrpFby4kYK4lA2Z4yEPg3n2lGjzWdgd
KnhO2yTNgL1gp1aabsbQ4FiAQmPxofAA5V37rKgOLidmW4ZSnzhVodcAjaJKyTGHf2gkEV8+d62P
2oEJwT3/FfiQn0Ft88gMctjIpVbYEYtTzof+fJGbijHjF6TkMrXxgvPzjQh7pisTQMKE4kHpe3wV
oRAwIokzT0Z7lB1hPm/WnHtNHXi8omEYlBvEfxz+pxcPNVPcmN92GGYoLKBe44+MHKw0grUjRFil
kIaX/1OUMnJmDm9cc/Wfw6FdtTEg1bv69yaQAR/LuKSsvoTBn/vDk4VQ6AQROoVgtSWrSMQsPw8z
K/bNxrfmR3ZsdEFCuQ6zQDKqYIcq7cYSaa9fuW1bxfQeQArMmMK/faaw9jnqLHwN0JJJW2f2AC1N
+PVDmDlH14eBCmAnATcxB3R5vbHfFJYIfvaRMzYXxV5Y6PwvMVxPKxedm+FefNUoXgkC925drF2+
irg3alwiSoI02zLd4fOOHfJ1xmixO5y/jZXMVzfRGbayH5xbPyGC/XsKX3q9OgDJCo0pMs5mbg3G
/gyQfrxg4X9zbDQ/d6dM2AgmWZShSkQJ7VpD3lC+vMTPozSBRYhVjlmNyeLgnVBTsKbVnt93hkho
E6b/j/tcMvfBI4B3Os3k9Tl70JccGx5BqQYrf9mblFAS7eQ/yxN4vNHXVCCTphupyHpwGKguOemz
eDUS+bLskF6/JPKdkzVufpsgfQ58E1UcaoSSlk7cbYhIcbml1DSt7ZDOpN1iFLyNckdd3Zw8S5S1
aOZ2Zj2lCtapj47JSb+Cmrz6ztwm8T70e7MaNLPOkm3eGH0OCGqoGEyZbEYBO3XSgmg61dincpHd
52vljqOIEmxMe/BI6hkYsfRT1tGJ8B3lV6b/gh0FX8FmuZE6uwJQgcb1YDLm+JcHVTSCAeBWifig
Co4uRbYsE/xBmQxh8ZwTkeN7t/UIO2ZMJKzNuh9Rz2LGNyvowMIX9iGLsm93oHeGKRaIX6T1K3F7
6us4Wbtu9uSDIS8WJkACykSEICVULov3RTaXh0/i8IiqKp6L44d8/5ziKbRm/gHQ+MIQxD/bywIu
RV2uiT8hsVJCrfMlGYcrbQ7CpEaQHtUzcUppcVVxMR5I/lvXDDe0paRnzdUbgLnJNLhLFU8TjnHW
ubCBFkrPIgf06aS0xLzUksSzNyQpCm+QzwHNt4Q6P4pRlT1jrU/wKg+szt7uUKcmKFtZw1+gvibJ
aV2EdGe9j71UzrYQJz5S2HYEcgfGqdtbksVt9bfbLeeNxTThOuDl7hPMsHLACAf7ZU1HFi7pedVD
KGjkwX1fL1iF0uA2AYz9jdjiP7+C/uiEr8V48+mgvgpCYytNxXoL/RXX/sL9yq6jzWO4Fr031Kjm
426N+SeSQY21chQklGLWDLeeeyqJB4eTJO4JhzuOlbFAuibR4HHBU73mqzmdqC6JIM2GGcgQBGGL
HJJBfwfT4iYLf3o/MYMbNv+keX9LKTCARMkifuc7Drn7UazO9gBhF/qOm6bKVrkGCLtAtBU9NC1H
sHzWpl0b6EfKBMpYhRQD5XqVjRmdopxHy6X4hEvBkXyQJnsN2hlYx+cZnUIXWashdYgY5d/URuvQ
dezpdTwLa3i+FsCzAfIZgjR5aajhVXFNWCHpZmk0aFdG9NlJf157NzXvaa1clkgaA+SOjerT1Kts
iGSvseSF2TpjOyUUgo0+N5gI4ivjOa6mXPM69wf9RjBWNbl63zQy4Ytijyw+Gee1yh7Yhdr6NzQ/
ThzYYyclKnngDts2lMeeg3YTAAoDfl6WKTxiKynuKqvP31s/J07/XXFaUUvur9gyXflxemS5zciR
srbLNJQbbxa0HoNlI1JN66N7GfVdwkI2KtcvXLUDxudHyOQZTj+E5qri8KGp8zq6aVrpYXi/hI4Z
/Jb5c/tK45mrHMk9w0XYodBli+SkF0TO4krbK9QNyLQnxdwgH68Pce808xKTwZ2hIt76kFbMkXSZ
zcl0py8w4SNfFUhpo2XNHwvMa87bf09spCpHPUa4kZQ1X5+DWFhRus9QwkcDyVhjz69nINABBclM
fg/xPpqR3P+4x5os2ls2OIrnJd0WPKO/1mghs3+HzzvNNbXcehKW29W9cSjLxy1fSb/R2JKpjOJz
APLlAui05jUk8at8rEvHnkxRzZ3MNcYA8MaRsZfPTl+zoqeX/QMh9CXxqD8sDW8flYIR9DPGs5C5
UgiVN55La4ce2zm16vX+lKkbfEfdckK2xSThGN3Yj3L9tFjuvfYGTckSyxxKEyzTqE0gUl92GiKb
ZZmR+o8o7jnXNf02AnOJoyEMp03AwNqlzEpiR64zX/l3V7fkWbEY1B64o3hWN44lANmWmRJmEFrS
8lyHwwf/uK0Oxzgkl6UldFK5qTJGnlPn3BjHvJemO1fkcFwXqK+qngTehcFqVB7gkqshuYK88Dzs
ttgiLDH/gwpiqtzc8VA0pxIOTWmuYwoGPqVvgtnh0KsAh1RXFhtILcuFlumeDvjHuorkcQLlWA5S
ex/7NXm1zmD7hLcLOA5cz4AkZ+cYwtTXCQF/HsiAtgn8/bquKUPddcAvx7vQGymrcsfB+imxIkgF
6o2OlDRggVRlARW0m8dKUYGjaIXiOHhFwi2urZXny70lLBjYzD8aXz0XcwOPvJrJwFk+fvZyOJFf
ZqfOqoEV1tjJi7cndDmVcRVSIpQjyvUFoM+L579a7vgkSOWQGlOJwRBGOvD+weJlRDhS0CnABVdO
6b4gS4kQrjlj3YVhsoGiatOj4w7v24sL9c7QnAcBuzYHj0bHGbzEChOXvVHeUnyoNmCzQ6BbSJIi
Uw6AuwcyxO6v4w6C+e6kbefP/iKnwbbq+gJ1qDsGdcfK882wDbgCYsK5PusJi6VH0htZfH+I7pb7
bbDwclUuSM/UmSAiw3UL3kAdjHn3DWz5U0Eslb7zLelj7lcKddRrIUvnuSkpN5hp1PG9V7l1mCy2
6/K23YvemJibaYceIGTmd61GdTUhNldbXK9FwlTltbV6mxdwjTh95bpHDZXDLge/qPBudV1+DjD8
cQhmr0cNhj2+SUZfntdAi2kEdEywR1IGqGJHqV4HAxQHMv/qGK68lObl2geeU0kRyRFATe7dZLCS
EHxCSQBEH+SH6HvukFIzhbS+1XHJvvee9iUmedEEXbyeCi0qxkVvBxLL8vM0MHOAOhZO0laOPwAQ
92BJHyAsa6Wqzd9Fuskd/IC72xRpmGoBGMbld/wxbExpwyDiVSjB3QshLkdHS7J0n4LOrvcJBqAn
Hj88fW2YIrf97+ZkahiCdDb8eIiy5m0oOxhUlinA9lzHf47unINXUtwvYaywf3ts7PtZ6iPyVJ4g
YAHIU7jPBE4KcmDfnDQYghf8kBzr2vPE6m83eKjD68AHYrV60Ee6cc2P5mJaH+6ng2eSOToLc1H5
nHLmi/SliXRIz0tQqgbBIcUmJgIM1JYDmCye/e6zuRZDNvWfRpdY/EKvsJcBKCWIU7mJhxJbClOz
B12mZEy84caK34onxUvfdU3xpE6S6UGHqLzlJDRBlruwToqueFEGw1GYi0U6uST+y6bFibvEV9hE
1zjBx9uwMePy4Ru1b5gMbRcIhgOleXqaT3/5ANpzlaKheYHsU5C+LxKbfRrrsfMZl7f93ci6Azm/
b40UxHlWFUB3FCmhVQZIHfhKjLHo3/I8AZPsgTZlvm9GlkVPTDiVFmK/m1a2NLwEECSvMWkmzSn8
EqAQ36/XEnCcgibpufDaDE4tBw15ZPrPhe/xMwc2uY19TavTSRseVfJx78cBuMUGe67Dpp01xSue
rYuxPOHrw7dy8ugbTbsn5gu6qZ1GGEze0r6n0xydraySv7WW9mFZ4k3pOnHZw8u82IE0lu6uixbE
9ouiVP8jcdh/0JcGlYEDyUnHafdZ4Aykz2tEP9IBmQNQUPdehN4rMoHrKYH0sruFBmsW5uFPHded
AEZ3gXBEH0EULR8CHWHD1pT60Zu4u4YgMXz6wR51ApRk2WBxnnqt1xnNhlO5YRHhlBrHPO1svniI
nyy0NnhuQmLeFPzzWuEKSHqaPr2tQ2/HNrdGtr3PeQVD6rJDQ9Y2PBreBXAqJP8YVgbs2thf8Zv1
nIjvDznRwA4jc5bwesv8YTRT81EG4WLULEH0E3OwuCf5JANLB18HLcSmYpPBXFxKDxXaE3lyEfmr
cru6Fwz5YauQhJFfG1KlibjiPXjqy5B+mb4F4DrJ63k4o0+cBBRvN2p3scwDUm1cZ15A74mN6WKI
nN2nuT/rdUi7j/iqc7NBZr/6gjgxyRlXtro8WpkSLlP6Xo11LovJIuxvUjlXbeHDmTbCr+I8JywA
kI9FZMAc8CDK6M10OLLUCedMWdzOg0hFhFJ33XC4kNFFZ+8cZvJiiXuGmrxgmXWFeB4xLoyLWSnX
NVEOUJH6gkqiViHgcOGQV67Ux5haz7PZb/VezvcHdXHdcR9qQ9BDTPPnFZsuxup47P+EFJAu3dfv
A/nevQd+2n03eGiV+XKSO2vcCfXyQi2S5mZ91c69Y4cDDMdJjsfJjzu8DbRIRt084kJlt1RLtrmC
ECsCyCTV8/BcFJRJZQWYy4s/i43a5Vx1qtNXHNqzXn1dzy5qPW4oOtBqU2UbGk/2T4Wo5mTqZBi/
tpf3S6L8OdJK2cK4bxYNwLaTvOVa+myDT/z3x9ayRJPLQZwGyNGwNagTVVI9fkZNYVzV86Zy3auZ
gFcr3wWFMpp+Z5jgwupOShz4MFnuUHSWJESieOIjd1fsOO32AU1ykZnbH/2cOiwEkmSqBO4kuxOY
mDiXk/0KGiw/FK/xsM9btJCanPrLWnYmqvZAMY+tGksmjMbA3rKKa5fIseB2Re9gCIxtVCjMnC0W
YQHuwZ7/7O3n6xpMDwxm6x2LSRf9mzkLeT69NAhRd7iJtLBdWHd62iED9NbrdsC/erkKmGXxqAks
ERUhp1UC0h4Y6g3nlj2Xd8819UwYsTj1T6asK9feBB1FXvbVwDJ4UWdgNKOVde2CmPDbL1CwUBK8
TPByM+zt5Azes0R0n6lr19UTnaXMPvaWMAisF3wY5cH9ykFjIwq3/1Wj+P4s3UIEq7ceneCokvEn
Q2EkitSEwbk6JLTSjrzE1TLPvsAvwcK5WyFyomIjZdCmILFKja5LMtlA7aUG4lSMLtTOXPxOGc0Y
NJIQhR93fDlaRFCTpDNT/eVL/h4sBiAD+zqreUIqD2SgQJsMuN1S4CciZxnldFc7Vu9dPbWyxt5x
vnsWZs8dfPjCtm562iNm0Volzh5EI6IM8JepV5plek/3c+a7si0A/Fd7eehyXU0onlMt8CJNYRrt
qFmJp0hOiMuurnnd1RVeDYWIGrSMpRQiea6LQ7zNlm13jxka0WeM3VWytjLL8F3kYXWz8xSuGpRv
LY2sHTrz845UV0R4mKanx1kHFDijOuh4uvjQ6rEjKKrkQpfc5biXl5JyHdLU1IMpR+qh4H/ec7c+
ByK4iHjPtxjpAzajpsEmtKpP/W8Bu0/ZlrG3uRI/lhWa1uEtA7ao38JuEF2Yfix6dQSM+sU4QeEa
qosq8XsM10WtiIG3+a5LaeexE7pRatGCOTGTRKFvXmuaQZ0XnQQC/DlFhEgmYbud3HWsyovUuAKa
g/6ddzHKRbLRbx7Kg6aVHBZEghDY4LnDDavR0MEVnH27TR488hYBLDDmLwYND069/N9Nq9Fd6OGc
1tpmF8GqvDdoeAHPKF2kzCRZdWGQKUJYqOm4csEMI8sgJlY9ucK7YH05sf/nFlt6xRTI2ICmBcw5
DT0q3YFuAiEiGjBJSLAY5xLug8rn7v06J4KdLTotaF6MVdWgeBo4huLNd2hTF5CJlS6R+oRoX6lV
I9YzVQF04dGjlAys8OaxQ/bAl2p0DdFWO/ZsOCR0DUi/TwHVScQ+4IzFAFkBkDgvuE6oA9XfZE0g
/dJJR3BEsPNN6C4+RY7JUzR8rKcjHws4bsNISIMihfxC9Wjo+86boOogs7R12UiJY9ZsPUSGYKOu
yT2mKLqLqMs7g+Uu5ftANnVyfOHdsWnj6Z115gXWXJ6nNyv6zIZvzFSOKC1dQRYCjXXTSUK44Jyl
2YpH8alTvCRCD+JK1czrQegJAbLfXaxoF29bzpS6Qa9nw/fOW8niHnybL7OK62ko0K1XsndcqHJ8
0EU7MyyhoJronGEEaXoysQVnld+qe6SG01P4DN/GeHjtuumLbBiuycmLPcw6n+rXBq42ErvKXVu0
atYu9BQCeNiYDf5YizAIFZXFhAcMzzUtqxMTqv3ZawR8y+6nxf5y7xs3CbJwRvwksZte7hZSrL7D
tDoqProaqcmZV/0uPuH+Le+ODi0z/tDYXReT1peFoNK1h6HKfsJUFm9DLsCmo/J8WeAINPQOg1iy
D2te/hyO/+5mj4Otk+fT3dql2ifQik/Cws64qAQPRT7aiIoTskIstxsVpOo4SSfgz6YiVXDaKNG1
Ld5LlywKooDA8mM6xU3smk83w8+Tcf/tezT+JhLyPQkodOQZhL2FYGwk7R00KbXDAJEFBpvFh9P0
2k2vXJ46WvrSFz2gNsVtMm8bAD/FUgOvdCbR/Y1+nX778c0B2oycmg7J7mIqsXmQRx00OUVQOrPc
yQJVnFTypDs56DgJvYcwG/1V3UHSJxzEt1P0KRSFVBixO+kzwCnJ6/zlZhz8W5ghNm0VhBMNh+1Z
kSW14MwbfFGBiG97bKWX9G2DhctWJ7LYh//h2PZAIBjrNSpfe3lTTdHfl6gzGs6JmF+H3VkJ+VeQ
dXZ0fGCD4fPScRmKgQfztoNhrgGOe9bajgtj3bUxHBtWauH96sQCGpsR0VODjdezAxizGe758cXS
7LIVo9W5qfxfQ7gbCVrPRX3fjL1boa+mL0gzjL23GefuO6oQpLXeGmauTpkY65v+5SOCL/KiKPvB
gKtX7aukN6F8irR2DPnq/9x6FMIYcEgAuXHFNbhhR9HTiKBBt5TRyCd7oyXpR/kqnCnifnuIPJEm
EIfTP2d7wt2mlSq9kpzcUjUlMIH9pdZaLITbaRcZBBnFD/FZvV28Qxhb4ZccmMXo7QXoph3+C9aB
2leXsMf4jeP3HwEzHizWHln6/yVuPBnbNcYKjW9UuI8vfLOP9KqjSlTuLhlL3Xgi2fFm6NzUh1Wf
UR5w3l4F0ZPVEHU9VCyM+NPKjMTaEnqEtP4b8uGBjnc5bbRmxeU8Ihxr6/0f4Wh1Mv2VVCRZMN/Z
ta5nex2244HEEq6XoIxnTju6jWbDReVaG0Y96dSAxPLPLqPqtjtv3qTRi7G+3MDbEy9RKRTpfUg2
ysNB1gPWR5nuQqZgDjKeaCw5OnwIvXq3wWsLQLFOrzhru+tPvLr+lfHKcXAT9YnmzRDJnjigDssU
56F4sLKU39ZZWQM2H/xl+z+H1OGqgsjtgSoPyYp3b18IRb4vMlDLWBUowLQpWM5C+qW1KEDrlFqP
u9FjVuRjcQ76WqZbj2e1Bu3GbnrKHFZ4ADnClhgPqhFmco/tAReF3mHqAghY+eDrgo+YvxaDPisX
k5nYGG135VjqIHeKi1W6Aj8WlDzkrLBzt2lWWkI5qAR/TlhaPzkEMVaYLqYjK8yj3qiDpJaMyLBu
JqG4JeM3++WdXQU0qd+0IcWpVaVg+tyexl8XYmjRNWf1EeuT3x1sP4sfzCfBLPvV+0LZjIgjyqYm
trokiW58HRoorJPZrH9aHX8Ov2FMNGGAj5eVizEpRTWHT1EoMPOYV804wl5veXV/gR4U94VfIYMH
yYh0LZkYXXt3ckgUuFILuhKMj9tNV/uMsxlOwaa0WrSGUS3NxJdB2pXpRheEUfvzxuYj0zZ+iDAA
06wBDamHM3uHCWcN42XXXKa0rnGoANhevPUVGG5H3iwnt82AE01uF9LsToBi2pv0LY8My3h2qFLa
VfeOwVIvLe0tg+ivRKonpKo79U+2TonV/nOLffWkOXMQGgwQh78OrnIvbnOrh1P3KGyAc4DVs/L7
7MZxXGP9TKeFjnjCBgMCWkqXIP4n26sJg0OH7q1zWJcWdjZclRcHiTfZyHOYlcaK6xwmby9pn99Q
2dUI+fMKrvUSnMZ+HnJcA7rs9pV1DSoZmRJuyJMUYoM8Dbp4cWtSfkeN4SX9BPosSZpyuhZD/Kt1
GXFejT9FcE1znsSGULFKARfNvpBwkqbW7VRS3oVmhwKC5M+wqYKT7kWCoDXUYCASV5oHMqwVe2eo
1aX8TldoU3U1x5WjRmRquOEegz68Gih1ZtzTibrWkvcvuNPebRWMKc2m7c1xIB5n8h85sTI4MnPW
GyApAE8jqqXCcixfizKNNXRN7QotgtptGCu0DVZw+8scT4iOd8YWCelWSfPRLjLJTglP2XM3b4NN
pYrv2IHIiVTOlDbc8QjW+RHR5t3er6DVTfXaHMIRBEVdChHL9Q9J2YqH/2CV4mxe+EeiT+bfXwPv
rehCbLgmdJ3X1v18Jn20O0NzfaLjjS3qAnKTly2iyG1MmF9g6hyD22oNXHrCyZinxfxGYSHhYKcB
TysiBfSVp+KBw3MDXnstSsdYOmCK7NHPauKFWyMadbS71S7O8jzZSCNWW8t8gSpSwsglnA1P5DST
KZPF3NrB80L9HbS2/+fR0zHtvHa+PnjPnshWkyFgfPGUO4G8fNsv/XQ4cfaggGOLWZTc/j4To5+k
ZMx26qTh+parp+UHrkDH83RZz2kEBvd8RSEJVa/CmgVsEDUc3IL2syYIIfENEmA260L7e+QRYMEA
L2Qbqv3p6ZBgE/VSW5n87kc68Kk/xqLvwpuN04W4VbpDUwrsK02qWzQ0ebkfk/PDjrUnBcovsPYH
nvrvu/D47FWqk4tBbOpcRkCqgL/QU9SMrJkFz3r6iCyqOhpJJ90mjo2EPwjj+7L90zsRylTJvAlg
oGxxIMHybaGYrBmoAzMAbN1AtpF76xZDc+/NZLBtORDZWC5bLfVfpmptVj41+iKNw/URc03vCVq4
xukpyqB+MnCeP87bE+eStQnSxfh/nGnC5HB4hmQ/AdKqoTdtnHYYSvdGK+RVl4NKfDIm5W18junf
EUQvaQjTowwBbVbeguArRp81ObMaNcjV6Hb9u0ZGmLELqEEvH+bFct/UYd7Bxw/aYW1KFQasgT34
EkfhCNgdoginf74ehbsfHFTJ7bqlJVIpJ+N+UbkBT8kmndQ8BRiHYXOlL/gLfyXnGpA8zazHO6/C
wBpZzHs7s2lrvspdODl8ROsVP4oFPds0PhQ38VIfp3OOHkgMFMTONHShR/Y7QqyvfFJWdbqw2g88
f4kk7jtUS1+LFqLeCcuCaTMNCBfF1xiypCxCZN9lD1ZxcXwJY5JkL7dSdoMMaSJ7twMkk1nppXMU
QAHCMIXoQipXtbpYEnR/qaT+HgHlFPy2chTujquxTUhqY9s4/rZuWSBMdJYgysND3TQfnIlyyVP9
+PrSdQeQaGsueTnBc3h9qSXTdT9RT0FKmcxR+c0WE+QlMHSPYunZkiCvzZPMPN25nlZCFvjBr8GK
QX+tw4cq53kCxiKfHs6rTxhbwiY7dcq/r1GorrNeMBMC40nFA/y7tZXwYe+0roE+U9cOqEm3ym8e
oSzDA9MPvV/AJySD/cvngrIEfBc8ifPSK5Ak8E9Ky1uxPnKPumUkgPKurA95EznpOHhoxqA/ocHX
SWcq4Ng0fOdDFDIedJ2tHwV0J8/C0TqbRsTiPxFujntyIlsYi1cGvK8QfjRtK0ZdfopYFWI3s6c+
evTFnP1k27DwfbumD68l75lI7CKOmdGbMRBxt6EgV2P93WaDDigH7Z515CrX/nvI4rXAXy/Eggmz
lBqJlNXaxNSGcWdkjnnx838usWDiKSnhQz8p0HpEQbe1z/MTdGZtOgfvjZvDBpsovxsS4llyMVMw
QAOtC55y8MrrMPFbD6KHB1o5crJl0syWSylNy1VzYfgklNIobq6mEohTKZpdfcD2jkT/Uco1L47/
WiSqIRtv5MO9qNqdiYVSWyUvv9kIWWp9yk6g4zYG5q49VaxbEpmK+8l+999IRfOAsk8G7luxpzSa
m4OEcPDFobJrjUrm3eEssAwGlhQLR4PWEDnzyCmtbsRtULBGsGdZJvPCR0DVfjwYbtis4jSSi0NQ
zH78eml0nACqExDUEhmsQl1GxUZxoTxH1kRqrqbSrFfHDj89DzsgufywI/ZaYZzd1VJfNfMEQbMP
3ILsGOGzfLklk4JuPsV29PxLhagAX8hqWn2v+wTwhOQ19aG1fNyBdTeaEOpYjzJMwNjJO9dYsYJ3
YtoXpkDG61LuwtFS9nuAwiUoXEY96k2X6sTuGaPFi3rQu7y2BldIJv1rR35kFuQujyPGl6T9NPKB
xX4rN6f3PFmygOjDkKSaBeKNkvFb6Y0+UOMu+HWUQure0m7G1xIMscG1TgwYq5tAnHHpNnnIS1Pj
xgRhOB9+If476NWuDPjzWouTgfsdFQY+9asGquMXuKL21BlJ2ROR/8IMw8m0wbs5KX6bHFZY8JyC
3M0PyP8nDJkaqaxMDkKAukoHHZDHbOMZWcbxKCkeOFip0Hy94DVDR1pZJT511FWR/wce+ZXfLyE/
XGOdbfrb8gUqCH/gtnazk0DoCoPsU3QCsjQOSdjrovHz+rEUd4OmTNfbKgtNhu0sPvmyyOA5b4gC
NAaTgN1dBr63/lW+5ngXCQiNYQ064RiJOecPx5SOa63mcXDlcYG90fc0wH2FSILWE5FVhY25DNrF
9E/Xy76tXN4wjJf/hcriyO5gDvSMMtjLNXFi4qosxSi4JiF8NjCfRqWwPMFsNOIU3evui94b/9/h
yCXMNebTAD3hLCSx+oLAyXiHy3Uvdxwqc2iBfip+Thzq7/2zC7Q0ZdECGFAXvCac/xHbDK3Pam18
OzRrbH4/GpurSgcIxyi9r5NGnPSHeBrc2dEk3zYa3F6rKbCCXjt3IiFjw9HwEsQbc7I5SpfOQdH0
KHsSLGjZb2DIFrFVx//opiBjUdEFoJ5qBZVfqn+uVPcJu+GyyeI4jsAiwrjQgQEGAci2909iLCOj
B6dFJdighXKpnIyOQ1e7SPpfwReqzwoV9SXdbQYoSlxMMD+h1ltdYyH7W43JkczJBwjBjNJuv5gg
amWWrLkaboEQdMRONnlIZI+WTVJ3EhhgLFxJOy+XGe2m9YTXAMZtxyPadOqYJEwmvXEJEw9JK8HE
DV2sa1MvMdTihyp6YiXXOEB5UEgZSk7VtVRnJaKxw9gR1vvtPEOtkPXbZOi417FjYcsp+HI64aqK
+VvXESVXNyCUnHuhnL7WV6EkkYxOR0cFp4fc9kmFgpo3jPp3duSNM6zHN7GCjJFUgkb9HlQmvimi
MWKmL8hy6Bld3fbETnTbBoiDpWxsIwheFdwm18wirI/4R8f+tuD4GCey39WglPEFDz+OZSFrMCGp
NyGkX+HxX4EBsob0pusaxSemUBAWj6OCoYEoDiW/gKqYfjYsVIaN82crqQa693E1K7bDJp1sS5x0
X0qrqCd5F3OYrWizk4mq2WLMzLAz+V65uQHktqeg57EZkPFDuT+I0JcVq/xX1/qZxu42rX9Ud+XQ
J1alL9T2xNkFymSUfF8PnBMR4A06Ni8qH7+8TgeFCc91GI17FgErM8mOB3jiOwGWzSyYCO5Vd0JH
OoazAHwGkSt1S/6XEmKEDjCC50G70FkTwJgmBn/A/LI7epkOCd+Cnlwyw0h6tXZ/sMz6RxsvZ1/T
V8jEIxuD91wF3aXrj1fknDV/z5DOTUGavS41F6rN+59Mt+ZiCyp811rxXeLWAmpVJB2fENi02fbx
d9lg2x/9UQOsHvG2cBj2o4fxXCz3tYk/4LNDbQzGY8x3dMPWatAJeQOv9iOHgvhdtBxyb76ev4CJ
mNjn8URMP79E/xLG8nuOQb2KxnsNBTmcQEfyJ8v1fuWODMscJ9RTde26jEGOF7HoKD1y7PMxLn2s
c/dA+rC5iSXJI9W+/Ru/zi2fkZU8Q+dGx+Rfg7xKSppabLRU5C4WJfHp1aM300VpepjdsCInko0x
mavnqshbi9s1GZlDcHaQY/Haqb0Wi6pqpiM0u2fBp5mldoDLTnth/47RT/qJnMaOkVNjtGTW8lR3
70RRWlWv9GCefVEQI8zoHEkw4vCgDeXA5bWX3bNAs+1PGcXEQzZGu8IWSgojsSjZ6JhJeisIvSd3
YIs3154t/zRpBK/CAxEO47hgDE5841oksfnC6uoegTyLmV9kLzkBNZAJideY26ppzt9Cu1W01lXb
qdNmOCynrIDhRrG5UuaCrC6HW6uZJMXh6ITYaTs7bSwuou1ngwuFVksc4Y73nbf9Rl5QO9Yo3qWA
jyUiXvxeYCnrHXJDhyWw0ZazA0UMr3QAnZLI4PdV2h7wV/AGzYAW6TTGzQGJE6bfoxyWrLL1JJT9
8fXXJG+SO1gIA3WzWiW226WUuqiKDMIjY9wNtVdrIHSJhdt1+4Uy2mFx8lZDPNlO7/tEHptQhyqE
TFoKjYFBz0Z6MY/xnBeypgYMRb5jxmTr5P9CQyOzGD1ayjvmPJDN0ZO5ZjvJlGGw+39nhiIVHgOH
GdMc/x+swJq7rZVsioacqrmyKNdilySOajVhgDQAIwFoqqeyCAlf9o5zbBKPWKZcfQ6Goej8JqT+
6h83xskWNdu8iwM7eXpY4Qd8DjtrCnIIehLkoSamvIXyU8Wf/YR7Iq9MKMjj3oJY30r1TOLPFxOk
Hf3jJJQxb6Z2SxRAg+0wxZnQzkLzG13baf8HTtNC7SkoHExKebRwfuc/0f3K+g6chEi6RUayBD3l
lI5EwGa0yepcl37xpk4LUr7TXitV/1k1R1AzP1hfkQ2Lm/smkyurlyMLRmoBrf6uEysvUQBOCxZ+
zWHWpz4Cn5gFWb9EkUY+ys8hMviqi91mqBxSLOhba5aMohB/5yYlsD12qQ9OZAS8/Pkt74lWCURK
3GLnSVISTxrtbbhwoA5pLfasGV+hLUp4eT8mreg/s0lPzgjhC+kU/Vr1jiqv2LMsr7hg+VcJR6hz
cgJsmJUFdNS6N91lShSAb6Qx/HW58+g2Xvy45pJh8uy1KIaN+BXq90LCLdvVWYMesJhvFTYjO8PB
oIYKU+oVRw3Qreo2EdfEzDH8gdfauLkffz25ymRFAlCVEzUcyB5GL6z0v+2FZAG8zB3yr9Rdmkrx
KP5WHQB7BWlkn64w/4caIFvg/jV264PJTyRX87enP0TtWwyENKYYvyHgsB4/dTN8/G3Ux1vJBfXK
ka74pyHJ8WHI7qQfYPFjAbQO2/T6cDk0qb3cMEPdSo85dFYC+bWbHiGW6LqB4LrVninhmzfiPUzr
huwJi9oLqPeZPsnxDLtoP3VoC50751IfGbLkCNeq8I1q3rjL2CdcZMbBo34oK3ho45iH/w+qRMr3
U+VzPIOjyahjvgxuxPcDq4wGfFikCgjat2oTdI2iZ/4lpfYpsxP4MUNyuBr28WwW+CE12eUCH40v
fa1pqmZCKrtUgYUZKzSfNGubUQEjkNiMxE2DcWTookcx4JK8Np1SrMkfTsSj94fnigYwxGiek3g2
2rxH69C7Zlfq1CtojqPo85vsMwI0BBdHMRNybAgm64m4VW/4XQIX72SPU/iDCT3Fqh1KhY0r8SuS
0PCeM0oZVI7AwTk6jrHcYaMDNVuK2aqUFO/tPL+Po7NF4LwXjAOaxVLSOG9NkSEDsLTj40c+yA+Y
IrzLSk5Dw1k8DNmZLWYqcE862VoE7l4zJFBwZi7zFFdy7VxoJJxrZanZl08pcqTeMoLdUf8+9k0+
dlCCry2lbhfsXYMn9Xi++NR/oMJjTjAhnQ7qoqrbQUedz3trzGrFcKCq64PCH9BPIrU5BUyQ9mmL
Ov4rkbHGHwBIkL0lwEYsFlS5zTYECyGnPMSpsM8NzefdQAqozndKNn1YrLY6nLMDsuuum7cK7bWN
9hz76mVC9CR9xlviXjNLldbzvYafgEJAC/1BFMuYMQd1BcA7TmqcXlYbcZXYAa2bxHTiN/gZvFKr
EPcxu6O4nKksFtNcECdJSUylxRCLX8kbBzV2w9ZB20YpbVIiiXsZpY5vQBs85to+fkRdSQ1GfP42
JBfndoKP2NstCFX+eMkJ591DSIGl1yau6PDjI7Zbosz9yqRBq7moYZ32HMG5iCqyqaYGPc4Qx+7G
PU97xsSA2iq1bpjO3bOuhj4nu3VyC9HQm1iFAZ8K3CnWOC4F9c5Fhz8oCY17AmEFd6rzaZLmt271
oGdj+9F30wKO8XUZV7M4loT0WcTU6cULBKkPp2UqaOKGWlH9Jz40iktW3oWOIiVEWC9wVsRwhfzo
pbNLNpkYWdJiBjx9jU7OtP1CvSq1ilZf3HtMwWY7f2ts/s27SH/Dhw1BJRMRaqYhHsAM+zIqZGFB
WfExRK5PFerRkY4LmHO67kRZx9z5SAd81mUmcQai7LvGD9b5pbCB3gx+9+WYdp8wCcUW9gYFXbS1
DM2LPUKw8CtKbVziBnORiZHkDF+gzkkfY2aQBlGEpI8DNaEMu1codaBqQyHtWXYIlLm3xmLWHAQs
uYfpvaA8Bff4K2N483KojvPciyfRyrlWtF6EoDk7MGTkbO1RXix1B2nrgTjVKlUKnlWMk4YX3xO2
tS3OV4zQgmGJrYZbI8Hop/G1q5NgFQYfAF87qv3++fN2hpTMCfzZ7ZwOpn4yDtSuL8FflvmRjKdN
EP0RbiSbdaCx3SVllR1zHe8z+Exowpo+MyJKHMvJkRXTbXcNkGPZ5xaUKV5bNCGDvTB+A1Is9o2k
VM1poV1+88vDlIzYmCkiY3e4sJY/nr+S8gPCdpYhMkneYNkIu6PkmFl94VYlDVsPil9rV1/1cVxU
tgwhCruQ2EtWNilE9Al2TdYqLENdpN9wQSSbMPrGzsuyhgMvoqP00s7WIBZoY4mWoiRobcpDQTB2
W+wtFrLMZ7NYIfQd0PZyVi91ktijdzLIbj59+N0FAtaXFXbZU8hK1DWKOZs9ofdf35eMJV9SXttq
si5kgDa0l5RTRMTKoXvmnRFr62O+MimMya6GwdXRpM17KPq9wqJ9k+a2yBnAfCHEoITnW7SD6req
gC/kV8QccsQWjB42Ug/FE3YP8C5WXER3qxS6LtomM72555ynw1XmEUd3VUwYKl8gLZ430XcR2nPu
FddyWA+NYS50kBTmleOkytlJ244MH0PQqgQzDlwU/1ovKvUFfgkFMDhH4z4Aq0ONI+EEelmUz8t8
+H2BOFvw1G1k+l4v9kiyyjFu7o34iFNYgkxp9P6QLruebbZLSDTMbC9WrnKo3zlZtTnHKTuFdsIN
nGAwqWiEcZY7KIHFKhogQCpwMHA+fGUiPwbJyN2mGeKMJwQB3kT+om7iEm9F9vf+Ba/nffYJsfY1
Iv4EPsfgVRrs35h3BOFOFWwoX2zsUw4JC3Pci3gwg20LdUYbjWQ/AZmZJgNVw1nCb+sUTfWv9yLs
PDz61ZQDnR1HxFWd628FHUhczQ11EzqGltrqEEUyyIYGigTXQjPK77n6vIR4tUiJpQXzu5hzzVQY
UZb4w2mpFqRR8aIyHig6toxL0+T7kXK7ztf24K19a+uSt18pZ3aHG7/KCk5U9fs0rfm4v3jMztl7
ljz/JmFAM3haziOxnnsCXcROBrZUx2OCZMoRcsEMp/maM+lvTeHwjXENO26mpms/ugYabTiv7eTd
OVDAt11QBUExwo4cA4vHSPlQt/67MfCIJt9MSPx4Wi5+KkTRDlYbe0YAkAbBWEQb/foKGKU8dILX
fwg2C4tgeKHB8o10X62EcuF/mZpz70+HGKnnmcM/TlPT10ES9ZFhcdDCsjVf9Vl0+1/AlVn2cZoo
0fH+paQCRQFQVVwhO2yZL7zBpBg5JrQ2+9HRAVeRkOPRCjP5z2/2OLEqDo9xrRnhPRCTghoxnSa/
y60fgAqS9DKhdT8xd4oLFQ4BqUDonoAR5bfCt1I8IHDG2Qy7+LgSYCeoVDbnATP8DBp3uxQ3sGBR
36yQ8l7eDlRavFovIcpL0DLvxaRzjqE/ucUPyM/AgEA6S7kDH1RXCPaHvqQ/MAeKFVdJLz+uI9QJ
gTvwoYkfU+94xJeIMy+scSXhQJaL+BCwxEo0fLAC2Ia9OMVu8zlCceygwp5YgUKqflBpthiawsrs
ubcsBTg22DP0KlFe7zrsC1PIZqEkHBKsIrBNa6U2w5G0pOdM255goSd+OMKKUksPwoMHM7FGfxhL
kJN2llF1qmzstZ0AY2cte5uFpdT9i8lmzufA2FBCOlETdtF+JH6xPD/mpiVHb+8PaV162itiDP0P
8kuz6Aycq2Niw4aRWsB6GL93fTJ49E10ptW8jfuMRL0ZZRJdGnpUF1H6k4kKAEcGRscWoxXeyIDu
7sIZYhT6cel/tNzXONvglVRbbn3GL52EjSPS37JKfxcjUSk85TVmlDrNVbsOpw/FhL9AGZNZcwOW
Vn2fOAHK3x/l/UU2h9RzOAwwuQCFy/xJ4DWMp9GiBWoK7IA4kPKpHbEOW8H/CmJSdwIkr4JsiSvA
Lf2+OwCNWpIuxyagDOUUkVr7zTbz5JvzkKzH6itai3M5Mwdh7E69FuLFGDd4uT1djB5bz1ZI5cqL
/YylMwTO8fknhzdURVAbp2u7ImZMNgMVOxkOR3+em6s0NcCUbjN8Nm8aX/FEdjd/qVHooqWWz79/
EIUkLp+gniR5T0FLbPAlNlTXpYsvbLnrJzP9KTT1k2uNEhWsAhJL90hBHBYeyFm+pgxaCoFh+dj9
zAfgcqc1LKuGflcwn5bAU+Fhzvd9+5eDRt46z8Tx+ks9xhxxHHOui/aGlluTq5bcljzakskZeirc
bzEMkSO0pYmPr2EE4egG89x0+MIVvuaPilPZCY0q+t6sxALYfE1nq+JW4v9KzsWR7pukTbN1pJfE
HsAmd8ooAHw7AjSgilyzouBFIigJJfvdEoCdYWDKqpkY/GWfySl4yOvWORMWKVaJMTEZqZzAEg3M
vw0lGBmOl8etf3jSfdndFYxlttSYwe8Ye5x2IdMIfmT+NzurGgpdR4fAHQtg48f18SJxpO305eOv
9JqVbNFWxnebREiPEkvI/we46MT+w5w/RP4j/CfmYCi9ixssS+4nnVcNlv68j2sm5KKkEBIFT44I
TPYuakXeixBwRg2KLL6fdoT2FPOS5OQ7fgDZtw+s6TAYjh0zDBbGFDtFOW9ZaMHiBo71VI2D21F/
d3pUhNiFK3+o4GZyLPrbo1153WmaFGQP4BCPU5nBeRZsghGmSCGZRQAWerdhOh65g91er+J+J3DM
PFAy0Ghv7hQ5kqxT0KwNOJb32Gf8h4ofC2QLyl455CupAttZrKVbiyU9FdhtYR4bROlnwMF+mzYb
grJSnAic/01M1DnrNZimGJXEuGCalkkT/Ogiair5WaNDAfVjbb6gS50KljjEMe+FkIAFIfZBkttk
+tAgg4L/LjkvOYF5+tjtR5/SDbIyfKfna0iOzJJA1OqNbI4iR26rI59Q/gexD+YUxD59xGRAk/5k
SbCk9ceEyiYYG1Tiooct6ppdhw9umsNEbreJUNLNe/0qdnCctL6Z7d+zHwrWZghleDDY7HBFATzS
cm53L5ksXmShbiaf1x7CQ3c8Raxkd7bJv7KmPfXxwgxaTw2+5O6EC9ZXFGvEX3ZI5TH+GcuxxqrD
y+Cdh3L8PF+4cS3LL3tPRPa1EoYtr5ln/Vc2M/6fN5s//C6ztwNWxIuLPpxfqjbeB7LGPiIsLyW3
xj+Qx2fSSNQAKnqtIR3HRirZ5H58vqNgceRorrxZ4EiD87PBjwL+preZ63DiUKWqgYqit/eAYlP3
kY8bXYh3KO7294y0BfQQTZtsmv4m4AMGOCMaUiKGKEqJRChMhG48tXlQ9hbemMEu+bv2/r7npNZV
AnOGeaF4Whh1VJaUOI0RSs4+E0ddNnjQcmI7NV+z4EqqZbTbi+0ylJvROvx7Xn1YiOzHAWbSHxQe
WPovoj6yV4YWq17hapQ1lfX8ML3wr45EWI1ih8T8kSQOPv5rkK26TPk+rk6kh1zxg+kl3yd7tKOt
HRk2zHs7R1AC/I2XOnOp9hXJx0cQGVAxUyNLwVkrE8wTYS8kjZ7sHZfDxwbSuCOdyDy9uTE+Paaw
ZfJVsF021oVIYxFAl0O6tGyjBwGIBvUNzcfaJ4GyghYs++nOQ0j/rMp7J8BPBAiFx4O18RbMpkqI
nWkHtrumosBDVpK5l3k/FFYZBgiqBsT4qaDn+wtF8AkPu5z4mAg9vCzplWQi7sNajYIhI/g8i2jk
QJgXavkahM3fA/GJVeOGs19/xDYwP1LeoJ857/1lUYubihw9lB2p7v1szu55gqk8+1Vo2KhqDUPb
nLPnofxtUSa2aawjh6wKJL4rfqf6+0hL5aepIrGLsmTAnOTWyh32lOs8UZ53TCQ8+7pbw79/Ke0E
5yWzdhLleyZfiGpGxAcMWujYN79/jD3csGDvQx7z+ZrAZ0YpzX9fXw4yh8aNr8uusv/Nj+Fw15fm
MfA5hXUO7jB63l9NConkJuxMmzESo2k9gs03FFM9hP6ZX8CPVPTpdCCNkGZAdQuZpkGmEf+q8R9N
TSs+f+q1Q8bujTV44KTEUyXu6IkHlQCE5mtgQcQNJLUFo0e9TZYdwBoCGI0ySVZXo3X34QAwgKrf
U3uv1iWd+vHNVk89onItuUVd8B+PDimM34faK98HoZx8cwfrvmcQ0Mt+WwtSSLvzau2lGam8vKQT
Uw5zjopgjIyZU9WahxZBSl2vQVstsdzVYqPuCXi14Xyv7b/EpunDHzINqQ17VVnPp9Nxan1Qn/x8
4OXitQpjpR8CGKjGMa9KVbaZwG2AJGQNnXvwQFCWQE9A5o6F7JanFl8RbctPtJ9SKvmXCULLMlGh
oHDclRgYS5jlztRQhS8BRnVQhe50Y9j8JrkiBUtq2hTzb+PcvCe7gFi3kMILNNKRD15KMs4dM1OJ
5arzI1ubRBxBsJKH3B0Lj95XB7EvfXSXMkuZRPx7V/1LBovFnCDjobQWn4vGM2DIfZwjgcQBpj8N
TcGW1oDLXPojxnpsvxs+K0MICBiGn0KWfRkkQhBWAYZpjND75Ivl2oBigpIOkIWRHCPqbLSvzClM
cjfjwqzCzAoHit7nS8sPgfjkhKeK6qpgmp6kwMt0P7G0LEfdetl96OZpfqEvmytgBg4XnONxj1ft
qSncWgSNr4YncKiI/W/uX92ftz4/a3bik0Dv+IH0H1ge+QjiigCzUuZJTPZTZsd3jDPLTOjt76rD
bZEqiWTmQJH/SSudJFJCFE31O9EZZGL88JxT/EPG9GIAXELZagn9fMgLRhUZf+H1a1XYmcAqBp5+
n6xAQoRRctKvIXcTeZ7yYrBGTiA6xqNzkw3CgwIOn2WekYn3C9L1TjzBdC95edsAz+OK0YDhhGeJ
Maqx6DvaeyHUUDn3STGHGzbp71nnT9NFa4LbFXCtJMruYNE7rT8+TyqNmePuppvvui9sfCTKGarC
XV61zWyninBQUGj65TXteWscrMKeml4PTi+nf3EoR+lwpNJbb9XKX1F52BE/fjv3wpeERV5K/9sD
oMBcv9SfW2ehvvWqtyt3DIwQo5mSOtt4JJKDC309mUIa4CLOe5LZZkl7eQBYjpmYzwP5H42Y5Qp4
Tc6PBjK5V4/i4VKDhdHK9CzGkhKUJJRX1dg3Y+hKVHnhZzKf98NLrSZiOhVzEZfe70W6vHLyRdSd
3kkFa02cJdfoWyav0pxrx1gP/MnXNVxPIp+2+H+1D818lEQIQ5zttfwTL08slp7QRWUbUFpn6EIu
8Y0XCT5gpbh7swO9melZNzg/KEKsqgnJWrFKQgTmqcMJjbeYsNwSqdm1RJ4QQ+tci3P2aF4eO7xS
vwNpnH4O0PbBnmwhO4vTRSctHywKByQSSaxc3Ne6Z8Fg85LJdtC9uKJwpZDqgDEAVXxvYBxRoaa9
71cmIpveF/8VGD1HXl2PHxGYYpdEJuB7AQPXGhmn3LgQKdqCNtvIZEl+bCLrm2j5CUBYGrRzGyqu
30BJdfWpxD9eoitFSkSA6tsMfhxE3RU2dl2q0ikGIN6wroEzKnO80HJYBSz+TL3iWr3mIhcDTMr6
Wab/JWHExFhcp6UZQHxW/qPfv6ewmbv/TiIE3VnUueLp/BJXlUtbvFutXaqAz9QHg5KUEGY0PdS0
LJbRp2vHwASmogRXbpXY4T7qOCOsB3DBUPDCBzro6pfg7sfMI/+26wM2DlThLJrad9caaXNesFdu
ZTy7djnpcZJojWeY0S2KifQUD0ansP9/X5p7wo9g1VNujnX+bmlLujlXOMoFSSa1NjgKuk5Mfkhh
a1QGKLUKxYIQNtIjaVrwhW1F4OrM1qr7FdGExX9Hmyn9iYCrQe+Y8eSU5Sx42ihIuGg39+RI4oYQ
nmLyiMc2NlcdURnxoLBgPv/JzU1DJrOjXhmNayzfuK1I82XlHovTACDxe6jke8p/yAZZ5wVNbmbp
QppjOJzvqKX8ocbMJLVSH7hoiAehyeEMequcFJASh5A12C2vkeSFy7NMdsbFjwXRRZjcab4P9F8E
OifUr2yVfrFWAVXq1IO4Zb8YimwSfQOOnVc86oPg9v/4wQiC0hzn3hAX2ZkLMtkpTgNZi1FMGq2U
hY5eB/M1UmpJ1oBmE4VXjlv1ke556DCe2fIcjfdEjdvb2x9lqUp2ze5xRwitOyTKAkO/IUw/0QQW
wstkQtWFWV3PzJdQskgD9FrYu87K8kZT4Zgr37zqOovN7gTPkkCPUanMPgFXf/4bHZcuWiYeH+8v
DOwu3lgotMXflxrxT1v/Yn5EWMV+pIAa/ith1y+8DDdRLs0s9fkQW1mGYzW21nC7hz3SgkpG38fs
6qs58tWf+1PfY4R/TVkARR4nhVXFFI//m/9uhBEQF/zCw/w1h2Tr6ha9lbJmGj/9mQC/LFz5kKwJ
HbqBqVnvi+1kvXbfur12r3dmldiNbbL+5IETg/Dse1JmXzLiRE136uEDj6oA7WMdqvHpnUwW2s3L
bf2tuqtSJuR15srGeRgBUul74uyVzKS0az1OY8yk5ygif+kDc3J5T+0XDqX1kTLhePlRz3W6LiVi
v4howsA+fepx8zOJ6r6hz6pm8og8MClEPmUhNMCCRIlXAU75gaCr3g27Jjnkdepy5X2MjWXCEp1s
CgVptaAL+FU7qf/7dTcDnVf2+ZF3ivl5E7SpztWbJ9gfl0k4z6OJKlUbKI+QrCM3Qz4LSbzPdDXf
lyV8i2E3bpEnPOsAESA1iEB6+MRFma1PjY7cuGkPolGMePVTz3SwZxToyrAW6Tjc8dtJjinMmCgd
R7OM+CEd0KOsUy0QnrQK/qlA9LGzPvVEI9pNkOX8WkHStA+B3R/t/ku8NpQt+5VP9Tnk+qTIuIxE
3kYlm8WeMxD3pWMUWwgS6U7Cmy/04YY8IxCGyCWWNQzfvabwcys5cTjx5M8wgGLuiIdXgoiO6kbW
WBKLNqRh6VirWkgVM0AOTmWBjbhuSr6Nb75mfLN3ygXdRhRcMK6CT3ZKfrcOiSb552vckS7QeIUa
/taInY3FBQVcYuXC6zXGG8ubiSG0LuAhVNl45M86kEPh9Cj/HSVbzjTlDH/VKo7RCT5kRLUEqLTk
ECxUWDfuqI3qZ62BkrLDKRpMw992N6qFYhmUln+5LWwRF88Ow0Yxje3ZCKZH3aow4YwteJulK+vJ
44C2SW5FmBHbAFKR6XL+0GOt3iiCUXKoS4mH5ftwQ40xoQSvvaS+zMWqyqYuHCrHW6VcP+IxzxwZ
fPN+XJEx0uwvAcI2lf0J8yl+AKnQQWPmI/2W0nvOQXq22nefWKWWVkh8Cd+dPu9wzZRqnWXS6vPo
zGSiC6sywiCeyhI9QgqAhWOi8WIdgPCnH6YB3Qk9d2wf1Vk/qcFPKwcvYv8HZMnt+uE18hQ35eem
cRIgeF0nJ4yLgGu6EZaVJsgvjYIy+nulGXFd1NRCLUopMXbO11BRWzbz3VEY0O10FRoann4CQZ+f
0AQ79Vdg3GsuVZuhTYjKMZHmeIjnSjbJuYzv4KD0twjOowFPCeidOSZzdk+zrDbOnpkzNfft+f4P
vmkj+1OZCLnnzLZDOimN4hAz5BPPjNoS5InlYBoWtdyMlvT6tDKhKIWdEMuE5BMhE2B1y2uXvMXI
5Qn/chqXTyYRuBtp4DolfVfpsAfy6Y/Dp0ZelBPpjzqV/+YI5R/WG0rk1tsIlREgwtWtDbZ59v2i
seC4wu6fOKm9MVIVDEanKJ4j7KEwjGVGPXwmUFPJ+ZRm5cfBqy28TBm51gFr+RItL5wsosM5FJL/
StvdBrrPPk3KSPkJ6O4Uo6JCLEk9XvBqu3r7Pjo7P/IjFEyoqSeal81fWdeS87PRSauWVzp1+8BB
LKJe2ycpkYcq+tHH89d85cmCTnjdjTt1UDV0gvj2ojOZtnLbio0arH7XiDX92tDt7rsfAdH8ltzj
Y5ETdCpXbSZaNIxKKlFqQgvLNkzwaj20nLkA+vetUqOG6F9aP9/UeGDCgtXT6JRv6d2PIWjWz9f1
G82A1VjQ5JevYOpFtJ9tLukuONIt2jkMAed6p6dMxlbltm38m0h4IQVVAayajGi718TXBKCPmrdC
4Bm0e/QWEcdj9sZOhY+gANUdMmRkonFyM2/RoSHJAVkj472zSjaAddCXcKycwLk+k+FxCeoNirU4
pbJL2R6hnOWpv/CK4CFdKgC3Y5tLcHJivOCSoJ5I9p6EhsPXnRrvVVeHVrol/qkOlnq3h5FZEPyh
yjPgv9DLuZe3Sm427U0fR7F+xodbKFdfKG03jn0rrm2Gw00YJ3uzbMn3/QFminmDf2tRsN4UNhK2
ssI0CEIHGScxH2LxLhmbL+KIxFmafXcozURUwTiSLXb5IG1bMtY4SRQaix7KSp/D1oSFGrMZvn8k
d2MW1hziTh2LuBs2XfgyYX86Oxbu1wsD/VrakL4lwbqe+HdrYI4Pw8cQbiGVL9rN8by543hiSzN1
wk1l6TWXIg62giK0qVDcl7zNbWhyQ/CF1VYb6m8nD8XR3uYNMavKoCQrFlH7s5dNGEb+0Y27nV0x
r9Kga0nTnWSo8k9GoDZMBGvjlTyDmqnzaqkT0A+DcDShVdt3F16cRA4Q7NEhY530Ibk0iAPPc1Oe
eIoVS4Ws+ak23ZB5IrLR/jGD64PUXPBhhDuk65inc3PO5sUNkoT2eslVv1wVXU+XeAAF/r635D7V
1Br2M2l3CPqLBBGIcFebMq7dMDnwORlNnWmcm1SSQJLz2ogtJDYLzH7S4ujqBzvtc1dTjCdafVcp
FwFlvi2y0hl4lxDEv8lp1i3jO+7pT5cpQvgmvpZAbF19DEnJWuSjTPpBbrXF4tMnm6WUkmLwgN+i
/2OHn/Uq9x7GgZnaLvnDBuO2QXQN9xU4w5gOORUH1LHAbNpXBxpTT4NpOjOWZ3VIW8Iht2xWjUkr
JdtPALIu4G1b5VyXcFVk91QRzWF2VtDbDYVDM7Wi61cPhA8SSXCZqJiAlGcbBkdJAFv6yXhlgv+P
p4ycZX6yB0WmbCj291Gyf3Nhhmk/fGksYMnWAc6FL0m0IG4A0WtrLxkDTePbgnZszSMCo3X8Mpl4
y2hNtlWOlxkgXtfPn8mdJUnToGryDTPyxMLcfkT77UR6lAMWxUbBF4MOUJwXoDKF+nQlZoB/GJGu
LFF19JJpszyRQkuaG+tn03Sol6eCwcOORRtWMc2RxaRL8UhqhPdcky94xIEa+qvLpgUIyg/94jdy
XnRXgiIZZS+ZtH4IkxwiVzfPCvygMUbZJyE3izuueXhxOA4KYuUVWkMzfNzAExYpzRv1LpjeqIkB
OtJy4QTSn3QIeVMjKlCBo7g/1rlTojjvuFO9reZs3b9nwOy7FOE9zGKZmtXOuFVN8q9iESX/JM3g
pSriD4xJHG5+eeeZdl/3rQ71IErQt4J7z6vn+UejIE/OZyMI1/Hi3mCHec4s2XdLrvMMp0/ypoqs
Wo8iH7g3W8ZWaC9v9NTGpFh0PhwUyQNf21gawMuBmuLod9rmKMGT6L9whbRcZEavhOaw+cO1+8UU
zmLJ/ULFhn57fGVGjcJXmXa/V07/xKUqzWIsNDwwwnUky5x3Z+HZBfVTxgsc5YIXGzKEb23HyJuo
GuAswBDzJ7J8JMrx/AcKkRkUbvWe0N90750BYFxnj/B9nJ7moFbZd16VrALwRSwLC8YrXLG4WIUC
t0S3AP+nbeiw8VPo3aCzHPO+NXEvV6xm0o3yvBiqymPkvqyzOdM6tfAT5CB7Su6zUUT9ZjW8E5Pq
K/i73C/KGPAA9gEwysVI2rucvTsIv7xY6/Hhb/zkm7GH7dBF31hU/xI/YN8Fh13FNSuVLppDBlra
yIOLUocB17L8M4UWJe981jy8ILvo/V9DJwipQ3BJ2q8UK+zEqOXQUoCFwB3PI267pkbTsfT7K4mT
B3ztzaMdxX49Zi0FaSjZS0Ye4Z3vT16ATLgD5HvgGt99CBrni2ZveeDYCnDvSYgZJ0u/QeDFb3tu
sG0o8iyES6eiLzi0FMsdyH/LbRVNmWS7o9QwHrZOBBYWFCXzD//HM6h0953qgiB/69lohLVRSPDR
U07OEnPQewG6UzbyOY7VNcsR6ca/8TpNaR9+Jp7/cfhG0Q/skyJRib4qYLsuaPx1KJaziAArQ6q4
UzmXoCwLrOh9foVWbq1a5p1akm7Su5cNIfQm6IVMH/XdHKl0YnbvgY3qFsTWXGX5LSB9nIcK45N5
MkPPUl2kzaMacJZFXhj9A+e2qXXvJzXnynb/4sdp61kxBRIS0gcD6DVhCefhRmyEi3OaOZ1gcBsQ
hkZzzwurs99JJAxve3MPsOHt8mOFv7RgSu3ZHkOu4mp5+qRzXJFauT+xxeep62wkhpjjBtxQuw8V
RTipGfZBEYaIaEGknlZ2Ypr4vj4yjOAT4v35jPbz1Fh8Xf6l+LO0uKt41QaOjgPIe11bQdk0nhiB
Jt32NVbocyO+58a1TSrhXrrrNXhXe7BaImcqO86i7zZvtjO/TiZjBmXgryJFy2bI/4hglOrNMoZa
bZ+Dhf0Rvxk5gQr/M6NdWpFNSiOXWNaNJp/FuCEMQ3QKR61RhLSlSfHaaHcOV4TUrbGtFaprLSua
Lm6uVKYiiJf7lI0F+Re1PnnrFEiF2jRGAy5ODhtvT7vaYnDpWm31RgX6Hb3ebo+p+/DQ+GTFzuME
f7YcVbffYyk7JhFGCnidl0OV7Z4JR48zXHjsf/ylIj0U9Qu6hBHnF0n7XRgaIgaWp2Wo7/443aSO
HJeGFFfm/5hJItQUrhouclu3NmSS/h/GkMJxVyPwiN9lZw0JFHMD6EpNPfFejOvTziw7K/zan2UJ
KOCCT7SGfTKBwm2+OP3juwmM4QuQ4krw6v2FII4aPK57Oovrdc3DvHkzIRE/r1pAkBfFuKHek51J
3y/kOqyPYFH82TPyzJCBwsIDRa2ogi5a5KHCBw0m8E5Xl5/HOZ5fykNsywyfIXkYritcgcIXaXRr
BkGSxqtefape91Bkqloy2F4HFGDNP6/dX442ImdssiJ0ogXoo5adN8plS+e381snXziSTngw2QWM
vJiDjhAZM2qYY0F9eNs2qokDMKRjg7KqATLfoMVzkeqHsYSJsztK/KgHryvJxbesspxHlXPLxBEc
lX581Gp5GE5w2GCuV6NO6ETw2+1M90HI8IC//OO8dciXRi2lBMoofVX6elGFptl8GGt3p7YfjWZK
fM2fpWCbAU9ylqRtfdB2r9kj2ic9MzGOD7o3UAH3tfLMadHuLBJZAUrOnqUXTfpUiNbRKG1VgD0h
vlI2STTvGvfBYo6wAVdytZVqSJncUDyZL9XAwQyofavbORnVaIADPVoljECPsE7uGvC7d1TH/YOX
1chEWQl5qXHVAIT4HxlDjVM0kDAZBl7bfMGLfKghJOEloZFjkdRjFUf3kz2YtrA/Qf9nOE1hUW+Y
E7Zx/TVGu+5F3XzAn9iZovy5WiA8p4PH4OKcgt8m1Y901CbupyF2VGpD5o7vjRxEJjOXxBeHI5uu
PDQevYlDKLmtqCi03JnO+W0S5to8M8lZIFjm8alFRV7/jXVCcLrQbihtGiDTAQxc6UGKasTmsE8V
p8dXfSodKmP1f9ctqHvHLLbGrEAJ6tBzXWqfqBdhUPVfEcCP4bN25KUWdXKNjpSy9plLU/s243jc
qQydZLbMGWmwormAGI61+uL07HArMidTSSJRcdLtn4j6zoNPThbrlktswA4MoTeJq1INnOq90wDd
xWT/uC7iHyQ87n+atbEz+8pL0n6Ug5p1bMYinavaG5WOXxkrR0RAYivqe2CU/JbcvjKULjtcRijs
L4wCUO4D/fEFZH2hy5+RzLyd4aHhL1zwAh2GEDfFy1dKNUOiIJpQKahtWkkICKKJvo1s2wLgEqwC
Gl+ftGU9i8aY00sy+fzJnE2FDtnw0NOcek7KLeuCOE5Y1U4PQZ6707mrXxq5+/27mXHD2RaFRTSx
Kn+rRDZa1i5aoqsDOSPkjPBfj91Heq5zwfw3kEc2CGe2KIsBQDtfjbSZe2jBrorMz229fmsPUN2V
b0dGReKr1IG6wSyjJhev8R3ZEn1cwVN/rmNfZIi4gUF6z2wa/dmAcVv0yQPt7VritGbCuEUT+Nql
epvc+4VSf8uwN9Ao2CBvrWKeBgvudtCpuwOean2++UbQvwCcVbGUk5teFzDHXsFKjFsJ/IMNMcF3
//DEElyEdFjoBUJ4iKmGfEG7tqna8hsp65jDVHVKpwSmqSTk5b8VpI7IU1bRn+xdL4yB4nG1cKJM
Y677QWiFmMTjXpRgX/inMyFDXbLpRwJQZwKLNBPiiscn8q3IjTLaimxRAppdC8e5Q77Q+dIiQyYQ
PNBxsFeakQz7OBf5gHBpJkFKQpHtzz3kziy/t3jqmcxU5q8UcJhWZb4FSa5wH6EQnpdPN/3UMv/G
IFirSD2oarAT+UvPp5O62f4WAa044YgvQsSaPYlh9I/AvWK85oQWL0NGtbHsswZ8W+eOQHDh+jDC
n4k+lJhVns7bk5/WjQL7kfH1GZSQHn0fM6D2LRGslTFekKGm/uP86nNhAz0LSroRvEJkk0tf96/9
jQPfq+e43fATE94VFU+8qXgKGak3NH/DLbtSP9TamBNg0OT+/h0TRXJqmkwKzAhwbLD7sUYc6w8V
7SnwQzI0MKvLLyRs2WuewOEJnjV8bmln1y4226yhCKqc7srn7KQyddXZyUNmUuI/HB+1P0kg4Imb
+QtX25A/R+Z1zW8+jGZ/3YJrpTKxfm10I7Fs7ZtJdc5GsQ09lr9gR0pZim3Nbpcx5UzDOMp7+B8q
l5Lo4ve61QNwAIVYoDpxioEsuMn5F73qESD7BAnRT4WeU0/nhtOo2tqJOLSIua0jnEQ2T6fHV31p
hWtPu+dtBk+8ZJ02cBmBFl3HRet64e6O8tXY9LJC/ngBwAsUBeEDka+4/APEJVHXxRrmoCzyTMIm
84WG8VrE4I1Bnezk+/M2hZ9LtCat7l8kGBAFolxz2DD3YUjLqvlRTukAXE86J0DB1+k6SVPYc9qV
d/gUfLo9trRay+s7iecf2fbZOYPsD/7AZPoC1m9dyP1M4tP9GNyerOtL/GaHRi6vr922zXAuyHie
FwhZ3DjwTtu2uq9U83PLbZJ1c07wCaE1U6FnnezHNqEHGasf5T6NcY9lxQsMJNjwDijCWacgmWr9
aNbp4pJZ3olMKzvX8T884wNaHUDduo77Wup6uJgzrpZCPPgjRVjXMcdlMomk2AWJrrGJjdt+90Wx
UlAtsVfI2D0pLmn3y+mhjRoxms1KX032pXrPqEqUVkFX+SxNsIwx95KOSMtVa0AXkqKW59pZ5I6B
JUkvqoR+/VpFtSMQl/3TdXwzEciwYVtPk9wEoD8kRMcJdb+tWXywe/GmAYmBcP79E+qyu+ZiQc9r
AHtlg0Fev2iI7hJq2Ib7/uGhPo4PsOTMtjPyRI1M93XEZA/7gwJOOSknbiOv+SvXr6lWXig89gPv
Gf7V/wXxO4WXMGSsQYAkqsNnAHiHHryyeRcOU4i8I1KKWRdef8ZuObWXA/UQNAjfFUn2k9lHhSS/
aGftptYkxusL26RJZOcuAeQnkdZp0f2yKIPNKHb7RyYI+Ga2BcFiUs/ghwrGTONgGZA/971RS4as
S4qiwAq6k0kXhSiLqdKuJMsGdaq7dP/z+iRG2KaEx2cZWyQha1wiL1cvscVGyls5CkMYyUbhoAlr
Y5OH5xGSVhqQN/TY15Qw98XHZ4ruk1hybcbkfCOfJ8CudxqD7FRMEAnAqT5izC7/UvTWZfBJQcJg
NtEGEZ3vWlvAPEVn1oNCQSxb/xINmY4FIdzYBUU+FhxF74I9d//7BAj3eMTvSAg6hwNBDuBaiFKB
8bpvtakZ5+h+ts9O8Xr+jb79qX/SzhDlhzh5RZtyCZXLlD+ULm2AuRdq5fs66P5Hkteqd9cquv8K
fi7sL0lPsUWCwirAbLEcfU52eJO0iiAe5KTcJMUG7FUSKfDOPzl44e10KmSibcN0ALAtR1d7hqN5
kMx+LAfl9rn4XRAdiUr+rDGSPqdpnMU6ViuDySn1AZQBW/ot4cE5Eua2hVSx4Dst5okhFZ6EawCD
W9lttJxI2c6BpKkEPHPsbU1TnI7mG+uZ0OmFey60dhN5qbX38dR7aB60yOOLwhVaQ2BtO/viJFiF
sGE+nTDiYmPvC7Nr4UF3PwFaf/DZzfLPXyc/J5zPjfUw2Sk6I8ZAZSsu+N7+gRvswbCLymQ/8pEn
2vbN6oK6bdIA6flV7uZfr4ZCi1+dKgFaK65vgjkvAZhSZvpRv89WZvYyUXSyClYJ4Ubgqfih01Sl
rEnBrai0lfPl8hryJvSTBvlEB81sYBjILxoGaaLui5+OdcCTMlHpsgTJhnohUpJxh3KgFJQ9qbvG
QROnjr/j6ADv2k7biUMeGYZ/+GuWf9EAPnzPCH+q4iss0MS/kAaYwkBAH2E7HboWNUrCjFSwE7sM
lXF8orhsDkLDcojuhnoNxYJaf7VIwWLc4iHXNYPyyWPRkFDM6YiOmAoclb+LenuixXTsgWuo5xIf
4RlvH/B6vhEarYJMUt8NChTySlGt8PyxoaoTXgEprfVy9TBDsfUCkjPliLKZLEQecCWt/hGVRQWJ
18nzuR1GBbuKrcmMDWyTDxfBlLoadnYVkFooWUzEgouNs/xV4vH4siJ3eq4d4Yj3q8hiyuXemWJT
B2Fn73pmyhdMSits0r1RkL7fRXMOg+I//7kd9Q5sz3nuQ7gRNpu3uITzb8xdCWh00xWILPqBSgKz
uaO270U32Sa84Mpe5x7kCEqHYthbUYy6FQ/9c/dM++vHbIWxJvxwV7j/1r3eUIwjs4S/epuD62JF
ET1IUClPiFWoyDHnodDZ5GEeU7yDbZ3XR+fPijuQmfxkX8us5o1p1WjibyqyL6Lr1vnH2h/vmAz4
LORFFfKOzUgFHC0qcbRNBH/rqrSFAqLq/c7n1qD+wQ1VYHcK+ctdigaqPtF0PV40b6xMTp5C+kSX
YbvuqJW6ibZ0eAL87RH/vx9rCcJCV0BgnMrz7+2c23BWU9JCciQZZcakm6CdUI4Siy8aYcgU+Rt5
ForzBK1VkhSh2s88Za72Pm+h5kVGaIIZq7ajD0O0THEgSB4AWWEUbFpECjStOxFaCvBY+Yh+hgDk
wTSt8R9KhBx3BaVbjOIF3f6Hka+9jNO9tXiHazbIqq3Uc5UiJ+k4ybMUtowkcM9gUcVnGMvUeJJc
AykE7jPFA/E0yE/O8jYT85PwNSSgKWNe4ApaABUkBTT8elSchOOUKNhqNYBn2BqQF8FCZJF4ZbrN
T19nzr32Jdm+kqU5tAUHbUW2bHPrm1t8RXl+JgS0S1Dc0JHVqjWmt9PKNPopfMxjKetNfR7HETpH
EqKfEH1CRm4eFbqcckoUrLfc1aEv8OyDItb98CLuYnh7eeT+P3/FfX6ZTQNe1V4gKHhErIOHzLKz
5dmWkr7kEt0JwXW9897chiUBpczd39hihRsbkmLw4zVEjVC8jeI7u7L3Gum0NhC1C3zZMDW/FdfW
rsMP+js37C1Yg7TQGW7vBcNO7/gc3/fHduWD8eyrLZgDqz36DGJd6Pw1wg+lLZykSUhODJQOp0Cr
dhHmH2wj7MsRcPUElMR4Az9h0CZuTOE0JMnAgWt7RXJ3om9eoy+MgEgeXJl5lpshGGIQOPKFPj0h
7RgOlsVgloqrIzcITZZPqBuObvlZ7Ah1lUJJQkci+ieJ7P6K/2yAsdRAobnEjhAvnmL1cW+aJ0ja
coJ9O9JGYJ/VbbZArbU5TKXvIuMtOtnfbstLZdYQkPAyJCQT2ZfCpeuJYC+nHbxlOY0kQPd/SpNq
i16u6KyWjkTOo0KKW68yAqtIEmtJH4+pvUCPSU8lOx7pEkt+xsSk5r5NX4gixtkI/T0cpQoDzfcy
HGkDVngUISNAj+mv45KPVoCs/cploIumFbzyAc8b18riZ8qQG5gnWM/LbJNv39ae9duru61pistx
Jo3yWMNUjRkFa1WBkp5T9MIC+Ss+Iw/5SgKey7Vkm5pfpKcTDSoy4vpSJIi1F6zLuz8wMstqINOh
ev8/j+8HWw/f16ca5UbTR0ZmIFcqQrfVZaskOut5v07vtlUYcPWu2TNz20cvQzCfvWLDmbIClPiX
7RKWP3vKaDDRduqVf9IBUFCJ69B/Ua4THqqGUMRy5fKUN4sBYNQxR4xjR+GOXl9Y03ON5YptZaRW
mET7w+lZ/fG4qDX4vk8hgm00D7WDe78nJdwVsOLAOlPgURnxvD15apOKSJAlMSb9DH7u0MBosenn
H/Dzart71mtn3zz6sNziSOKhwuDA6EoE0cncIjlcJq/SudQufwD++AKmAb4HeJhoZVxMw5KWBd2G
VRcNUcaASqxK55VRthgZkb7F+udjzWXnEKR1hX4Pdl+0OSqXsSj7jabHTNbmRzUvr9/TIQ1kznTa
OD8hVIZMf2qrYXcEvcIR7W9YWRzXZ36/b4MXJ4atNznkuo5KKWTYBcgMnRwQMdwfQm0TYGAdt43j
I2nnDzuZl5c+mg8Vs/tRV575rgBVl5KuizvvQ+0vnOv50GAvJScHA5O0gz232VyQyVril0gg49/d
z47LXcASXU1cXC99bT1ITc658+lSi76kIV8Q4dj1tGrFuh3j9/y+on9M0alX2WS07BnqxRroEmaD
00YJD2Za371DrqMPXEe4I+ECqWJgCHoSIY9hYD9IWkkH4IE1vmAHeF5Dj8aXi0CnJb0y1lhoDkMD
Muxo8q8FevloiY9k+gMveiduWetwhUI8bYmnQtguwxAJWwqfUPp9s+UeAFgRERENN2X+zfgAWVNc
bInAkGvduk9sf9PyhZTPaHtWlQ2yXOc5h3O4bisEOIQOLx0mGXPQqYOTJ83ILnmsFKUNiDxjG9nn
g6Fa/FcaHMVh8d1NrhaM4Ta+Qq4dh9xwH/50VKdXdkKu+Oz+mIglspcb0Sqw3BsWHb7toKlUOui/
Z0xcjDgEePYe4fUmw4d1AHQS9200+7bX9q+O5v7UMTUMIRuPuBXy+IJgUxZ0fuF2C+MWRZziUQoO
V677qWyETeld60aDpCzQiokYq5Grxf03imPpgdj1kDcgKHMKH5mn/R0zZNiwYm0wtOXV9UUuarOl
fF4jk4WaSZIilO2uWdCtLtk7/EgG52QPM2tSINrB5XCT8UY9cGdcfNqbda22B4tO8gOUJNOyNgqH
B9p/eK/RKNY2ETEYG3WY0JJxTZ6hktgLCZvF3r9iyDfywe1Jeoxqsg/jyAJ1NjGDDlxjhoD1fcHc
pcC1JfSg+YPxUh+cmG7Un2HW1ryySIeE+OXsi3qiW5I1eVZYbBWZKW544G2EEshovEzT351KT/n8
704uS/R1YEcF0SU7CKj929zlaDylrMjkzRupTV4o+qq+gEn7Xe+7538T1ynY0xUCn3kibLgPJYQc
JsKh9gI/tZ4DmVDmuV7/lnElgT52CUCJDPMLCkAn4z6zlX/vZnkXUZGMWYhfRcrSiapVi7Ddu6qH
PiAfCxeYxLNhBkvLxtmLAys3SGV7bfgK8MLmyu08R6C1ZV+EJ4rdtyAqaryO7gOKUqe3E0JovAPG
SRPsasU+N2Hk3rzEQcuTpyc3gU4y1PLpMCwKNVIVesAeNhT2AC0/LDCueEDOKBsBMLSARG7cOZuu
PoXL/vXFUey9czhzUeWHo3ezged6+N1FaIjWjv+SYm6fai8fZVp8g3jqyDyFPZuCKOxpq49fCnj2
Gxg6iWT+5gzI5geekEzyzfUaoDnLdCWTAroBqFyO7vGIvsjwLzOdG8RTWTqaeJmpKDmqYhMfWhzr
WsTsSpicLPkCehxdu3EXEI+B0FqRPFFxjnd2W0IIDIByacopO6hSCJUEIhD/OYfv7yeocWruacch
PTwEe2O0IvIEbn9GAzBuE9iuZD+MGthoYhrDwFk7WJKtcKJ8Ets8Odvy2T+fI6amdnJhvB3JBCHf
56kM1VX+j2P97rFu/HfUc4Dv42Iybx2KSBebhAvHW1wa3A5N6W97nI3OO6ZIqCm6sAhr+VgKO3TS
38pDo357HNFAppj7tpH23PxR0RczzcneayUYCDkz6ub7y5ctZnrAva63ID/JE8dpiOfPzGJxavsE
KWWinbkGpO7T5ZPTepjGacFOunDr6CUwot4sJgCJA44lWKr140sJA5g+QyQ0saQ5J6iVWs6HFYUG
BNgg2KKv7LYP+lOD+grGv2ELFgFHCK84ji1geSmfl1AX+yFZNwuS/aocUHmmxkB8e5ZJygUOMqED
P7OWT7JN3FoW5u4zQg4kjF2ur5Pq8vC7yDRXIOsLYVHeMV+v6SGFh3ZqUVc6ZqQdh3t/QPG1dkwj
XsNWrjeoFydp0B0vvNRTb4TrnQyuUgDM+cUsth85LbS2GagHv0GYFJGHjFNWrLqXV1GlHZd3pR/S
NgOCBQdTomqfmBr7RbVG3p+Lid1eO9vdEotsWifDN0yw4WWVDaU13bUCguCAXc8WKWQ8DKqMxdvi
VRjU2vF3Wd6aVP0nPgUynamGyV5tUPUj6Rx5fw8IPlAIM8J3R2ha7lR4slxXHcoz5pKCF0n9jt2m
Jw2Q3JFhAec16R+4F7KJIibCjtCji5ZvppBXhbnDI79GFDOjnQAZZstVeyOWJA5fINczUOJLBedZ
kTG0DdkTh/g89QuqIHNo1D2+srYNF6kv0HPmmB70B9+S6cPyGT7c6y9DNT73sJqG1qM8+3EMEPNj
HP/HX5Ls7stE1wXkj7y3Y23EBUTz7ZnLrUUY98FGI8loAGARqJKreiB6y6xqfZs09N3XXEgjBhNH
LFVFS47z7Rg72Gkf0Hipn24xmCQ/mTIIm06kbNnYK4O5lLNru9yA3WSwrNrkH4ZehWgjdrw8ol9I
VTBwYu3ANEYVKqxVsE9ckZTevbBP2oiLlggGzpUGXVd5PGf+t1lRhH4MATVdRByVNcIi8tfPVfax
t4uD8ZoQ5TT7odt8HrSkTGVAXuCqFMWzOYj6+HZRj2wQ5tttuDHPlGlu73US1LA3wspW9MKM3fix
KFHOXNkF07rn8B0xXk7cBHi7Dl62087XQmBrf3SnQK3Z4SSV0XEzQer/4jgZjdoCSvVpy8hXeOoF
9hjI7Xs/vJXnPM7CJrpi8PWr+YCIe0BQeZyc4UZHOadjCFWZvOekbB7/EWf1E9emh27vUKdNlXcV
KXhdIFHBzlz+/iNsdm7PEF3YN04DAoAune5kdp7+7CsgGe5C2MjtwwtY3HzY8tjqJVGsat/jts5c
psidxaMLqbSO9qORu8VnsT2ErOhcKkDEqQgWLckP4WwfPZZbPMM4dmCMPYm8qZfrDrFXJsaB/+T/
62JZ4D22/LQHiPJY/nioRm2XtiDcV6h64Rwib5D2mZv9/pfFmVq3hdKvNP1q3QaDu6+aA1Vl0jpF
2Yr45oNd2DLOCoouS0/0s78BFs9Pv4UruC5u5x9OwFppDFdscR2aNBS6dSU3oUkxMYxeQ0XO0WEK
6Ts8PWybxqJIB8Ku7vYT1aw1g9wUkPuf3rnkqUN3x+mzzP6OllUMBhY1mk/G53WueZL2tuqdlxI2
Ne6a/WHm500X9nqhwr+ppf+X0xosOSD2OkbeytP8AMfKVzRPSUjUZlf4IOE8Q4ylli/abPdbp7MM
asJYFmbVETs4TJKX8NBk/4cordaewNncyKDFrrRNxQX6sqvbH2TW8itOfQcpQ3eEXQmEwyCG6AWh
bMwo3TS5Of/uBk2obGh2ZieMNQWX4oJgLgDnG3xjK6dcFfyq8pYGAuY5qMSbwNSH40ETSgOdOssA
m2mLTv1OXZJEG+ELrlqPp8/Ejk6nhSG4xr/ePXMyBvcFsSH432p+FEMGZYFudA3X8m7arK4yJl84
8cTvO/LWQS97xlPWLEf0+YrbWuPHDHDZw43Nhr4vMWL36dWCTeYop9eZwumSbNAc/oqgkMyjkQTD
rr4Q9qlqvKp9xSZKEL+9KWj4UJ/jLja7VO65lLeZZfz0tWQ8XUxlDyepv/ia7dSjO2ZTv3RyO+Bz
R9lAh1yUiOSWFmzK7D09TuZeohOqCjMMvM7Ox+uIF5wayAVYg37Zkm5nFIDBgU9EGrQXfR47GWD8
VNZ/bAzShQtpxLXiyKH6OwSVvFlvqXgJxU0ysuOfO4eU99IMcCM2vcaXySAkOZEL7uHz9uZWUPHp
cxmq5/A68hmPeeWPQlp+SiodnoImdKFMFNCJTnYmrXXeBT93vS0uI7J08Cid1NcJB4RdRrKsq/21
Ozl9R7jYFj6EJ5EUBleBwbjOjKEs2oTtyTRRvXVzZGqBZTYnEO8cUxdCi7YSvEmMbN/6F03txEiV
KX54yzzaMcGrteJwMh6tHntys/8LGXc0fR6XqIp774P4MNspCrx/uprtlWakIydOWsYlulHmXnnS
0A89oMxsph8SngGLp0ZXF+2siWVU0X9N18h/NfmM/MIQYs7HBkEEtODlRwIo04BJO4J4MUnF0vs2
fFpd0y3MZ8EvdQYYJxCvxXHqsP0hX/v2fAh/kayNWWxohnNII8P1vMOxf6ExY6vbU8W+vb0vA8in
miaBs4lRJQMStaSMHcKBP1t564DukaiwTDyXdzzxrvCEHg8sM8WgieZE8Rjz8lzHPABJdY9SXNyu
u6AHIU+MOeMUVjRa30RJg4rko1vwQwT8F/qTPE5TdX4xkNlKJJdKPgfh3Pgh+hAyNoxd4xykdCXu
4m+rAb7u1CN4VGVI3nIwJMrMZmrg4TtGA2m2UeYTQ9xreh7HF43aYY9ZxDgJQl6sOlZF0YCZaqlV
0m1yAe9lkAs4mlzRWZozd3jCrV3rmdeUAdcV2JgJgNihKm9FMKCDafi3e+Ul9B7TKHAJWinEyByO
VNBFrtRax2H6O613CWaQOdEA62IWOe9kT2EJWFBh36itaI1BfSjgunHac3Ut4ZTm/ZP3pbD2/k6W
qF0zk4DRI6eVBdvKoZXwVJqRGGotVIN6ws5K5QztIWDiZuIlag1EQxMiQ5BRyw2TOde+D7UKB3op
JESp+LseGOwX8x05FrSlOQK8Zpa39CUtdshfuQ90vG2CpM7EiST1PABvzqJxBrHVXQKH/Wn3nZ5/
+/WSKrXTprMwwiCnIIU1O6Ly2U37RDUUSHC0BF82Q9PRqA7xQ4eDrtCbz0wjDVT2cbjzdKsIdeGY
H9i/Tdb5Kt9Pydy/PQBPcIpHnCspSVM35FDnQsE/i35A8iEeNfcc3r5p97iTHGO9pwIH8lMS6XT6
0qVE6bIDwemHB11g2wrAbQbxIGhZX16dLvcnq3D2ipGwXCxd+Z7h/LYJkqAOTJ2EEb9tkAFpDdTh
xGB8FHw1/y8FZX+SZv8dHtanP4ywxKRK6RrrIKtmEAbEhTAnlbg4xeBbahLEtQErfson4X10SUvK
mgRgbkE9PsJMTZfrxhTt3aiXf9UXCUzLms2P0kFFmNiPIB68lgC7yUe1e5iyTIDoUW73Js1vz4Xj
1hI7q9ntvqYBl5hD6CICzUpK0+12LcD62FDJe6k7RO2p7geIn03GzXRW7x2BU4AS1XvtBp0PV1I4
/tKOH2BcajwKgwiquZffuNcA5Thq4vWYhJRB01ID/CgTtuVn9lf8WWBvzWazw2OfrFI1jYKi2+GA
Je0kEnIg2X8awDckkmtwbgGXlpcmUpG+xze1NAlvNEMIAhm8DYdfh2h2Q992Uo8Aea+SbGd+jpQm
PjgbL2vK/y0iRBvS+ssTAHEQg6Fhg94lgwl2fEANVnEkXez/2fzkvZMK54rEBL9tGIt/2H+R7Ych
mahnDNLsAk54A0M0jsTtlAW4sL7WHQIzlOU143enHOCkQAiz8x6gh6PgcpTGNLRlrBHoR6wQ+4ux
jNnL2waVFaCJi3axUPy8LazKUQ4852Aqw9lGJxna/qldUFnsjOpezCnd9D2BmV51gXCO6LqvaJzK
sMQZXheWuAP2LVCqtALf+aVvSNaY2eHPNvodaSvFjlTnL6n+P1rxwPfE8r41MURXZGXwmUSIDEpK
tL3KlLTOFYrUp41Y7blxnnhmXdm1M0RI0u/72BRAQsxPgrxcoXufMF4NIJxTFC4ReQOvoF6ca5ZB
5MtDTNe13cB18qnmNp59pRL8PPjKLxngS76j9dqJy2eUaH/EOir8z/uSbTNubSvuG8C3TBT2QrWX
3Gzw88tI/3YVPt9OHiZes4GngYPJlAIw7oa9Lu0PTWQuKNVEVLuAjW4m0giWJMIajB5ObUV1d45M
HR1mv8/1s6/ajgnNcgbKZOa8N9GfO+e96ixhJNHYb8VTDUKrCYF/Hb0eKFZ8kpSgXyvRBYUOaWCv
MWMwDpuCEnHk5GucR/6Dp3Pdsqfq+ZX41zx40zu3JXTepes5+qmhoi/kFblHkF3ahmR4W2e609FG
Sa6UTonjqqzjzLNc8aJsC5GlnmzC6RQv5QOrw8L46ouoI2lXLBfmZ7IBGeYMt0nxvrKyrTAEeCMk
tU7czmrzUi4cllMQ8rvVnH1auM2MI8Xc7s3j2BZ0zDJ8XAk0OQ5NDK8iV4Dd9EGyRQdUWcVz5Q3R
/lIZXMyeO2K+Dty5p53XcUhnJZEAfO5HcuLzhj19nBR6UJo7vxFjsMfhN6cnB+jCo+lOQZ6sG3d2
zLoY60Oi1/01tkPiIcp/nS+q4KN3Pu2QM/8eTqRwT5eM3vafegaIhnpjL6hSlO2Yd9pneZwYNBsA
gNq7uTVoWAJz3GVV+ApMAhOSvmnIA3VUmLV4HvqqUx6nnLAG+kVFgNECueXiBkqu3zUmXih6o8og
vj0+kULs3ib0iA2R3Vq/fUXoqx29/yAWzUGJxrvsX0U0FEdZmOdINNAJEOZITeg2mRNxmOu0jQ6A
oU0bwt9SNMmgi4d1YyLAoC9QMLR15LI0y25EyY5dMttbLjgbndmyk1g9YKu199OqXv0la412rvYy
rKmrkTxnNQsEQz/V01mivJrb5EGo9pU3EHzFCKo7wCncObJUU/ByLlvoOdQDXEXEhGoFxOnKdvKp
JmbZ/tl2gThQVOTP5MVt3udIY/EspmUE87mQKN4OBN1HG/wD5quNdmAdTqYc8xNsd2egzRn8zBxZ
NrrDLIOR/OXs94fh5n/3XOQr8/ypNAdAxFSM0naeScoea9dNSHY66AQMA5ysA/eZGjULHUvDgcz7
4+gP98JcSLFNkOufaG3F5xlSxP6m19aKvwX43ZeuVg0bYlyM9wwJAqA9VsPn4Nghvzk5GBAFaNRu
FEmAW5jEdPmvlii+g4LYpHuNrWQQCWpYIzxm/oaod8vRdKYkxc7vYdTdsHE7hIq0Hw36P8Fp+lGC
4lv0EPAyim7a8xtSRAcx9IWuXyAM4Nmk8NpRuz0ZSSX7qAODgBYd2V+OMFrbrrxXJpwiBAHeLKeD
k5C4INZdihjlF7DnAN5MSeLLhD8+005s1AW8OjB8NvQIamQPLDcgphNUhN2+T4TG7lCzW9DqhZUk
B7Zs/wZ4VDxPQLrOfvaXL8BHq6nVlPbsqx6jhrMaKWzsYTAKyIgIZPMpXSiy6EffZpwtDiuJyznn
25wNvyH8msqMGrp6VAoTmmMmqmZis4w3/7PjarskeVQjvQ+WxQBxtOEX0rBic1XhqNErq+xPGgFh
P2EzCRVjZxTmT+9X1DQW/Aj5ePoLGxnYSKmu6j/0BT7LMT6so8mBDU/34O+Gc7IvwHvxn9FYPZdl
sHrXyzq4AUzmOGdCPwXl5Y4918G1lEAzCAnO8dCrcjlRKCMaNBbrudZBSPwD3onaOaPHlyi8QwjU
7wkHv3NXyku3fkcigeOSTPsa48VMzIJzmr2HCRKoMQaiDQXrVw58eMGmDjHu8UDP8VkWIGX3tHGn
YruhSzXB+6o88teXvP1wdQ0aZTzY6mivki8m1Pz+syRkTfnHY2m21OpjGyomO6+HJx8cR6LNiPIE
3nH5MtTUUyOfda+WwZjC36ouOX/Fj+u+UzVado9LhCvAiARB2BaoWK8ccszDm9/nQFT9MtUxCSdv
BYG/UPwYgqe7bTQh32KTZux2WxCjF1w0h7aW23wRyXbGGyGIXp47R/EBWLn5A9xgYGptTUbD6XXG
v0w9DYdL+/fq8nE+MALNwtJfkroEzL+n6il5+QXafPx+CGA8D0991rflzeIcqxCyyJFAr5fONiaf
baTnd5+FtWY079vU+8+0tKlB6l/jlLzC8z2IH+INCOT3+MS3cIUr/pd2HRmr0vo0HrFlE7xJ5zKF
xdSQYyJFRVq7HISCWPnz6Iq8QZqXAcMp5Z/Pb0wBkDRBw3hcxqt5UotJv2QdxyC2muAkMPNOcOQF
3Ih6Oc+DV89IwsVFfgV+ugLP7I8feUYIC3hgSGFCvKilr/4TV/ifrYE96zBuO9eEq0NBNB1wj/qS
xKN+TXHm/eMiAMzVQS6gPI8CJ9iVxidyr5c0F0228WAPKCo7BEqhh9+BxiOQqOn965uJIGu2dtLq
rSCAXspSYlOvGYbB8uWO+CHplrDGKzQ+f/xZRdBuN2i98nANTW02UPfKOiQgqgu5lwga5F8sieEh
bEZ309ojcXfHvleprIkR3OnOMItEtrlY4z9lOWbcgAwXRuQo+hNQ4vzH3lrbRt5CATgGWH+BBSm5
hom06Zpc5F/JeVYJtKOtWF9AtgFNNApCQ5hp19Z9qO0E+fdY+GfH3V3MMUT6O/WcQShrlQN8fPMW
3uDJXeb4qdDamUYr/ft6B7nS0MDemJsDqh60TfJjGzxqAeD84owTLu/C4553UV/MYDnTv8UVN+lm
KBLK+PwceOjI4T/Z0EzuOpHdQORcBtohw0zsyuP5O1aqkW83FNvbbR06dVjUiroLfLWw5xl14vc7
L6hAWMTmmGVCyJfjqEVuXHZqt45n3jg8mUC5HM+e6YV0jk1zVk9Q3pkgblhC/x2WKsmDvRO1vp5n
tQHsrfPdYjrnV/i1X8ITEsKKJArUhk+TmRHcBsQSjDUKthMpS3dExMEZAHM5qk561m6wWtAuuzX6
Ps4WLsqVR0twHuiXLgZsaX9xG+9KCZLDyhoM+WWtFFkamEYOubVcIIPH5krwncirNNWAxwrDH3Vw
iXPXOzmaVkCJaJalE+pEKR1AP9ADfPoJxS9Rc3PIstg2tUyXYyiwDyMT45LNsyEwnrUcqrhHc03p
rQEKx9O/qAHbDZOECOvlD8BbVZKiKHMImNm6/Vr4IMD53woGfZ85fSLztLOyw8D3vxPDhyVpPytS
+H7EgnxjN2bOhPvzbXEmxnQXu8AXI7Jqpz9DypcwT3TWnOLKWXvf9Ld5fKJ92+WfCoqHQLBlN4rA
NMgIOyaMI4cyQpn4LbseTiYgo5M+jUrYqymgyneTqofVTssuz1K3oifWr1xbqiBekXUetH1pZ9Fi
WZ4LLb/DhYNsEmmOqvO0ZgjX1prPAju0OCiHLUjkdSbNoE5PuEINPAzW7pI8+9lYZFCa5NY3DtKt
3bHYwEquu2Vjqi+hlIXTan9prkWxlKeyPraDx8f1DYif/DZKS2SjV3Bqnj0K+CmuMqwzHTKYGdfB
nP2AwJ1q0E19qosbJTorgz8mGPUSQqTExI019B+j+CzKrjELFp79BTd0rlKZK5s3p8PncjkbwoiP
xdHv0pniCHWb+R0lm9ElMwkUwTwnrwLO+251ZoRAcH7/RVokbjGojy2UrlwJ5J/Uv5Serbvd+4AB
TUZbV9nfp7fKj0makGXg9OTnErXTCpBuzyqdgYBgBpzu6UJcuSoy2JfGig/38Q59L0qQ9lhsS20d
k0saRwQwj/eTii1MtrbEaC5AkX/c6Jf7cgtk+KHxN4Yh/YaeuhcpoF0KBsyWkUoaTi0A7a4lOTuI
jEaeyKyohAzDUBK8BMJCtoi8MQ/Eh7q2yYnUb9EzZxy1YHVSJ5G81l1YKH+dOU00ZXj6MzmH8ceY
C6aMNxNfmI8MhcWD4vybuYiKZTP6AOd7lpwrhaVrT0Os/pgDtEt4pzh3GYT2pUJMJG4TUzGnUNmP
ub74oYKgdjjEJvAIePCSwnMlnzZCHfuhC0ysTLaHE7Ud04IgxXcs0PAJYRoQiGp7AMEiKpcfDCkH
t3QoFtnYSK5fS6J3h03rh4q0dy0Fzcm/8XLA5gsyNsQz9f+mpXglMOnHaDKoZPhIu66Xb7Vkxr5c
KjQpwHlj3OvjbhdIE1NcK0GUnl6lpoMvaYsA01Yzf7rwdc2dggEUjblEEX1zvz7aYBZcBoXtM2ch
WRQSgggPeJd6gdzm8Yt93mFDpL/M/t6Ouj/R59tlT9C5B54ZwxL1jLIRjeEm5mK6b2xzlWRXc5kQ
fhDc/hN5WWjSMxqIwEZTfvtBF0tJwyhDzg5pgpFm6EDlZAA8TNNbLdtTrAsFs3J6lpi5JgR3eRFx
+GO3+Wxx+Hlx9/WqBkatzh83AuISjUYq2ZjLPN9ROc/+y0C7iQVIHJzt/xud5rgLVI/40XURhxf8
Udoq3zi9B+I2ZK6oRyTiC7VNLpr/H6fuWSBxVmHs8sl4bAQuaAY9Df00FTki6PQ9VkggjFhiC5/d
SK+l+jciDYfjceiCJ0yY72fOCKNfE1X8C29MRMnrRxZ9G0rHG3snkFQ0g5bBlHil1ZDzYxGZNkGZ
bKR6sZYAI9v7X8NC3Vw0WhyGVVdrp0TceGHbwKSgvfCmLVsZ/Y+u7ggexLqR43k/WZVxtOQNON1e
0J4awpAkOtLl354CeeHxljhE9Eqv0g1kQV/cQLTjn3b40DCkbaTF1jHFG/URbPZ87H/jOV5xbqEw
HWVYopk7pKGCDTgi+QRqTEFmf6/kdCDKhwnoldlWyRycMogmEzT8K/6Jh14YeziexOs75LIQTeKb
asWcueXGlK7LWLamNJ5n6XOF8inLrk0GecI7exOUdx8AAm339R0wZ64gNO17MaAlTdfk0Xd4R1VN
bh8/gHYVS+5PAa8QYPGFltj/sZ5uSBUQQD9M5pMmj6vJcuMmcwqsPzTOWEMsV2tuECKk43nS0UGk
/HsTuudqWYXqwasR4MkUCb+7aUeaxoRD8iPkoR0Pi6eOSABv4s4KQML2sDYdNTLKq9PfF3I6RiYX
9W+QyTUAd0Oo13Nt3JA2ZtG8aoiIo0IA3Q8QN2AM+4/Uidx3hC/jSxAh3CeNauGd7KZWFS5rj9Av
lYtS3omqlYVf9m1OfTg+BkZSzNWtwzy28tmZfUIxmsM/Lodm+mEuKWTRfKt0tOGpOzxF6Ky+KEUu
6ssOt+QPwbCZpgexFVxCbI+/NN+sJX8i2tD0Cka6z59qbm0WdvNdL5UlHkwrnca0DDab+R9zPnZ0
AN/EkZ3EP2skjpZiNluKw5CXolIs3pHcE9S2qOokfbbzfVx2TYjcPoXIcQY9xLwPc/igGXEJDhVe
3pPqVINPCGHperVXBNFWlBnEyUZNfyZjXBLx2MGJR6F/IXam43mN3ZWUtKe5WYXdCyJxaHe0v0D9
rAvIRw5EWE9p836dRIsrlwE+jvtsyVCCbt5opNRCsZT5XKNxuyVar3Bwk08tNvHLJde75Kjlf/nf
/UrmPN90VG0aYlpHcb+KhU//xpBBW45LpPtqhhyEF1/5AbEUkYH/qQWogESNYL5nMdU0zyNLbUJv
d/r4LO4j0CY0ToP6sEQckRs0WHSq4EORBoszUM2ri7D2yaoIe+VmQ2T8sW8+Z4tKRZPCFttkjq2s
L+su7ZZcuRCZG1Kklr0NQ2Ite0i2ucj/Y4T7dp8RUJJhejTNBMN97bjmm7L7kZEiHz0UKwhXKx5X
j2B1iWxYYUOTjmBYM33R1if6HFI42a3No1ZjJV91ZqYu10NcS+j6bZCQ5TIRV12/O6xncq91GDFl
rGmSjAI5gaOSiyHkoajoh9O69DLBD/0aVB1e8Px3X/SKt16xzgmQcP3fgjpSpftrh4pvzq/aQ3Al
DHh7lH8KxXCB3pzYsBHhkTlv/Pdh4jqNvGn5gcdoJf4Nqf9/oF/7Qqs2VBbP/3CrJSwManYMLEvl
w/m+XqPGF5lgBRrd/d006ZawB3Fypf1TLqfUmbaT9qopuhNVA6/8W4skcQF21lXlUUQ3A4vkSg21
XAHW2+8LyUHRYf0mfhNDDkxACfviit9+M6ZowHjFnbZpycux8bS3meRoQTb4/alVksNW3dG6exQX
ri8mIkjgHcrT078O5tjwSay9fYieuvDgfSMu5qggVFo2a+/sJ5ndVriTm8iEmF/I4eQTaIQhx6+I
N82Qld4f6hr/C9yCShAR/ixGkC1b6ydJQp2CHtxgpRwY4w5zyYc4+yNw6be8FrBVcp+mtg21u/Ii
0MtRgMv9S/8T2X3rMWqn/4/GVPVAO7ZYyiWLd4RCqy4lb35yGoL/Z6OjfbNpIh6QuMe3dIMJKjri
rXvxKw07REC3sDdAJv6YOcxtDIJjDX/WpaoC5rIDZuuCH0xIARVlMKpXpx1/X9zEy3iKKPg7LnuM
rZSr44JOjksiJSd65Uud0QcnPZGsnNSCatpPweSLppJygxqckuysTpUEhu3djlHu+iTShkcJjbgH
YgElBMFEBxhbmypUkvsI74bhbcd8x8IGgxuA40dWmUIrv6z8XpEvDPv3YwwFmcjJOvxnu95s6b6Y
3rNG7OAS7gUv5PL7EfFd0jPb7ZUywC+kEcR2J1zXrvlHQwLrzI8tUj0qGAGOh8irF4EVOLW2QLdK
bVE9OGCp43lglblWSEuL3APp/gOP6Xpvqf3X+48zEjRBkUq9ibdCPb7frhqDBRLPn3QEm8UKdFjD
1c4Wm4vKYHylPujRkhgn8yMov+zhGrI1PutLLs/I7+fKFDFpMVWMxsT6WMiB9HrMFB8fLz+O9yg8
i4k4eZgFxqoGiCEz+kXzABJ320jbNoWTAWP8Nik87nZy+odfrAbPDLDCRwgb/FHD6pbRZSnd2Q2p
VAXkOagXoJk/NW1HMMHdsQFrBH1QoGleY68XLDiMgKJFsj8Zj0RC/HcHNeypgPntU37kS2IdMrPA
HAtdP8z7G4JK3B7Z4s1jFZvGWpUBWFmVXhPi0gZat2AAOrpgkme+9f/msLVpxG6a8n8aCTLEQNEq
t3H2F8nKKn78eEhBDav2L7uJeH1JHBZwb6xfKV9V0K8HjtvzCGS6G2yMlpRT5XrLe0EsbTsJ6HoO
Ak1LH7JQwsz+s8VbGdz7VFIU1e/0BIfNesNc/Vqg/E4mq/JIQSaUw/EkRaYJNSSahZgaIwYJougr
taaYrrJ7Md3f6jH7p7U3g29HqN8L9Xpj5QZ1KrkTjQFxtFL882u+EuRcV0EFtIoU+EbNfHJcxlSE
glbnMiq8JMd+023H05hhafGRbEHTIcsFYCfC8wHZ1g/e++eTcKjXJRNfSeDMKzwkCVPiNLV6nno7
BPTvVqSod7OsE1RuBYBqQMDtX36yjzkYZ3SgeHlJffxBhLoBkZpDk+vOiHpvj50oYKCAYXmPJ0vC
9vk8mAcsPHtO39hrXOkpdyKKw5bbLRNuTEEol0S+Jc1m5qW+MR9NapMvW79Siq7wyw6aH7mXKDDN
MVuKjnJfl97uBBf7muGTAQd0sxYinyPF7SdW51xkrT96CWJ+fMA5bJ/qdvsADj277JE5jLo/6HFj
aFfJl6eFhFZ19tc8XUVAQ9L98UMYEaRh3eXuEVUiGVkhT3steQaoTQ/HyRUpIE5qVsP4Q3IsBNeZ
0o+Cv4Yh1GdlA1xI+yIPo2nRNlcMwxuXgiUdij1nszMwit/yWY0/assvPFnjJhzWIrS0nLDP3A2y
yG5pjWWsi03Ed0+ycBLINRLFJq5g82f6PDbtFRTkXAfw4K2zmERYD+IyOZaVA5v50pvkhUYCCkwG
ys+EdLT1DFiAfFfO+u2vNq9P+5z2a+sevKGiUu4qS3EJ6kkroOQkO9RwEK77QI+LKWTwl2aGNUy2
4qQ8+bf2eW3xtOCKMzQ1nYuaYZB3JktwWlvU+5czFmM1bb/slBgqiaXBNDfemCkj7CeaMLcWRwIz
I5Nj+lW1b1Cp1+pyFPiDsNUqGL4r68/44dR5EMttseS4sP46N8GIwM2CNurcA5EbW9SxoE+Zw7kR
nMpR00tXl1v9QqAHGnOgzuJCuX3aaeC6UmNnqrkiCsSsTRswAeyasjYF7zOzmrnz6qS4wOqbQiCZ
cMFm/cA0ICo0kxrqBxwZy9vLVzhAav8IG0dW+2NBTag+nVjrzi0+hX7f4hUSCr6A1lcxy1KjLNS+
4WX+3Xd2Df9ngTylLKNM86dESi56B7CJqavQ/6u7nVYq6QkSMiTfQzGgnMkveggAocYmsxLUlU1I
i/+rl8sJz9RNoYE7yGLdjLTbnayOt9uBuNSbNK20J6r7uK0KcoSAtOEF8Zv1Rgm8pVKsBRUumEu8
eP137J5r/vOSwEAODKnpMn6SdDGNJbXUVcx5UNBqgBIdSCxKFDGtH+3QDpi9iK1EHNJjyh+D6/es
+2ntE0a8psdPwR5VxvRg9PdpthWZj1R6oWpjynS+ZWKBgkaXlTzGRhPnmRevBXUcbsyp1Fw98Gww
98t8I/AHylGneB5DWpe8xlmMAZ9vNtycUhFPN4XbVWQAtT7NDH0cYPsHyvQPzzkjp44nYnH0dymj
7yjoXxJ80kUD6l3LVxTqhnHmHOJvxgJxtosN7Qqa8w9+ZnYwLPoB1/CSRH6SCo+V+ghVEdlqyGYP
zHQds712GS/48XDKqclOhnEiSSa/QomljLcA9opCMidacm70RiGjK0rV6VcGwvoFem2D11DuiJmh
WZkN3tBE+z4N4y9p2/ik4alBrYZAmef9v7R0WCMzyPBhp6nWeuIdMcX9XL7cpi3NrLnvvTbIIeNm
PGZfrgiuZaZ3XdpwK0tVt5skBovkycSlNYtWxzHPZJuMI2BhnoCnZhfoMyGn5ukK4gcqwlDyF7r0
NJ4aeOhQubLBsLocDj+FecPcCFnm2JOJuYVuoTIuyEG6L810h8RRS8WSeR2cX5VyeRVAPBpUYtBF
d4cdPs0Fw4CSp3FQMAl0odiccWAdR05m8A3+YKhicpxWGJiWKfkMKXzPFXYfDBMJ4TFIuBD5xkos
FBdEuNqLUd4N8R1/oGrWYPiy7utQe+5PzptTVDeoL24frHpbZhl9sTaYLKo+A9K0Nf1jBXzO1Y9Q
nHoRxuFhAcUuzhWUmP+aMa9tmEukU7dUYNkKtp/nggkHP7eCq1mNeW7Dr2zY9gy/V8lhsY25Lu0z
JVAYAUl0OL01MYiO79814j3kKnTVFSFUfO9EnjZgB91MRItnm6hDL9gWZOO7J9qJw/KyMbPl4ZcH
2he+OSAtwpxfdbHWo3Cqg15KHoQDbPAPSOnoUma2JrHGRCOvWt860NkCsINxHd3uprvK/idvq5tM
egu9blScl1YtV+vl3tdbEsKwXfWwlrNZxBQAlHG7u6MYNZm44DfmVHgXY5c/src7JYti/Iqk0VHB
XSbFGWnvVK6Od0n1FPw/pt9jIg6Aggtgv3vOPGPkkAUWTMdM4w6sDVp1qjNl4SvWtdD9wT6ubhym
2qmIvqRAo/BRkyZU2ttFxt6YTWRDKPEnLCcR1+kxAvreoJ+9apAca+U7wD8Km+GAHMU+KhLxugWG
3WAxrnEwOKsH4DgNxoC5J93piIQCCpA+av4FI8AYUDqkufuOfs0DSyDVkogSILLgvQwXvsiHRncL
wVCBZoy4aKSGCRQj4FMTlE+LslzqFRWCd8G7iGUJlxVmvDvRGEhANi18UP2GSp0LJJYMIJDK7/de
Dr//K5im637yzoB2rALSGUMB9xHMBprpbBlxFIIF+1wpyfmG+DEdZ70jofxzYvi3c2avXCo4rv4P
l6g6uB84eMnLB6EB0MuFbHAxbnd9Xjz7c5kWBhFDXwT67JYAje5jsNI70gwPaColY6d1kbUOXtiM
xirvBlsoc8g13ECcULT+6ZyF/i18HVl2MGj5JDoRZfJCZkZ2WrvyMYVM59ncVTcPH2MvbN/aWG6c
pFSbG2rAiJPz2Z41/qVB+zIuuzfFiB9C0SWdmqs2W2fQActH90g1UXmPtW1/JlcdGFx2tSx5cfr7
ElzYs/JgAVL7N8eausF3SYEGOVZzO6u3ULNtsORe8B4ZKq634GOvJY701AdM6dnoDyOEYSuFoIye
1EgZvMe1OQ3WV27ZTtbCwQn3NO7pzPlXQ5Aut3DJLVEQgF+bc2lzAqYpCR8vaDZ640b+9y5FK4Il
DdzGzG283BmU8xUKS2gGSzlSBCY8QMKCAH3P5gCY/abkn3C5XZrSb60+QH1GQRS1kbyxSPIA4d8K
H7LySjKP64g4YAMm53ecXMd7aqbNbeXQERcVZH1JlXjRPHSAMIdluB9ez1gIjEeNq7mP87MGSW2m
tWeWvJBU3nF+GBoz7qCzg+aaGC0fs3tMGGC492tG1RSw5r+VLIvwM4cg5GMMLzcT3QGSNK6YhNCW
D0uIKuJSzVlGsLBdH1aQKLqOz0xdTpT1kRSuXj8U6mROm0aAGCNzKN3QERtDrdw2PbdU7SsFRNZ2
PdeuHKrMWQsPT1ftc8DA8VfJGgG+TYZKjNoXETMACj2UwPEcCcrckPMrydCKCk5k3RfXTezAGl5h
mNDSuUI6j2Wgm1rg96Ox0sq+wUB9pa5fNEf+nlAyABBy9NWV9jU9rgxOZj/WzyhqzYGJK4GWVLX9
H4mCP+BTkvVq9RudzXw3YWStm3K9jT4Pae7UkinZGJyZaYDPySLIOP3wYqVxacYaC18GfNPGs7SN
auVuO8QV4DC/IkOxR1O5JHUL63TmXMDdGsriVC+6nrEUG+gd9ApYPPMNHoVWpgz/aHIYJzhip4Du
eiUTAHZnCaYPMO6hNUYOPimCk5YLKuB9RiGfA119hb0uNqvHQqi78OJCfSbeKR91GPSrUkvT2PiO
CLqCyTkUCEfEX+eHF3DPHiyEMTlf65R87/pifzNL6Sh0n3qe7aJ66NBiEY5pELfsO+niJGYz6uMG
LI88l4Ar2lZNa6tdoKtQIXG1Y8d6ZR7eBxAP0YdXjoPydaQ14AZZNoFIdaNAwMxpCXxlIBwavHiz
l6mCASjgrcvaYB+EXrBzxfwyxWE5zx2/wpF7NHNzQ0tVWwQuW2qoy6Nb/tOnjfCxo3JHpqnftIRX
UoYHgdKw6Kn4WdiOPOfCOg7nC0JRtuqCCDlg/KQ0+FiLVkMseLSf+wqeAdFMAgqZON0qQQxIjJia
YJrZJTadTIO/GL4xH4SihCU1k65ltn7jHmwe1/0xKzxmRvivNPmgSMCx8zU16D9dejgnZpa6Fs6h
V80sdWXaRSaLJoWH5+Wljg62YjPgLzHnkUuZ1JIAUM4nz7tEDIkbWYx91mcuaFjmYz8TdMXyJr9B
lGbpveoqz61B7mkk0D2UW6k+LPp7yXczlLoiP/xLmq3VDcnY33Jj26gTOZ8SrHWyGjmrhyp7SGpI
UOWw8z0A7hpzgIDlhmkBiNIbZ3txcXqh1v2tWQO0p8dYFfqSfGVxecnfx0ckoIIAO2Ot7QdJfcDi
3nBiXntwIZ4aA/hSRyrHd8fLzvIBSjU5hhRmFvy/Eic33/4QMWYurm0Xj/UO4e6LGlUOWv1oT+33
N3KudH0C7mFJ5913UiAThsTlfPVYuaQsKpKAnNdUsQODOGMtSpIU7phfX/dNJ/KTXrm/rFBX/6T9
Xsoo6Vk0ar/Lqn46xJqB0eq8W7VFiMw93D9SrKroJWdCEaV5JfVuY5weMzuMhdWHJFJ/21hUdvvz
NCQSmCIAqGdXJn2k6X2NwfLnkCO9HzUKX+0u9u8JcpZaTNY9vhQs/gEGV4jbS2HP7WPLXsWPJdrb
r6H/e5S6lBOWyiI3I2TLX1DssxevS3hYV/FMdBR6LlcQo7aqqZMfpLyIGR9qJz34qWzi1r23CwU7
8i7nJ73RW5brr9biAIbeUWESxyTdnKcG7QXQGUAGvxGu0OPcZe52cLE3qjx/pKbFzI0oIWKS7EWn
D/YMPdoKF9Jh33T1PLj2FNzWAC6Xn63XtcEQlT9yd5sHpv7ALt0hMmuwoa/rjJigxHLkIH4/A7h2
nGUB4CEC7Lug90AGRNf/nUw3mFlIvW+oSp+rv1EfFI9eHzFH7ojHD52vr0ZvmTsT69eBOm/C4adv
OEUWefTnHHaVDUReoDU8c2Qni3zBG50A4EUQnj+nFcZpgLX6EOQKDjdgGID1cgqI0clbxld2VKjy
R8rqBkc/te32RS+zsZbduWE1mbbqFBeAQIip4gOj967kEp4LvqbJT3CUShE4vSUUTXqYQcSqqdCT
BZcNbIHXaUFc5pPJl2mUAM2cNTW3snQziZphXVTndWto4PcFECmgipgukzcZMxfJ7E1nq/JTg+UV
Prq/hOaX7dZLWE0+FRwsES9/hKQ6Pe2iyDEeswyFgINosL/ffOtGHXsW8dDxdLwbpKuXlaRa77nj
h/ViNEn7BHIkmqIhw3oPgQzACwR1Cxf31EqGaTg0AAgxO5NtD+mnBacvMFd3W+oGoyFgnGlJrIgi
T9XmXFVh043rsehpFsWdL3sus5F7SuRBPeCpO2Vcnwx/qWzW3W38a/Fm1f/vLQtL5kqx9mjxVjcO
Plt+OFbf3HIDWPxOk6MwX0GNZcNUS5+FF4hW4Tu//PXYRSBuSz0TxLgPA5pFviWqvDz+kqpIUrgP
Z3lKoePTnXwmkpubJDftwocRAwE8XA2X2QSJjy7yM06LOr3FXVxuXeuPDGMJWygwYRFW3qozLxIu
I9klZbxotXHvbBvJoOCqSouAdBZQwhBoSw0DyCXxUdisYHy75gCqimr0US2bOS7iFxVobW5/sXfm
ihskBvylpSmahQ57+wloZZOaF5niKgeKtW+gDk/waBg49uDV019xEUg6Vy0YF7C+utQHX+WQebg1
AinnExSvdoNSCh3IDsHx9UCSPaWns82RfI9tBYyyZ0NTvDJo6qv75gVEAnz16QkYtzRZ+fzbRnt9
k2jIMwX4jC/uiYT/yCmGjsNTjTwv5XKQllJylc9m7RiJYjOQe+4BFZV885uJJeSg9A4XGoekFiV7
6ofCGiC5lyhWUp8CX6SA2f8SQZfSOM1RF5r+YOgZrtitmiqRyqxlGC7AsSCEU4AxSuaqB1ysOVAW
qICopnoVVz9G/RDBmlaPSewZ28F+B+Hjd715GPC46J0BrdfdQ7FDbKcTYs9ZO21aRZ6rqzRKyOxN
tgMDkSh05Lw8cR8AVKqxMP1YGqra523bZ8ZoeVaRb++wm7bB60+xkWdCO08ky0Lz+yp+pNz2plW6
j9QiH2sADRUcoj5MjSjiDfCdNnNpQztuHD+SC/QIdE+w00QPEPvGkeOdwOFGndiygLQVxkFo4IqZ
lvJsulwiLGx2Kj4u8NXar7HJz0KepBVaHrQfuZFpOwf8wONf5PLEeG9mAFBwXyDkwReXcgkW9Kfa
ugfVx/VxSDmCBYa7/7IIYElVDJmDnLmLq0NeiAX1TzX24yNZGLoPLfG+ZDKrDpT5K58YQE5RAOGM
7ioqArGYLtRAGlaAdYUA3AoLt3nKZnOakFt2GGv/ldV7D0qGk/oUsCf1opwJD0GUR9+Bmnl/lFfm
GqppIgP05ehrbgaTPSze1oCeeFI9XHpvy7LROnFgMep8nsvpShpbn2CxXvuizkG1ZYDU/k1ANAxg
QD3AT6JQaXIowBzzAiRgiz+/gaLYY6yChmAvnaIDX4yqvE6Sp1dZzi0tOOHrelIwcPZB7AmHST9e
f1G0Ju9oqiHDYCfG4tIfrO2axEWXWpvzFzJ5KCUnc2nHDlYpv8ifqEZ2Enk2UlNljUiWSVyWJjIN
NwwbVus+F4G8c47j/W43NgouCUk4/+eN5FLpsjEHrU+Zd5PI0coqxff1OIDXXBAy+4zr3GFGMCcd
Aon8eDIP4NF/UXWEfdV+W1cVsNfnMkbx2P/qjsS5UK3DYlhOmF2nuU3ambaXLMT8lXKejQMwa1oA
yfCFGfKuMHKyRH2f1XCKHe8TBYP7dKP9jVMCVjwkUgOvwZHStOaadqFV8CPPR661OaW+dgxKDZK3
3nJUgslPX9Hrnj5KrMhPETDpMivJXUprpPZwOepj2LPWR7Zz0eEwdlZdxAg+O48LiNhNKg70k8Kf
/vpFlcmlolbxlfM6z/bnlRqj/Be9ifRHoRtA4pzWNKbAVsGZdY4QuZHjkA5nuPMGhrDWmONJaZ4Y
T5q6hiPgCIIgOuL8zCDxZAlmH9AM5VG6R7bHWxpwH3/yOr06WlyDFVp33SYEvgB4cuXbfAqwtC1J
uXilRoYp3xCMv+v5Ql6JDbjzDuuhM9b8kGecmHP+EmREWEs4FAlNH9IJJnDG+DuwB4gkS4LHbcyw
YL0jP2EVTS8etepfSyRsPDkucx6KWR1kkM/LxjxlZJ2KifADwMa5PbtGjzg0w3raoYXsjjIHvOAi
5tvCYRx7FCgmXIgBIksZh77QRL/dCLa3DxVmWGLlXf+WKfX1bQOgHMyKWAGK2wT7WSvFrSJY62os
LyRw5dSQOd5xxgGSs/39eZpc9mCPS5c7I7/8GwkdZSPYmP7hP9/3nJp7XCi23KNKvASkOSwdD9dk
UB5dVc1medju6aAy0qE/llQFf4IWeGlc4MMSfjhRbJmM1mct8A2vOlGCjxPoEltwWP12ATMlwj7m
Rethia3MKXsL7J9friQdxEs/hHZ3aeEEFKwTEun9LtlhJo87XSw4VrRXH7KvHcPr75zq3b27+WmT
TE4EZNFsm8Q2aDP2NTvD43sCnQK+bEe2dVy26wjtNe/lw+AUYz7PSotw6w+liVwop+r4j3eV0U7f
0cSEax/J5nEhfV8lT2GFS/FuqseUzRT52nAL7EHzCrb5igkzXcd/Sk0fLOAIrWpQXu7st6ARA8ev
6za+S6vmDP7pcIAOEiZbX9iMSW/g3rkx1DKWjc+6JSydZhE8xdZlPL3QHLkipuTsvv3wb7+lhgFB
ZzMK2pUS3li5awicDJYNkvnxtisKLBsSjmhwmOifxIjS+lz56GCm0F99aDImsCI10mAvAXKZ90IV
7JCvEWuzW1HEGBYqO6GJWu4kbuj3ZeCskXpdwZmw9mp4qiqzqX07fbOgwzilAUpcOmlphiBMEXCq
EWLZKfboayDMwuzJV122c6KaFwl7O1iN3BmTtjH7xl45Ku95Nc84ijv5RZ2r/jJO7xdOzxcdYCCw
6tCTKD4lbGTUNiWd3S0AMOsU6NVJg+K5IsT8+N4LwAvYqU/A/FBGHKnJRNYU8VSAmksbzVLNDafg
OTMLsCzdO05vSkLp5QpcNykEMtDS1BkfykSujoJ5QeUGRu6qnZUfIp7vGU5BIIvzKndVTDW1akVo
rVx3FUVtEiYd+4RcCPgzKmFwxV6HAH6fSsbrZmdcaabSTNqE3rX7wlKwu12RSlRO1VEuMMFGxHul
TMFmlUiS3TM5rs5mYvbAFWmqFTvGXaxaN5JcIWpxPW2epam3d2O9h/AoRgogGsdHYVZZ38Mzez6T
JCFVrmeuycqgo4a8IFH+g5EzkWg9mEjv0a/Zy+aAF/skKBmQGBlQeiRgESrHN3WvqYjqMbcUBRf6
nbK9X502BbycxEWUVlUG+JeNz4aJnYyWbnI7+5Rk7k0FHPYiWTw9k4DQTeDlRrP7l2kew1EKDKco
o00IE3oA8DSqt3aDA/7aU/kvnFL2ERQUX9n3JakEPQgjfPpMmwaEfer5C/fMj5iN2f89pPujeN9N
buyg2lBD/GseDtZcDmAGJGq1Yft8sh50TppfQVxx0WUU7iTEAbdaPYa5w7WIUDn1jWqWH4Qdf32s
LgnPeUe+TZHLkuNcpqqqwE/WxIAcdOdpZxorXaj7wnlvE7y9n3VqEsfESCiMMqSVKlcNYvBApztE
fGO/2qUh96zQIU4uVEDzlfSTwp0P61VP8V7w0gTc+wC3KwgTkoUMX+4LO3ns5hPN1krZgRVyj2RN
M79JO4FNWsdssrzpBLErpnWI7DzqG0sbs0unpRW6RgQBxhhmJk7j5crtTDwENVaO46s/xgQkwUo/
GhWoU83QQigbS9AigEsFjf2wAYGPPSdMddI6vyycpldyiVL6jCx+otwRBUANjqQRt7BBQexfi0my
T1MEI67BsXpsvzFoFWBUeGxayIgYAnF0F1uqqtwCKW4Gn0x/1zGGiqkMJ1NlgWuzwY7wdDAECve3
ii8zNGHukCzykE6m9wYbNMYDz4/DvJHp8BtOaAxDQ1V1dM94w3Z6cEDPxrQSh5UBUSVIriB0y1kq
UDZ4svRRtX2u0Sy6w/ZDIxUe6VEznDp6kj8YChWVl44e5caXuBDtA0rTw9UNm2/l9pEum9tQ42cU
c3r21y/rpjI/I1GpEBbaSBwL6eTvuxKKWV2Pm8ehR3S4fSIi0EtcDRNnklMI6R3ZxJO8W9C6myFa
KgqOkHI+a6n0drNrwEV/spCqtF5Gzfxu0n0YREnWOz6VVg4AwnzXGfDj224ZV0yxyIN+0nWJdRMJ
juhTfd/KMi2get/YVGBodjxEhB7PTDGQisKsihP26E0f0Dk/7tfkvAWwHt1q0f0s0cNrRAOcZ+/Y
KVWw/Xe4mr+Opz7r5vddQ2yd03EcRXtJksJcj2FZ+QEho10OFCf+96ZgYjP6uEt78HUfqUcPbe1c
TCIgp6h1Z94PygI3n5RuSqBEZNdj3N1C2fImJkWd26cy7EhUTKt5Ns81x4k564Q8bxEfM7GN/uji
LFiql/ibHFDn48LW5SsU4La2buI35pdUEDtMCSpsiZQN8wpU6ZcvRn78PLaIgxVP4hRuy/gonfBJ
lU0rp+iJhUISDr30rjaqswW6ThikXdCYu/im9W7J5giWH9aiXCcfENKsPew0G46FkBh2JNuF6syr
1xLPhvGhgviKw/AaWohxwJ3CexBkACGhOKxrSNcpNsqo2bXpuoCRMTqzip4pFvb/odzQxKVj6DD6
QaHaR4VKt94LXEDsajeeVK3eWbmtgdVAK1SJpAGExbesBjiq3JgCGGOtPOQEaRYp9xkC8xuV9bBW
dgLCDqPS3drm2IaRmmE1+zqbFAFbGCXS3ZQ/wehe/z97ATKIlcgtA4wFrQrinOfxehYt4Mmd1Djr
Y3FEWh/O7vnbrxMuLa5BKRaGRijoZsi1r8CHQ5jalS3BRD6SooC9eedyC52qY4aXaPir5hER73Ga
a4rgyrvrVZS3RUfX/vsP/an/FsTYdASR1DHfREGOLX1EoYEond4AxmsjnAzpeR9vZ0Zn9GILH0k7
j7O9J+lp5ERDDv5omYjM+5tFtc7k0Ox/FzZ1FaGgIPNdgKUFxLIK+XXgBfzbPEUN72V+Zjapot/O
5J4Cs88zY9+SV0lYtXrBwXz2YLYyhrtzBhgkBH29DoS3e6FhWaXeOUjA+G/p2UplpGGudg8DFWrJ
dXTdOWYTaeX+5qEw+z+ss7gIYQYYeT1UkYWsenL55x1BHdL/Fap8sAq00zXNJREaEJMHCTvxKiql
t/tV7VCjTOliY1OM7NiGFcEkPwf8JprsM2YxesJ9IcJAa1ezI9rklR4aWruLV6cr/vYob6jZyez9
AYXqDlSzwXW8q6hjAWWzjzGS32m7Th05LUJIpmLouq5mO6zD7VQ0ZtvEbKdXmbTus854VtRGWdwr
lvLvgFTxlMjlguMSOjTI8H+uz3X7NZE/o0XKIcFdpgp+cpI4FzrZJlypsZ7/cBNFNdrGg2XSEa1V
sV+kNLpB+TP/B8sbHwcNOPfZlZ1ADUFUEQXdE8V4bBSPI50u8Hwv/ETnLXHb+TISy7i0RY1F3aMp
iey2aOufIIN2jy+8wNpldEbb3CUct2PuRL5t8J7F9oacJ4cfxiHRGA4HrnMMEv7BlkNO2Syg53xa
pCoj5wjHeOtt4CQ224Yi2DQ+DjMv0YBVuVcINi0lvJwbRCYW9kt/8QqmjVlSio62IJZpazvxiGIr
XzqeUJq9UresE8OanIWlI1Qrk0ckikbHoSjxPc01BPtbs81JApsKlzs2eIwmgs558dFLSQ0Mv1cw
1thZdNEG5siKeiHK4RUb97O2Bltc8DwHVLOahhK0o+UtS8JyU0bgyJNmHVTskgwaK31fik42z0Oy
MuCB30piWIPi+kwOibLZLAFOApJ7YvURpZICvt2LNMgvJ/4Y4+aXynOlUX4QCU0xj9SfD/nTTa7c
lxKWg0kxwEQA+uKWTDjkEqp8snaPauQbhKAI0TGdEhIeLd+KkRbkpioffgIijy6aZsKwTzFY28SF
GccdEZlZRwQKT+TcbpjPYt4DKBMO+GnTo3IPze5vH4AyhVRJyxsUtE4mlFiHN39NNG1Swv5cWVLC
jHsda3VXxBi4uW2W2ScYEPqwcZ1zG1Kozte32RxDxW+kT8ycv4o53t+haOEOZc5nVYOaLXza1ZKj
Uyc4yvX81XCO3rUHWRc4tuD2xgxsTQguE1GKk66gFwq3jdjY6bNwBBhGj0Xs2E5q4CETbQNvshG/
wQbwquyMIrzILQFrj00KbVNysZl2kBu/D8BYMv7cekJNZe662rGxgtmtMpmqeLmd8dCnYxu2DBlT
ss2ByAbKf+vfm0TewCY4Qj1vWYOb+Ooo7ZXVouRttHFjEpNpTLkIjEwhitvNsdPKQ/DnMNPOzyMB
byOg05KniK9i663lRMhhVyTGVrAsRbjm42hRjh3diD19+h3rbVM5P1BiU9QeyrZa7XzpjjKEUqJx
MglJPndS+aVYJerBuGIDbKcI3N1lazK5AwQQxM/JuUDEbaKe2QJjhgptmxykdyWqsq0euZ7mNBl7
P8QHtThS9nAcKLwxoDdCvY3CcJigJ5uQ3lmH6DSBly8jEeeBAlMmlWOGh2Cr0xzFHfjGJWb2YAo0
JZ5kZk/B6puK0lAMyC+Mc4rFIeYIKh9DYE2ZH1HrTDzVe1ksc1YCT9yTgr7ANjb48cbaRI0RyqwX
Qrn3z3bjhccU+O3yEEW/XWuIMknKCzXZP2vxNCiO0LbYd7ZcM/2i5dJySkjrfiiAiolDNUEMfs1U
EUSDk7OYWGKetRq16QTDHdL4AyssJTzQAIcZ0huiuDjdwWmVCO3xuDAHz1eghwn1L7mi4hGx7i/s
fsKKL1oWLQXByCPuR+Kn/sZ7XDTSxhp9qMn15as2zamiw5p0X4rX8NkNV9MryChRTC+ycvvKA1LP
KyNJkk9UPIF0zdxLdaIflQOzVf7C516MXD++2T/2oYJrNytgvKYsua0GdS2VqJnjMLA10Sxf/0yy
hzyM7J242NKsCFdWDtK+d52wA1O1ptuLjKPgdDoDWFC1oLOQ1VLTW/caNe/BMr5u3i9MfLmogkcH
KR3pJTvXpchWTHLxcprV1Rcujh6ByB647blO3SbubfTBsPjo9QtEBr39BWY1SWvPK7szQWOGNSs/
40xzUVJF/A0Dq0JSzV8COAP3Zbj12HU25O7vx4VhLrOOAzDEy4/AtawHOx6L4jT+Rf0Bx00oLk+V
7nFK7LpzVeGeipNZ2RHYrkDSqvvZ9pyvLv0iIAJfd43XrVaBzabaMceNlTCpHtW6uK9iSskk8BsX
qWxIrAWejizQ0bQ+QcbCXJJvcZnnAxt+ZZl86uCxaWDaQZJtvoZA7UbBNky57OInam0tefuRnvku
WexWR/0tt12xDfjENFWqNVxU04M0RQ4t6zaCWqonusLteF3oq3BDsGq5encVlSyO7fdWzraqgbpD
YTEHYBBTOO5p1sYGZI+qsCad5XXAs32ijEt1KO9n1fMuikHzG9BXkTMGsLhzFMmJgTwmqBilU9Ku
ID13NACKn6VpZBYd0Q3WTsErRCPLJSLOLK+Tk/X/qt0HifFYyt68I1WE+CmcUeEPXc3SzDaaxvjT
a/p3RvKsYxcN+AbjuR+JFtQch2A/nSWTgJCcHXm5JQK8i2kPXKfzDDYBJR3hCUsEyuINwcv/wF40
bd1ZOk2RVoYHS7uP25OAxkQ+1E4xcOmY2sCfi0cO9xmUgsqq5AldnHjJ6Hbq7BoQ3bk1X8GBK2Tj
97KKUPsRb0YGwdz38+kIbUpSi1ZpZRh6Wn4Q8AQTXRapnTGdThR7KzyQQdXs7jHaVQi73Mup6Lau
AbKrjGb3KjvrSuAn1bYOebkxDlJmrTJPCwlpReMjeZXlpCeqixQct2Y11uf80mqaKJMbKsKdBKtO
RO3WBrud7tNeFLn2XTqp69ljYBgLaazE+MyiBIZHRt19zMEuD6HivYSnBQTEWKSsQVdBMB6l10H6
m2LwTsDR7cN3UJdWA6r1ulePZG/qcxNvjgt5ax2B3tcEOLikkfoKtbwybqZBHVjecIYZGB2sW1Zb
m4nBFCh/yH3xJ/prAZbhF9X7pXbor8sUS0XfGe+IshnW1uYScOpcZIGl2lM9BclcpQB1lfC2FYoY
vFzLeaZxdJ0VQdmS0QTevifNhJvkRZ7KYjkZ8pky6vjiNo07xu+a9ESc0ZNeGuH//6a2Wh7TAs5r
ZuUCsqwZCRceWPIC0pz4ptLfSRWqqOxkgo791h5DbaTXclxVpG1RHVp4W+/aMW7OvKwv8YRLCyQY
MvJHgbpG6W4z9y3re5LXGjnK6sVcqB6Zn7uHUv2cKyeAaAuG+5x+29bxhoaBaUKUNw//Y9HplDbk
kkXle4w0Y0lJ+Qn7BysIfwsljm9EMkzk6rD8uuWXbuAyjNbwoDDLNK5VCvXen6uMHYUAyoc12h6Q
9c1ZexUPYdWxyfqC+Rq1soW/R8Og0JGWxlPo41wBf6yWCkPZLe2meFwdCWEF2fcIsQOUqE8jxV8J
szmuZIxN1oQy/1PvNNp3igBMCk9xxTIvSKgjaDEJPXzA8HC6lLKspN3GnJv4WPAN6A2w1Mj+FAhe
peMZNQG6+1X0v/7RrtYvpWNfws3Li8yQFMWuXHNZkXHUMHNWyV5lGlkdgHwnYrO+FWeHRAyAmWcY
isakkn9O+mJLJV0sy+rehmdwFPnsbL82H1QelX/QyiQdUuXnv+yklHbTqHrd/kB/v33q3xjTTD7s
Tiyw1Iq0DoNXTg2IIn053Z6GEe1lhc4+fIHJ+P6vNW+W+QJyQHWINqupN3wVmXY47Ct+Jn2jvFuf
V4GPLIWsu/HIIs1nD0ojZsEZHwofnSihH3qGdtbFKBaLKBHpfhTqW3v+93OBKoq8mRuMe1DL/6iJ
uDf+AMWId0RQ/cgnJoyBq9c4gG7N7PBuyBCwYNwKDivl8Q/ysJTBHXWth9dGfqA/Q83gel8I3mh4
R/ZJQMNWmzCKAnYF146ZooCNeMO/6apBEpTQP4eADmc0Hg5wViJmeoyo0BMe8rHSA0Fpbp8k4EOF
3jdxLVhLHTbaHuAdlgwjIxOCElT2qi/JPLW/gqNaDCieasgZJxd6wjD6yHnwFjI9Hc01RkGLz2tY
hvpR22s5eoTzeeJW6x2prihuO+xiVLn5ZeFzMkWtnhWWe94OwoGoyFsgKjimDDEJ2ZZKGIvUvNtT
Elpvdt7Bd98a1vyMESRv4IUxtmvaUeWd7UznkPAbqQS9RZhZXAZ0tXYjMMjZpreCQdnUxnn1x+JC
JpoJXc4RZHl6XskiFu5OkcKdCo6i8YWmotSoR5ieDMsfl1OPf/oxgmG/vYaq0Zr8WAv7LAMNcC5X
80SF5X1IwBUCMxkmupajawYO9M4SG50slvRk3UT2FVPWGbfveNQNnh1Ef+GQEZPWdOFvCpxB91RO
skfOM+M5LXck9ale2OpSHWwZlJ3Y7ukok3cX+2DMa6GqTSIE/FT/CKbFjUmG5PjaS6OyHlWFsWof
CCyt+B8giGGV82CaaDMmViBgq2fr3C3COLRdxsI0rVCRpQUmyAXtuS6cMkBJanCdjHteCu+4p9ji
aVlvnR/b1nD4++/mFmvub6mpsc+RJDVMl/9z6kXZNxr30BakX5hdmBojpKadpfjec4yvWLUAR/be
SOVQIGTWg8uSqXBAhIEmQDrBh7EBNUPLUCqmu1r9yhYS4MnhuCw9pzPNKFh+ZfwVDY+Wazw9Z+vt
19FPuGu15nTrKxeYVweiYgCf915hQlQsMbN3tAbHmxq9Yrbxnl+Qq+F4hcxaWs6l2xAW4BpCKC/y
YdCPOdmf6mtK665qj8uRJ4iHcUIjSiIisU/KBIscoYaiLeTvvQRf0oUPaqbJTeg6w8ylJ6naBAIZ
XcY1owkre7rDidhogIdA0jXXMrKJJlgEoSM6MBxv+K3XqGuxJYrwL8cCl1cHxPIUMAlvO6cw2TTA
o7Q6dTShdxcGzvTTV+4xcF/Ab7uVy6TNHlee9hTSGYSPGZ/4hAXrQtCMhZbacb3wWjT50qEdWTkD
JwEFtFvB1JYXrpTIsbOOcHeTnrOkvt/pVaI4FSrdDEn7sdRgmJEKURatkZe+b2+OrmAda3X9L8fl
5RFv6exTrBsqPIiAgMm+MJe1yrytwhBgAoHd4/XIA9nC064ZIaJV07GWvISMooGxRFelZLuqaXYf
BGtbOlrENbna0CI4wW6gkfEUSu9hiG5iBboxVzuE04u1gre67rQSl3kzxMDTyqQJrOSZVgKW8+F8
PkezxV8Ww3F7nEKvP+hfgdxBrd8vuJ8zsGf71o5IsyQzT16ufd+ogzB4PSpHzSwt1iw53wHSyPFg
+gUo1l6KekEyD5/KOWNUTPKpmnFToMXcW/gOHmeVnNJOk7e0hvGuRZRXP7hydW+vG8s2V322k6Tn
/UTaXURvamPW4148oLhprpUUZq6vcIcao6+GTyGjMP3N+9T5z+0xQmkOx4ViStloxxOLt431lJfi
KWpbsB3wKhPlx7yuoojRGCAEIep0XI/h2z0BwZK9Y0V0LRKqZrDgOSG+DaEwS0PkUSdrZA0ShvBm
iN60Ea3PPiU+/IgdoTkPknFf1oIfHJhVM0UcGk8xjm6jPRhq5dEAhdiOT1vb4C3JONDNkNhVWYw9
ZhmoPDZU3EP7k1pXxKhUEP5HLhvBDM8u0EOFMu3NHXbM+1wn2AZNitD+CA7P+SHOBh7v9Ds24v8h
oGNLeIs3lT2AvZp3WbOLZ3qNdhsxxyf3yVZTq9NRqNr0OxNqwL/KTuC6I17elJho4AAri0BU7j5h
sRK6xk8sF1cyb/3LuT+VXl5+B1aWQEAcmgyWCk/h2K5TovP2oLgrU04mHo/3enTqhvRaFCFxTGYh
7q9S3re/E/dmAnxsDaJ/kM/MMc4ApvSY85e7XbfRCtz9klY+DRhwgbQDkodIh+p/sTSH0cqy/YxV
nBesHk86G//vwpVHHRtxew62o116MBj79IyoRbyNnSrvBNXanXMGWqjLdQ6YNA+bgZC0UvwvPGn2
8zp5nLpMjIYf22VwLcIhztsg9XVfebIXsv4OivZWkes7b5fT3MLil9axZOvbAtzrht9juC40LwL3
xRhhq1SVTFo9dSIlBQwWb5hM58YZVwtX9sIRmVfrhBwvoxQ7/OACM8LXT1d/NPOvTqg+ZzwKEPRY
oT1elFXsBcAJh3a3Ps976KYRjFfm4/N+7KKDG336OtSnei9DoC4/JJRtOpSIq07ZQcmYBMT7QkAL
8xJ0YwHC+ueVCxSrdqsYu0JsKcpaCFD89e6jzS+lQEx4q+spL5osicuAFt8RWsD+vChjQpsvuemj
wqwrFLKEInAUx8YJGEgtUQLf3R2TcDcN9vb1p1yRYAyqoGGI7eO7uqm2IgY06kQn/nNXr2tC+jOh
E4I2SKXqZIcLKRoOTsPlUmc5uvZiXqu1qNFJ6SIQlYvpqapvQFIqRyr0uz7X8zjs3IBh+0TjKNmI
DuL1DAl0HlpRrLkb/4D6OqeL/2gQ07uzVwWOv4PKMyYvS1nST5/rRaQ4JZu8NRUlTV7deMfsYLQp
XhVqFtaYcLsThmkJI4bcczp2oTMBlh1o//Vbr41fzA2Q1YfoB5913XyhFdkYR7EAOXdhmo7Tv20X
4U0B/rhLenUDYGnCWhwT0HonRtpNxQcSMkWDQa+KyujoMhXhb93qFEMskpUDZJ5gGaAWnRbk0qEp
1WnnUPYhj1F0gNcVqtTnQEcDO45zto8rKAfSyxE6K0Fb7S4wQRgr6qYcUlgkpWY+/RxrVLnK2nG1
lp5ryshMB7w80wpsCQfhdEOeingUEUggwk4y4NU4NqmVcs+rx0VnLTSNhOIyBk4K/S18UvX/Hvoy
80LxsRcaz56x64zJKPFk9/xp8klZhn5Q5lNLI6+NvJ2ivflocvt9HEUakXbzCLl3D6YRYHKzadWg
tjOVvHmKRVKXqK/jw3Q6ghpV2jshZiRkEV/2MATrWwWbBhqVQm8SruBUnsGcijklWJ8zTYc33cGI
e3qVLC4dFGvvEy9LX6FfWrgL7s4xJE7XxzsRrpTG/J03dCleuWG3Ip7oN0pzdjBM7hZxC6XgSlUz
6mDSwgxfDcPP+PL49efIaVmhx7bKKlftCoRs8zpaDz9dtvOpNH7RtSGsIpoYbLN3kX+P74XvwlLx
NOIA5r7e3tXsz549TzNhHEJkvmNu44iLeokz2S4N1pwKbAMFLS7+qf5G7Dm37KeUO1liXF2wAqnu
fcldwej+8pOad04Munr1jO5lcSJsbIEDBoH5U8D9pGOAk4gQwS0IQlQRgfgZ3imLOLexEJLtn+fR
4wajyjvM2fnfnyUkfS/O6Fmz4dj4KvtFO+84RpUsT7XhWOtTUypxxWKGQLBca7HOqWH4066YSHaC
RZnc7RP0YDggjscV3Tb1o1abajKFH4qyvlJaEf0zMymElDrvKM8d58Zmzxc1+C94lVqcoO0QthMh
wsr4hyX/wC36jgCbuuzzBOw5t1GDr5Cok9io+KtzzEGhQG2Ok6w8kutvf+vL4ckRAzcPpeeEjaHq
SU8ErFMbJxXfwAyIhtIbtmqr4gdHY9HLkfSNB3lAyKBeKD5RK3OIanZkT/bJ69KDO/XH/yBC2X/o
OWxwRKawiS+o3xKimh67RcVwxE/zfz2woGy7ZNWRcljemlBMFWz2oregHYTM0GxaxzxwXTrrONm1
7vMM/UD40dtG/cQ6b2V/yagzio/rGBSBxD2vNrQ0+Yedp2gLRDznNZSEi15RFStHmTCDxsgHjvEy
RQtJdwB3Gdfg9PPyCHKUTx7CpLeTNirjKYEXpqADS77J2BS/AKvtWUv1bz226i6UVaYRTRZoKbjo
7t/dIfoeDjtyIf1BfKqU+zTF3ILrLL9ZVZNTCfj0HnxOg1Vi0Ff7YAx7eUtDxZZg08gAy/3OThbC
QhNGMZTw4DfJdu3K3I2cIaZy+JIcz2IEF2ruVgP7pOokQXM2fc99B3tCQg2i9/LNG3R2/mjAZNQT
DxJI9mIHkil9KG7VmM83g7dIHv/f462rh0I+K5aNGs8S/EZvmKqEPR9T7tNBu10qeWkrfsOjqJ6t
7lStvvz7QHuP0/9LIhFXlhWpaLvnf5K+d6tQzHeB2DmlPoT9bYK711gKjl77oA8YrIxlkvtQB6qd
hIIwKprZwpVP3SGndw5IGIjfCBf5AD8qeEcS+LK3+4NeYjP+/iNg0Dg0nSbPFZJeH0gehGPfqIDL
4+KhVfm4HHb5pMPfFrPYRzUlADsEZ2ryo67CRG3ZR0qnqdTBnvjehx2sMIvPvQ2Cr25fv0S07uOG
Q6xjHbxj+mBr75Uug7fVgjzaztDHKPqBwGZ58W/aYGvkZWXtsJPdpk9WsqVYrEAjzLvAd7bxNdJb
jW/9Aie1Ky03jCkNilfj1fL6hFfH7y1KDjoWnIkOZqnTKwLSk3B9yIbyFc544g14bseNEWTtVp7Y
NZNvaWjGj8G9eEwTyVXDLrB+RCcGyl68Y1iBzizIt07bJ8r2dyK2W2di/BwB5uFROT9kcEloeRF4
mQE6dP5ddoN7zrWzNYc2gkiEXtK6eemSSnRmkDEKP5AF/NwB1fTLB6tYT+i+EtKiSLIh7VNx8FCJ
fE4ndoyUmhU0m4xdB0yVDMkYdJRZjTwLTTW9nDT52HJybQAQ1NPh08DJuqFGGcRXfO810jqItzmM
3xaA8mS8M267zcc804rmLgbYQAl1VJVkPEshPXCa+k+y92nM0KzES0y2VSO/6fvUL4Ow+a1LA0IT
yhOATmJvl8DJuJfihZkiNmq1buZq6FFc849eSeQZDOiw2DtFYys2HHqB85FPOsNlQ6ccS3u1oU9e
PWOGRlJDwXaEGmx4mHVZ5qRnkuItl792Z8vZXU06evpmfMwW7o9X2LpEEY4T1gr585or9kuWLBXA
iIyHTm/1eWbUjDkDGg7llZBnBEFA8oKYK4ZK3SZhnDg27Gy8OR30boiwg2mT5TKvUT+VmN6pzsxb
ikZLbGKQwhwHc7mijCyHIy3qfweH/7yxndcfLpRhyALH5Wjq50rDtDXpK3cWGx26oV3OBCYsou4x
962r0182TIzQpHwuudm/bkrKFhoXS+LrMXqrJZ+qIFQTTigGhAn9xZPdhtgCDK7PuXU68fEh0y3U
gg8Fm4qqNfWjhVbHPV0yoP6C+TezVJgECHNzHakfclGIHv49yQUrIsNRaUv+yh7aVzBtpXaui6MN
ByUyTP4fPEYrL5ITv9p2QdeK71Qtc9KvML6Ar83qkALOCsk5gnLUl/TBmEn1WH9laAkpCdxul02g
IVZK97yLwDA+tVzZW224J7J3MOPE8TjMuvnTbjZxUeu+P5Qy2LZvOyqXwUi2G4RullmvmC0sWhXr
ecXc0lwq/Agfn+vom93SJet7otvmsAjPkEscrFvpgTHGQulC1PvOYP+wj4xKhyJ5WaQmj/4KgAQn
zxY3f2g0guSPb9ueLpA5PLnuig6myYFVOTDaEKiAuj2e0Wn9qJW6I3YQ8wwuA30gOZYtNQZmrz/Z
CfcnELtsIQ46vink4YT3bXZO5xL/JIkgs66P0JyjWIWgBbPfvIwO21XOC+1++/pz9dILazpiNc9s
INQMY+QQejDGfTG0fR36xo2cd8D4TQdzseU1/EtjO9cQ1ItfavIWki//Zreha4KkAQbyqs9wvkE9
FTEBSs62GF40WbugC46RDbmr7aHupLY1SabBebV8YPNUY2TW8pCeVZkEPyNEnwLt2+mWIAshJrSn
oc6vnhhmVuyK3J6ThZ4iTAXhbh7A/D4PFGs6Foshb25o3rMw8NrKlmfKqSI8SelpouXfL5kLPhrd
YgyLfBtOAzE6BUdLL+0gL9WsL/FsPSf8aqOpowXBkxPtc00yNwi5FKm4loIoYOoU1v+cC/oOvc5P
uNrGJv8sjASl8w6Vp6RoLoFzLwT/rWXv8DDkRjujNkwhfo5F/PeH3CS15pBcfcFaUi3bX0k5fRmG
wFmO83KT5b9g4iVizZfH10JWinXDi36o7OGcGIf4fT9Q3WF6nSmivWUmBuDjkoCObmGgKMSgIoAR
CYhR3FH5YPSC0oKcKqQ9z/5qyqUuZ3OkYi8/UmaTHJ0PmkNZez5Q2OVDsA80sNLs2WH/90NgTY+M
mCJyrBU01J36Fbq+j2TvqAv9wdKxZf1byZLw32Ztoqb6hoIBklWuup1LYUVQlFRg5bADtK8crZPb
Dh+RQwp2t5XJGr69ND11FVM/hyMcYrtQpt7BHcSDyTDzwR8lsmJFcBQHFwBZ0IQYbhnXWbNA4iOA
7hdznz46hsxgeAKWRLu//7bp2CzNQb/Y/Yhayv6zXB9/I6F35jGDtenLHgFWfChNLZfEsM8vdAyv
1Ul6NJpwrtPRYOf24k6bG6snAzPrzB7dZYYTNDmelfTJ85yokAh35ZkJDxyMsYUbgDvTq7PP5rQm
SzdLF9I4DLWZ643bOZaZcdA4zUzNun754vhoW9ZkmarpuHH4q58JLHS/pFjNEZTUmZGEQQuJZI74
MydbL/bYrvR+KIODLn3GTALphwxebkDl/HVPQsxM1oDoU/NAWDp1qid9sNh7mvg8Sp5bqdRzGP+Y
HhgY/v8ee9SxUGhRyeeav70YfyYkcEft8Q1Nulx4gVf9g35Ji3gDWZusMKdrsLPNTyXosmThUWIB
8PTYFbyMYKo0pgGFxlYdMwXDK/tOLOEXW+XBY3K+SrqVMChiUCzSwIZS5dahIgJwxJXxLajBP0sq
UXUR3I9bXOw5PggA5k8VrhRzO0F8biFkYgTm0p/UzRGX6Nl7/o5Vqa0FaGjdNNCJTJLivx2gpMtr
fW2DAXA4mfMZ/RwgimzeRkMaD/ZPWQGBy8C02f/ZCX2LqUow7X5M/elsGG+yizHxfZ/uNuXchSKj
iKHobMQOZuf4KNAK8c0fjMbnGjc3sOAxt6r3u5wQQECYjB2weRFf88bp4jW9/mR7E25v0yg7WUhp
X48a0grE8UAXL7RZM4tMeaxALH1MdujZsmiBaE+VrXbyQ6cBYqtEoSn+DBw2JS+awAVVfZmqBwbT
PORHKQW6YIJeXHED65CU2+mo/ShbS1HpddwHdyrNLTeXGINLnWS5OfGy7kYU2OjpMuSd9U28lfb4
lW7c78P9KK/wxZE2Mi5z3IhKcxw7MK4K2l39Mi/DQF90nLfRfDN1KhciYUWJA0ElL0CUZ6oPeq0d
4CsvxRkxGWHyua/UWqAdMC3mX3V6NGXCeVS8uSgNx9g9V76Iadg90yjZqbaLvDCC7Afe1TUMYYR6
ZEwtzIkTdaA97z7Nv5F9YBa5sA5r9aKbjR/zJMJna0MGTjGTB11Jwwjbgm3vBqzOSosRp2P7tJaH
IPGXNRjW7p6IdtH1VSvHGkWLd6wA1nhrtX9lLf5b+hPdUArBY7LKLcg+aOe3XhDXlMAlNxYXmF35
0Hu2xN7yzXAVry2kuVZI4YdvRcOapsgbUWIflszWkFEN54ke0vwm9UTzBedkXttNVNBC0FrGCfVC
XRw6ZKxLNb+b5FIzGt4BLo+wa+P4Ec5d8IjM9MZHGFFYthIIm14Od3/hc/yJbqtTwowUAr29CY09
LQZFNQjUSBGCWotMInUUmkXsXM6SLw1lNMRaW6A59adgQYEAHARNnxclS7QnhJ7+iB9WAugXeMtb
bq1vIvu7dF3PcsTQdMmQTjsY7g92DysLaicqsCjc5YrtVLWxBkXg/iHXYn/Reh//a7La3EI/kMii
9KJE8Y3BwoDEM55sKN9oTq8onPc3KFzFP9nycgz4dky6CuoPbz14Y8AvLzmJTu4FtV0eSxrlrbOp
NTTvJ+n8Tjspxtp7WMm28tfNgz72x3sLXQTo3XA6rvyQBwTQVWPvfzBb1Zu1YHOl7FmeBKjROkIL
bPqtUv8DXLIZ8CYpGJiDt4Uf6cSy98TTWLPdEV/b7Ly1O5UMbJFLx/ZjGqkzSpuiW0NEdhkjtKqy
j4IM/WtUOeka9vpw840tIs1hRo1Vt0lbufNC23vU9ie20zpZ0XGqjNrBS2VqN886i5QGzU6slcmc
2aVCYA8TzXZRqGtO4fWgMdlDd6WvPf4x3px5E1dZ2WFJlH2Qf1VrX2d+c7j+3OEAruU9X47rMpoB
cqbyL/CgPy68qHbXwx77kQfZvLhv29wy+4vUeljOsEFN7pFkNl25TtkIocidq07P6f6CA15Y8Er0
XcfI0m/mcdL80azn63zBwNpmmbYTnkv8bgWL1yz5GfL29Ds0ql0OaqBoMOJtAAvo6N2bOCs+Jmzc
wX1RNaTQuqD9Xxbjx5rnbmIsYi6792L1kRRiTvQPUaRixnAC4/2TiJW9TCFbu1lP8NpOOTBadCZ5
8yoUXZ/2D+wKYJ0gsKnbFMzXxjLvi8a6wiQTBX7uPkDdsajS027guh4uHCNzYd+boSs+Y3RpGOAc
Xgg1eldubcNb+nNtzAF0ot58rHrJjf2+vUvk7t5zacsQi4/j/Cm193AAHGP9ScQv+0hrpeRHQ7f1
ifg5sWJ2yq7++HDDxco0s7baPCTdfFIUFHQndVyQu9ufj8x6RE0ow6V8zxP/cDPCl+uLB7siRASs
+59TI/6Bu5tlOK4QjPvrm8inxPNAw86wEBi0AVcYILjldEYQA/t4eBhp747XzopjE/HgnASnya2g
HJD0r4R8BoeP89P1o0Bb+mRAxt7k5xfkh9rOjvUmNcBsupT8dlr7/8VmDPY5tL+ORrSsaABoBcks
LoTK4xVNrcdIA3Ivm4ofsZW0pYwLUazJhO7p8ivO3Wq809U5dBoGEwgd6NkMmBEsrTOkc7th1iz5
tLi/oHltsnGEBUCBHbUHehVDvoiic1YXuWR24ww8rpU0HadgTR0ndPsMU6b3rBKI7VyX1fAtWNO4
AlN14AMcTS0OSphoebIK65oQ3QCwDAKc+5P99D3/W6kX516+tAjJSGt/m947TiOvKTNEbKEuDQoi
vvv2bi7ie5F+WqcsWXBOXj2Ny44cSnIm40xP6lD6xlhmi0qBkCWhT2UJt2XUZveWXDPZ15ipixDt
2wOYrlm0dUNqhR4VyX8so4ugjJAz3U+Ja0V37TakjktzpOJ8Oyi/UQmBPNzUNoLPdiQMFIR9f4Vu
7skj847ymiAJNrhRD6ZsHKf7h6Wgb+746mM+2NQOy2JUHC0kEG5bKCTwnyUnwD6U2s7fHHZOs0T7
lTUTBbep3DAikLvvzlTcohYDijJ26mcZ69MB9WWZ4G0TCIj1c0FBBPveBxuI/X6xeR/CfcxSs/YG
DlX+XsKTCUHsLAiJmRp9eiqwcR0WQDdrP2kGROMgC/OZAVJQxngoX+f66tCHEOJrH1kUU9XeID7R
RJz5Bi13rjlsLFKzRqsE6bL8DYzihmQBC6COgb86S7JpyknUHfeUMfYnsQelB6o+tq+ZcR+o5oc5
aKZJ2Zx6+fKT+jednQg5ve7Tp8cUdn7lTYpDd275xZlrNR8sZFJ7UtMOVrtU4QhpUWSly2J0vhmS
/50r+c36tdxZbTtbn+ctDUhSKFiQk11dxgon7hhXDNX4ikQOxTgvsjBqSrbRNCrdiZurUHojHmzG
iZdtzR0oJjDZ92LcMxFXMH1nkFapAJ9xIIRoUN6aZ2Wwgi5WbwwG3YLg6fwY1poff/HerMpnCHtN
LMu6Bq94y27ttWXfV3pIYTgadTqFQr/t9CrfrYTTlSNXjwrehAHLaD26hAeKRkDHv6rRyt+ww56Z
A5wOncYOO6whr9hk71dtb9ua67g78g5zl+/UPyylFYaCpWmanFNH/Qk3fzzer4BZoXZCgeZkIIyG
CDtYXTPivu6oJ2ES2LVxXpZQqxY007+RhxLAlGZKiw1zLzjMvrgEWkyfhohc5MBwpT7Qc9iP+wZ7
qtA8MH00G9iFD/bQ0f9RHp1y/+t/0+270CDfozVh4aMPx/t+1aVd2vSoA9SifljjoryXKMdBxHJ5
vEwm9BsYq+yEDmTjrvZKQp4QzPih4dhyvUueCK9FgUy+owIgV5+UhJ/U1rauSywR7aFS/RCpXze8
weTQOBeH1y4FE26n/C/5D8nvPZfSqZZd9+cz5ru4FxY+Hq8/oqMptWjqRqaG2ToTqnxnkqe4Fa9y
yo1E6/xAdgRZMDq0lUcpspBzSgQ7MGy822QuNCekMm/LUmnPHiF/04e9/i5geyL2EeeOLAxDzYsc
3vNkg0in1dWj1pSa/x5qIAfYicfmueElNwPcx78serXbkTQQrHkEVH5N9HhSXT7qU+4Z4uM1Q0MS
tHf1eWzREel9bj5yBxwxwO8puhwM7yADnAK8waWc+ptkOlt8iG8cOwUbXzCBOxu05HRDz7na3aZ+
nJwykqlFhR2TCTHqHaxfCWxdn23FmrWko9bnI+VxGY6LCysFjismVdbhzZDqWTDmJNjzFZhlhxwj
ZQwX+be9WwBBoDjKNWq85kD7ddNzWsBxf3lp2T7/5VOjqmpMMxG7C4ITRWUHY5mNsLmfY4Pv5BfJ
QzO3WWvXQSpeF7a0GqTzt1xWeqlCb5qUbyoehaVnWy+OjM5gmTfeuqa9llLSQGPIZ1sDFqdqI//Q
INluVvpvYC3PZ+MCNEWt3M9Kl9qst6Z91uNWXyeiTatnyzyBRuDw5SgXNWEpZXv6C3/FzBQBOcbl
SStKA2SUigkU/9oNLsOVnHDT7i6pYakYrU0A5XgmBSmqI4iarvxwyoe7hSgnc2AX52xu4u4O47yQ
Y2gW2WTYz/ySMHQWq6lCzqRBuHDPofMcadAQWws3iPAyZCV8fUNMfpjNvSev4RRPBGg7zt+DSHOv
UqGIrPi/koAAXSvRfLZUVrGmATLCwnKpeq+e5/bUM6I68qqzU0AEUAkhj9EEgzsa9De4rJk1+ocH
Fk2oOEdw5yW3tomz5/h5/v0L+ddungy61bKySXQKEeNRNMBqHmg0m9Km8iVVHx1ew8xeZcUJKhYK
ubIUXsU2K5gxQzmol1QQ0+okX8dVB7PGF8crk56lzizaGCAU8GNzuOTfOHzPMoKjaj8u7mCzDkgd
RQBKzC8gZMpG831tzTYeTEd2NakHww/k1Vy3gg+27GHE7XLCpS7PZI/3bF2Q9EOiS7Fex/6mYXCi
jRNY+FLI+Akk9hfHFFo0yQnaRfoORRo7Nzdiw7DsgyjpLGU9o+ytYA9KbmZWUuxlO3Q91vtOSLXf
YlCIVRTrokn2TNNqeiFG48uGFbtYlHnA3aUXd3UPBTnfI65lVRjmc2Zim7AUAa+tBicPokq0iH3s
IYVzHlHI68joNDlB8IBEOrBbmcgpyHIQv+JRnIS2IE4/aPn6VnD/e6C+CeIocmhP/kQTPcOMZuqd
hKyJ4KCLGBIX1F3CnLMHiXBglYradxxlpdmi0SpN/xp/VgghhoB62bQFBBE+84Z3TkK2cC8goWI0
OAEZUGvvOPbbzgQl0Evo46lEVH5DOeOrXbIEEGO6AfDrp+CBX1B4MYB01MShcik9pf81eBNbd8sa
megS9jeNQYAklDpLJtXU3/VWB9PEBicJqm749GQIRgIlVr4zf04HTftw1DZoBMCG1n5sWylJxxtZ
kqyI55m4NPImt6e9/O0MkHe9Zn+YTnsPtBIHlNSySMuT1vwqP/y6FgbgM7DmX5y6t0X5YfM/ndRZ
8D+o1qNIwzvGQhve8VNt+tdeTYzVNYVN0+L+S0yQDBv3+uvEFw5kfTLwQ2gVguX+/oRapqCnsxz+
35Xxw9roY5zF1RtxthILcBa8777Lwa3ypfVywmwSVrfEcBPQAOOMD6LRIGl9OLtyNEkAhmgsALAx
nDsOcVqCKUrFv8HrgJNr/VSGB+bYs74nBnJqFGKg5GdaHHZBXQvf3/slxpy9fv6vFcJfyiSqPtDB
uviQvTPuDSiaNLrAKx/iGqva9rZC2jE6InCs9fbKNrd/GbKx9sRTB/lA1FpidkSfLgg2yYaTuOYx
WBjrRkK3zkXi4JXWRoHXyM+zEgwfuPp/3EEAi6FimaFluHIiAJc4cwJOWWl3qeXpxZUmErsaVJu7
GyUFL+8CHvZlg508kS09QodJpdiqxK+vEUTz+R8piwAyWk5XGR3vz33z+e1kTxaO0wv9RNl9s6hb
RR42TncJm+2RLxA5Ft3PB2dmrJ0/5OHw2sPriUmnaNh6iuUDbAvoWf1lTiwXR8XwJTZTYYAshWZG
74K35qyterutggQbAk62ijJj0QR5n7FkxjZyyBp04HY0zDu2hXGR3Lj3R1ZsdLI1Q68YWaAyRLY4
Mn6jPT3LN2v1kBomHqcuNZY2P2LwcKlsyeOuxAXlaQIb0/AUS90NIIS9DprMIylZJGWQLJR+UFYd
2NlU5xe0zIX+BweGS6aZaG0tw6Hdvs+q2vtxQo6Ta8cw/N5ZSXxOqthQOx9yXvGZDBIUpQL8nUR4
kiN/tnTCLF+C3xNPMP7bnWkqVe36ZJPirSUhpoQGgVTNAUb/jJltas7SNlk/mwYxSRR+3tOQHiVu
MO5g771Wpg8jLcZu9ahlJ/c2NONRErk2m+hfIkZSBRtqEV1X9HyATm3Ux3+80k6patCEnuGmb4tH
RHKrlQmjcgCM4p3X5qBaG7o2bnksftaRHNZQqF+YFIeDfqReuJG962lcrx0TbfytTUS8ce2Yr2EZ
3aIJZBM1SKCapwv5sb0rrbL1f3h5m9APv+bmuAyz6wG2IKDI0eUz3rzXRhY7QiWAykriBBfiGXHe
B94oOkN0H91t5HjQL58HiJvvw0OmflFrLQo9wu9cXhF2yYa7G4fBeyZh6wBDfisPGZP7HRSVoxO8
SNZBp95kO+RFc+lNJ9edycCY5yNJURjCA1yyZLscNX0mCTgkrgZCIyzmZl2pihD0FsVpKET8eirR
jx1wq0CGqNOkt491ti8s7mxSGeNCKeGsnhbRvJ00l9UbOCA8CIZ49MsnXIfFyXADJcjYBgVAQ/8j
GO6lNkELdjZggzGBTQdrFHThnRSwyqcGox6i4KUU3qqhHVUdH7rKTbxdAy6HxgerNoVqAlZIVBUd
IofJbtf4PoqVz73aEJa6FEriSFJ47cBKC0hfh7ZZYSXr8bIyXJqgwnfE1i9ixctqekmz324JwYNz
QmHLPr7HGulKdtjHgRINnaSW9aVv3Ss3RJKVNqPNFxilTxJdLJm/hUQtilNqE2JMK2yDTITWfvoq
2H81mVJqZ67kR4OBA0R75Zyajjybg5TNq9Ns/FyPzmbQdsfjJ4wxd48vjJYvHkNxqoUNVeKIqdVj
jptaNo52MuYKjllzvd9Dnk4S7FgS714XSvSjCc6noGiyu0d8/KQvyAXrHN8AlrC4A6hy2FvgX2Ux
Xc0HcIlWna8DbkuOog077iB6NgUhm6HjHDSc0JK9pVis3z0A1xI6n9/L8UVzdyPjNc0KxouaO9aZ
AZz73kjRl7jlngP+2jsHlVGxR8hllHl3JC8DE9e5UE057OycMPvd2HRAUECEv+zrnNg1JDxG1hta
tcl2tXKCt2ZseSwgJPNjG+vflpPVdlDgSGbY1MQhsUym8faOeu5JHK2LRhoK6tR1suILZXVHYnRc
8kYwxRlZEyqhNkqWT7IUiFZyXJHDAFZCY6Yqu50D+r0jyDEBLLI2as0An4r2198zsY5bObG6MCuL
qgoaLtMzHw6adIAGkX/k6HqWrc02Q3ITzoC55Lqpxg3KaOL3daUFb/+O2zjkPqjvvQXW+GkF8YAI
6EdhNDuNbLtOJItHhTsvJXkndMx0/3F7RC0Y1XQOYWp2s9O/aoRWCH3DIu5EEw27ZFOZlMnL8WR0
CUHRQNhtSYFmfE3om0hp24431YuO7iisoq3r1Lplh6I97dif5HJPCw0xmnBhbw7HhMWVkTCtzn7j
eo5Z5ImRlRTPjApBuZX/tu0AOQVWGtZfnhPvBx4RJrS+qxlp7R3NXvnD52emkZi3MsREIXLfAhdw
F5b81pnUpb42KU/83r9n/43lGXwDe13ylctHhFkp9qB0PeMET3zdoINFTyyycwcPS5+d8EEM5ZeL
c/icJTIGTjgXKjwJnZFMpDwxZ3CpJl036B9hLBhuOmaj3kDanz+bx0KQaskVNfHxPitDde151H0s
6db9zKGehWlGWcs6wzAjT3cAnnbzSPmJ4pz6OJx2sTmASVAy/r4opxdI9iBySTjFZksRpcnVGfnk
2/NH6AwiPbA26/YFzctOe7fWtw2zbSRYhO+RqepJahSfaZx40BcqvEI+ZlCa4Klx/MbWKlcH1ltK
X4FETEOq4FsrSiXci5hN1oZ6Cg+v1lOtu51XeQZJh+iFU2qnC/RRY8cEc3x02lNYyypkUjkVqt8L
ajgOUDZMD07RS2AHO3N62WN4FcG7c8TYqOgQAOs95loI7XrmoGmFmYTQ+EOOeTXzih9F0aPen88s
MbKp63Fg41TRtiOREB8uDJDwbeL2nLTnQFhexxvllyDlYaMBTjii3CIGNibhTSvyVMgx4ume/7Mf
/XE+jjqbfD3oEAyITyo4/k1uCcnRD9O0sU1+NzYiU0EaqZedko2BWfluG4SWwR+1iqR1CkKISRRU
YbYtHM+DDBoAx0rvgVt7iajym4H0nzc7Du4tlVgezuqk8uAe0Ria3ijmBl+7Uz4lE46uvTCkfUHD
/vebxjXcgGzgfk5DXG5tARYq+ZIqH8HG5/Ff7s9GAe17nEGSNjKIOz9t6p6PAfIDdMIADMOqb/q/
nTrlsxPkgTtpmVoH1DsqSoEGOQMgEyrkkHjrEw/QtI0wE/YpdVDSg9/+evREy3pdWO4RKEEppSgq
RghQjfsyJaBdBYY65jUdWa84qc6C7jBfrjWHXY2Vl2ka2lJZCYt3CDcglBuNLAI6DlQo6FvSYEJn
elV5jmg62W27uIY4xYonsOslxnSnZ6sd+lQHao4M/WM2HxzqesHM8xRV463vz+V/2EsvL5wPYpAC
Rn5nv2kjiAlmPKCg2qLKo5D1uXxckV2yZwMl/L5mjDQE2bsyuQot0o8gVaBEW3kH1wF8lJoRVmts
iYmFlVovKxFUVsVMjh/Hx/87f4clhNtJb4r2go0d/L0u78e27eny0fSIHGqzk+u4xKSf9qPpP09f
01HvBAcVWwGBwrs7O6XVolfPfDXkFxC4crZlZjmOmu98KzcX95d0c6QXiCi8cUm2fzp/ButwGVi/
R2yNRQlj0w68IdGuLws+lT8AnJiQTc0S2WspyMQ6IGmqX9tYoUjVGcHbud+P/E1pNCp948h79UAZ
L03nHQwBjNzTKnFCBruM7jFU2Ho/QM5gA7slFWj+qK+6IU+J5BfmtUVqPeorC3jsN7AUZn2MKfk1
moplgdPh32vSuZO4vB9dOlih7whc+9q9GPfwq7r63hCoGpix6ChSdDrkuICyBPxO4VhXNriVro0Q
gi246IZBGMya0xVteXVKfvEt206g9gJHUXVZNSOTy6mryxYg5B8ps12PSCwv1uJo/51BpBqq3yJI
pSO9DiEr4rPNv+ABNEglcs7I5/Lq+amuM1i0MvklLhGEiP+XKPpl7CWWTByQNZwPG8RwEjUgF6rJ
EU2B2nRU+jA4eyzkaAuT6QQq2XpvvFzfP7642hm15Qz+iK/+rLxy0pw/VN43AUEWtU8C712lTpPL
vQb23aCMxzzm915MJecvjXFv5V6cSaj5GHtIjPwCaWDhHB6aSG6cVkEIVx6tXvsG58e59F7rEo4A
jJ1x8xXNrt5PIvWFi1Dl3aCiSogpHDA6iwcYmvN2YB0eRVMOQQ1wQXMNURX4g1IJNtG1WMP5TLyx
1xd/aTiwM9ZPI5YJ4QVDrLG/Wi5VNSno20Wa19jS+omDnGInSwYG/ctJTivmieTQ+/IFGgmD6kaN
DpKL2bfrgPoFDfJDozDIFc8s9mzuBSSwIASMA97+/mLbiE7S14rnpU/mxyqqBmIkU3R9eKxT4aKT
vbU5iDvASGy1g538T1g3pkrhJZbe5FLlMWSicwfB3yG8z7D1Xa8U+re6Qs410KdDGQ0Vl0rZP/L9
SjslBxTrlRJm9Gp/OmhvwsnfaLVE2voDTYBhXOEqN/7UcfGpaQ7NwoaKIj90j0IwOiPUtaHzuUuA
R1NnA5yQbtIG2of1kMq+4k+0oW2HK04dDjzOJEWq0d0CmtcxxRUr92oHCCRwNqzup/iZp2hLaftg
1Jj1Bo3HJtMeRGGTdhMpb1C5WzUGz+xSDQ0ouXgH4gf3bFub3AsxXxxv3fdaW6hAX2x2NQx4JUbu
2RcriRgj6Dsi8u2xB9APk8jXmgSBbMpETmiZhNP2FtruUq4ani7WTNSid4Ue80THZTvkfb31gidV
BXShdlcJnYIKsfXjdwExgkT74PB3bPdalezX50r9enXjnBDPr+OFei8QTDa8MK16KIrxpkwfvFk+
LrvMAZGVAn42Y/Ie/fFa66BLym0Xve544G9JaBfdXC4Eu0r0/+Yzf2/KAajtSi6r7B/PyUSW0fyC
BC2vg3WhOko/+h90ECuMTik6VDpzKTWhYjArST/sd3uv+gStoGa4pRoKP9kfpS2xtIp2npextli/
rev2ccO+YbULgGZQAys67FXa47djPa9qzsukrjwyRvyHI6cbT2x7pBFhycSC3kewK7CGvsi/MyjL
7jxVDjVqttdnnNHPmNODtRv8CvEGbjCurN5nn71CWYV0PLfzUAp1NMsCyTDJtGhIk5BMhnejNS83
CKFAbr5L+4LOmt6bt0YfYVgWqfa+qXqjgEkOLGWeCueUB60kSPoH49G7on+2uICrTYMP/xxvk9VY
j5P6cxYpb0OFWkdp791a+JjvwAcW/4bEE8fu8SVLoB0Z4F7CXQ2iO52NsP+QckZ5UVShNC3+TzsJ
fUIqwr1ou5W+XzpywHOQ1ibS1MWUc5+DDBrE1DVXpQsPDv3ccrY2DeYJyVRzuqg8nNItrkSteqrv
pHqQ3ukaZn4UbXknNMiMGAzIMJmaMwAXCHxwcbNuj4/E5eaRgopJPHv6RHSBifH54GAUKIUw1sIk
VQvayNs0kdTo9v4PR03dYocgGd8wLSYf2QuPzDnuHer7+W941JbHtQp/flFwp5H/SSBYfVzUh8br
oOZUeuV1RuzivK6SK9OKXXqE1Dy8DBNvYifGDXw1RLfPONTck/nrCO3a9j//KGJMhBcgtT6HyhyQ
dRJW1i+fzjbp5BRa8jWUJ9VlVz5MoKDPhAtmFpUk6pUmkeRZQKtB66EQHTO1xUac39ToTudWINzK
uIPp1G2Syld3FO68AlBj+lnIY6NlfSv+gC6rhI8beOiB9cCk+5BFI98liGvrjTKNFlag8YrCjfks
hOVhHxaOIoWc4t1UXh7kdYqpKcptgdbMfzO8d6Xq56maLu/duCdKYSv3UNoSvc/HykPURnZ3FtH+
lAzMfBgt7W6GFpeChu+JtN0eZeBb0fUywdBKN5RqS9wNWMQ85WeK8ETPApHuYOLUSAgGyghfb9WZ
4O144UueIbMWbqAFlJ+ap/SgeOvsl+7+GAb3KAoLi6FOLtBNGfBHGqzVaIP9qlmEEfle7jWMFfUg
pgzHs9uQQfhI6MU9r+vdY9wuCbk+YryuQutyGrDsc7TyUAOKVFnNQSqVZVA9QmahLz1jUb5603aB
f6ipNXDD7gEzvwQBQQxtHBIdC7reeDaGStfSXVv6+CqQ5FH/l9erEPGul/qLLO54jf0020Lt8lE0
ks0wx73CvWqbH6obcjSMmkJnLsQ0P58eNVHQB2AG7cBJbPdwqlG9JY86qevEx1awmHdbKAcfJ3Pz
/yGHbeiuh5WYoiH/AZzoCsgk08nMOAGrdPtro8ixsPhI7pRo/Gb96BNDPULbrFeCpN9gRIVVlm40
sbo8fhMPHvuBzSm44rDIhfBSlXeee9P3U6HdTtuu/n3Bf+J1wWP+ii5SXHs387lsbug+877JtJld
DAcMDXw94t5GXsOVVu/XzfW7C5BWQX0o95OK2zJxfj/GGkIt6GF+axjEhgnz7rWeWeggy6uSWx7o
OOXZGnfLFvQBygdFvarnTe4svtc2ZptXnbmfPpFtTinMRh745xdW3W7UUYLTFpcm/oUIZqaNtqrQ
Jvy7Y/5SS8wzgSsYMGRB5RTkkDYWZ253YjwoHddg0VdsMvJ0jgA1JIqJsq1NU4d2uEa9YS7NguE6
iF+EW143q9gXT2R1AlLx/PmKcIQc1lW3MtON5y0CxbNrEas6R3dHs7ZproCOpTalGKM/ETDQudfn
8eLXe9iJVy/bCRQ7GOJQLSQE3a+E6RDMuYAU3sc76drrk+RrKjHOXDvpwc1PDGDF1wZ99035oEzE
E1k43Xx6ayl+drRwx3LMSeg4CFu3U0Uyzwn6rzWknaFfkke+Uz+Cd3t1IGFsfse/xnb+c2g6L4Fg
euKhjQ57M6MZ57p8cgt/fEWmeQRngqfWBLp+t1odYaIRChqB85ajoWeHvbZvCfETIjEuvZLvcmVC
8wGR3cU2r9l0GsBvMkng/O8qDR4kPUOIk8st8mTumfJ1r1Q2xUWXY5ahDCqO6DmERr95u1kz4vTR
V9yVgvEt83lGcW2H81aWWIB06a9NSPfNehDNfW+EKpGW/+cufnHPOH77lokT7DRjwI/rCVTT1TYk
QE3qIaAMKSzLqWOhayK5yy7R5IK7XFEE341aHvwsNT7A6PavTmdT1sF3rRYZZ8dJHUAzCvtM39WR
ptgMLK9rWhLQKwNSVF7KIGJB2/uqSQ8reFJt4z1NBWUXLUAIGQBNf7ykCefL2EilzMcAlatPwCq/
S2n2IEeqIb1l0GlOdPceYWufxhn0pxFa6wk7q4pXpCskQhSoDPRnFDnke0C4jhkqVCVuYNJjGp2k
z0HTEj/5lLH8kMCAiWGgkUz2mPSYa/NFvRwmqNXCGdvg0kvezmNQeacKxlL2QbimYz2SX5ZbQnDA
iVTyiygqLBy+JCscCxlBVZ2Q6SHCqT5+7BIz2LP0JbLGjQQ3nUR7ITZgLQSDhMb7DcuHEs1pykcm
q3SU7EvXHQxFVOGs0pGYHRo08Gw2NvtvQFUDmc5PMpRP4GCwSc+QZf3pGX1lCknuiujCnXCjUikL
cTPiVbtlsEnG/cbksGrHiwYbgFSxXpftaLarq8MzW7zWxU+a3X+rNPSe5pcaJGgbNEZN7a2gX62p
+ioqDkJDhouabjoSaMgjCuJ+UNOwRBdZKQJpbxmAX5m31/bKKE/AlFhWQEvMbpfPrAp9+UiS05RT
O1MvRJcN/BtYShZWJB/m2sbFPHaojvKEUGkqPPkImqcS3Jt5gUmjfZhnv9yZMgKSZNSFDzWwLNHl
96SxZRbEOrV1mefU/cBI5voTJEN3X1mETfXKiHqB9TpszGapS6B2yLGuDcyk0ZOM7cCYZQshFzxs
eZX7ZRQF/HLzJ1gx15938nforcZNETCLk1FKPeV6+21sjZ3FWO/mXmgBjZU2QjQhz7bzNVMIckSK
rLqjO9gm3yXm0LgxMFD3/K+F3aqEWMuwWjDnArYt9cnQwrcJL1afFIP3DHlM6PcQCYkeyDTcChPe
cXt5+dwaEH/v1pxNEXg72AfoGgRCHB1IGc1HT/QhIddN1KeGvheFy+wOWZ0Nes5GWQvRmvLjNgeP
pe9UfKOvd/wUxk1eTFbEn+LMahEMqg/wNqvfZ78rzhgs0opQ6k5whlkYRIOtMDoCMpa6Gbm19wjV
hhFyW8/7/0eijzdSJp9HM7ODhvhKEJAA59yHIsAW9emAFBFTMeYLmyTEYdkNqgxgEOHHyiLz7m81
hpxwGyJMJbsBJeWQqN2GMOm1AorA5JR+jFv1RyOFc6/EaWtBmiCZ8autR1np+yBkWuSkGb4dFJZQ
jKy+QU6eJv2/YGAZi1/sKb6kslL1tic+mSS/nWI6E1zZBCqX2hRHlQaTo8REee8sm3dtKFAS1Vef
FYNco78A1v1l48TaZBpQ0SKJKub1laT9y9Z4mo2a3vaHwlf6n4iBqxXfE2X/oazepehaiJKcF7nV
vSS//YWVQ4Qvda2OMLQxKvCk1Cb/NV/vUZvu+fdI0DnDgPHJ/D80UYEHKxDatEa5LoGmTZb/GK0F
qYlVF+TNM8L5nBablMlVOsYu4Wj/ihbivSmv7NxHCIxdOCQZYaYmpy2fJ4rFxkxfL87lIVdKC56V
QCOnUGZOEKCfSUnx2zwspvVrXbH8VCJf1jZW1L8lUS9GoWB3RQ8+P0gJhFS0dsG5AMkzbCQ0eX5X
2FCo6eax+p3EjG4yYN87L+oDUdg+a3y88IzIk240+xmQ1vFmkl4jf7CvcbHMxx+5tF+xot1qywxp
Uii4qwVAd6fLSnhvjFr8GI4bemwTrLBBPFcOxRNsc4rrJZO19424EbKSdok5u4fLLbgWGr9HRpid
OnKiQhNXR6jSfHemHg55QYhDkl6nqy3ConTCOdSHCz3tQFvTwSGuYFd/LtglpohsN1xLD7AXu8SB
VJQWKrz2cllPA9OGkW2EE7phPd69/EwrAJUsY2VM9k/9FZgvwfwnboHuJJd7bgRjojVzux8r0Hgx
FPRUsqjO4CXZ6TmZYOGg/XFvhqH+5eg4g12mqu7mN1eXjSNlXr0kn1LSDXxs2mR6BXpqdu/kwTne
A314dnhUQN6UKjhzIQpbFaJNHVCJ6vaIvwz3jHikirth9Ulw1L/lvHliBF7jHTU3NqnkPJsh8BuG
kiBswxXzogFxFelcEH7NE9BiJ4U+gNKuXPxxLGm0ZPAAVLeFiAVpPQ7DdnxE7m+cyFG1pyCai6nx
m1XPmIxAEdwKP1MjIESllvTc5K4VLdut6nbg0IftrB9Ib4iQOLEV9XCzsjA+mZcPyFteE83DFTkv
R9izLC5EG3NwZR43qm6lVy6VaRkWC5Ygb6QDff6PIYr5yjOT8I+o7hgVVMKtZbsc6WkE0XM6vamD
ezVkvro45XFdaFRr9k89mt+CZriXJQ7uD9PL0+2WCPxA4SX+BZKNOkPJ3P23Wb5XFQKNncEiiz09
iBz531paZ4cyXBYe2q9qRH37jMKwCS7hpirexK4VeXRROBj+DgYlaQihjE1uHAzB4YOEONirRJkG
GgGBnynjLVrBcEmWl2A5neuywNQRujKTsAAgsCnU5XiEJ45HqvCrTubrpcmr0MofqRf1Ba/sVO9M
ydTIUQyk1SLTFsl8hEEp+fLNl+3cROOdFWHGdLahuGDa7emnJjolRHo+LaR5vN8c7/pj9Ytagh8L
FRqVFscpcqbnbjObnw0KI4zoVnE0ByORmttoqXVjspm0J8QhT+7UBt3iIELWHsdoNEsLJZVf1A4l
jPOerPMR3/5g6tEUwM8VtUP2nIXWryWh4C3nBQryvYfvc3kyUTVVAYU3O9odjJYH1Pd3yOedO8zx
H8RVk3OVy9n9A7BjyBc/P1FkZoKISt235O5Vf4MezSqtkWkpA8YRdSwgsAlopgDuLYpoF93Qk/S1
jN968pQlsmkS/75UWB8TDFvExDmmDppV2ws6xCtKcjGOwaooXWY/bpHj+deHzAu22nkKkwaYSvho
nhfsUUx2m99tjyn3bB+yNkG8MHwgTPIdq5C4KsDOvkuI/MUj2CPHcTVX8KjdF9V9KEmH415MtpI2
+7KcBK+lOyYHihP6Hfr761zzFgdcReMCtvc9eXKxi6TEAFyrV4mwrBZkAOfjgNTK29efql9A9gEb
j34/vDn9PFNx9hrijkzX5qXP92Dz0W3w/n3QT2AORmi9Duxkx1jQw4dvfiKhMhUa+pXrjzI52I31
Wr+oBwEK2NiKtCdMs0ZVFlX78x11F6viBmwfnRSkK4c+yp7907LRfdCyGObz1qAnlYVr6BoeNqi3
hHCE7qljEzlrQmUbapkkIhO+vQrFnFQLxvq5K9Nsdh/j7MmXrSKkeD/cvJQS0/snJwX8jfqIxkR+
9tbDVkZL1lsprEjIOeTNw7v31+4j0GmSqweN5X7A3C9HSY24+yjOCbU2Uo3Q+lQ7jOdU6wJngdW1
IWa94AUAn4VOnE1E8k7tUWn95ZmniB5fl0AOOWXzK1pS2O847vassiZXLPBDaIcFvZXsV9BF/YiG
VYzbVOllc5vbADzPoDtrtaN8611HixhYAHi87+gUG39Atkp4QNxSq7oeD4g2+WlaRaU+RhGvH6+X
V/Gxr4SS8xtA/VvcdI39QseUnJk+rakkBZskK6RF0vq5+Nn1O+ULG0HzgaeVJwVpdKFpPRzqb1X4
6PeasKDHes+Qn5NGxikHN7i0I9o2gDlh90uWLRqCx2y2j8M/RZfb5c4WSJ9/35xRBE0lIhdcgPj9
ltTyGuMz5KPysi0gL+JGTynuFyRcZujLeSWtfju2zfCNhTeWnRI3rae9YW0ObZW4zeXaalD5jPOL
gRibJyghU1rgIlXjGB5hsaj5QSRtu4Wm/2bFGnWsdM+McMcqCLiDmNf5QotrADLuTuTAeYqYiL0y
oLV4+jrnqRkJJEgdJKm6KjUv1vGnoZDV9gm5253dxkFQ2hNIAUNvgUrNdfO6j74S+NxA+yhImPF6
dSNiJ08dNdBU2/Yyto7++sACSzdK9Tf0QW9zVIwMz4H3ylX6+aJ1LDWGwWjfTKynKzYYNhxXurXm
HNWXtB1VllvMBhahnIXZe31//OcMv7Oce4tw3a7gBOGdUicS8kW8UV45SC9frOIB+4HSf1hVrPnj
63ZpProP3q3/ZfSu2J1aHFfl7IfoJcBhF+uGipXgiUhzp4+LWvtIIuxdA4efmg1ynRVOFoe+9/pc
Xk6c7GKHkyPCNIZC470bJjBWVecdzBX/Auf7v8685aVRtNNTyDtRsn2eIZnd+VJE1Y20c9A1b24k
Ym1oOQV71N1O9MK/YryIeKPG6+vHkuiieDP0TJ1BBRdZgMA4ol7V+4b1Q8o1aqSOpPbEZC6TJmov
BCrl9PsTmq8LjRz/oMPlF+nzQvGk2DS8ncMcIFtLS3ZBE4TLNrWpRxKRN5p4xX6tNdJhfE/TBpQ+
scvmSHgsjqjRl/1R2f9TmuInTe3ajtX093gQb5DL2WwRqJxuI3JORwumePLt5SAF+Uj2/zY5olMm
phg2t7qZvuIF1on8vGw35nypKb6l3Ux0Dfmyi8gO/x7YeI1UQjWiH3l50C/YgSeuCzYD6LDv6CAF
27++xTSvhH71VThQdOjocxiQ3E8tFwhU6eNCSUYaqFchBq8k8pZEY2NO1RfPsNsO1Ta34eLWZQdl
heNxvKnw1BOEMwDK/vTiwGfnztlwH+oOrm1fgYvVsdxU/iqTPh8FUdJkVBlV0fM74Mxy/CgI4itX
KqIpuN7QBGFiBBR7xboXnlD55oqWfJZP18mHflyU8kDsgzCOJVivOh83DTUioh0kA9ydeHojQu9M
JaAFr6BrVd7hrvsXYz0sSxav8pvIoRjV36ZBAgNkQHxBMW0JeOLoOnMXvgstp3jQ0DEGLipDCUfq
jbkpuOe6CeRARuAH0Ga9jv/lWeE1CvMsknlOiQ24xvbdit88BC7lgIEm4uV25iZkcb00scskomg7
3XdDDxvGX+H4iiwZaxwyBPmNCt+G7pvhaYpyCYnT16qfNqqfIiCYxHxBNzcP4E/JQn3j6Q7cTc54
hsLiVQyujkhtRkxYyx5ydu5MPhktNP8t5LbzHK5c3pOu7NfK4DNZu0jbSMoMedPLiO3YhR025EGM
OSq505JNhcjdyarw/4cpXb2Z4YGVAQkQujNreiS1WPktv2M76D1+VvawmFFtfXFutNchE8wHyopg
XFkI2ByNdqB/Eb2U/wx9Adg91ykrfosKRrHLU5Bi9jhX0gih7V9wiKaWSp18IKQM1sRbXTYBNzxr
DnGIusds71eBIFCzNHboLQkdUBnh0MfCwt2vsaToWQOzdiN3TyDB18eMydWT7nBIWg6nMIRg6wyb
b/j4XQ9rpKorehpM2dSgVFxjiaLFE3kah1wsbR70o6K/Z+6ZltmK3PX34gRZowahSx3+25CMf4KG
5/yLUSrsj7h6/iQg5bGLMKJmVfVFoxc5lpIWGi4RnaKYCy9n1EriafdbDgzqZ1s2cAn7uPN5wgXY
Hy2RR//ZsSijUd6tgnsbRfCN1AExZ8EPTb4WF2rGBa0F4WjH5vY6hGGxY73fH0c41uZPYwZKiLbl
rCGvH26uE+hMHvWLqvu0+absdYdKnBnnwl0LtlcGrTYCbkx99TF+5feVc5G7Jze42gGK33xi+uOl
iuvu+ziOyLQ6rHxSPWRN8wufPm1e/ZX/pegt1LmnQRwGze7gGlMfuV0qdqfZhRF37/4qwJen3S2L
HOkIVxcuW518b4gdEWNq90xfbQ5fSOmnG5JHnijiuobNMKK/E4sx04jU5cnKkZx/VvWziDXNBeyX
xy4lIVrCruCMYAmPYVrwspymaCP4f1HbcNTujForHsRWh5MW8HpSuwXEONdGonTi/LQDYzAVVsrv
T8hHd6xiXAeU+bbceUbkbeQpnQ2O5RHcJaU/GxHLsdt+MTpV9V/8vVRLdlcY1NlC4uEp0vG7H64Z
rIemOJ+4izRrKUqGNdGkwP77iilq8tlJpP8xOqm+ZTbwvIyjwwxXLtrqKn3CQUPJiSAYYumxMoBn
aHxwGvacTzTS9Ac/qbSndkzwm7/kMw5kaUlwau+AXHkuOl4BALhiwj0H1KoKuSJ8VQ38V9/kURS8
hRTrrJAG044WKQTYuvIL/ERRrKnj0ZW95jP5hloi4JB97AP30W7/Iv3B04mgyhRkjOgKUDmRpK0z
Xqpu1pJY5gh4+bM8Lok9U+zpWowJd4VfN6TPhb9Sr8RkcBJhTW9RNbBi/I5l7wKd3w0UMzhW1SDr
2SNA0SQ5aRV3sKQhJS9hBaxUNfHdipLOF8Ifpn4jj/un84oDgsO3ZbDrzXtuxSO46WPMT4LJSXVn
XvcP8rFcI2qY68NSt1l8ppYdXAbA59K55pYq8xM3oU/makR2TZBKr1IKc8HKHksJt/M4U2eXEQ4h
lKgAUFm+SyNIPsdCuISfMTygNhorTrZYV3/txWS8kY1BDawfE5xzbbqeC4ZsyzzN4PzqGiIfN95y
P715sdxpMt7vGO/iTuEHOizMj5tgldR6DkNGHwqxIZ1Mm2QmuGi2fozNWp+pbhDyrz0MtYhydTuO
pNi8399QGNMRqCd8HWNaU7XIx5kcDyZMaCRO0G9V7/FWEUN3ilShABF1qRbvMUoKfvGxq+3YOnpn
Faw0CV0Zrmb+1CXpJ1Xo/OOrtYzzpKsEp57DMe99yYa8BBtfawlzxqkBrx1yUugcgTLcGTJctIWK
4+Jf5a/Tt2v1EdMxldy08gSt7uUH70wv+4pGB8X2jfJzLUJn15F26Kjv0gILNNpLnpHQD5hzjia1
FnsHhre8IRZ0yVmJmLsShoNqFkII7vpriRQzGowdCLjOf3X5W2+XmbZx6H9qKbcTLfxQWtPV756/
6ZpX92OMt3Dm2qUUdV8kqqasoEafenjdXC0Fhsnh9vpu8aPPp3u5SQfrChvVQbgtP5wl0OO697YN
bgXCwr0B7JkeTgC73ynXR8KP6EjZq26x178tLTjlP5CVKB2WcBmn+Jti/ivwxPl3/yiCoiEPW9X4
IXpA1fF+hBJMOjJzCMr4bxTWettsMAVpRoC1UHVvAGtgCOPHnog27MCMpeo8kSEnwLNYSTGmZIgV
tJe6KBH0ecYJ0hCWhCbqk22tsDnhvb/VrfSE2gW5bDoiYmuME4Tkd2X9xK4rO/bTDQw5/HFaUemB
0bnZ2gFnMl26y6LQbWUw9XUxSgP80KA8o8BLY9gnrAWZPETAWpOz8z2MncMIfO2FaGiFsHMzoN5y
OTY2VVJ0at54iBC/8ZIipSfDGj3J8B+3muGscIg9nmb5TvBVyWEkCnIqgxu3sjGn3ibORciDNBUm
KGat/QZFt6tqlzTSUuvLSFP6Fk2hC7YpB5+sPoVXu6Qw9swjfyuFUyU6sD1Hq3DN9By21JDAJBv2
oCA6ogwpFiXL8xyF/V12k9k4jCjqNhf+Nq+OzHslGhdgjLfg6AGftvMg45+a3z3pQKXZtTPCBS4n
G6CivJZhmMsb1tOqnw5eWx/G/Y2j+8gpQYfOuUzFJbh7KoEvyEUQ0osgtDQcf2EjmicL6ENTClbQ
opKYsBdGBW8HGjJyQPUv0ANFMyyFj7V4o15p6jZRUhjvx2YFjzpkQCJD5BtvHwpGExZpVSZFXSUH
apkdrWLrMruiTc5FqCwQ6TOhNRN1zTNrgrmdtTgFSyynVummo2hBQTxbk1t5omPSZtR1T8U/LViw
8Cc1jJHmfhqvnc5YiI4A/G6F5eftAD+kq0OniRGldk04g879cE42PG9E1/8FVos8k9PB7F68lifZ
W3EbBmzoJUxXaNZIEwM5KQnt9xr6JT4uLI8P6SgRb3QMJSbP0FZ7jDHrYrxziAt7YM2zfnepQVIY
yIaUTpdGE8eAWdXKN0KmlpdpKzR43wOnSFURMzVx1LEBkS1ldAvzl52BAJjmGD0hBWoxOrPYInC1
ih1iPy9S102k8+UKg6/x/d7/cc0JNa7oeyQma9Ir/KzPd19sU1w+CohGBfg9kVpC3kxH3x34LuY1
rzVg0X2bHEF2ABFdctfvbe1ShxhxvGmnBgx3R65kmzt1k6tjf+YH5tGgMIxYGTNKNrMH6PUvpqw1
oyq5lfJo60c5EqPYY/bjobbUti3iWPsXbTzoK4A9FP9rvwflUIDnQFNzQha16/j7oL0P7FdYIlDO
IiKoYmJhueb3KIejxXiM9m4jUf4uNQVQzcJ47mFfqit/cHX2VFzmJWqZ/AqmWX4V3ZL2q2tukA3K
uVOvTNYRuMLzVOcAaIANMkSuvjETFeSTMWSCIsUXcIMW7a1ep8oBBjq+il+2e9CvHH6ouhWIk4jC
espH/cGD36RsMJPUlP9gy0J1b+55ENO1guA0OhQANE7gSlBDzc4DMYyaFDNMOkFSWruQTp2YX7RG
+tzGK4zP2QLLLBxBKCi4rjNmm1q7zyUE0MuviJVDsBPTJkIoaMRNIDA2GyRhT635HVQem3WLC4h9
FVwUR2uy6TZVckzFS/UpqXupzUJa5RGCFJziHwHIbFllDIt3RvuKl/nMktu9B/7sftsGF1W+mdo0
8m1P/scb3/Se61a6bQiVHBz625f5xXdewUf7MKNKv+3V/OjzKhV/omuD9r4yQeVrDZwRbvtcYoIF
WhDtQph5xKzIr9enGBFrZSAqj1MrgvC6dAo2KJENGlnkrMkv/FMFtl1wSJiZc9XE4biRH1b07A2T
x1vX3nm7L0qSUMROSy53B4R2wqcWt0tyOHIjImaxeT5QpwHVYNKOVFS0g/jcoUFXjqHBth+nzL/4
iJX7YgijKqWzEGcoQCvXtKBMMOPJySxoaC16Yxyb1ttzfbU4vzK9EsWMGDJLl+D+Ljl3Tojlp/hn
FFqJlEUP+tMx5klMUso2nS7oCv+CcE5Ox8FA8FMj4A44TQCBVd7S69koYz8HVlJCP1Sm4o2w/UNc
f7WwAyhKQ7lxE2OqSM7vvlli7WV9pa9z85aGlDcJlqGosRUVleJNVgESUR+EIBT0N0OMS5glfGWd
9pmfzW+/sZ4cO3Mkw4z1pT1K1iRDcS83N89suLfTzlcxIgqoG8aSOiou5b2qNUPtCvhR8huSHMlh
1WKyq7dXWuz7f2fKHgmrkuM9PNINl0MheevP8qyYVPe17JL4yG3Eb8oRSJvrzcWdgGmnSTwhvG7W
Un10fz64GBNh5usbrTUq/eMsuFmFnd1TlgcUtR5T7Gt2MCP1boBjP3chI+sE9u/CL+sDiZNjFYNt
ooN8KNr8msc0fGnBBq7wkBwd/QgeRnAms1grZBEXXzNyEyk3NFfBkhOoDdthyQIpa6cpsQqUCFtX
0CGgi/dEQgKkEBoNp4wUJlT0vXoFtGaKoys2G+fIUPyhhINBydxz3yS/seIBvoLYAYstfeUfBu23
yxmswfkO/T5q47WEHoN6LZy7k3LDG/Y4HAj+KxV8ViriwKUuH0ppp/2pE0LdBZjZaLER0f6WpFsM
HmStSQ4IYB037qVN3lDydp9AVFYWinfr24aOr68PeFZlOOfzcLqDgCAUV55hJGjzB7QTaWzXExJG
FOweOaSP9msaLaUUZXRjCWgGBDvlB1PChMaNptQzLBy2c/UzFlwFFhbHmEb+JJb6AXW/BlzeCJ4k
8yHV1LMXgrXaAwL8AdP0z9vhvi0iAvf7tFf5J/pGLt6qDDwKjyZXqxolv06ZPSrlzYD/DU4LGcIg
KiQa2gX+2C7XhtceYsoa45l/PopzAfwK6RQg7wvG1aSFkeoJbqrJvmM09M+Wi/cie+WHFUDH2KCp
DZIWZVTCfnHEqJseEWBH1u4GUqetJtZLWmABcMYKCWanU8KyWb/FrHmBgF0IarlOZKUwYoMe7fzE
WS8ji777bs14z9CwKhBA9e5Qin4RCpk1BhfRJRWgdwlMSW6iYxq99fnRz/ZvxRqpSCQrxLFsyrpH
XeCVUszlgUc60CnKmp5d34wwySLVwtOu6IgpBec0gNzT3pNwzWBWHLzKhWROra9tQAZt1BOU3KeA
hsb33C/iPXPfGKy9qHrMBtCVVTuO1yOiYuabo+24cTdwnsEvznAXUSkbMxzphy+eJ4KHcDPw2H4i
4CkxdKFFllASXJ3yyxnlAr1OIXAEXdwdbWmCpa02jiOdrHXav4/Tg7AdkBdQ+WxBwS2XnbvG9sAV
Sk5wogAD5pJkw4eiY3WAAtOqE+SaJwJPe6neme9L/Qk6o3c4breiGcdd3yI2I8wNKP2OHQj6jeUX
C0uWyD6quOdN51MLuWzWsJR4unA8y5Hib3VuU0F6j7XFv15xZWPZkX7i9mt45NfBMJOYGjV5eFI+
OXnuExw0pQ4kY7nY0DTnfFwEvQELq++64XCxsmeN4GH2pUSPsIyTTU7qiY3Nqs9d4BG+JQQcP6Gz
xeHSh49elP42Afvf/ilY0Od5a4jgSpMpicF7LxUsJqkYiW1mLcYEx9zkXkrxp8/4ZX/Bmq3kbC6Y
MBSkDJDWK1KgrPcHj3yKZG7u+SByhjswN2GnV6EBs4K7xpn0jLIrOuomd04JcYmyAxp7CS/nACM/
eXPWBbbCWEn8iAyfhM3E2qpo8O7+KxfNDY0mep3EDce0mbNfWr8MDKVaZIc+vzVa7CJhiIO3X+p3
1TDejNjiNiDEQNS+i8ZqbiiQmvu48b1XIccsxlSvdcakYDOPaXfPijBWyp8UgmGkcbzFH+/I4KtK
EHqEF32iZjY5m/g3bAwhHmoJVHUPk+CS9ghoFa+WFD71JM+osXj/5uFVkiJQJcBpW4Cu+8+BaGT3
p22zeR/L7gwUlaFcdHen/4wDJHOoXPXjPv2tww0OX8Z9X4H57uMZexCed84jAs3ZL9OdqnZp7o29
blCTrjZ0R0bcRLaTff3lRLXVegI7EcRsL8a02HGxEBr+zmMlew65aI3m9ASrCLGobMGCiiAD7YCy
XfDA6P9dfubsII/vrsu1kI7pHk6ysRJqD6ld4B6Ztq+L3PeIZRI8Fa63YmbYxV8QYOwqcYAHolqz
eCdz0GmHgK6IA8JfS+bWNnXqboE/BObhCfIeQ87Feoe0GoNHTOgY7j70N8gzlw4Z0VStK1v7p0Mt
QZnoBz9F+jrgj9/CvDTy+NYVDQDiBNuMzZoGWI0xgBCVuOYBUgWXKv/cJ746InShLrqJO6ZJLZUF
9daQhQLcFnfW94pzCeLIjPwN8I/JctZyozTs+o+X1mqqMzSNJ8xsNvG9OWN9VQHoDQlMabEmpSff
jH3qjV2P1w9AKk18x9tiPbFPzNv/tw+TOzk+pyq83rnLA1dSAvGJRgmQwBPAyQqpu4smXZ5FN5xh
N87OBs0GqxsR2y48ARP7AqBEfDqH9x8Pv/tmw3pyMRUeQpUWq6UxR7g3muL4VCfjAElUoOxrXZM/
F8Df8ZGbcQFTDjAPs62i/AD/01IidgBJIGSbKVyFbdfybcOlZ/PNhSIwxv1SPF4grk6O+NM5vKYk
RrsyAZE++DDYo1r8EWhwHoYBjQgswMVZ58CdHkT6oBj8PIVSHiwQ+aZGa7uYYFKz1NnOIdy2Db8h
pCr+x2uCquD1LnZNsUNSZskzplIoEriJUNtBa4ulyVqGol/Z6GDtb6XYdkOkBLT68eCuefr7ESkP
KXTF89CRckVyELihiASmVQLV784NCI4GitF+yhSAZGrPOocHNj/DPCKWcNVZFusGb5kwM3FNAOLO
GmIvsAQ2+cDKNYR4EY6kKHCMESw20gYToB0dbcutkj1LY2SirC/mIut+di62S0B6Hvn7OI2N4CE/
zL7oj5En7i75axS3emCh/UXt094q4Bd3ASfJC4Nf2Vm0SxhjxebXuGcvsb/fjX7TQrHKNUtW6eN8
ONYj68dPMHv/CO4T3AI6EVOX7xI21wDO4639K2dnyMsezLrCV/zvIKYSVKRz/yZMe/B8hyHnzIYy
VX3RUs+GmFT3Tffv2uuUin4ysi28iPfGpCvYA0Z0DPeWhQDGRzww70/36HoRSOXvkE6E+E8ciNpo
dqVjxxhNfGtwqYxgFv1mY231eEcSexleLPUdAH8FXAPRg5Lnc8gcu4CCRdwr9Jzh+dkZgVu6oyGa
Vd3QUroMu0qPeozwZgXjLu414zAhyR5coGKEwy6vhq/6Rs7cHQcTonSVdrAV7a2AuawlW+F6qxWY
9yHZpIgOap1QALGr9eaXpUtG+E0rJwJFUlnBycaB0bY/rVXx+0yGPEOzB2+k6swAqgZkhAQg0gsv
+SbWK6hmOMyq/aam/l+UZCM8TfdXtHNY/htzaUEPswxlyzpReT/bzIaYSYPtdEQDZQW1P8ZgsgM/
4fQZcMuun7O1imRAaw1SGAWkW3leYQQ4tgy9cFXOo0oPu0PDskDdTuOvfFw3/40eVelF2zOgFfcd
k4kEbEYI9eVgZkrfnDYtmBFtjv6xzifHjzDydBRKJBBEPqd96ediBGTi93OCRiXfH+QQg4RCRuox
F1sgbp52G70if306fPkKoqyHDRn7fzKp5RjdSgopxNfA6IVMuGWMS+DouI67naDRNBMRVQxSA37E
Ya5uw+tsODAQ9XSFtL0c3Z6GWdPoFvD3mcR9cmaERrrBDXF4rNKLGu+HNOt8zTDbn0h5u9Hd8GpX
7NShNpEZTZ84mFSed6wP+NMbrkZ93FdH9wnmPuTt8aIVwvAg8i0uv6sMLBL+xZEdVpIpPyEcwHKe
Yk9n7T6EM2TbVBJCIM4jTnCYeCNrOyki/4vKLCOQELM/4ZiCQEtFP4lVGO+UrX+yRKxyhQ2/o+0r
zPi8ZpSl+MWHb+DTp+cr5NOX3uMVUBnnxD/AKecDYUWio58KDNpk4B27mevYHshbHpAYQ8dNgDGg
6WpasYbTOw4EEv8HHP8tkCoBfVKb/qO0MmzNZ8u4ngfGRKhG63SrUIJX5QyYKzFqzBPwyrRd6qKT
emTyTChxWAayizT7RWVytIF/pcyAsFsgWykLaI247pgLKvDMiaBzq7soVf3bNzo87XprrXyQpuxF
bgj53lR2wTOAEiJdaLNZrkyIFVHZLINeREdyphwx4BoKeEvizLbPLaxIOD7la9kh+zNGgAd6Y3/d
5zC235a/HcppN8i8ohAPRLRHB8JUKxDvtX9j6BsB599bRN1rTGkCR22rIlbZX5VhHlWGsSoBUVJd
q17EfB+s6N539/RIqg7rFauHSNQQbTsri9KaCuL0oQnCaQO06ZbHnl9++AUF7LC/3V4g0dGd1DSb
nrXeZwMR/F04w7T3kibJI2ZRq4BwX/tWZbiD0c3RCJ3uAGkUluGgDHfrNOGGuqXP11jOa/cZ9THM
KjXolG3JMrPQY/15TQMaANZLCN+y4HLX3HkruwTT2DJRetbZvVYgV2RRw5eiCeczFetZtDoFDwmj
xiBwtCxq5oxdFgYEwNa6nrUu6M9pCBPLN+1uoVcrrJdUfyNVrI05wG2qpavhOIxojuaNC7PSS2K1
E/1y+koPZ4DGUaOo+23wTGV+k81f4wx6yy5S96VPkV1nu6txwGxXUY4CDnUH157N6MNj49349vjJ
qiOwW0nBm3L7qKzS4Q0QyQxQnvGhKLBjC4cZRed52am9GkV7ldf3hOU+ZmbzKNw+2ToBlcNiGs98
4vMGKbGBAZxA3QGxUHhDLrrsA1OP+et52qe6KbCm/YuLRjb+TW/gVQZEPEVUTrVcOQtWyfxSlL1U
06bOVm9A8mWcoHNjz3xHmfHYPUB5rDLI/uXW0qTFmcT3AFDOQ34ubXNNfS8WWMrHa1/2IBaqkRGJ
NaRr7bvEehzJYQSTgayM3/vGnzbxvK+d8iHKCbNA9oHCRFIxDsU4rgq+dT9gU/94gZnZqm8eLP8J
qPp5ZkgcKWrs3FRvbCO/F7L2Wou/xh4kH8veSL/gLYu+bclt1uIG8/gWIhds+dzHvkG5rEnJTRA1
7b2S0s7RrChmIKpKjAh4ZBlWGIqmBJ4rn8EZUdxdHf8k9g1LDaIy1syqoklSupos1fI7ILneK/Yq
YVHBiE8ktKpnDZoTIDPguw2xIYpyl4inR/egwq3xeDdJMpcNEk9AfI8x+uVHrz3HkcaC/VmzwYzx
Ki51/HrSsdo/AqAc1n/+deQj/e4hX80fhBOuAwIy4JnCUUFstPwvWzAAACNciexsFCW5yjsc6Yd5
xZarBm83o5O8aSam0KJlfN9rponfZZagIGYLk9wmX1xlWdj7aUpyLh1x9D9bmPABZPwUkT5Xsn9/
s4JDqO5JkEgLj1n9D7ShNamMm4rPcAf6O6xzU3yf9UUtBsm90/Mim8+NdtmjkOev5GvrOeorHAq/
BeDc0F+uYhqebWvNWhivQeX+x2Zqe5cSGi7pp72nSrLdiz1hRrnSJKm43Z/+T9XknnnUVO4sMGWL
2u7g27Dm9Gj08ORVgaCGez1rnLKJA0BYGrPpgFcM+/MmbVkF7UqrnC2smdxWivKNnQSl2i3YDucI
721HZUcV4z7gUI0l7FsMd4KC+4ECKDnvBcIBbxSJgki6HuTS4EkVvcqwyqUGEicRC0mrzXNBRw8V
YSZ/WAjG7Q0klKJ7Jp5bKXfiB5i52cbenNSwchkn9y2nQN/BnrRyjRuewgWpFz83V2B3cO9VUQKz
Es4fZzp5dBN95MZfVy9+GBWpPHFQ/CTeZwrT3uotF6BhcyugxuQ+xDfeXc/jZBiB6G5t+NDBtkzz
rsR6f/7Xd69l7BoI7rBqt5g+rysAnnMyJdiPN7cZ0Sa67ITUulhFGiCllTS9hM3YHmDFqHIYwUGy
JNOZwvNcw5Yk3UKwYttmAc0/mFFqEKwJ+4NxqOWXsQPHf2UyumaN3+cPBRihqaEcVj4cNixQet8h
Nlkv0F8P5Wqz1Hk90KvM2cBNiWreuRlZz26hkMc1K7555fVIS9F5O/UJeH1/fJB3QO8b0uI1VsOv
M2yJ6Cu2cknJx6JJsDzLKpX3v1M+5RwZ6fBI6oMYim82OYoaao2Xiem2tg4lQvMLRQzjPaFrns0u
9GwSrWMglf9JWdAjI7CfQcWdCVgjm9e0AsO6D01DOyu+RdX3fkqN0X52csrBz2wyAsH+ewCiwqTD
nN+qU/v8iTdGoL7BLUl+ypmjxh60Hf33m1WiCOluUwep3+Tgb0ls+PvgCwdZ6mU/nBqY5c+haQH3
0z+Sy8cLPsKwDaJyfsQ4fWVq5s0/IeeCghFZ6QtmAdnPhBfSkYo+tWqFqJ3ipWIs7DL+jjg0jAWn
4m+b7I+JWvgdqZe0dRyhFGAlDZo2A7D2tIBXypM+ZDbqVIa+tFqnw4Xr5LSkrhV96/SKeZUcqgx3
kSE12rPesA1j6YM3db1wv+kYEoSb3HF4yNlFwsuqxfA40Ur3cdPZnw2lX/EaFOCThTknC5d0jAHR
VdXgkDNliMWzOhOivyBqdZx90IFVPMBhprhWRgTGLng7iMjcbdi8AOX5gxAhe8t9JCiuO3QdRz+e
IPEEv1H4cfY8awCfSb1qijKh2UiDtbyczmGIgIWV6QgjwRVUB1n8wBEwhavqdR556XIt62ZYujN8
FSGeJaFik30+6tjF6nceyE8A8AOKX2nxPYF/xOTrh+OPmdKkTgdrGzcSo85LjR9JHK9oybCI1ETB
a0HO85x657+MIX+PsrtCjvnFRrWKEJliXAPH/9/EruAV6+rKzlUY4y/R1HPdiEpetnm7IS84kMcd
NWqaBAI3Lj6Ub76oEOw9b2vxsEOfSfn8nuzo4ev+7h4s7FbWlU1IXGNjuvE8o1qyo+3Ylj+YIaWc
gu3ftvkH16zkYCvqgPirzj2fwQoUviYaemtz+CxcmY01KrRUyX06Hgbsil/A3EXYe5N3NNnJ9qf/
hUndH/X9lpS/Sp97Ld3CMY2LSlo6zhoWbrwZmBTMu21RW0sXTI0V73Z8gY0r6pUtSgHn/elmm/su
bvrnbHzcB7C64utmIS6M5pzLDyiNSWdAIFGVysFp5o5iWjmiIodAMhXLqmaWcl65KKJqnTw00dGH
NvFUopvMpRNY82OSTzURgvpHN8MueMJaQTp3h3nC0Zy/L00PPvsdrMYIU0v27wqrVTdBpCPjq+IZ
u+FVYZeQ4FJAM6GShTAGSaIVi7QZhblqEwhJZrtNyO2QaxeQ4OOXG193RyaCO3Jde5hPjCxd9rBV
C82hjFVn43vQ8r9ehtPHUYvb9UCXpPuC64PIaHvhFTJw0ScL3xpnevIpeefNZX97+PAYlu3zNftP
VkggTvr1ndC28fmp8s8AsYRAdf4G88zIFMoUQ70zKbs+vBP/bwlvm+NuzFUXc3S0Wieq3eB8ucdI
JnFfWN4IJnF7GQRHg2uqGSoRqsKbLMxlDHnFECvvdnlTSkSLNPQRsfQtE60U2s77n/FL/w7hpqAU
ZGPlE97O+5yQFX/6X0InKEWz/Jc9McsM0ugI/wYbcgWc//27DkB8+udOl2IdYo1BwGQ6LhgfnxoY
XTb15L+K2ySTV8iHTAIx5Zi8kGjuUvVWI4k623SkCtjJuRfEOi8Ty+mHqpILFX4jY9aRZyGdbMDi
7PEbKCK08GIlS01iSTehuIe/v1PT8/thPeMVEGh8BkBr2Jqv/Oxq+O3GchwmUSjpFX++E9oN1kSR
WT9cnz7FmmdUTIMBc2nM5g6WGirhVBmocfTsZTUSJDV9+rA8Cn40neSr8LGoSWS4UJOpYeK2OZEc
FvetJP5qSx5mLSfp7kUZQbYHcU3ZJmCbF4f7sf8Lbpt3PG5EAjq8USnaQtHMZmva1jLom65yCRco
7pJGPhDdim0hVQrapwU1ISuhNpjugbOpXB9okBa9VElCerO8laZe59IHMfLUJZd5IhsqYJo+WcT/
XLG/02fNonp4TBK1pf0z/dDhWWzJe2FhArAofF+aOuTRMr7GsCv0auNBiugdSZzxSQYQMh3j3SvG
i13URUKUYKKNkUCjNkk07/C15YgmlqSgh0J6tgXfsgotmZy3v8ujYf/MVvRVqCThh7bEoKrFYI/6
qdl2mU6RJZfgUnSeORn/eL9gf/xYh24Ct9DFyTMUvAEbEwaTUz1fpwSbamY0YCTxXeUxPWLW588H
IpkIvio+Gdxe+PH0pbcpiufbCO8kftfGxrxMpOAahxhqlZC0+0V6y5MiD65XTBeeA0lUGyUmpFtr
/eWV3z2P589aS6rNHTA6BXsHhFWcXvl4Ea7vWNeUohlKCo4cA/4T5VbAr09WMVo0zDoGQcHE3GAN
R5mDq/5/UjRRLwJvsJjZ2M28gUbgXYz6emUKVjKjBrZXCMIfdRkPVfRL4BcaUZ8NLDGLJdUekjXN
AurHbSGga7zNfMbvo9eo7H0VvXa4XUls92OSRiE15eIdxYAdogN4ixZBep7TJNrSUkSNrFT0K723
R5Gnp1xQPPaeyFvKohFA1h3RRF8E8ER/Z23JEeIoszDJNTDEokYfo+lEalOqjVLUrxxXqAgJoZLc
jXW888LW9DUFCvgGUReFRH0vK/13LCOFLuFMYORN21VnPecF0+RWWp+d0Os5lFEcIc0at7qIjDaO
fkFDpQ38v+SJbxx3LZ5vWw5LQEbAq1r1VVeHOrwgjPKwo0+JZHHEGD4Mdv92xnTZFU9+y2arTcle
7O5wMseSzmHblFlcN7CLaiDFwqz1tV0ymT0C8JrlTsP2hDcKjPqwRbVyG0G/k0HT0AFYXja5GtUv
KCslHlH+ZfAj08UcdyG35k3D0yz9lF55eHIizdp3+1aPenA8mGH5K9efjWovlQt0WRFbwio+jTe9
H6JoPcL/X03bkAQ4GZB+GGfjs6ToFy+E2Nzuf4I0cOLdNGpzUj4xQxchs7PfZXTL8klDQAqcuvU+
s36yX3ekQCsm/1rtL/K3sV4dvKRpq5H1Vr82SiPUHi36BtWplxDy0HdnQouuCUY4a+ujCFlydf0U
qeVjeIAg4q7i0tUb3lHu7Gcj0BZGmFGpnOhvLE6dq/U/3LHn561SBAWASKaoMyyIkQeW+ftzDFEL
xs+WdOdIkLowtrKBEJKAVvNI3H6+GoeGh1z17ZJms3eP6Bq9w/LJ59WttGnLHfPVzmmMk98Y2ev9
flewdI/NYRONl8tOsyKhsdj78y4WAkZEgpWLuPqtg6j/fVjUjcqE4CmLo362DQSyeFSuTHc70RCN
MSges6uK3pQA4HPsywoz7Ea4Z6/qKJS++T9klr6xfIBFf76IiTWxPAwWn5yD0KlEu7woSDZxXvq+
q3Xfu/9N84AXePmjysR1d4eWCbTp4waAZX4SU1hSpHJi/4yKvXviD2zc70+TTuT9HD+mYZjvwtIN
P1qPcuEyW0fMYA++IqIBb/sTNKBNaJbXRV0BOTt/4yAil5fwJqmeOGa+V2qGFkGgd6SCrao5bqxk
hM4h90WkhCt88bby2RKi7CKiDBm7NV9Qd2kMH0Q/BQDhYAsGy2ruPnCikmQLGt/md6jSSOpo0qLx
IesFaGRMGnueuUjpZ2B8fzPAjRVR7g5Wspw5i4O5hwz2A/7cDq8bUy0Q4mPgoWSosyPpH5Kf39f/
3u5JtAAmqEV8I/fwbyAit/UfvML8QEgyVoM4kngUWDfLD1VmY3wy1PaB7VjH0HSGTz7iqhZQFQRq
FlKXaLrWYN+1WHQWiWp3Wm4sRCjwdM7sTf4aGt7mi+2nmy5PAduWJx8l30+vc0FblKTV4y6Ng3R0
lwQ32SIXWoGU/I8T4GdXoK2GOMbUgyialdbEkh8ZMjyno5HKaTp4MBKvqP0KfOkMcxXCJtsO4a/y
aEQzj/0aG8fIQ++U21qNfNC1ad3UwB7dM7lmFhCtl5apLoV8V3zlfewcZ/+5kWz/Ge8XQ8K71ivk
MSeojANe7cy9vrYOwrMTY9N2w3E6V7r52XPZR9R540Q6INzFAPy6unfLAw7PNTrqWnOL2V9PJSG2
wOVbQJUPFtfhQEepHQF4wsFnMgdaS4AFhTX4YLJJAl5Vm/a81/R0WnHYwYfNDiJOtG+XayQggOB4
krg0LIFvD5+rEifFrypXpeo21LWMqxlvm2PnAMLWA8bbjECCxmVRfA5ZLNTuzX9Af/PUHyn1Bjpq
XCgvvcN4B9VGa0acxQFS63ESxqaBsrp62D7bf9ywxZS7suROa155vU7UF+GhaFMHrZO3RsuYhHQS
W+ytgK36k7PjdhnQav1uZ++853vwm0eDZj0LoDfVu2LMU+T+susVbP+5fOFF5Ar/eYdPrLIgpsHJ
6UfRAMk2oBNR+cCKeweAJEQp5X6vbbJPQThEvNypMKfjznQ1dnoQKAajoUI9v+q3rzX3KKPH4/0A
11Rbft4GlEXK2deudbBFXlebp+216PxmPuSjJ4+QdYqmz8RPR/ijRhSuPBR1hKAip8g7By54Gpbi
onYIZxj90iGmKowPJQmS/Ke4tinV6kEMTxQR5l+FOvBJ0FjzFt4trvgqXndE1YEz2H4V9O7qq4Im
ZQtReQYUx1uP/DX+9bF8CrzgQIyEdqCxCtDR7SlJbY5AioBzFozyStFiNAge42nZqddhZtEWHAjl
SI6mros/Fd2RwV17v1nFBOoY4TmwY5NMfKW8sGNy6VCJM/jxnq+HCauw1BnV7EVGyA65GGuoKv5G
0M8S7w47RnR7Z2xBWQhAre/1woxILrwZf8egktRqBzaJBQisdR+ILEGLNM9ODgIYNh2OAtLkb7QF
IC1er73decDR9VYVsqYkynB6JjS20jmnLr7pTETj2SU+3V6R8wZ3+k8YWXmDrMeWGymxWzPL5WPC
pY99Eot8CGmBhZemNPazq7PCJ1gfRTyt0uPJ5McOv4N95sWogBjriYlPZwNKlwIFhVL3ngm0B96Q
b6v02GbSaBBSgSLAEzoZWQLEF31NbyYPdh/goRXtUI9fhWbBPV3nQf9U/9/OwjJjI0C/Hkze/muL
n4saRBylp91XAQqyuO/gbMrxWtSsPK0PVj/rBGrAhgPhGofl+EtZeRDAiFVlhrNL877AeK169/Pj
zojYO+qcBd3qvaYeXtJqjlcV5C1rzMZNV8YWEtdCdj75XOi04WggCOPQk1tpQa3YI4TdflaxOaZy
tv0Yfe7JxephfInnlXaXVnvIsbUNQdTzZUfE2KAN3PcFOKn19m/h0MYW9mT9MvRf5vZWw6kCVk6s
yhNx0lDGAuqVMVbZtKkdjV82U4IYgQvtYBUvtmKF1w7tS39g/ty1O5eIyqEMk7MWCF26GWxmpUSH
8NjfkkAPZJ+XYiGTRJMMd7yRZjDCCqKbuszQlw0Mux7BQbne3ycCSvhfztUNUtFQdDzTIizMnqzp
OGipWJLaU1k8pGCW1TK93U/qz4EbJAjoTfawjY58S92MQ3MicPCDavVc21zAndhv/yhk+k01snrF
z3EiH4FQtG+EH16fvKi74DEroL9w7qovjKbXgpd0U7ptKBersoErTtNbzB3wlKR90XxHmaWPHES+
0cdOLFiunMp8yLAA/pvpnBtUAkvAgTCDcGKmcJBpiHFAxBW4ThwW4EAjOn8mayTpFqe7vx83HdNB
gspZGTj/ltN/0fAY3k4OQLkDifAO6xoLwo+C5mDyeMdQzTtwCIIdySpLLjYEs0A+Djo/mXSYI6md
VHnzun0rZJ6osoqomevyAoOmYk1rDHBLc2ovgQbcGIpqpU7UkbLE7h00bhkJk9LrCujRTb6sFsKj
j31VXHoKlvmIyzwVzrIqx26IMnqVwL23zvY3CLOAaKF/ENfOrhFSSh5j8bfZDq5mBRlnX9f9Q5sR
mxFxjBzrnfAXgNZ5XcpNwglKEvRtMMW1qUk2vPUie/T7OGE26s98RuWVuOMMGVWW6ekAxY4UmhA+
yDXngAiRUma/wiU+g5HZf0yREM0dlvctXZ+t8S+o0qC2OnYBxwhrLOG95UFZCUT0HfUJbs4pQSDz
cwUJAnE5iORw4GPDndS2prQWcl3fhaXYlUvPcN5TUfJQkGeKPLan2VHsz/w4PTok0tA50fjV8Fli
puwV1AYt5GCghFM1TwXR+BIKrqRZdpw1cJYeu3xLgynhbl7U5lbh7IhkaH9nTKbd6WSGEBDa9ALs
5gtyX4ZZNA3KCytB8gichq+ob67LLu28Pivz6y1GZLGs4oOHOurQYeHNM4fcGTy3Cs5mmF6JUh5Y
EjCP+lI3P+7hfly/4gV5cSRqFpjlLuAq9pNIKuXmHYDuSotdZfols5nbAfMbcRXRgH7GHeLYXRpj
SyoI1HIDJ4Xt30o1N9Wrv0oTnGZ/Yfis3E/lt0RRAo7cDG0AbUH1j/oDoug9ZjYxG1CQQOzVQtVB
3bd4Gftq+S6Ix20UrhBWlUwHsPcBE0wwYCv/uDy2LkbEByEceOjJT60wnfkV0LBCZdCVAiplRjYh
TetiwfcFiqHt6qBRejD6PjZMRN5J/ZQYtnHaqgTm71tDo81P1ZkPoSOLy7hJk4U2klx7d9oVt9U2
S7cpib4CyhuhSYXDIGPrKmz4ixCi3NKQSN2oPcfZ5dMXavVddaP6OCiARveGUi2pTIqee78rBeIG
EXsTQc3K9UjtffvsDtoH/D1QV9fHH+51+G+YU0scpBqNcU1krbZk4fjjJFlaaiKDI33CiJZjt04j
2l6koh3BVBgM3jMOMcy9KQfYnkh6PjLIzBijxRlY6uZn1wVqRU9Uqqfuu6xy4x07rQMvPpAuW/qE
66o24yxNk9Ar0WDjv6CrVLBWPibDJeMae5WoewwyELUQcBLIGYXMsmqbXIIlLK/QnKYG/rqL08/j
rF/qAwr3Rbbxs5BiT/ir0s54GF4SY62LDdPy876gn65Pf2If6AJ2nBsqLCzzN1a9C5f6WvD6lYDk
pV2NIenq/Tv+ZBCxyMs0bcKZFJosHcgSqESUz5kvGgOEx3/DbKsokeSRrBLmfXGvkjfQmm7dwJCM
gJabHtyDv9B2uiF1Z4Tof9Y6xgQgwGiChZzbyKtFUgjw6ShYZBer79DnF7IeILI4C36W1Fr6oEXT
cxp30oVUQYDHZQK+yTUNiNH2KvOzBklx0d3L1PXyv+ejdF6ITf8bEkYP5c+wgHHq6QX2HQlslnJg
2QhEZh00aP4ZgV6yWez8N3qBUZY2yloTun2YC6I+ENzHiIlkbHC47PWAtnpx+sYHE4EhlNWL7wUs
Y8FO+407ou4E0WgTfszskz7yVsk4br5qrXBmoaKhR1M5XcD8K3zV42wUGeIAi2TcYO5G8Dxw+C6V
KxyxCzAuge0e1THuk+MNKixiqnK2PCOpNd8EJRc8CKUbUWHT0QNinI3ZqRHMVosF26P2SIuIXH1H
/E6409Oh40s69eTN66vk61cTw0Jn/8cdaz8KiRQ7xA5jMMpu0K0PlPNTN6RvtertbeNvXwgyr9Rd
OwBHBf/BnyvEhBqmuy/dJpbhptKfPW9c5GLos+YR24v0kU13SaRA7AV7S760puvat3DKTLipO5Us
07tYyWLFAloawhoAHqFzOGwlzKkgGO8W4CXglRINxuAkAeboae4eGvFZSBBWe+PnteV4eeGckLWh
TIHfHnndx7pN7kq38gMjXQ1AJx9pExtklRl6T9XUz8Wum5KbkQUOx9QBI8lA/Gxl37fuEdpyCGPc
c7PjFMutshZAK9YShX3I5aNqt5KjC672AAHyemOOuoULLFzFMBEqwLA0jUpwrSUFmoaJoaCJdTE9
JsGA/i6LdmYHAHmpMjTdJMvivliar9UxtWZ21Ve6JsxwhSwzH0yZcJv4NO/sQ7GhuIzRLf5wjbx9
pJoUwlNa1JRxBleFoSq8x2laVn8av3xrnhckLXYLf/OU6Rgc6WpHQMMtgv09KBqs1TlkBnnS2wts
9Sz6VzUrSFOQZJCd2buAOXqh7DLBcbrhl+EZO/ird9pbGlngcD/vEPBMTEEKjVP2AlmIj6uXq4iX
1C3dELxtFvIPrFJjKEwg2976ogp6v01ds1uX/kphxQqdnsCrtizsKxFVGdAg7K1yBfl43Rj1J7EQ
dAFNTmhjHrhUehDbP5tnzI1C+PLL5mOEPkYK43NIloz6wWMTUTqEBJ6+S3nBre5L2ThE4q4sm3e3
tJatbl1v1ddfhTfq/uoc/thH/yy6PvH2iN2s0UjuSDK3Z2TH1pjiI7FDVV+L2WDFZt0AjeCb9ri/
3ZdhRl+31eX5LqIZgcVTpxI6PgaTMDAbTHK4Q1HpiEpJmQawls1rk/uxPc58q1EUL+Qu8K/Aj+Lf
d9AYCXpVcExYgZ/8mKaRxEwIbiDpYRmg/6q+cu9QTpeoB0W4GFeSqr6W65i0tblcL+/oaXyzr0z/
Wn7TWkYlXBOtzBye/AwL1G4gDNTgeP4IebUvcj4neJvjY9YlZwvQoz7K1VFJ1hVU76sAMhFZHH15
kFVJvnQr2/D8IBm8tYJGerNe75hzwOQJppzvpKUw3b9vih/Ae65+invy/qFBqLXd8mhTbU9Mlsrw
FIv34zqSiyGB9f7c1B9c5/ctyM2j4yX8yPFR+6DWmetfZAG42RLLMOoROUJCygGN7hjZNm18qB8+
mEzJPEW8mjClvBhKm65LdeCaysje2RiRk8PE+lBCqzRqCnzBgx2gNvG07yB2SYDR0OQmQe/mKNIc
JZcGMsUs6uC/PGqV7sqsAKBVb0qfZlcLRwwjdJ0SKU4pK3OwhNyeX3roMd3vpUYXJdsU0BZ1nyzD
JbG4UMl4lEG5IQkGTIM0RC+55JFq6d1T6gdeY+Uy6g+okMIQF4yKiaHw3Wuq0AwlaEY+qw8aCUIS
uFXixmauBCa1/24glx5FvD2Cr9v7AdPUxsbuZr2k/S9mCItTBcr6kZ/iZiubYsSkfTA80L/ivoSf
4f5vjlAOIZ5fvNS6EHqLL/NHEPDk9ss4YyLDgHDW9g4lM6xmrbq7nlu4Dwmw75KZZ0uk7iHM2joB
ye05ZhvZs3klUeE9eMN+aDWQPjMwbCvsXwkV4dsE8lLCAbthZ2jAx3i5aDZqWF0o5UbK4U6N3BSz
2b6GZKtxGk2noDQBlHIH0LeZ7QKes7MVpwVAAv2S1xchicUipunP5Kl4XNWEYCVdHNNhDZHUX9kV
zDFk2y1cnJyn0eXbXxN/v8Q6AK0GP0ATQfWWvQfgP51EvLQChGBmqoAUzdnWL85RQOLBAAyEk6YR
OLQRzCKPDI3eMPE2Fs5iLx/JW2sFKpogCMIKZAcwkdOdohe6oMSvf6scAZ56MQm+NkM3pHtBAch6
70k/TIPTolbTKloWIOykiGp3L0YXPWEytlBZj/RplgVKNChL2jI9j+rTEEOm+aZaHLA6RrOaw4sg
m6l5bO+ms3IzaC9OWlbgt7LWVO9wvRoy8EVzSHtu5wDlcAs6t26euNthdlCH6JhnEHgdAktdV/jK
xCbRZzESET7mdzXMQJhLaKQZItj5RoYpNp91HZwz1guaJk5v8tm4ZDG20qWtSXHxaSorbDFgJys3
dvghE2JyNz7oAZy3bJVQeuP1NVhUar0y1JBJEoxNXHAP2rDp7nkHXGURJHCmfZDzZWn3jpVcYfol
v5lJYT0EJ+Wkq0vWmAbtm9DoTALpuAKVWlwIpBk7Er95IUge3nkP5LvnM1uM3ve+BMgpV2+Ho8db
953PcNojEvBMqT1y4y1oLRgIo/zxaiippdivyJdCil+FsCIzAkBp8GXQ1RMZBprt6PhdAW0bqsB6
YAmYKmMyqfRT7m/nSWliDZRCDkXwV7gUrq93rmSY8h/UEGV/MUx/JLEp3umPlXke34T3J1S9fpve
dILfukJwSHjWRetKNPPFTTsmJVW0ER0oLojhapeljThicJ9yKW8OZU9L7DRm/tuH5x7+BsBhCfsz
NQvNwEbjvTSydcYpAqjUuBhsvk2aoG0jXh+7dXarfAoN0MoPLcVSQoJLAiRrEzuuF3OKQ/nerYQ7
GR4Zq1tDf4P4VE8dXhPTnRF7Z7aqwQi7g/qMnhUA2+oEw80utZMxqlQz+ebU7R65Ui7+FMinyd4E
DuPLYxF6YAt5GhXRvsP8+xNoLX6bQp1HXj9eCKRaTUFS+U0ife4OmLYZHDV1G9Zk1/2oVReQrNgI
fyvwsbUFm8H/2xr7vk/PKEdaC9Op1s+2D3zebCUYudUFHDjzNN4LlWBzCuFHEwtgdGIEXqJ/E2r6
7Mqymq4iw44p7qzT4py2ULWIa0V0GUiBj2pFhFFo6phU9h4CqIyTJUlhk7ZSEUgD09A8Qi+OVzVe
D05+6/7919L95WZPmfQfde4tRZVcS2784ny4pb4j/h1PvvigNa99Iq0oePwBxPUfC5Si9n/NnGAu
3xoOI3aRNWuAEldQDmzEhz2C19YWpd9cuY94G3/vxwR09ET0QsKaOV2Z8jFH4BHwJCYfou9GwlVb
qUKEDwbuyMurddb3xVB7bYRLZ9cCf+8NWpHqJ1ikxzVJjpPIkx80tNXfzc/cm6E2n80+CQHhyQ+X
DXhbjfirnPyXo+bpnaK8ahQFQaJKX8MGEi5LJadXonPCGQKjsE9hVE3OZccwPKXx2nNhGtj1uIO6
NcH3ECksYCH3lorrhjafqbWaDwxNo1d0FOfBJzo0/J88VAq2QR9hFuH7fxPo7j7o8pbfKrjqPNy0
6GSjemkyPp4ZqoKw7WpfSOZutqZEccvAKZLlp+1pNijE/ebTxI14uEiFFQuUke5B8wLMoCj4DE0g
nV8IZuW1pHijmqnxh5whnuRfEB7UHr0d2ANQ5tb3QWlcY0zRGGL66jS4Gv4MivA49dE1eLAUvP7K
TGGVc9Ux4+c90gDd12fFzTjhxy2bl4+/0IWoMwWqQKU1y1Min6M/jFYsiPJi4zkxn89s0uWRk6TW
R8PB/7nQvToPBJVkhzC0tzuM3mUU7XCY6j++CJPZkS1yvQ8OglsJE85o2oe6CPeztJyu1MoPYjJZ
qta7udHiIJH5lw5tfVFKyDKyxwtzhUsf47KB5gxCTJvSliyqqGwME7HAcSYyGn2iTIwbtpOLG8fq
p4uwQyDP+IzvC3mJj7bdR7xgLXYqKTMiodRaMLfM/FsmwulgfYfIH2YZQk1IsrF1Zer70XOosOC5
W7UQNYxWA6Ik62dSQ/L17r3tFJKZbqmbikaiIw1JlIpZ4wR+SN5AGavGpmmNfL0EFh3N0MHdeeT5
+yRyrBN+pGk6mOmz7TSTW8doJJqpnwb+wWYfVHgcxqG9GaPKcCm55NqfVi2nrHL14MuqE1+CCfRs
/cdEmQRj52CYGGpNgpwIuz1k6SX5J0pMUS2Zj2nVR+eCHXt5VmMGmn5wxyaXoBv1KHcYgCO5uZnq
qZrM4Sj5g2Qs+qB2l+GK8EH2Em467FgFUHvrjnszQlqylgH6rmxBrIVcIVUF8tforI/qeZHafeC5
kWOJPH5oYXQV0HmHCX8NRsRkLhS5M055WTU6yTboMXrIR3UKugv6cLqvVzcZmyvTScCT20WWJ5fI
9ISfQQoB2Ku4TBTBSFUrUSJYhN8GjqWrxA5sSwQ971GfDj5p/U9KH+1/RHCqbpGDxUU15FhzAHTX
fSme+j0/xz5ZKgr2kncXxMNNWOjXQVSXIjPVG7VW4DLKZ1ZJfARXysjaPSovi/bdr3FFM8ovvTY9
gHDNJJCzJbPS9TUGCSs1gHo19kkX/wFsTV4OUif/wofb+oNADySg9XHbsNsxc1zoPiMik9beTDoo
RCmocZhuWKuf9HxDxFW73A2xzJe6KAtT9tcyNB+eUkJ8JgKAPoCT/qXN2VGLQ207FFdPPIwRlj0/
Rgat93Ivte2aFI/mbu6yEFqiFFl9CkV4gMJNDKcN/k+5W5wMVpYciW55YIDI0bUcuYmirdlSKgmh
kx+ejAZDm8BcUwjPiJIXy+ytxqK5FHHnsePO1Nzz26GhTpg/y+47iNmNFTprwKOQQA3rgnW81QGf
wsttyfQd+4P57EN2lo3jEmHJtsAtNIbqZtRagLPg54smVi6diKsT6OnBoj5EQlX8pE7Y5Fcc0sZh
uykE+75v6ykMeX6Qab6NR4KPQCamkRafBj8clrqLlctdtVQrqg/oPG6Nd63QypAKUbm0t9AFfCmJ
EWFHuo6qWp0KBkWrMi1m4Guy/NWvH8VjQPkntg/t/jCWX0kiak0W+i/tehgGk1h7mBYrNOEfe3/p
ZwuLiJZAkpk189Aod8PeD+peg8AMQJT/c+admCGVWrEUnmyEgQU/6f7d7Scy3vHNDQdsfvDoPVTk
fxmxVhAFLebXtX4RNZ2GzkGzbs1ZiXI0TVjJhMFjtUl9CvUmJf7a8gDjZc7ELx2qqCFkk4a4Y38h
Bnp9mSulP6SVAI36gkt2HhaFuDJ3/yjJF13odwy9MpBM/PCcBYfH/11epIXXZhd8WQ6MlbDbyLtT
emMPDKjrg3FOB3veN9VgrcBTPHf9kp66OFtpifzaNbOMtRa26v9FjCrfeOudVJafMebibqhWV8Nf
Bb266dwbe9Lyv51RngfeAdIV1vA05JUZq0J7NpVickK/k/VlVJI8VxwCLn/yoVK2uy8wrzgTON2q
0fcrVXyabhLozipM1CSChVVaPnzf8BYyA+OBKk7NNbmCR5XFGx61IBtEktF59eRjLjnGrDarljnR
6/uMtYj91dE1KiAwxTomJlAK4uiTwC4MWP7SBQGqstGkzE3v3TciV/4ETD3WHfPpjDhMAR66uqKi
kAWXP5zJ6Akr+C8mteVuoeqmCJkBOQrPsmwMTpWYDQ4DmZOv7cyvEk/jDM40ZCSxT8IF6K5FLE+c
gejiQbopRgsIa80LNsPOKoe9HHtgFn9ok7zLsmUeVy8ax61cgNR/oWXOrzQibwG7DpwU/eYg11fg
eJ9DGtiAiI70MaQogH+75ZRyABIXRB0nsnzCezaesArt27vWqOM5g+KaHuFw//ObTNQtAZySSYOI
FqloVDapmS0+uIXAKDR7jgjpYStlg7NIvyA1nQyBGlnJcRjbng++sZy7q0zvAS+aIrcly+1EGx6t
fezVqJbx4Aq4RuPepL6KvoGYapNRD2SkioNi8XBybuRHhqyYq9z7aNk7cY4yZRiYveOjNU9iwsuu
6NS8kL77HR7jH+p0tBd9iDND1YoachqesZXRjKvvT1O82KpXlIZDQCDDIUW1ZXCbyGqvWefYQtTB
8v16murddKQMqJaB4Lwi+nZpk5A6vrD8iUGkC15p8IP2HRofFUKDfN6rlIruLjuy6lvEsOTszQ/S
7QJB81hS5BcHJ/Da1/AlJ5ssbLffk4MmVeg743ULa09YoSESXz/KkqLrMmpJzjzcAh0CZOhPsNxd
UqUxBsHhs830iuwWQo1JfgxlBb8WVZiVeB8rxCr7WF9hVQJwzmqrj7fgyoG0mrVVs/n0WLAG4jH9
vFx7ph4wAwu7fKbTnXnSn/B86Z+GAtlkt5nCN+KQdhcSEK1qukYobNjQJ9y6TIIiCenkqPNBpAAa
U5arCGNobrwyv5XOGNuZuN0geGix8lZV3zQMbI52kTuJtmxlOlSRDlzPwAM37HhtZxb2PFE4Dcrg
Qo6O9tSmFxzJoa8NPQi2+4eJ2MTyBdHb4b7uli+H8PopEkhoJyFjaY6QxSVx15+Qa++0dxBdz3ht
ogp+g4SUIqAP0ieBb/3MVICc57k3HoLfi4hv00QIHQwNFt2/V+Z+3EDqSS0f+ozt8YE6hGdClD/S
XtsBzp8IiDaCE4/OUouG8mTtkWjbwX7JU+ikaYOg07SJ4x+P+e7bEB2QDq5tQLXev9pArBGHdzy7
aZ1fSi9evBVWzG+QTWbvUwbF2TG7J/Nkv+y/GAlSg0XlC1kCyoWChf4CdY+HOcd36ezoMj9TFlm+
v0Y6yCE5iHnghTamK1en/c42odAH+z5XrLIU2XmzVU8gtbkfXJVaCSjUXwS9ONcStpFR686coP+v
ikh8NJ+q593yKj37dlvQVdHt6LXPwVMs1INJ4g7TjdUZqtfiz5pgZ8bJO3kOn3KTCiuCndqHIly/
xaSllDE1H5Ib6pHLCwCECHfllXUoB0EUTOaVplNxl2xhroZ1X/McF6rI8N8z554mg6Gf6KHk9asH
niMpvAsVdmpIvEfMoLv0lvss4K0wo7NvgzxfA35Hs3m1PB53YsqZP5JIVhbeV/Hc5ROyNlXxUFrZ
9ipY6BXO7UzF41JsZVhd+ry3tWJQUCw1WvVtIsmQt637rwq5T8Jzy/ZrOHU3NWUI8sYQP9Y6c2zw
zGKNOakphr4YWDuwgyiUBfaieYM33MqSAeim8QTHAtix3zy27ny33/J6hc8lsPg20BnNFpp0Wtvv
NRKVU6nK/+qFvyaFupsrHb9fxFBHuGOYr4wcIHW8jt+lOgq344O2eO7+tzIFXj5zVusjMh4iWFZV
ieWYDrUhRYt/tb17YR+yx++PviupyYtunTSKqP9OsWKQQD3PKmf7ILAltnjyAEWUdCAKcBHJsA0m
KPEVBXdvSdexoDoxITAFdUENqr4c+QbFvMYdjb1c4VcwSF7q2bIx1fkce2YXVHHrhMHWyGZVcH9p
riTQGi+rV766DACBqPNXqv3yqzf+7HvkHqk7VC6V6Cu7Pgva2VpG/uGgHhdHsAlS3gCMB9ScFlfL
rya1Fc76J3lbXCdapu68ZxZhgVL+bqZ02CXAwkNstf41oB7m2w++5FL9Xiqx2SggQlU+Uc1942Kv
aetGc7AdmOzqGMnSPy/THUGuZeFWdIWdFx9DfHCu+gnGM+vS7u0cMDmsqyQW+vw6halm9+wGLkWn
hQosk7RTqt9WEaW/ai9DnRWlUsoUORFjpvnqtncQLFAQAwhPhM/OPCDpfLNQvW1rCOaGq4ePX5Eq
FiAxjOdNPmM0xn9N9iWE6AwDzNv3F0XH721zD4pjhxTC1OykveFaRQSODRiWjwgsdD5q9UaOqqr/
VFKjtgnw0y/wqKn1PdqxWEoP0WhrYWdReyNbYg6LVruuL0V2GJgW7uO14YOyBoNCqxi6/jFPRt7p
uDffNEIlCq/DNaH2gkLsRDLowxzv3egpruewfagQ+vDiJp9vH58vzAqSUQSBzP3S+r9IhZe2DB/5
NQzz7s4vm9jup/pulmByCt6cf7sZliXjSxfUfy03NBIl7pvB+X6/j3flr1ILxg2MW1Ka+luFD6Xm
731FXjcLJ2WGIZ1u1RC8sI31scffwA7K4o7TiJK40m1tPUCEPBcdy27NJcjktoV2/7o7KReyjeQf
h16+M8c8jXtoIPmy8wkgZCujHm+FzMVVfIz32BzMaklAiLqO3TwUFuKbcE+pbCCbrxzIXLZJIykc
Ns+5F1tXjNKKQxyL7+n92WxAGPqzM/HLFrggNGFJ8g0SgdXxoCmMs5i71STSGGZFO+feyu/EuW9D
I9rjsfnxRlXEXO2NWujWgfWlDhSzn4zJlQP3n0TCe6aF0McbA+lIi2YL1J+GLCwgk8c8ehWjTd3b
O3ZiH9e5+RiO7Zsb+hJVGA1Yr9iLjinO/n3wFJvTU/8DWFSCeRJDJ6WCqWjjwVVFEacpQUIxyuFC
o5vvStwgNi+LXpWCze/b4Fe8N3ezGC6TnVth+Zs55nU1Dahk4q6YAS5uLl3BW9N+076dzbWxnG9i
98nt5ScV8yzxfhnCfFN8M9H1FxV5HzkzKNxhRNJYtQuNh1uplxSBgH20H20Ff2W6vsynS/zUH4S5
rudh9XCjn2JNVmgbdJaSjFci9ovOeU9gSK5o8DlxmMsECuZvju2QYrkRMYUp/HBl9U/rn83/y1Qq
eoj5hDbOkrvWoemRwdCHvEI6nymoxZLOJe2vHzGXbweUm0zUxOiYtCoRgzywzS3LIzkTR9m6+QBQ
F89IWbqV+jdxmPCWXFfIZQL+PIU8QQJKno6OBXjM988l+7GAvB1fHX9Upl6J9YuA/8FAZF2gmXWG
HKbiKmXBeszDO6n4qRr0slbOV2HRz93z9dlUt62PsGY/ue90zxeRjIeIR8yByDqP+f/u0RsXDxph
tM7N5MiRCQIwbmMWAw7Uu5vd0gCK9tBK5aRE9Nl0fbPxOaka3cmmG2hMEFUppU/YqbPRDcwawZIR
HfuCyAKFrAse2ShbrcURM6q0iSYORIWK5Gld1r5XDLoi0rKJsxZLPict/FkoPbz7TlHmz2Cv8Omp
hwYq9qm+1xZsiVVf+Yp5Sd2fUyiXjucbVSxjno8jB9jBcqCXjdGylQ9lP08okGzdXpAuqt1cOvRf
tj3aO+4+8055E7H5PJom7eNzfv+rFRsISbUSNQ5sdpu9VADr712vc/qOzfZ2BC/yLshSt865OVnh
6b7NWpmTeIpbHt/jH9aQgd03Hj9m/rhhj8M+rXHOL7riP8NKZx3B5MAmJvLePXZdaZi3wG+XMBfT
VVTivgRuF89TG7j/x55myHqmbROBXx4zLVI5R3+vhQLCRKCqAwnB8TgNoptVXkplqX8RJnpQzPUo
sAi8XXUEEPVnLW/nQ34dcgxA4UCfSATkG12SYNHmuJmneqTvhCEBVG3Uv/6LfDBliaNmB6zQMeXh
KyMqw+pmtmPr5kvgD0DZSJrkJQTNh07pXQptxKcypf9YaezLsCC6T2zbwSyJR/66rcXpmVpZalHc
JECnRPVxWCcm6zUH1L6HRG68lMVPl1ZpzFc24bUK+YEjsDhEqj4DdFCf6atdByqr4dISJ0L25dZs
RjkpfHHwSETHqTmVwxpFLz9OOmq1DvvXTRiYZ7m12+gUiweY24Z+S3WYBz0b+dL9VOJ7cC/5+70P
R+ZUHLRUjF9fc+Pri8w/drMfGNYlEdpqKA8zW+hgQdN/AycHXqdj19rqSOZNNDg8PSNl3jCUgg/Y
kZuqj2UfjmBB1BRLxnrFy92gyLjhLVtLpGTmO5Y2+f59YJobxKsx4P/iCGTfu1A4MZ0xgkldj07F
qlAQSTG7pPd+NMTc098aCc6p1/iTzt0b0MoTiKN9/8W0TSnQYbLQvJOcujbUWBATCzkxDa0eQFTW
eGuJXtZExxsw/zuwUsW6F+zKAxMslS9k/mGkfRlwKviRkylpU8HfYA1BkLaODsZGDNiNScWl5BQD
51wae+7iIO2fRfhXcKW0I35wejzj8UU0qq3aDfuaFnXMqwmm1fJcQ5YmGTTV6/Eh0Pk2TH7pa7Ba
gJxXaPiDtvq8I3PtAx3If8SoUd3rUumBjentPtpKBtyxBGHOQ/MhJtiEc7c1CL+DxVtr9gYd8weB
RAjjxJsDq/AcZSN0vaE+W1BG2BhtT5JffyM4HpL/VhpqDSrV2k6HItotEXdPKyty819mdchWuNzn
TlK6+yO2Cm0da40eux9WxBzCAEggAhB1HVpiMQdQja9/jNqY1ya58Av4sAS+/0nTNogj5qOeh3uz
YHsLDT4qzjq4+n/ghZCgFHXg7isSxFUaFZt3uqPFOvBYuivaJ4zXMJ9RhbXt6pKvn62a++r0HBCt
C0AaafJfPUT2CoOjvideOooffXtd//wa3behUN3Erl/uUIRXNDN2lG2WGFiuiZoZfb3nG9wzAe7l
qOy2+BGGpllcrouUmto6w69bbyAKC4PGbOl6bKqN4HlyrOMZ+lKgEJuo3DbtThNOJpSEtZRBSybE
mEV3iAMtAG8Zv9KZFj9Vk557nlQEAIUhsjF65ZVxNdQdAJouVKQk+VTuWJyOHFvmOHkvJoK9vinU
Q1vwaq4QrYnN+LpW3Jsg86qJgZS3ViiNW+L4pm5lhbDkjjnQpitSUlt53bPyI7B8bZnUxvX2Mqu6
ax2kSDlu1c4VrhgQkIZsYOGvUGh29eJRIeVkIJs94y13CzMRkXe+wr5kRNPDE5uLUr3hwd8kklbr
zfXQLit9RazOt73+Oc9rfPY6POCftryjI15Ie4+Dp8xaFS4rHa6v3YyNuxIGoRond0FLNPHntnat
QC5/ebXf/3q6wJpH3B8jE1xEW/qW/iNqNaEr5Arpq3j4c2u/Y+nXLYAnWSEgJ2TLxI967RsxJCtM
4oqQKVdQucyZ0DbSqIw6e8BLUTvr299P2iTEry0LQR3OH+jAFDMYFQogi9LpAxnJUprbpirGpVsI
t7/GzemydF0cFIybiLDPLtKAa/CaC7omT0S2YJseEkpyl4D8eqNA8sp8CU7rwcwNSE79W1vwyqRJ
EDxKMLkWDdco5Xgh2IN8fo6LXy+azI4tbjeLsOtyV8k1q8gVHhpX3uI6iutFOhVTdszY6lH9mbI7
bN8+dwxnmCnOisRWC400bs2vx/648RhmHZxGvi7ymz8X0q9gondYCdz/OsZXd+n4l82OcLFBx1uQ
3nde9df1SoJWtVmsYA8UeGxks4boq97bijnmInLELdHJzOVI2wDQyalJLnPg6JE5MO1SF/isKZx0
82fiXlPSxg+J0YpoInj9okFGNkXfsst899WRMcwj2TSgDfkmE3pWULW2Au8YnG3VbUISMRUdeB1z
6UyMNbMJc4bcg1VBiBi+j8kRG1zqLq4/OeaUuLqr/WXhAiX5vyWXS0fdCvPY9Cb15deK89iLB484
y3H4N85xuRmrAtyoi0jcidtlDvmxYJg8begfqBRUtdECBxntQmOi5UpoPr5CsvZRFbBfGKidHQow
jH18XOyoKPkEnUnyOThjHHGOlrc3oo6V2xyFCeulShYfD8tuqYyrfPH9ghtPO6ZU+WIFnabuJnSc
Gj3bQitceCWqgFMHnZL28PcKoPCZL048CnjG6B4mEyY2eYWyar996uB6xiKjIBFYPlcv1S6MV2q+
7v4ehCQ7b7WSTpc5ap+hYPrHlIZMcSXZqSQwxdlOXhB9g0lPWGEsxc+pzpFUSNFRIHTOH96KJb6i
mAE9JcAGXnrkNvR8E22p7rHvR2pcXBWFvPaxaZ6GUC9mR+qodT1etsCiBIKxYUVtvKlelnKxNm/p
i5Y0rKnfTzdICjBnOKJjwNwDjf2ICqCLP2JpJptzKXI4ue4ZC0Uf+ldnwNLu0TWl/0lr5KuXOPv0
8JM4hbeUYejyAOmid2yuZRJ5Jw97eEMTbhPAqXr0jWEZdxYZ625Z6i/AOCoTyD5qgTNvJN37BCYB
0e8vMRB2Nqgq4vfS+2T9xCJNiGg8LzLqVrkcUJbIFZPoKLil9huGrr82nTS/QOOLDG8yf3IYbF1K
4rS09ClXq5BCkM1W66q15NWZ3oqODTlYKPGrZK8P8e9qCidb+TCd2t3h/BIRel+QlLBiuJuhiSSd
m7/jW+uS7/flvqXKYCkpkl4mZl/3r0THIngh6NhHitYxDsk/3oN18cqeEM8bhtIRxwPZJVVnWTsr
uiXewXVggcXeS8HF4QhR+uqGRd5zC2qGq0EA+bt4qid4yudDsmHXrrZxALjRBsgmat4EmDdt9eWe
c29E4odAyCDk9tqQeQF+k3UZkktTmgdUfXEHewvEnWLFvSG4bxmxZkqQq9RwzK/TNbloh5EWO8ya
5VaAYoDjJkZhe0R0ha8f4+cmuoRex2Mt45FyrPzo8Dui7oTS+gZg7zRlwvU/+c2enUXqAA/2OTGA
ATraZN5i3h1YGaRIDPc0v1CEhjxxDoo2Jq9VaR3YgdOtMDGALzukNnoj1nzU8wC3S0K9dhw8ReR/
pdrR8u7HFLznyl5veFJFPu77uLelR+tlltsEKiOWULfSaDyCNH3DGLqPcJvpkupIdCWseHjMdGn7
v9JgyGBJHuCzc5A/58MBaMcPKCRAZ90Y7cUM7yfcaTUv3cLOKnfkXXdEO/xqJoqfvIAX10Qt3/47
UUtIew+DtKra7bBslMzPNtuwlKQFycoVxTfI6KrHsGRq/owNRKtLyAkgcTPAmQlz3Eq9qx2LEVSk
A/SW1bSxW0r0urN81tbZcEjOeXLQyk9Ua+fHhCDSjtErDtsqICXJV70Q22PeCgWRrd5sdk69Er6D
VTvunLnwm549JhxrPlv+8a88zy7yoLR8EGS+fGOn3vZFJuwI6Zui+wensxKOweH6Der9JLaoqLuF
icRJsYChQwZasOuTlfJAdwpwD+A3teYLGqPhmglw7lFvaTwxLqFO1bzx8fqVtmkSU5v8mXdKhmmP
LXgcOvM74FwXlSUE2cT6MsQ+NyA6zkRsfuChfG7Oti+gtFcvPRu6JNQMpFvLiU4qDBo/ZU97FEAG
iz68FeVhXU9BPpxApI6s/JQm2EC16Vxaha6yzKXvMM8wTHZ87DoyVFU3P6q8IsCzkSiz/jp/B3IG
o9yI68boKA2LOv7+5pUs7FMenXU2NkTINTR+L6hPhOlGJuf9BLMQ9QhKxk+Pa7H5O+FAyMeP1ihw
+ubOrVDgRRTAzxSuchrFpCIMNT4D7qKjOALTBHyTKNQHEPd/nuLNI1oNutuljcGfEls5OH6bLTb3
izgXuXhWEnJVc/0pJAXCwCHsjN2NKm0PssMNs/N9WpgnDO+HiPEtJBsq4SG++ylRbJuCDdMrdGu3
6WXudQymc4zim/p/LUk7rrz1DaAhwG/ZZXfdApKH0JSTUdXPHrBY+5dcgYl2T7TPv/OgxtLTapiB
okZk5B+iNtog2q89yc+v7VbRChShY1TdT0YP2k1xEcZfocLAbCGMYtjTcCIRbbeB4rFUFwl7dKE6
IsxiY00eKONmSwf1CZ8GZH5dfcf8i7/k72hJgU+R6K2oyDYnfNjqziktom7pfP76GvSDhcSK1Vl0
H0pJR7IMzuyiCmu+GdHY3S/Lr0dsBaOvsA1xHeLhybTxzhLDy9EQc+3aqGR/fduKjjLznbFm53qt
osVqCjxaBcOMprApFzabwWyc7+lHUXJJD2fJPuj1sCZYNwPBqTFZ1ALO9rcRdztlJ9Ezjl71FN8R
NA1fvSwRwWEDd54IEoLgFY6M9uaBsg9aeu+XaW9Eot+zVlLwcy9yZcrkBGI3QhYfJkmKtLSkiRTI
OzeR+SC4YAOd7j0yHUuSHYzH3p3PJMRME0rpiRdyW9EpXSGOZUWpC2jhF0pm3eJS1zUtlrFDOwnk
PsXKx1jrK9zbfFe0MPRVEW5S5LH/GJKlP79JcGpPPk17zMAdYWgiAv0DMk5JOSz1RnD67GKBEPCz
x2epdzUnQWg0gREooha2X5fe1JmXflMM+i8tgXvikDlCbUV7BjK2nYfLgY/exGAcQ0uepx+80PpP
pWiTXcs+SOcTBF4aUbzkVhl8P5xczLK7/t+5ZnUimoJeNRK6SfYtrzdxC6v5xJBIyYJYzqalsMtk
l8lKSYdED0f3N5Wur7y6FNsQq3Kkvq5xYWZYMIpsp5uVun61/W5SafAHDSjUIi1fizqkgcRKl6C4
7tnIU0YziAwyMgoROyRdp/ABLdKiRoEkjB6wxm81tX3VGpugVLadwgM4XZW0yNm+Se7TKvf/VdA6
vD8wpl5K1kYZdO23NoPodhZZIz8Cz+ej+0PimGYBxII5r7yNbLmML5K8X65zAAjatWD3ajiUeaC5
UNgPz+Vkqp0A1xkbHe6SMAUrhrlni0/Ojp+1QoqcYnler4YWDPoYMZMAOwsHzMj/pdELA6Il2VMG
ahELtbTuq52MNNeXoFc9GYeDTqfryGWb801iLKw58/LtNVaTsfK9r9DNoda/revSA6G8e1j1F+Pe
hL4vqdvxj/1pzYlREBQ2PxYkAqT1E01xIdBT/nhlFbrg79gE2he312cCSg+DiFmtIQFAmfLdo9ol
8S3E6+lZE2xUg3e+9dI3vakvBdH/FOr+hy+l2LrdaPVyCMqtCFI5pUF+NPXsFwKqLmiQsNMh+aqM
lXi9gw+IhrrelZAzsWUBLO/EO7hjUl8rSaqDiHLZ3dCj+fZMdxYq+bvcErCQuqpgzVIe2jNTpA1I
uoTWelOWtNaVtRqIw7qHJ+Q90gSp2lunZxKEjBpepjGCPQoT9lJJOQeqqCF3ldwQrI00S1kBsic8
rPOrKprcKcs7Bcvmlr+16loBJZt4cNlGkDmMJG0KU697YJAJcohwMwIFzoERcRzt9sgC9QiKTiha
46sSXUTNHcWswtIM6jYCTg40ryFrTcTG8aj36mgu0AeIzjoqLVeP48otQrlrThK1urt4pWWYtYri
M9pzZizaH+KRDRx/1sFWNOInXxRUlLZAO996zkVcU6bWFBl3a1iqB25YrzF9AgBehsvgWpTgEJAM
Lbt5rTWSVbZdQV4yCqIISW3e5HGIWYo4YokMVvzkkV6VDAsbKCAbHNRQJ9CePzSC75gaWt46Mv4x
Mf81MLC/FEGRKqQsd98pzqsnXC4UgnFbp9jw74ZywW/uYYJ2suexb5DBzDOH5aFKWlQBD7eVibTH
RVSROxPzdGhHfGCJB4SWwiFfq2SrQE8ffxOpcyiHxVKwhubDYPvtpbfDHmc6A8pTjNxMtHJ4Xru4
lAchG2+0dugb70xTyGMV8YdLYtJO8VflwCabfeQC4i3daOY7saY3+86w4l1x3zwHZhRD9mhpovBU
RTU2aDh5MNpm8n86jBepBoRkrdmTPBUR9baBCdXL6XtnStjGx0XB02xO6YB09dsC6h7By5td8CSZ
3YTkbMmtrkJ4kFuMAl4VTE+UFIP3hnl+G4I3p4j+ZWIb95hGaZB04r6Tb5XDFJ2vqekFxmwxHnSo
No1fWuBxafdBg0Jh7tt0fjypIgRbzXhzq0HHVYSbrmODHBqa8iK1+j5rgROI4GCXZ5q6/RNRVJMZ
6+OV/SsONuPKCU9gssxM0tBEQlN9C1yuLWclJrm14JKv8MfHYuoEGrMpaLL7ioiqyCv5ZurDm97t
06FhDKgz7OyeOS/096exm4kXWldOH/znaBZ6seTzNkENAlXPWvoy67b1BE37RXMZua+rAHcVlKwx
by+F8QwK4eBmJ2uJfLmRc2t6DB2w0iXKogeOoZlOEYxlKkoMmQwj9Y2pXlIoD0C4+DLpJ9TSzz1i
z0OYXyRuJOLc+Wc0+rQtsZgaR/pJATgbiwd+a4lZIvxQdB360E32yZdlnUsyeE3tV1xlDdZIPkDB
2jb5qNtaG6vdRR+1Aq9xoxelSzAkY6RvPWMWOVTfyOPlTWy6HpPm9jSi79OafqEzdtdP23bqTXq6
BHW4nx1jZQ8wKTkR7iDKl3SB9Ola9UJuvQJaKVUJ+7D8mJt+F3S2fk8zwORWCYQsJ8hkJCgiZBQ/
1HvtUTQyocsSQymh9/xoFUSanBIc7/BtzC1MofH25jwBLNSNP+J5iTpmo1G4OZdMzHz4Ve8yNGid
0oUq1oRMvDiV9+nHqk2lg7WhEMcDqy4tDrahsahWcGZjXA+HShWE8UFdr/nSvxf/GmUv+CbtbCma
m/Huz3Xqvzh7exU97Mv0xE5XJYbkJcV2h7bKA2WICr1UNg86rxsXApYQI0emNcHpMOptR/w20U4s
/LygsCQoKBFonyny2jutq7xf+sY3AyQERW/1Rhr0j8avBYLFt3g5yAJ68Qj+uMHtmpCjxXB5CMTz
XPtQP/88oyklgpZrFlAqVsNhkxwAZuBqRiZJGSK53IsJuZF/uUna1f9sRXcJPCeGehfm7Y5A+MUz
7US1Y19cr4cwvMv1ZnDIyxDta31SrjjXkJ3fJDuJSGRHqs4zE+vDs28DAoz8Z3PJ4fC/c/AppQ8C
fCDSUeKZKDhJv2IVWcB4J/kmILfvQp/+zvb6QHi5yiC1hS5Bfv8kFfQPsafYiSCxkdayXYNRJDwP
uxIvPCd4xRM7itldsuIXb4pZRmSDMFOFl9OYeJaOGWzzCbx6UM4qH4AalegKIwKPl6vxmN4tQiTf
o9xVfb+s4z/VVzy3U6Ak8gF2yeXn1I7DhS5Q4pfqZBTe4d56tPldAgCF/afGgv1Fa0SEIyrbanKy
akDnY392MNy12LiaL+y6kjkbxqR+ZkHJCOG5ntNqz5+OqWIpNKRoLzHAXHxPoFHsIGLREvN3dLtq
8rIn0NmnqphfRBAsEqjNDb40OhD1I6AcHRebgS6b8ys2+uHh5RGJ4IixDA7DNeZia1qje6O24rPx
h8DsbYc+38rkQihBXWPua2VjUH0MTI96Lor26TQgAibYyALW0FcOpJ6xc8EA6UR1Wqz8hZr1MI2M
bPj0v4VHaWC4Y04u/JNSX3lvCcaaHfCsQfE5Qh9O4Hb4gymPp6THsVRxHWlE7H9A9mka33jRcEsm
kCMqPc5UHpxcU8+FQ8kgWZoLMNmh3QIp0h+W0nVRnvVwUSt4AmEPexQHVCBCfoH89ZrFDQ3W+tdd
iT/0nuVub2XSXEVGW2Eu3oFqFV5ZubX8Z5u4wnH56BYk0e3a30DhZDKcVAVFJqQM06lQq9E8gMQi
/B8o/k2D90w+TlqtIKxDc6IpoFZWOMJTTdzaFYt4yrF3Hlyau/eMAdPE0vF5RAl2eDftTaQYDOhi
Vb4LUX5G/Igz3rYGh1B3E+psJspCIQO9kqriocrPR5jKP3k7qNO/fivzJgBl8g8Au7OSznXqAuKn
N4KNoAY7sK12w+Y4iYpUJmrI+ZHViUrx8S685SSqYoya4t73/urYtrlsiiupwBVt1pZNzySXwE0Y
gNPlkodxsDZs/XtkZiYs2ceOW4SltcMHv9I3EJO5R/BLeWjku0L1wovWtA6VLK8ofVrMoxrqKGFH
OXFbDp/zf1gJ8YWFZGVAFDVVsnBshccZa+HeVzdykHfca4/AAoUO1cpvppiKyWWWgg5kpZbogiCI
JREnS3rq7tT89u0g3H9W4wtODFpVG62vBsZg8AAbYtaiiFLVmOWowZkT/rrpuLM3dlZf9Dzfp17N
5A7eXyg6W6E3nLjw+IedRSgkxqBU4xx6PP88z53pHvCky43QzV+LEMaHImSmN7J6l65R+DiMVNkE
eslCzGZlEHyCwthkogmvn81/ekPG2+0mzEMP7TOxeKTG9z59UhkI9+pBvoY9qJZUnPgswnPvWTHc
S61wU5HxQKOBneTCyk0BNjxA8TAsKgNooJ1VhVGZPdRsVIzOS8Ty1h7Jj5k3CfKdzNbihy8dy0vT
Bo9Hdw7cLMZSZ+/tSANSec4VBVI5K9b2ScdvUyNSlZNWfQAGYKa+9xg+AtCVYy8V5TFd81Baj3Ez
DLNIGEImLDXZoAbURXi5XWtXORXz4j2K9aG3SbxWUuKMlOZUh3NaGYwDcNazhm0jPFRTWqu94JfM
1pvX6R8IAl2GvitXonh73hSa2+Qpx89XrSDBUjPv/4kLjUNEPwWt4StBoFClKpOxt1NBWpIJDQDt
tZPjDAfJQZAdL085GxJX5zShU8XeOAFJ84hWbrLbL6nRizMjOwDDZbKzOj9UCa8F3cX7kWvnLRes
JyPLxjtFdjLqUiy3nSh+RGx/Nd1+G+p8q7zeQZpoDo4knQpLZ0BtmDFpcedrxV6jsdblkM5HeFGo
7ncAQdHzJQ0qxKkWRVEHq3KZmeiRrEPtoio38Js8aTaeddkIuJ6RBTghg8Py2cvOs9+QyqUQoyL4
so4ttL9MvYf7N0TaJAi8S1aVt9cNhKoC6wqo8udzwsbWI+ypcXJL2aHaoUlpeHhvp+buSoPAHpUm
HmP6uDhGXciv2d84ze8Jypq5VXwz2ddKGOTulLNE85F0eJw7dfBWhcBfXAX3ydzW3w5xo24EMXTl
wzwueSrbasQ3uNrpOp7OWZPDuU4+36uue9BZ7NFBj9+/LPlA3TOO0RZK/d+62iFsfWRuJwUv377P
0jhyD7RGNLWF2RLHDLr84Eei6+TDkseg/h5GaEx2qwETrFHX+cM87WHjfjP308vWFfOdl0bqiiUa
RFmdyZMW2yx4eDDq1D90cMuMktRaqzy6Xe49zrN4jW9F7PvLZ65+GDCWYeAc2b1saXVW+H1hvjk0
Oh+SuERFisvBOIyQbOFCp4W7VNG0en1dDgZp3+TkOjkUb3FlsKUMUGqLiE2HmO1vPn3VUogouIg0
ELlDEshdAhqrK6ZIcr2sRomsjjWZwi1KsLQgEk0QXVVQ5mheQ0tbKTNBEzsyPtskLvqJKFWRq8Bn
vzMtwiaQifHQbfz6Ld0jJ3dGkP3binJVDaTHl8jSJoSPWJrQqAsUUMNc+fxbESjXO8m+E3AmsP8r
o/QFPmdx4EZVTAkYNrgjSf7Yv4uKjTXu/PrgDsP9zjVjgiVbPJoDT8SZn+Y2VAyLyAOKG1CRhfHx
fwHRACsRPbNL7ifJiFhfkdaBVR2YxJv/xYWTXYXdqrJxmIkh97XaOQX7wNaIjwioyFlSQfqi8PZm
I059WNeRhDBNxg88TZJ7UjdaMhSZB35Y+grRmWiyFv8e3x2mGHFA3JhXKgDmjF1t3F0aZSHurxfZ
zKwJlOF4qxrLwqAfrqHtSumbhwGWz9HfcFU7KJJbkSldf8zu/pV4Ej6UiNRb3mwbsS1H+nI3gumy
OywN+JfyT56TQdL+SOlWfTgZ5P0kX0VxHs/kca/qEAzXkgt2g+hjls7wxS22Y/bGlPoBPvfvgkeF
0Zp+2JwaydJrB6G1FPuUrDid06kGU/lwj3OtC3HKVgKFILQ4i1fxn38TBQ0u1pY6xXF69LRNncmi
vUs3hGYpBFqUfkYyBboXk9Iba66SLA3xYCe4CWQXlQFqMtduUv4sbwnYybvvM/SGiNePqaPT+h2y
0Fufx991ieYocWQk+NiKdya6YQjrqQYLjybvy/9K0pzHHs6K/y5ezV9CPd55BvLBByY9Qs4+GPAI
M7EZQsSxpN165NczJ6Ixej9HSd5xxptW14fA/duurC2wEJIdZuS6S8EqhOpoKDlLRpzhsSxw0lqk
D2PklSeP9gmjYop5G/7g54wvdWJbCIFl4iDofkzGp3PFqdkJ21Yl0W5If4/v4ngsi7ewTCKsqwer
6NqdrIqWDaqNgQfs0EIZg+Tn5TjDGbgLLnnPKQFxmQ/UuAQ52ZcM8zHTCmqRBe/PWFsGNfv0zBtE
5fwvo5EPon49pCRhln78vUw8t6bHxzeg1cCA/B4PAQPXXV+QhS9c3XuScjyz4bR8gP839sjAhUvT
c4FmrtMddc8hCMWKD5gMsJuzXRtiNU+fnPAcJViZABZ6UKpTwQNetMEi+wKjhiT38Td4aFHqQVsO
xJd+n4VftJx3dri3UZfiKEtmzJ/4NDEgaPFwysYC6wNUFeV9gogiZ5psLerQLfO4lQFquVgTXd7+
GkGM7SU7TCqbLQz4KyJKJf2HZk1K0POG3ISQ1yXH3PpLIGeA+70wQiJzoS7vf9IUu1toLHjXn2Ym
dlWhM8ctko8kgyi5px9UBXezQIFgaqvd4HEdMD3qArYC04+6LvVgI/qVPp9s7ldGlVe9UEHcS7CO
2ehVXki6k4uuJMJGh+/hvXEAjYAr57p/RR0nhNKlgky5tkNRQMnto6In/1Q9JNR1of5bmiDOvjr2
0gIxO3Gq3Tx66WhYkJh/ObUtPEhNItYFPd0aiAnGitn0YR3/l7S0m0sXh4AH+nxupQtRdVgBFzdc
QYLVFm5r2pkVc0hXQgCxn8R8QOK769MBicW0w2FEWqYS95HzMFa3jkJhxSdKLPsc3If/6BtkE8eA
m2jn52haCLkjbQ65sZgGTc6N5Qt08i31Jahh4WbO0JLnA6usrt2ia6DdBllWJjNr/RlCRb8izUek
hHIDgL7tmLGAF4eu4TrklxU9vMflf7IhJX7y+QBVnlyzpA5lTwALlVrPNuVaV7SwF23xiDGnhmxU
Osk1sZOwoalKGu/gqOUJntZYo71JRryqbVClkkYApm+XY5ZIjLlrUaKAi+70l+qGOA6fbbeeTj+8
SQWjc36gt5ECnVHomJOUUtOBUQQYwvD6suv2NXmP5hzTLmwA33mukB0Azy+el4xL5jnkURH577S0
Cg6ZYQOA2dfXACOYbWimWPE3hO+A7a48d8diU6vlHrOb9Kp6pOACfJzCpU5HHZvrBCUb0Y3bh72+
0TVpMwRqJ6+Wa7Zy2WgUUXNRi+331gfHubPN24DwCFD3ts/CPKSVL2drJGQaQHmKCMNvY1/dIDFk
/P6T6nWicHiMqtIiy0dev3OSiquHHUCvBN3n1Fd3zjdYwZGflIOCxln2ghCG76S4ku8Umb9uX+L3
dFEGwu/2EFNuuG2yPvMUzFZJqdwkhufVx/LBohtXTjbGvMViJRHQ5nHb+5ijbWtzxrbTmXVXER+B
+g2E68JAMcBQSRDReZXy2TXZSFOlia9YJgP94hf/aivYccco5NkZP/J+B9zZEmcpjvL2PAGVlNvx
hxV9Fqr0wyOFmZdUQYdyRXOWfo8oU1CI7EXdxuISd3dpiNPj/VfqYSmjDq0wzHeup6XktokVVSG0
x8zEkc4CKs/ZzaY5zjUNwQ4eqlh9NRkxcrstphnCR/+o7pERgSN4TaQ6vmi7sGED1u01oVa6Tq1E
qGniK9uu9nJP/h/GEH857E9CKZXjwdR2NZglwYkmebcDBWBjicmEni1Z4d693EC9x3dfVdKgG8ad
kNTkpVrjmUs2ia7YCqwn/HEhz3z4MHhWJR+LJDlJOOMphXCfweI4hFHjcjeXPSZcTA9f2RoH8a8A
7IhuRxQXvmRwgJ1XxXnB713X22y786XEqpkGRWhTGck/CutOCXmWkHVTplJ8BtcRS3uiKpes+o/u
avyZXWZRyoJFjZbWdJPrACGrdux4+XAhbtVUdRUTNqs38VLWumBWXgLhrTHK7GpT3ypSyo/+CVzv
Mfvc+tKWf8nPs4M3iggjJmSfebqUcRUUZSpLdwO3vkv03ulpRJshZpjFHJFv0FDI9aCQSO/9MUYa
GNs9da/Sh/BFg+ed26/et/geYFPmOhiJaN10M6mm/NotTOSuZvZvPFT+1uS7oGUeq/X72iKY9+Vj
BHBfmfFOMfB2TNjYzj2qaW8NRTagkZ9weEcG3EEYWbntnM5SUPzpFwlEKFpuRVu7WptJuw4c0ckP
BoNQnTn9V3SEeFNT8l8jTfccteIwR/yCT5jhpHk4Tw6J+NrZkmo1a28d6WKlBOc0uUDmk1M+J95/
Q362SKtl+WivX7lbKDi0zGM0vmAErJtKCXxeyRcJvrqXEyh+uGW9r1oqiLnaSYWH8FLUGwoWnEZ0
WW/VcBMix8Kq4GE7POFLX6m79f/UqC2nfDo6EMF/q3QQCRcAcOifEHBzF4Nb05l50ct/isPeSsXr
yBfguP9Ztma3ZIViahkBPpAsRFWCyAL68mR94YevIUkEFQkUza3w3duJ8yllRW2UsjTIJMtBat5J
lFawkJT5p8Z3UDIx8DyHyyrD+zpJ5++/YSG0k0j3DOvxl5w08jWJ5ohrYVIcaniSqPARODnOEGMr
0JExcWI+zGJ5E5HWlQFYh88Xgb9UZJ3Omt+jrsRck5abKvA4/K4zWS1G7wu0hc7SThCCnpGX6fv5
0huDAqsM0O1J8ftNJ2zFQ/z923WAjwRNVxEZH5374WNeImnehbg2LGjpZjht5tKDxdAOzk/XOqDR
gxfIQho+cI40X0fZGpvAmZG6JxiCpGNnlxapL2TIGY9AWRS3WI+lyRhfgcNYdVpfJf4fboROGHMk
g3JxpqPQArnuxvPJGf1kAUAZYF/HK5hMoaXgwBzgrk6KP2BtcGcLrXxWqSTdQNISzMg5x8O1L2Y6
KkzHYgQcvLD2S5+kJjOAED00E5kEANACXwBaRdqQkv2DxBjEOg1ZvZZd7ceVohvv+4Tv0k70y55P
vH6RFKWC2FoT2KI3eXwP3IH7jMVsuRTjWrfhy4z7uaepsQ/L2BFMaSKAAmHZkgd0dDkaX4ycVI7a
UdH3G099fM8+focJvHZt7AU6GqU6aG+BKQR3Kj5C2dQr6Iw2UxtQmee2N9D7KIJzdkC4SBt/ihRl
oq3te3EXcJXVkCbULkVwIvLslsAjlOUYoLz/7M9FKQtvyW9ekifjrEJ+2VADWqdP/KHnPXjgJAqP
ECh5w2v4C+mrKcXsGSG1FSzir2O9e2cB657YgYO6fiTUeXV0TAQrkOgFz80T6i0SHRHt/DFVGFLN
6XZRE2fEuf70p0yGEjyptVDPOQoMcNhHsV2iv49DcatarN0cmFD3xNIFJ0CHeGpjDA+4TTgSyBL1
nHSVs72n0iCeiIRWqQO5cURFuXDaSc8lIec4NzoUZwoocjSMuVdq6wTYnj+mwje6LwvwsPnLO8wt
zKkGW1E3Lne49PBQX/G8f4gJqb/4c7LuBauOKp9S3Fm478fkvIlwXp5zS7LNVc4Tr+gbajUO/rzA
TYOwBTYc/8MNIvmJ7IUfgnFqvktILb2nGC5MKT7ZMs/qtegxZ67B6nzJwL+TCKFa9Mf66AKvaKyR
8EQ4RE2j88kW7DAtW28O9PO+FMeU8uMDXPf05r513AY7j61AocvNcvyyos/8vm6NdSKJjZlvdmPz
dmeePsceuVCsT7PhwoPICpWVdoT3/PRxv/Ts2INhmUkdwyI3qIVK9BxMijVodAvDPC+4GVCu9yyM
3hVx3c1Y68uhbTE/ScSGzOvzsnev+9QIPpW+AZadKy0Ks9fdDnCZdTKUKUMFLR6FNW9/xs7W1VNr
Ntcm7kvoQPAwSTrIzbM69dI8begx4pNPCZDHDjTEORx7rjBrJ4BSHvyV2Vr93Nb/7ktQ1sBzbdzH
P+MkCdUQwLWW8uLaTM/R0voxl2oYFBS87LqhxBO/mKCMySVghF6krgXx/Z+qDT+Yey918qSxB7gX
rUaf7N5UKvtFNkvMf1X2j+mxRYz/Vyt1Pkxq79BTQiD/D27H3/Qp6u3qIjvugupdIP3i+/xdvT+m
1PkKFlHIhvk5nKs8Q38wEzORPpWbXLqoHPMQlK9y6VpvWwdOx9NpcufBVVfE8lDJJY6yN1CL7R/s
a4f3ZoRtHSY8AcC/ab/K6aF1NJUXkKqmSAzsXbjvn4N3wF+9iBGCjHYXg0hXQbewwM5tZoOeRwPc
vyjrEWPmompnrIbVp8yfZRpRMNxIGkcC5/w1vEIpczAnNhVJvCQ/X72eEkLi9GonOMQrPKQGyYAD
LAvlR17qi6qiUKcRCGMk6kq4fb45kASLJJZDNaC4G2ePSrcVufrhOQ9FboN48tBwap8GShgM9AlO
W5kSUG9mkNDrzg1/7l9cbC5VchA5aOGuVwOyhVDIDzwck44WEJK4BG1jic2DEXpFHsXT7l0y0A25
qIWR673CjCAU3WkXPOXnKbBHP1f0hQjODZ+wBauAINaSnVS2RfvWy8RCIw4cgNK10CmY8PVQw+v1
+rXadIHRySEjZegvQB5emYkQfNG1aHoa3MPFNoVZdYpo1zBP/HlofY1DnMBsEejGODVs2gVaaLn6
WbSTc8Hl4PVMRdtxCOTPEYheu16e0S4mpo44gqd3vMRHa5UfnyN2/s7r36C5wcYGlV9ZFbrNFpqS
FfFP+ZOCdnZh4wWvXgu2sIoiIuPHjo3vMck+JzLbzhMHOp3ClVeN/qc+R43+mfji1ne+DH0NLCNH
tBebqsHfW+DhrSDT2nfDzSIxY+hCwSerE4JWrF03sZhDWEBc9UbaWFrBidqgGHeaNkHgM+e0mjdb
XbE+hI6eT9l64IHywvU2fzODqWDYTZ4t/HZ0wRDwhH6xsCqlRlMWSSDP7dg8/vBtcl+WwIfa/h85
yg99DpqqV5H/y0peu7O33dJHLRSt9lVQHD/P0ZpP3iFWU9ObyXjifJjOdWmweGEowHRLOC3WJL8g
w02OuCyzfXH0mtbHRx6TS5K2pJwYysndGLIx11wtAtmaG7t3VBEN5xf680XmmgLfQkm/8+6DT76I
jrzph+oOJ/xdzY6gmCQM7cEfpoDXJTpCUsB5m3Ui0qPKH/yYvrbfuQ3Mqr5vW0M9qCk2+PBF7ihp
1PnAuUo6sAtiujoI3jRzbt7maybSTIcgPOKtMFisYsizZoDAhS/Cbfq/zhLuiOkWN1r2QvyDjKNs
fkhjsvPsuAiGtoAaedplS3R2i6zfun1VTj1G+SdyOZJ4UN7utoFiN6t0WOwL6xR4kfUvjFzg1h/L
sZOJyrBQx/cXLrS1sxrh9dzVXcMn0QE/HI+HoZ+FP1+scfvklS2mZXoes04o+suX5UGDs+gHwh3/
+hujdGMwQTcMdzrNxC3N363h73QbPAtrccdDzll0IJk1Z30wxJFkotAak/xCcIj4nbCYXsy+dqRp
kR84KiniOVMz8T9GIW+8j3SuQtfLsCNlPekPc6j2MmjwiRW+A4TR6Ea0HyVgSAZsyvxgvdQp2vCR
hdW2fqO4dpp5XxxE+dGfrkGeR3F0bTywpPR0MnG0srXXQBKAo+LsMMNRINKVAZQbHoYJhnKlpzXF
xFPG2cW5VTsWI3zelslfYbqn3LdRof6H8S5W2iZaFxxSTrsHBPxP8BxwGD2U130zycsaFCcwmRz+
j7FeO+t2CCPYmdSFQ8CX9a7pN9jDZ+VjCQh2Pz/VnQNaWwRM2u/jU6qqfgRQY/KVncnXZ58r3ptk
JO64JjLi/kS5Z/kN+A1F1SptDaZ6bCtdMv12NMTPPGIR7otd8z890P4jJ8HFNPxKR46d7y+bUicS
bKHAWz9f+S7DR5fpTFkxOMQGNWE9KFxJFlaN2G+2TIJVWWI/K+gjSP50BipXxI7fbFP+zalJtOQC
XP/riNGItfzsH0VUWn69xkBWy/xQSk26k5xtnu4RBlJ8pUYpZcGwRJZ50ejnoOHNSJbBQUAaL3US
X2Sjmzdh19RgIJPNKrZWYvVHKYIncbebMQ69XG5kAbahHltky//X49gGpdtG34H+rUZNThup06hx
OPC43+C8RAeYTaWVZLGwl49Djb/W55TEhdjViMWtwt2LqHWNBuuihHzqsx82PvAiOWvJ5tIFZra5
QVOyGPtm1s5+s8jKzUlgWI9HMRCqMWWz2ZILESt7W3UQmVUvhR7v2uH50e7jPaiYMqikl9FHdLT6
d+v4CLwduD3PAcu74lpLouGFNMDWySwty8PKPKkMgHppcvlO8S5GPUiP2gYEiUL2WlYGIroxMIZJ
dNtC9EJARSxd1YLdDRH4P4bsRBVA5WzUGkZLPcTuCeFhHB28e6PJlzmuxjC+Rh/gQpJP/FMjsNlN
/BuLHe7B6hkDEgjgy01frFFGQMs0kdXjWuWj4g6YErZ8uP7FHtEP+XkhOHyxkLwnSKXdx0uiQeqF
cWrvI9BLb7Aj3N+jStlBOowYj+UTtrrG0CY0FzFz0Ua1bOJUQqSRvjJVxWXAk926WnYm6VjUcOBY
O47lnzazm0p2phAZW2RkOiwvdQCnEAPBW39pLOK4dbC3UL7Ke6oPxK4VlmLElUAEnOWi6CT2emHX
paVzMqgsDSxfl+h+v22byXlsXHThWR+dl0uANn1RqEWcWtN/IA5Byz33PaxJMcFaHiSdbTMxqSFj
NkJFeUJ5nfUEM/pjYUgzajPxFHe6jcva3ALlcjQmarog0eq3TYy6bGXm2Vg/jIzakylvpQQZUPsi
JzvN64lxJvLrFcCdo+907AKHb0iqFp3oiIRNhS2726WSuSceN7lB/h7RiaunlncTkP4GvAzxvPfJ
e+NR6Jc3dxBjzZd+yTjNcpzeQxqBy10Ho8/tLKHacQfcGScJhYsffjPzjREnTpdkKKb1y3ulpNma
aQSGBuclUFPZ3eZU6cDzwHjHyv3IBKQcaylv8TQR4014NtZyiOYo0FSom3bEC4Y05OH78VlwHSaK
5htyAA7F6mm7/K70v25sce+nALGKuLJo99FrRIeI6xc3WWFw9ik32ZTw8QOuVJCS6sjI4zA9VGea
MF+Rx3BvC/GadI0Pe7wYD9cwoFX6D2isClduU2HFmhrEDaxylA1NQ97NQiqzdC+9iur07ooDkxjS
7aPcFGggRznUep9+gjaUWeYRM2S9fqoDAfUqQtoW+y8WeHuju+iPcT98FCVYA2n2eHNlmif7Fo08
kscPG0imHj3QIXbO+yscOx8/CFA+YNg+wgqbBXryYdnHh4g+xQ9HDkPm52U+DYsM5TaSdbe0+1II
qOjFLMGGFCCummQoxiNYhLDJTutaPsynVuf5j/FZ4trDjz8pbnea2YPNf+lb6j9Pl4Ee4Wj2SUzn
N7K47W/ZGUpmkPUYSvMOryXmMFrpkUQyDNuUjC6AgXTywcc0cqT2+hxC3wtQIfvGIEEo2KSRUbrO
6zipyH0re9xkItu33SVkEXfGK70ldls0iXNOqtAPhBsL/UObvAR09vrz7purLSU86K+tVOSqt5Eg
2RoCvrChozq5asGs3WzM9N4yZM+LpU5rwssU01DEytNtdEYAo6XSeJek8Mb9yEiWlyGnBlyULQ5H
rlJm3UhpfDUiPHzLOn/Zur8Crl6iWpq0JW57sSpXnLS6Sw60Yeq8dxHlXBdcHuw5erTTYG5GUt+3
oFcI1mI+XAzKR3pjHCFtgiLI705CLSw1dSoz9q4g4A6whP1PzKhvImJsfnbWaixUDseUK1ThnPda
z+xYdkLfX40K2g124cbJZwq1f+/waYX29wEBTjRpTzscH4S7kIs5r0D6aQnWzzB1Ff2Lbys1Yhmg
g24xjqZOP4mr6nXBqtnGlW4V6ODTd2UJ4QIOX7+sDMbNNXauQjNA3se7pwHPWw12cRZiFr4G8u2m
DWypVnWCVJSChneM0wBrIGjHjQHXZ9R34U/31AkNJjWsqxRQUJs1mqNCt0570oswHH7rmUU2E0Gq
r+SPoNYDaEsfnqZcD0yn+LCcL83xZ9M2WIXC4ue1Z6NmBLEd6QXGKF71Q/clAi0kZwx3btUC0M3R
YGKAnPNAjANzM+9s5IU4pMC3aNH1/rHEvsylAF6clLeggCT5jafDjlWmKuc6wL5biQfsRhmSAt9m
JSLaczT3BrLsC6jH0jaQKzqFLLfx8NkCEb41twcje1osgo5sHVvtst5vFwrm/Uef40OovW+QMx8r
D7sfc4YAKSc1+l2Kr6dTv2NHYIr61E06iTqA8AbKYrxPWSA52drVX1Bhglwji3qlDL6y206gWzdC
T7MSutDR2+Wzor9ptfM7fyn5Gl7K/f+G7w40JHy8Jzc4y+4IH6qmDNnIb1SypgddNTg2A3cB+NXq
uqmpRMJouIrf/J4/ZYPyvDJA0zlscnj8gFkJlGkKY3KvFpVzCRyv7u+z+Yi+eOIRoSbi4n+6TUgb
lMaJuejq9okC5k7Faw3Fd/QSAfRdH1YV26gHmUEBSUvRqKt9dSxnJrBOapxnG1Tary+HzypeJ+s4
9i9EQ3X4V03KSQBJFbflqEuIwovwuQ/OPGvr1htWRSEv6CO+/FSvS+gRw3sbWpvpzbHGHtCJcjl1
Q6SbqyKkevGtpNc9v7pyqRDJllC21NUVW9uMdEJCFBN2qZ8+Xe7RDXnmzVcHAXIMoQAmfcQN4l56
om2hlz0DI75sQHoNSt0jz3aw6ReLUxpnLSuxWYNz47Opgl80mYNV6iN06jCPaVvMK9BlLcJyrymm
VN05FMQimkrP86gPvpq3LQGg7disKtrOKGji8v/iqWXc4cHes6pFP8f6o6XbK/ah6lbnQH1ElyyJ
wReXI8Js0YGvH/0szqPdQl9RcnUhdac4T4AgqFeYloq6WT2p7iEOHbuwhR5ROIarOCxAj1c4Mdqj
kvMWWzop6ta2nX++Do/Aakraf6z5ppAS4eOeuw16oHfHcMVjuR7IWkNQbOlei2WPAPiAUqX8sSEJ
bU4IADwxvapE8bQojMnjC/WKSWuyKy3jR/SekLzByWaCm1b0s6L83vRDGFDOQpCjQ/Wxi2u6Oevm
CvgolERIY6AaR7Z84iIXIRjJpa8JfNkIzG6+d4l/KDwxFMd4u06MjjhG0bkzrrqzD+9HN97KkSpO
zwIVrTMPk44s0/nJNU5kErI/AmAGVYYqPVuR28PU+oWlooQLyvEIFTUzmUKPizCvB9HX9Jrgjudx
GVLPXeoOpOyZ5LAULblwOu8mFHnAMIRU484r54fFnPFvl8cKzgraEvii4Gdviw9VFKAFdVDQO0mA
noLH0cjETnIdaa8WC6mmEBvVzaQLLq9jM3xm+LQTqx04wuH5mS8gt1TpV/PMKzLBpe51UWEeQldG
nu5QksLCoQ6GRY2+dNzdco23d2Q+GC/fYK6wKTvnswW3Mq1iUHIjYeLRKMsRRE+KeOdafSu1Tx8G
Gl3k71SP03zYrbYH8Hq4LQlTHVc5Gt67w1Eyz2EtcKy3fndSI+SDlTGa6+qjxLD6rq89oOmo5EqS
qqg+fIoIVMftVTpY+qCBLMtg89JyqYRVgFMp647cYxMQMkmAs3rSvbJak6MseBBHGM7oBvmYJTEo
xct5M80NKDbEUpbikjx+bBMvUryYsBVpJ/N6gsi5D7HWOcpI+8fLJWezlw+0R5KD/h5izYhCK2Du
6cnsmgpdxqZ6467sizSvw4PxpGn/K90zvyZIANuIgZDP5RktVH5biG7j7zb5Mm2i2xg19i3mz1Av
l6oZfV7s/vIR/GTYmhLUgNLqRuiU152hrg5QpiJB+ikoMQRnC59OuwR+Gs7gcFEtTCkiyV65bCxG
2lm9C3AkP1Eh53bh580Hg3hmLt8lwvum3Cl2TBbFYaflVu9rLEr8s9r0dM2W/fe2Bz9MvRMMolsm
ZSJmcXhKqbG7QF/rSrDOk/qDTWC6SCNZzv7oX0hXEJg5d67BjF1W89JWnGyN1sY8+RGAmtLNc64J
Y8sRzqjYYDBNosqY40W/n7RPjVU3+qjIQyb3Mxjdywh/p23zT7IdH9gXAuqkqeqplLq0t6WA8Wrk
j4Xr6kGq9wMdwuGnDXBV4TLarhX+usnS/LZqZYwvpVBRsz4MMXpDLz+d7sNMYARMXKgH8sPBmQgA
rEBOhZxyMAO8nGMILcCG6b5dFZPaFoYUHEdrAfFybp8M7WVqOqTl0lmoi+4eDfh+qORD+tChE16e
nAXT6PLK2KtDxsDcg0ih6u195XDxxupQhNSub74pv2CCpw12l4dcIQws7YFtqx+kKmXNN4X5y+BV
bY7N1gqbQQRYPMsTZEWm1YiFN7a6Oi/b34lC547lJCgc3wlmyn9VjUBe+xbJRjJBhx6gRak0teQZ
BwH5B3YQErra0wiwKDI8vaIR9LWQb9cE3EuTa6vfgEVpGIJGv/z7HevazW376g46H6+corGcVH3j
5JPTG5UtQhQiJH+SCWKW4kIniBCA9wBs3PmYVvjtyVtxndH+XRuh7yzQOPETNqMisRGCezeNPv2n
znBs3xk6ugRxw7gR4vWHAEs/rta7PQG5zJCa8zvOcK/mWAbjizYlKIV8JS7pdFduDImXYe874sDI
6NjR4FBjv2tCYQEm8pcoNymJ+I5X6x70wN57p7z6zsUbS7SurMGAeSoJfhHzJ+AiAkBfoxy9KgPK
uE49hqO9Xg90ppP9IBEiyKsOB0bBZifclRx/GPsfscDzLTnRi0RLn/pehoLz26UJJFbvtes5zy70
UJ8qd6GEYK7ytVIIgU9HNf2D6qHQ3BiLYTmonCuhpwfX0xfDSZ1iCT2N2HfPt1w0VNtAHpIKI9DE
ASsJvohErKHp1xjXlNFflzCZLD/H7jFkQoFhqK4FBvJkHHDg3MryZ3tn+N3DmCPg6YaQCt6bxqV7
6FGFOy3IfSHEtnnwYNZj4X/AVzGO2e6Ae2yonqeMzcMQeBQl6ceK9f78VJqov4/Qr7G1zPwaJmvK
qHaBT5vflkApBAyuWaIsQ2f1Bwt+H17IuPAOWTSOiavjoHIJ3digtbvwZg4L3dG7OWiaHbWtPfVY
Se+iCTTqpEXr8+0kdNTOABbRmLoWEyJ7R5/0j9KhxeNHBk9/n1g3jDH3suXwUV0y39lunvgXOS3x
It2K1I3yFE/WsHb//8hkVDwFZoIv+UaGj+hNQc6GrIor/Y9IcuwahY31UyDHnCFreFRKzO59e01Y
p/1eeblhsfOmS4Di6VgSqT4gV+tjVruuFbu+lBoiz57Ei2BtQPosvYzZc8Y8ACP4ku5cBeMRLlTl
hEk8auyGH9asiOj7C8YO4K6uiZoZEKlG7plb/KgKKlTqeSK7k4u8D4UcZeaBhNMdD27mMFnCWMlF
nbiQU1FiseoPJEeFIqa+hVE3marzdWH/4p2Td6teXD52DN0I3vF5IWwv+8rYM5eFiO9HN3z3GYl8
EZHBhIGpmVcYQJOznVQyFRR4GGX+5Q9Gn5BKgZk3a5Fg8zNZYRoeid6Q1/jItynOiqz4IBFpaOEt
EkJyN7Hw2tFjX2rr776qns0BxIRjdg6M1oxBLDRnWQ5dXT0zuTuuBaP+udGWc25TYTQc5QJTgxnq
Htrup8nEFDcJhcHSRNvh1Jdo6g40UKPM2AeD52Mwuy0BUNquIMOI61wi6ytnLuGPOhOd2BrwjIDT
B9gg7Y7VT2GIjyVSH2Pu8IDvg/wJVwuyzW/ZUVzKOSsRwlKB9Qln+FS/pNln3Ith4tfIgEcOGvE9
SZj18qLdpkhyxZ0JTStXkNiHemaN93bbdjuE77N2uLkNEJEZIk4PSAiZqd12dRqjYfgpNNFvnqYL
6EudDG/6+Hjy5JcoIf4EJEajapODfzYRjskKl15ATpcihkFPnsTQaLBA8GWYrsrKi3qndcX8Txy/
dvX5FjzUmkxDmzeCUaKqmm9fMuy/LUGJ7yv+3q+l2n2p+8F3RiroegL8o6iREe2I9F95vtqam3UV
JvNelYLrqDR8j29lGg9c8y0qvZdj6vvUarNHKzz+6Xr5zLmPHkWQXuhU/ucTdatUxhkKGtRCxEgK
SJI28S9hIeosL8YoGHFLRh0dlR+ZDnA3JnJg99N9LJd3tR1+FTdyWhGXKnO2HZHScTjqpDrGaTzx
/0u84FKaBsjvb7WZGfwhz3wVSrURjd1vwUap/c219zMeAqCWEFl5gPThfWLutod9N/ib8+8mIJSd
sFXwN4nu5vVCBe2H7+FhE5ZSgJ3nbD7B3+2DIwbEthW1nqsG6Ifz3e4YB0D/VEfl/6eOsXV0M0+6
fkqykUICfibdyHwqT0i+/l8DeLZCw+9OF5ql0m7EtKU2P8yGL+WEpg7to1PjXQPESOPFSUD2i8A8
wLC5HFbmQeYF1gZlmvPWn1/4VhKnq6URnsc9U1tMvHiylaEQVQSS5cDSk8sBZe9NQgeksysh5iNE
9F293dp8Jn+DNhHNW6ziipgsKl3ntcJ49vi4qmnhOLR4X650PFQ0DfHw0u9NguH1bcw2Veqsjb/q
hGN5h/HC8LW6jJ31BJZ2zOQIzUpBxRy91SxbQcXkWbBaYS2Sx7rzncg+OVoXlz0Hsre25N4lkOIi
Yu39vGcD78Fwj/jBKefWeYZzmmmJ0co6LClbWNJWCgXY7HVScUpus4aI4ZJ5Wb9zXf4HySS90bWi
t4+ZpWQiKLpHSTUJ/KXARI332+5q8CU1Al977bvCExjzxpLzGQykTMPA39c5cncH65HQErd3PNzc
UtT3/Im1M84+gQFc3aydvKpUxzNPaYi66UYvS7dW8yN89xVUwSRrZ/RnQrw9aoUBUwGeIKb5GpiZ
fJTgUg5J6+lyJf4xualiWix6ET38uwU6iEPwUJzfF0oAyuyWawqABXXU+KRsvSulFBZ/fIBjQoXG
Ajj2YKKMTVVbQzGYAaZwTcj1SkGuyVpXF46wJmbKbTtze9yyhYvjoVs7+UTikI4GbQlI+5L5jcRg
OLOH4uil3401aXGXFvALesZKqx1oAKB08LhpMlhkFZyfBUq6ybRU2ewe9S3lIFcrn87TBP5wJ7Fb
HJ1UF/pk63Wx3ijD3n/oUuoYZRYAyunjD/9vExBxpyeLK5pOe0xp+7o4XucJEWM+DBNrYshsoOPa
SAgZ4+7biwE24P0rOcHtd5scTzbgOW+Ba1CFYg5/brCLNYKz5guZ+5x9bHH8O9jwGyUS7W5NhQKo
kpHcgRniFX9/YbflnY25MnpHU1kV7GprrkR7S6D2YuLytyUru/f1EgZ7XQPRQ9icEZhU9peO6Y44
LKDI9V9ujlN7EZMLISx4hnskKdvjIxxavlos4HVC0G02Ly4rzwh4VC8BFmm1XuE83V3SKoKs8DN+
uHYMfm6qybDw4iQyslmHFs+GUw8hUmDGzzeey+wNsXdR//qhoG4md3Q13V5m0stOQP/hB0hfJGMw
GTiVMHO5R/e9lAJY2PNq2OgtaJ4gSfFstRfhOVcjiMzk1tfDTrRRFDUObVWUOyp1IsdYjfWXwtWf
chvFH2vV9AkUzJqKV/VhdznhtguLitQVWgx+8yDFuvkhlhqIRyru5Fo2l3sCVyECdXWf3S+Rx3oF
wVN0xSXsquXt5oIyi2fAwzf52FaJftHrdIevh2RsU1qRr61SuO1nF/74MElheWxorkqhPiVftmET
HFY4pMbGJ3u4568aUkaB1/oV7elaD32E6FwcdYl6JeBbE3K89lxngpUiYDbBLutMh8wCDJjLtVDy
Co15YdIRNHssAPzuAR7MCh0j55KVpb1uKEa4jRbwOeASV9eXPKRgEE+kvqh3EcbuFS2cZPCuUIkp
DHih8geu6JMjluhFbFJaRoXDJ+hTz/pzOimaJ4uCsD7Gmd1xJA8zPuMB1pbvwQiODrtZPxGlt7S/
MlBV7A2VgXcM+TTkGHsKTrcn57UnDsaE0zCdWY+9PyA7RSRw2LH3frKNa/WngD4CwKKhIpajc83v
qjcTdzDp958Vnon3XtUGhMJVpyair7Zmq/jMsBlYOq71Km7UHY/YBbWN2n6AuBg3TYugHHhD9SGb
MRU+JTX8V6/v1Il8gZHdr9uTFE147mmgizPsBUYkCRAcswFOV80gdTF1SvG2aoiGnM2gL+5Mwa0u
BeKS99JTe78+lp7qhiAs4T0Aqn7vB/gOkVv+5I1UYkmvG7TO7t/BpwmThsMpzHS3SZkdJrpBMl22
c7rjCkGN232RLP/9QjLn317Z4H2IkRnx5HG63l59VpfRhKeOSFzewfx8uFGU9CC/DNeRk2Fe0Me3
DEy+jh97TSU1QmX7gYX+hHRoKf5AahIUy4/d8h4a0Trds4Y0SvHFsLnfDR/2M+TZNweOTD90JFSa
eNsRHflWev0kk3aMTIse6gT/PhBLPi68SLgF869s2I00jmDsLQ1P7SM5XQzP1jYUUD8MOctOhJGP
k5TwH86iiv+A8F0023eJXUWervo/HmJBN3xWSDDwHb4gqSMNBEWOz4BHaBa30FP2k/Sx9IOpIa6T
QvP9HUrh8aE1k0PR0ZfecLSOg/MQo9jHdUZ7smIUKu6SYBjU5GqRsf/sNCEXG1VDczgS+/lg+YeN
ybOlCUNT7HsVbgRPy8fTI01U8kxmhlDoc9CU8/IowV5/8UAh6TpUQSNhQeuGRdQDRWnhSCV7CfBQ
Vq14BdNuqL8zdACVazWrhWhoRR1AtkE8rc1jlGAdZUaFLg2OKvyh7QDq4jry/XNAX4QQyFcyhtQ5
6uxxizJMXt3Amq4rOMYk8C2MdKDRYZ8fDSuxLoghdrfqRdJHdP2zGnkmZ2weia3MxrJdJKQxZNn7
NKLFLlaLbm1oPyP7UiUlzGTNvhUQ8oLmZJBMdjgwpv+3ejDvQdaCkdXXc1J/5CU35cEyyEQah7Yl
FUg45Wo8SPwHkMSn9XmSH8vHrJ4JJ16sZP3eMNjCCdrOp2l6hZFJWLuoI+YPvLE1jVuJWgUZv3V9
H/Vw6yGRcNquRkSQN21OOIyplFJ/doQDRW9PnRI2ogIXY9L2EXJW8YReafQFZfsnlwfGqGd0Wl/C
W/QaeTWu2LuATwSW8XyK9OjvlWpvgr8jLEwZ7lh9S0Q3SR+3aWmePUE9YkHQRZHUiYxBEqBdp4nO
A/ZmnV7p8xd6Z/xeIhHHRqb9oyHc87Z5Pefdt6dAOvLfYvFIRkMCeD3eGROlkE0FaL5e2SqJfok+
YX8uYg+VzvSg8CFyUpywH/vkxlPZbbOpX/+eT/79uLHl5MAeyO9+7n5LaBNsDlkkZT1EzYe6wnIl
FO/SDuicIVVxQYIZnmqvhuuuHvOFPG/S0JwvckSgwPeolG6c/LY5YsTd1a45Aa4bYmfb2AoLLXtk
LZC1FW+5SUiIHTFMFaimYniPR3bdpns3vrXNme7C3EODOawyHyfqgOaxMT3yQvr97NrkHb0Oo92x
Go8BPxFz6XQ54BWRMTlBJn9jzziYgxxkMLZCoqG/rhsuzVYwcNAjosGXZrKWYe2LEuZZAS/c3B1/
4sZ/uzP51uEqwHV6V2EDseXr4lPQAyEZaV34vgsvIjE87FxT8gr21YnL2FSJ96eAXuFyWkar6eMW
gSlL13UFdtSYjSFgWSjPofptBBMnKa8Fi9IDoyTmUOutKAPnNSi1Sc6fj0RHyPPYuDFP68rVWhyp
IPvrlTzf+TFaKPgj0unZWPgOP4CQyrp1+PDONToIU2tCVt6zEQiux+zAGeC7dRGvRIbepetsmtpZ
stmJv/U6cOl6kHx+B84rGTwggL8HDL/mdMdlm5UINdi9diqf1aeFYHvZLaUZ2pgMV+rNyru9bn+U
wbKIEfnkiHcUpO9WPfvqjwKuMIWxYR9hJmoveeeMi1g2IYkFhMS6N7pwsRv3tFtHCxOLj6w0JvOf
2TiRPVzjBvmwtynsmZUXO+ji65GOtzbPMBxfpLHFgSHI5EDlJqbJYLFBOrg3CsfNOrRLkOIjzRQ4
uQ0kqG7aS2yc/EGiBUXjySC3lSSnuXFJT0+/X9r2ywsUrHmQxZFIgl+kM5eNX6upR8YmEd2dRlg2
DzGXMMTRaIfzV2NPMKH3k5bpXFZ+qeC2oiOX3PaoN8rkHGjjy6ieSTpKWsiGQLqaD0Ew4UPTWBK5
BoyCtdTxIjcRd02G1ukULtvtdhcytIsbUhrgCGnprd/f1he/4L0NUZNzwGcytLqTGxrPqy8Xe6Qn
6pd4vmerUwb98K66ihNLhBQq9TvuhnWkVXQq9uNyTd7m5jrshLhKbxKQ7849yM5AFpG7Zb+jaXJv
IVERHQ2NYLY2uiCvoukFGRfRFATIL+kUqOGOJ2RzfMji1VATIOM4R7SiV314zayPrj8+x7C7Y15f
uNmwRa2QFuNGeSTlh0LkxvKrsrExA7Ob+LVJOt/9lXikgFNMpWtC7AXXyqLS3I74C4HGkBaKF+Vl
bS6H2Y/Yc2zXidoCX7ZLOYBtF/XRiFTrBGMWS6bq0X/jnhBg45g+Hr6lgstq/zIBp5Cbdtj1h0jh
d1xNckH0VASW7FxOmefLeKlHMZDAShKAYrU1BtJtekl08GAqna8+hLKxR5md3jzhgNtyxNhtedjs
fgOX7TSON7f7kpwbnHMY54zAyDrzRoPwInzPSOH7kZ+48oyC+ugG6xkmppaMUYrQ/AoSdyskfR+h
GTMeZIU3n5bbLjHLyLjdTvK+nsfnUg0f+j8K/5TJRJ1e16psFx5myZzngcFH3OyV+7RuGzpxbVsF
O/pfEB0o6mbdQyAl6RWPlRothSQUbGseDvXyqQwEDD4b6u/UZW401gCTK1H0q6LFUlodj2Wvueu5
CwZbmFH1G9bUgZoIFQxTmo3CBC4Io6P/V0SHWnjdWSmL/db3tYZgS1v4VsRgI7E2qxhEUhJ4x0aE
1kV0yO9brXiIliUaq+bKXrryTeNyvb2H9QQ8FYdIgEx2CYP5EnFPic1l4GBFD+EGakPsZ8GbEhbd
SVPVXK1XY9QnifdulC9ujBdH21kU/VnJt+M13VCOMCTfVNOWG5jw5XrqEyURhPFZdsDyFoxnPkjU
/iGh7NDcox6SuDhp1nbtEZOLWtNRCY2nFwG/A7ZYrP4p5cafC2zoigva8SqyMlWWJPaDEOyecHLO
bcXSbXZ+MqpPe7DR00Ns2HNuylXG9+Ju9t0KwedCnCiKfas7AnbPm4nQ9cHTlbelX7P2TVzpzNeP
IgvsnyMKLRoKf4FOuu+KoWvR/9BlhgZCAufydQf6LksnpLGIPQY5i+i2uJKmSBxcV0V19v63/W1n
7LHZrCT3pmbt2qTyipDyW/YKGZBBVo8r7jzPAq6GDB9V0/ZOTwgpbI0/JL7oM2HtCIZXZYltWGcj
oTLtG5PCjBEVSbX1uBenvuV6unOfgcbJeDbI2g8Fh8z3pg/sXqRC9kNzmYQJdI17pgjdwSxXlZrp
Cz3D2qnKKpaX4gcuqjTUKWpFKXdysAA9LLynyXj6qYprmT7QW3I4Igtj45yDZvzqeLzRlV+clzY3
TJwOaNLnwtl/Wj921tCUifEbmPwtNxsCPTrGRB5eAc99amgv6ajrb6EYiudwzlsvevdKAwzpYJzb
v/Hyrd3CVsCbGT+Ge/dE3fM+qm+Xd+9l+RbmCwbNP+lz6QKnk6EQtlcjHX41B079Jk+rYrWtOXxJ
C9wgNbRP04tO2BjNu5afybLviSrQBoZcCM6WR8TQ0RPYa0OPU3DCPrMhmjq9YMINYE7RtpuZd58t
vM7YxeeICW53onAx2uHnUZ391mn0xfJ9YCVFLOHDwXp2Bz0e5WrEhRen2cuGY8Jodi+HcIyVSWCX
SlYS7UBWsUE57AD1bHgG4DQQcsW3dtHoVqDJBD6IG/v7tOHM9y4zOwWuWg5NHsMit/Bg2O6qBflu
pUFA/998lObM/trWkS5z0+CLDem6qW6w7Elobh+DlNUxKRsbmdc9CRd8ay+P5h/d9ujK/X5F6SS9
RBECstxWQWiXvEtabLCCt4jF4/lyiZX9cpxI4EqFw3lk9y2Q/NZWaplSg3QHJL1QM/7wsQ9ep0yQ
w9/xOcmfXv87E3bXXoXw6PLuEd8s65PJeaPjkmU0PYNsUlYd2ufabXNsbSl7sgFfN6fPSoNFYVEB
35QPaRpIQq+UKumW0B1ox+mV/dZWxcw1flK9a1j7KPhO2C2IzvJrBXYtlxS2WEjzP8RLAYT1y5JS
5ajuPIlgT6Q9R8dY/0LqkSiB0kC3FoKCUfpIOr4LuXdAo1S9YUfJggmp1qcbCjO/U2nzZ4rmdV1d
4EKgCvRKsoiZJE+yWXC/LNzD299C3J3lIXDhjAavFhk5AYlydWGK3LCzASGzHI4HhBAUeh2ViUF1
ahZU+mIH9Opf23VwvLAUw4fuk0PJnQ9e6+ClAhm+xV6LNt+NqLlfU0BjoqUYcgCjK1C9SXYr5jER
lHNtDtzou0B7NPAKlKWb1ktlZa1narLTdZqsfNur9n7aAcK97fMuuGljIeBAJ+mawI8ly5LB7OQp
m0nGZ68GNH78zztlZOctkyJ9sltxxcvclQt7V34bYc2Ar+qW4yJX1D+84yhvJe+uigsNe9P1SkaL
Zy2Oz/tTpnCSKHdB+H9GXbaIB4otNA6iBQDI/8AD0r/j4Hk6x43oUHtqWPtT5mIS981fznkcoT60
/UuorXS9+66rr1mF7ffafuxz6AdEdtJt3vsp2Ftm7dzgPjm7IfyTuVvTjPJpj1MCYul+8TzZcQTp
buIeBbIZIAqKBDpK+EH/alOsPNIVLkOJA773AVjjOEbAzdEQFaOX0EOTrOy6oPCYNAu9orIpJLYi
8s89DVc4qO6GELXg3+Ep8Xxn4zKg3RGWAnm/yRk5sEeyWS8xW5NXodk0P2KZwYp5344XpOaMjMVh
sg/rC2hKScMRZmV3AeNZOfRZW6veSeLKvJ+LV8QR6OObGXGNFIefvZi1hw+Mi6UgI9diUrbyL+vM
SmDqc32t57zTDVRMljTVOVE3119lKFpgGs5rflXGU5fQg2aMyl6ThFfpQr4jXjrYX4+0LnXcqJbf
TpYfXiEqnrisYCoGqaK0ZhpPRRiEetYS78SACIlUyLospYiaQuJ0Xnc8eN6leApABXC8zvchLLIi
BSTv4NEysE+PARTiWZpPUIl53HVUQle1IrVwK/l6xH8Y6AcclHy7Vf0CmbqZ/yrQ+pKupY59p+z2
gZUZ+5o8hX+y9Pj2bmCQ7T9K9QY5/w4l/MNTmb0nQEmSbsei6IizC39TiC265LtjrdR/Cq+MzD/5
7+E8XYXZjBxYr/yJMjogzq/wnYnyrtwK9FNxDbPXxjPx+owyxrC1AqyJfZyEvsYLJQiaP+hq5vtQ
O9CN1kcp4fBSU/OFjQ1vuCVQ8BX1tQ9myQndxeRwKineeNQl8d6DVD/V+zOV6HcYVcu/GhXHbvJ+
8HohzBRroXjy1NBokAcedDklNOZdK693IeGDoYtUWMx3dqL2KdaA3h4Md7s6iEVRvzZxqjkhcV0o
u9j3/tft+TywetW7DldyevdI7Jsw8dUTHL4O+liVwVsXMksoxzINa/1bXHwh/v1cHPR3nwNYMyAJ
6PU/YdMtvdRfmz0l5O9pCzXzTTIJgb1XX/ATRTn4NKqsalsN9dEYBDIBop5WZXfk950l97CpPZ6k
vttKBb5LvxFkVp1pJhl27gBYoE2ojTjiVslR4g/gG76Z6NeyNR54wrt6RJ4uuDHBfwSVz1DdH3tU
jrYaDSTKFY2QZv0F6VfGUhzQUksGp3XwNf51BXr02+CRxwGdxtxz2Igc6XV9d0j1KXBmqSyWTzNY
0rP5mwPVtxWEonf8bkZmsIW30daog8QfhuHdIPPCqEURrVlwDGjgQHvzL+aP6FDOsLjY4lNVEhSP
6hwlBX5nLeKX+rHuu1Hd73KNAUqtcHLGoQmfiCUKbB6cDNHgfiFzv2B/HOlkpl00GFTcR8HrnWXf
XYDG7/2gWe19NJFW0P9pdQRJyhkIXgQhtHy++repwsjCcZ6UD8bXSAe1lKwL+6aFz0Rs+5+Uopts
aJth2gRFR/Q+3I+YXLKo4oRpxmbNyu/TigHq1HVBm1Qx8nY7hS7zXR6T3C75Ai4SM8BLmRNYRjct
WOqt7nk68zlXcO9Yiaw+XD7CnY8cRxN+lkCWwMeTwSvrxGgJ+xuu9PFsSZJbkJDhXPr2NohKPBxe
XgF/JeWAOVbo5Pv7AF4TDIQhvQPBJnv1KBBWUTXk40NuBii9dy6WYCRz828yswImEZg6uGD24KPw
W1l+AgDZqA4ODVeDHtd6CNIoydptPGisO2bALcPzQSrUHxQoS1ImNqLNEE/OKNki8nX0FLP+naFe
mZXQc7uOuRIPJVTyC93Rn8Vh05SWJRsd2lcvdneN5rdzVOWiNGDVT3XneUTWk77E+d4TjhYyVGDL
MxOsL+X+lPuLH3AJTR8L7VN1VVUS2U35LREDHuB3/5wy+Drhqq3uhejyW/GsGbKFvKiJuo15KhR1
LwFhkIoq9rIAll20ZKCd1yeFH65cWhKSs3yt5v3IvhTBr05iJrxyiHn7I2EQQnfGfBxZKjbV2o/W
ww90ob0qDEMW01TC8dCkqdnvxVtNjn+0mjYPnX/Hn8GGkzkGy76FjLGGD6PytaEIerKEWBSiEtkm
8FeRUls8SDQxDLAVGlRE847TIAPfBQnwH/ZE3HuYfAI8XVUzGkAT7Tbw0RLZ3npheT1w1sZo0yYo
dQnS6IJSXF4WRHB0zaAZzb7s6BJGx4i+iGcCUN1aT/YpyQeLJjY1gAtXndTgOv91n/v+lbgJlra1
zs7Sxh1+TNR4DojPl78lz2tx71OcrNDa5rUdMD9wmScyF4TwJBbOQ6GjhdRqvqYgFd7LV6BZ04sq
oGRNpZd+XX2q7i/R2fv4mSiDGObfZPu0kZBjMGbbh7iQZAotzMeTKtTW1D6lVux99agalyYU4srk
KcBTjdP53gjfbDM3iP9mUCmOSZI8p2o6ohDmtFFUIu97PZCANA4ESz3SeP+SFZnXs5Trd6rtwagV
frxoXtg3RlXfp1OvmDmcPx7pg63iob8c/xO8sLOtm0MphR5nYh52OGYFIGyDAG1k0Bk2BOkJDGMI
l238nuKnuV8gsXSXxBwasqEsjv/QMLDq+ydbWnxTBI35eRR3HQi3nK3N/BN1B0pI+CpKj9VXkCmx
qIgIoyZGrb7E0g4WA7fvdOIDKq/0OK2enl9i/DMmYgYyeewCxquKNbqOuQCEScrdalnqYZeTqJ8r
k6IWcPzq/27JLqSXIR97icTqkC2BnuCYgye9pqvNgq7l7iJM/d6X5NIx3cVTxg8w9n42A2Trgt/v
9y3qNWr7JSanC5exl2bh0PvvWrYt19AArmBJw/mockxYeilclX3WdOw+i2ExyjwXvp3XQBhLl/lw
D7agzgmh+p3dK4V03SdcOWnKBMYdr/hX/zwj2ywUpjh4R8MDcrhV19LFDV/B9W7Q1twWrdY0tyfD
HY8PRMBBmEK2deQfQbv+T8XZye/UdaMQflKT/3BeMwC6N8Zhk9BNO8utC+kBQvJr/6v7XKLp+/Az
I4RGT/4mlLKpmTFk798r+lLyj/jJDBA8RXiCOK3WoG2Z8rYHSTuxcdYB9JFt4wAK17RT4o4ZA3kp
xMl3vDFF1pDO3eKp4+TxnpJfi76m9+lL5qqd1zy5Ikkr/NwIlZtnW36XUWHULfi4SY2J4KzN/oAY
MU5Hacft8o5mPc73/Cd3nFJYxHlLX3XxIXYNnVxu/5qTR6L7TMybfZp14oCN019NU/ygQkS95Ofn
zEvV3IAwsvX4STTcVAy4XskeQfkNhKZlBQYc0H/99osxhlw8WMqAkM8d3lWs4GKyjuQhEhTo5Xoj
Y5VRwMqSUdmGgzxx8m+84SBmMIDX68q8/lkjqELx5UExChJ0L+/mHLWmc13JSR1uu1L6ENwKLlFU
EQeI2oWEnVCQLRiEg7MY9sbTTodORiyGmVnvyhrcFtyti+NP9mLQN5sa4dwL9S6DKnZksxL0aaj1
ghjILtK92uoe22C+kugvyXE1Jex1B0YSOSyG8o6vrdIEMO4E4BHd/L9aepTRk/DnYGGXzZvfFZPN
b8XS2Xg7S4DSuddVvNlWUPgw9fj9vGJcitohkfxuVBbYui973N/JPf6yOnNKtXvk5QuGI8MuQgP3
EgB8E09Kr+BSkczUl5pq2zCoMo7QFBKO7ftjJqMk9zLg8k3cVZOXzmRuyk0Vmp0xzpu0dJHyrk1x
fmIxdxycyh97GyJkmsuEnQg7GwYoaXnAS/yoz7iLsFyIybunk1zl3gkuSUIL7JvzkuxD34QjB6ne
dwsPa7UQsiGWdXkgvZMGGSsUUp3PsxHzPZ+8RRN5gdPSrxPD2bdOYT3bk01Mw0QIKNeW7cCZEB1X
BVCFqccIC4OrHXz/j4YKFip6uxjQ1sk8ysD/3h9WbR4cb/jx3JJLS7PsThLOLk9tDo3J5hTuFmHk
2092HYRSv1AH1tDMEHeoxEF1XrAHrxBb0hauLCqnL692i6HpLrG3k9096FdvyC24GiFVoiyWxyAd
8R4KzW9EuQBOGQ5vimGwjngqauEPJsHt8GbZupmtMgOtpMq6VlUk7M8PKRHtQZDC5ITYLl5u8JoS
3pKB7rVlRuvDIuNZRKKSbJcfP+LEyUIgSqTWd7dbMDWbkfhClyRltsLUPsFDCep0Npa58dNN9mUX
KNRtQzLBP0saWGbW6qFKO/bDXJQ2NkopBT39Jnf7mdxFZ8s9USFqqO4MrmDI23bjo8gE1Nyh9IKH
0ic6vcTpnDNjDr8CoYHQuhgziJgKVprrivhn1sXGJZILX+syPpLsT5DZ7S2kwFILZwo0HRR7DIfH
x8t2Sr0puxW30mTBujN+9x4yyqb2M0r1SCFnGM//rl7W0GmKgMnuqMO10VR6aRnqUCTHsLM9laXC
QLzDKP7Mw2HggCtTYmrkwAs5RFtPGL2keHOlbKVl6ZI6HiooywJz4ygc8QKH2yECL2KoxwBtjvW6
n9uzesCjCVbkOOhaB9GSgn+oa5xuYS2zfppiXuQJdJIfLCjAtPu9FBpCfDWT+uYaI1fZJB0L5jL7
DKUX1aFSIFSqe1frJNgrAzenEEUkKdj1ReAjbhjxtaBjUnpwENdGg2a6BCCgE2ZliUHtS6p4wcAm
5a4gx2EM2FIMaujGW6KW2P602Y7huaRxCiJ+gtzI4fwdAy1vQf3UYIFZfWAS5pRZx0N0EqTvRgNB
uo0KvmB2ZtSBIoS6NxWkacIdr1SovBEssUL5l7mzdYLf231h1JD09tEPndfvmQnDqoQCbEMDSYnp
4gm0VzY0zekcDkHEVBX2MVN6mRSeog16s8uQ/R2cUtChcnwz9iAqiMYdn6IXLwNyCD/95eparMbC
1jJXnIIu9iOdKxVA/KQTF5RHFq4OXS8BYy8xtVXPtrZOBePvQNSZlwIfFqWwN/t42j09tByw1HT5
/fDL8Bv64933AXf/y7B9H2BGJZO8TegLtb1VQy30VftAHwtFzC05QzhKuihPefh8D3hsQYjZvbHH
czrCnIFABtewuckAAmWhwM1+XanTwnXwHS+IjbfgXvG67pY8qqxyDoLfNCA13rGOHnfVAJy4tm3d
NoHfnSfnVjX8KOtWeCnbv2pwCzDEQ8WjtCx6+L5kZWzg6mC5KTN3TIA4dAdfGtt5jlGSIAYg7pjr
XAFrgBxklyfwUwPr4bKReB3RjCEa12S4TF52ZAvluXuKt7rohHJ+8eRxpzGKiZyO8cyWtNJnw4Pn
DedFzUTUpDZyv7KQqRQ+rRyUoCTN+7DVwirRUNWQelcZ5/SgP8ZU2WS/B67SrSGvUYajMrDfO6q1
I8l9E9ZyUFqndKqriholuy4HsHMAHA2i2qksPO0O98WgQskdqFEeCyVg/eIzYvQaA4Q/2GiI0Ncv
/+Xe+Ss8sX26TiQWohEFaygIdOHf1VOfXCUsaGi5Lj/6XCE9yWBEP4zWXS7zJJba6Txdd9mpx8IV
p8OmxvIGz2lkY7pbN2w76Z4j+gWATlIZJt3qBKEag7oqmG8afA6YZqe/KhhmoR6iahZqge+K8qiK
7QsDh+HoM96pWEMjURgOIPlMxkc+9eda2JhUBnaqwWUUVL1SRLraF0PhqAYV2p2TudrmAd3juo76
zaerfWO5jzqOmHMjZnqrLyjXXAgqZ8+HmsP2yFHuaisQ086C15XgdYoYLxX95GArS5tMhyJLBZrl
DkAIMM4oC8DC+gnPH8J7Fyc5mvw525bTG8jIkfCQhS5PpN77ygRFy5D6OtMK7wX5L0RmYDTdrfb6
jFErpsHkpGuv7Mt3Xp4W8KP7U5db4TIlBysy+ylB0BB7RQFEVQtfDfKalPBdefXw8tELgfPBc88k
MMUqqOxn8usUVbaFz0EUyoDSZRS6YkF7GG4oxfFE2uM8LrGSy2K2GN//dM0625YTwd/TuXrcZuko
bXBmXW66cIXRFe6U6ylJ+5+xs76A0Pwa28ggQBC9+DhlgYh5XAYnxPUMnbE7ClKM7e6wCBsgQis2
QWM2oxDGpq0UcXgavvV1H3aWOC+baE04KfYHb5vvyQ9nDSXLqF+c60F3rEOh0gXxt74xxnFwSrF4
Y0v+hyaZyCw4rKoyC4lzhYA59RtogRkf0WNe07PbsfWkJQz+wqpMHC1uTxtfyIHusy0XWRaO6yZk
zT5G4zudre2V4Nk/vyYehC/DgoauFNHRMhXV4CahqEmB9QC3skfml+rSPJOEBiS4N1LNmqEZdrZm
x/BNN1J4LgrynPxFwy+85tlyXk2KemJOrAIjzemsVyOlVxKxuRCYByRv/Z4J6CQMGdic1+yqEMJI
g3nBUC66SqmnKv40ZRARP55mUf16gw0iiKrd9B6wNDQM54FB7AjAJaYRJaKbtBRQwsgFMh+WhUlt
lC54zYq1EnRvVI1yFJlnyYf68JPccGNMjXQBVNzU4ImVfLGg+uaiM2SF0BLhKLY5atq1ImQejcD+
oiQmf6sQW1Ra1SNRnVv8jzqhrPtftzOjZV2LfVsUF8/gZkM40cGopnDeq7h/EuozETkjqvg9+XD+
jMmdNtaQTMf1JI4omoSaF7kRZseuS1RXFVcYzY1meEiivTsC1kIckyVnXE4jXDG2Q5+81v416fBw
tyoYTCZ2/5DHFpn5Kjlq7L6ZXx1JVcs6Ie8a67GBU9FgOjyTvGF+3zGob6krdX8L8B45ykv+1ePR
Tj17CBv+0MS0gBryBhi7titGhERwj1s8RXrA1xrRt1Xnxum6l5QMTSj27Sw3VICBph96PYBJTLRc
vdvzhEKWpz3Smax3aHhziz9Fn1/81weHDA4Ej5YPAfwGL3Af8vsqymsKavznS/UxDgz86s7RqUZl
fN4WoQ3UDy1rtGiTH0O3XwDoN8kMHI2ig49g3j+bcTlDPerNThUAUJ4fXQhhKczffRfq3D9n11KV
7Gc9KyEH5Bh9mKD3rXAbgntIDhhUIfBbFnFmWTadRX+Pp69FajLJobOKe3BA9EZnfGFEVt8qGPvI
LhltX9ZpSRe6H22Wj+vnAnsNXKKayVlqdWyLqvFPlNfpE4gz7EV4C7vS4Truvq/MEg/yqx+pHE26
MSnOAq0ZzqcPf7oX5c0Tb7EOqUPrSBXvZE7Vr24czgnIkwPRADczwmKlrpJVJDat/vlW6C/nbusi
oFJyqCfqB9fkpYqyyVO9KYLaqPZmio3/Rh5T4Y/0VS5ZkfqDXH0MwknT2nGj/En7CPivOQy0SiZF
PUBUXp0uqeMYhX87ceCo8GjrdzFCkCVEo2KyTzn0+CrHa8u4zHc6tIh+pWZ6Vt2owYMsGl2pMkzr
BqLLmkC0eiKXRfi5a5/xKBRskC8Rj6dfd67ZhUFJPXbegqE5fU5vAurVFe6K36jlzHRsRuyu8Zl8
CvdDUWc+pmViyfdvuDFDIplUVqjqWXPOVEGYIe3YKHWN3SXpYYLHHolMVFcIHHalVXgMfKp2NAAz
z+8AgXIRTfUIMrbg5eo4GpwdGlZyLJSLMNmSfX4/xTU16JEYcLvOkBi0Lf9uFVi9JhxdPkPmiwbV
/dxht3tr63YCEFfLwO24VH+bBOQ6HLJy4b/qN4xiwsI9CAZK/3/jpSpvik2WvgJ7FI3CCao2zlFl
AFTcgH2Lq15d4+foQHGEj1YtVEyr6ZTlL83lG2mLSvtwBxe7MuAgBQmwQ3df5BRLeVYcduRqpiWF
cXn8beWHBKxoE3S0+zLL03SN8sk0SXXw+6jsYzrKfa8itJy+In7Ug4RD/UcvDr1gv3dXNhbwgQzZ
XwqVOUd/nhgXz7aI1zqHDP9ya2we47seVTNJ4Z9GlhlB9sDlM59vgkEhvoRgN/3YM4LTkDgl2lNt
ZGu0hL8lLqCXyCVBgbNIFa8TKIZ81v4DDfG+Q1znri12MFyQpBTEBnA7YRNyGHd3PA5UpG4vc5sr
CxmJFE2Xsc1KlWZ3DSw7p+j0kuvDCFY/YHF1dpumaxat32VEKirE0CMgk983UiTNLjt24f24EqvB
kr9I9IRWtUif39hCyMwksL3C3WTI+3sWdhXFXnDusZrSzE2zwoZMWqH94m7HXgHHkS3ozrwpN4uj
ouRlZVKL9BFPx/j6MqKIxhWLJhjVQmh6EFwPTAZbuMOC+ujDherz4eyq206ewGdFFavufDrR4pvk
Crvf32I8kziXh0b9iHIoJKv+3wTc2WWbTAnFDAieokTn3yg8K/noNWoBpZXimu/d6EW9hd/6wmx3
yjnVKc3vJByZVvgTOgC9I03WhfQTvVwixdz/vALQEk4xFhkuSrMbgH6hhooIVsIzG0SGRAKxcNwh
Ejz8GNwMsTz8jP2WSpXAzPQjUB/ozvLU3UTQun4LvpaLNauRBSGzSzgfS8mLAv7ayU8eq42SNgly
FjwWp5aTr5Hnq+hHIlLPnik0j4nqAKM2eJNjwlKEWxBMcX0IZwNB2D/uWJWFNgXscKL3OzPNriDK
GqdZOcFb/aCWOvPRVUoANlviR5OEjE5Knyjqyi5WijT4NNs/00XRXNmBhSrUwKYZKyLHDElJajUT
eyCqSDFrghGNcHMDGYgb1e6+MUG3NMHnYPhFU77NhPHjlNDf6FTr6EABbQqX9g0G+TjFhJKn6/R9
AJ/g8Xz2xN94X8VuNS8BKyNHFB0g4VKpPpoY7b+5RuVw+dxBSWOZ76FgPAHSSrHkqS8QbHVYcN4E
Axya+GqrqGxSrHOA45+NpCCPWt97E3Ano5Low6uY52ly8hH3/EajVzDRmKjr2x49vBwMqDwXZ8dY
4gYUxeRrcHIh8helfDVcPGZ5IdMnFbJMPnLGAusB6W322yLm5VA7p2qqyHrd1tGeet1KtqpBUGD7
2rFXO8DEqYwU+y0Mk4kQD2J9h4CL2ZAPr8pjCZo/NZ6XvyKHmVC3m2BN5mPhHTh3aM/uA/mTlzCI
iS35eXqdnKxly6ldCFLLCPetFC0CkP65t1vXgHvKMoYZ8xUbE6wS2It6NirmG0HQGH5cBHfiYOg6
Gn4hhBQYqtf6kKxHv3JT9HBuz2vwyT8STceHMkUMjYx2Q7n13qoK7SD2hRjyVjaviXY2h/qjz6z/
AhjWdboQKgpu1gThRL6qpx1+ozW0OhTDuR93YBWhIsAG9fhJp3vW8qmBPpVjCe3mSA0YyAGNIlGg
eQrRuuN183ZALckhqVIOXN1L+0L5k3kKmHTGRfkliNRtg5opW3P3IOZ9aTK+Wb3w53qufIa/8uEP
Y4+cqJXLQ55v7TLMWpHOgs2iGEl46dX9W0LV0Cl0UtN+Q5xY+yWAm49PK4ckDRprSAUyXpBJHQF1
9lZTRqCV+v15m0c5ALRheAS7uAidMtUxlmQz3atNQjlyXonEskJQ3JBH2tDEMlOmU4xm2l09Dh+U
+gX03Bqu3Bbz8eiShazA2U1ieYcgN8089VM3lCDowbB2ZjYIcXD1AklAVaKEDOinzR8RF0ZnCN5/
7k/JKKVcLkU8cNZVNaIQuBc81e5jqCeb3HFV7vayG7+0PYb9TQ27opWuKiMKwy9gBRXiHOOX9jl/
cNxWDZxpZqHMQTPPBWvSZZODB7tFYWOf5WvJK7uUmn9gY2y3bRz8GcbfxKZwAypFcSkuTrDHpMHB
goMgk2Jvrgj/ftYCRxeQJn1RVM1JgE1TWzbGJ4+PugoiBSTBLyiMyR/6GyEo5BeDnarulXdBBaSo
V96oBDHnVS00ZcW/2dcY9WdPJ3UL6xWLlP0eLuS/oJF1lVS58VYGOs0cLQyvDiMTukg2A/Q/fmN8
eIQa5b4tv9wId7G+UMhrmR1o8l/Njo7wTcf71Enu9TzBjYWYzuvv8bFbk1Oc0jdtOlRnK6kiiI32
vUjQTf0aJ7bzau0NBYVAJ2iXbzU91Ed9zBzvuEG/qTt3+O25UWMadHTZOkK+euA5BM0192aG+iCj
p3/EEhMd9q8T/ZymzpJgQxsmFA6JO0kafz13tOU7QkL8PMbZlvTKlr8TfkcbChasR7d1dEkPZhku
p3Dzn58PCECuxOad4lwFebIwENzRVfqgfuxwSRm4iEvq/QCq70Pm8iKHbQfdlI8N9pfxkK/X6Fq0
BTkCJXVMclRA3JsIVc5rLKQ1J5PaiU3PmevsyOR0If2xTotxGCknZYpfOFU5LxhHKdMWJj5uesBj
BFrTyOxFoGutG1ZI8roTOQBig4II3xNwL3PdWtE0Wfm6l+8lwENr+pQpsSSJF+RcBV/NgTKfdH2u
bilb5QXJP4KgQcFumpP71hsKbW9V4R+C978b/+kWFu8wIoPSUEhd+JteLE7fWdyx5rxQ67gECVmD
9dvUSybUDIR8VyjYxZUyrDRLxVhcYIiqro7vz263jYpXrtf46pQYcFrZ0NE0eTCK9hRnwrtWMfYy
PaCiwEB3VCIoewZX5NgLR/KrReTyECnbfHMSGNXco2ai73WgSIkgtUjJa07DAUIoEoGg3GnWqxec
NdiRZqS/oBm4nLXiOEqrXEZl+jEVFBCUAIbzUvO/A6mF3779rF/Hs6zmHMTNc9GUaMCRkysxVMdh
ISede2scIvyUgeR1TI4YkicuoRGbgstF/EMgDNo6H4CSqOyslkXUbzjBhUmT29ch2CMp6tdnmsTV
U62e2YtpSP4pxOk1ClkSrUJiR2kFLqYrtqhYc70cL56QgAL7kcjOzywe+l/NJt7aVbNJira/UFhl
l1PAch/BhopSjLlE4sy1LhN3lmLeqObO20eExU0Q+sH+HAOsWfB8swaKWtKgj3Hai186t4dhhare
ftaxY5YszjvjKom1ess6yc22d1YmYoNaRjWdJALZA1GTjMXC5cCFMNCB6wJXt6e46VRmUw4Rg/Fy
lWDHywkQ2F6Xmn31+SUe4xZosRnsGB44wun/g5v5woiQjXabLGBKX32Y2U2+RoATVA5nLLF4gnj+
pHNv7hQhlntrMn6XmNCFXPJ/WP+BhbMo6eIY6q7/f0JzcP98Box9PewHI3bvkrN1n/e4fRcVTvl9
L73q50Ar70r0M3qZnCKa6gxVDcacRUm41wpZ2/Pq5jlcFLZ/OQKwqFqBj0zAHRo7LReNYUkW5LhS
C/dA4rnENiyOWe25ZsdgYZ6QKL/vlDIfjtJiZwYIFphU8MdB4de2RC5TFSaoUVZBFd9KR51MSZ98
kFgCokb0Yii1j4Mv5wUNuCCUQaQURnrVoczwQ5KpAJSHE7RJAD+HGeOVA4yMMAHiuQTGwHH0mjtt
ZsijQTjM+lPbZu1fo+EpA0DXq+6gy5HxKPImujTNL88rkeCBFfAjIcKOL8YNoqY0H3zTqGtrlyh+
erZMBPxhlDMFMSaUqdmb19vtTWA1eGpB/iUa/K8lRQhkf790r+oZ6cNKbURzPi0J4ixo2ATqCho6
LvBifeb2V7LL4iy25jsfTOPvxphW4v+G0QZRjZ/xqREoe5xVeQZ5J6E6gV7SPP5YeBvBWsTEKZ2d
vKg6pmx1BwvlzyRVZuF7YGAJmTMPs/nVOAy3ezA1aVpQdwBpz8oq+5Hbi2/Q4IjJIDFfHzLZzQYS
KonJVokqY0SzVTc2CqTTNqPkbWLX6Aca45c31JDWyfjAlYSXcNfCkFhz8Q4IHMFJjKWoUtwJksxQ
8+krhlBqNxJ5gckHr5dHmt/A6ELSeFq0iDqnWJtHcs2unYxjLse/mVKkKtoAPm+Bp3+dXVBK6BI8
ArxQD7EsVXO7Nq97fdaCxY/DbPLI9F/kJhzryAId2+3636Ls3DVpSASQgzFeHLGhK1Z2s196Aawr
s0wjtmVbbHyrrxdsPmPYbscQq3gRQy3QHl3YtT9Knxi06/cWFa9yBbobei7E6+qL/5miX+8eplbq
ILADrVlpQ5EVVhyKc+NHESYcuixOGwscVMjXXYcg1erxymc69/w2Ak0yI94Pk5BA9BTXhF78VRaA
tq5UpY9H88Bhq2jUICUmaGDssnXHsXbA3KKDsKbxGIsL82Ew7v/m9HBYtaQQ2A/639pIO4rKaVcB
g/0XgayD/eN2n93INAhytkz1GdxnFYZhaKss7ImYK2NzxOpGyxsFXUpqfyMG5APPOKSbi73NKxue
kHNBcoN/gEEIlb2mxsJfg7z6/mzXa22tWqBvfKT11e41mjOM/BH7o9DjksWvjui4t2W6VbF++qQt
ffgHd+nIIVCJaz9FLCwrtt3HmoDrWKRGkI9Cn4Hp0GdPPT+b5Ys+ESW9NOVe163zHRdVswrhGtR7
F9lrrW2BOiMOUDo8mKY/fBV3mSR7wd75Yf1qY9OwfLyIweEAm0iqfB2QGrQrEe2O4Cav4kLz93gY
2EKLJHXp1p8s0AZlDOdzQ/dLSlXKsSE6hK5zeyoZhXcTshz+8MWtOGwrT7wWIjOGQgyQTxj7uF74
7OO+CWfybwh2SnfzEMKidTQ2CFtvJqOQhLMVx2nVAg2Bj7dvOKy0Sk/vLlk3TcGu/iIW/QK1j4jI
UC14dZQ8Aj/4/yQYYqQZKQpArLuHPP+zUWRvL8kXNJcXD3+gVkUSUpWF/oATZ8926D0d3b9pLlfB
0RbmveHxvnbh+xbR3173g6qNw7nsf90dO4F8SakE1IyTlJUqC3g3xZltgXN4Y2MvKy+rGsP4aE0Y
CgBUd/8EuCyEteR5AcMwko8WXvybu5CKkTCUNNUzfzUNMgVc+Y/nX6X5zcpHvGVNbUKxyra2S8MU
tw9CbYuizsr0bMn4Vd0c8ByIvLMcHFDh3EA4RYwzcQeRFeVxXko6irz+xI3okZcY4jg+nOrPH6y0
Qg9bpDL1j18GZc5Kjs3QOcdmCJzNLgW6AkEhVIF2f/iGa/UC3ePDGjSV4ryJv3Jy1pYRTlxa7R9r
9kChWotIguU7G9W7Q67VmHPJ928MJ1OMLxubDenRgLxSEJI0wi4yUY3sc15x3GTe9Qd6l5CZ4N64
ZMI8Ek06ej8M0ME+okDaeeci+Troyww4WH0njRmCapXMHYOVVvlqVu7WTm7lPigEhL9qizKoN+hH
LFhXQMMdOkMeCOb8oisnaJTFvyBSiXxoFd+yM0ym1jLmzfU90yU1DVCyenInckFR0yXJijLA7gmC
JAgkWucNP58rm4F7VkZJVz3smcY7QoZaTy9rH8+xC+ftHprIs7Qrvh6+3POnuPi31uK1WFV5wPMd
fnqTu2SrFlmUi4sITmKH/+9fL5c3r6TXhPhd0sw3FSfCbJ8qKPe8wNjG2uk3j2cIVmaXjftjpkZt
zoYHKYYYFQktCOr+s/ScNQQ0/4zrZCiH6P8JAKkcPIHCQu5NmpXRL2j/C5yNeVznf6DyCrISYJ94
ayr5mYIdSAixwFVNh4igElv4d7LTEHsdlDd0dibyzeLNnL6YMQpwgazKMGAE27Fz9tbx/29DRzyM
16I/AaoXp1Wxa6HXGYmlSLz44U2O9jTs1fJjkn2Zdrm+mK8waZr+3peErgRQLuuyuu2MdevRx9CI
WoRI2RuGXVNfjrM/muVG2LZuY3kOjrP0aWK67hTn26Fks/O8jxswgsRz3e7VPqEbzA7wuX0UqHcl
mrCr6NXNsccFKWY+qNJ97sh/230bkl/78eR14A2qlreFWDhQKdg0pMtDF+7IKxcdDR63bWj/b047
WLBbfqDw/MfOdAT2J7CmPdJlSLhcsc+UG/jQHwdCCvZt4iR3/8yhgzGHOnNNN1EDi1xvDJlY1N7q
vsqHVVzPJnDR1VT8VT52eQ2sY/7Y3Lyz8SsurbxOSgMQByyJXPevZLSNtAGeqV0yQ6H5Yl1dI9JB
wz4TOBfhtCve739NN0w5CyFahupsN3JDb1k4r3lwXr/iGSixMNlUkrdy4fr5NUMu3oTCcF2uWZEO
HpCIz+E+QZHuo0alRFW1KjW9E4zmR0Ivuh4P4iaBPQcW5rpXv3U44/rD4cEPdPjHHW4/eJzn47Lr
+UmTWA+XB/2wBCcPrGGI7WahL76iH0h/ur8ASkjuQwH+Nludchnl/0yRCsbBeN3QZe0j+Y8nfHcK
HAlPQHX+EJGJhG7H1ixMbtPzE46g5u4OGmjUkBrgRsNd0n8EGkBtFh0uOIpmUK0bIlv/zH5cFU5c
aCd1+5KT3w1he1JVDQDtcZjvlTUJ4StKap/nSVVPoKu4XFL4sRmIlPB1eU1XPJEOg5cJxZTUgJ1I
i4c6AbBi6X2edNq9AOgsWVwLxgt7C98XO9dx4edZKUiup0CksV9ngWeGnaE8d91+RMkTN19lvYJi
twEyOUy3yZEiVwUQbINjdx0NgCfPUZ2OAWPbRGwrFBVqRqzqMXKEEqTCrmQnPP8JXugaxpbFks4L
7fzqxYWdzV2L+nkJOArxCJNGR8ToPbRLd7/yCJVQd2ZkRmIuEPhf2/j+Yr4hEqdQ5XF8JQEDffMf
n7vKIFNL0B1LAOYxBstDz50q+cSnVlAWHeZKatDjcub5lRHiYTBXcQxSHkqImo02VbDlLGwn6Equ
FBs+03VwwVXVGfsgxAx5Pls4uQmBe4yx2v67Tel3tesufEdMobZsTcVAm/lsqPQWlXc/qizwVKff
HrpcMvRITg5vjHgaeu9Zdr/ASUIAbdwYExgFFs/xH/Ec8Lk0cONXxgK2azZSHmWepVUNGfqW1ZDJ
4O/y2zfWY//15KXrL0UznKxtPTag8bYEwiz3Dyyj1B1KKdgiSE1cAKJ0BjTgPBtGlVwze4TGVZSM
rJbewflm56lbpilGNQQnTF/ApNh5BUyoeFpee0QJoKAN0e52Zc5bi44ekYFA6YTcNUYsxFsJ1Cz5
ioOZvk1W8nhC6FRlkjb8I3fnHpTUprf5YQjWq99FqqVhwoQmnn8/4B/uw3XKh71Tz6hoFTywpjgm
ZuX6oBjPMaYZommDAq3JK+IPz2p52VGQRt5BZ/DL/iO1+BsusCYl0WLShM2d6cgDpe6pYBuG2vHR
Ai15tzJi/UssbNSDqO6Rmjw7OgZ38c2aehjL3NHHUoV532Ajg1M3f3vCi3KMSmami9nXNi/C6cSp
CbnSLGmG2hBMKH0XtgeG1Q5CpUlGfVxK1O6SzYRT/xGHKfu5BAjGwUMELlPba7iZQce/mDctFs7g
nduECfylpYhEBJV3C1CObeTHK9k2QpqburNOAU2kItb46jHSh3wuR6XXxIKwg0MT2OfOHd8d45tQ
7LWIFOHs19S37KrMVSZ8yYqksxE9QtbQdVFiWTsmFx3fjzzCfa2pcR42j+uS9VJaLyC5pUyK8iv4
MmsUGlUNj72LCXnCYiIIi8v4UwphbMlj4/gPMw4CAnCTEBxvViY40VJWxWuuva13lAkDLNZnxBvL
CQdn0Btj/qlqgRR5nsQmjHAJqlLEmOE4DKYgJnQN8toz11i+Mf0W7sDf7rxIeXKVQmgHO2Fg6F+h
3ejuJjrlrtFyA37h6JpgaxtSDCjxpN91WBf/SodLLjEJrjWD/jh2tV1Vq9ucTCSyCXIySKaDdunY
WLof3PukvNXOW8NxrBToEA97KkpOOw9D1krocdWe6WfW409fJnYIA8AjzwhB21NQqNEshRbh8IO+
hngAb9kt9gMyb75szRL0OhTp7Ove8odBkJmnuilzScWf6NZ+sZ2WOhKKgO6F6dLIhRTg9dUkyWbj
x1SZwumQzstH4cghEBzTXgzeEuavIkkHfFFn5JCm0wApJoWJ5oSlub+69qPS8ojt4NzQ+d7zaT0F
w0VsNmqw1HZOSdjPCizgi7uTp84TmQ5OHlpFGMowJhfqBYhpIeRnD4xD7buVjQyv3tYeTz9WV9R1
jbLWsDL7wlITpaociOF8KtvR32zC36sAPd4rg68eCq4FvCXTO3SRYnJHbCnl+NSJwFp4pSc95qjY
u9hucPGWoLRNT7BX0mytxVJitp4eF1Q+EIiRK9mzKnStmP6sIYHFB0hLEvEgctSsgJPj/x8LY75t
Racg+uRvoPvqfPG0FmMdGoYuGTqsLnsTompzZO58VvUxoWSNqrmrLsRnc4dj9SRYREnz1r0+tmaY
aBbQUcgOYDT6Bz16C3lYbY+TsHSN3B9YeZ2tsPd75hNRzUt0OfWL0YGQfCa3Ywy6gnYx6BuJITiV
jbohVxeYoq972l4O1F1gRJrzL2xVw77r/RpNSnLwO+eMjTG2lkyTjFym5bT8fBZSrVZ2YbsUBbdw
6IxmuwweT+NBuxllT7YpMU5CyNjr6wQABm6gLiLYU1GhNZqh2wILEBmbWDJymGWdRM9UTntsxeHY
eAlnmwuXL4Lro6xK4N3JcMOaWHZG1JIB9S2b1KV5gJBpLD+S8e2mtnZC7L31XXihbkPwl6molw8v
nIHHBjrhYqnkMPdOTAEPmQZezkjHu8m3CGEokHMHKnlQqfpR8QpJtXLTi1Y/hAj7hh3frrKJP7wi
nyorgXuIIucRemCmSItb5zir95SKacdekm0LJa1wSt+4FYRKTOugmwY5ZtoZ0hpNHqpJJy/3bXqi
s1sp9ooo87vltmgiNrARP64fT4fzGDg8jw+j/f7vSicqnJ/TGvcLSbzmrlszArDfpZr52gu+dlX2
iJ5Nh3SE1UBKOpYvQ5ccJ04EnnZgUoDDTNx7ncDqFoMIgRJfH8cFNt9e1UHKoPVaNtAL9MCz1Fqr
aGBH3RWvPDJPJWQvCQDyung48veGOWuMhlOimQboxDU0mn/KdlxqCkkjdPSaChc/xuGboW29p0CR
9Z6K6hrMnAI6/5BbIFpZIBbJTbDH8zlGfgfEmoV+AyrR9/x/y7nk5TzZU098GwjtWynz5vNr25Ia
eVfnULjK27JKPMD5V7LgGF51Je5rZnNFxyWh6VIZ5q7VzbNKOOKdOsNflay1Jt5ZwLb3RdvbLKtx
tlbCAkRUYTab5OEPLwnvNVvBi4h2dSqtIYV9fUgi0hn/NRIC0BpN48DDxivldxtcRm9DWLQtz7qX
mcIUuLTaGW/5XIQpWimGaZ8YnutO2F6wc4IaZSyBtSEWLpT0mDCWvk/ODYfZSzgHsORBYdTDcdX7
QLnAOcIXxhHdQGDpE1EBTvVaEZAvY4Q3h23MTELDtYrWxLwhruX3cSaUjVDKQ8SqdpXGl9fPiHWc
VX0TW1uTQ/VBbSE4lozC/W/3oXUjxKgI91t4l0hWcTxR5o0QfX2yuszdbzmqOuLW1fOih+ZJUh3q
nAyNrggb0I8xnMJDtGNuaow5MDThGG2TBxqoz1YZJNyBQ4SJfGZclCO+qNk3UEDs1hdpch127Uqm
B+5uCDyEaoR6EmMih8mqA2qq+EhPkRAG/QpvVILJbLUdgVkjF/jYDYI1C2Zpx0kBCj1iVRQ+vw33
Ittj+aNHcPkIKR4lGLQNNuKqIgT5VgF9AyWoNfEhBA/+bj6jV+GzGAQ0WG9HVXB1coRr07zfNnDs
p9n/UTpDwNC/NZYmU8VO8B/8yZX6YakUTcPjBJm68esgraYQ6+2oBGk01Qd38jhq6EGUOyltVrr6
dWVw4mshXhBN7UnL9D9V29vN1HlCaIVEk1S2M4vcwjcF3YrLOz1sHIyWzwJJWhV4+c85Io+eNmUh
UoVsmRJeiqIgFyqv9866HFnbjZIIAPnTO21mDuP2PPiLaxfE+SE9VmmFofM5GV/Tz94WhtWZ27FD
n6UBJU5ZO7UxrFASXQOfalwcFfE0SlMAsZs8y78Pfi6NBf3QE7QzNjxBcKVFRankLtj0/UvwUx5A
8/0sLKnhDMEncDCxN1PfOB/s+KmaZz6eiPBHNv4zJD6MFt4rBwF4HHiNll3i2AHVR7hdsj9VIyb7
B3kVm8WRpzsP2uGsFD/73CV2QpkuEgmWiLcIVdaftdCpKU//OH1jHzNd6GaOZoXBDnh37QZ61e2x
p9qdLdcLrZlHrUh44flazg7YVsp3cScnSc75oIYnC/ubaxM5mj1ygcOavgaOx2B+GnQkTA3Jp5wL
9tU+gMLYg6av8FUQCSAjl2unS55Jk3O+o6RirxArmK2PRkR5KNptxHCfsCDUSyn7YXahRNTDOcE7
tGYWULdBrUaNJeWxugoEOavKnTVnk+bg0w2kVMWP0inHr6eXb0yOEGi9Oi6pD+a9Zx1EJpTosE1U
oedhra1ZL0PPjhjSSnYneZCt7DSdvwK4lqIlTi5ujDJjyVibMXvLWLzYzVUE88o/xBf+wIU4orQd
aRigbfvxkUWnd0jRsi/t/QMLEMtsUPUyS730WYr9LBBG+Oo538uBckFoiIUWofF8Q72HOaTQQZHP
HBgoTGProJDpuc2WaOjTeZg85dE9qxonfBSCSCQYLadp2KiPk+xEX+xTOaS18QFC+R32eCmI7ekz
O0IaVoWWVoMy8EIbln8BGgp6aHn5Sru4qxpaSY1UoAMRRbnRei7DPdzrcVhYgemSDOZ7wwKweeJ5
q6d0dZmPIrBi7WajWJkFKVLDY369WoEkIf7Puo9AXwwxYwVzr9oti8pwJxjMiiiTAvmN7ZerxPJP
ll8uX4Bd0SA5CKf15ptFCTDds2NC80U+gBzvak3mwCu7vknvInONKAHBeQgIfeXkmKnqoA2lercz
8me5j5AhVldj1xQ9eWJdP/q8pb+dzfassEN1M41L/BnGYDKGCUZc9ijn5A9T5KiKHUxwW4lg7WdB
bVPf1RBra86469rweEsadWzMBYesHLR2R9lpEPi/BiIVV52WavaHPP/uJTbVVBLd8YIDNZ1tuU6W
fbRs5n6vwUzmVCKose/jYPCwXz9bnBlzOAp1cUXZmxE922p4d/IMP4n7d2knuEoGMo6ENvbgjWtq
4wMRU22RLm8GBPxLDbG3dFva/qt6Kzk7Qjj5Vs8LilAlK9KlIfrQLYN+ugeAgrY3hCqp9JU1liyL
7FenhpZfmWmTtS/9aOjXHFtuoSmg7/6lQiBXpcG+QBsN6ifNBU4GSXIcqawnShJ+qFX2Gf8I+Qrv
wO8r2rMy6gPPFmKlPQ9Ry5F4F0zUGqroVNJD00HtCEFrxJSMTEZ48tDffKZSXe408Lw82h4FivBI
YnV5jd54pTpZbzcePiIC/wr7kaKyznPK2aG+FKov09bsZn6M3J6afUlPMcnWcMj6jF2ZJ5xB/XOb
SbcSAOcM3P/LaO4br5h4M56HU4IZtlPT1Cyh34Pw5oqUZB7ZS4s91xAqckj8DgedcJ2U97GNcykB
uTWjqrzjowFqt8P98h5dbtFZ8G8STkmKulpjg1UuFDD0jFzN4EQxNA8B7YoMS1I7Lz2eagEuQznL
eSlHnqTP2x4vvBImsE03E0JyJ4JhoiCRRlUBVh6QPq9yLVpfE1PnhHc8/PZgAlGit3MU4Qrwbayg
5yJ0TGnQxxt4gUziBfFtgp5TlitRePohtKfwWNLYDhOa0rT7cTkTXCfgNG/KDVjYP6oIIjO0sPuG
1FlwOJL1t2aXvto7jWzBxgKoHCqyQVGhITjCmvis+2jzsIqXbZaLzZbdeSvymhgTXlsE3BYiuvZ/
aALgPuQMlQzDgLzoqe7D3L3ZsIx4IB61UELxllcXi/EM1Tye7v6eJc3JM+EL+mtQLL7I1DpB3GQM
GKpSwxYC6mzn+DmFLXRuzlrcfHpnfHC+0sq32DdO0J+lOGwcNkxo2s2cPonQEjYBWO2Wy0Z6qgnz
bQ6vRb+u/vQi7tOyeh3H9PnNZF5JIzxKSBGRmvcxJdYdOF0vsax/jPekfWErfmgsBsDhhT0X0hpI
1uKFPpN5GtD15/pcvfwmgyPPn7TSbZY9HrhHLMgrikoDQWj2HlKMQDSeJjmnQHjo6iNg+GLQUCaM
Pf0yXrH2OqxdzsHETRlz6qjl2o0f//E4nN8dSnBPG2Tm8Z33fnNVZG534ILuCJebdzzWxNWRvGqp
q02F6EMC2NqVGRADSTe1IbZWVPhlapLbVVZk1liozq1mr23Wwn+RsmeZ1+A6+dV6bvlW1DMn0aWZ
IWvv7m98NBb0Tgq1IJZA8i31YAkqhalnz6s20nggGEZcg567OyeV6y4H7qVNgjtFegYzjpnEOVP0
c4lVc8ywd+3p7J3vanlpPXjzR9vIz4NbZ+AUse3ANVF+oZXDYahxAv9t+Kx+vVATb3YTJavU9Lu+
RUL11yKHvIa6m8JzP31s4+NIgcYrG1caYzNhko4bdIRe6zluGBIm0CvXUEN4hWXrQZCGAvfGroRc
7t5KCKONE2lWcvaIirHvRWEWXU5RZfNcJYkpdHrxnRuHqETv+ky5/Wz68YQiyZc/LSIubk+9oVYv
9CrGjeQe2CK9hBnEzL7+GSiRB165VtybOOvew4itLQoM50lEimBlGZToCixbLz4BRb31CelaVgqN
FhFwHoqqD6surVVO3IRSFtiRmIM0DXL951tfblOsq9hMbj0/raYURFCZoQuP8Vd+2vbxMtylXJ2K
TJMYCQ0YvViXu58rxiswuTx0qKqFcX8/3NmMUgnM+r75K5DfTPwbNhvxKkY6xu2+W2z6k+NdmnWB
QHMyg/XKu7sE+4VVIyqAgGqFMrp2r8I2ccdPiGv/eHnszQj7R7kEg+PVPl+Et2eWHsBdDu9EhlpD
skb/9J6vDsGp6bplgSA6LKTo/T17/JnDqjDuD+VBGqBZdZ0t/3msI1wrWW5saLpJJ7Zq41lUsycf
4cv5AvUKxAzI3b2SEkOe+Oa7uDCV9vfYsMRuxkl+dOsBgClTYVKhJIdeTmmJ7WLS+lSYoSqTu8oh
VjiFnEERo+1bsvp8r3QN67ZW695OecP/NeJAvZRBAqvSh8mh7ax6Gb1L4YF0ba7+wXDfCUuVLavf
yozS2z8i6kO4NAQOzsuODej4IaVMvn8wjuj24Kmup0zHP89T3Ljw7EYMqPDellR+9UYQ36V+gqTr
Za6eba3SGGcbBLRq8wlnh1fbX85OYBlNod+Yqb6DQ+d2hC1WQ/Ufc5gIh5NGcY5xjS5oOZuWs5FZ
Od8ToEWw/EMu+0HukDmjfMXBo+FsAOIUiCwLj1NxGb2GDBkgKrnp1oDd/WOw6PIWE8C3iWERUKxr
fyQ7tlhPkS0KiSiVhKrdFN9fXlt7ke+5tP0hf0yiP8anRhfSW3PGDtdnx1EJCCYC9Vh/uzaWZZDi
zFFp2SqPB5wwlyVeN+x0gLOedWBIOvdlQ72Vlz06OjiSHsnABQH5a3EgunTPq2VXYnnRc71M1Lgc
jZnA7ttrMUrHy6glPFsJec+7FxFCnWpcMljRQbHryf4jzNS1NEUhiD9nGp6uC4e09RMNN96uoLg2
QdQ0nS3TehPZe98hhhxFMIy4uTsN68DXTWu65ohaaGsy17fSCVmTaFo0C3SmAFZ4PfgnCk/hjV0Q
QIiilxLjvYo5vxouA5taPaa8rQWFonUnn0PWahk4wKlqExFhnZtcfdoz08lqWMF3mJPcuHWlQ3dw
QL2uNSLznbESFK3DkjTbB4IEjepuxD+CYRLJeDgpGWZoE6kYS2NfawDIO0SGh7Z6stRMv6XMD317
aDK9FwHD5w5AcJ1jA4emvcfA9eMCxv4UBIf8TCjCZJuAbZ+Y4+jC5ha8cUmLHuAyK4gX6Qk6tdBC
3VyiTAKmO1ZFeVAbe1nJb4G3iFpA/46UV3Fgc5fymmmqrpJejx/paC3yaw9CRR23GOKn3f6Ished
ssSSRyhAZaLDNwqEzael+kli+AuY6xSJh0DWV67j/DHegrU0saAY0A8fWnVxZ0kW2XPQ8RnUdTBb
+XDvHglNmdqHU2oxVOF98EdP3VS7RtvQX/mMfp/nX4557/4bhMhIf8pQ8xjC3aTg3VvBhUFSVloK
lvaUDtV9J8J8pGiUcBTF0k84+6rfqK70awTZvPfEJUYZvc4W/5zqg31NeGKkj8pmi48WRkb/Yfno
0PuZb3cJQHcDB5iTq9LzR2bXDug1kJTdkyfwRpdEN4VoJLmlY7LiOPTBPik0KwSTQW0NWG+hIxkR
lq6t/lcMCTmlPuinzRAWciJHcyVYYZKAw18SwpAXS4/6F4NMVnwif5wnHQi0ypfB674BQcAEKXOR
vkDO/2NQL41OwkTNOZn0ja9WHu7DFQk8TqKixKHE7TsovjkYEY1jeh3aREwhqI2eNjzduHd5HLQR
4gEZgfjnLg9xhpTxtr6Xr/pvOhMLbJQBlvpCVdhM4u/tBL4PXUu06sAnlgwQOkt9hyYIh8cMNQBc
Edo6Q77rkxWDHu7Cim9PnIKZDFWyd6Dnxzgq8OjAQlkPwcxMuoMjZbo5SPLoc/EETGIp4D4cEPOp
d5uxRGRZiB0unbqs0LF13iKQ32CScinn+v8byFuq+nOIGMeSgGSLmj1gMkm7j3VOexIZoXVXQPOA
zT0De9HlOIVEYn67NgGH16m4OzWEzIbIo7FzKHX7Qhc1rAk8AxzX0/w7X7jADwxnz6nPR3A7utNw
b18ssXVHB41W8JtcmwVMkuHCuVkk0L9ULUeLMJnMJ5qzzNAMtNe6ffM2nMh5oeG9G+q78lNgXgPr
bWRTLGQLyfkuG0fBOVXIjuWeWcGlFogctlxaF2AC+km3LkOWQssjuiQU1l0ythoHwHHM8r0Ohj/1
liFLV2b/SaIrQ8bqEfPV8JHsDmQLfbgQhuBC3ry9nsIZjO8l4PssuArl60cDXMHXJA558hOBhw6s
i9nSIw1rMxs4V4WbdIO6VM66ehzZOUMFuLE8+L68B/a7excTiuXUDowGyCv7OMgsbFmR0V+UlTfg
QPRU3DD46wd/t1H7VKdyacqFWsyaXymQ4yZeha4U9plHMJBUm6bWv+0FDGH8WEWkM3+1/f6wXt6V
JzlhyN6oP2KO4q9dtSOaet6OzGK329pIO6ANUKZjTPtd9h3eVkSQ0VpkTnTfrhZEFYl/zdB1qtMb
9SGuPOfPpQz1LRwbFKhLQad1Ss/saRbtjaq98TJFow0CdIiT/9ricIGm6rpHD9H5d/ofVkyGg08b
wTQlbO/Byj9Gew/0brDP3AoQCv614wyp9TTrfBrMowdp4OLYrkuj5bMUQ/az2pUZrQmVrnpwx1D9
1O7MJODeQm4eL05IQIr40gtJtu+6L24fHjUFCcpmkwi1eh5GEypitP++QzuX9ugoLmbW1mLCCMnA
Lz3td9FtATw/Gervm6enCHVVY3fu14aQv+OdduCKW08cUALTy6CsKHuE61alslUkt0vstHmFtvzg
DcWVbwTlbqOvDTD1FbPGMo3BenaEV0UUwnz4xVP1XSogwLvmtmElHJcJvhxsfT/h/08fMZeVD9li
ms9wOzQ8QYI6DEpOoOjQt1565Zt/gR2tAb8nv2lUbe7J80UkLt3LMmNkGOOd7v9qMOgBTllLqKMb
Fg8TrZvvDYr4o34HpPlTLn6gURAsFwKdHHltIP+FTBDWla7CWee2ekpBpSvqTChUehHWeJlkgF3o
MKkqofxuM0fX/Nw3ZWya8YD0OjYVCyI9pv+NoIxUXefxyddtpuR0gXtQzkavTh6XJ7SEi/jWZsPV
G+pEF1gUTZ+FP65umY2frHMVX6A2ISw4m6zupFhNPRFOBhwOc/BRxQQ5RPALk9zxPY0kNBq1f2Nc
CA/pN7Lc+Vy+Yn2aK4D4EMKHity8XCZT3qaHbtUklpmNHIXb6uRb2N0ej2hivcsORN64lUTm06GA
OzLKCNRzY1WLhEx7HfJVaSooGUMVij9bq+yBr0hRfOmV1b1WEOMAvnJ7dS9oYaqZghbI+RYYmj+s
NVxcuxjDguvgFTqlNlwzx7eQuSlKpuUAH6qtHkABI3MOamIcgiJtPLGaWKWFGNhaH6PQRH4cEaux
8bjkkJO4NDviC3UWtd7rfhIEdMMBeK5v4AnsCRZziv3I2sYD7X3Votco37SL2Z8MyjNGxIPbyUgM
78oUhrRmjc0TDpdmdYZhafRRik/OoksATHKjRkUOJwaZ50URKkzDyL1vyqiWsDlM8nOW0tnXA7DE
a/Bp98yc8fQKAIFBzm3A6JDp9LUirnm53opRwLMTDE1G9N7kRLCRW802z3HnupNSyKDwCXJnVffG
fxyiffwfSBFi1syokX+aaA+/bPyo3uk6FYO78cTTRgED3Rjf3YOW2nGTsEJ68lPi6guItFwAAl60
oXXrhK5V4NU88dymn5ajO4EDtOlaIvHxZormdQmM+Eu5WAi9jVBJm+IQghsgPqgI/QFWNogqJsEc
dbcAlmpZLqMb/oAo8exzJddAaVHe2VhmhWy6mSSr6exBvDeny+hG2En2YfP4WPfoWupy+ZaWrSjk
/PeBjvneDYd86JLQvwbfW1WVyXo2AjrIJHnlyLCwwMqi/ZelxkjFjs19cr8GrRqdxTbNDGluiFjE
N4gsGyQf/COW2448hep3Ggf+PNnJL1ywThSaCbG5CEW1r1hJaUOtDDn0tirQUeEsKQQBxCCshJTU
oa9xXaAvVYDXHw7SjftgLQ/CNLwXZoMFfRjbs0v8Lssa2GWZvTIlNsfTR2JbcahgC71A/vVrV8yj
QjxXY9ds+/mzJQA7vn8McnKGYQmuNj/sIClvGfIhusnAEf02f0IeGMwjvGYKtiwzOLrlQdKIbRYc
mWdI8ae7YEX4Un8tzueQJnkBRt4UNo+Uzx+Z4JutA+DPxFKdOun9yJrcDU9vZ8oVd7A3zrXWFwWT
TLSEZ/2UIqRsNAg7eljqv0FSP0wqbwjqWvL9oV0E39+WrJveAZ9z/g/01NHYVgxYaXOz7o/vZHNb
W//EHGBtTOJF1bM4pw6qEOCrs91jZhr5WpSfX0iLhyOoacRUI39UmIDoahN6hV0JM0Akx3r8iI1T
xwlc8iZynyGBztSzLELXygmrS6jFyP2q6WSN0Ryemw6EpExW4pwENKfAdVR+oO6jydDrjALNbZNg
mdShG8XMu6dwIi1Bk2Ye9bBveCK+OGU8NlEa9iCWivTrHZ3JfqnznwJ/GLs9BIll8eqTdg8u+HlN
J/cDv0MjZcTNPSoTBtj8RNVMsq6OQM3eliXuXR00UjYTwYpUsIDEiR9N47LuzMGdECFFb9DtTHFg
FH1S9CsYh+6nTjBI6Bnz8Hq8GFl9MASLxX880LXVo3dr5q52m8wokWEULYZKJV2Z+MDRNl9h1n2+
Yh3X2JNdg1gvjDak2SiTB8PBiYdvBVaoujVTZ645aOtyEpH45PF6XrHbYDkBbmLh809S+SuHNhes
Tsq7VXt8h5TDcmJ1sw5clK1riG3aOBXqTyPmaA6wTqcmU0By2nkkaDI+m6dRK059XmTMqtX5/wH0
7h/95Vet3Vd5VrHfMBrYTd0Z5xYADEvtNCW9XeJCO+YN6YYnLL2EgC9PVo7odxM1S8Ba92gngYTY
pao4I5Cp6wdbkLanh266Phkrx79fwY7JIMkHN9mHK9ahrJagzxlN7KpWMzyGo3q+5po9H7TwmJEX
sVJYTCR3rGbP+HicqV81JiKCCJ9yY1BEICqGB5xD8zMTLVASfhYo1jkz8HAhdPnrpqQGIDPcEcoV
piPxD+bFkiKRWjIFVTvcoYmw12XXjoL/U5AR+uiMeIob963ZuDeP01746iPpVZv7O0ipovSmLLrG
vWYALtpbZb6BeXnjm7YustmMzur8pF3wX2rdCQFPVZYWwvQ4nXGTNGr6NvNPpvxkcINEqx3SLsll
SgzMNIG7PUMyVHdHg25sYHgz8a4Q0kY9uG7PAxqoTtaRcnHknrs8BRmLQpKIcelUm18K/mm3cRt9
n5pbq0+Yb5JLEowe79pHDAzvSknJK62cfzlqFivo3KUQ/lXpKcequRaS3koI8tCkYWcrNRx5FD02
pgXUoU/ikHnt+XnXbU9VB/dD3Z+EjwBWsJGL5qJ7T+D1zigs9oUBzz8prvuPb1Ar8C68GetbksoV
KpTrkAy9JckQueQVPMya7b3yzwehFM2E9mbBYMAj5rXk9mHx9huCTpOok/UU5V1A1ACt7eY4X/HB
uyWcIMMmdmGbbZI9m/27gH+JlN6TUvBR8RmSzEQ2FnrtoSXPQspuXFd508jgrrAtfFbqRJgYhywg
xJ9B+fO9pu/6RIh1Vd7ZEOQfonKasBMDPEGHIMQ6lyDJKyLQGj8VEBZIy0nvnY6BOn4aaXA2u5iQ
d8I6kTLPlNvgKBiUTkfOdzm5tCrOcgJfnfxereZbsdFoRM8APKR76w30e74hZe+nlY8fjHLsveHG
oulm78/SMmLZ6rcD6q8jkVi6d7zy5n10ms5vJy+Z4dXF8xqRD7cv+c3tIfLlIi+KjddqrGAzAPn3
NM5SIqeJpSmMx7Y8hrmCrp9kPweuOqPDQjSs3uDsaNlshZVU3uT1ePZQkQ1B8+jJ2J2Hokav0yOd
9PJXwTQyfHW7GeQyN4hib8lSHwwQu+WJd7wkXU9cv4ioDuu6uOnq5Vd6i/FsdP8JNmx9qucNMvpl
m0FPsHDoUaFx83lHOzk2Kwajm0yXc9DOnVqqRgBLMERtDrzD46YX6llSqCY4Q0VkZvvAgXq1BKHq
OfaJctPyiNBnXq/OZQHDxWIjr7S46qppI14Q47QnHJf+5/UrsygzR7fu0c5hjAHAjb+4TqZj8hz5
6X+uMdi+/kB+LrgeBI6fOoE+tMz8WQZ7FxZV2tfYszmNTSdKkg39Ie416IQKp3hcDGJseXr2v7kS
GnRSNNMAvFh4Y1dPefaY30iRzgncy17/Ch6ZiAB5WUnzenNeovpRe/freEpQV6eu0h+ue3G6LyTa
N4fBnxJH3IqvR46en446CCGVXQcAFdDqCpXnpghflUiocdQDbEd62FIaAd4rQ890p0fQpd5SQQw4
/ls0eQuuFldL/j/PMdt43T348THqHacg72Wd7npGo37cP+Xe1BRCKsJEyihZd/fVxcODWBTKeKfK
bHMpnH/3iFJ71hspBFB2JHER3pqnR8sDqlJAzPzFpXUimkzzGcyJEh5lAAag7z1tBC6IbTc217Zi
UFKLDv9i4PKjb472xaqYok+LgjVzTMgQ4XXiMgHmIIr0soj8xiblQ15wo1ZVGZOT8NKGJehvQ8tV
VMPCyvcnqJ3GxLi/vW1jtld/Vg1i2xYiTWhqNJ15HaN4GeOHcBKgkleZXsAjB4fPwDCGNvCEdKl/
ch22JKDBBv8Z07dXthU1+ExzeFCwup4wLcUvzgKZMXzxjGvzJ3aVgRZolcbjIvdU0jnkIm7xIdIt
MnC6NeW8oqR4ufulP7mLiFmMZKdImKMlDbOWuKHWmzi1xxhzVjmrYVurLOhWAweC1HYwz9APWZFN
WQ6xNcKEiBKsqnG4Y/1b+OhdQgjw9QrP3XcXFv9OOCphS4MwHOhiGon0h/RhqBMeKifKWVb4VeWu
rNduk62KTGVzplTihzshnKNxY9QES9yHnyHQSzP2TMdH7mLkLKl9INoIFnLEjXduyysb0SzHCvmr
vnMCqFJtqoa3ceFT4bQTcSJCvIXKppL6uH9N3J2qWgAqUBcOZS/8FqfwpIhcC3pF1HNzd9YvMowd
xDwzPZo1oKnDFOdWc18aq1yIMv+eByruTDsmyo2klRDxJ62x1nwnWWmeb16w7gsJKvC+kJR+aJIj
AroUp50WJorE2/AXiB+5z2TR3aEkrVw0KdvXnUrHeae6EmNNshvuddpVg6VS8oh6dWhJooRYfigi
xAsOo0jVAvxFWx9IuzjECFSylgy69MCjLLYA0jp7bNBdoTNjKpAIp7eu+lM8j6B6F329pNHCJDl9
YnyJFKvx/z6SMhm4MS1Al3cCIdDX3ECVM2L+XwM2c/7zzAP/7MRG9ADyePjD9ZW1Kw3d/922qh8x
kcxV55g2XHSUpQTDPr/iZjjY7t9d8a1ZUKE5RFz7tVErr06/F3rUqjbwGwPrxjQmSn8gYRzpO4hK
ixbFLM80Y4qezUO8EDpqBdMSwH7JID/MrDRljl+yFjzDw5uT8ntrekAWZpnOdSBx9MYBKJ3FUre9
G4epf5Gtemk1c+TbI5js5eTttmrnbBZVREIAnX/LEbTiM+x8j0WCSUIQDHsrmbIhql2hS/o2U9FV
+DPBrSo/8h/tUGKvSe/1s+mrJKN9OINH0A70L5o1O7VQSmZ4+lgkdYMqglR0U7a/I49VMPS08bMR
zRv1NJlSeKSyQh6AGbolVu718wolKIPkBoH9XSLOKX08sdP/kY2WHM+Bo+wv1lhk5aiyHRDE1dpj
WMWAzCOPD4k6VZCnYV7t9wWjHyVlRmuu26JGmRiONvf+jseagnKsNDAvtdtuVLVKgSKkLObeUNqP
KWMpvQzGc5l0aaJ1gnbyWSj6cbjRCH6v6LfuAfbk36tvhn1iZ9oPaFyCJUP3CBN+qzb1/CwWMVJw
ntJvOd8PjcUETdRFujrAT3pAdWLX7cPDzrRkEUw5/oolFAybzzeE+p9OevjXiRV467JgkO9lGRVg
eHBU4jHncGuBcdCyIHqgAtF9qK9/jZyoRzhc58leT2qNnGNqrb56SxtCoUe0Pvn86v4xhwl8qe/G
/RAYF+pIcF89h/AHFnmUfW3Vbl5hDrU9R3AzNthTZwkgBncX0ROmAJS3rNwVa+oJquJft90qQ4E5
5kh5jN44Uen+zcjQw2I2qkAxLb+l0N0a7xNiRY/aqcwEniVUbz8jtL1AGJcg2A80QVgLqQ1doYLZ
meEV2/ZKqF4viNVO1aaShLZttZCWX1i1JOmfl/GYdCqDCARcuZdt8or0XkxMlMKSH87ggZLnYaiS
PvPIUNVgl97JibtHvTQzLkSzrvFRWsKk6slWq+P14Z7K4rfcjSqsZrwoDryTdZ+LNGGlnfuQDWHs
UtJGR5Zvm+voTT2eURl9FsQq3zCsqRPSXr+SYBSAvnhraIEqzmyAvvQeuHPI6dIYTZCA8FCuxmGX
HrNXPdIdTY2X1NhexL7miL3QdZUpIEvPgP1xeX6l8/P4cCn5OrOpLSk+w0KO8g8oY/lGJfQ0GBYt
1cCY4nWkdoqSDvJytSPy6Kg6J5BGchZHJQ4Pq5LjTiF8/CEr+nYOjm2Lle5t0ZqOI0TXUTGkO9Mf
uNO7s9Khc8e2ShqJSCKPUSDz/ybDTUGByY2DqiQC5y+mwF3kWMPjTKm8pD82qQ0Fq9G6HGxVN8QK
BGpapwHG0M49L4uNVcvaUniJEX8C7eoE5XMt/kzI74xk10RZslXBnc3u6WJ4xp3LbCRsmj6It3G3
s3oR8DQyjymbcbBrDsoEBvdiBKzHGDyjMnmtsfLnJI34NrHzknzcXSWCvyn//JVWTBBlTqcW5opi
RwchWyZEhw2B03K1ARYFqtD6uDEYaGbtQciQNVpHIJnOoZgyrDy2WDYjaMuKCRsmX/G0svioJpk4
/SIaANI5xR9NwMVUakqlEy6jM/Jw87rnIhgMg/mrAu7kfdWhSjHs4upUaUf2Yle8cLU3ilRRprcN
PaXRmzpf6LdyU07fRU0eDnRyRerqC5QPuRx9XzECD0Jw2ydwUym5IinnY3pEY26eh8+HFZ2ejjxG
pJSobG3ovTBZhJvFjDHRy7aM5ltFxfCe/hOnX1yfihTTxIXH/eMwYy7Kxx1jWygGTdaOTkXYAeTC
DmmS5IALtT8zmR4rQ7kl07g9sOq3f8pt4ErhB1CxvQ5Ap7V2F5kGn9iTyarR6Kgc9pghDnOf9vQq
SpQfig7sOszMJmGHPeWTyWEPm6CpPRiUdWcCwzrI1FpV3sXdknx8XT68v2t7RQ6r8xNv95fXGzgw
M7PS76urQ8rU18rxZJbkylOLPjRcjPBWXFzTFmasgLoc9/8QeuuDB+yZ3pgiN1eZwxlK9D8LZCLQ
FBqR+WotYKu+WBDPN78v3nFYkLiBoud+3cTpIFemk0qEkaXdbLXMVxSx9OiuYmmIXvsphwHiWTKE
srdIin6oRZXBw9YdvvOjZFEJuIBeRdmwgt3i5cd8YjKPR2qedyJabaBVzkf1dGhF5SjHoqgscQGZ
ISMzAd7l0UTQUlJBGYO/RV0X0JdE8J0rB3vzzi+IJiPFAKfE9HqMxjBNyXEJNeKgqM5UE1+EM7uO
oMf5/ah7ieQUJcV2tsqNdFsRGM4ouOoIQfXCH5SmiqiuRskXyKzrx90pMGBR+/x3meXFrykh7LeD
gtwxoJtotxGhKu60LaWZInD791GskzJXgvkAMo7fezmy32Ncs+AqFr3tqOQ6YfNWIAFH3kmmRsOV
fmRpC89wWx44mab8sVqtcZHebznqOb4Y2AdglhLX3we9gpNZAVOmUW9Mg5+X9CmlWprCPtCrNNes
A7cF+bbx1TqB/sjYRsZG3tEoA6nkx1xZ0+UT/EJSgXzBsjwIacNfsAfg9zY5onZo38ZMmGUTQa7Y
UdZBxCe3kSDKriONVjW5YpH41OBMh6KbjCcDpAbcq6Yf3ZtgQ97UVySYKQS81Z/gJHB80zDXBJqQ
+d+l9R9DuVxoyjA6ZxJKWhn5MnT5ke0akW4hQJV+AYoSKa70Be7NJNjFGSm92LQ2i5RFifKQKk1D
ECh1coxAxVhbas711d2KQ/IoGceTjjWCU5C64cPuEKU0EhzIJaCoW2yc9KAoECGeEBUSCzLv/Nux
2X8nPsY6KQr7Li6qNAGAkyWw6FALCD+gE/NkXWn9PC8kPq0bdpvNP5/5od2DDWQtdYklLrCRibmk
R2bYddXxKmcviGuGqIwL+9eLZRPVic15/+oCKNHHu6pzif6rsxzy39ZOnRKtAFo8q44PSuhyxUXP
14lAV90lcZfkmCtoheiWC7XeP6yQ9RW4tu9vNoBYC8MEU4AAd7AY+jgeV8IbJAzs30vpmEZtmO31
3GmuGGOk0F26fk0ZwdquJDvQuXj9jhgAXt0/ZIBT8PSdpr8m5sdVXvAyx9NOpxAkMEDdi3G+aCfX
ObA5/c4AMeKB23y6Koo3lRieNo1xRn8jOjVzdHPGLKp/DB3OGpVkjybcG1s4s5gOEpESB9bE1QWx
9j/tBaOxjlJF4DLlyRQ2nwnARrJpIqGO06DYhuvLnfabFFUj9FFABDjNSQNwrf7V+JRDfckz81cP
aOST167aTn1Apn27vbM5C0mOHS7Guc3aKd7D0bFRa89144sV7s5l8qMyTHPXgQ0fIyd49h80WOhR
9hzjAnTCHlsVvcKvpjzoDX75WKzAXhYgG40kF7IUlrqNA8e5eCdlbT14MuYod9wA0v+2M75FqwZU
zbL3lG9Zn6V2Uq/BfXazijJpjJE269Mqfw/KqLF1fmPR1kfNgcXN6jlOHByKz1d7DmZr9018doQN
c2JUhRQGPpq0vn23yahh3ooslz6CmB800YjtKFjBjnQ4i1j2veD6HBPGDNfwOto5FQTH+3LrpcR1
dULlRi6f+HEs+G5Xy5cuP59hKThgHlJKdyP6YB3jYxoJ5ScQem2yIdjy2nqIvr+H9yT7J8rBtOg4
a9Xcuuhah80yAoOQASABWPrbTlXvaACnZla7Ytz9R0NgVUAJU22EVkGKKm5BxaqICoS7hC4KFQFk
cb+qtB114xUGnnFENIW8NkGNNbveHg60u7Vu7f72IKzI6Cm/APrw77fAQjca+hmau7tFjn9FNRjB
7QDq095VkaDgtancQAiMLpK2fTSSB1SpoaWTZQhbtxBH5o/A91c8W+jDFxpm7DSUtMLImT9S3Gl9
ZQ/AADPo91W9ZlGDa4UZGpOOtuShvAyI8oP9wHaglg6PI+N06EHu7X58QRmyepjXmVz7Q9+hefBc
xj/RuldH4N/xQ9/4SWLbuJGBVbxr3do6L6pF3myDGpOGx1qQWk8xl3dcC7KoRGMzHuYW9Qln7jVH
oaMZ7Or499UaUJziYdJFpkGfb8d4nry/Ooup/Fj4CY7VBtd1gZzttnTKolQdAKXMFtpDYZkC3uZU
eBCXsLv5FmuAAqZTGnV3Y+Si9TwPSDpnv9iuzx2DtqB6wnmvK617zXeBinvX7v/yHnPaC3u4GI0i
+xu+ynFcVrH6s1kdkH6qXDPBM3vwpASLBtXf7LW9+DmKlJAp74R3ybeLqpA3qmsE4bJ5cq1qcQuu
jrbkf6JD0YRnRCAtAljlWhs2x7JpI5NFHoQjf0UsZY343suE5qqYN/EkboPbDhK1iHFy9lr30dac
mPeHMKP42eX1tod3K9BbcoDtGTw1V3zBjhXxjRrlsrxzsbVdsG5pqWqDpZfDwdbJ6m5mXvujHAqh
3iIG9Z7IjuYhEs2VqZLm2oKmVqko+oKvNCeH6GHc82zbLgNqpa8obRIqlAugFuddlSQpW3n1zRQO
UPxnkgOhedLo50nMWSYz0CkwMg6K5PP5j1+wnMXYTFP8JYxwLQ1joBAXTOBpKaOoG7b1kR3o5WyG
kbVgHJQ3tCxxUUGGv2VctavoY1pA7PHqmDL7fJbp+Tw4DJE6oGwVyEokTRTl6VVYc0Cml9xoIpCl
95CZWFw8g9UK47G8YawWq2iKYZWsacC4LN2F+iDHvUnUtG/SG44y8gdWuodIPl9Y+7vpEQqAHwsF
7WdpajbTk7/BFlz2ecgR6Ykqym1NrCQKVX4zBTZDHEdQeLJMSvHiAqlWUPG4RUcA/bSm84oOQDB0
hTMFhlKa3pEzWVB+uQOeCKYL0etej+YuJd0OWobOhjuB38ByhwGm7Z4VwER4vR4ylbyiTZ9nbwVp
9Ew6GBZ8eryqHPgc2duu2VDv8VeGfh4rG/y0Jw9No4rEOxOMcFi0cpXBn0PP+P/ukhzir8y+P0tM
9V8/DiJlioS96ndcqT1H64YLEK0LKMpE1pjztZFnFeMEBBFZhc3sgHd9qMZ2GYLCJR6+lrZzg19E
CYPHxfl178e7CRizKOA9GSoBreobSNBc0YIeopfcciI3BaIgnIEtWotDezAXaq2a4ielcaPBn4hz
qXX13DoinORS/2Q4g/Bx+LEBxWCUuPH76AHLLM3fwLlFs9BJOZnr8OiaGilfmGtGend3re/10UJN
pi9owCQAL8HEUOV/cJ4yBP3iIzBNVCzsoNRMFO3n6MUDAJsmNHpUlz/C5M6/MqqI3bfQ5cMAgI6l
54WMGU3eFi5O9UXBLhgQep4p+TOQm61oA3e7aKsUBQjUO8ZOEhMLccX7xuk2aG7RMlTNHa83Orf4
cW9cjDkGygvzniPm9p8pkfc5Uo1jBTHyw3xkl3JGZedaMJ0O65NcaIGFbZzT+NIHWZR3UG1O3QUI
LHKUFq/CbEKvVZdFZDDlJC0nDqcZHKe6V5N3NOecZ2FIRCnUMS3HyjQS1LA0omriweb1L9WnJKD1
LIkwwb4YMfA86+CJVe37ncMqkc1x4oE7riEP31iRWE4FcbNtrRXL2l/xFTDDZYY528IosbkvDFqG
haqxflePe5SEVQl1DzMkxeDDFDp71Iu+A+k1BUgCgznwOJgMMjbsd9nUVn0WGGzj9t8E/NwjERAa
JkaWuqmlIksULU8ePrqbTxHWddIiToJl082UszVsQeIw1pli4LokfC7Q1JSIF9Tjrls0IIvMEkUw
sTyC6y+B4dHeWfBgn7nxrbACakjAFHFWPALHRC3kjvPE/I0S4GWgoypAH92PFv16ljrOrBDtiN7v
3eBBNsdEXC+LG3/5JfphUztiyVNQXd6trViNUbwDRwt2B+Ke7VDHZbpGrAohYeXl52juudSmYsor
NulBUzQzyfDG8nldf0KOQZx4GMXUETN4NsrmB1EKoKbh34i2WbJfMLLLKYCXUDYNKueIUzhDv/mg
9HtdJAoXvDU3NdqZ+FalAp2KIHuG55biVPxUbx+mAYoclZSu4p99+HLmbvDiA5pW8Yj1zdFn3/FB
Vt+Mhq1zHzxbwa9VEdQhrVjaDhE/FW5OxQWvmIhf6zhBycqCZPEHjTSC6c9uIHlorT1QImmmsLDX
ebcv90MT0NX//n3j2Uy8cWQbcokDZ6vp6YrGQFa1iE3V4Vy7Xrqkm8SkBJ7vsunl82sLVj8sj1Jt
VOE8ZW0m6s3Sc+0iYkxJ0mhBzTwN6oPlQuL5Q9mQvY/te3JjxNTyZoL3kA11YjXLksbL3RORYS0r
0yupk1kKoI9mc2YfLJZXOUprYl3Q6STi7IsU89IUozeoyHCWg4D1YCBWhql9JkiV/px03S2nj4Ws
VVN0f1DFgPKrDo6lSip2s9Q6JFH8mSsRpi/SSU1BSOqAZmEIOobCXOdfT+DjKWyJBxb+gKuPpe3d
ixgswYF7ICNY+EL+qUC2f3ttCDPtqXTxI8an0bUAeGa4epBI/10sUTlm/wEQVe7QRKn0QK19VtKq
xQUrDHYowwYFbKiYd746t6MJbBmPeWTmrv4399PqGxp6PnbE0NhOwGHPpa0eGD85XU9LHfTUWRBI
58hOUARGTtls3r5+6qVlZXLNST7u0nXdSUZbv0jd7s+m/INxlI+eXqVlb20F2talhr3tzOllbowE
DEWpjc21GpkgCodk69aWbhceg+YefP6B4CwYrY5lcA7YigdnNvr984r06MgXhAORPP3qDRyvszS0
NnvrBRaYFAUHteEissvi6njTbS8a7bpCFVQng04r5kL5B3kOC9BzpIzI/AsYtzo2mrz3h9tMB2vx
CwCX8XGEtcdXg6Zi9bGFAdpJ23J3FsDtZ0ylRPlnLCTqjjD0nOfKEZTXdbbcayVqXNvhlqy0QjUn
oYjwDX/fzOJbBja+m24I6zxUUGMHS39S0A17R+AQUtUAr7ucmSHO9VFEqWDKMxlGRyJLs0ocJG5q
kJ1qKLC+tFWPep1rHiyf2bbYvEqzh0bO9pgncM2iBFzi1RXteVgVtKMFRxyBSL4Q9EoRzEXi9Uwz
rbuy4uKRYrr4bIHRTQ8iNfADjjFkyThggt2Np4HUxDUVrQIeOsX8aK54fErk4JHBkBYvPSNR6BCn
pUT8l/ajK82v0qNSZmB4SJIf+BrzTp1CdIYPCihBKtsE36qBhcHVMWqnu0HH0KE+6oucWtQxevmH
y55iHWPrdFiX6ut47QuUTqjmZ58i9QVTJznqZu7hJIn5fwdCpa6cJxZHyHdkOisPkkux7sf2fQgU
B7fQlOQQlY8+YLNytHAXXEhWV1ThTDtD+iodERsHFM89oU+YkS0udOU+yPFr0MurA7FbYSyxAHhK
ZlivDwckQc3srPHLN3bcnBRjsl4JK/aqix0xMzyaSsii1YXqJFlKlWIOSCrKzoXIvtg4tM6ApBmx
flVf1qeb8RpwmLehbZGnwOT8wNBLGi/2r7/901Cm/d3AOz8mXs509j3B7gs4dzsIIR9rQWxcAg1l
a3MSwteop7k/cemi2idvthRui+C0ok9xq7+5nLt5CXHYUlF3EhOJ6FiN11Iei7+4jvNBD2BWrCIq
crZ/2Jg2m+BcNHmjk0bStRiKthR1PIUnfHE/0YcpKbxU12lzzWuRy7VvAAnIVhEPy905NFezyGdU
y6wBLp1t6bNvAnY374LsthUG5aD38Zq1Aj5/q0bXzicXvshSAVIPwEUSysZk728f8ZPjPIbr4KnM
LX77Q4u098u6NeJDZ7amohSdLAbtVNhCpidNz0TdjbJFHvqnORWgP+NcL658aZsQRR0rAERciQ13
SbNF7taI9aCNEteFU/K7Vlx3V1QMs3xVHz8yzptIQcMTVvXYO9QPQJhjCeGM+ejBEOQrJRVY9JBg
gCF869onnjry61dCSF3SCCAvVd/kaTvNrbb5j8c97Pu/LVgWKlOrG6tWZWiVcHgtdm1DcW0q11b+
VTbtaf8R97fH5KwgkaWaExq3GdrHbUcTYg5Jj2WwrW/UwHCqW/Qzsm0v6X7uloRleBLb7r4Fu7b1
UNys9rshEoC2NfiiC+mwL26rf4vBAm4WNUbnv3jPYN/Qw16Emd2XF/EQ7iBWmvkk3G1DDCeoIafo
/GJNbU3T49sUHwqKbtmZF1Mfd1XwtUP4DdJDfSH+eYCbI1HBSPGz8U6bb5eI+YluNNq8iejWLZ1E
l8qFXL424KjQfCW0V8WHtrv6ZkDlBgg5vw8tCucdTS7GURDlgPRnVkftKEMdPhipXN9vZWiCSclS
1WwdxAORakVATCE5Ac+fN+KZCOnXMmLWVlGxi5y1GtXqbnehB0a6ix8NUO4y3o9MV0PD61Vjr7g/
TQYSy9ii6JDkNp4aGaRENJ5ZuRjGQBeR2LIwPvjXqeBJ2jsuKglamV5Uk6biYulKRr9el07KOiaq
yLsG3YrHOQttckKUGsJQxfQZ0mRxejckmCO36OCX0Ky1LBW/nT+ch4k71iAeHJ/0ayiz4pZ5Ikhj
GsGTXzZ5o3JOooLEL2MNME9nz/YdzG3gOgzIM20DqQVZ5wD2mBx50EmqpGXhIHiNFiPOe5TA87+T
PDiPm2AP2cCyJOHtMAeeCYpnEfgvOZudP+P8mHPVpsC/iNJcznIy9HoOHnf5ExlpLCNtS4yDtBwS
gbEFx1IjFCmD5JI2VT3vZjH+YQrR8VyL1j7sDrpbauNu5Nku9IBQNkrqNz3Mg9hgy8fvQBsnLhDQ
9V8TRhBl2/szuMuphsHPqAitFRYQxN/bgSnZIEjfbMx1gpRfPwRqPLJIoYA//gHY5uHD8OQ7SsVs
BP+d5ByqzbYb2OSsR58enn5Cbw0IalzT5DGefBPpv2DoMU0zGTo8sxobSL1LS3EGot4EEo7igBes
WSFVMk3sfZcERGCj4mrhebWGi9n5WWgTdFoyZov5xEfqIf9umFIhxQHDjQXae/iUQW0wc1FXRJep
i+TQpP7IR4dZ1FuJtM/pIr/d8pXvzO3xJfdvA/lss3LABf+H3QJa6CzFKGN6b4dCmkVK63gpY0pS
QDyjLpqV8aItYH7GKTnOvqXEjlR2j4lUPm4fQVdHfbEXOYZMCQtW2x6gN549oriz9oyPPYGiZwv0
Zzi9N4rBvWkh25KpO8hwB2YQCOmtT5B0RehqxVtEK5Be9bxgca6icQvysxgvwwVyc6DmKiUZ4NDb
jb8OG2RYWMARyukX8Aa4NJrPu+NaPNf3KaY3tWMLQy8naWqnsHy9O4/7gT8wEIh/+9pYczOl3+9c
L4DZxmAknbfZ6BtW2rg19kecmbCtpJ4JB+XuutXXuvrGBxANYGZXKweeqrCAiPPEC0mGSzkEstQn
ibKgUquAEF+V0FGPocxDxg2rxIsph4c08Flo2p3jdOUUKvGmimnAoiDoJRdR/5Ek8HoatKDFO6+p
HtxHL+qZAzYWm1hqgxq4KvcvI2l7WnTh5jjnSRvUoPzElFy26OpZ5YrtvEgYRHFeR5dtYqnLMbGR
YuIsMwZqOjkY2qsyq9bAQmBUlu0f+JEkQwmTYkvlcXBlo2RZ0jnyZxniX4Qlo4T5PQJUdj/SbYDY
9R838e7CKcrE7J2OHrILQH2AFmYkHWoc8h4xbY0/XRyvyC1oWNsdsU/93mJYE8AyVKy+96qSa7ic
wdgVSjiZ5qwSk/H0vt6RgcMHvqwQi/OaikwpibxbcYgLHruduhBkqAOujRkrwnGM1U3aK1A/p/Um
HpQI8QN5+BahI9QxvrIWCdZXyppPbG0hoW8AJS/q3RCpQUX2nMOzG/lzH4rRFMJfep2jEVPCTNCV
ou9tj3OGA8gUYOe8vIZwbsWC1Jo7bhV9YlwnlNSjxXBbPgQ0zc3lIjI2R3+khe55ArCaXmobKgEA
hStiLUQVD17Dpyov6QxeZfOn+46aTnkBN5pPyxOiySdEWUiszovri303+VzMqX6izsDvap2F+inG
XuPyAhWRnvBB78+uUbn6OE+AD5OXGHuw6CpoKVvMnW7f9+cMu2FJTJicraaGkvIJFCx4iYcjoCTA
ZuVZWEK1mBOT+M82ivlFJr03X3cW3IZ5A/+J4Xz1730wkuLE0iY4LfZdjZskfZegrLlC7UcS3bmp
f7vN7FCRlzhqHRRTrR7ynhEXrFn8ELnMZGka2X+XA7RK36XWtyzGmxPxiRzfSecbQ9fLStNt/xkr
5JtjbpFx2T7hAJPIZnGVmPhbW6axb0FE6VlyhTx/HivSGvNEUJSXHgvPga17WiIfJNZzsqiSt/w1
zsV6aWRjrgoKqS1ALbEOcC48NhYTJGR6PBWcpyEZ0slxI0atno6iDYW4JoMiDb5MvDWBfMI3IwHu
TZRwao2EfNH52rQAftSvUa8jqBUrWkxa5Nja4Ja/wQkiVAlFo8kDsZ/VSvaBlA7opSPhUXwewn0e
eKlpcUFV5aYVma82nMVXUMCJb6fBQP2TVkq32DJ9JG4Rn0rWwGurG4L+/2X1cc1QQlflA7GUorQw
alp8er3maNX4FAknQGvwtRNgpopS7y1noFmTMSdhCTJusgD/UUWS5v1PHh4Uum/XB1CTbkRikOkF
rVGemj2uEA94x9S9vCNg/5J0y1T/X7ZJD+DMmqQfSq1eCkZwWhpSU+QwDPud6wei64UQmhFRjkhi
hfPuBCkHxaaNsPqavt/cn+juc8iAUtXO61H0Gb33VxZdUgiL+aKK2WYpDk2ZLJAkUJ3qHznDTnIr
Wo4x+FiRW+X32tu0XJW+N8jzNj1hdFYSjZw7BZ6L9iQi9hubuQN5Kif2jzJ0PqDDVuBkq9zWZQWn
ZgIkj0NeYEOZCeLo68Tp9oQxsQRRo8AyXmiVtO9YCY5OtLEF9DeYkReUATrRQJAIQEPnnT6rYG74
k6/+owi8ggnf0oTAhuKU0D3ip/L6GbGpL64opRbWYG/B1x/rqOLzzKqYOsFtOgWdDWZ+6BgOzCFk
xW59AQrY3C3A5hxqV/hNt4aZH00MnSImokXXraw1wFDe0DNLhPZrZGQFloeaQerBwnDAwCCCJsCV
nxPyzwKnQ6oSu/vhfrin2n5GHI/e09tz+39pXM4d70pVeONqao1K38gZSGYBphMwl1fHvhQhHEvP
ZoI6lkiW0GxYPyJBc8tNYdOejeKMxaqYhFara0rny9m47zU1rpwniTjJLZbLOtWkt15VIkKEOita
nLJm74riBJpkqYFd9xqt6Ofl+VfOrFgI679+3NCASxK76rsrjfxY5S8HD+fhJYFeUcNh2pmR7fMn
jT3ZYxy0x3UByvahyZyr7lv6Ys0Um0rhhk+iOYq2c6mwVkA3goVMn+e6zAJXcU32T2yOycHNdnP9
DVmOHR7sIN4Uf+MP1CWFyLZqOOQTzdpr/bmXLkZ09W1qUnfmaE4D/HlM8oYlj8rtOA5baGyfWXk6
ROYGryBkXGmZeMo3fzjk1Q1PTPPVSrnmpnSHCTYF0De8U5e4Q+nGKeqJDnbTe/ZMcQtz+D+sPzQ9
b7IEicL1dHo0P9Fth+740LUn8JlHAln54Mx74p8+qXa5y2a4ynot2pAz6bt7syKLuFj/TVkWk48U
0rpVv4mxBGlWBpgr4tiRo+UpgzSZUxbX0ZXmbriXA8sGwD4Vlt7D2GgsgMGWBQf1avxBOvorHXVu
fgqhjBsWp+R/YEW9VWruTTGkvEXiqOjWVVeKL4k80haCRCdw9IXZE4cNTf/tMu8l5rgXSjBX9fb7
8q2/ZhZI1xISZJbwHcC2zgFJAZdXhOUWyZ11EzAkqsuhr1roMptqOX+TuRqAoWxrhdnQUX5JdQ0U
iq7f1azzjiYMm0OaYVDDzPZDHQVDnqt0z2fHKBKckLWt8tp8QHlBMm1FeuvR+5aAdvkw/jj/0fcw
DhObY8GhJb3r0bX60/lpMgeZbtBhpDDu+W5WQLja19ImAb329kPD3TGgq1YsHHmmSvRYMt+nmZ7x
MMFn/Aedpq+6SWRxpDe5xcXbF43Jb3ymXZI/ObDgCYQ79tyHelTCH2WRpPmuE2BE+XBBlQ7mvXYu
e5tRLwE0CLf0KS/oF9CES9wq5/y42bYBd+RzYfdPNcbnIP0m95dt1xNhFmqA3QgACXVI7+c3QU/x
ysannXEWuW/sQcNuEkV+ls8BAEL+0khw/TBgPGiu1Kl9rwl8d4fjLK5ULh+reGwJ3aNT5JpYwL02
Y3s5rVtjOTkENv4gGtQZRxJ40ukifO6Dbw2/Xc5TmQrsaJaYat2KO77l41fPVLC/jjboHdbHrFYK
zaIrJVxRuvWarr3t50lmQzo/yqqVcehxUcfrxLydmef2EZE2WE34SKoalk+Z2NYRcF702oqno9OI
e00e4wVw1DLTgpHR9ejyDvxldVWxk5jA7ayjUv2HDp1RS8vqhy+Gb8Qz543awGJG97PDLJaMoJHr
+cYo27wB0gAhSaV1RWHQQ/wWox4MOug3n+48V9PzGMySLS6qiu5tqcJPmjmX5PSVv8804LiDDNy9
PhJExn2XFq3UmUwKO1Ho3JBiWNWldcn2ekhSBQE7RTJawWdKh4bpuYFOewrs4s8cypi9yxTd2v+f
2Avm/YRankWmjseo9gmnT+b9UOUspzrddG3jGmjAyLdZfykxjoEYX2ETcWMJsBwJWkQtQ/+a1HhK
VjlfI+/85qO12q0dG7sbY/ul4eUCVh6NKiPA8tq4Ie4S/Xe9QheoBp3AEqReq3MAPTV88xRsWQ4h
6wQA0m4j/hUABIbNak5UVaOjqu5+owDqDDpPlsaIP2/LqzycjG321qDDIGDmpwc/RvArRwZ5IOJ7
b8SEnbMAQ42r//QPHPIbLdugcEAZbp9p/6nrpiMRAmXQu37fFK1HUG+00eQCPgeviZYS2aqPWUBo
htqx/oIbapso/u4YRAKDPMo9T9KFzxlTZmsD/Cor73+Y5LenUalUJxBg1sKJfrQXJ3UYEc8bBvf9
TG8rZ6kcWfaamdyRrQzndI/5c77ndCitUiZOFTbzIdqs5PcKSWn8d/y5sh0zAPkQYREElgfxqGTX
i4Ab0v5VD4LraxJp0PiXjr/Ca5H7ph3cYbx0U8GRxHINflnMB45GeWdvES0Z0giKrgda4S1VDH0E
D70klr8AQ7/wTFV99u9BV1V2r6tjgJ3hHMelEnLPZLpXJUYpfuPG/jNbpRjETOg3hd59GS/ajeHr
vwZyhZZno3h5c5VeR5pqjfPI3HRZiR2U2wxMmWwGgsnjOly9Gwj0jyPYd960PMCPxLzyoMfo8eJn
YN79oQsKyV0qzDyhFxI7Xf1JM1Tn8tPl3jf/NUHPvS7sCgHcAcB0OO0b44bNMwo94yn3euJxBtlL
pwteJ61cySS871P3jjIE8qxFjtA21kPooV/N8HxEGdNyL/6zjAzZTsaYuWa32tLh/OKP5qdaytfX
beuRG5OkDXBfcCk8rTVWoaCFgyQ6eqWv7on9aa+P7lTjINjaYFohxYFsbv2mPCjbFdhWDMIh48JT
khTgki9e6nFgMP/aJoWLa0eYNjwFFjRB5dUYEurur/I1Y6O3YBD5pj7isS/G2V2A2b97Pa9LCFcZ
Bdb+syW4iFqUMs06zZaP47S+5ygmsj9fIMl9bU7fCIx9528fSXb/hwgPizm0PuPmshaLXTA0x1R1
bY0bNZszf0WEQosKUqIYwAHjxOOc2pD0Fx6vJY392sB06458Epy9lilHFcBvYP/awOfc4x8CTrur
y1BW1nxWAZH01TC9NsyExJumC6OjXtbW6EtGmf21ErVlZeAWaLQ6hmUJ9FAg40NR99f8NZafGIYj
zoMfoCZ0sVmR4MejYkvvhPjFAjY46IFp4/Wl9i3CAtX0tczFzxtixeANgeoxKqaJ4RHLfNXnCSVv
NhShKenMv9iFIjd9z77YUynknDnVAjtnVnsY13nVxvISMvZoYaoMcQ/wyvfLQ4l0iXBMy77+7FpL
1H2J4wfL91R1JQFZChswUxiZtfwtePUFEX12omlgA88MIPq3fvaAdel3iw1pqDs5Ublh/HBzwJQ5
CYxL4XBJabVzHg+y+nM40NScvUHDjxaeJxqSovQ1e5tOZFqCWSw/x4qrHz7wayU5KKp+iK9h6fvg
nDsU93ViDuo6CzpUoPXimhNUnnuooYGureODaXJPEHjBGffveN+sw8Iy6mj4HiHJB5AS6RUmbxpv
ZlKjozu8+XJeatcc6gcGkTipGJE6zcUdLee6t2KcmBqt1i9I+ui5v+254ugz3Zr9QYAFbf1dq7Bg
V7QvH/RRKPwTHiKqKPrPCFOCO3mni6CN69Z0OScbM3HqF57puToelR68JQasFlV42ucUfpaISXAl
JxSf18+DY3RmrrAXX1mpsft6jROajev2d6u4XjgOoyc9bA4xy5/6rHv97IO7JNrl7OyciShhRZTo
6VCF5fX531WsHkqw+X2nJZ4Bs5pdFOMaf+Hyq5KyTPEVNseDDXdWObf1ehv6WGSrByE5FzEcK+VH
8BxfOY/wP2bh5+jfevsz4kqLgb5t16pDyseaRE/jJMTq8LwLS3zqaiQ90tIw1FjMWd2W2rhASXW8
PJ/3xhr9CLiMXhWxaKseG3fP3PXVTOUTotizMqBqMklp7RzLmKSnksdvT98+JxkLdqpkMWsSOnF3
Af4rPvmZiGaB/7KAugFxZeN5nRTylvEQpC31yQe8IIfr4dVnPdDQG5tgVAi4QYUhE1/APIuPtSX0
Z3AYQZbcgXnWGceY18hQD3Ub/6laz4eSmIRqdx/i7sDGCCxVnUU8NqEHKknf+4m9Hwzyf4Kpw4y6
k+Nttdl9kINp69uallPC6CvPn2aBbbOmnS96dpUdCFVENzo0gddDpzOzkcpKScEOQiQtlidEdJye
sG0ix0jet3LFiE+3r506BbrIPAU+Ssb2ohkXMFRNTApyW4DovtaUbwghLzM9jckHipuLtPh6hAAs
seiG/H2GjE3BNWs3ivOyAdzk3R6Qgddk20mHIlTqX/dCGaQNZEf9y/gpNmAEgglH7SEM6b4eyqnl
Q/33YyumqD1JCib5bQmbcnwb0sxVzNY/+whNI+sxirdGy0HUeoL8OGkFZLlgNAgomppRc30lnLuU
dN7L1Q4wgcdYMe8Ps47+oFR9d0llXzsrV95ZkipgjrkwHLpmX8yc1I4dhkqVnwLJUgm5fW9HBo5q
IZDrUhPEP+sBJmcjDqjCL/DwPI6nZMT9IPFuTZIduNYAH1Xo4TiDovWJusFDexElRfaOdCFfD7WO
ZfQ5Zet2dv+zdNf1sPpzyRgWADej5TfMKyCDc73IL1qWT49oU5u+yKISj5HahNpl+QiWYGhYDGgx
d/H413NQqtGSNjtqP3FNWjP7mjGlyDtjtq8rnvGR8CmwmdjjgaiOre4++ogy9SPTME5EVksqHY0y
5PS69znMr2ZMpUfYLVIXD6jYYK7r8hO8ibF4/WwvDNnWTvCV5cWFytXIDBbpU9iRASgzQoWeVEAt
mqut3XHtQ+Q4wqRG7xQ6neVtVVsW90yyLBF0MrcCqgYYKKwa6k3bl7R4DMYaeKYbjq56ioMd3ten
Vg8G++UqRBoY4vi+trb3FfsehXqNIjb7dLk6NaOrEUv5mTXf2t8p2bz/JHixRl8QCb+G/i2TAfS9
0X7PUdHDB9MLkoCgLyo4d3WBI6cSSgMo2mE0y3a+lYQCTzMGzG1KSJ4Ih4LjQZEkM5BdPUMmwVu3
e9iGcfgz+vsoMg1NqeMIogtxaRKSZD2bSAssr8f97WpunLAb58RhY+5nhA4U7OJHyS8YKRYY8vYu
2CN5SdI89d+UarI+s2+SSrGRGMwYqoD8167tIAyURYcm7XE9mR5dQ2IKYpJsZtGO9YZCh4/I/j8e
HZGTth5QLAdXE8ClmD8Om1e+vWcTlw2p9DiPB40Awdi5p0KiUUzTLYZE5W36mNpRoUbwUIGPXIL/
ta/MJ5rTOmBB+7wRTcqF/cmyVw7+5WBasgu3qYZab/HDeY9/ImpBqp/M391sg+HaWIPTy0gb9jX2
zuszFuLXNQ2bEVLvEJ3YBBMVtHOYPakQHwUJhbknFZNgxrDPhj1jC7aBl4wiok7WgBfG6O/qf3e1
TQr00z6QnrMI5hx7uiXy8Nf5p+ofm65oJAxNpGaEKhx+vtWtqvITvgwjrwHxmG+rLG89CdJRwP2g
KFqYOQwVwUy2l7bfHOg4pOFmExuC7aCXN7wRuSo8skqPqrplT6xrZWjdmatM6ssRvMvaTrXTF824
EnOt2XxDJoUmyoGU3kut66Obk+oeMeooZmqvsCirPmiRdXd6f/VJXuW5yfQomUHRFZXLp/7TtXdY
40+nxmAjv7wU7/q5syDIn7RLa1odUaan5oBIxavK1pNGLvEmUO292IsnOeBglT//Dd8WVLk/gXpK
YzYSHOB72nMsuQOQTMnPkS3y0tDt6ygiToJ1yhwvXci1C2rbd7rD1wCJEopCg/l0ttBc1rP0fTkr
c0hMpe5roG/p/FTMf26Pq5DFGoKpqk1/lCtuJghgndo+2jJi0V2OV+S4pCGTKwWkbmTG07I76Bxi
J7qvcYQj97cD3MO0Z7T3OwafwAQZZL9ty+91/vPRhqQESatbBh8AZKx9SeOrTT1zQL6Uxp3tYzCm
1ycrO1Ls6Vsc5JkYCNRhkp2MRD9m0/8NtbK5CvNOZH85Rii/ihd3OwPYx2nDoAnKoCo4tyZksNo8
4fp1yr8lu6yEpQPVWDiuZJNSJmICj1hxljo5+Ka9iF8I7X+HzZ94DhKM3j0DRwUPI9kcoPf3cW33
XYB3KGaxBl2NyZ725bvfGwYzWONjWa/d6uS8baNHXAkpqLq/gUPCCsQ2loOF66IIzmBllCkA1EcI
xvCuQLWWEeNN72gg7GSpLxoVx4sbeEWGG0Q8HSoctBl8iyY0UFL9Eu4N70f+D+gDVuEMdptthTt8
B/68ANUO9oN0gl541Qpa/Fn7gesF8Yl3YytjkmTYYZ/1Ykfd1DtJrvoU+KVEN1rg4KDP87Ccy1Qr
jDuMgdmDvYYdRwsNEMpgp+8eEo0QJbYknrbuSs36Q7Cn63aYTg9MWKvjWp6wjbK0alJ9DFy88ZWR
4a7eKaoPuTJJoLgPJVLIZfvxolPpcnlYLU0GgPaLKXe5GfQu/lFrDaq1AaJig9XdoLrmklTYcqDU
o/+aQSGQLofth+qtiR5gFD4umA85E1bq47K1qGrTx8l5zJI9Fxnim6CBEJEDqPO0kitGfvNQ1qi/
Evd3vDNBhO/EynTI20nOsQuSAeErcmbfCuRUJ1SbLw0Wu2k2mEgPp7XzOmajnAp2+AykQ5lqzBiL
KSCcTl36a5C28sIzKhCDkW7arxU+eiDVEWR79Vnm6AWyj72SEmftHdnQ5oajtsfoaeS0SHxK0Q+Q
umW4JdGVUZSRc9nsTYsOVWq0IfIYfQWg7UHLAQZtHSJSJbkgdtwsr74vfFCPdHauH5LLOtzLrsHr
OdCIN2pJ3j3KEd6FRclVQp+dy7qKP/fzk0/hpsbC3zVwawnXSKNqiwChoZmRBiuFQVK2slNbBM9n
HGQafX6T5d6+POEtQr2Io+zJx0M0AuzbCBjmZkim7rJhB5Wlmyigb3freAbR53nZb2nStzEIIYPe
5b3DvkPexsG+6WRiju2j+CAe6aC/xI6qO/ax46ATR4huYgN5taRGjn7Ft+ssD0OvASztVZ/UpYV0
KSha4X6P7kLcWMygQvV4mFidr+aLlVmrzJeUDzgFjan+or5dpceacgSBbz/qRlRmZ6G0TiAXGCoN
M7SkPXBtaCz9T6rMnTGUmal7STqCPgj9rPYdGNG1fzZhM3/lUw5xNRNAVDn25MeR1IRum9LENS3y
Xp7z9dkSdOQdtroGVUnK5oXXFNcWED4kimMJpGr5unZrsaMkFjZLt9QBVhrE9vpi2fbpudGSAsFl
zz1LCKee3cIdiiFq19TaAW/0J05OdgQWjS8/cdYxwAtt7PgnWaxuWDiR4UoUdKvl2I26Z9XLMYCZ
khN4cdXm1ZzbnYWbTprwXaurxr10BNQTzaQ23hJzj7vRroX0QAWLG0Wn6iHuzLkivgl9GGY8i1kn
UxopjVBSKKom3u+0PvAhVoJc1X+8Lf2L+X2P49JuouikodWvNnYMI5Ken1mCRy/U10VjAYakcwkO
iMWPwSI2dOA5Ep007ugbkmAY3/c6gsnsYFmrT/Au7sJUa8QA9GSa9arFsHJHqoAY8MB7fRo4QBOR
LrJf0Mp/fev2WMT2CBC+2m0BTc526wDt2IkewgrrOsd5RuTvMnqy+jLDTcj2F1RgfiVzo9iFHcM+
Nm0Zg4BCX0Wubd1sSmEOzByP1cxuglNMZggkoZV3oQYmWaW2oKLxCPWWVCZmkUJ72s2kFd4BcPGQ
oMI4eUfqJlNwsOu44L6mJIEGxD5v6Go3nH+i+x+GZef5lRaFfAyXsjvRAbz6I+AlsPVAY26lzjDq
srXMNewPWe6kuTbVKbjNxeS+qH3FxVmAQQteJFLL5xUlwDsiUA+b83QdR8L/xPoxprTtbsnL+h7N
yz8Pq8zjHMO7cZV9xINFxPsGxdx0Hg7qlBNWLc3hI9MviiAJIUJzfWP4vaYBoD0cAfOVPTf7UcCd
b15HF+R3BeodWoon3bgaJlAJsI+0oTxAtkEHBhPB1FnLbumRfOjkIudbQNffkuzY2br49ZCuxSg9
w+wD1oBq/NFRYVBHBWT2PtNlTjrkTBsizZtHe39VjOM2ld5u1u8rDPmGmjXbrAgtYxYN4VyemOba
YI1DXiqbGG8MjatwYSXmqmJJX4OnDWOgaFKyUn7gNcG9Yl/5ezGj53jW8RaIoMyG8uLlApc8t43x
OKhntzs0i5qau14Wq5FMIKgPSQIK5blKQs2OzeDyL6BWVqBa9TRTO17Vi6a85B7v9fSYsKg/1MYj
n3zzNiwGyYNoAhyXemGXjsKOgZpAamEL8GOj1V1C5+7JyUZadhYiGromjJWSsqiARJPwoG833p2+
uOgmWLGnwjyoJabsCZGDUQRr/JbOyS21LjE11I/+fTvDKPtIO7TAfGuvJZeq8u9v79NdCDdzFbuR
Gt8g5bMURyo6F00IbibzFaEzDSrSsBCyCK0wOiEzmcGlTtloJdC+n+L7b1KK+qSefABLZVTcnRKJ
BE3TMmXnGfHA6GPFmP0Pt1z+RyyXHe4uWc8aQ3QVzaiyHN3ODNP4wvY07tGPIDSbh6K/OBCWc79z
6oA03BwWIcKwiRkOUlAY7AMGt/MXVwL1yjexGxbFRoqjMnoTRVOAPJ+W/DUt3e19qEOe3oQ72XzT
kdSO35HxyDs4MTRJkHIVDFVjFFLi0MhSBqSt4w/ap1gb1BPQViJBmv0HWUAWA7brd1MZiht8FE6y
Mxa5sG4a2FD9vkTWqNJnRN5lvqXXO080AtTqxEI+ys9/d3yZOIM7JPuki8nhQ1ElwoY1Y7pP+m75
stTTRyT/2+t02rNQ4YZmp6Fb4GjqqNaadWpnhwy5LdgN0jR5auwpSDpJibTJ06YIZ1sMtsS0TlPB
ZaiIAiu/fgwjaHisSoazgcCZbAOSWPY4yt6v4F/feNEuu0xhV12nwSO3jzHN9tg1mrrNaF89taal
x9rnu/RzI1Wd9DljaMppxazNTZPadkRKLkKaaumdHbpCRN7ToY9utyfqn5AKxTDis3efHv/IAHyq
R91e6Mh9twdde+flZ5OxtmiGWUY/uFSFLDcTod9yz2MPNhqJ/uANE4rQKNfQExCZ9H+wjZJ0g1Ho
rs1NNvAf40Jx6qswRrQEDC8NyOPY8K2pQGG38VLsvIRcNj0ogsiKX3pBBP5hzvu8HESCPBea/8Xk
Uz3dYfOVqCR2mAohGGWS/IsXqVrbATfWxKwp5Xq8aXGDTB0+oJHjswqNe1RbXp7jGNl/MuS8Zf2y
d1wfdFhKxgkq+9q8lWZ+lRZ1ZlCt5//Zs2TgAa4lEyn14DghY0pQfZ34dtXED8mwr736Li/Qvkn1
Wdf17NCVv0fVZlcfNI0TOnkf1Kr22sGUgw/P6UxsS8KDfj5IjkrPioHaS5M56We4z5mB4yYoKJRw
nimUeV274N0edqV+e41bYzmH7edFBSDimYtdC78ewj17EJ+FyyeGvZBG005M4IxdoXNY0ARJOJ9W
nryXktBKdWDUiFqX4eUotkzM43XpfsIjJAcjX+j9Z/SpI49otLuauH9ueTjpSmGMCZyTA1tWrmD2
ooXskGB+FrYzu19AVTmH1q6xlnGb3LkPh5bDyaNsy5AjGc3qHulmNNm9ViGoeWVR5dXZj8Ur54Yw
X/1ccmiGJgc/smrk19Xlvxh7BnkLLDkS4rxWE5M4WRKas2V9++Yk2xfSp2Aue5C5Qu4ZYGzMwy7X
sfF+hI+LlyjOUeyDqcN26uMO5dRa1dx/6xEl+yTyZTIpPdXj5Kd4CjKU7aF2TdYlnT2IfdXFPHyx
saiLPRm0T2K31ORiJWhsEdBdJphazZ+BH7a0LJn5M2oTR2EXjGAyV077JGqlJtiqRYosR9A7C9lE
oIir9ulQT3pwhoUzGiHwctHUcjWNZsYVYurkOE/4ve3RLiicGi9HF68ETWLW+ACO5sCqjciQcqMz
dQcXMzDNWHLCvUWu+3R9AIgGf9AqsvnclW+W0ef/lULUA+0TVEjhjoQpGhCUCNHRw+YJ+M6JKgUk
P6LAxaGNZiKAVATJdlVhPViQA3uNGhcE21wP7PkbcNHEp5KgYn0WiIW62Bqy4k5KhggO5Aeq+95u
qki7NR/jDojRfxJM63w4aZjO34q6AptOI61zxSFaND0ZHKoNHd25HoAMN1eM0myKPg8Q0VJtmCjT
S6LQo4xd8aFP9irbvf0UTjyxWDefMdrNI/J5kU/MocGvKIzqujhAV2tLl2q3NCpzHhIJMuiWoLiN
l/YQzoz4l+fx+ORaEALQSXhh79fWh2QbcCR1WnNhxGlm3h01ODwzj8u3q/c7ac+voad0GXtF0tjU
2OObIJkEieIkGHL8ZbbNX/xTJZEZ3VM2xY/bvnjeRXXxkCPXSkQuehepmnVwaIYkSG6OgjGiTiM1
KTPooEo7L/Y4ovNARx1nJfYGOjDnR8RIoufrOm90QUSbBfBtoi/VKm8nXGmevHtT641tFO3v7xL0
RNsIh+TEq9cf4CkVe8mGodiC6hL5YU7brQ7xxwYwR1zoo6r8aKsWpn8a8MF3D6XTH8s8CiT/vQ8n
y71i5wU8uIAbxEN1PZ2LwxwvmYoIUjA1BjfAXoQEzLBlt9g4l9lITvLbhzc56xtTAaMzoNQszLlr
H573zi8NgrmQuN5Y1XhrSLPToxMnzDR/a0JGYEfJfUG7YOojoNgotBn+gVAXtvRChXXZZUI56pZc
S0X+uH7SYtzOUFsssMnl4Shu8fNIt2YV8Lg5Bn/jU8cF7NEYhc0xHY0xMpAjZOBFUc5YbkMncE3W
mYtjbMPhggufh1H/+ZCT1yyvFic/FbCE9xMMUEeieeGH/qoJsvcZv8jYOLsqMI9Py6N8iYSDYgbt
g+1Z2ORcfQfZxJencJ4aGtpIF3QTTD4C8n0BWU+44ZvewmrgECWEh+o2N2G2BXnAwvebYK6YsMj0
uekW+1vV/JblehFAg5slkKxUbEiEtG7owaCSMv+BWNaEMDbqFFPrcQlgq/CWKexozmVhxV0cSln+
m5qXbmJEeZxZTfGy097/8ktiSjSAu4RWobGBE766O/2kWxcYCvTYi1F+YBzWQhRfWdkzVgWX3fKM
RN6RZMg5sFKhh8oh7tktubj/Dtqdvtq1ViyxL+12Gklg+EwvCBdHcK77AryW30jhxbV8EQHGciJT
5v52/YOLOd3Al/zuywcL0xMDt01ESxDKkXUag2Why+LA8tgnpz3aJ2GxVg68IzdBFfPmEM74d1Dg
+emSa/RkiIYJOkEem/kfY+OCbGzlL/eBkzt2bhPsMZ8QdW+x2QHKiGHIM6vTL0pEdxrq2Fvmt37v
hdoKdELQZiL2U5HVO80HnCxM7tBbwJDFsSg+vYGiPOQcZ1WkHnunw1mbUGoqGl4fDD1+8CAe9EIM
y8y1OS1pXzmNooQu9HZfkH/SCaGCC8vZsMYVdbQtXn/7RDzCmIDDDe57X1naCQXT2ryqgI/D94FE
tUSJF/qOvdo4ikhdvddUyAePlaKflpaax7nweS9/wtPIcoOgCfg+eSynD3N5jQ6YbGUv8NRc/s8A
5kmQmWUboVv6u8H9iTvpiw0UmuH2CBBp+SnvqYU4nZ+4bwO5aJcFyXSUbUDPZIvQz9rFKjed2fJd
ixOFtu1KxMqUX1jK9qxlcr6e98+BJyWSHCJKWBSsVaRyD1QDLtFzrkDuGkzhwQN++ymlj7GYelY1
0NKMUc9+UFhg5L77EpqSQCupo/H0TOmsmisSQpUOTkoAF8NwIfo0pO8o84qm1LHvrJzzr2hFpaqn
tJzIeFCNtTDkXDDhZ2b96lNetHD0lZMol5SqSNEi0YuxO/2X3d9+fOoH0piQN7YaiH5MJ4SvFoeC
kK5CQ/GLw/2vTIiTdSDHtpT3OgAa2MREg7bW6+dAa65Pf+ONT7hkPbr5gFhmlXvTeWFEG6BPFPiO
xbTF4nwX28RAwGwpyrfLUyzwR8Cpvss3EJ/OdPw2KokGJQUI/leajkhGnQo3d37F9zu0QWrRasIJ
FZlKbfTy4BWwW0u7zxBIlEx8PCrkDy0KTg7fQUNV6NriR9TsGm0TERmP8CfZfF92mGO9plAewvVr
pKqAY0IWwy9l9T1/q7aRFS0Du+p42U8puS3beAhfXl+NBbUbRKdiJjb3a2qw7WLdRaRbUtsSXe15
2H1mi62Cji4CPjCzWqtTaBC+F0vjJZwd8qKJBWzWRQcyKDdJ5LRL6wVSL/jM19YQhE33t3vUBa1V
LPk+RySMPtd3Syu7pHnGKsLqYT2mhnMcONJ6hIwVEs7t2w9BpfHmSIHyQ0pk6bHethpgH1QomX8Y
wKFZV7BVkjw2IMMdcn1jCsVuzJUTY9TJKxafh34+L4QcdPzE25dcbxaDG2iVeAARsgvhRe0jjWhQ
mXdX776jzho7h2kaDnvBAxLnt7JMTRs4mTkSi6+NdRyqCN6WYZryroootQ1o8Ehx4bo/gmpkELDR
waFFWkFNCb+gKRwpb2dZ4tTaJ0ZYUKp0QpdF0AeZN8kviDNTrEZOiTk6IIbUw71G66zvmmpqv53N
SVPYym9yUAWNRlvkB8SMQw5IJlggbX+PHaHGoPod93AO3zN871LtU0Ln2qhiO8ay1LekrEQMDLct
M06i2+gDfVzRD5QD9dXN+lONYvfWJe7tRIWeh77EUpOlHyTCmh1t6uYu7VPj0HTSkV/EnLZ1NfNi
r5OToP4vPzZ5rvwlczTJMfZ40wlw7S1ij5tfFiwprFwsL9fy+e54wLP+qIZpseWlAW5VCatuhtph
5KXWaBW4IYj2nbZdRupnsjtwve+qjCo51ihX/vSWoILvm/zx2HfTDlz5SQBbgqYYIHQyv9MRA/+3
Chf0jvhCzwihwLcXI7uSxSx1DCFLhmurSfpfaVAxDtS7hMDZ80xhHhk4GQRlGO+GWbjLjAWX9Z4r
aeOnbNuCWoOv5S9kGanxEPpydOj3NpT6W2NZY+XemkJ5T0dKh8eEd5l2crz4+Q0GdNyYYWwHD5uG
ikAMKIKo2X3UuIciPkt1X0BaQp7Mp+HvqtFAmrblnXMeVQU7hCEodnAlWTVbmQN67dMLdcljUsmy
5nFX/TGVlLXXK9koDlHnN/sNjNcBp8CS2N1u7RIvBVFQO6ys6wZn5AMJ3SFqa04CXi9y9GUDrp2U
QztPi5aKPlej5Bm/RXlrSdu3A67be5TOhB4pkhj9njYEnZgt9Iff3xSgYK9HTTcS3wJvA71J4J1b
xAKAeFIj9eMcogPrfhcumRK0VgByq2NEhnSTNalalkAYatvRszXi1G4GK0qLSqkpL66KBy9V/wmb
05SHxBub5+s+8aj9YOLQYrNh5OI1avjCg/A8E0yRoj/UyHXzPh1xUEXLI7bMcBvG/ni13K9Iw7Y0
+UwI838tM92eXBJSIuX9vKMB8s4TCIrYs2moqOX3kHxNeRpPP1dkTHHuMARg/mK9wHgP+35X4wKB
eEMAsyf6gmpeflK1E1MmZDdLq/IQZz6rNEbFDe90YJ1gmTElzBkqPJEEg7enz6arRdpHU6QSGemI
4HQhniCqkjLPt54ZiY4/HSiIOYi0nXfn8P+alO+T8LjhD9jEGg0DmRKL51XKwq5LiZkD9OKD1bxd
sWk21Y6BlE7MG2cZwqBYG8Njs2XxeHMwRwj2kcA0PFmJxCmoxH+H3/O6gRamOwgCVVRm29RhDf/1
+/8FU8vEywsuuA0iq0KpAEB82RConsmRi9wyXaHINsG7/9Rp2rWBD5HP25FPmyhIUvw4LnZ8wEqR
Ae4S95VFrtaFavJuJpsnpJ7VOFIQQPdKHMiPoC1GcR3HEHkPS1SQSBDSRIt/wMBuUFdi8cvNfhfL
+0apq4dPz/sfu56s0qo++Pt+YJMarxWIA1rVUzCB1WaRAwXg1ox6Nwu0Q+sPpWA9+nZSGsJZH6IM
2UCe6cHw71wN09EKycp/6E55Qlk4WK9S0meSH1fNquDC7ZM5L4BcHLqDD6eVlzTROICVRID8sqDd
lFi+aVhNZfc6O1JG6/huwD85Gm8YyaOQAfrhwpPl5uXGW61Qqra/bG/0bvxU9pW2TrTQGz8++ciF
EV9xmEa0gsFDwIkwIm51EsEm04ePV6dsDUTaKr2PuRUHLmskU3YYIxzs376BSSiLOtdI8xXtSc1q
zTFIy3JDbbkZc6TeU4GGt9+JMNbpfv9TzBETSRyzOQxna9+9whrJu8SqdnFV5GfCPYmPyh5ZNIQa
+LE8h65SdGxrNtqjKXTV8UOBEw0GXYocW5SXwJChlSeDDDhlsOGzJwrbLl7Gs+4RmTrB85BJaL+p
5/AAhLRsiDgkxc+5YAHUujZCHyiKNj8N59KEBQBBunGX7MWseDCmTlpwrAIljqurJfujYdSXIloe
NSt84Son/eu+iYjqLQugWV+9102Ml7OUCeFCOhAX7jyp/7JU9BX7v7RgFOn+bahBB1HrSX8uVghN
/T2veWCDk2TAmV8JnQm7rzP4m/moHP2EudJ+GnnWSQeh+b80R+hvYBNzD0gXj8TqaC8YDR/+x+6/
tfMXO0Zkyk9BDBp6ZC3bmZe2rnvia3KxQXamPZOf7moSUeWdfBneRBaeGDJz6iA2VvM8xX7bYNPq
NkWYhCHKAPnofQPuYeURnlbmlSjPWcyZuIb8he//RzkXWbL0ZetbsK37E6Dm2Jn8+9XadKr+vzKH
tZmiDqtvzumzpvfewzFupeR/djtaaWsSlQNlNrHnoN+Dfzbiz0C+S2ZPlD3v89CuMyuvyOKYVDhq
M8cpslU1aKkgxhW30v4/XR4LaYQOP2NYKcIBZHeyMqtaOwhP3a7DKH34/Q+wYBQUULvYL2VGvWm0
JgJmUUnrFs1G9a+8djUg48tWc1WIyEHQq36MlIO7Nu24/XR9hSXHPzKftbzCAefpHbwU0ETJROiD
RWEKiLD1XnSbWhl0CU8enUZhVD3R7rMkBabsGRZyAjfzsl4P2oPTVteMiAsFVWy0nW+Hx+/g33/C
ZEtnO9EteGyfxeXDqrwks0tSXhUaNdwnrcJAr73JQbI058sHY3fKgmknLqo/c0wcc1Jwh2rpuWxy
hyegyoeLt1s8Q1EO5v5X9erbOL7Z0iE8//3iyyKdh7BCeXWsYkJMTpDmdi7r5+MOM8eXFjLly9X5
32VN+Db1xjvQJ+Jhf0Gyif9aLS7gADwZPfFJjRJD3CzXUZCpd0CB2D8Dr9WdZ6vAvcfEsu8tqKyc
KWwffl8WIEKIHDyCiGCZ0T5zACg1HV48pm9HACAzugwdjrnXCpjAi/FQCUHPjabcbbEew5dBA3Yx
ACP1ykj/5ZHjH7xPh/pS7kQn7Suefk2rqzImV5UA0LpwprRzEUIKYrCN/hsvYmxcs4BWmQllSbSm
9UcK0JVd/mj2H77fE/KAQNbmQrwRthQAM7FMrohHaUwC2wKtT8H20WiFOB9llnTz+reoX75rt4tl
hBFMmtULok+DEs/dZHDaOBek/2GCqmfImQKOqvxM+6CUPEK73NNLH8oWQdV+ZaEmxAYJWCAKoPdz
Mojh7lr6RxHsJnAYTspSqsXdDVqhdUA3LNSAvqSAMK4vjV83XMkDZ2CRUiisCQnj1z8hCvk6nhMq
WBs8QZJNw2caQU2x/KK83fYGZksff5gN/NGp9P5pkopqpf6JzjtFZKB17UKI0b5p2W6pI26ojpQP
4p1au1RXxexbZqWOAto1q2CrPoEsYeB5penp5HeSnLzjdH87O+qG2cP1biOWI7bCqIKk9agBVN4d
7laJaMCmWmIZ7bBoeI+MrbER5njVrluL/hC8CwVjxBnubPJiM9PzGGyz0U/zwlZugwRAHGzMDh1P
h/Mbq2aInprHnlWwWm5uDbxyI7recKA7e59ezEYebqYYS0nb6PhTehsQZcC1Ljmbll/XB0zm9vP1
vb/t74tC+foPa0LuJxyTUQaRC5QH38qf0ln43TFpIPbZ7Xqe9i2/KYZMJ+0IRdNQkycVE53mhw0B
MZGgCCOJxEzXBQHg9HmSjDAeO0Y8abo3Evq12kASkuoB1XvNINzuBrRYyT5chrodQRt2cxPsL665
nealTXhiHWqRgFJtsTyZZtXWOph0/dpmxaWZzJ/0SD/yw/FRm2tIJxxsG4pe6hGRAKYy/6YHulM3
wrcGwdp8ptJhCWuAI0kR4tF98tZCHiSuIIXsYq0CQtqFB1Ajt1RheEwLwVoYi6PBx9z2b6f92pIO
zfYarQkxYPsOu7bLGZ+RoL5M9FyZjKK+HB9eq9NV2tadExnqYbTTvQ9NefjrNcLLiVYZXekBxMb6
wWvTFQ2capRj2ZPHqAdKMui3WA0yHTbuiDNBoL7tqR2fiy++DOtRKFfixAPzBIZEobuc1H+6u7/4
IxCIGg9xoO7KFVL8PbFKwIwyWIS91H7O3mleU2VrdYUPTDSP1b/776t7PnFCwnIJSlFfiMt27GS7
vQ6vdZWBcDTGdjL3D2VKwl9UiulWwuPezycy6lYJzN5AszFaszMozVKOP7V4ISz32uZqwsu8ay0M
cQzeRz+QdyQYVmiDTpOF/e/VmTdXNWK76bCGier2dFuUQQVLf+xwaJPCoTZB1++m8hvVKhlVYUH5
Eg2o+uM09qqgjdwR7OrFvfuLXV5+mutnbD2amDbvyKB1W5/rqrA6sIJxVMBDOyqW106kdSKQSBz2
/YP7K/mrxxxkDeYTBSyeGPkwHFqz/b9LoBBusJ5LrAMZsF9/0C4SNs/z4y6AsKCIzC8ArspswVr4
+twfPAEur2BvBk7IDWpNawnvGYXILxzDJ4pH1863apXRPJGsog6EYIrZ3mJZOGOpgxIm/Z0z+nZl
svltKfIr9OvMSvIlKi5wLObOMRePZbtDzCVFET5nHYhHp9cbD0IBoqiKf/GUhfuJZnmgWZ8OxheG
TLb2nW7xap8CMhOoTEK5kUsu+NXsms21qVR661BZ2yCOLJMC8lw1by266yUMBaGly1Ad+Wl7JL67
kMP9+MhLCW+sMPF9n7Tfw1jFCNS82bzV3yGOBRSIN0qBNFpmpHQzXJ8BUmhfjgZuU6O9QAtlDPZH
diaspB93tvJmTNif2myXHmcixTTguyRVKdrQp80PeHVpNmwoJB1ZSXKTK4yLg4AsBmKseoe3cWqX
O1uPPB+SaOB5yjuMYE5kBQhHohi14+eof7YMCcEYMZmHrV2H5kVP2ftwB699k7PdgoTvERLSptFX
cI0KtxF1LNVNEKf8PypSGqHOWckPfJZsCnTRnTlGATRA8npf+isPOF5mT2ZbYDQkdPXFmuxLVnwT
4wREBvnQKc3AZdJX6ly3/hLPZ74kddkpfL8rGip4zlcPt6TxHAq2PYuJg6NeYpaypL9Ym7kP0fNo
gEA0+yQkm7YCqz8pySt2O2y7BAWe4H070wiiPjcTaIGQMR/QmfrEESioxDZ1zHvGNudRxSK0VBYb
OUcoHM6DsShEVACXDUi7PU81usW208u2NhIEeUqpSrQ2nWwBoq4Az7nv0+SzjvKzwhqAl7xgM6hJ
PdNNCNFaB1PAGT2Bqd20HjYe9dh21D2jrgDmyQiCAZ1051L6TEkKYPS31dn/oNicvArT4JZct9pF
RjXtV6uqsbBi8tDXQTdouioI9q4tDAzOjNR7IdFOzf+pnJR7PmSgBFxqRhLMazGDVfZIKuo+mh0O
884gFe6MI/pu4P7An+p/fmOCc5WBUMiI0Bnt38jUwpBWNjnIOnxjqqrPpyX/dcqM3WHF8Xsp4+M0
RDVhAH/vRt9Wlzev/Etn+lslPeAZjbGXqfM1NXzUQPSoQq6AObaSdFKC7n70/igZtx4l0teQip5r
COnSTi8Aj+Mt2b+wpAG/RjwXGsqmC+OHTLFTOOtyQ5zHQnOsfKAVo2SLKACNILe00S8YpbVCh/QJ
aHbXiJoAZsQ3t5jPwM3zMk8iSmwDmEirb8G4BMaSyDS3A52dvM150XVfqtUlL2IaFuVYA38TkYFc
/vg2Tt+i5NulNgAtf8Mz8LZA2tbEDZXYRqGvk/ECZlMtI5YR7xQqd2pF/7ll6IGkOAq2VPDBp6HK
QoSP73nZyydibdiO0oRwonYo693zp4EZC6YTyRS3B87Ni6YZM5Pf6P5t9SDABp7nJ6Ytc9QcdHFa
nAntlJurUfm8qLyetlhvyO2f54HtcQO/QUUbRfDNxc2jjIP3socnbFmz9as/V6CTC/153ZgzU9KW
3B2fuDvN3qNno0fgTCMmegQO1xIr6F5VuENXxlxz6SMwd7QBqg//0TdQGeiIw3zuUgCs1O37hZLT
pHe6n5kThJbB/krY+lLR4LbxxHrA2q1PYE7e0V1ddeStIhzeoHcv7opTaXVyhVm+PvchvTh1aSdX
teNifHAP0OyW5KdlaZEFkrdXpdPIjMrbSZRZsQjk0TDdAflnrWrCHJWtflm24EhQyIj8Iesv6fSs
PHorxX1hWRX4Od0m1I1Vh9lbHfMrnKTuwAxhI/XfFEKQ/WigUb8evv/eMp3qielOe2mKb9FwELd4
2Z8r9rvO4hxNFCkmHAvBrdD2KZSJ7pHi19wWn00NeKvfkipiNjBw2ag43LsLXYsJmkInwAWRQ0he
Gn3Yc6ut+m6HzW7Be0tEkbpV7fy0yeH9CN5zQ5OQjA7SAquW4P4cwp/LatRRqE37tMGsBrUH8xN8
CWxSIOmjYfLEaNE3reIKfzyfxr6TnAbHv2nDlaERXrmTaOoNvF4L6SZ77m1VtZ/eGQTHrgKLFp9w
MyHrGwNckl+axPNtHk00CVfkexK6s/csNh2ui3ZrxuqHRzklroGaO2ysGJDqU7cSEB7KlGl37eSl
TItEfY95//c2LbaHWfSmOdf5wE0D1qe3g1TK8OpVbV6/OYmzPEP5DsS5dBxrkDy/5QJsRzBDcq6p
f7JRSdgTr8hO6YRLGvdjF//TCS4XucdRMNuLAcsMzbp/hbPGuOW3Uz+xvUSb+pMyGuny9+pemvnJ
tWwx1lbokYJjS3RYI7jTOgqyBxc/IPvNixuBo0xA6neBcbTvWS61jF57hiU6vS6DGNBgBECMWNyF
1adX3wZyi4Jg37Yg9mpasCQ2e7YvnVBTYAx9Y55M8uw/lxmHDume5KwEZBGGa9zWXgU9RaB5cAgR
19aCV4j/qnqgEaUQSpl7jU+GWR9HP+e15KP27wgN7P9R2+Fi5sS7q0INlbmt7a2B7lwrTUuG3h/e
OFJwfByxsqxfZY+XdFsPsB+8Pf9MhjZhyOJlZAFbSCwAid4EwMxmjIsjgnk+SRb8lslBt8wgunhE
gD6yE4pzQIwZR9wg11Wt2V25ZcLj4PB44hnTj3PBXk0ktvrGNSIbN1fndphpvaLgtcv+gJVQ/iTk
+a/CafYdAmNSKZRSJfYMeNCPLMm0GAlYhxqFR95S0ADYeTP1LxybtUQ6BpdZZ+BuurUOHu/yPvOL
yj5MtuSO+K9ezAFrDQydNnSc+M+auGClhUItmbwWhyYIUvz7KGVRyrhvbghykPvuiRbYQoS78AcG
ed60j4ZnCaMg/7lPnKYqD1fVZDxnd1tVZxz3Y9n51nFXFvF4jTIOp8EcUBpF+fEsDqkMYfeIiCnN
80t7ql/k/cGwsC/F7Fia72c9q2DHMRbbIt3veb6EhRPaY7q58HjAZtRstuox2GJFiah8OJ1GJ0H4
HgWflEepo7S1++LAiyPgGvAbVEnDlFIAeWLxrtvxE4dseq+0CSmwrf6aEWbIrtGDOh9VsA7iBD99
plTsTujxJpkjZxGFl2Qou/2MsydLQozHjsbz07D4gKb69FyQd27cGjAFiFEPIRoprGliAUxipi+z
8Msj0/eRaQ1iTVWQZElIT+4xUwOtrYpcbCd3B24209LDai2lQ8yms5Yeq5DIxnXGo75mhoz8mqY7
8DiJJNLETXyDVc6goONvj6HsDzZ/UZfgYxrdQfvwmiqsZKdRt1DE2YZXF4KI0A+afaJFr/GoKuot
hWw4fPL/CjpigGd+zJg2z1VNH6WDmmWHOHpQoPhpdMh7JhvsbCNgErUTQhLLIU+H8wlMBb0RbQ3M
Ma865WMqJtiJgTkHmfE15bM0ckhTN8WdSFi7cqguD/q/EyD/my0yAMrAwoSOAlak7n71WthZHjXw
21LgTCwyeo90QX4a0SDMo+JFmgFSxkaex+KY3+BN5pv1iwZC9eCFDjbAzmclrRvAI/5xEaAHyy1Q
9SxVBNkTNqg1JkZA2sEyrnqFNKsvyJA90dw5+yh1VqpWGp53lbNspGpiEG19p10h9/5KjJUDYN5N
hfmHSQSEboEphj48jQd7HUGaTBcE0vw35Se45UfB8QH3l/D9HvF+3hDwRCzqYIpbI+kWYWXRkeZD
EDYRZCEVZQomVq4plIQyAkZZEV5Vw+9xI3CYNb46ir2yNOTGFC/nBqfFDkzquv/XZR9064Lt7rbU
Cdc68oKcTzz6VXJp5ewBXE/+o9F06i6eDsHkqSqbvYc64TNZ7+YCPJVbz6IFwqY6nrZ9ruopQ88b
SkNOvGpMWFmYhrU3Q4YLoj+d3KjAgwVHngZvX9QvuxxcpDuEk0dFiZ38qERsqwztA1rtnTVrVfr7
3dus+hSI2zsYTu4PT/UF2dG187tyPoQpK1w3BD5mzQIwL4WvnqINBbQ/x0dDiwAzqfdemafT10o6
fAHQLnbkVaP/2pz3CQFE/lncgbBUTrnZiBMlQxzWeqSogjDYwP51Vo4nmbknV8xOnE7w2AJVVEXh
MB4LlheQwnat+i05zoKY6KA1RG+hm2zz37kxTVYK9aeyuZUsrWyWbNUo2sLJPaoifjurh9e0FiEQ
uvisnykGGGOJVTKOTXryQk/dbjsMOAPGSSNm2qqj798Yv+QM/Yk55v7mydcaXP9Hh2mJXNKODW7+
6qzzLTyXaOkwwhPqz7sqzKKzzZj9FVDo/2C70X1OsMUzU1g0KuvMJ5ReVRs8t4MY8tgXrl4zfbuq
2BRCcerTN6DRAy9c4Zd+FpcHdDegR5QyRC/gnqmypMqFQVOYCouGm77AGA+kTBiUgu4EympMddgc
C/beUfSJazNq9keSNfpwEfIbv3K6T2yZKoyQlpunFkgDtuh9IkMStjRK5EEURLfKNiDnotm/cAwh
SHRqcJ/I6mA8qymBI2pEXy5csqqWw1FGKZ2/Sbg5PoN3+XPeM2r9A04Uy7ByVvZy6KnePXhzmjYo
BI5RY1cs5Jt6PGoKFkqxDTfqeQkY/ZOWEZ13uTFjE+yblPaA9/qL00kRekPkc+1APV9u/K0gAlXd
eiaJvDldtZ4W36H3cBzsxSdZ9X5nZz4n4SgflVbYLHpS3EKzRueh5BMEoJewm1/awVAtWbLX2mgO
q50rnxwOPvKwc+vIYuxsoeb1lx2KRV69SpXX+pTnkigjC1tZ2Y4m231CUNs/vrt0iFv+lG7/J7kC
MuKSjnAzBvfLgLrJyJjPA80xpGXdafBdzrIBEwwHWpZZVkcKCjuWpZ1uPha/OaI65F5vku5FqNCv
erRgnxA7G8nAc0hN1sIwXxBHvmIN5+hr3t1rLRn//IKq0tdL7EixIxsyaKOg3X8PPU+AKv/iuz27
a5iuU4vbaIezY3E/usPgwrW3RA+GP7m8iqCHEkxnAcCM37PRgiVMmoTkbt2z2xllqRl3xVjgVYVk
rNkeQidkerGwwpSl+HQVmECKueqbmFfjA9cCmegdo6Y2vHjiAvCAf3Jw1ZwiXDdodoOe/aZPbn0s
P73TemNRk6A7L3XWe5g6E7VNkDmzMqyPBqxb6Eo+pjeDnFNfH7T9G1tvpiSjMIUV+0mBuTESBLtd
9KxKMgTqP1AqHU+op7765zWNHXfvOhPSXngtXdyEyjzKN2KD7aOwo7SuqIKprtd7S3QDBJzVK3gm
fmcQ8VA0Y+Fh5oce6AbNZliwluu4V9aaqsHAOlDd5AC3uuNq+fXsPx5BxY5NsC8S6+yVEGI3ciA/
datnnBiD/U4l1ggv6c6tKOD+fZyhtCqrvPlBU4Y+riHCR1S2nKaqjcOEQvv4QKyTnnwh9/q9+ywU
Jw4MDLvdKc1Lk8sx0kXs0taDGnTTIvJndC3K//ON0+pqSZc3yQmaKLp08a7B3OyLYxkTC3OtD1N0
Ccxx20V0kUOn/gt6vjLhyIwYyp/kAlb3D/Hm9f3116NOyIRWmuDlY9G0ivE1JGR7A3G7u1DLdXT/
JvCQB1G5fkqpHAk/D8nHRLTaKzzggqOImYLnIoxi2WkS+DFeBwI8UzBvk/zMgX6bn+acnSaIyg6x
p9UZPIYON1z3POriWEPIXbgZFKGlms0jc4N/ToVOBbq+MSjk8NF6nl4yJzvOOICLyLOhqdPqRiRS
uTFJTLwyKfwtkqXLCDVT8EbHGqs6fOXFz7rAw5WYyAVvRWqpKd3vPAFu/SC/IeNPIlVjO3FApfTn
eF04vxYXOnJ+GlezJCeQIRYXa1R4h4JCC79QNwgf68Nil1fS1n/f7Uf+UQmH5ydYc0dnMcGjzR2E
XxhE2GMLvaxN4YHEj6EJDIO6ZJITY2WTYZ2YbmgX484a6y9fPkNSmiUxJSjYa9vAcVPEf+d4wQ26
BlghalrXTsgM064i8ki+oBdzfMs3zF2ivDxD/0rdACB7OSczujsFp1kuDE0KrJW4sU1fsSpieQUl
kjHLd90vmEdxwwlumyHkB8CJ1m7a9MWno9i4VFwG8lbipaKaI67paHFWzKiMtmmEV/TOyqdIj5rv
AGB/fXgiKA/kSGbHY9E6NvTug7/49ucrrLJcFu15nqQsY8Uf125J8u2YaA/QTpkTQVUFFnEMDSBV
1hiAXABAL3md2qrOSYusaH+q2KSOo/x3gDo3xfCUZc1TPyzvr+I0V/oADla3T18mvnldfXchNHUv
fYGgJQ7jn/TN8wURCZCnHwB72qYlVaFiYaLZp8FJynLt2Qfg/6dU9WIDR+qlk+2gVnR5BkgrZRwA
tjM7QpTpcI4kja5VKWBLZ4+TbyNMiAV7ESj5Croi/J0ApAKp/49BSpzfCxFhzmyEdKoofONtTAiF
TEIv85T7u9anmNqnt0oteAPg2JrzZweOoaveGbHTiXL6UUAFlARSLFqxV2H3l0MbLCeQmaJZ6zgQ
vu/U9eVJMCbr4c/WzNxowybXTAdnXgi7LupstFikt0blEfj1Sz2ckkHXS60n/asZ/ohKnZTxnWU7
lA2NwuWO3C3sJisfEftlNqInd0mKLsX9y3DgUt6DIx+bS5oeStC0j/+gD5oOSfKELd1sYb9QTXl8
gJfBvSYzjUwZiSeXQVWJK7Ru30tOD+NP5LDRYnScDv2zimtne2edwpn62cFByBAjvnoRx6Vns6BQ
NtypR9P2s7CglhpeRRqB3B23TD7yC1/+VX+erYDGy8xFAjsDeat9EYhfn2t9JB8s9imJRjOuRVq5
2Uq2TCSt0I5O/CJA6CcR35Y009AoZUzIxAqSnxujfmL47FWGWN0PlzE6jiPT6ecxnDDWgE5OGpKY
JeRjwKMYvjgiVGuGomLzFMsPvAqFK+JUv1DQdvB7ThfQxEfTBmTSTKPzq1EHah9v79FqVbinZCRV
22jaUNfpUOzwSq4ttv5OnfYwyd/MLI+wRRm3zK368xtGn83wOvnW1yHc2kP7926QK3cKZC6xhCFE
S/jOx8XHeagYXpE7FOw3qu7qvaWpODCHMLF2gKsIGLQ0Jsm7JSqtpu/EOl8loxKsGEkC9yEVKQdr
+RcJ3MB3osKSvgI4ojMk/0Eho8yGx2W9hYNnvNH/8FwtaQapFFRIkIVRzRctED19VgAxjI3gIYu7
eEP0o3aFzNUnx591JH+vEcuEFW5Nj0GjsI21XVoiYMLmB85YOQb+AIfNqqHbx+UItITYbiMMuHR5
3uQwfZtzfFur7N8BzbsJxzNHgyezKszgu/6AnzeDhB6/AsqdOYXfGYDBcpKsaoba28aX2vUtltR7
8OZWTcoMOX9HQch1oeJb4IPv60tU6q5FMHhQkS2UuzFnuYOPgJ7FaDuhF9J1NSy6MmDMk7/nUGRX
mpHwGz3Rh4v9FIbBEawyoZzDHb6nhuSNNIOo2uWia2bdm+JzJHVtkCdOEMAdk69U9rTIRltFAawq
5ur2v0OBxr6ipGjEDbyHHy3qzdekRRmIe/dzCd6dwK2xr8S3ZJMZFrjfa+ZxOkBq36CF4ugOgoCt
GGfqX6FJsYwAZrQUFRTiE4sPr+z5fQlEMHH9mx7kE61s7hI4PsERzRLhRrISUtxExNULMasiqft4
1Ekd6/EFit8zjatl92eqwjJvZ3GoXFKeWTAwFzz1inCbBWJ+Nuy8+qyz0qOOHID2zRC7C/goY6zp
14Ch7HnYSKBCpnuxdJMMRjU0qXHE75LtnR4Y4XtDjRAWneqVCC0VGNfzD2btBo0h8j54CwEhjruQ
CLiwf0UGF0RO8sV8t9fBFfb2LwFXugQmSKRiQdsrLJ3IDW/5QI4+MYDW388BzRTWk3ieYyYtb6NE
T2TvxYjC97PuWARV/ljeaNXDegFiPViTy5ny/3BfCsJ7QP+wiEBQ6hMGWHHK2E3nGgnbpgwIpsmq
TsKgTt7kKbblA0PhG9DMZYIFYQm1XuQLlOWnj3xCmYqGU+4J3jg35zQfgQ9exe8rS/n4GrBuVowQ
4HIoSCfEfG7eS3OemcDxo5P2dQZyeVkQjrQAchn66hnhLeSDH0cjIX7uLpplYnY8t/8mFZuClI2u
7N6xbN92BHzWQp9+RlSYa3bcX0qHASwEtE3Jh/H30qH4kbDGLzsxi1Yv/kdF8dUpXjyj3NG9ZzFW
eUX087UKtndOjd7qniNdh4q9NDnkVrgl6QJm1jGBbHuqYtdNeJLEvfZtbud9t3osexdd1p7yDXqP
/aGkI0N/1ckUs52ykPkISn5qmS+VoHxGGnwYzdPsjw9nArrQVZLdpDK3EDSyxEM+CD74RaSOTBYs
/MBvxSUs3D/IQLnBZpDRchCqOQv1iyYUf/JmiwFhocxcGAlnpRJW8R6ult9dsno27bc5X4V5umPJ
4WMfeWPqLF638lrAKgjMCH/SjnY0X3hXBChQUBnC90nHSl5Kf2ubkhuTEbRs3MUFE5N/RM/tJ26g
dDLJBzTE1AOeyqbDnUg07OaEdtDAkf9TcnrnQ1Hv79ipnaGKz+abTJJvEw6QIeqFuwfia+ULzGGz
V1wl77SFZsQANzhIdntwYeNj3H03KjLymxt3vTrC1zh2+UrfDVCN7AGf1MY/P6oLk23D6QOzTC22
zNW1oM3zXWEjtqRrtw3RqYmoalISjZC3Kodc7Jl1Obpd8KwX4lHETnZdGGrYR/pk2TqCdFxE4j/8
1Lw3InIW/CQ8o839uaBTkJ8Rx+RK12cAoRz8R+s9hseJB28DHKUtl/OufEhcuNNsviUvgLTrUW59
2sORqumSH6NA47rWO0n/wgHj9SfvwBJkgOLshPbTc9dwmP4hmp+7Nb7sfGb+ZTNmRYEplKoWqR5q
P5XhLjTzUgqj177s/kPiHilVb5Omw+RKYyN06vRPPCulAATgVj4KqRZJjXsEH/6uhOyVf3BhYDaP
LbGjEjFnaZQ+jF5qmuAM9s6JwXk/0zGoWkhmkKQejJf4+x6rr5u2pytaZ15FTg4BOgrXasC8J4hq
Ak7GTFZO9MFMbkbwwxp0ZnLHsnMnAqdS6aG8Cv/s93sPU1p8Ms12hcP7ykkAlKB9BDzifmEaIuTu
PgGW60Qk9zVcwwrFYO9Tv9pXWqaZR5pBMAUL5Vu7WlHz1774SwBcJOZsu2T7Qi64FGzgS0N3VOYW
jMpVm3libG3xD14ppT8P47EmyXsg4ICFs3LcBIxwy3FbneWgah+20YQ1V9VhyRkl8BtzJUTfgOkP
uU9gKEy/Vo/SVLmIdcGvd47jiyuhuaXQ7h92UaTQ2ztyTSAGhTM62IznjJqIepwYk9b+hHB9DaxU
cWUJkALG0DASxlKQldoG8G+WruhBmSa9UCVr3H1q8mHU13gsYMoBj6co6+yNzxB7psQdaiacLIA8
HFQDa7Lui4+9m/kEkRX3xTrWeeEVxVO7ck96cqCRsyIMbC92/m6O6rrP0ktz0eNZTbHP0Wb66APF
EFLvHW2kACE7Qbz9tOAF/HHRCcs0qKhW5/+7/BuksDuZV8uYM9axafMcbKQzC3Yj3JSbjOKVVhVa
j77rI90nKBjDBM3C709UxTprFn/SSu1LyVwXAF4fXclpJrVKQfmksRca10VB5YDUzIyx2rv3LVdM
UDHeWe8l9zBJQ47wFXmlUymanjIv8sa7C8lpyEeffVlVWCyYcgtu2mDdp/WgtgTwwvlGVSvdynJ/
eZf1QyGNojSqnNRirDCEPrbwdASrmD/lJ70i3EmidHcNLgiqLU8j+jqjRn/9ejrRIW73PT5MbPNC
YSPX/3lCaj52nzxkWFM7b8FVknDffx9966kr0907fKY5cIlcDy0xm+Kv4GkE+HZn/4aScLP9bA/p
0xX7Kf+xI5a4IrD/8kVgz3Xupkxh7loWKLLY2hM/nx2qKpD0GiNdd4aliHVvYv2H9JBFJJVx6xyc
1dXpxL1603NuUvoiC90b4kEnN9V8Mt8uOIwMOfRqyvZJwy/PbUGGuf3eMkwIKglrbt1JecGnRQSb
hZI+dOwtjem7UpjqHywu3iILbiavgQErj/2EU7hBuMfYkbvFPvsH6P2Q+rrM28e5lY2IK+mNjlyU
DM7awKXsoy3xAr6Sai93Fg11u4TfHLx+Khsn2489RAtL+5oAe/Cx7dZ0qX/xjG7tc4ni/RDeVjne
kYARNblz6auAvIVblrxjMkz3g6K68zapjNv42NsZMVrCm+AFY6+cqR4bnxSWJ/6B+32iHrgqGIRc
i5d9YEt1hTglBAzXwesj4+B9ufyvVuS27Ezite0DWMPJxzsi7eK4kxR+TQROHQpJ3RJTHViaNSG7
WXlo5q3jN5KHbbJOnQqr0G5uDQur6Dt2HgCgaKHn+BESxOqQ/XrBkvddFH86Pzg1DF0Nt30tCM56
0Q8L/Nz2BhO+ope2K8Woxw3fXg7d03I6Si6s1WPE55DcQJYzX0Ib/FhmMo1JSfEZAXBo2ASHbv1w
FdkRpIvmcUH1XXX/COwRoDr/QE8L+DSPB5CFKXmIevVoNR1I9vMzrrrvQvvPVSB1yCGbbTDZyx8Z
R3A4unw5yoBJx2950hJmB1lRGpViNA1uoEbdeIIp3TvXIlhNOKbRbWwNxoiwIB7y64dVkr0FK3kY
bmdQZ2bwg7YXtxvOSdZI4HbKEuGAWfddA+gyRboekDYyJy28kS/J7EYGwrQ/kHKQ00wzgk1xa+PB
OUjtfDs3HqcM0R1qNSLb0vDj9WkWWL2+EPBQHG2RBwvr1RonjfUvIDg9cpmKhD9ND0inRym9rhCq
5pGs2HUIwmmgqIlzaRWjZ82UAIgNv1+nGGRVzz5lRDBoEZmpCeOutAiP0LCXuygAhFv3EQIChUPf
ooYNG1L0T5Rf93rK38hYrqYhfiPLaHim4nU69mYrRNSV9RSU0a9RF5Bq96yGN4/DZoMdHY7Ef1PG
apFtwY4YDSCNr43k5sQ4VihF0tH9u2g1FOQfWW1du3LlD7r2PVRTYWgT5d1QXW+CWbq26Z5wq38S
/VO4SceHu5mvuUq2ciPoo5fOjI3dnwkxj8QgYOCu6osBu6VLawB3Bhi4KhwNwGdD83FkfaMkKpKW
5KTtz0OF/fJXMWfkqx0z4h2Xn4CKbCI/8F8wQXfBsga4+lNXRK6amQP0vgBEC0xa1e4rhJ+25wL4
tao03j1rSP8TXRMQdnIfKo/b06woYRoJQsDZeBV/ej66PW8IopjUIeTIk5NgiMsAK3P7uhC+4aik
MhoKTPUFlyCz1oZK94tm7ERR9WMV8+c7r0l4b4tHy3WG7ODg/dU2Yabf7heWS6Kkq9bwkeGKj/Po
3bYi8HgoVjQ9UQQ46wxrFs56PiFlig2P1kHZvWUySFoyYg3zvLgx5AUrg0AhRz+ZhDSG/h3RrILJ
2mNTWIQe0rX66BBC3N3c1ovBL+Q2gGW5L4YHb1ifhEAhj5gLdp47TYNoZtNEu+jMKtywuWhdeNO1
HZ6p1omLIr9uA14jPh9Bmc9+c03ZH98BXmMDVZSdZt1il1bvi6lJhS4sjqACCCm69PMpebfaUgMq
PeeeizGhBRVBr8P+mxunzWXDFegz2GUuemnUKseVrLiAFsuzXWWmQzXl33kRiM9j//fb/vhbIXEO
+SkKk8kvbQ4KArGlb/kdyi1m5nf+GDG2kJq/fJh/PfoCEOtRH1j4K/llKo+F6VbnxgDAxVNaImku
V868ew91nR77Kb6KzNXAKBRVHqyzSc6sRWrtRgoU4oAguKCsrPZMSu63BO6R8ii/G6FQi0znOyDE
tbaRRSqreHFZVbjkQPwSR6iy9AmzlcidYtjmvE1R4rbA74DJG62hnioPSGk1EI21APG6/qwRdYH/
cevIsRHz3efw6mIPInDjCubQYLOiZhhct/899DalzKK7IS5fR3Df4AAWAB3IVz6AhlItoe7s2DyU
7KScXywv9MVn/ZECdku+Qbiq13klB8VUJr2+onbPKz1pRcpyubba4NaHE63zI3j2+KpQTWq6y/se
qWEdWli8XY15ixuAhq00ByFD9m8wwStZJRmCz0sHgyDmRi16X1VB/ZDy/qcdxFiRwGvzaIzLOPyx
2zkRaacB00Epm0p+iGxhU1MiDW3nhQ5tOOzYOxyfntDzAlVyF0O3YfdyrbUOQ4B8BMYnGwXB10Vp
dPXuEMU6LqDGe3jF4OJnp2m4ie3tw9+BvEWMDynyx9jDlu0/h6T81a/x15DVWijSOaZEuJMqwNsn
TgKY+nIs+PI/waaRCc2CnZ9EMyn2kft6M2He6a5rWgD4xzKyCPdseMe0zgvSR1LTrIzBU/eHko0n
hJN8wgxK10XnIS76t967SO2VRypKUPeTsbyRVn4u0EZnh38MInUqQykia3iAEW3rb1/oyldXyWFr
O5qu2hKST5TmCoX36s8gEufdHoElHww0B940+mIz14269bt7y759Et0voAPcBhXCIv/+uHGf3lq7
azGesJFNcP+0DTlFHqgXGo8HI+ezuaZUEhTXkCP8o8f7J6FvtYInN+rwVvY3HfY3lN5XRCYHTzC5
3A5fKebLhTSUC2dvhIY/TgaA8LsfNr5gw+4lHqIJontbMUzg9r48RUJwvP7kF/lj+vfxZiMZoZdc
2oMniDGY+Q4OQiHT3f08GWdVWaJ3EdoWsoHGhglh0ek3Waw7F3njKSPVvPjaOx1MxCiTvdLsKBd4
E7WDuJfkqlivkr60gbQHy9EtYAwRbWCL9sR1vGWoFkaLLdR3WgDgcjZcuB8/yUzKpBSDIeSJbbQw
zDSWXBQWxBZ+rX14A/SvdsTPc4DWFAPxdMH4KNrtP5jcRIMPc4BSkBG/ddHv4RHFm/NLHuVe/j4n
zejZQElCPGECGQqxStI+MefoWFHsneAtJMKBXHtDPN9mtzDd7X9jWmz5k8VQbDmoCmyrO5aO7sxZ
zHEiPrKZUTM1e24HZTmovULHQpDYmW010w0O3CkE54G277mniLSs0fo47uVXNnWOsAM/ywidLqEf
xziFXYfAxqDxmICYbvPLt/GF7Kubs3UpeAh8hzos3mRSPPA/eWJzt8DVx4r6j9zMygs5ovNO/eLw
Gt/0VEy5FILqZnBreZogJEL8P7okZmedXcDZjvn+u6978hEAt1GyHVBg4psP/p/OsIfYA1So5a6N
biXD0ltOKXc2MOF3gwhPR9RDS+YUTPhhj+uRsmSibEDm8ygP+ldSDRV4URPJC+//p7mSAUtJ4rzi
iXYCCuVVd5MEv5CtrbBfw8+t19W1GYnPBDQO3gtB6YzOvaOSwMJsSDCY0Mhs5/6/tq4PiQJapCMq
15vBtig8eAubCBlbGclDLdHMFX5kCc2ksFvsIrV4XP9qYNg1EshypcBppJvg9qhpFu2oVtgBOXka
OSVvUExff+AHAnPeLYIPi/MheGTG7xtSRXluhdHYT5c5ACj8tri5Fdxu468JI0XqUmKsmtkrIMZQ
pVcS2B/TV52Vmsm+EWML78gs9WSJrm5Zl97Z9NcrnO+MM+BXFZhnR3q9lIvphtiP9MHPXWzcnWGv
bMWe2x6PcW4bcL8C0d13I2As54Wivgy29S/cRScbOT+D2hSadpe4aYNm2F1jofXZoBqli7V+/rKX
HH93Rsf9c4Ch8Q/vHRwZ9H54C6j/ohOP8opjQK+oIyavEJUJFpbdQbLM8nb8jDhg45IYMLJ7e0Qa
jtdtlkqFXPw6CjK73KFfdceRiXJ0/wP/blT9Y27rd9uqMU0dEmL8GaqQZO+/9QfRC8+cQEvi+ie2
opWIt7Hz48N7tkB5ZeJ3HCPEu4yk3pV/ua2jp40bEigM9LsjhqPISoncqEQTGrGideIbmMwiUsp4
lLbQZmOV0Q06N+GxUamvUDGB7ESTbHPaZ4hfqf4zSh4bhqYRPIfaP9AmcVjRjRnqxVVzu+DKfWPz
K4rE0aBHY2DDn1kjJ1kdSQxHEcZpJ8bqdvIsRybFjh1u0aGPK7diF8M6mK+07YigLy5FjzhMWPb8
9Y/QPmc3yc9q6t2ml/+Di6KUTgVxui9ZelVcicLv4jMeKUqDI4L8DGHa7f5t8nHls/qHtjRJP8c2
UznsGdwiRriDJzI1HU5fusmfHDaKLiFSSzGgt3tn3Ez5DJmHfsvdVa05Hh1tnppQ+WQc/zyK5Vf5
+gK0au8JEVb+fAr7G3VMrLJTNrMesqTIhC3u8NtEYq9aGG22fMWz/fzJ3MVg8udTopzECcTbwja5
48HSX85Rf3WDL0XremwOR/qvTEU5de3Wmp6nPrD3p4Oug5/IAqSiw/uoAwcgVGxZ9XoBg7fDL6Tm
Y190PrNrY1pu2LANZ54WejAKVC85MPpfSjneY5POtnz7yqW2Lgffr/qCz5pDk64F5r50Xwk/ieXV
zBDOECWUCU8mQeJF4rCoZ35fVnBJa+D+Q+kRsukcJvc3T9kqFwzJPlabs+xWp7okp7CMg/oOuC6q
1LVC6EsN/ptUruRNnQYH1j0FAzcE4508jc5rsBxuL+CTtRNNDrevri2j1XCzna04bgEszWJ22Shi
FIbiOjC3MMDRBgMIoNjITFW6Nyonxe08CWUFYWMn+VtBkEdxVJVPHukSS+XjewUr97PT7p/ruCwq
tlHt+L211mAyxVuxL2Ca96u0WsPvGiPGlXqLq2+Z7H/THawpk5MDTRyxY6su0/039CNktzdSKEQt
18TDOunmTTGU+6L17LnkjfJGFTW8QHRHZjdCkk3z0th70OELa8KzuA9suRW6naLj7WykYHQNRPxE
lmAkXpOvT46RUId63HxTR55SNcnVXY3NUocUiSYAy7Z/VMHqeY5UJNHKIBvlP14LGRfvM75/jRNd
C5wG+WmUPjv/Te0qkMbbBfP6Sng83/71T3ZVdqyf0k2qQHj6WW0jyGOU03nAKg1rIxruApcq6MXI
et4p+4ILs1OcjuU8SGppe1jF/15vhXTEhJiz3JdrzPcPA9fE7+M5HNLW2trUJjlAuSy648MQNDmW
La8UNor/h95PS/22VcnD/MeiORjfDp6pgdppo48+B50I2rhq1JISQj/5UXAoa7F1YvNDywDKHNPG
XhcasaK3jBbDbrMiAgBxJ9MPchExvGtSuIQ6/T9qeLugwLicRMKbw6rS3TsmMtOWQFHJfcNKzUm8
ohY2rqe6qjWBVmRQ6WNQHw70PX7bjjwJUUyfldN9fTAfcHxqxRZ2CIn15GfRhKNXR8EVxFBh+Rsa
4SkRkpU8givb+LHybldBaBpstvqDM8wMWjRqXtxCjBA2VHPGaZ6XI8zq0FXUK8nzSYkamTUprVjT
YgGEwCxn6T0vFBQJJ9FwrLqIsx1itJKdBh65uuT/z3XE+BEvrih2wh/fFw/BNuGUdRVhWabnvYZ+
qKxGCsvnqq8cvA88AYt+OJKo/Vqa2Hq31UOCOp6I/dAmXb5Fivpid1cAnH0ivcZ12vYUPS5BgSJU
Zj94yYKD81fD0MD5lDRlrYHn+BS53uAh3JVUHD985WtXb87xc7b5JBwC2DgJKfodTLUaUnf5cPU3
2BQiDryVcHYd6nZFVZvBnI+pkIWXfr57ODl5zQtJtL8h2Ne3FO+jKXQeXXaBsXOzt1r1eorUpq1F
GZgvWooY41qiNjq2oMGeINoLnMMlQZwkzAAwWnDluFLemb3MyJsUzXjveZl8V3b8k1bQ5yJvL6Br
uhSG2Eg7Ph8i9cS6hQUgwadiRmcUxtum63sEJZXYxcMOkC9F39/fzeX+P7cZHI4CaCESBCrpZzxl
jIDtXwMONUq84iF4SgUNNF9pYCyp9B/LssTnSu2BYaoXHiF+TaXuqborcWqk0Wj4CxyuTV2pbLNb
zcpbvWABafKtxIyzjADJGRaSob0rTtQka1iWlG66VHe4aLcnHn+Ay+VlvX28SUkHdFfo/8Wj2rYO
efZkaHHdAeExZ/20XKZflnHPu0oHe8PLX/coM1MSkVUEJ0N0euijm1N08xPWzeJ1RhncXoKmGqKy
mIABQBngIxCgbcUBbohUwIJhyDiRaEU4skButBVX673GopzYB7I4tBFpAevMKVcas0mb7AqYrIv7
hl+G2fdDaWWehWp6Bu9T0KV/gaDRyduKXrdU2Zcl7AHvaIzavYnT68qHkSgW1IMFM/EorKoadPP7
BLxkx9KqNvUKLXA4m2MAcpaOupCaCBHrSG+b+Hq5kOjGgRNhI1PS3loJjUnK2i/isr9HfE2al+5A
B22yeo6pT1WMW4eAOqCCVMoqSGS4Q/cCWBTUYUbNZtsaE88SK91x1GABzYu+idopR8JqUIyo6Ph/
D4XAMONFVBH4mWs3AXm5TRqgb5JUiLt/NnFeRoRNiNbR1J7X5ZfDTF41zzEnEItNIyfzxBdvMxoT
j8M5+nj0uvX3uXbwZNkqdoUK8GxYqNDkzmeS/G2tvrhbDCxmBhWS0ILhoe/NRlIJbc6QgqPP3vpC
1iSzjsUQDeOOI9pAJq4jHYGclk33rnNPHK7OCY5SzafdhRFzAd3qT4+5Q3xE7zqCp9o4E7mwiZH9
ZnzuN7eqtyxMphCXZ3gh5SyGCmew5IJhv3BJCCDvvtqPIP4BNAywvF/QCetpal8fJ1ocWTSG6DBR
SIyD16QlVlQdGUXKtrrzRrdjTB9pqm3uwvmEL85S0kLS+30O6dKKH8ROxMsZ6Dg5/TM0cx6q7TO3
G3ABit2/YPg5AMXE9v0mmpqNFOHY5pQ68rMtnZux//Kp8eDmbWvH3XADm51zGN4dSVCJZC3xx5LD
nEuey0KttVBKwB4thla5I8tV2Dr8juryiuqI9UX+IJ2Z2WYTGCm5ctZNhsqVe2hl2aEz9TmqJTqj
Bxaqj09Yq5hDcQGvCOgHtAFuSrb1snm+EEQhTbSHboS2z3hSmwYrKA1VHEMhh67PF6n5YdIL/wBV
UFJv8COxR+wd6el5CvXrrin5p5NLE0zQlKUdzQLlwIp5SRho3/mDwYa3M2hGCrmpHoRIi61HHlkH
DjeIWMusJw/23TuAWQLvIPpkkkP3/XxxXqJJpfIVp55SbVUhyjoItmXejF0UeQ9uh8lSVAHKoJzb
U1+Ia2EjzIeVDTjuLwJIJjXeM4kRDWHO6eCGzcKniOnog0vtUV90zCZUcDHmVM3y2MFkzBkI8cqb
8WWtDYgORD/ajirSucGuxSKShLuSG7q80NAvneYsH67ilbS0tBhJltG9MhJAY9i44M8QVrdMczKN
FiOU5PMrutgfnRud2Nyy02dctR+eFDv96ghgX4XObWLw0JfikCIr4HFGiMBuhN1C+Xmwl8koSKv1
uZR6fSodQyVEWStg8GxePXNkAmRv/OvBpKKXNDNf+DUabo+dmHkocL/nPR6JgsChKcd4pWzAdTLm
F/lO0/GonKLtGsKVAcLGmgHxiq3djlyrO+/U0ZqEBRGSf5cNhiaoh7BFMGunScYUgrWKjPRFUoB+
eJ4ltdDwI/ZE3ouAV5I/QF9u44Yl4cDZa6b/zCPQ2CpltIIBEMt+XtaQBJkC6/Oi3YtmI8K2rCen
h4WqA25QteeKxMNVmHHiMc1N1SaWgC9t67PcV+dyP9NbNYAhpZaw97jgxZYM/1Bn+8ig1q06+3H/
LaKtVL3Xwd4964nne3Ia73mwZ16vQ9P0ZCcjqnvQ7bsrp0KmVDH7neGseIO2q+KtfbankQkci3F2
9AM2s4CR3gYlqaU3nvkTCAqoCky1Ed+EjFNGzqhkEdddDd8XJdc26EU0765lLzpepyuBMG8ipCDf
BnD/MV/HAhpa6EehhA/+x9JE5HlGwh5fEcGGEr7lNRnzeigWqi8MhSigmFhh99ypSOgAq+CzuEuw
3SjkxvCamYzXC3i6gb2HduDfudVicHJbfszTeAjIIYAG4GvcDtlUuGqTt6v051jNZpihms3CUoML
ax82a23ro8Dg00li1YLKx1rQrzpwqsSd5z0qqNiSUYz1iBVRF5qgVFN3yFYQcqELYUdgA9WVwD+g
B7rqP6IWCJxbdP5pABsE5OkYRr2BHeOffmKi45cJdBnSj+xVnHEz/wR6QIQ7bhitTo4fe9MjVpJG
KGNc917WhgYK35Vo0TX1a8mw/tFBnHYAM4oqf1EH3vXnKAb7s4wV3uaV8i4MRL5lmZrFFkfWaziM
sGcltYvx2/7iNDMZ2QkNEr+XHY4hsOaXdg79giMvkDXfnTSKcqE498+nWBLs7+x2477OnbFuBbI8
LsxjZC6NLMDFBubpwBtHdloFlwwE8HgTzNvHg+GRLTlC/mPXRcHE3ycB/Z4g62NtzEkodvfZtlVU
5rVdl9Uos2tVMqvKn2PYoJGfr4joJOKbNtvjuUigOo+BpnW1qhEW99hl33HlpQ4ljGavi9B5+66m
XeX9TwG/Br7z7KuJhosniiWb3DxoRzLvM5dfky6eaAta/0ijVgq5jg2v/H5QIHzvmwJl7vn8Qj0z
7y/YcYJnzW+doFXAb06Z8PnTgadOuv/tbkE4bgGtXV+M/KxK4xvopvSmIp62YRUAAJ3068raN5El
wkXqVVQQXpscNvYpgz4lbLdZi03cnYiCciDR9CLy5fXlJwlPMuzPpM0zs6BkFw3LY9Gwv7l8nCgb
vxnrNBAkWW3bCGYh8R9iKgESZwU0dtX/1+o/QadDut4EfUx8VUJRVMLu4HSKIlvR6iuwdcNw0KYE
otxyl67tQXG1IHc/drZyxtQrHZx89lL0ywK+p1bXYFPetg/2/ysMbkkbLGDgksSTgWfZIuDlRuaJ
TmFDoANAV0VbbbdhgjUJfr+xvEanJ5BgwMylM5yUELOMZZV7gwJ7muldhQx1M5EvQLF3NtHCh329
nKE8kXtz/468GzU777OYvpu6n6Y3XxwUMVzX6vdY5OzUAdV1osI50YpFE8OVWUKOox09Xpxk4gHs
BW0yD+xdTzjRWxwCTWdmzdwHjVCegO9gGxDho64ZQumO6gZpMwdtd4MViVW98UUI9QU7ca1199g5
WBSYN0SLf7L0uJzL6QEkKcHm+N+D+3Ybu0Qg0qHSlvUtaG9y601uC0bku/7i4vs7EdhKxH1j4CqO
P4ki7TIqjq827u6ghArJp8KZPyARs8QqPqYSXp+UlRqnrmhJNW3PKOX2An5YZCt9qqp+xmpTbgs+
S8e1JsOpAlPmIjmjdRweGjr01GumWTg25vWzc8zD3U5QDu+S8Uhfj/pMl74YrN5ZFBFNX4hn3eTJ
B3p13SvDwZ3c/41+4JKsSOVy/QugYRKyLRHxgcQkNTsPN/uF3I3JLzehy8u3dAZ7z2Wulh+W+8X0
R2exrOvsOX9QuCLzbDNoMXO8i3W7qhiprGH7VP0VrU3LG7WrId4Ngo+esSi9Yq8w2KS5MFWZoO6A
MStHVTMnman11LcjD84gLDYqM/5XIuRUvPOZbqKkm7BmIdGojTpTH7yM4MqlnyzmnVApvlLl1WEt
XuVfvO9ZuDXcvcT4ZvoMkr/tZm+glYpubb5HX7oyyTZa9/3Tpl0xymvgcIDE38cCgDpUoijAQgTq
FflqbrQQvxSDVAQOxqqb2fnhV1ZpIdUM4YihOVXz2+1NSfIYAoEy25GVsOYLPNpXIdOdBluhbGB8
3qWiBtNzrZ3thMerVVdZCGkosI6nGQPenU+wiUIkVL+MDG+3QU+LDxGiD1S41DNbWpJhEkcB13mu
LmObxPr9bbNPqgDA5eVWC4nXkTdFH95BgocPRv8P53ObhRjp9bcjs7AQstvxdgFqUx0uhxc+HXvc
g1xuumvNsv8BLYmxkICBxfgSMNlm/iV/esIWZF1bQhrxPNRW40w/V+D8+qUDCM6ORM1z4Hp7qufN
dBcRIdC4pT83m9Q/Wmls7v63EL47i+K+OOJW6rtv+IvgAfhu1TG6g8qSVxe+E0ztCQmM99MyipK9
hYOfl4s6W/epN13YZGj79Z7fQNKN+0U8lM3KrP7qFA3PJLq/5vNcYgi5VT9sZ9mwJmrgdVAiQ+54
h43Hr2HLuYn3ZqDQbOiRhcMJ52iBShmdNkg/0BBXgim12B9XU8refjSJecW/FwQ3PD5uYEqgILEP
XrXuSESK+hVBEZDjiVHu27TDRG6qfjPep8eCXRJIN5A5Wh/5UokbZgizhz7NVqBShVYE3XxRFkEB
Oj0hwAuxD7LtEx/GIuL0WBLasa9B31O5kvdxcupBV7vGqG+dKR7Yk2NlfkoFV2tv1g3K2D/hFIXY
7NdP4ilnGsr5q/fkE5DyKP8aLk55e9OmUFmnnTZm7gx9b8L3xzFBZK0WqfF070Bu9sTfWkRCMyxF
HglOC37QAy7wffNACNstnH80xTHzGJ8kgBjj72FayBGKvRPk74DFbItpmLOBkuy+J8+MPkg4TJL+
F2Mt97dapqgIN3fdVElecXI+XxapZfxGy11obliXsCswl+KHm5/USpnVxFDZR4J2AQHJv+3sm6e1
zcicr2/WQ43rDxrQmRJ3AZrqFE/q0cCqA6TYGBil6WBrMqbhUY+2xWee0IuWCFO8EceE9hlmgjWU
oJxdzJtONmcgnJWiNqeeWqFzVbdvn0tTOhkizGg82rOVLl5JUb35OMdN1zhnQ50nV0h/842PitWu
/rm/mkmUoQ7DQ65ZOuNtLNRZHu6ajFpzSnRLFvbti6inuBilkiVWvuCTjKz5Mb9wftAqAwPBAQKD
9TI2GOHKXxjTkInkBZyaRwCEFgXHVY2O0U/rU/iMFlqYirQ7OvetqD1pwNhBq6NVnXlAiu7g1LSi
tqPyFYkMW2HyULiS37jFcg2J+jKfGYhBDKDUhNiKur1pgylUGt5n8sYqcWsmFx9g9YNC50pniDyD
pjUYaAI4FT4pVpliGdav+46EraL5M4RxWTqI1jHLMi8cyRWR0+8tBXPjb4ttzL7qQKpKksGAIiFQ
sj/3Eyq/VnJWZ4aLsDLJqP8SuXoaGWVcfy5y8+g/0cWLQoc21ShvWogrMoyECIX7GsrLWdrExuH9
LVUR1gBKZTdDDKuuwcCcHg4V3Q+5KFKvFbQRdm0br/9qyM3tZABpy22RgAdp3dfq9jSTnx1m1x/l
IaOk5QaBlIJUKXWYr8oCe4sR3E3lZA8TGJzjLb7dRwDXLEQK4DssjiZE+bTd+QYxlbGekX8Opl0X
ZDK9D1+3/oFoTRQn4wBdie0mxChu9cIeDUl+b43OaCJhkT0Tl/EvKOZhL2TDURD6kXrZpFRWvX//
GX+DHhQLgqxiLWGVl8qZHgHUeizT9hfQVTikCed/7TnNRZjtFlXyjd4iGHJuHV1m8lwGsu9npLrB
DtF0CjL50/Ar9FKFd7/6lHtCgCe50AaXh0qFeE06uHcbUuU7A+znwZJvSh6kjVYQad1mJKCmuG3d
htYoQd+d3hBIksjtQGOsKdA1niV3bI4UXdgclTyB1GIL7cu0kjlCVKgrLLx8VFaiZhQAXoMNrpt1
uXUUTjGJyKz/bz1RE/Z5o2Dlwb8VeabX9QZbQh4D45V5uzuStcNWJg5BXy1Pf/bkVxr2xM8tVDUn
tdmiVl1MxsGlzNMUgbpVz3lgnXkpDm0yvzq6ZizUnwS2IPgt7d/9MqyrJ9xz1AdPQTnTGBEOxBWt
JCrLAsL0zXszaJceH5QDYHC3VFPDiPmtIG/XFr6siFRtV25kMlnhoRcs8J5n17Y3FACl9sUtT1Qd
HqX8gUfrtoqh0mPOUl1GvxMRnYF5ijsWS3tn/OJ/LE23pLSe0BuSFTFpVaCXc0qBaKV1gVihsHKr
aSCBvE/G3bF4ukytbYHJNnnUK9yZo0JVLDmbG8jqF01TK55YGeeSsOqro1svmXw3mvPULAMxaRLk
//js+yr7it7qdVY98zB37kdpd/5A7UHGmwau/H2RNYHd2e7uqf8myRphcCYnkiPWevLsT3osipzx
zWsuHg59sySNXA8IYmWVm/9cNTVWQaOv7PyjYfWiqV5K5jh5djrlrMBtOkdqPC2AybaqejGkLNUr
VekLZd8AC8dih72+XmGH1Aj5Ov1hLSBOrihUJuuCiwXDlGsYhuoA5LXY3qqKEAy+4ypKxEBqdqyY
FJT3G6H8ceij08WNQ90t7YcdFkvkkLCWN16IPWUYyBVR/IPNuFKcFZ7SAJcyqKbUC7aAwp5182na
hRheHVNiniTc9P8yD4CSuHPqYWPwz9SKduzGFOAIysIhfs4P1KKOW4gkRjZPDu3swcCss48rpg1w
3NEYOe/MaCC9x5mkIWLyOl0c9ROG3VX+dtQ0HOtn8eszG84vx4mW+NVjE5W8RlHW6eaPQCti4FmM
H9gZ9zDHaYkzLL0UPIMLApix56mKNzKIGBg47BzvznC/MHQiJ4SmwYuWdVScVWcEIotsX2yAQKjE
IHqC4wiMWwdmWnJBSeic0hc5hJG6z5XcdenCZWZ/FfB4U9qzFWk6nmvErwKYQFxuWhcuUHlyvEMk
neI7k1fMUugYQolZZ6VyVL8zJEcbUZHxdo5D2h41isuMQjqIMnrseXKAhKxx07Q+G/lftoeqOpSd
Xs0LyU4hjid6jKB+5YzTbeZeJ9n9mf4AJOAtYhVYy7tUqS58jL9p3Zw7KFqKKJLmmlDaIJwh1BKM
LUDym7mmGO5EHJ7/FFFV+RPcgevGJCSFTHDql+yxQOOlQ4pDWolXkgrENPbB+Q/JRkAwsDLsyzC4
WTSuxZSxLct8PDSptcIPozkcriu5ttU4EcX00WUyBRxRL3v7yqezGYBjOyWLP7HAN2cGnMCMhTUS
3d0gJd83U1BfkIu0SzRdUnyUprFVykzShtduEu/w/BSGyUh7zajuJUfm+T7BIsj9ERX+ZvPQk67O
BVXIu1iQ9cr9KBpL4rxvS0YS+fUtHlFQaYd89ZG5JeY5lWdKu/OB9aAUV3i8V0mPWw0Gz1pM+JGe
4UbrQj2Pdzt8+u5mjpBGLLO+AkZjqqzpmwD+m7RG6ZaO/0Rr8CGLrbJ/T7ZkCkDIXXz802T4gPzm
tSZ/lfnSXMzF+YZVHU9qC6x5yEAm8+8lKXgcHVScQARfNTffWryzQZZItAcP7d0rrB4fTFUPr8Ol
m0+YPJac+uAc6Z4ylbuD1Id3vZJ2sRGzFOFtDcCTWYYBKBqVi4pK0FpabP/xvmKRf/gBKWqbv1fg
lFgAbugoAfim4J3lmPHp8q2yDVStnCC46kfAPOVzTK/1x+yksa57V6KecUwBzTaHmavadUXuIfsM
DGk3pQmV/uI0v6L3Uixps1oqlFHLLg+Ct7yWVhVbUz7NmNIHZcJ5r+PBL3S9zKI+KSNzqB+X4maq
QyNMu9K3+Cz2ghiondwHs39SZgGoeeEe6IOsdUUNh27t6k4qcxNJdM72Q9h+6OHZCQqEJwc9nVra
Rtqqf5VW9fx+I1cSiBTgld0sL7C3kuRHYoBP85b1KbVefjcWEExYXTiSnN3HXvUIe/JbHcxibVXI
tbTs1BhWFE94UD/5tpbu8YxW+esPlpIbl9+M83Brq+hd5Kggl6eBIPWsuIhz5QggOBL1YsteOTwS
KK7ro51Ua1xpwxRF6UFr9Bk3xxyDjwGslwfmvKX5epCenA+Z9QB2y6+p7Oq9MpaRdZii9mMmXDLA
S0Rb28r6Bjiyq+LNiMeLH2OdTfl4qoeZYhjVUnHKJ8dAbdyg23XhA6/XqQpCf8hSjvRYzU10glnK
SmgxrbN7/sqzj1OjgPe1Qhl/eOMFzxdybUHUamT2Q/4DZ66vSzfzt69zj++67lEWWJFatuu9AcXo
OK6w3lcBmpLc9FKWwEjVFyKzUiJeMPf9FtGnLjjepxyRYiujE15x7K4pS6YegL2znzWx+snEnJn5
s+vROA682FDuK+W/fGGev0Ayv48IshNwZzNKRoPRX5zyUu7R5dHYmvOUVuuaAR2MHnGdD+q1xu+G
vcnIlPvWnczz9kGxC93zyJwBh5Jj7T/nXuurbHIyOVh5o4CyxgP444Pwqq43DzwHfBDlssJXSo5J
ZZvdCpESnxJVHKE8l/MfNrXUuAq6jdxzGsIyR9lQQPk9FxmGx0KT136Eh0JO0w5GbStkJM5FUenY
V42Zo3YNX23UvSH+Z3rY3XdKZkfThliD7zIECcqh9F8w3iVwyKAr43gwId27fDvn8/UcSXWQnWaC
LBqK1L6D8R0qGPTGTSOD2fUH+wfL0V+b1gdy0cNzzy6WIqZbPxkrDR0LhrI3c+cNZFDWOqe2HXGr
m7c0ctEfxnXp/3j4v2fbrIgm+DSUMZD1G2ow9OLy1NILTfXBBYPMld+4PnRFQbkv1zUG8un3d5PQ
Ot/NHcMiZr9w0SIKb49FSbtk88PDMoZ49sNWOks5T0jrDHxzs1eEQQ8EBc6dYKGVdwsWiaoTtkzM
Fo9IZ+tZ7bEniYiBlmoYUseObAoHT4P0ib1C998lNnKn22ZnL9KPUGan2dV+l7+1zZrQgjXak2nB
O1mWBx2xkfFsZkvlH/XsfyF695TrvHbGKT905sFUbkItdUcNx3IUOAVGYqr34u54dLP6xDFK/cpN
CTaGWqP2G3ZgcokZbPbpm+wuuNCUlvgrGT1ymb4zq3aY9TlomT3fQNsGWiwKGvEIorLNyGm0GA7z
yYrnIH9UBjg1DhbtrdkXUqYGiYW5j3py+9g2roRhSsJ723jIsnA/TDwh66VsCoZ0jR27CILnZHb7
OOkAsXZCI5TI2U34rx3I+nrP7KKNLJrZz7v9HHC0Y8ozUq2rzjQTUOGNhToE/1ss56kSr9NwlVRF
Oi7m/OJ9m96OWcygzhD4VWC3uVTO8XYB3UtMpq09VH0qrW8gJMW4Uv+9/D32grfqN0kxQAE6YGSt
BIs02GIwyPLBX7d9xYJ3zsrQHX9iRfE+EKYdE1izifpBK87hFzCcfwPxghHFZvc8kSOxisCJ09IL
ml8CScbB6pz+C5aTxrjT/JNfDUWT493AiDfTq+CKHR/KvQPM43eeNb5WFiSsJrcyS7dh6JEzPiKk
fu1lJ01ZYkBI5KBsWFcA6hg+9vZWpdLe7u9QBIeIElA5JLW6WPd3RpUwdWbMHLruR4p7YuPCUKXs
pjfR9G4lCyIllOiXfWvq1/biLzUQG+u4K5PrrT00AVZ9URAQLU9FfUx7JgrD0+iwVgvem8N8V526
+l0kesDZmtY30KyxAMYXFr0ESThYbXbhNEZXoyqQ/C/ogqf8M/xbsqdXXV14CEg5hGmT3aJ/nArg
F8YXnDDX56Am1Of9r+SXzXfZydxjnrKP60Z7RDCm6B0pQANeGPcMbR+PXWypadLGdJURED/s+rtj
00EF1N5UUSJEBfp9iMBT1w0HSZ8qOijnGSUeX3Z0DQA3AxUnlJdGjsQuA2teFollQdBizmq9agHK
n+rHrg8ljondRcptFrpOKseKoZ+IIMGrZ/x+cXmnzK7RSnHpLiwXE7AlZAzWExZvaHVYVKoouyLK
O97e5qGa129EZa17DBV/2YfwWhbwrzLeZ9s7NfhhjzhJKPXOv4t+iLIDRpc4i4NV+fmuYw6eRLoN
IL1tBTrbs8UVDAp8ro8TJzLOCTUVppJGmL/2DaFq0jjBqmlC54laVsUBznf4jmSgl9nUr4t0DE6K
lc21GWyTePwQvojQUyNkzlfBEzFk2NJWqK/1KMhV6e3heffU2wPGks5BBg95EGmYP9G4s2qEXTqR
WKLnXrxpQE/bfax/xzJLZOaLaE6H8Muy9coZNe2t37kyLnT+A5O5UeNz1WGeQcmEJojUJeZmu4Qm
YmZVCqAsmIY29Caa+z6k0SZkvshIR/c3tFsHc96Jqe4SlafkHGn71KZZ1puhKCJKSfrRESSAMAQU
rDl6M8W4HQyc30HcV1PUHdEzG0hlK1bm+4XEoE34/zF5glKQsqYBbMdv6ljuLiAK/5u67YS6+jKq
FLfX6KCtzc4tJjrjUJzLQBiIPXx7l3PST6CW79yZix29ZQL/B560Mt+/wUo5n6Y+0FkN5iYjwnE+
kquUeIskRcsrxK+FJlFuZSwsLaO7BveOt/PofK7P9C/tlYAGI/z/mCfWgfGdCmWzhVtELCfskcJN
rVgqF7wFsiQEqxYDSJFhE328Id456CqKaF0LjeXrZUt4vkhu0/meROLW/szNkqKpn6RTgUF3hveU
6e7dPTMdWQxNJ20RCWW07rDf/8H2HriFspknJsqplrX7Kgn7bz7Ub02ON93GQa8SbNTDEmgr/1/i
6iqFmNWWnoDlvnt+ms699MPyv4+OBJ5ThfA+fAdrXILpEjji9yvZZfZYr1RlFHXNpK2lQ+f1M3hd
NdiEY5ANpy9qGjiD4fZGICba6cR3jjDI6nnbprNWKnrCXZNVzcSG89NThm8YRc+HAZDeFgzeO3Tk
7ldjcVGAkXfHMEJMtaLxq4B6fnEbaTO+n/3WZq04hxFCzQWXXu8Q2t/wduT1HWjsOa4PCpte+aGE
M1O4kygiv/28WOfob/WdqzCueqxe9uyxJj+yUCE3ZxaV6YophKlX/38JnQPS2G14uk+NKVSkjTkf
bSvixB2HmiN6hhCitr30tKhW8uD05kvpCbhqZ4EJburbKUpnQf3kBInlyYnK1nvHspfEH5wmg33p
0x6QXewN8TCgybElnRGd2M7H9I8nDD22IPYm0SmRcHSaUI0U+b871fCJNPLuuaTrBGU/GQneHom/
9JUUY5DJKfn9un9AybHhh02vg+3mYIgFHPMheeizGFd6ojns4NTiw/CsRF6JZ/0Ys3AonLNolRkL
JgRH813OWefK8ezRuLmgMJwhgE6+1+vexu4+gdyOlkbLzTOdmSkE44NUmlZrqCvBDGW30gj6jtX8
Tr23Bj8HamK4jyLQKLEZjqoyLvcA43ToPSbTprLGiW4QNgLwsXfaLRKvbUiKgcSLN6okIUe0bBmb
69veh0yFaF8j8wJoNL7ZohtAiWfUJU+Vu7k8CO9DLDcxz8A+DkIrqIxRBhHS32R+SIoqb6fKKr4c
GpqjjvE8ZAN+lRE1nM4FJoB2+n/OL0ogGnBW6ozH/RiiWOB/sOnapRTGdLpwjamno3xMCZdc3N3o
mccqSLe73A2OgDz0NdRZUnPuvpsgAzNJ0WV3UfOdosDysdEYBl41NRy+f8J/Q52LvmpwLYkTgU+x
aZE6bAGWXhjO6Ceyu6cHNDVS8JLbfe7FUCn5Oy5bhNNFeSIExBX2044o5uFv1uR6V1BwLS4b8aNh
FHEqbhkV2M00Iw+NstUL7XhLAjL+ymYjUDEBsws59k8URQKMbYJBIzPnqTsit9KlrTGbUrXQGko9
7uszjx731d1RyUSLY/k5h3xi204jHrBeXjE40tNOp1+pGvnAZPKjLgR90pzHIpVf30h3M9b5mnFc
g+Jt/3J0x6CCfdLem0zCvW/diqGx/eCUiU1vLHe0U65uHUnugT3y5N+zGj3NhrVIW4cdSjSCiwqu
QVFEt52WgwBYUVzhHbP0aviAEcale5D6362GljJ2OJ0PtIbBj92NkuhyKzMouonMNfqEkaNMu6cO
OAonQYZlF2lhQSJXN/XOCldeejmYFYM8r0VNaUs1JTP5MTsAiO+YRe+FFIYbA0jhSHbSm2wfD10Y
PXJT1WDpZ/mwLAg7+SwQMPulHKiau4RziRG4PaT6ysG/UeYAwaJiC+hIm0HC8KbN8Mtlb/maJsv0
XoHthSbzz7pHsSGlGEa9OVKKeh0mnu8ofAyXLY97XTgMhcUaaPWeDZ90xLEFuaAsdmQ91Akr3zpk
ZhKOgtfT2vC7Fb2s04GTZYSKsmuSBojFA5O26cVK2GBOxg3s5R/QYpLN/sQr/He2ZDBN7zyTlr+y
9cC6ASdwoOajNmgqt+gv1yaN3anBr9WXPWSVTppQcUEKYVKp1kymco3p1Q6oXteeOZS07cIsZwXB
QdgMpw34VZF+nBWFDw66a55QninH3IkmkXp7nBjfGDx0LxRECOOrNY/ld1xdiYUbSiXimZINcjtr
kXrbmwnfCBRmQQMzrBekXMM4NQ79rvTExmWVovsP9JP/jap0Ptxmcnzdqc2Kz0x3m3SkeAT6SEug
zmZaX9GkpzGJ6i2PvvYpTY52prYb1ajuHDHOhA7SnAjW+PgMtlIiXPppccqDshDb44v+P+u+0rGD
AAdRA56GTvvJIzXjHcc7hNwk6hf12Mn7qZRJeQXH46srX4yCS+hQvLmFbPFwCYcIo5PzMnYN+FSV
pOI8n5LwmXlf1GzJ5KuXpQTsK+J+nAC9GgtHH/RLjvMqp4nY6BNaEPU/ink4hkSEmJXL8GzEkUkE
+x585MnFXIeKEu0F/PYkAdd6EBlX4wxGiSqUxZACV+gM+iL4CVcnH+a2cvc6ARt0FhBRa+a878Al
Iymzto8+ZSCq1CRaOwcFyJPw4JCd3boZiFfQVZEzAmiiw0eabNchpR8avmb39pEPwZun6NdVjXP/
4BoIf28GM5MH1M+TctLpJAFIeJbCFF8d/kVClCQYJlR9kwFPsmb762T5MBV92wp2cEKKBaEk3H/Y
aF4Kj95HlZ72u17kzHCybAUzkh+NsXGMxJk1ocbhMGUGQwgTpwleUNPNaAP84OhBqe5jB1Uv8BeS
CjSxAPNIU5/GS7sUUVcL7DqxkVnnJex20y/m9TBpUYQrBb3xuh9NzSz6Oiu8pBtLzODqhbyv6dmp
ghPrbcyoecrJlGzTCdnc8nujvo6SJP+sFuEvW14sWEEjhTT2JQ0DQiHWe77Uwx11JFAObohqW0Tt
semGgT/4EV0rpYSKe6F4QJ3GCqm8PI2JsknfMpaus14Kju/76WGc0JEW1qwA0UzzOUeWwitzrNFP
dW8kERjPyefFTiKnJD/lMnaoFMUV0zqjD5l0Bh8+xDnHJ1Q+hjxo8i6HOjvHHjrTkRourWMDnL55
qce3/tsptg4FF7dowR26jcqRu0D/1n9JhOQZk4vU0vqhMvloCqAku9MP10EO+22Bz14ZFuNMxrSg
Or57J7dOwylYY7wLI0/SjHeC/RGDsPsaBX/y0qztTfmccTW4JJ/H0K6z+5nZ5HkaLYbK4aafnV1a
ClfTk1PFrp/DpUdcdaGiM3dBoVOBJ35YKNcbO3qbS7fP+rGhm1NGzzTsECpZvheh2HIY76mXNgJL
7Jp5iGRQfjwsCYJn5eQneZFtO57fGqedkbWFf/pNzqD0A7eBHJWuP42C5ZNviFp/b8URtBrImVa9
AONaR04IJkdfC+FiPvpnWG8n54OhH59CabZ5j10XfoiONnz4oYujy4NA25hPH9L+IPu41LOeM0lQ
gRvDaLsLmP/NXeTdhki6d/hsSrfV2gD+UOvWW2O6mCVW8KYxrpgcRnwu2X96QssCcyRlusMEeIRZ
Mi4nIBCCe4CaYNQtg74Qm4Cginsr+KM9H+fVkx1+/4ZdNwWrEkiiTFYv8u56J8s+3G1cdCc48Akr
UBTcqLZL6f4PtXC+fgA6hn3gIc1y6hfPxPxoqBE6DuTsMWIvMQv116+PyLBnb8fJpd3QlFJu5rwS
2m8b5po+rAOpCQp28OlQPXLZEle1p8Ue31XrKJ3J04K0F69/LXl5MnxR1B9f4hQD+jBmfOVKAfoZ
r7R1KaYU1iESDhvGMeDlKfuTYwT8QQ5oVroJb7SOGpLFYSU8wcCYeJR14ZWxKLIAa1nEg/qF30qL
JcZvWYWcHrwJME7kCcj19jkis6284xXaowyZuDrgQVHHdxhSPvQwsHf9Pdzg6j5ebP8ASey61GR5
Qxry8/4EdyQWDIyR424daBmBJg2izJBnumj8msTSJ+bTaX0k6d1bdMKPacUjSBP2jDHKGjmjaKC/
88IvNWz7zNgv8E9nGSMFkZDL259DkkplVav0Uxihjl1Reye9TwzjePQc7rxkIPcPlAmKHDACRpn9
Fq+l+usQ0AxcW+skhHe+cQI6BmQHI18YksItkjPN5aF8eRNKbX0TNfYfI0yFtW/HRIh7RysOWV2j
01iRVAs61gEnRudeKN8ALB7XagVFmXceFDt18dcmZd77JSpD6BZDykr9BP6kV/qzSqUKDvieUVQL
w6xz+yrAnjdfJ3HYqvzspIGZ38+451JWjM59m+oDTCmyQSnAdKuF5yKL3CWxn8behfOCROEU+rxM
FRJD3l/7FpB2C6VXUwC4bkq6UjLiBsJ5noO3O2qx4wg4gS3N5LMes1hPkOIMw68FoD+eCIcqsflI
q2zGtvORu6KlcqfbBoq/B+eZNgzl2dRiiODwqh2h6AukY10GlIPsC871uijfz0kvvJNs6iE96nYD
EgLX0Ge0nt5f5rISMsxTHiqFReqfzjLdxRRE6OaLJBVeaORZHG5kWopBULorJ1+pQh0vrOh6qmPL
lgRhWSYzzXBD4mnk1CHO0cBUw+xcHKX6Pi6O+WyUlFe38QEJbrTtlMYCqU5hoKx14ZWi36/ioDXW
hY8NaxS7iGAQ0nTQWUmMCeRNP5gnfLCJ57I/w7+IiJCUgLAGZSodVddJmZrCLO4oyUuW8mj0Tqlq
02pyMOLF4r/mk5qw2rBhh2m23ihGuM0fyDQVYBfLd4IFxsmoqIz/UTIcqU051ZO2hILO0KVj+I3P
UYzl9y1jmA/A3jI8oRhJWo5E4g7D9SoKArEEdHj+YT7yP3IBOlHBuxBs4O7wFqLl63/LKANIfWI7
0jS9aYrgKaauJxrtZ6cRZbsKvP4WHhuhdGQXNBoh1sqbC56O2QtuMyFWvJpPh6gOKSBNtAgnMHFr
pj2h244tWnc8fSaJFDQCh6jDxGdeALX7A0wo9B6/53CghjD93GuXC/fL/lGW5DbfmpJnMyG6cY79
hvoKrZeePtPcu4k14QQUQg+MzlDAaYgoWeD4WWx6a7n4OxtqROPAbzJ2tvZOs+YH+zmFMujmn4Am
w5CWbBzdyf3+zaX1CtqyNC1KNTwRnKHWxaSEpa6NR3DZGsdQd8X9LkudoDUq/AS1rpcu7q6RcaPv
Wb+2In5I+XAY5Afz4iOYZuTxtSePXExoCb4Cte10o5d7sYpng3yytEJhV2c1W6ecFrJJAjxRT6yZ
CJzBgrJfvP4zfayW1gizox6orD4h6WzHwm75HxINJ5YjnsifGvZfDHPLR1kOBMi2ZJ42rQiA26S8
D69VLA69HJZKY3IaTDXaU4IRii3WnTv2NPCGTWC4yEW+1C5SPgkNX0HdETTUPRY2Lp0/LQnLt1Mr
1oUqzZfKxxEry0s4XKDkU1RStb+U0Zi+MNDHmM1nH8XE9W9GBaQx6vpEtMMDinh+pnZKTttOOls3
VApF2ELkRlJH8I+oESX/3vAetwI9RsmYeSBCP78vdIdCywiPrqIrP5ydiojoYc3XH3yJBXA7l68S
cUzHE+o7XAfEOmPGwvudpSd7yuFqBfsep+1nCQeJQyeZZmo5QW7ZODoCogNYhu8bCxwSyeRi7yPW
dRZHnSD0DcryYS72CHLaM3GYwj+hDh5ohY9jkgsXOg3UbYke6Q5sZc22iyinVRoAB/H1qQMCC2Wk
C2g/qG/PanQxB+6WyhA5IxdhGRadU8L1CWWoQ09rQOJI5XgIRPvELZ4/akfcRxxMF0MgINd3c66J
RFxh6N3iRwE7MVTMcO4iQO+U5YvQuOQufn5CnsbBN/Bfh9NT1DJYmt2Y4n7O2Cq3rCg2x++h2crl
KPZ3uEATtkL8nC8OfMd7B+dq7Ae3xZ5DprJVttQKtXWfjFNtxsgpp22WjXTH1rGNw/ojs6xmSkbo
2Y4UqnkK6luTez86399yLDMGjC0fAV9OWbILqw62HN/WvxUHh08DnHuG4aiBOqS511ipoQ3oWdGo
Zr0PWbz1byZ0fEXzG5zkOjGEBREnUslqxFBWwIl0yw6LYwFu7k1jGVRyscCoLRyWcfDHgCJAohOB
2kjJwsripdgfPFid+S5HVHq/Iy5D0ueH+XdBUNH8hWibgaBr/hldO8x/ogJ4LN1Y6tZv51wBtaFH
qGKrkj+LSPXbdhBiFMV3UalltBCvMGFN6t+ReIxZVsCM1sJ87Kak5vyoLkwEmLMA5qrggx0kngfv
U1UV7ub/jfhZEpqY+6dUKDRdKjiEMJ2RaWBx+oC4TnA/Yt6DkH8HrgQ/jMyzLdqwGyBxc6zGXkWw
wu4V/MudTfYE9mlYp+q2VTyqgterjbDLyIuln3MUwZW/W3QjIY0Aj3+4aGUuNRb58NzIQE1VESTD
BFRLfyFrNM44pgoRkndN+IOQUWBiCnvs3tEABjgVo4KL/rx2aEUrlWhkge71guF5fqRtcsyxigCb
+iy08Bv2zwGWq/L58FS37Dz/WU9Pgo9RO2aDE0rVwkrH0dB8LXl4DzbZKn+JVGrz6jhtkH758GLa
J0VOoJGBxXQCyKxo6xFAA20UBg4vt4tueL6zGMD52yGlUEcS3f8U5oK1ICdd3sfvHvuYXwpEHsSG
yV6tzaQA48FPTYNU3fOe54qfcEf1pUoK93EsEutcf06TXRlWraDLp1JjuHCg15h1nHTEV2TAgFfk
F1HvMmC3yI64+qnyb8uRmpUK3lKk9xcvmPF2/O3L/NS7PzV91tQblF9Pk+CgJ8OKF+Cw52U85kKh
Sq2k2wP6fJUyNfomvOYtjbMNP4SGKJ/ruPZOOJDdg4djZNUprK2zRCSYikIVHH1FznpciP3Sbbmg
Nd2FV0htaA0jVf590hvi0aChNJboAPlkTrz3MFwgcoha4uwf1koEf8apFInPJCBm+P52BVsZJHOe
VvzjRcRme1WgXqjGVdpL92rbE9FZnoXDN9XEJL28V2QzphCZUFiDb4XDk3OdXpj9t3E3xF8Rcjnt
Qut/UJX5HJ166HaGkTHqqUMpDKi9DVnIymLUlmcj4F5TOaHhsWOdhgCJa0VBVUBTspWEmLzFcbc3
d7Mu7OoTOhZRJacAnPd/fXCxdroPyhbV/KMQkfc3/FdihJIM4wv3U/LK0Zo6ubM7AZEfXu/qlfFx
q3b6h9RgsvJ/vzjQ2WM/QPIjESyxmOydViwXYWB5jOTD/piP6/YJGy+9S/7exr2crawJuXgOJJFC
PxCoCKYNkDTXml1+it7y8LwnpXOfWdQL6MC81ZoZJhdrsY2Hc8fUcBAi9SYogDaQzPn5AQQhW5QB
psxJt9eStl57dQXH782DRFM69oAZ6fae6mbHdPUflYUjDNewY1M3ogNd13EQDDBWVcKY1iIQLo86
tdCdDIiaf6Y9CLLiA2ak8beW5uE6FGD7dLPa80GbHHV+prYrn/+iYrOnDSTaZTtBcStlmaBJK0Mg
SRZio6GJYwaPMn2VzDjQUYLrQ5m+JPQTvcVwHi+YexETpQRZadMIFv8fKI5N0RPmeKLmT0tCMW2M
osFhUW3/qU2EKrcVKoEYj5+XDTZp8pgSlObv9n40YKa2W/PK/zDC08UhfPh+ig16S5Mi9ugOoYnI
U3vwpeLmeI+A2kK2w/jw3+z0iYh1t6oP2plNLwe9rJBkvIaUrd71on5d+V+BEStccmWkdCZGo+fL
DM7a8HL1VvkJXIE4H7mZEvmLGmqy8sWmZkIOL0CZFX8Lyi+QZzxJRQRnQFW7COJsGWvu9jV+tLgI
0m0NgwPlpHY7ENJNI/OrO2bTF4EXiZiY5hcu3u8acSHmoPKnb/EA8waQotk+Fceb5lX15CSikIIM
LxyA06E7Ik88MBrbz9M65ugyjh46aw7xXwgxyQCTC21s7S3urcHTHDE0Yfj2460iqkt2NHIdKkgh
USf+XeNQxRmOzytK26Bih8db/EOYw2JKq94ikfvAgPOXvLTXFVM4gtar0/AxJEU6WpDVavpfQWsD
01MzbzKDuw/EiCMvdc5u1LkB0QfA76z3Nx0RAZwz4pFZ9vOumLhGGy6QdGk0zDV6N4F1ytn69vFr
IX8NNKAAAvOS1P1997WGifjz5xubk3Rx4dkXxpw+aoKjtA9XarZJcJltg+whM2888+MwfaDal/Ni
BubJWyxlPwZhl8Kg2UOdjgYAB14SGgL3SZGR8sICNwJfMUxfzfgykDWk9I46JfUPCkrYawl3LfPt
Cm50A3IqbHAFJvkprdpn8o2+RFvwZ/pTm4l+ka+4clh2txXYTezp9eb5Pt9V/gP7wm+qlbe6BXy8
pLz+DnBJEczpzOOpKtuQ4+rvznE7zvz2Z9xbEDnQPQ4kn4UD8BC/M7D4ZRzKRYscIeJM1ohnUZBF
pdH594Bt4IbKITZkmgbvzdmaCEmiMqGxdrW5JX0Q6Nz+TvB6PuTrmLiiKN70z6QHWkszOklwCYb/
bHGzWnrnuf90puv/Y3vYiYedmZn3gMmCklKsMNLfYwUYYTmk0L/kmUd7DQtkVlN7Ehf8wXPZPt5x
hLNfgfJ8+OWRW41jZzUOYxL23xaJWJrMIdhwAgXh1cs+iepfvax0jf4PYqrG3HE/rIs474sCS/MU
Zy/w8nqd3ck5ThELuy96O2JD/AIKy/mA66abFnHaFJH2JoTo2PTMZBB9Dl9LtR4wKrvuPsNOR5+a
fGHeBQ8Jvj1lGQoEAT/KtQJ8obgA4JO2IQL/tGwAbVJvTiRJyidOw2TPjpYpekQWLfjWwX8NH4qS
Oq3aK1vVMeF1W8O2f2vyrwtsjEloU2bVGuRQD1oNo19pN4epXVUIeir9YAvjaYvIDPMYvQDKmmxX
2sfXWatfJ0kejQqYdyZej1eRaXW/QX0nlvB8yijpvlEsCs+WnqvPxc5MFFA/XcSbQMFW6BAPxTkB
fioy9ufcpjTJfbWetwP/AWjKGTD9ObEbiRIMhpgbLUR1cbpAsj/sfdC8j1Avzn8/DIWQoRQ2KKvP
RwwdSBiYu3kj8CXXHnHwPmejZLCjYOD8dZLb6jEIU5e96vBkLz7Fu7N81mNLRiMeo8bB5lFNGMg0
e0DdKy5ffX5LAosSrtroU4QoeFKue7TOV/6zGVpIH8boLCwAPAKRdnFGIjHlVW6HXfjB3Y+zmz+6
wbSuMEMg0HxV2yWYaJhqyKvPQEjXzPXrf8mRcGvxtthWbfMy+0ujyDpMIEpQFRShVVoGfZb91uAz
HCk6Su/vgpJK94ao+1uqDFgJEQ3TrLp99woPe9wu2h/9MAg0Gem1o82SlSE994JlFNL3g08/87Gp
5m1GIenpdyffckxB1x05/6Uh05ElMUP6jdUlJuT8z3KSWO2iZIUjjiVtuNQv47O0LKyEPTCgXmiY
S160BuSRhZV6ZVG05Vtxh7kwUJ28dZO0fJ0hnps1LQAjHfPiAcgAobRRPQiDwTK53LtvctXmvSzI
n4VcR+/2wNKX9Mub3wftKkDewYQb4Z0qZpQ6CTqO9nf496GkZQ7w/sGcktjW1+j84GPFpQ/oTyRZ
ZLFMXP2McMP3QAi40PilFP4cU7oxpWGfAlLlJdTq7X6up8QJ6PLr8a6VVsMxMA1Cw8/kzqiSQ/lK
dt6z8r3/TvtPXDXkU4uHankew2Dn1o8DOJGCvLtaSTx/32EZ08VrPlF1fOfIodKVeXIP5CIYkK/M
KwMkLgHPSg5/i7HLWWFXzXMVcmbqwZH9YMLoUlH6aML8IKXqKaLWiFin6DpjyBF8PRqsTArm0FLk
o5JnG2ZX9zODHq+UV4oZzwPN+cfMlLaKjfaXeHv08yqIyu5fjD1lGBZFUjtifM9cmjPXmhBUkfiR
7Y7Obdwe3FF+ddliRN4ZLWv1GI+fIRyyH5BzZ/dcKu9x0uWjqnF5l6gsbZdIoSpI2h0DVcUiC7Kk
AnfabwXpJmyoPujWOVC21hR+Ix4OLd+WOizo6iVgHW0snZBiWihrNS42dGPFXgeRAF6nmMtdSTyp
kofkaf2a13S+EaEsxWjgSyt+ht/rmSiIswF5EogyhxQSFPnl3Lc7NDqFc/YbDYRu/O+UXqrDnI50
ujFreFS4DGyAUAA0+BfHaF+9Fl8rVuz2joBtEJIRqLRIeKryNDED5aPV/v7nnlOpZDk+7f9Zb6n0
3BW96cTNISJZA5vP21vNvCBd4ojmlhzSsOqfVe8A7HY98bCdFdQiUTLTU30ddgXA1i9PkXW5aooL
x4bSWCeSEHTwRoN0hI/pA2hPd4muKHva+IcaumzDgWHqRPNIPZM9KFSoqdQtFu0k694opGf6fJWi
OfzHnwDqqLHNXTISZSQ12cohLapvN3c0CK4TmQpv3xJ+PsGvtEtwl6p8gzXQfg9NGGbsTld00Ooa
ufkS5Wh4N5QOHirstFw4LC/+2iJQYHRn713eY9W3p5YP+WYCijK00m/YIPqWM8o5fY0R6mePwgnw
90ddxlUFgPmDe6NDaR77E9AQvKa/DMWZgrFTgiQtO4R9cVbOnpphbr+50aZbKYl0H6GAqdrf4Pg/
lnlmcX9M2JJN0cH7+FFddq3s4oT7Ivqi/vkUYyN4OFj8T1Yh9MKA5AZf9tXW6nEm7tCL6K7bZRqe
9UaKXtwZY0x1xNONdmOcfhMJ0rclcGodCeqrk7/WLjWBirAamm0GVOkKJowpd6JHdfSR/LWUUGjh
bW6Llzpdc6DeOdj4+aJyMS0J8YFIp7SvMIbNkw+Ywkw8FQ8EwJH5mo4eVTe0cC3Totx6jRJ3f1M4
xNqFx6FHYRXeSpORZS8bWuIKSPd2RLVZhk21Oy6npFI1XInL8+KzGdehRQlxtBbQHwkTL7vR+Jo1
vk0976gPz+9qBSme3erXwoNPNOxIvtqGp9EN50kgoOG8XA9FUEaBTievuo/Dw2a7fTq6LcikzRkn
sc/Nl2ySY+AmQXe9n1171KuGhdc02r/Y3OQRWZDNGB6ezEhzSL4U+4c5iGczUBHun9SrtIOkSW+8
vbENy+ja6zWJm7bqFaSgoPLNR2LGI90sEWbZtMmXr5/MhHBOZf5jEFnqa9EqhSK548iL4AO+uk71
djSCMAH1xF79iWepSw8y2avdRxWhl36FJHhNJLP49TNbxrDQAf8/qqqSFpIrmuo2O10FZbFENbMr
v4pYdqomTUw4T12Gev7nt+9sf22CXmzi4S7fKT3VV15i4aZHV6eYnRbCk2kPcYhPCam/L15jGgbQ
qHIYly7NP4/2pEHu1xABTpZRWbmr3XyFjYHZN+mrkAH+Yeowu2dE/B/QM1dN3b/aDxNcNygdCP3U
3/rH3GoRq9wt7h4QJAVKi06Zf95Xbad7GN34gmmiJWbw5/wdWRM4Xb+Boy0bq4kvme6mzzHqqGkw
qufAFrF8FkxlUCl7BV34ir8n1d575dEUlZm3EEfyaRHYG0pTnLl0P6xhLo7PZw67eEFc6RhBYDmv
328c0K+o0pEXc1Kx3o5rI01na64jOrqnRkYezd06/jmwlsV0x+lf/i0M07VHwKvR8TtwAGvEqSXP
iCccixSoswnGLnfBnF317BmWx0+Sv1GCpInFb4eM1t0KkUk3DCuLf7kFv5WtY2wpYXot4OP4G61P
Kun1JcX9iGOf6qRn6jMkXIONvYzYpZysITEdUdCkBWBk3t7ofq1Z1le1qgmYkBB+T5q4YcMPUgJ3
QJNjE26gQQAjlI8qX7UfMVjg1KAsqSi4xW4c1dc3TMTGNx9y5QsE7pCeNjQDxQHdiywm210a1KJQ
bbNU9HMPZwSpAb2Fs2SlHqRryCM8hNz8tKcD9NC9J3DAO3QRO55cIUmeTfi+iclUIwKFTFiz53u8
R3PSlAfE5dl7Vpxe1PYMeS3TKp+XE+k9b90sI/jmG8uEDWB1DDWJd5ZEPSRdGM2Xa0KNDb9XmI/+
E/khA9YPhZG07kZdg3Nh8hCfpv1F150p2xRnUUBSFXvsX2jHDDJ8XVtx676xy7N/OcK/UhA/4r68
z5atcODP/zFoOwojF0Hjze4zujawnxUDa+8qnOm82Ff7fqxfkdj1j5jXcLFhf9P1xLqBBX3DUXVn
Srixnbp3qIQYR474m8k6USBvzuLz6Ab6ZjnmYxEjMv4yprUg8iqo+sOCm1TSM+U935iXOJUwRy+g
yS0zse5gSv+s5R2gM5+2fEj8ZTUnLZy1LVDGx41aUUXRhDWurfLgBNoirQ81jz7SZj+MEdHspEt3
Js8HNyKdipiy59kum6gG5z9z+8WSGu57GQx6spX6tnSFKvXEQZ4+8I4Af308y0y9IA0t8VY21Knl
eT3pHPcTuDDmYZQS9fgljxxuaUooAL5uVbjP0vQDscpSbCcdzaYK1vO+O9I/MQeVYhnqPK1J9UjW
weHxerWjBmXmz4VHd+BN/eK0+treOB9HMbzAjMf+1NzH10YzDlz62nmVwrf3ExlEO6DEQPQZDpyq
ixRC8By4hXeT0QmA/VCCkKfwhbIhsz7ycH/EQkHLQJXusyZUMueVvT4JrmZZIvxuRr3ayZuH9wfl
6ajvBRkoNCVqAVqgVEUTsa0iREsM4GbW+2gKilQlbOV7PnVNTzELp+o/YJZaMIIeF5Q/Xk2hL9wl
MBrIr+Y4MkA++a5g4GvM2Qacr6b0wPfSApmmpg/VShMn4bjHQN1gi757L8Vbo3q3D0V2ygheaDXl
JtF96zhs7A18nFUyh8FKy4cBB2nRgP2aHvKkT3QeTJLRev3jb3xJxZQpSBENJARDbKIKgokX2Csp
IoKRhroAf1B83i7emVlXtV4d0MLoaU+Cs+hRGWFAml4NX+dB2hZ0rIghV2vexUcmVmaDMSod2qvC
ltKg8NnEQaLqQJpVUY+9NjHg/idTxLang8IOkrHN+aMeLVLVKCeui9vB1i3oMEVS0xndWWHG2U/V
4T8FiBUbip0tK3QWvsbUvVIdGO/v8/It0odO5feWaj+LMymQ7dLJwXpZXNb2RG8HlDbcpn5N4aHS
R5Xn9WhKNb7bpi58eiN+MQG2oFb6tYODPjc6Jvcnl3SuMe658QWDR3SZXnBO3QSj0SDYhqpoBMvE
f8D6t0WMMpHVh/a+fHEaXepQpiWpUgHeJrIGQVlp0Qm/9MLdBOTJEFAY5wlxxN4CofXCbsl9criV
0G71nJM77/Yh5PnLOyjuPzrfdHjxqQqozPIilGlN/AarnRtuQcFxVaSzwynsNVcOruNTjp9evvWY
3vFb2+3a1Gf+uEpRsIsVpDbTkB2NRyZ9iUXOHmNsvcQVUDSeh+XnsV4jI/XXwulAsONQr2ZX4beR
4Y+PuAffMlBWZA+8ompBtteXPJMXimKGdA4ohJmkxnVC4A8b6LLkx1Lz3mGKO38nwwx8SlJgeM34
lMSqZnhKBfcp7/M86buT0Z6H1jM/vHRlPzG2/8U9TtLQRqysFJyHQUdLOx/In0bRvF6DzJLtfZhj
zdkg5H1wvHMDsfSr+uEupRbCmM8fJqPeAidTVsRrAkWUO3hKu2X7g4wTgHxHEnXcQVo4MwW0AxzF
y2ph/TPvgzS46L/fSMgg6PbycCaiNHrQc/dKEQQROZibzUPEtyYwZZq+rj60rcRgmrt4bHMQeJQD
klDpgNBejcjBE8sc6Hz2fRauHtTWyx3KfYtq9H9cFKqqWRTO/NxHdf5cWB52ymc5ZIlOkCX5O2dg
Ipe6/pSDTBSmuRLiAYTZVuuMFM8mCPFbQbPUb+0Ox+yO/2N8hgCddHX+591ETq4gMAOhbphgK5WG
1QXB3aqfGdXFGHHqL7TuHdqiObNrsh3Ze2gleSE2jdziVrwMjfd20bFbWMHW99uuuSglkykyytXm
M8ZeL2hLy/vLUy1F2usv1mmc5LYtK8H3UMvfLqVTFjg93Y7c164DSs5DDRv8B6NqWBnIoRYdnlus
c4HWKGafIPD35HeOuvYc7hd8Hkl6klsG3723omqMdxYfuINUC1/ElUVQ8v8HIfywAWV7UC/SkfgD
RIgUzRcXc+1pTUNe4tAjekuLulWHvicTfKAId5qc+0m7VHvIE2p+DlPASsbnTuLKpRiEHnOQTY0p
pM8eEIPv6+bDiJjks8zy8w2W1nZfNry55JclsLQvvKx+8wo7ThL3oa/1E6CrHhvTPFDHC4N9PY9r
Mq2VZE1ibA1Itv8AEi4NHBrX7b3USacGrO9C1WlelsF5BWndR9vtXOLx6byHd53n2w27i9G8JuD3
CyuNd97HWaQfJvqNPMRhtWDfCM6jluZag3GXXKOBSVz5Y2D9N1KFd+vkgVSCssN+ELmaW1L9tKqp
aea2CNRkOAJbN45Wo83tz7PrhytbyGOdsag0nRNpQ6cplz9Vms986hQ6RGo2+PuEA6/q7ebz4CdW
HDW38pLK+BGJLz4jSD2hkK4Ma/pYc68ZO6RuGSeCiMxxQHtobOx5NrBfV3MxfcfhMlpGqAPtwE9i
uGi38F/P2g1eJYZZgICvfbsRf190wQbM8mrS7aLmnfshBF9eyti3Qa4OfY5PyakIOFbtGGJo0So4
lbx60UB3Egd/cSTTVmKzz7fyMWRaQee0eie3akV1gAIG/Na9mjtXU3BuHUc7dp/APcqkwx3beZKk
YBuM8sgsArjvvdvbD5dZNq6nbboPeJLpzEMhYd0w/vA5kEO3MqLN5nIV4FBs+Td6X0b7+U7aiaGv
o6OTW2AzeXwSt/52VLXuRdd2i2OhfPEn0zzzmgJcmWY/cYOnOF0EpXXOpF2Vf+MjEBXW5qS5PxIk
rsnAo6F/RI5nKnFikUTDSO7gvphSfgDPdogHG/c24ymxlOzO0AifgmAt9sTsoaJ5ZW581KNLQMGM
JUatk5y5s6hYVhS3v7Bketm66pWH74h3m+l5Qzqjo1VsAl0c+W4FkfQ2UGgGEKqsW8MCZomlixYc
oRApCdCM/HgEFMuiVebyLs5I74INVPjKwdaVvt0TtxmEDcl5PBueNg8wjccpxgoFlRiuH7pSEAUZ
k2sTcqFgBaEd6L63kNgihzc9j9/ruegzZFPnd+sOM+t4fe2Xm6ZQgvvI4kK+x+8XWxB3PWa5hu3q
7/YYdRrch53pfstWxDx+g1mP3dqbHuL9Vi3AqTKXJU3IaURQpeRmho4mtCBLU8OWYGRnlMRjDMsN
0D+PNziy6EkJy+bgJwzU3n69XLp+OHaJiTdOPYeE9n7DQZpgbogEqcZzWKZik1uv0e6TKRNk5zbU
8BcY/fpjnPA6MG86MWDdb9gGFqpXoU2XRWmH6waPOll+pd1v9UGZ7PYe+GNpTAeejI4zAXs9LJHB
gecz9ahHQ0L6+u+72rQzp0QIVYwMgK0/NNf+3d6LbXHXynPv5z3OZ3hXc0okkiLAcQy8GAZ0keiP
O/IfHOrFc47bJQ3ZreZ+cIXwhR+wLVLbGwUjkPV02MX7ns7TCjjlFo6vtiMX+/eDtwEVHVOd6tIu
Y9nuyu966dJQz89b2i6f7IfmywolAPqChuEJypsAB2glQJ8f4yr9U85LNdJGU6zR/eqGyXgl6cBk
wmvb7Vy9Gh8G7BhTJmiXxNdC8EJlB270DUCeQ7eBxMuhpLWQCYvhkmKFALS57ACZH42h0Ax2N5wu
uSOn06pIqge2tRiqKmk6tO22AULN6xbrbA2P9HtLDXUDq/sCXexyDsQU/uj0KqxohKHsWnjR+NV2
1+fiFz08YgpOAdi6f8ubfxz2r2CueuO0oRGDXPBpVgBPkgaGjT4aZiQX6oyeMravjUDp/9qj5pov
ff+MJGOvnhXt7fEUted/E5O7Z1nBpFFNdT3q+htyZ6Y/ZhZe+6Yq1sGEsbAhUh2wIoAhEwIZJjzN
oIGg9afctoRj6Go/wHEDIo1A9tawwR30eW7fecNrv8g4kQiCSjDCCHWzT66+WwWWYovyN0VZnq9U
lgPUnr7JcK5TptrbSl2hoiH3DGi320wiOpiKPp0Ig7Gzhg83QoVipSaccF64Wy8dWaf+J4S7RTvP
z9HaH+Q33KumUFtS+RZTQ9Lv58uF2Tf46htRCvbv2Thj87+a0P3RdLEyKEEqS03UGUhF1tVFteqE
BklcLQ25mQqHKCttS6VvLmUF7S4CLNB+XZ2MArRdOWhw0cp6+y+zyHIj4V/D/JnE/r7P3TkeCVKR
bynZsx37ksTbuL2PmtJm6S6ZV2DKRD5UCb1+ESO1zO5KbhhCMFh3/G23ITOg63osa/ms6SLGVQaz
gcAfErrglDXJCD+vS3FtbDcs1tkSRkjEo9cLrh41pq9Z4Tm0TCYEQNj544EJzyZdGw4aj9u3dr0M
jj0RSqxq3/DbI8lKUL/VFbn5zagIzISfMn9QqB9WUrfz4htjGll89CR8tFvrAbj4TZqhGNCIJpw7
Zj/9frcFAmF/XVrLqPZSM47rwAiQ+KsUW6ZAvaQ57WlDH5pjez/uOVqYU1yCe5M5dx2hm3m8kdNI
AsG4pJGECFySq7FmxiJNhtQEDg2HYTcbgs1rHOxnk8mY+6h69TB5jAJqLrCtfp7xHq0tyGqm+mhF
sv24cqBlN0xiOo1ynU+R67vTdIqa8OmKX4Ok37zMFe/js5DKASlsmuBZMj/kRtWKvnz4fhkjG5tS
ffszZtVo38+ZDNBkYuXmQKev7EUjCr23EZS3BNWWJUvgxi2R2JSlTy13gpwJA63QL7IOBUNDcEvy
qGW83YkGMgCvxqTyX4prfkcKT2XNy/grTWUJghHTOBD9Ygfm6XQ7gLJUhuG7y2OMLbKySwnx4PUX
W5aeDdV23jvJt5LTUNgmX35zKPDcUDvzwvfAIG6ghj8i4KkWc/CZrUEO8HxS5Nff6Q5nigC2D6Um
rLcFqseuICju5BP4aGLlwl+V7Z9SgKKPzGMwtI8ijs2rESXAAp4UyjdFP7IebHnpol6XrLNKebHQ
MXsQIigR5gEaLqnAUaC3KTfCal0fcuaot7QKyibn4MI4V9vthViQzWNQKz8MBp0yC24n7Xa5sm+B
1fl++X0NyeoWe1r31zLEefmQwwiHhE2Q8a0Qo4y1Em3bZk+nU9YfZvXK1fDpL7uqDIcX5sv/atHc
2GGuzBdzSUb2h7Oa0nM+uD/UYlzTY1k0lb4ONAhQ2YGekXuQ3HV+kjfWCR65dzZuB7s49zu1x/zr
1zFzcZZ4NAsLtUOohxt1foXpj9v885/WSbmN6tBrV7OeP7WNLmBygyqcEuf92tR//URphYy9oWk3
6E/FS3nN83qw+muijjLe3D/RuAcPxgosAEPUV1pTm+fBmlK6PVlyERfCaix4bDO9leU09dqK0OZ4
nDiVo+m4tbv+vGgwvjKuMjiJhOkE9ixy24jNG/WVuPdSHCmjlULnTUFU1lKV3q8OkFAlA7Ex/JeB
tG5PFGqeG2hpZ9CCSciXo8qPfB0DlDrWfaTCqo/7rQoZqnagRHD1QT1Le65yipas+AHAk0WWNub8
vSNoV7iJuhbkpGV25l3szlIZt/yZp6mQPxWCSQSrKB1uQ2nkayr6ZygJbissgAVHTEzgnGQMiFNE
wC0kDQoCAc90xUmO5vabIV9BxMBVvSPrgZ5D6+Y8qGuoZIK1NXu/7pdoGEpY6f4sxOy7lzup43vs
TspeSGU75aKGjl5Wxd7Me+e56aOhh3CgRCA6f47GXAy3bfspNERkk3m7s7ZfLpCUM8sY9RSpxds6
/rPQSL6X4BbwJXprMaJnHdgTBLXWJCPA4X+UGgv5U2zPMfTxwzpahiqVwBFnzyoD3QQxDMxqnMRw
v2xhXYwtiF0nDBIPUeAMppQy5LqS8P46aMfEnnVtCDRjpZCtKzjSQQuNmQf31uPSMOxN0S0OW29T
gp/76UrO6hMGunMEcioscsMyDdDJXvLi6j78K8puVWg7J+jqYHBaEpS1xC2WK2Xt+OZYDBbHFOST
XDMetiaymboEDrpQfzENL/h9KaCWujlIXNJcrkMcq/5FqFjFkRcCZzG3usvR6N2bWUbfQ4NbvWxB
CNwG/EjspbAXPeOy8thbHcy6pcbDpKnzMpYsOpVwjUMiz87pMWpj5Dsm6wglV486xTDqxHQlM+a6
aGLbQh0YutBy880+jEQUyQinmce7H8reHdfOQxY5W/Is6tfaDtZrqIzyvYAHN5tc/cD8DkmbCDLp
DiF8dJ4MUTc/Bgz8/CSusbo/++WdiUgMofObFJVB5QVOR1DK65GLV0mBGu52Ocdbh0EEbAyMhydm
T3EwdhHXubSY1gEJ/yRxR3esyJCwSJHSHDjvApYuRuwITyT6HUayNesEdW9J0yWFtGIIas/f/vlG
8RiiYzcH5Pn5C5+wOoU3Dqoid+NDG0JWKx8BncdJQ0vl4kHW9q6kyfeP9jn1cAvS7xXAeq5EXsSB
Ht42clvacKaIPsRVeJFKhUgsMNrJJ0FaQrrxlRhItHUWQ/aJohI0IZ5zyfT9CuxAYU2RYbPPYQX7
j6cfbrsXKgmoLYkgjXEcndqbDSyUhNkTXLz9glnE4t3tHAPZo/Q7Jp7mE/rfHVzQWiHTnYmaNh/E
jj7hac9RCk7fmC8doSzG3QaL52VpYvAYTTswVNVrb3HYcqJNCrenAKQNTmN4MpMTfm3wLAzDi6Cv
GsDYgoax7bTl779Gl7QJmASf/RSiBWHHBauD+wh1DBKur7FT0dumTLfoisIyRxg0M5xrbhaAGE8l
QuEC+zwoZVtB1mcadADr99oSqgD4fLC6wjvfSvumBMzYKQfOIZAFZ9yjtYG5sQuVxGwyV9LaJ/Rz
bqtd3Psfuw2thVxCGSTlnOHWfv0UohAP/oQo/Er+nV1rjwWwpS+kKyrifuqqid8hp0zhG22cPTSQ
ewDuhS82nW0guIbsndFni6MGsMVXyTXEfPOJ89ARu2iiVswCvG3yYF2Jr9u3rZy8221cd3SSSobv
rF2QZINkUWG4XvhjjCBM055vEqolAUB4xvmYYbuTibr+paaFK3qoNCfOYlpEuUXMUGmkSbcCDbqR
wrzyCrpibnfxuOINhLd5HV8nCi+X+Lw3NbWCFUKhLarJ59gZsjTEBBv55eqLEr+dzKqNNxoWkI6S
OSpt4MUGzB6pOLwnZGqH/Ch7v71ZUSmUA03kdj+4K+P6CFIAmQv6kBNJAer0qtNvBa/0/Q4sXUXa
1WhQKQHHHKkpw9X7fgKwS9ZQNH74Ysd7Z78+If1WzdNZedyQkoldPmQooPR8AEDxwwd1nN1voUdI
cNOFKhgP9Zj1x5UuovY4kqjkD7vir601VofPzABJYmMXev6JOO/9sn9rxslaojCTFG0Vxw1s/uZZ
CG3wsSO/Py7LmpuWpugTJmUjIfW8yTiYW7vuuReQkP6xchc2Q3ubyrkuCKMW1yJA9sX2/CLTnhnz
OY6UKW7kDFR+g+yK9AnFvexCvHaHs7qEAz/EiUaLScdca9gAZwU2WM/+dAn97cKlkwwdvTgZ3R9y
nKFw3hAC0TxlFxIpa1AeADqlx2BboBXNViGfDOLFG5v+dkFE5j0BImWW6tTm+1nZOtxr+hFKn4Lm
fXdVjBuueqaBy9/uaNw5psdt26dYPTCIlgYYZoPTUNt583IrVOjUKdVA64N69aF4ZcTHUr4in75Z
afxyQIytzWQFvuIZCKKBEbBCUtZWGG/0ZFV68BxXUWW0EeWy5oiHwP2fMKE7F/yDRKQ6fmZPa30p
msvfwWI4QFoCcZBh6+X0gMiNm2mtB9KP94NU57QB/7leCdx66KKufi/rR3CQIIh5zMCiyfPPr7Yq
nNqkkemUfkUYQCADXKgTcyD03ZDWtgs2f6Z8dLRdofjkEkJhehsWaocpRIAMxAl7sYUKFMO48rKw
DWt9bu3/JAgK8otqVINVtDGtDS+WyzsKath80EpNL0RTGDijhwCpCiPJ35ydzniduY4/OcVlbewy
lo4nXQHeYINyd90m2OJEq0jbmfiKU4/NAGtKUKOsOw5MqZQevjG0X+7sNPQ/4cDA87KrdSwHhYTU
9cKlkAVuCxb1a6Iakrsd8BpycyJyAIWaZxjREd0HKg6zNtjEGtXFmGLXFQFXmKNeWHOkQYIu3jA+
paFWaVbHtXwN2VfoM0Q4sJEavoWjN3dUa01XOlW0ZvLjwap9CMNZgT1nlCA0KiNeziTHzUW7AoXb
rwT2RJXSaKOoPVNXZO43M/4yRuIIpnlCqW6wxfvlBbmlOV9B6ezUDERSuhqoMx/Wl5cDXUQz1Eex
brz2LtfnxGoxgGAfYJLmXV20Gr013+uI7UCirhh+EW3q0aECUe847AvQrq82AOZ+jqg2nxy0WTJb
te65kTzfmNnZ9RUUswZE64K3+M9tb0AGaHaFnCZMhxLrnkJhmWTtFN/6AKlAy64AlFxShrxgnXwt
UnGkWsyEgjlt0DviWj7ShYjUBEouarosH15W7C2vj7FTul1GJSGyYu9KYVtDeKJMSLhhCn5LrXgm
HlVh73q7abB1/EJM+rcDwrhv58FE8A1nBjDoevKftHf5cABhBwG4qqA5NIWVNQLCi6TuDnwd6umo
IevsDe1JTnWFwR87wGhXXhiKAcl0qLnKuDao7+/dZ4tqzzVWbmvJeeLXSirVJWY0tWZXdxOGKLkA
6uYF/iIOd/B9DI87QOobRGk145nmKhV8oCo36+gFp228ftmiJKznvk79VL+22rx6/WogWWk0Jacz
raRLpfrt3s7RX+e7oX3N/SckGFj+YRW/ObENmIBg/PSrJ+JUT/kSHBrMcNLh5oLD7wdNOp6bR5bJ
oDdpQKf6bHDLFuay4ffwXvcIV9pGvDm0Aw4TFwDuuBcAFVxuX45wIAhH7+EukBXgFxZZO4aLPPSA
gRM/xMuz3gpqjbZuQJveA/Xptkkphzkk8d73m/RNouUxvvik9yl9D3XQHI7p5vml8DcjWB15QhlY
9kLFLVF+aP8Ckh1HIG/Hb5qKJG/+jv0N6jR5Tnc78ZinwiWRj2eQnLg1dwqFU7TfRwWfktD6x3Rn
24yV8P2pxXph8OKnL+Krdn/NkMzLwV9t74tNATJ/X3Wt+oWcISc4mrQwWhEmHbir6RpZLZVTPm0O
kHbz45QivKUcNRVl2P/qm8ALTF5L7EKk8aCA3EIMejijufIkzwX6lGi0KYfmimJKQ+h4zG3bNXqF
ADxYizR+zPHMQRfpoQy+UTMsiAkY9Ia8fcsq9U1LweL9IMXo7E/P8bYo7BpNsGZVh3Amaozd0RPY
UuVbkJp+fz85DtHHga/hdVvDwtQBXV1J6SYXUSjk2Jj2tXRnml+ZpzlVL0brumhxl8FmXSB0qnML
p294ksEb7K6mySpHIxFq+SXEUxiOzZOaNVY2n0ZXcePmPika7Pj9KH9bfkW7ZNOOAKhRnDBRNkeC
FdpGdH2P9Cd2ehH0XedS/Ji+2MiAA6UFQhGhmLhylx0sItOZr6/Othg0cXMmXWy409mIax0GRr8R
bxGXX3enB44hB4g+6DEhQd7ZKZvNUPs4zjb5aP2wPRxk1jdhkziHaLskEzdLxEW5bNJovY187uic
hlDuAPA04yPUr4C66EpB+yW+YAWN15l/BJTfUVNLkLBlJ3S39IgMGOMqR9DtC5nRwocQ6Dq/ChzS
y1M06hKHm0VyNgfG/3+6ASFeFtEvsYcYHHrrfxE8OQYtMhdZiAojT2q2TKMcQkPh91gmLNCSBLOC
eMs4gstsQ8eLBYn80WZyY07C5cJ+Keb0VFldBr/FeusD0XSEliHq3UOq+UpxHGdBGK4mzUnIlm7e
gVTYomFu6oKPLeDOUDxAfYQoiBX9x25znQa25ZOOaVUn9+/Nieg+n6W0Tprf7+9TjSHfSOfIZeNN
FYXm9lmBmzUzsyCspmHUGc2YJiKh1ORBPc3mK9WyNPPomy/6cZjwMPEgwXOZco3hY6IfwskcuiAu
wLga9Jd+n6RfQ6AKXh2AH2RbP+eZ1WgkRCJEZDwXUhjxaQ7+mihdgZ5OwGwJ7Cn0v4afh3RZmqX0
SgQbNFN5v1zYD86iGq3lv8pYstKX53cM7qDq3F6ZnEKtIDFLwbsP017itvjQecEV9hANE5tg+pWH
p9DMvVcMt8kQ0oYIHBe2aSErMLnpjaiPGp7qzSzwko9rECegdjaqvYV4r1aBnh+thphqv/A+uoEi
W8uZoygKRYnRlWqhyIBy81zQoXl0mRtXjy/2w13XNR8GsSTkxFIKq6o8IOjqGuBqG9h+i/T/8sgL
WN4MUncvtcwqEGBHGkxnKE1xwSpapEXMY8SCbYAeFpe5fs3tPXKQHhr57ZliSacSJdGHu4Op/nmZ
RkqtelduiNVcvxKZLMMf4kTW86+8OkZIgtiuw7sDSR75zNJHP1zQuBVzMlUO4g45JzGxSHGKzqMc
594zHtlgRLvJle9vQpEFsqtK2cS4YOcEhWpE3kawMOpYfuasKG1aHBNWDbEdW2MHtcKNbt1rHfez
cOvvxUWvsmL7ZuScUxULM2vwhJvd2lIlmTC1Gv8w6itAPHBeDQVe9Ayi81b/HkpXkYYbP98pqwNJ
Oe721LJTOWqgP2sl6VfD4ZUKLzStLfct57NVhEFup/LwHk0JtQschilT5LZwvwXlzyK9CIyVrJZR
ixnkQ2mqumw7Y+mCgawuhG446zzEHgHOsVAPc41WcvZlsJQ0VNXzo5XM8tlRHjnsbYrAZz2qjt3X
ZWJOukX5Yop+sgfh5b9xCwWsBZOmGM1K1O0Bd4E/z/b+ZZ9Ve6G/Drjjev1jXhLj6DY7lCsQZr38
p5X+FwUsiIPrpGU6VvAkeLpx0pAVQh+5CV2W3JhINElQ+fI+uVdk5oAXxgabIMR9lNjlQpCNkhCU
YI/ZBqV7179Y4uDBW2r2JVV70+FBpLoQpn9BpH8bI6iMKeMuCArHcHfp6NmuxoHtMZVSwO5nJ+sy
YkIHruqi0gUc2RubSDFvo67v42WFVP2XLvolGdXivN3SVh5y3H3su4cyvMRAwBrwgwJksg+8EncA
37gI+FYn4CFuCH5bn6RUrgBYVL3/+gwXpc0wTBETOFdIbrroHcMfTUPYUQkwiUXp7LB0xEQbPVRn
GzAKqGQUi598wgzhpRea+8qNAmhe0NGjUgq+KT0A9TmzmpGEGH5noDQx3x2mpTBycpzivODdYoTn
BlfMSj7c3kOQlgWSpeo6XHCzei+6dkQCvM9OwGemErpp4rZzX3P68+7Ijs3C+bu1oYjlcuN2ADgh
cbPbevS3vsHY6/WFYCygSxNAzbFBgKnlgeuiPkqknVraQulcSpBR45zbIeM/wREzAQAWVIFjyxXu
mYXXKuZQ1atlW3eYnEFT4EeSII6/4yR9u21V8jQou67X2PBRiNsMzpQR935VokNUugBGJYp7ZxB4
zSx0j7Lsay2uCTpjJtD2lRppxsnQLwvkzzxK2PMmEdwgEXJ2HF870LZs2xsV4BJ3s77ZyWMBKS9w
7BAwEIF1PHm/RGT3x6fQITPIlM9LedLjoTWKwMgVvN6GUUp7PiKUUPmvE4sBZeTG/ELTWINCqnPB
OVTgns8XMOpM0Mf7BJScLT47EwLb+VEVrKTEgICGRS0XdLK/zIa8+RJIyBQBHBVym35O2QrO5nWo
FrAL8EnYBwl1zfpydngNru+ZCSYB4YCgYRU5wZ8PCbzUkwMsH+vTCTZJl1ZIN7hAcKXaQMCg1mma
C5oyjFANtI1YTa3WJqPoYwLRaxuPgU9yAycvjkRnVwFWVMSgzl1YKKDblE6/bUGS8qEBKEC+9gQa
pts9tclDNmzGTa/G+lLvzxYMR2DEtFUgavHpHt5QsqP+omdPZF5eLzkHYP0Y7Qq5Gr7mGVmhx0VF
oc9gMY+rDMEPK3sK4lxmm295i3iJBNGvLrxmPD2IGSy0kS3Fi/grxFBLa5FqARdO3pR3RAOj5VOp
xv0sQIOmkiqCgbI+IbHlfkHjfjadsfR7tMYZwpG6Irrq/sCNU8fPTCjd3ABslT4IwjPKh+xrBGVB
1PuAHpdTXU40CP5LtMnVTc5V8n5bXnvGMXUzzPVLEiPADoB7CUZVFgZ9OY/zFn0z5qRhzl7kqTbJ
u0gY/0W+EtfpAVTI4oEVIt7FJNq8QzHHKZuXBAeh17RLjL5+erRmFRX3akTlSw4sDPO734OrQeyg
pI2Lbz7XXr7nDTfrnL8lAPwvXfir3MK+A9tmT5gLkGLi/rju2kJyj9UdTy0/ZPLWQchwZ+oh87Q0
ZAXssHkIwhe5Hx6rXG7l86WknQUCzWOqnJCCx/Mb1OcCvOAoo8rmQAQPgbwS2je90mT7EziPIoMA
fcCWi+5WgafQYFlRwx4CRpQFLP7U/BYdL4+FYrR8pYk1TY3lAgrO3G3W3KCC0U434NGgjr9cuOho
T1IcMSNDAn15mNz7inXfVisocIC+rR8jGig4QUsBbqBU7zEZ4wkVabfczwiIH9yZFlfBr8ZCeaAy
yoiyM5o1yy78Y8LZNKuf4INzf2NrOu353GXMDzQ3WfXheb/D4wGrsDHVxwJYmE4QWbX29yjVaCP+
GbtutncydYPxMouHH0Tme0ywlnEabG3Q4RutkjQuTeiA/sNoQYi9UWqiIEzgFljZVAHayP2TSq2c
lfY4dCtE3Fw26v4xejyWuksb+aioqfLPAa5tKJR+LmNLqehrbG0q7tFn4KNkdYHMaqdyhIO5DW+l
v50LT1nvozhKj5ahRvro5bdRguR2ums4k+b/kydducKmjyRm6qrDadO9OT50lAXkJrrOfm4wdBku
DiDBRTwrMNNdO8coB0YWB2P+q2Z6lxsvHkwOF78k66QmM5uiMkBJNnMyS+R0DEJ8yz40RfMM3aMi
lmzIzoe5bWTk4IAK/UnlQtD4uIR01Pcmp/WuS6TrcY1K41va9ZQcf0Z6iJPtwlT2tnyllQ+jJ1D0
4raSy1/VkRQ5u5FKcKLPrznuyGasMNknuzKRK3Kin6CY1DReIO2WFLjy+GBEVAIbcdCNpFNMZeFB
PUThomJ/nxLzRDysGGbjtRUKqFbj//CfqIJxHA8somdUNBi07XTnMEGFQs9EdbeVQB2LFn8nxs+V
N07kTwaWIldneQ+0nqRt60XH1DfCXwRDKOowGex06lUcifcp02DPWlYnAQYKPtGCWqDa4z5oEvEo
h4P/3AMga0hWNLPtC1ItRbtB49Gn7BP8XRna7wHLobDxatudjCXdlauf1atMrAsJvBaQTwm/3F/8
isX9I88JFK8bAZvxiJ+DJWCAtS9Ytmqiu5oED+Kem6dOBScC/hWfrd27SJXMLJBPH+8bTIW+nLUW
HfVIft3SjwWku/zAs1zRA4a/DInHOYPf3T7e8krrPxhtL+1i+Ak4ucaMXkhUMhr2CWS24c7eOEmQ
ne06CLQDNmggJE4cp263sPt+eHiQpe2phhRjC+DtGiy894h9LR9cr/qk1yMNKlcZ8F5sTt5ImYEM
ZIoJXIoRFRPKG9xbT48r1CeDDVSvquLzcGTeFfHyw+RVr1Op0WqfivROb8zvRYXr4vDPVMprb02R
nzhz+IeGwBkmRFstb1waZz4rd+HGq2Xj0jUAxRhy6gmZytK+yD5rNdQF/oCfAzlfrx/6FpBkTQZN
bIF5kAh34we4aTNv6V5GwwZfOQixAcY6YRN2SJtSJH8y33lrZjhieQjSa91NIs/yAPc1fq1GAVIk
mmFDA4xjVHTMPukcpZJ0kCAnEkJURo8PKA58TpDbfOORm4HDiy/albEWeqj620iW2pTfm7F8TLWA
wRDniQ13Sg2TfluR9mx5+QyxAD1RMFAG3cW4Aco1qUt48fn9WbxlBsEv5znYIkLtVUs0dkh4eVdC
vx1KyAz6tfE6Qb1u9C48G3edpE9MbekwQSjiDcy0FNGQC1TxIYCoN+0Muy26DMXv/beNKXPHf+u1
5yPyRiTAXF+Tm1rjj6KGZz7fS/ua/8o32RGvOUoWuegWfJBhyfhYeyQGgZGfIDnfYV+n3yQ0RY64
MLt8LFpifymq/d/OgCAK0WW6IcmIdc0qyHbhMG2mVtrbQHhNVazMy3qXcaWGjslYkf7ko5nopOH+
zkwnNzRH20jyrGO69hkg8oqp8ycbmSofNTqJp7gNgKVLCUuq4HHtf7+2HFY22LgYTZs62Ujp92Tq
LAftqdMvYGg3ueo6z8vHs8GM5X0GFUjRhnGWXSicoObQkT1RxrqI/v+9oGnpXcMJc3ADF9CHpn3/
BWRiemTLDodFfdfKBPWFeQbfKBgDw7a1O93gaiYNao+yI/o5QjtfSLbLI2xYPP5eGpK0r27o7/6O
JyNGmzqbGgl01jaBoZqg/eH3Z6Rl0n5uYg81jRS5qlQaidHMtrZsPTLxrjhHPVriL0XhAu/Xryuc
vpOpAGXPM29QEfqPjNT2UmQZskZ2Kwz9xRvUwYKzIJmiIz2HKhfIYKvVlIP6qCA00jiyNlZu51fl
lvPClZMq44zEtrPBffd582Mwg14/zZr2kxWxG5sGPd0vEbUTm0cZhXv0085SUpMIKnbHMNYXy2ej
QhqfYDpu8RWo+aG1lu6nTx+jHeMF2OOmR0IqERosIzlIRqntfQXmjtgtSLGnerhy8rC3eaSFTvf8
1flnjt4wVEtdPDBwUKKk7k+iBDPgkTvfqIw9l9Cq+KfmJXHRjaEjtMozGDtUlZvecq9ikqBQz5OH
68N5brttopHskLyyUZ/wGC3v76JrRKyba/2Rsr3kozrl3uKw1wRLmrorNeDjdlMMQiTw1ZZSzsDO
EFikKk8f9HNRjgMU0PZmv/6jMoN65MWuYyurSioz+VxJIBqp6TvgvGTK08XlDAtSBlN0NIym6zLp
28rA8Z+EEcnbsDzar1ZU4zWTEaHIQIdALHTR5ZUh4bdqnBD1oaz5bl4dxp77xBrK4ujwfQ/BF4Dd
AhdBmStI+Ztn5qlA5NE3rdSd1OColfpgedK379RkiBOu1vcIFYMg+PQCWYQAXSm2O0q3fWVVqMCW
SR8VLghH2mQgB883vyhFi4B/aXwrJvr9zF6+a+3SDxx6C1RYlvBdNbJWSgcB9ESYhW4HV6k73AYy
noAnId7aCu5ghlhraPEkxQX4lkxult2dF5cOZKBPc86IRFhhPbgmwTpbUlwimrPOJ/np8lbRBybH
f975aFinbFl3Klkp9YrsXmLr+r6hF+3hMEQxFEde57Nni5CteBDAHgUL6YHOtGLKwSCUk37ckZWN
fwjvY+y/u85fJtl6OIOfsCk2KIXMeoHnCaqX7ugGLLemk9MjWgWOTMLLwUnAWFRgZAcMvEXddIRr
0THgxestcL7INXdn8iiYGU+xm4hRoKyAovFlAQ+dbNiadaYk+2Arp57M24cclzhL0uQ8gh1yKLTq
Z2GwR/mtM5LCKV758KZCLjbCm5njZ0GX79NxMuo3QchaTjhfAqzs4BfUbqkzn28FPSfSTMB0gIL9
XDl2S6hJAudWUI4fBAtqI5CboGM3sXXIn0slInJVeATbdOD2MWsH7LyINNZ698eO8FOZSCVnOKzp
fvL9Dzl2xwDcmQRN4GQiJdrWJ/oU2mIGHPbbz/0lOURKWVkHWh3fPVLlX/zV48Ix5GbuhVhOkPiD
7jzLpT6jrjfwdENm+ZBgUS+3WxayLlrkZis2NtlDUP77K6Ijl5xF8or19A1fXR31bKhUb8qIBFNB
CtS10Cz5PGheiCwFyVOoORHLDbAB7wPhAhVNdMszdIfCY42nG5vTc0raBmQaoTFkpGjz6NErrR0i
YsubzfeiLF9QFVBGmvPAAMQnIF7aXkxgOiV5J49ab/aWWk9hciV6OKRbISpmCc16g3mUzRQUGgZ3
pZo98roE1efXFe9J2ev8FtltdWHbyL63i8XSM3zp/fVK2qTo0yd4mzn0KsuWzV2Lxor6dFisPF00
4yhYtJmH6obMz5LKT/hUQ7iyEC2l9vXZlKDHEQB8Jl3UkA01+M8hxqy2xItPjE8e0KyxsJkG07TV
o7NI8LTsHEZKKWYMOwh2icz2lED5quxMFWvU8jecXRhO8iSwUCfCnci0T4R3musL3iA1W81cEv9v
aQDVsm32LSira8e5oIpAScUXGh5OOMVyYD3lFxVOZwOY//cydBjv1gAFAknbxQ0LEVNy8FaxtSUI
sIxjUDggaJWi+zC0sMczdi/yY9XM+/QeeJ6IpXtIHfx5FGl+oWIctPq+pFW1Zx3JF9SFf+tKYFie
iMLiu29+zsZwL2DpoKhO30CPVcrkCjq8AHwYJuuHrLazOGrONIVqgqr9tk9TaMXWDurb3FtNEL5M
pXqp/ssBAKUjGomMxyb2wj3jRGDnxKkIWDHKMxT/iAdIerOyDyaNEblG11aZ/htZhOtoec/jaA02
6auJA4opVES80rqXgBdcuZTutwZYXqBQ4KwMHswwtgKmkO7RNkxhIqGZavjA9eIGEGgGqTb5vVb1
LwFl7t8c4Qf8p90bhLsoCGcrd8rjCklyLTzqLJSfABpseIkRG3ZF1sKvdZnnluctmHhXFosxAe3Z
uXPqxLe16WHGEDxoAkKK/usg8tEGIaj0JOCXxSCoAxS+zP1N5YKF1BFgNQtZr40JhTzEW93gA0r3
Qfo1WMbVRLfYv4PSpb4wgekidJU8nn9SuSQIJceont21+HwEQuFA+qSVXL+iNshbLHNIq0vcY+5k
7G9jnmFxFYdnU+kpox+x+MdSCSNz3tcEj+B2JoeO1Pw8Iqd6xNjRNppLlhtDupSLP/BW0AIrmmLh
PqKC1Ko5n0y4YACVcN4k8bHLJFnVH9d3OVlJLscFmp3JQ71yID3cU4KWO08ElkwcLG5GgxymOX+E
9goYwFvBmbWdWJn2DHkW9Aoz9zNj+ej/ItRnEOhUil2dcpOcsuDJnykoF21lat9/SKUd9LqWqJQL
1GrAv+Vk8Kof88YB90iric9F68gu6B9KjBnf+xOlrwqsKG5J2yS88lztRWHZmWCk4w9dweMbn2cK
mEkmljFUBCXo/u2pUUf9nDYTbWiPSUc1UEy5w8a1n/NFGzhYBylX5BxkQSuWRVR7hUyHohwj2FVM
K1WsQhk+gHUwqQTjzI9nrWO5Zi6uX/+OYmhoDJ9hn9gop/kK1KwVS7UT5lHWtnpxZ8BgjNrjW0si
lBgjMyHPdzN3GDywGfl4u7YXnk+gX8NiJNDqdrqSIGYEwbrV0idfYYotp90jH7j1Vpubjt3y+ve8
2GOcqaoUHLXPM9ryS3urGliseh6f+ETdILvm0k2X9E3LXMQUuv27+DIg9GQPQ8O6Yypk1g/k8ZM6
aXpR0NiS9qxTAaYXVY0XilinoruSMgcqk5lYgi8KS15eWmBlkMAnrlQQwqAu2XmubJi/bnVNMfe/
npGHkUS7VKvbeSFBxp5YyhOVUSHqTHdmQI2a8u6SJV3wLuY2WxOa7ZLj7dK3qsECHlbUUaKp78qQ
wIAOhw7/g3LmkQC5T9Hoqr4cZ6HDRSCfWkrIr8FUkFnYOu5IfmCMRY9/3apbSsefdtrtxWfMS2HB
rYOweBWS3owx+7prDA3xJIoEFJSQODbrh2eGdoJpAtDDzVs2SgoBfGBl+4gchzbMtnmh29sFEu4N
HU5V9JLm4dGSHqpFIdmYJFlrTPammhVP0DC9K26Eyf3MLeunf5Y9qVZATLGPrTfw7/QSk5C2HIR0
Pk/E1eI8PbN/ZKFsiZMOOcEG4GaiZlbGFGT/AFw4EHOBktQEjMOJhp2qAXXZV1a5zXDJeEXEOQv6
RmBfPvFVKtD3BuAkR143wVd3D7YL1/kGH4QfMjpkdiyMCQqkW3X8AkM0CCoCd5DkAxcJKaFtlLzh
Z+rhiEU765ZKnZeTO2Y3CSjm4Ac6WNXKVKDgIiMEso8yr4pWtYRtdqMQTwZzzEqARwaDg/oPglUO
aGXdLn8KZzf4P4J8wDvbO3ghC99Fn8vQ0jsGZLMu65H9MP0oFuCpSYDtTFeKZk5l77hKtUzEpXHG
un7paSSNdBSBAjrtlBu64Iz/LXv0dnm0QImDPQxJYyZtcX+hGgUaZlU0dlFH069txtNNcC1jATGq
v7CtjrRedJWTnpbzyJw3RFMgukrMDRZAOyXOG18HfuJMbqKPNniBjrkuxa0T04G6v88kmAILF33o
dzbjRH06Gt50iwF4YivPrFiNhROrx647CmAAALBNooIJ6m5q+xl0kBNPNkuE/5h6n+Do7tO4SllZ
bWd2dcL7Lgw2FyLMf08lZ1vPRhjRCKdPWdVQGa2SSABS/edZXaTWBVl3ByH3RQbd59xFrcXi7df7
HQwpAks2gA0HiH5cfTWtQIzs7hncqSN5TH2nEUVy+Rx8EsYXzYpKtf/eH95o1xthv8MPAXr7PB7z
MqJO1JDrdFG6XwuUn82+JHGdqYWlAzHn55nyE4Q7eL/iUklzfpFkFIFFWePpJh5W7MNrYsMKpZtf
SBTicVb3+3QxjN4EZiX3niLutQJPQImf/Ew7tyKjvBOCrxhZwrMAGRbJplITR87L08bwTPdvjMd8
QCQU1TdxPT+GcCLrd/4P6kC4pBldyzK0STXtmoYu4WwIfFPkhLcZf2D9mVwi2p+NSHpX5JM6vmy8
F5DcRkNYnEj/br522NP0nBp4uCNZpxOa5OzR7nGvF8NSEJTD9RCWXiAhtgeUYNhILGeeEIsNH8pT
FrgxVITXAfv1SaTKm+BivT6YjlVFijZ9aQGVHFRnqp2CgeSaF/wbMQlR2SpqFc7iRYTPPRwBZkBY
MxWmu0IfULyKn+3AzZYRC4YRMskUmZ5GRL2ZzBbCQ7D6EeitQGA96ZZte7EtEwGVewSJSfhGWSc+
kT5JmDwDL9E6Bg75VUFCoYLYO59LOEoZDlT6qWKvo4GIUkkiZ6nlD8fIUBlF5JZTN5mdPNYHqpHp
3yRYk5zxZoGNuBnnYkqvJRBK+FUIabu0hk/ZAd76zAmHA1ByktHdZuMwQMnnBSLfkSzn3VMbvz9w
9zuiNPwUx9eVOQKsg2uBzGFAQ3RZUWhZBNE8M1sj96xePdeQoyzct6nyNmttCpjLCafFXzXiXhz2
OQQAgU9tWZe4LqysVVmFxa59ahANPqoc2qNe3iAvy0ihDpr1b3Ctm/VnoOaq0X0kwAYNwz2D5Nam
MSfho+8uxF/L7142gxbmDKx7NkBSENNiOunCHylV9nPtV6iP34Dmts/1gCtPA4zdTT+9Ctf4tz/9
DPX24f7yJNM6tG4+hBk+Cx7RsNjV0EPaEHjGDd2kO54QSUXVbO6jn8TVPJn+S7U1d31NdmxvPyf5
fLaHbnGILaeW64M46UXdbiAE/7KdEE1wNRk46rzn3P8SWTkZXR86PPjONorFGrcruu8GDdnv9rlL
iOBccSy9EKPpVbEY/1kGoiaHezPLf4rmwQQCMf7mQ4W4F3NPcOYza5dAs+guGsesiqOduzv7eK8e
noV+TsP13nlZjrUXYzw1Jqo0Isx3Dhh419za1SraIcMTCtsErXiEhd7ycTmmrNOAr9ECwSFPsTiE
oa3E6FNJtCOlAUzC0WMKAdyvG7e7tB8yzr1RgQLsgMH3MlFzxV3mI8A1xQ6rtFzQtqkjz2RpTR8z
GwgIwGNLaZfFxvuVy3BhLBFnBoktdYYk2u1w1UqoxD1qSvNJAOk6AaB81nElSKhgd0qOku5H2Anw
9QwWB2kM/29S93qwWjk9D8im+vP1j4W48T9miEWK7izQwzKtD3aNUZD2SqO5lCJceCD3Sg3ATWpp
DIAfj+0BY2HiSWFNzhn2nkJRbzVYX/RtvljLnn9imFoPXYLVQZawGb38zx0P1hlQiE7mTfZ3foLj
ob4eo6jikA5a0C/+KmQR/GmPrG6oiepjkwKOOqQxqJlskVsr6jE1OHFSwvhkY9U3ai3hfF9MT7QT
MOd4j+YUk2DB0IHcdO7gvRhmxzl27EsmKBmrM61edsMhH+7dXXY06ouMums/3dDqvNLqwHhB3xQg
nUGXevhY3PjBLGHkActHacUjuqpS8OFklACArPeLiJTq6L+ezcIuQzSrx8PvVUtoJhG0Q4QaBkP5
BFRK92lsEpl8ME8HEq9JYlOwWgpILVuELgHZ9IBe2H7f1J5RRIbTGKi2JpIre2dH6uVU7LMDMe1Z
mAHadZ59tvHeMKooqQ/0BS84kMqHxbZgZPh48vmfzI0a0fVwQrTtZCHUm5UTTaKJdHn44MWnLK6/
hw5tiCw7tiq21gQwgYsG6C7+tfYCUhrJMgNy7XDq+o1wk5wZdgWuwpt7fGPhaGWRE0bFXeP1ITn6
GoTn05qEGltW60/NyOzNYjSXjLb3BbV62qbOKLUbQ6VHz3SYArErH3xL3UxRJKXM6kJ0fSOAiy2d
WGeRdI8InKYwHX+x0h9D1m0civoYJ8HHOOElWaO33JpW5AI2v/30TgDS7RqU3zPqvAlmpuWpkT4F
XkZciXsm28egTrjJ6muy0zGPxpAWZbJUC49Q1s034SVyCO8vXNCVJWPOxZDy74PhWEBVwvU6dJjn
1tPoUm7UkEwd1i6MSEOvOT+fpzHxI40xCH/U1PNAh7ph/7xz4bGyiX5JSJGS4vgEIUNSj35o3Kpt
qmwoxhfC8qeeJnimbJgUMdTcLiTmxalxILaeMoszb7bXCX1eFfxiuyxi8jjd0iKrawQob2ANIUSf
xUmQ2wgrOlz64aVaUGsU1hMWD3GQuiIf9nxjl8iEn0Y0laKZftgSkAxCjVmj2EIHVlJtGLg1oQYi
9hsjVsyo5pxVVe07t3VdkckxZKZtu/iEUdgTP0QuAC8kGgkB18DmRAqF4OREyvOTEjRqe9XXoFpl
csXsK4AGUYucVfVLHhpahlX+ZX1Si//xAY+PElcIVRm//MWPPG1Nv52HLyHsmpuDsNLSNtYcNtCa
HRJQVcoKTt0IuRp6URXPyp6o+wMwuBANtW6jADK4bdHkmXE8kW/MuU1H4QQ7Gd/MUD3jUGXYm2la
jldtoKujeu0ELVU7WwTK/mkRxxoidFbYcorza1v65sXKI5XO1RZv1iObg23Mu+d2ywKUmZg2/un9
RRteYqjhzD7y8fBCbd79DuAocUB8QJ03XQoHnnuaijAFruzK1v6ZwivOI32Qt4RuLkcugkZ8cKOd
Y8Ru5xR1+ltGovrybdwF7BJM9b5qlUyMcS5UCvt0RfCBGk95Q9tRg3n+W2VKA3SLO+XaU+8ddN45
2W9z9MnYIGex9aIceLyWYYYx0ZgFiU8T7jCW7QEUbmYN4rnwX4PszuwNaLrRGWVe34Jy8DBcOAOJ
tsHtTygg8eeoJ+kP6jByaHTQ0I0iuSNxBQVJInwP4HKa7ljeBCpY9SV6Vp03teyHImqQvNbI/kff
/Dt9EhSzORBOzOdvKSlIS+lY4/9vcJdCs3o1GIVGD4mL4/w43lZp74X2N60O2EfVg/3h/BTiRoVp
47SQH86arYRqbP/8iiWT2oT9EJIDPXqzinx45D2ovFKlGXbOEFTqNGph8PZDw7nv6lcLbIeluibn
pOo3LgpOPMp53ZXEcG+9IzMIj1sZnBRdlFMjfQYdwu4AWyg6Br+qsZFiJW7EtQl7gL5NAP09UTjG
FOt1udcydjcVSHRe0ussbpXlx6pp7ONwo89aAf436dbR1eV2ZpH2NS3UoCjHIvnmutZNxRNtUDD3
YCJseE1sWE5NmWYiSqrRGsjG9RX9L6eG0p6sdbTRV0FPp4D4+XaPdxwt0dSQzEphV9J0ElbF2y6y
rE6bzbm8fXybj+pTj5W3Td+Fr7sSff3fQ+5+pbd+F4k3KiHRW+2WWBf4OceOM625kO9O+mpgC+UF
56C1WTy1LpDqNVsVbD3YmRpP8g9ZIweY8dPooZpfAGOWiIefreFMokUhFiTjAlxM+s00YsUWCEg6
mX3AngnWwmsIkDKiG0zSO9wC7OF2UBpfjLrjXKm94qQ3wCbsB8pwgb+11y6ZDrxCZxcXmXt9yCeH
p3gbdBa9xHwxhN1C0Vlnxdf5XNCxx5/TxCfhzSEbTi3qBAxxoN313257jaJ2EI98H7AqVi9cq/x9
rYzGRTYzxEPHvYlTWWuCnnbEJKDvan5FrCC3lMoupLBJBpOOUn3wRw6W16lRrPlEbwU0xzTH7cBH
tq9Rne2cliUt6u4Wfiy64uYfmd6jwztx5RfXpp2SV6Ca7n9PnK0By5NbPbflGBH7iBsnQr5dmTOw
9kKPvz0AzWX90dvw2FyD3iLgkfXjNuL+5bxHnAd4tb4aVqD4XpcITYAL24G6nEWMNqWqS7cGlrHb
AQOgiNxGXf/b7bd/QZL9XUXMBYwd7SvXHkXu7p2FZwPZQLYQV7QsmGaFGiaSp2aAkdXFD0v4Gav8
wgqK4/ukzI+VLQ8x+3aqtuYfOFTNthxRruf+qzDNjUvQzDg6EgUzDaHnd4jMmdB21OVItuWJoYdQ
S8WbMONVRM0f5fD5w8POuePaOXu/1hwR5aZqHvwmdAmPG8yiXl29xxaa5BolIgyZVnpzQKUAHTBR
HrGXrBbr24ETAs2mioNMgRyY5CV9+eCWh9kxuj+1gB8XzyOsZfb2UW4xjiqy0iBOuNBlFJNY8Iva
ne9mkdBvVS5E5smv2ulR+QtM8mWqljydqxDVso5kMuypCoibHUFKEHwwwqhR3GlLhj7IB1ktLJzH
8lIamN/SibGYtDW+41+vRKhaGriALz1PeoYfErmPBDbW0SAqhgm7tvEyJgH+6Cj6pYbhtEroJZeb
AIqFbC2lfSgK1xh5O4n/bgH0K+8xLz2v1qtxNvquVeQZ+mm3m+n0TLh8SMfdYOzlWvta7ELFI8qr
MR770oeNb7b2szdtiNUROQEY73da/7/9hBcs6e1GH4b3qU5PBaeGgDtGGe5J87O5TBwSDhYia56X
CU2+j/jsaXxhAbAcGyhk4rzTYHCnQ8caKpLFdSLKHyd68jlNok5XQVQaRnoNdCaKR0vH2rA8sJOS
wrwBCHNFy1BROcjiQQLcG0hyGHNEoYtSurTNG8BEsr9jTAjJ5j7vYimhhEaCfLes5Xtlnllu4Tqb
Y6WeNCpY1iaAMVeYweBZaSsUN1NNLJh6cRWiDkEF460cKdE3fgYIU1SeNq33eP33r4j5WEh9ADEm
EkV1CEJvBwblrQ01xZf6cpFLWkDdP5OHCOQHV+kxtu4MVn78QWjFih3eq4mKotY6Nn1Eg3uSIZ8a
EJSfIfEVTb9cWn+OIb83a8uUGBZyPxfdDBorF69i3Hae282nXnS+eqg14DB13UocNF95pyCUbS42
S/9bIYCjUmwdtgHUFB1WeVBh9pM4tOgkK1ZsGyVdbbFfPZJk4ewvPKDVJH3SkQDIflRisYOLn3Rx
EMRxAe+Rm0YWBB8fmfkj3KTf4Ni9Yhu8rTT1A1G6FDM0hX+ISkKeJynK2BYEKrhReSkQrvjhGuU2
ztlwogy3cj102tuZ00a/J/LGWWKg5Xdpz9zKJoN/spr5WcCsi/n07Ib0zJhMREdZ4z/58aOPpLRr
kVFD9fdSTfM9Jeu78DPdNSIt9/jaUtHH+ivA2Wl4+ONTZ5McPebLOybBppNAcy9UAIyVnnhMfS1a
KJFQ88a5AZnuI6dtaFHBLyvREKIRN6aZmHBmYgNtNR3mpsKB71e4ZvSm0eSHUJJA0QeHhuq+JEGC
fUvnsXtblQAgmyCrmIpKvK40bwbODbfHNNK91OUuDkm63qZkpKeIpiCQLS/IeP5Kh1cnQuTHrnxc
ly/fQ0ZV8B/fI2f6elhjhj1BNUqcbq9hfafAniIGjtvMjbF2dQ7edP2rKTrjzu66k4oe33xN3DTl
JfnuvfcMk6LCQCH1FCkYub3zohjFime+ZorUGDw4vMkA9Ik8ZTRJ6ew/8w9IBf6PrS5Tcgsx0rH/
mKWRRweQiEJZB5k368d/VVV23VDJIYc0CNU+IdK7be7Bk/CjE0jyoSQ7KV8FvtXvkvp7UJ/EBKR5
cWLv9ovt4L+MpGp250IpPx0KzuSAQnjuXMN5dfQk2hQtdtn2I9h0B9uc/2IkyU9ZgE4J36jQObXC
aLx/xiQCsxKECZV6F5tnMYHNOEIf8jiHGp7zhYib4e9GZthx8l5guUiSkUfpz650Vupijs5wiyAq
cwWn5ZHN4mrkA1mFA8XeUWz/BaArKrhonG7T5EXYDZ+RU9u3vs7UgrHhTvgzKRctkWkL8+5xfFTE
c+2QDsj0alGDTht0fkt2xOauGOpaBGsvyGA3R+iD0SSjZa1Xw/UOksHNTqA14NqAEzqY3syGYBmv
/bgErqc58BQXW1SSxnwPQn9EoFqEmYKSlJIKXsqBT2x+i+OjfWhNFg9GciUPEqfCRvAQYApSaLb4
u9dQiV5WMyfoDghiquaY0+0Pe2RgwBJvwOLfaBJaY0eG2WTNVXt6Va9PM9dD9Eq3Ku98z/Zc4csB
yaPfbJ0HdKu3cAiWCeVcViVyGpkA+U1LQA1jrKRf3yvubjTXIs/z+2BYe5MHF/WQUdaSbaKZzmIp
M7DrnTTkh8bmwHUxxf0JK/9pKgV3EJfZwFeMo5NuOlCkLrPzdB0eYt8nmDIB2PSbZQflrhJq4zOS
ukp3/AxsjxICTwsAtcNgHRjCiukegvDUtmbQl6ZvC4AIjxbXCyWbWs3UDfTok63z3qOVNh0p8DZd
ks9Af2IhV/dQsLqASINL4i5gzlaZA/vM7dfpP2Cr7aIeIWUXmWlDIS5G4bLWTo7T5mlg1HFg5vVS
9vp2wiuSYuyWwQeEpodIbh+H/7Gcy6Wv5W3SVVz0wTyP89RHznt8nBn3lJ5AbmvBws8o5RMLsHOr
fwl1uBChT9ONBU5JEShdjJvfPApJK8pXpuuORiPoTzb+XsRu3e9MAFvAoMNoHJJ4dj4eQWjD5rKc
RyS0izy0ktwLS5Lp1nIxyXpQBe/BJAScVCKqJ4BOtzd1+C7w22OwVipHI+kuX9B4pHizozAdpg1K
vM7kKrPVGLJCHBqV8pobDC+Dg7/sg45I6dPSY0hm+7Ek71YxB00N7EdQ+KdqSgygB0xATjXSncnt
flLdkbBEhwq+mRYVvAZsi0s/aTuLNN5PZCKJ7maCmTHELmP+F0i7hboQL8ezHvPA9TDAeLTpBIR1
QAc8R4T5AUMmWyRQvErfCwDtu+j4lfc6507CfFwZ5Xm2n4BjpzZxCx9QPIoBfXDZqqOR22YEo6zt
3kuQHxwBNh0+6Zj7T9lvycWVolkWyCZGwwnUpHqPZCf447eb7yLfXBREATrG7VhiKZ17FgLXknS8
xL4dhroeo0ooXjkwuNSKUud48o/AAGKr1AOOfgzUpSS8QDfr6SrP1yx2lU29EFUrld2X43zgPCwc
a8w5wZItFAUY1EZLAIBE8hFvbFrZziZhyNJDrwsMXYbnPH9g07nVOQEkOELnK0jqLO1QAxPXlJ4w
q2mw9qypkd1xUNFofcNGvjLMJH/5FQvslKED9OTpSFMORFXw+AZtGc6k8cP5fzmPwMVZR4xPT72K
Ch6tmhkUSqMZZJxWmclB3S4WGgisx1Aw33WP5+p/b5toTbkswLYcC97GDlwAx6Zd6L0H7k5noKsW
pp3cp0s5/DabvcrwOjthcSqeONwhlxIVXFuE8jXlyRxYobhy8zFk01UkZ1sMDe1mhid5VBAda1gV
G2nJi0UzhnkPMheHCKxrwi+21sFXCHODQCVD/Sui9JGzHD6BuNYQ4GYNJRncOXa3slyMhGlIWZ9D
UeS/ubq6p/5G/jux5b0vtGOl0qtewPkhx7CCmCbxVoYEIqLIuEeKwWQXDTfl1f71nyX/iPGM1h3u
V/Uji+1Aetv2swBXtEiimLALiRsIqgDQc9Ti2vLVE6Ce035RB+203WyxyAsSyUhX0ILMon0NcZUB
shmxU8rvirCWYpGoZporRj6SoCqMCY7iIjlnMM5qdgow+dPM9/gQCQxkp/BYzThyo2HzeeC+oKnB
jBgHrx7hGE7NGq5WveMlFjqaCbpbtKsJFMoWM9lWqsMOlcZIwvTrgDYw5QGvklv8AI+O07CE0dHS
TDLodCFALlZEIZVb6ofCaaurZ0cL6bmmaYpitMUIHh81YI6aVEYVhF0TQednnSnqTl41ZcsQHLJf
9GnlmIdpKSyxvM2RB4kUosgH7paZk3WLnge4mwSDnAJUQkE8rV6McviETDsiO5pODtjMtpI7z3os
dwRXRN1lsAoE3/WwJnyVClASip4a/GlpZ6VJUt0Wo2SXtI7DIYZNxoXyf/UtH8G8NYv5W6KvoQph
K3ehoq/gIYKoHOEdAa/0qytNrEJz20Rs/2mjwZdiMroE/jvpfzu3g69uyGGIoGZbOhRYDuSKG5S1
cp/GHVoQ0MgEUV0Hu+1hX4uoR8VnkjjkskHq29ujtMsrG6296rh/VaP4baCN4m97+NFS6A2JpQAX
fxHAr4ARNpuAo+LoZ4YlXpqEVBw42OV7MByUuAoI64kqLrsFbpb0oflBoc+B7Ov851RUP+7Pm3au
qEhSHB6CpdyN2gKapigOHllmrRU5ds2MmslLfdbOIV/qIhdLS/dawC+tBK4CfznKK2CrvXaKIlqR
chzCkKHQFlIm1zXRFaQ8eSIeEtnXxATBByQzZN1OqqhskurZCkfinKLEbBDEsqJvTOpwJg+p6KNw
cYsBd6SNyfn79eTZfvFFuaBx9A3txbfe1jVMayFfbNDWryvMl1x1+GAei1JFxtxPwACfZfjuaunJ
bfihnGDkIbwGkRuCK3tPChcSI0Pr2By09F7vfEvr/ZZr9v4Y+mIy+SQEb+iofuVkVcy4W6TgtAXV
jW9zlrxfiEaDeLBiWJ5l+EN0zQaqDRgpVWN8N4hlcsuA3pQvThWdxOpWp8IbjJ0IDakpypVxAHj1
8EuotpTKw+wl3iVRX8Hw0PFjCYDRNEOGox+1M/fpSjZFrk4kJyUTHsrF2JhPpyFNvW92Rc8dKYrf
n4csovDPGLKpGSK4o6N5ChAh0/tnmmdCrh+FqnCUYuXARHArh7h9ENEFIErmoRk/F2WkD9i4GUzr
ylNvDXEdGzq5QPK89ACNJ5MjImr+x6MPy7VjpFjvtXEPF0qGAsLfoIiGaZTS/HioevM4DWQRiQ2N
6QDHpQLO8ZbaKyEGNEL8y3mlsdMkVMowpymHvKk8JslSYT+JSHJk3GIrhI7rvfOgd/RBOGQoeepT
TT8/XRnWKhvbE1tLpUhsh9OOdjC0sugxVpbtevxX4tPg6HjRm18tyoMUB2xZOHd3pzQbAyXRmAea
prPXZ82vrICzNivG+ZLtO5TgLeN2mhLsCzma8vJ3/v0t9VL9ghnWENiBAy0IsGxRvHrVshTe7X4W
dgx6qIOjW8/LMcuNRNTiF7lu5csj0A1mMKjHvDKtyDV/MDCdJaSxiBL2bnzJW9isadeIoDNhOCwf
dJBBq+vU1HRVH7q7o0GELnk3v7O54n2CkGq5PSf2yDt5DSn9itnHA5v4zn4MsKzaj6+WFyqDwydj
DoSAbn1j2N0XgKVzUouH+I/j+YNq7qSrJeJBoGGW0/CID+/UZl4NcdqdcB5yKrg7vWc1CIdcF2+e
GqPgfakdX02zyypX1I39pD+Jr0BYheuMxjv1imrGpC11t3/ru6tgiXvdXQBFNVkapeSp/wrZYA43
ISPA5NBTadxF52nku8WluYbQ1SLb4hFkRaQeAm5alZ3xOeZy68j8RofOamIoFyYqVx1MxKJGCLM1
FNOwPqMqLgGbiTVMCoFrh09gZj4S6LZOOOmI/cIxzfb3zvVYF/HfxyK0ifqGD7jEv0QhisPL9kjU
mJf2taD9Z4+HW/EHqlQRKDAulABrrUBbIE4AwDZcEi/iiY+fSxJRfErzkns+Ihxj6HNILHgreuWZ
3Pa03pf/MZ2NlHiSkWII/KFd7KwWf/SkeVXUO63kUhL87tsRMim862HUymSX5RI3zMjbxM8MRwTc
0Hh/RD/qOsEXcWMmfr8gvHRt3DZSMjF8Snu2Ak38jM9nBElVheuREJV5ITNJ6F20wf+gcNvkut5G
Dy4+c62cWq/sBke2aHV+5WRw7MQ5MY9Raj1sSUhcR8RCdJLaJb1xP6j9sijNevmqc/G7zbKZjZMv
BfilPgxyWx2oN0WB9Tv2uLf/V8VNZxjdPT6KQ6F8ZpfzVmA8apezAXbx/Vvi5sHOyco4adoqfufd
X2hM5t87qKknuMf35mkm/jog9Ubes5AufLiuctc/Cic+C/3sPmIuvM2UHGDJOaUOzpzZ6EtbZWEk
TMiTZbBJPdJb8+CbCaazMOL2kAvINvVieco3YeKM4BvZu39beX6x0jLZgh7puDHI7JyMVjZAunuN
zPL3YQNRMXHz0eHfVuEFMLPNLMiopLZdBmBMxBXbKtV/XZjvWXNmtYK9d3DdBU8lTzgHZwsxADvJ
AoMma2pRNrLyVYI8malOFcx7H8jiMgHpGX2Lmw4Yrit1PBR426qvzRxCDrKOqD9G7Lckq2ohmNdD
GjOtkObfOZaHRCgv+crGB4sV+iEL1j1yxOvwGd6YNMNvJxzTSp8Mb4n+OtvA7pXjt7x3QM678mv1
2nAShw+vFSE87nvTzR6D68vK+IaQdlTWc9tZgiadRl0DpvJks+WaYYQx5NVHxgZ3e2dUuQVfLNVn
CFcxUckPnpWc7BJdFNQJfeGyI+d68VD5jDicT8Kv4crZVTkB1zzG7AmnCTqQLVWEvYSkJ1JNcs6C
zhtBuscUfCVLhk87NPLdUYusKLVEDHfkiexaDrsHvWSA+nRSYLlprI2wAccGfkp7VMJuhG1oO0H8
eYJACmGL6bYURuqgujpOcXc+ql5KWQCNsFtTlWgzg38QAt35E+6wRwF2DRd+P4x4ZJA2RRLfHmhL
RAIdiP3jBoa5cFXlST6PpPux7lTaaBh6HMyD6betf4Mq5zF9TA174NJWmZliP2fyQoph1tUOMH7y
t29ec0mgZ2az7zhjdaTuoKH4Zrz0WPESEWXVJ1TzWwStOAy/RVPgDcUxvpfZ7zS0I+sXFht3hPsy
a23Uf4FM/Sr+iclpg4BK3alk2TUYBLuWr9/H0GQA+64Q05kXAc0D8SDg7bu+xEbNV7cAoetUFmYV
DRASXqCV+IJ0Ut8z/yo1zmo4dnTKF9IXT+auGd6AtpFLAy8i9e+vzQaLCRMDPWyeQTzz9IDc3w3H
6Uk0YQh4mid/Oxx5iPIAHR7eNUgzK5XLQSHyTXAv4c4qyJ7A3ZtPjXt6iDTAunjg2Gwy+/9xu9H2
mYWfKAVLBj8f9FGpGsO8JIzSDeVNzweJC+z0LMaECD2Z27zKIFoVH1iPIqZ4goTMDc8wQXUQSRXa
8eZ8ELyWC19+HhyIRdTejLIyPRu+7wPLRZP9mIY9H6vN9Wvnbg5gCBaXEu01P+9oLg6kUZJr4NqE
fgleSpnK50/V6asKwROvqirFFfrQ+aAGOh5zrLIIhGtmun3zQLUEVB2b5h2Z5KEL0UKfgjgG3woQ
LVhOMMHSNKtwXzVJq8VGcp3bVpboZVcch/2yR1bZnm70XegrnkeA941bLOOnwR9oNUoEaxjI2R+Q
lfgE7JJ70KnxWBtU3JmovYRbtKtxziRKC162OJKncKsVdsHKP221oGPuKtXV6+2s7xaNun3CD0VS
hokXxnu/9HhvHtun4SW4ccspFMCYErD6kYg6Udm4TTalk65lHHjwkl/u4axFJpzfijYzBBdDXVQN
t3Pyinh6XuGzDuyQKMc6c6ryzifTjM2WD1mMzPVSYde3qeK4EvDEI0cQgsTZ/FRKbq9fcwi4EbCt
+UpI+W6hvqSA+DQyrdaHKKG11VGpY8aUAJbPdOV1VNhAN/3qDQiT+4VA7hjl/Pr1YzkUJq7D1G+n
OFC/SS8Kuu7mGyr+5jOauIgK3TaHjGaVNODbzqdB1wbhKj7TY2dfdukiubBaqL/ckWEyBqnrqk9V
/uRxeEjvhu84V4WYJsHfUgIwbJe9GNmkAf4rWdhsYbuTJzuAmWzHwGwcdAnbeNopJ9M0Bxj2U3so
PhUXV7q1Jx3wlbY9YCPFb447dhmvxU8+eenVmlqwAJ+dS60sbZQsHNdIyohF6AWpEYcve1+y0B73
8TR0bXx84DlNc4ZMaLCqYZm0rdFydVMzs2Vh7b9LDlLLWWTWux9YK/ZslNEVptlY0OyOMC66vvY5
+HpfC84iEssdDWxzTlm1R6iIVENrYy4frWNkUOSR3Aecjs6u5afrBklmebFK1gHj9Kvtmn21L92c
6wnKb1QcrEKaCVrPc2O6AKQt1npBwCGD21wvgyvR5EPVBhOZMv+8fACPHxOuObxHonMmIAA30BYX
QSO/yt6G3iMIN5nsMDAGPJoTOvpX9LCVjVL5ImIQL76Ui7lnpIY+daXZH/XdOjlAT7NV7N1uj5MP
8BXG4YQeV6mdJM5D+KMa//j4TLA/jSMEHPvlBjuJUnRXMYM2WDEmPCZucaxX23/2WZSq6bO9547K
Iq2wBGXbQPR0390GmeStSfmTN+o1LuuUqH8cmhLvCP1Fxw1Rw6aZ07JxYYYZrTuQtl16WU7FUFjX
gGfR9ZalKFyp7BwuLcxqFVjNb05GrMcny11zM/CpmhJO+Ttd0VlqGyq9DL0dtV3OALQdBrZURv/B
pSaUvkDZ6Ol6Ft8j2y2GNw1E+Z4+ZtFmW21Irdt59MHFwziqp+eWePcqjQzQ8+DoL0UjJmBPCv36
359KHfyEQyQKaIl7o/wwBMXAkAlYJnGb0TEph1rXNdweTNtJPiGqIsECEsxosHMrIsM5Ci0fv9vd
kNlEVUJClqZwMLfzT/587J64QOg/TD/b6vr8DNXnAzZXRT+tfpOzj2p2rXD5+UJwOm/i7AmTaGFF
P9MEMK7ZCdBZvBqVtJzPnf5Iq8m6JlSnby+fSX38TNjH+HQYZ3St0F+2yVieaUx6HOnW/+yKgEX6
wa+tPwlk2jNmzFH9LZhaB+JddlTbhNAd8pLEorkrBBz573zBXyhAWPzey73s3mSFhaHjvRVMYK7l
m6xTUWLcpRwMZsb9/axO5dEbauZcGtHb8zVde8UgjMsegVpyGVHrq+jEysidpKjT9sWdyEv4ijyn
Da3241MLR6OxEktGxfUPA6VC0pTnXdTAOB1Yidt0UyFZBTts1TrxS/NXpbi4UI5Z7pJ4Q6hetDsW
0yuf+tGvflz0InmzaSZEa/LKok//7g4kFhhpqW8LkRl9tmqEKYQbF+5l30sCmRD7V+5bKfLZeV1y
ohrWOQrBAK9TozqF1VjaL46IXe3ok2DpPb8uraZJQPvtHn3mxOK4aLtNHuc5hniUCvJlTa/j/i2V
DhYyf7b2mzuF1Ak8NjQbhBFos/K/dFSrcOSpWMW4k9wiLtXfE8rWSp4xJUMHW3ePNk9SuxRQ5PU7
voYbtGWzcqS5lj1QxMPsfSXyEuj96BD4ir2RYecVD7hm9zeZFnlz4xhqXg/Yh/mfbxhhIOZca78W
LQfaqv4uzVoJyLyNHbVIU9Vwo4FZ4jMhi17vPVLGLz6/2ANBzn8ognEKFgpN1JWGok5RPSV2f5Ac
O8EuM9IxJ3M7FF/6FLsENG3CtqU3ceKi0Z53SIqiXPZ+FuS4cxhFztGbLFJOnvpe8rOVeMp3PCOC
mSkTDy44ZpFViaM+4F/35GkH4e1BHyAynWX9q7LXRNCmzoa88YmBo6S8qPNyUjbPNu/jLmQ2azVL
eg0n+nMaZCiO3BMp+DfU/S53Q6j+0AFo7acU5SdlHsnbODPe/w6Zyy2Kltf4DhNX0IA1kUid7OF8
gTa03DeGc48PeBqnlmCF78gCUzARKQKDk3PF310utQqNy80z6n0E36tcgyicG7Yx6ONcygxW2Sl4
xYf4OBtEj80bJrU5pd64K5jVeGMhrcz8qw1N0sa4tFgxERCeTbHQKrDc4IkrNPbLI9yL+MAeqzoe
kMiQZLMxCuZv+mtZxBkxkDDy9Yoi/bGXCc88wph6KBHveayYpEhHVQlig+K9Pa7qS2kFyVzWsV5Y
P6v7Rq7NrZzGyys5JBc2IP2uH+wpY8cn1Wiqr6tqhFqDHqoeMAsK2WVHlPoqGyuZDoBWcpk/21Up
XMf1SEuJ0Omy5Z8n/kTtiqycyN/yhzY+zGcVWKkiByDYNnAFoDFFIUcgFUCdyFEfFoJTPxWV0C/G
jUGSuHGokGf0DelphMQzD6/R+UtcGsz/SWpPF7GLLOjUf/r0W+thMuuisxQU3240UzXn87TAiD8h
E7SVtHjRs9zDVDKIicoe/AiUZkkkXFYWMvfv2zc+cOjuj5tVDbnv12kOGJ77+EMRDSKd0upUbKju
e3Jdu1g1SA51LvO1SgNbeHcxgAGh8zw28/jmgFksZuQiKYZ/OUCOKcGvHnrtgBzrxEf7o7kYK9sG
xUXZ9brDqGxTDv0YRR0dCT3W+7aJkG5DNoV7gcNEUSLMo3660vNvef4jDvkzvGWpkXKMDU3xKKxm
EwmXahDd+ndjO1xuO0U3oPhrCaH2pIC7lrrbFgCffGPhgHzsZtd87ge8c5wCWDadp4udj00+uDVy
A1SMF06o750V4hof98SgRRhPlxxoEIc8R7o7GoTP0R/JP1lAwTdzrwLZmnIvwveSHnZ60wOePuy6
EeLFlcDBVRFoQBMDzOUAwNIIZSjo9G5DrRT4I/auHT/13Z9KTDseZaNliCWpYhmpoAVyY221OWFA
6KCwgOvTrEapSeAFvHasmmz31bvmOVXDGZXR5VpXjt/+uAOwYuee0cE8cMOmvIsASBznVFiEece8
HJ35IpoUFBW9fp2mdja/t5+gQhCdBG2cEggiGb7fQcasnRsO7ur2e6C2LEjSwFZJIbhfTngNgL+4
K1sdKk+vF3PBvvK5I13ShX4VEjONxi/weMOhBXQ8bA5XfOH0ADgwtk8/FliZuhxpDvu1zlBPdcE9
T7yVAa9IeSAEd+rv7SsOc/tKNgMw1T34NYvDLWN/zz70OHoeQuJTInCy4PMv9O98KMFM18q1Sglp
X7dJyjQQeT+DvwuET55F2QElkr/4mWFsodTfYdS0N4LZyTTlUB/fFb1U7gm8a9kzZoq6H4zMsCOK
1Mb80rvIYEDiQDyJqNVMb+ShEG85tPJuDFYs3Dxp5X12YdEuLpmKIO0u5IVy0l1tfc3L9TUhVTEB
yhxHDCc7Z8Nnw5rWBblP8mj4rqsMpMH3z5l58i/iobq2Im5paLS+3DByDha1CDLFTiyMEFlHIiFS
yfWZFdwZX4KY4AYpJkGQPZ69X6/P/OhYYdyt5mZ3woNTBO5hcQxzFLF9zfFIw3oqTJx6c7kUqXFG
3KeAvsDBWpahapR04jrRMWJg2goUc8ffpMkk8dSMMk7Czk5XwuxXddDY21xSGGE8ZVcrjmmvRXqZ
4udXjnNU+W0dvhc/rw8Bd8YU34JPSfXH0TUyNtI24QSg/psf7asAujnF4uL18t6Tc+0LTIDO5tdq
OAC5ga3HWv9CswmuQUmmV4Aks3nNvbrGRTObZIVquqK5yTv/DKWLkbdVY1j6AXtb38fV9jkAQ+ix
uKv6DTV+KBUojEl0DZ/2uj4O29oxWlOtGitKYPkiQxiJAOmYPwxFdwrlFYVZpeO5lHds4kC20zSm
epBWi7XoO182C8eihdQevTf2c317hiKd7/gqvfzsZrFl52SkeTSCO9NyCQKaOBBdXVSC48ZIEkAh
MyeS+B95vmAWy1D8PWjW2kQJ3lR3OMYOnyfU74fVXHCUnxTywhg6oPON+kNL087vcYtqetPLUvdL
zQTqxYm7K1eBPFrmJmhm17r0YMMJT3QhltC4PiPwSq4uH1hC1P5oflQV4b3+z3VWgNdIqKSRzg+b
Be/C+LQrL6h/QQrKrewD9YWVGEo/EGLFO42GKvadbHKB5rQc1rgvGK6RJ4efuQoaUe2cc2xIveXu
Ai83Q3+sTFG3P8qVaXGQkEAifdMgtEKdNM6K0eVvfXH4LRpOBrGOpd5DHC7S8jB1/xa7ORsUlv9d
o9r+pdzMEoNAZqj7XsT0rabzH3bWvAxXFr1gkGRZwCi7BUOS9RODWL53eu7+hoTvHXzTDZvwczDW
HaInn0gdZM/X0gpTQYM/X2bhlOXHtk4hWYdX/VtqCkI4MBTFud+9pqRA2KFFLKn5BRsCTB/QBiVT
3eHkcDlXrgGgGkyJ8LoAxA/K30fTRDzTl6phDJqkT/Bj2hO2y73HGI1F0EI9m6bCjc+uXijN9HcG
9Sy9lPvUe3PEF6bihgN2S5FwEBBY1Py6YXAfa0XST5PNlbREDLutM8vFrDu4HJGTdbA4LUf0b6p1
E+iJNjfA+JTIT2Uo/svTFDydzqe7itHoF/wcfA0QNC6xnCjZvB/TzNdaQdgxE0YYrepZ3iDz6sgS
BCmA/1+r554rk7oDigochV6fFiQ2Y58IMRLkXDDHxBG8V1XH3UDaBT0BMqnkGZlh9rk9b12hcpyM
ROwKdm1a1DAb2gN2UO2S0PJmpOyKQa4oRkztzAx0Squme12boVLl3F1Zh5nDKDQkKmmgs4jgQVcq
ksNY035+yAfQdrtcsE3G54mWf1Pmoa5HabxePwsd9puxJZBdRSr+SPQysJQC4+SCLi6wRZGRqd/V
q2YyXpbnwdKo8xRBL7zN6gbDPcNn5b6CDw6xVDe16xxLKsW078UoXHtxOS1CixCNU6zeGdKYXVBP
+aanHCTizCmV5SRzQNhG/gMuGqWtmpG5A+4CwBrJ3+GMMbN2DsMARhnEe2h+ArSeq5UArTiNtzsp
CV+f3PDS+cG4gxWiJVBBeS17ECvbHgU6aCq61cEnIVLWhtk2ZzgEZv/yMSIYfyb3kgC+wUBGR1cJ
V+1O7QcpOfhb31GBpKGkmbV0p7fHxlD5iyLdeztb1bqg0d0lrwJjT174+/YVdr5uQcsi/MF5O/sj
myiqKlup/5trwZObhb00iCHwBHr6wnnbUAq6jOvn6B20g4gjLyKGz8au1NgMf1j9fJT6lfvm8euK
b+CUcXPTgOewwZybyR7Hzcqq7D2snUaBAylmpGgD1qbPv5Wrmg3mkRHg5jKh8nfsTrS3w3djeXia
Ybp13/PawvZRaI9wAX+ddgkCmk+xq/uGN+7BRPgiAcHJB9YdE1qBqFfwkGvMrOP3FbjNaVPUxsFE
WFxzcrgiQ2k9oSVE5Q6usvyC6h5A2h0Q/ibvRQUrcLJNrPT1Z6n848b4xd9YzETx9qVXnGkCyu28
ppq7nqaYrynzHbw92Z6IlqcFyQBitTe/jDL3pyi4q5MbiXPxDZ0O6GtApmkZ22jhKSS8g0EoL86f
z+1hAONqEiX4kyzWxjEZi1yv0aJGuA+66v0vQIo9Z6EmAIrqzfif2odhABxAWMMXoy7OyMsIvCSf
x8YIKGVqpiNEakUb3qavs7qs7oIy6F3/i60E+ia6bNczd6za8Z2m3a6YiscxHk3dQRDVlrSQeiZI
TQuKeIyq+lmPwqGeBnyOhbUj7i8Oy3jgzlGZ24HkjM4RLiB6Ez9SBxxaXaRPFc64RyPHZ4A6vnen
j557KknA+/132Tt2hJ1vCp7yPPShMw8eQn1A8OfsI5TEZZtRladG6JRg+80tadmqV8JIYSsyFUdC
HXeHqbrmzkB8kVxuU21jsxtymzieUCx5oZuoYpU81qHAguNmjXir34jghuepz5zQhU9d/SOYBa3v
xIEMZRE+pwNYx1bK5+gKjfaCVxD48yWzeVvaQxaZYuGgnwpOYTAMPVHunykGmjpxWGTJI7kWn9Fg
8oNM7yKXcjkxd/3QdYNaI9WChwLOsU058wgVgPNVfab5IwPLRT12SMuwWM0bYIYSi3yhc2bZ+S3d
mp9kc9EnFrEvWtO+ByqUR3jQCzIH0mXxwFtR4+fBKnSbXISJHr39+ljNA40ISJoJGgSu/+o3/tLD
aeqdF9Vc5nOCEKxH1OqEMe0kgP2eCPyDxLi01XdlsfN8vWVaf98iWeXNfIJoYYPqwGJbbEQstYqF
xLy4B1t7fSxIOyKVheJjPiMWXuD4XhpWzhrdsG9aqRB/UGhREdtWEgPdpB/nDJdI5+rENul9LJT9
0NIvcc3+b9wGY/Cq8IVBtFynhd9CEnrOhbs58ir2tbKoSGrEyVttfAX5j42/yV2zyYGKIeCuSHPc
X/ZF5ZSjFgPaNQUoGWAVUNUn7qp6aPgDDSVIvpVYTwQbfGqSpufuoUn0aZudWt29qp3L3pNKfAfC
OJSTpOqZhGhPnLY+TQHc41nWhoBjnh2QUc0VvFimvwZa5lURj7q9dQ2PQGB3tb/OoLjOPgYbH6b3
I6CQ5ea89KvHpzP3YcOmF/vIKSUOzC0+NAFLDNsBv2H0NXQdn3Vj4AQPLJuKqsqkWVeHfpNQ5TCf
Ginu+6pESdRSit4vRaNejfDzZmN55Ysku2Z7C8ig8OCSJVxe9QynZwYd78TRgJ2DYIm4PMU8i/tO
jTnA56THeC8dLo0tYB1fmkURpC3qjfqVwzgXJaguHEWnT0yAdS6OBssuaeOeROe/l81yL+9bCz2C
boTAwXeL7O7cw1XIMBOROaFYrQnbLwWBxqClmRrHvthgQGDFzghQT/5irHXic3R2TfgrZ6khbFhw
1k0S2OrJ3f701XdjXMoE7FM6nmgF29Mu2/rsvAYFwwFfzn+VruPV3MRaphU3sXew86ow7Hs3T1mS
lrJK/xdsbq7WVyNbNCvdzIJjfz8WD5L5rOB7uskx80QviiYdyBy+7fM0u4LxMOuW/UebSfndLdQS
WSCSPAKIfYr47RNsIK/k6qnHeP2HyEZUxEAmQkmnNZM/ZPDab7SrPe0789vsOmrt94bTYUX1nCEz
iKKmzGhHBj1r9MOs835pdMqn2OgzNy1ygAFCKNlfcqzVsLwBRQ367LwOYHPfwiw+DPF4r9Sa7OVK
Gk1gF684WxDesaoyEwXOnRailJAWgrgEKcnu2MNeANg0rLULZ1G/R5qtcbvKYIfKtBBzZmPvayjY
GAgaBnl/4T1AguS2DeLkR0Gh2mDb0W+JiSCdDXcKPW6ke5nxvSNG6+sqsGSohjKSCG6UkRla6lTp
dhcEyZPX3qD3s9+I/EIPMbNclc9172oRlAoUiSCUUvuyt8Rxncf0mkBSP0GrzEpSjRYKxrpZHrPF
KgM6O4tZxqMe6fwF8Odv9gUKF3ikwWAENrFWUJkfAbqzSuesjVinXcv/iffklr/CwRRFGU6LX1Dd
tVjAR7QJKNV7WP7Oey94D+OWpa3BZuVbF30ZGfKIOKuwYyzaUGfXcdWdxhXHsU0xqZZlUUbEyPm+
z29gSD2R/4c3glMvyo/ay1jFZ84wrIbCiYQVG2RgjLfxG5MDpK5nbbHJyNsh2UVah1Db8mBbHyPe
w66KSn4w3NDO/E780RBXy4Vj7g9xmwwmGj7ANeoNDEp/Xfy4uSG960YaRrVtf3BdwEd0XSQN7dog
EEDpus5zV/DVAlrKdO3BTvS78ZJlMdIUe5o5qaRDuWb5InKGQ0M31Uv1ps029tYgrykWiKCtvDX5
I4Z2f81zm7uPnHPwf9LnRF5oYEziZcHW4QujPzBcH0VK2rON68sN3s1ySv1Ffag0Ig42GnSxxKk+
LFsZFcLL1K5tNMN2ZnaLqt4tt0dRGQQPDiI6XFxapFZ8rD7v/qcEyGbQutHhjCtZ1aV9Z1fZ2q9A
1j+ekOMfjCBRGd7mtoVvAps/oWvrqmdt8toc8fUk9TJP0ZHS3usYtaVC/jqlL4u9asV0yky5XqQq
SvX7k3T/w3Qp6bPYS4dSfn8zCW/X7e4qHOZIWERCpi/no/sB/x6+R6oN/2W2MHXKIANPUjIa4XW4
WCT1beXVe+tG8QD4v6kY8a7XHvXl1mBuj0Wi5/zagv714MfMfg2YZnwO1VcGuApTz+tAd2wrdvJY
LWHtRjxSSNvXTBFu+pQyYWEiXH3bdUGV0RX8UZbrMjxTHfJsd+GuE5HsvrMw1Qd0edjqwYWmCi7E
pnfpNYThXdE6sG+byByaigM6l04xVk4YGU3VQd0Kk1PKNf2qvCHE9i6tkxxulOSQlVXzee7aEnua
jFBCXhxBpoKBgul2gjUhwyMtwDz2G0LcFGMliXW3Alhjd+BmDD+CL7aR2Pyeq3MmSpYRneOzJhmS
p4l2yRoXF5LKdDTeZFlAxwd4CA09WvKDKDQ5cwB0Qyjh4gZyO4rlcWobDdoqmUHBCAz073NYsxlI
uTQS7LzqwvYmPi5JYfQD3JWw7CxqboHqe7G+tOPv+bBTd4uDKFMKCyfRwuYk0jAM5x0Me9IlqlUz
noQchSgPI0g5tjo5pIofpv+mhhQkzQW4kCBtj5YmBLxOZmB3B4gh3UaDPio7Qa5FMWsq8bI8gu7n
kD69cDhUg9BAho9rQIrjFteMaAUTDL8oGUHnUob4/dpmNqWIsrkWnly7NDk0etzGxqyX/2q/NENV
LyABr8bJLbSITR1MciGU2D+/078kX9TZUTIH090PsXaKCw84CRLFe0iZPNAift0RyMCsbqq7bWo3
XQEdzDvftJUKBC7lfoIs3lHwWfRTvHyZA1XRnlNnSuIAPspTiQuCJn+smBd7kXz21ykiJZMhAB6x
YiWtq58TPR0jLiH1oYqm7ER6D6I3RvvGM26yA9EeyBwOMtLlmYEc43rz4DRHhejNOg+6jyKeFN8n
60fAbYbRdTzYiSpj4KlZ8mC73FrgH8jcPMOpczbWB/X5fKOh249lVWPswuk/ycQexWeDw/Tz++83
SXn3QUDq9i7RMsLW4C96lRpEJU4YXzRA584l7ruFNMI7JxlLRg3Ey/sOAkRoy4tc4yWZ88r/rsn7
EfjKfTeFrG4LkqsX9/decUgtYLeIjaC8nCMJc6jX4aRuwhJ5yT0JOR37jSm10mR2bY9+bJhmhULW
zrAXZrOlOX4P3Hnxv1szdZd3QdpBzD930aeeCxBIdxe96t7HguGBEJU0GjwKetwIvdCszRpI02xa
/vG3V2OmWvxTaVTNSCf9BGmqrwBJSjTSXCNTbFk7rbVT9Xg67cUByImAFBlMUtaccK81/NFuNGJy
a3tBqOdkUrg0p0oia6w1KqbXxSiBRSZoq+GugEQ63HL0ioPn6TbtCuwTKBINolRyb8kaifmjvvia
ZUhSMphUouZd+yZJPOq9tMWeziKG5YZQglulO79cB3eCc2Ov1dQr5JJHDM87PzcQzEtoQcpPWLlr
BQFcJm/uNIUq18suVAZSUcyXpW5WVDha3Ux+hRm9zFT1rijRSHyoBEBziQnU7osiZtikQAbH1BIT
TAHVUthyAFmy7f/ZQoW/N8gTFAakALShvgEU4kBXYIRTo6hOGijO4p0DqWH2R1ylNQl7oV8VEbZz
ZDAkuX9BR9NYBVptKZeL/OsK0uMUmaU0ltbOCQXuQzNhcMYXDI1zLkKySFsvKjDLtYdFggu2PSTs
AwG5BYMgA3owy+apwWvAXtWvHlSVazWttuTx4oBhEbz7ON1lntefhVg4sCgjikPMDJJH9teibcHZ
SXlhIDjE2g7odNbRsJr2i+SNXjSmJoh/cC2IH9+OnJHf0qooYae2lsDj+2m/xFH/fC4+urjEhLVL
yLtf/in0YGhATWFfEwSToW0O5a7ZZXcf7c3wolDyEaq5kMl2REUTsGpcjH0lXBu5HDQ5uoX6+H9P
k4WwKKjGsXKBZs164I3KLOgVKvxogVt5o5CeioAkIdyPLJxzZ2hccBsJxRp8gaZ0YupaciY5n3M0
VYxKCyruazFNLoogHbGriUoMZ5QOW1pwhMGmiXp7U1eS8v2jfvcbC9ldh/EGc5yP71I71FkdiEGC
1Y0fd/rwipOFQxaDzuzTlE7tNaFhjAERQ+FDLzh2HZ2OvQzPMxB0qVz2ydigyss4nlZYa4fiedeI
4bHqAk+9GsWSkSKciejF1qiygMMb2MeCtsutyLhv73W1yEEehKYlHNxStDlzO3VCZvuSJLqm6Kdv
M8953COvhUzqe0UQnkkFuvbxPb1PWBLZoMmSd4/gqHgFF9l1wmbn1x1mfSIPK8h9cFFLPgOgoUQ6
r7IqKol0si47fUgHdO+93r1e5aoKb9I+NorCzAi1cWXREOcBu141to3lLVcN2gnEYerxojdvVMla
wFniHBTGJiIIbvvaR54FyOMLwm9RFA4StDLP+Law5+AgFWjWPDq0ScHd/S2vQ5XF0xe0O7/fw5yj
YNQJ9QvqJm7DfN5wHXhtDgHsU4Voo5nu6zKtzRNrw9lusutbLY6IMkLQ/6zjG584PmKsIrtciJ33
ivFkUw6QjdLXvadh+iEwMkKjkOiPrARaZTUyGhI71YxgJ3HWRa48XSWo6F+C+ZMVfCJYAywXP77v
7KjnFJIgHdeKlx9mv+WNRIc9XbnDHZc64QWz/EGSlhxZHTWNOTIqDtCWZAEgikZzmAM7Me841tVU
ZV56X7a+YqOFAKWs3dnQYmguEqZU36QTwHbvlCJ0qXYOWl8qWdX4sVR1zy3zZZr920lOHgArTL37
yMsEfaQzpeKDNKLAqqjmes2jxcAbG3aGuvROv31cOXhXmqNl6jC59ilKmlZmSuIQo19M+fkscMk6
U0DmHieQlXp7EjCysdThqYfvlS4DeDd1oaktdBYbCrPrQI/i9paPfB2rNz3rUqtlAMaidjEQDwX6
ccezQHOBpHlh0x3aCF89GK3L7MUzEPy7rAql+yu/57a8dqQ2CfK9aQ9t4nAFKFCtKEGh/7YbD5rv
PaDsk4WBMMzklRo6aPlXw7dDokuvP64W0jkxTNoQcJqO74XpnZ2xcMQ1OH3cgtxRFOI/Hvctnpmb
gBXZxsYWOUgHUu6rb/pXhQyCcp8rcXrf00pQplrtaaSerjy120SXDWHoquWKDLGIEyaqWWPWdgs1
3nQtFHnmmo7SiLfpRXB/FUVZfO/eTu3p3tFieQnUGb6d1C+/nB3ubmGeMqRt7iliY0sMNMYgAkKj
ZINwOAMhcbkQ+0hUbr9xrbiNJRJaLI9zDpifeeYeYRizjLuMm5sa8UsRAyTqriok62XFq3/sQi2h
jzQiKcWe7vm9vPL0IGbAmUg4qi5Ld9aHa4ZWh+mS1ReyLGubqhtyw560WTwKKITbkP92FEtIEF4X
OSjGFS2fT3DKOPeDtRo77E1eo1GlaKI/RrMy2HX67FNi/jj8MxbxRBtnvxHe0t6Mi2qUr05J8D91
RY999g04lndW+N46qpUcHePT8/xb3C5bYwgKT9xRBhKPvlIN3SFaysJNBMPVW8wYe6bjzMC157Bt
OgtHhNwIXDsPFgPq3UptFAapesQAOemnGuOMtqmeZfIC/iF3XvgidJXb4M8wpipF5jI/AjDWa0ew
BGIEa1D4z5YokVeIq2NaPLs8LHZYRPbzNx0zYpiXAwMghP7Tvl0v8ZI70dsebiUUtdQKkaCOIhpf
CQ0AX30IFp8wS1cFPBusKew95Gyx33NvxjnrhOKByJYwd5rkhnntC/QtdROlwgOXo8iVJLkQEybZ
4jKy1izuphQfbK45fJ3g6eQIlp+4aKwF9+FIaAbgDHZ/MRvoE4mcCT4v7LRjmPx2BerUgWZXVPmd
J0uloJSvUvOYv1wB3iKafLTvQuVTqWr/V1Ym+nd7NLSYU136l+gSkPY8RYvNK6RlAzAzkQ3UvV04
/zEuJ/kqnvGPfYTzKB/RF4psBseEzlvC3xVgq5OzJbTB5v1mXcmSfdG3WISkNQILjNfawhb9P/EJ
Q9niLTJJ8N7CUTLFb6b8IRNhLC32aTb2DpAEATEyOeN4HGMlzMnrpE1ToO/mHYTix4xKDgueh3iQ
hkXGUM/Rk+vV3omo1izRUPblRXKJai6JtyTMqeWxF+NNoa+mQGQ9/iWhO0ZaXtlZGzbCmoxdVcw2
Wugg5Ke/+EWJ2WjTXNoipkBa0NJ5PtXeZQQYXnMIt9jfq5u33/L4vSekdfSAPwrSQpw9A54LWrjn
IhplFh0q01YsepsHthFgknqaaZiC+pPat0j2qNqWdRrmOp7u+cUnNicdZLcQgZ3Hwy7+b6+FmRnb
JTG9XE7hwN5tW77FThbMthNol/BkMardWsLjsiB7iuZKFALv8u1VWAVQ0f1HKUH++6pw7h+5xxfX
k/OajPJwOi5ljqSCADhuOs7Cxw1Qfj4a2Fq1x7S0nPZU8LLMpVEY1rXXqy+YT55WX3Ies9Y2wLPY
YaE6D2h+yQTKwc4YyvNAQLkCuHfjPxBeWaWkgNvud7zkOj01g4++BgMhC1IgtjtUTAGPby8Q6m09
6sj85FGPqum5CY6BxLBUM2Ew8UQVz614AoEC+CoMBdHCVNhaIWaseXZfPGlw+iH4NU9WlnFd/VBS
CBAKuGTd46qnIfejQWw+36GD8cFC6nPVMv4k88qOFcTbsWLs9eyVF5zBewbP8eaO/WfFVcDDYgZX
CmTlG2VBVYuoFpZiqfh2lPyhpLmhLfQ6Tal0np4QuLaeDsS0tH8imG2QpXm7RJ06YO6is5k5TVQj
62yuNSMv8pAGYPflQ0lJIZjn3eBfx/DCCLqmSXAtm1ZqloSaIekipEn20/67aGd+dAZSREQCY7s/
YNdjtepLCjrj4DlQD9A7WYmFp/w86JNcmoE3M/oHcexZEcjO1QImKduEUadqqHZDK+2v5TONi+tl
AfC3udv0zWquGjcIEB7pWWSXAFtyY1xHG6heYXTPXTq4XVTbWtlSpeNmMkwrYOGD73eqyCHQjZmu
yGevAwU3xx7wNkxYtjW+0t8Gdfn0+IFW4g93LVWfNFJBPO1WIm49d/E4YIeqX7H3MsOAYHeKNzV6
zSKyTWiyPrsr/h3RDBvzg+h2TeL12ER0G8UIHJj4/QM9A4EnuzAQdaBkxeaCqPJ4xhhJxTkoFiWY
pmnjmFRge9LIue4gwbRa6onQmSA9j/gIvx0UsA1+0wAGW/E6y7uPkw7IPmTrhpFkNka393qPNrq4
GPtDvi06oql6k5lhsux84pouI29zWSD9X7XsIa2I/QdFmGcVViXJLhrPKS8Cgho9p5rOLqfodZla
CeYgSgTKUsbvclX1LoiS10emfAAx3GsjMMcgGEj0BURupJFqTPij+dC3CxQuAmu2zB4U4HC3jZMx
+MfQ6eOSf6FsvF1ZjSNXu4CpqI2q02K9lfyjCVYScMoqsgoKsIYBGjMbyv/3Jy5j/FrW0DuS7kPO
emqLkku6UeCc8O1uCuDQdaEw+89Btd8jm/FBIUYRlmYzzDJ8HzIUD66OKtYkibuxJsnx/laUWHo4
5XXNy+iCPSKq0firacw8YwHBjs55BB2w7bWYvWrJ0Jy2i5pr9DfzEKTd/f0ihQwnY7mAhAvFb2MB
eCWEmsSqVWYIqLO/kl5XpZdji9qyTM4b1f69SsunPQ6rahI8UBM6Lw2dZ58VxsT/1hrd3onp8a9X
nH0aOXGBM/Ds2xhZDUPIWBFgHfEl1JY8xI/pIVvgqpfuKZQlq0PpE+35Td4A5+UHZaQu1FCoLGed
tgRzEdINSMR8mqVoO1+tqVF+yiaAVkeA2YlJ4JQZKTumWhbVOJXXzwSdDRcqYsKGL1bEFT7mLIL+
7GE1BUtbuYt5VAu5EsBvOY3ykZfs/7sf8euLSE3cgtLYjvA1DolGMhCNa8KW3hLucGegvsX0HdV6
EjJLs+V6XfXbAf7QjLGCG63byphj+cOV19lqm3mvePznYlJYS2BhVuwZWP194bhRTu4XKjEnVpYe
AYqglh7wpn9re3Toz89mhydaFhTSf5Tp9M4rOdzPwGgTsisg5aNlD/hGxa+478Y37CKYpPzDPQkk
8hvJfoF9daMJvMmDli+6ReaK1oCcRTgDzdqUhBzGCAIl7yyaDgVF5NLdAPAQHRYZKAkXPKmMPhBX
MRuE8/YMkV3oaG4b+Pa+NjT50fZeu+ZF9jYSxcduDMi5CJxoUGPGSpK77DgbmNgS0bJ7TTPCp2vP
owdKtNcTUQWhBBDKLUkr5bNfuoitcHU74ep9qh5XPtZGZLNxxNVLjJrotS/3Bb1W2aeG4hvzio2t
ohYZOAHbhTvftcSy7MrXxcKeAyMKK9GQG2Q9a6TAYzLTMbwo2Vl86F5GpOUc0UGFURUdVO9iPxzs
d1fn0/XIHml6zcuGtIBxJYjWTWTqHHpuWhKM82giRt026+5tL9HHbyuxrWNh2zdk3V9ZNTzzicel
K50px8eIBO6y1KREbVMVeVGqihaWzXezrI7D3QooKNdD71A6JHGAX47FDSXl1XIMmCE3ntTTPN6E
gHYvqrGqRcrI9ibNfej3NLgqeyHcRAs5n67RdnehyUYhlUtYOZrEpf+peyejPAmrwmq8atQdcW0y
IPd7hPKKmH+g/H7btqdek+zWxt+C2e7TWYS1YRB7KvjIQ0z7SMg8aKfjcPx3pmif3r+kZPrspDbH
5Ug7NJjuDkF70jphVjG9Y06Z9qy+08yp2BVDYSdxU0ypU8RqiC+s8+eFr3yKXr8J6FFXZezgaOMD
m48iU9vrn1Dx/gT6qzEkvz5xhPsso0A5zefo6Es14g2C/u7GkPF4NOi+cVIr1Z1bJ3UTzGnA4nuq
FqYRrP+tXOmLJC1eA0TwVIBXsTgOuh41X2imXv3VjsEmrHgi91ecv4oDgNSymq/dM/jtzOTwWRDy
mC1xxOLOd9R5OmqxmnNZAgbkF6Ubx1rnEs5smvYzB+wSFxZQcxbxDgqkUUQwoaebMd4hGbBugH7M
uyiVdwfPT7TPentUSq10lvgaPu0paHwCu8pRsdjlUghl+DQEoCUFV5kLo2zcU74EzaXR/nPavaHg
ETYXGjYO83LluKhDbn5n2uRePyS1F90H0/uTGweCK9s+DuFe/opaIs0t2xQXJGHolErTakPfft0f
tUaebp0whXggBZ2hyxAh+kPOOo/PQOrS6idhdv/EQBc0zSgrVSXUlrevozgExkeLOQ/lsJ3Er/dz
qXDq4iBC+Z+gTpLACf0M3RmsBsnMwL++1M/SuF/k3zmFaGfnZr5CULVyrUDzPdbIeb9L6Uajkt9Y
J8OxX0zL9ZOysE7DqoOQV5UjtVytenBdugpjvB5upCemM4sy9HloeYz6U0+oPz/cWsv+5yH2sGwL
9eFCEjWPaD2iCNixdAVfjxd6r7xbKK6cYaqp9l1Oo/n+bU+N44c8M9Y0+KszoMYJRgAfoSLtJAhC
4FBGthotprCikBLVcRSlJYDHIejPGyjp27Mq/m7qo1r61X/tUsIxHetGt2CQkZ9xM0BROgKWQAUw
8QTiWDJxWBa5RY/uNSfcXwprbNVrqYDSrxEG8EDYvA/IW6+QeZXdteXyCTRAR3Dw8e4DD2SYJX4u
kgklFeMS81QwEqzvOu4bWCtBWbymE1TRYw10JK3rgpRIoDHtImLdPfy7ceDmNx0qkZrphX0g3514
XYzrGwJmaboGNv6I0bKFdhJYe8qAjZZzcMeUFdHWUPLjUxlQVSSgmkrjK577AWeYGeV9++Dfm/AS
NMqDq5r/rjVJbWm0ek+fBrM0FIhyO/5RChuDWljNh+gxFphtXe9secxr5HKVkguSSCr/QfQlITDd
XkFU0XbgGojQ9Gw1XAvSWH4KXeVchBd0mtQ9ExTN1O0IL27HWXC2hX8QMfamgUeikIJ0hbsniWlU
iMChf/DMm8KKKkEVkffs1JkuhraLGXGZvg0Qo0KkecxqNuIsdQ7wBnwrRcy9LYf9SYVaLGWQaZQ9
wr3FBxqFPaW2KXsjeLQWBCcx43I89TyzUlP88vBunX/2mWZJgGfG0ujLq+XP7j8iBKSKis7dGgve
JXhyeVerg2V26Ujt9Xa5LUyioHHsUSTc0rXEQ2xbE3+iOELqMSAXxaId3tYVNKiix3miJH0kth2z
azO+N30iQakzohjSj8WfAStKrg8/lbCHKaKr2Y+8vptdnQw2BNBgl2wClInLNzyGtsU+uotV4PQO
zH0LlwNMqE7d9+Ok6vUfeNImUzACpU7H/3imwGYuz36Zyf1J7Lf8FD62OOa6okCBOjojzVASAB/B
J//UR3QrKNo48+Ilwu6GJrQp2bv2tz6hI7HcMYde/OCCfNlakvfq2MIfvUxO99gSh7Ne+upCSh/J
jXR1Bb+cSUJuX+KG7EWKLSqHJ+HEmSt/CwilPqjmeWemcQAGWxlOIbnMv/IgzKmlLXgOEIZO7cmL
9doHpfca8tS5thi9DiJLSLY3YXZqXKmCmW4cAYII4kSP2ReNPekR/bYv83ljtStYx6bynrY5gwIw
YzVHO/CM5x8bTclfgRjTIxnyOh2uXRByiyCk3h+PZoHQz/MI5ub2yynUQO6kdkCpdQbRB9cDfIYD
jOYt9xR9uYJHuWbLHpGk4EEO0xo5MPW6IUubeSOUJXQgd9P4M1xyV640BKfFB4x6JUT7AQy9O8ae
Z2SsFmkD2nyNRZgNUzS/5Ezdlxzm9agMjGO50F7CRfhNTWv8Rt+i2nKh3R7SFLdIogBGAVPM/GTR
NAlGNXxNIpMyT9T9uuu8dl06pSpyI5qNTIbWXqRdoHRglTdHkyZQ7ZRQmlLaF/8UTklvG9ay7SXa
8Pt+ntZJDtPsSS1W7Yjw2WpPo9u67y2ewSLP9tseJ+KC+jRAcKOn0m4bUDvxDRyVKtqJHzeZPJVb
f+TACGTvEvMkCp3ErkBEUuqUWmRawUXUH6UV3MUilqiw28HaP5E1biS4sX/ONgNGTfjIQkvaNKwK
IP/N8mvZS0H5PstgsH6Hpizdy1DyUKiHeb+NE3sduERrHLo/MT5+l2dORSlzuS0qHVKvNijH+hN2
BcME23elEnYEdYPaGqNLyOFTGPoyhXlOt1nOLB38M0Wy8dAtE+pyESEfrqge3j88vyyHDQJrQlBa
IzEB8RNW3DYL6O7L5DhOsYfFR2bWff4i/XFLUWPRPgIuG5NREEPQEEkQpWzXAnOzumA2xv80PD9C
xDl15nEyfGlxOxTMDbdIr+Zo4FYwsWsvADPeQAu7NZXmwuXV+299cPyEwdz505kSriIR9kEEqpMY
J2YzQLFQA/V9l2AKcmc8E0iN0gehwc2BbRAu51/FD64TraoDFePrpfl/KS8iWVn4uM1TV73Lgp+5
EGCRsZwm7fehHzO3jGc8HLRtfqvbN/2lJ+/+Vm2ynO+L3ka/F5rYIi4AZ7zmZygMyDUPTpoFzhEm
wQkXANe/M3L7TUznVThLlaCbfN7sXO/co2BySut4XXnv2B/feLLPGkhGmNS3qLm7Fnv+WhPFajwM
X1i9S6UEiaM9ETetL9InFigEUxwhRPmc/DIEq/X7qxsemIZdjm/P0rd6ZaNQV+Uxvx5DAbRJKAnJ
cF8QhFg1MJWq+d41OeHM2gzLTyNjxygJkwtedv5sXdvnBmOcjQMPTcyHSQFUs5C5GhThgio2r4H7
uVaoUqYMOU4ilFVnRJpDKVg6ZGtKFUs14XtbLltmpkpFeREd9i+dGN+udYyu0ksmssT0knb5949E
1VLMKmXGNbn4YfG41CREtkGdM1q8FXcVeCC6RItS7mWvX2iwUrbO7Ix+UzEzLD4QH2d5TTjSFwBc
23O0F/cm6X2u6jsIyefDx6FuEClO3Tg2pJAY6cIzSve3b3KJyhRYRmR9/wER/pVMcyNi0brbZwYF
vdr3TjQl1wn8ZMItz7ia4OZSv9nGNQQBbRQNJyP2qOfgZdQlqC4fNWQAAsxXqRX0NNagxXZuNfez
0YqmQtiR+v6D/w0lLOK42brUVW+TQFYsfW04bjwKwRZWjtxWybAQJujc4wkqV3Z3o8K0+MB0vBD2
sZgHpIWb2I7EAYwUD2Rbv9sC6DL9sm02b/kkA2ccej91zbmQhpFEPDMY5G87xXITAiWIooSh4nkf
s4MzcYeV6k5exrP/MLhjY8h2I4fbBEW6VUbJ1tzX7YFK0mHqT+ZA7HWn9vPzpNwozd7X/Ul3NCr0
nw1epSeYQRXYjCkUIeXIpCqT4a9mUV1Y6so/QiBCj6oYyE1u4ZSYLpBW5N1bCu3OpFefLeQwDxRW
HOaenDhfGLK1VPWfCap7I0iJwHvIqOLbu/EYStvgumU5faIfz3UNn86bQJW4CV7WzFA8AAUbnzVx
U/y+lm5L5G8EfQdhvPZxZH9FJUn+wo4J7zMUofsMM6qiM+1HtXVXggksMxCeHLudC/QBRupmFa4N
E7GpSLOTco8/5RD9yYroFCq+zw/efNI7xzcgWc5G5bQaGIB6EC41iRCVSnE4Tg4CF7iIcP9ky1QJ
uQtu8EPkxWL3NNzK/OMqSMc8r66ILhghAEEwuW5cXdb0Xw0Ku4SspivRg5bVDS1U5wd1lKzHrN8u
gKC6Djn4sdqmvKAUy1L0mm2W3unsO76ww55dRF8JlZtytummdj3Gu/IOruufhy4JqDmnVbsAlEbI
rntA/0gxZFQOF24VlOibLLQEQjXuXmDZGtYg9qh0ZF5sGSNdaeM3vTEgzx5hk0Biv5pvG5CCgE36
AhVBlYyVPMrsKyoALBsi9yQ0zne6TJJ5gWobF0+EWqax6FFVPHe55OXHaBt1dGSgvBy/cOdbzxfu
CIHssg79OQ0IDzJZI5MQCZw546vC120YXaDKGavliapYb8aJ6+RKTHnWG9F07JBvoSrEUpVC0Y+5
41Ct2lIqG9Vm6xDZnc+sTArPbaGmyCyr7Y5/vKVFTrCqg7euHDkkaDxiCoLQ5uHFmnAGxMezg+w2
n3Yh/5DkjtR5kfav6j9B5/vDXrLaktxdMQRXjpYePv2yB2F3tyRH5Frsc0QhdJfd78nd9J7+NZY7
r9F49wtX5F3XpXpjFgBv7n3qRrWPW6wzg+zILApQdPN/s0swcXuCk6vjD7ROYkbAWz0ClToYuI+g
NBQYF/+01p7NIax1MU0s+tWiHDw7DxsFuOxrrMivpiXOAZk15deU5zc4KAIxUK0EDQsEiYgHCkYo
dquJkjwUzjpIxan9PqMqoinKdFhHM9kU9XSN7wrI5eH3wPEg9J5kzC4L8E8toogFoO8KsiCbBYUE
Ixt4X95BN4bZxVwQ1bqC5KJ7EMdH1sH3I1m05TvOZ66PMNK6wSV9eiL6X5S0fkJDKOtDNf5ouaXK
mdom00kZ4NCY8xXoFMYXmJ0RmzENO/bvMEMg/QbhHyOu3V0NNsVz/lcLmmRp+5V4a9HTzIW4moVY
1Y1UrgF5lpwFJh8qXEETBtMoyXa7zqas1Phhs7N2BtlAiSeBDxg1ZF6eFtHbIkD/FXlM2V64lUqb
yzJzWIp4lrWVu9rf8RfdHBZaaWpdphBOsQ1ove0GheuN4DFfS3+FVpGADFRJtJkMWCE/tNC+Hy2+
mP3TnoQjR0GXAYo/vuSZRddRMVhnk0HieR+zSBJVzCj9uPULYb73XPNij1/ETEmMO7tihbM5FAM8
kdAyLsnF6E8RTdTRPDyxFru34aUQhiD6VsxBgzrlbJM4xfBxinlfD9z/CyfzZUhuG26VTsSI2z4/
Ag5Dl+mvMGpyFdO7v08mJhepWC44OQuv+h2hriNYIrrpmE9XfGELIiQ9Y8Q2Ea6PLoRaENs//QtP
kQvJePNwiwbINW2GYo2ir84dWUcXw9weqpswlykOhMKegyiV9+0Z8NLNQm37QmXtjA7iKHARQorR
3Hh0+DrbK68UsQZdm5ndqwpZiu9S+S8JpPDi3a6VQk+GekOT1zTihPgDbVdl8svrv2gzSH6pZgW2
Ynf7sSFKAG9tCRrsH5ptvHKG3CGqMgOTI4rLFwrs6BQUmnNMkmKGteLNDEzqNX2qqUt3azh4Mj2W
iC0O+2b39hOmtMvBOAHphhWkOZhUUDtmJlg9u7ApJ2dtfne8S9h/MKQb9ovCjdwD9Cym3x7CSa5G
w1fsjsqxD3+Plz2zu2to1SGxvT/qvoE9XYfenLVz1/Eqlhu1b9VcNT/uNCi0hCg1RijSPuKMYQ3R
ADmPkHi2Ek4nlpjTfLtXqb+vEYVp38sjZR4YWx7WMLCc3tzZk72buCOeIioTiIT84aY1uYrbt03w
axhakgtbnx8vVawfGGDHsOSW3DwDpYkU4/RkCCqZBJ4mjrFPKf8GEdKDQkzIewn3iIwWggNCBsXZ
jyOUpSwefg3Sirt59+UGhXjosod+3L26CyknR93EduoBWP5Mcc+nIDtYE6dl3kqp7NcR871IXsCi
0ZRV2oCFSPufAL+GxkApRAR8Unhn0mATqfK/PfLHTL/EPdR2SzEGMV7aZ4fxHzCGfoI2oj2Lz8BS
R1j+VwWEJK/E83K/MH05dCV0TegW950WO/4E0TC+fQefPViUh5P23B4UTa3q/R1y+O8Vyk0x6tnz
HBTmZLy0AxBQhkJIUlVNRG4ZvatNXwMT20PvhJBCmooL34imVMJtMeUFohbFGepUQ804N0o1lPkc
ifdKlaB5DUS0fbFsAmQ3ruU4z+/7cl/NON/FQgHSFPqj7f1N9Pu/aMvSIVGsSKqL6kxBEmEMMdsX
C9nktE6ZwHd3kd/a5WIThIFMiLpDAn82DrGie1/6Ui2VgIhmpAW93cwGQQAwrsC83DIYcYd7Sl3h
9MrBUMUuHXqS5qLFlKuXMhKd6JDlK+n3vR0cS1/h2B2eLfLGBQZkwjf/Z4CgoPb8dvn/WuKFzzwD
GvIjAFHb2uIY3EbRPTIV/PBeO7rjLF6cqGKp5lkyALz3lC6OPVXy76zFz/J13Wnke9BuuNUr3ij8
9nYlPMSwgF8UVTNeA+ZX8oXC4SS91Hzr44hx0xheK0o+xCsCxa6e3TeNvTLn/s6Dy0GmVlzSjPGA
UqFIBRnDCAvRrZj1rkBYUH2ZDXuujvi6/96kmNS1yE8HjPDyvPOnpjmXR4Sx8VlpmZ8ke34g+sCS
J/6vYaQAwuxzWi5bdiJVYSV+cpLdHSvv3QuaRxXvTe9XxVB5h9f4zljrDS54h98vPHVFmBRNPMSb
phqLBLgVAk7YuFoiiHKG4hcb3526p49UswQZWz/x6zo6TkOKf9viQLCtVXTGdJordIfib+p/8a/U
XaFlq4Qr5VSPeg5vz8Z8P/zJX1hXJ+MaSbYjqTt8mPkJycj6uiI8n/iHkdmlUDKZpzs2YvbA7F4d
BTOslDJRKFbgshytyxWV3xutxHN+YkuxcrfOdNq+Q7O1ils09PDA8Ry9i35oZofLmWVh/+TJBZg+
eKSOtYEhoiAW+aTte0MitOw+gPUj1l6BCqJRmePYLnQtv/xcvqiQ+BQCr8C+cV6DktnIlO/13cQs
htxVTt/4mdRi8qStVakxiCSmdxLGfxJDlZdBBXtonaqi1w9PBJsjYI1Af0pLjT9pXNgOpwTu98oF
FLfJx3F4iZ2eJ5BupMeCynOMHPVndKjipYE3O91IsDUmH1pZI/v7JlLC+SjF7NoappspLLMC9MMP
Xv7Df/72B80oQTqRZDE/gWqNu8monl1TeIPlzKm4Z4pU/gv5c8jQW7wQWkArLMf9FIV20N3tS24p
d/9eddwx9odr6horlHrr5gXU0QyaUDNqsbNrZVoCsBzBTyLO3kQgVTHSAwAO2x9/VyUj9Fo4X2jX
XhfwRrMmVTJO5X7NoX42KWMNaqqhyT9nHgTP7R1uuvct4ITRYeWJhkqn95qKsqTcFVW8ZTat9AY6
yZsm/4jmlRz3ASmXVxXSObcn+cupKq+NWxidDZXBO+fP9kk56RBcgTYLXSSalA+O5YBbAarzHJIg
WYWelq4O4D22ee68y7v7GBv0HqnaPUrO3X3/VK/FHL465QFS3lkm5pZMQOKJMhZWQUU2n2scgR2N
sKe0YaQGZQjhUKiZ5C2Z4YP6stlYUuGyZISl5egYebEQI+u6JU9Uhk2RZKEwlGtIW9G0GVpYjpS5
PRx1u00PBDw/b1iCTjjqRsLBcUoFTZFPABfFIoM8jg1n5zejLFHjelMoCJbGFUQprtN7B30+lN/H
MMAuZznPKHTLIBTqFoFUbXxP+mYp2Y0YIRtYk49b++kTaD75JrXCtgx641SRZ8eeSOq8uV/WOco2
mOk4etWaSGy755z321Iw0cZaA/mH4tZQwPfk/qOkkWkd5SPr3C7uGinpkuIq4zoxSXQuGoYJ9Y3q
VAr+F6m6h2w/wyM4eCHSf2VkJ0c6iSFK5L/bUi4zd9wtmakoiKTQukcHy7Hbo7fG2Cei1IIvPFFs
YPSbzAUXiWrIDbBHcv17N/ERnhMQhPkJMxH7o51q5YAjcQJ2vY4/zgFnlF3p7XAwe1W5fzp29Vz6
H3asrD8l9+3kW356uDEz5I7H6A5b8DyxIGWgbgJY7m68afIrrD447dFNwNExfLWgXmsy1fe2oLNP
/j2HzVTp6x6DdVhP33n3OLQ+1GzW7qt50qboHAgdCVEpi/aAi4XMHEiVkFbMbA63I+Cd0cgbMpSe
30E2GH6DidPY8nXQxo5wMmg3KXs8/pNgvjWmnObst5pg4zBEfvYltUjRBmdZ9Rb45Z9sxO34031v
9BYJ6fyN8VNO4aywp7ZkPIhded3BsZ8r/pkRFU0QBDAAEVCUv+D0IGC5sWPW66Q1Y/s2kQhPKeIb
LUsjUY/C7D9WgShSIt9C+24lJoFyqSBQhps63g6M+6O5QXTsXDRQg4RB2A3pI/bBlPAKgTUzTvzu
23zbClc2XTklSJU1Q/hBeDmrlGcRP8R9bejCPo9JHQ4/D4xLM75RQBVl+prDx+/6exOsfQYFfKQz
So+QvJp1fgB6POVensfzTa35dCmnL9qPqgaypAhlWSgujO/MxAn10qHpDay1P6+lZtfIY5MgY6a3
2ynv/Wf23xiIfyhuTzqcNEaJMcrU3DrIGhrtLzdNr3vyygU/FCVIvEK16hRDyA1W9uhoeJ4MmH8P
R+y6TONSkei3kOJFJLT3By/AD0wYSI1GHZ5iyrEQ/3/L9CC+Cu76JbNkNopzdp9/izeQbC+fjzWQ
X0NHwxD0GzGZ9lKw9EM/J07KbyRolOe7JLnx62QNyZJRfvVxY/jrbaawRYugGIWKMceDH4mpBvrb
A+kXjfjECGfPA62MX819zAqwsW5cdPWO37mlXAu7d+Sy1dM8/+AEYNTiGBLuNU2KJ4zjEFfflRGn
p/aVXBoyJ12cSYRkX23a+uoJ3YJEOlPBEYc6lKJiGLr27b2BCh9c43er9HPeeg8S8DKap1EfV57v
PmPwWkGCZkO6TZrqkUpUBIDJqNCGcvkjp76f03gTWhmrFNQImC6bh6CrrUEZPxOeDM/CnsFQxWfp
Xmd7xhtHmh3p7+0YIPDnic/HJ4leofm1ieWD0u67PTKgTkX1sjgWSfDtcnd7S9mr0TEj2IxeAF/f
GcgTiL40+YlxK6z/ecB/vTl2l/MErOLmnBOZCeK3vhn3yK2LhTwBjksBg5VFmbFS3jfxEEUKSBHo
m5ZcxsLotdcGaVOG8lfu2DCFXFZ1EasUVvht/FxBtZR5rhS0Cnda0thHD/ec/ncLc9VU7QUNFp3D
d0A+QzgKuGlrxIXi3M30qQ0fENqxRGETuYWzS0kbTn1AlR8svfw0I6lRhlRpvwX8ydh8aXMY/Gs1
v3BtDLggLqXWi+0Xc4MLZv0+J98VxaBJeZomz7T4uSITeCO9SgmaxVyQonm6m+n2p7C4rYGPCiaZ
7ZO9rkkVOPWLQf0XCXSneAzY3HlIOexPHfEzH9GoFWOz/nN74jFBhfBox8YKvHvisJGyXtpfQJiZ
KudCc5XRqL0ukvsZ0lKE4ZR83nZdEvi2a2/PHhFFRtMbvbJARGeKWOIHg5nJTfrQFb8viUi4BlC3
O8YDd7/cIH5g0r0bHKBy12nhpy0Ef5wXD9pkwAZFfTVvT3yybc+0//E8nBVBUFceb0PYKO/7LuXQ
Nsijcu3I+/Bl4LhmIOWgGg/fIXv7dfMm9LFmGcZW+j/Z9kquvwrya6bM523my0sv2bS/cAS2gH2T
Yr3UJl7UtVTvXBy+JbXZpBfeOSeU4Xi0pC3GoxCumKjNBeyCSaLB3ASsiXMUyKAlr325cFruUk0P
CavPV549BX2CPDEbdxTb9SOzlfwtPKiD1kLTC7qLGOmusE512wSd4ahXEjQVy/WHIo04BV4xF3CF
ARF+jYaRiyDcn4OTcTGtyoqPVqEIISqRfr/IWIutQ7vOxOgrZgdnmvCqDt2GosvA9HQaW5rXm/pP
NBjsKm6v0UDZfHf8xP2CZXG3Hs69EV9bMlk045pEY5LfrIeJTV+JjUHOr84PDUAQGjjqWmGYYBG5
AiCQAbuZzmgo+fKS1J3xPjmburUOB8As5lvtpZYlAm4Q1JOZEDdi///TmsD/qOTW9rtZsf2ZH5Xc
scgZWzyrNCT/Flf0hRE56Ht8kbGaKN1Zwqgo27ffZpgVQyau19lOITXwbQEmmtvMmyYU8IjIWvyb
ZDJjJ29XGST9oBZczbdhgtiVejm5WJQVTha+Q+imZY//7cl21B6p0PrGL3eYi6Afp7K06bnICmYB
uv6e9cwjwrc6NsZ6VAJtTpErxnoZkE91KyBWKdUy0/zpe8kzGAyU29Ril4dc0tXe2QIzdyYpKl73
jdnmVb0Jp5aQf4aIK1LLCYMAHfHySizuipgu9wRg9w8VkmIE0BUJ1arZnKM8/ed3PAqucEqtbTqJ
uL8N1VyQ/cRFdS2/rU71PHYtHka+xpsw/5bxOE47Zx+99Y86bxsw5gq7emP045/k1R2MvUzdTGRH
VH8jaYRDdG1OR3UJc74uhy5Q1PKDFwtXc4B/5KYmvWJifsu005lRkWa+8wSuWj+Tpm8BIKlq5bPq
w53CAmFLPWYdkuVG+ur9hZSECjeIwekV1+QGz/hqFVNY9jNED3e0t4bLv7pNZdjIcBL+7R8Va8AI
mRY9PIlzH0BeW0K9cCMcPRzLjv1qJRcktCLW8HpmqiPSTP+S+5vSMaJ70oj0UAaXAw5vxdzbN5Qc
JySddm10kmCmCBFOf5qs/Dlnss5pafcAJGDFGTTZs4VXzp/5FF9RLQIMM017uwnT18UzFFiCpl16
Bq+2/LNC6PzL9XzCNHj257HWZAG9Kab0A3vg8azmqpi9302Zja/HGdMBFGA8V7kvUDcnZpurmW3o
Aj5RE2Hd4mswz9HkqLe7ReczKjXOOsEBRhEDNmu5BNeA66mcw0kgJiFedb8Ut6+tPogVgye5oeF2
80TOyss4vQ0+R4fuG18tDiDNcfX9TaMRxniQ9RwRx+aSBo4oeDmBydyqTGFlb4br7851IEeWzsWB
mh68FaDh50teRx6bcmGzDlbGLcCkYpdWjcmSRYO5ToTkodaSmZ17Uu4BPLZjI2ZZ37iyeV47gRWd
vJdTkxYpq833NqqoJc9SSItKTBeFpyJ4Wc5/2BX3R8ZpJh6OwLCDbHbKuM/kcOkAVtWbAUVDmxx0
1aqJJzomQl9v6SpgLYgOwO6+5PAHDWL+0++m/7Z0HDM7RflLt0MJBIyQTm1aP2Da5j0+37FsNqAH
yZYkPZ6fhNUj+ohPXSB71TpXpVQB6xqk4mZ0Nf+/VadXgZL1hIfKw2qfiQed7hRX5iuATqGe5QBR
9YxnxeWbmEfFG5higTBhg0euHfmRN29s4Wd3BjlzHkdtDGkJVwUFCQQkyNXcOlLg7WadSVz7P+WR
CbGXPsSMg9Enn55ols2kzEHbJiRFtyqWCXk7yKz+zqjqJNVjrb2TjoSBNfYutkRcuk4XUw4EKgot
v56UizYD6T3BjGytdvKKEfdxLdA8EAuX3aC7IajMzB5Sb2kkH4pJeV45UDOmjirE8Qa2j3kuQodk
dl7AOdpPWrTVqQu2WF9dcij/E0XmJX6nmAWXjf6VvnA1undQekHRXWmp4NhYKc/4OIdjs9OqZ6bQ
PvISvbhuWOb4qSXzg62kZ6udx5WXxv0EiWzVrOTXKyYWtukvcRNKsCOXzyUYMv1kCt3QOpn0jlPs
GVyCBxrVnovhTJKgaOGWfg/edzZSpJ9dcYgQ3bQBjaXAE9z+eHFFXdLth5rUgQeyj6RqUHwAKrQj
2hk9f9p+lC8sNhhvNwAozJ0GjAumJef3Z4W3I/5neyx+4JTHbmXy/f8wm9Ih4o8rRYGy9gcBwFVh
4cAIxrx2JkUKbfSBAQ1n+EKBU7bTohibRjt06aGyNizoi0crQAbG1906Q2HDtLJF/2TXGmXOijLm
TraYTkw3UQP4ak4D5fLDDhr0aAvSyytd7WmBUA5v4OSd+XsMu28kdDcfiTZzYMiOQb3WfJA9eo1x
geFcYSz4jo6ChyYKSeqfjYUqO/EAvB7CB3MEygZaaFUPmyONWjKBaruwnMvxrfLvZ2HrUuzud9Zv
naRmpyDyiaFZ4ptUGbniZl4fs43fRD1OHB3SLU+9i1lMx81bklS6BE3crvLNKwE5Nnc5qi8QC7TJ
wPgVqPl5spbqup7qoKhMm1HmFs4p8w9ENPLWU2VdBYcCAjmy5fohcaFcNW5T91q9PGYNU+Rb3cRZ
rKcodT9OhcNuNhRp2HyMIsYteU1afA/zLJq/pQlMFYpR5lb/SFC6EO+VmjbgjMiBvXbpdHx/vfxN
Zk86LLYRLXXZCnWPU+nsAAGfWPcTi/6FM+1eVgxW6Dy1CfmS6+zvT5U+1K5+KwukzUJt8KsmDNiD
yWi3kyWhruj2qDlOkP3/T+u/ITYlbCcnzetwbTWgSNbKmwk5WALQfQx+65XhjAGuHveA1NVXynBU
YNWc96UvJh0wtmoOVJYFg2R/vowxNd1nJP59NrIme19zIaWhoNHIH5YNNrGV0Xn5uVP9npohHUVi
EA/5KrcmrdxYcktIsykxsrwIR6f3FaaKmjj4Fsz+3Oz8qAVY87JeBNtwg3VZn6zSHG/F9h1Hty6b
AwRw1Ra/7jrVMCR4GDVj2KGmbjwtk+ImJivo1klymjN9TEiBgdYxpW5EVWZoq64+V4HmFY7sgJa7
nqAsgN65hIdyHLOomU5NYdGnuIQjWFIfWnNhRgptrqjUd4pgcu9wCpI2myf94Jntj1T02yJVa+Ub
2Fa8CAhUza8UHjulWjNMy0vqbW3Zn9LYpBx2hyrsbAIw2Uu9SB6DQRtA5KPOsvMEXXLlGkI3I4xq
yGsIypxlgeZVa414Sy5ZzLvidhiln3nhwJVoBaw9sT2dDql3jX5PLW8dw8LfzV0Ct4JIEvqb3x10
N15HrFXqUbVOqUakF0fciXwyQz2Gbx3MgdM/wKFBerdtwDPP2/H/nbCUIl6cvZqNRU35Q6g0RIDo
QF3GHuwIPyQml2OW9ynNmwXYZ3634tFLzSHry6mNK5IHIZI5r8aljI5PVdf/rY3X4hvBbIJlh8CK
2BorxI5aUhpBy4io3VMG9vbQtLRRaMrBvkyxQnEEk0ExISHAuPpoAT9JAnP11LxI8fkY1jlAG1lZ
HQewV/xxnb5wOeLd6kJP0YqBUso94CpYHveyA4oD3w64p44jSYYwFMv0Dx+J9zEXjClo9w2cXbCs
sGZpnZG1vChv+BY48F7ePKwpdOeyFiyprhs14lbwATpQowvbNBwqq7iZZ6bjBTGx9Qy3gyoZ7CeA
i5fIefFSq8slrKQwerHWZxRvbpQcF0sCyBKUczKHanw3Gw9zdIj4jrOkkFQ7v7GBTISwSlU/o6mY
bLz4jDwGyI39yRRL5OV/vFIuTPsyaX+xnTckE82dTX6BxlLS2uLtWS0q42i02VYsChP8DLQbMe0u
oOncXFG25hkZsaK5EMraPphLKw3nNHd3ycdj0ipmVB/ci835f1d9qmctpLAxIIDJ5dDadwkoXWCF
FhTqsuYFrkoh0kCdAuHD+VaUlcEAjM8SYjYKkD02IVAFIvkbH3NzdYx9qdSiz8HvXiV1QrBOJuEg
zeeMz/dDwsDPJ01BfFdZgSeNcKbXCgcyZjQfrM/ZYltOiFLaJz/GhxfRnNo6njqSJkG+/Df2CctN
dwfCwUdTRuFJw9KQw72Dl5Rxtl3k9mYkEaGo0K31DBeA1YQv/IStp4QTg84ZYQARPFo+8Ss3+Ih3
svA64m5bl3tDCUdDLfX3BbzKI9rXIW6G9mF+ut+Id38yCAwo3hP2UHbiA7MbppBVBb12RrkRhO+I
AmJyYa2PV3rmohvwNhYM3P2mSFXP35qRYGsmYK+JFOyNMfSuhgRulElKy898bOd7tRRkP8KnY2fu
Yv9ndBMon2JQm1R5qZx1lE7uOfnkRM5O8Y5/pLQHYLEk34P80zjcP4t+aUebdTh1YvkLo7jLgw7L
pCj9Z8I3BuyJNeCFGmqOx/JiZCjvQn+ECI6QK/NTyo/FHS4/zLmW6nMWBmHbY0IdtRzT0AJoVMEN
ySdKj+vSOP++evqVkTB2Xlyd+F5yeXG/mK9kpQFEP0yKbLENIdD9vdBvkBAdnG1cB1gAeQI5Smeu
Z9R7a+N88xK2LOk5tBpKf4Uj0Auv7JZQreP9Sz+rEMrENbtRqZguj/vWIf1DKGEb1XivOhuS0bHr
PFHBw6VhwYV4ZzUwAvG0iVIUofzcos/cyXuwLhBNLJ9O+jCrhneoAo2IKqVobwO5puzVBgaJ4v37
BB8hRXdD1I0LtgWhghPtpw/cXq3AHPj5q14rmUpl5Js9/R+8vze6ZM6CaiHQFq/UEn1N+SCse0eM
ERD56dPJRI15Cz5suIW3+3t8gVKswXfLZuZOuasSxMrNXlc4GtLKGNGwHg44yQH3BpgWwaV4SH7x
BITStKQfxtzXd5a3r8teOn9SClAMxrlVCKKvoFQ1+LgddUaV3YObZFOklGpVgPxja08aAEnX/q4i
OTgvEERN+swYb9WDUjTDgT5fgE86e00CR6d2KS3yAvUuwh3S4m6DVHtC0x593PGJVcWak3rAhWzL
MPjD/BtNKHUjpfMzpkjmWEmi2buR/If4Sm6AhDlgyDFzd3qh7TUXOdUC2/DhnS92ve+VtUHV/HXP
0BTBM3ZXo4NIDZfODTiajgJ8RT0AnqPSPcpl76h2UHBFQ1oiDVi8Kmp1yaHH9blAWw3o0rcf/RxJ
W38Jmu+ggmho5mWx6EJgCPoVkC9uX6JehItg8zD61fR+WcthrKG1YoyerNTlMLM9GB4naeNFuYE5
CjEJKs+29zDaBQoioXRQtnr9bd1X91IAtYldb0nO+OZFXsjd7sEqi3X6WssYuuu01ibUnI6Jzaau
znTWJ6mQTCXJrE1wbTAmI9a/68iK5gbLebrqntJnTTc6DeJdeNRF5g0ksv1n11hf3khHf4y+3EsW
QmRklHS+if6X4sBCEIojlLwiwlBOSj4El7C7cyCc7FLLgfqVodB21upTM4O14KHQv5a+BfEAiKMd
k49WeCu1bVsno/5wrkoJueqzTYJcZ+Dh5ZCPZSSnYjC25Ux+1yFkAHg7pi/x8p2WRaoCv3VIayNQ
DTKeMELM1ZN9EJGs6TmyA9MLWPiU7q736FHYkFKxhORHyaBX7E5jpBKpKXCZJpb9XY9OkALytfpd
own4stfl0TFHMdpC6BzIpSfDy0rrpfMp8Y7EC9tHz3eTJkjKKup05BZ43zUOpH4Wb+qgIx4USMsc
shcoaNvzFBI29nSY/Hubh3R82Xqq2yuZTxt5757S68rFrIWsURd2r1KXlq5cgPDvyOlAlcxG6hTR
MjovyeMAO5nCM+fHGD3vGAzVTgnFEQMojnRS2ANr4CNTiwaZpCnLL/54WoB6qITg1CxHTuijI6fY
Kh08gttVGihf2KeS9q5KdXBqRJgkgsO17NuKiiBUTt+EVgzi5Un5Xj685X7ZWho9Njb+WSmWezF+
ouUgYoJlGY+RAR+4gy6+DBJYeWVdxkHH7Wkd7pz+XUQlGbBSgRwDS+0INfhoRKqK8NCIINJZBeSA
A4TyIzjBALKnTp3VLmtDK75ud39xKkJujsLWYEyfdM0KZS4WOhx6/M1INxfROhw2aGAW1WH+YwR0
ND3kMp0swnMj2uDa+cugOnyLRJn7TENeXAAXRbNy2ByRR1zXBXZVzVCxk6iV30OpOhpGfiuMwhXi
fClf3l8d48Q/cwzwChPRZ+UfF20/vtMjvHiO6QAufXRejf4qXuhpCOTPNDsRI++oPaZW+lbg9V3t
eRmnqyj943hg5jyzfl2PV2QMwcL1JazaFbEx/6gMjW4QM9x8iUfsKuoynMfNE3AAlx60/TW7igDn
9hYtN6GoMfkXyVs5/J5GXJsjuzByMcHEdW9Y6a2jHeu9NkuYiUhOEqfsb2BKvHDXnop+v7MWaTEN
FskzoA/frDCYul1onvOiCrhNSPnv7qy3VB3eoRgtYp6w1bkWBvyR/YYAj8KMRmndtgX1M9p3pmZm
LsPVLTW2jxgjcPeWJBPMDwsgGR40a3sHzASnbHRnblTdnKOXMeCTcEBkvBAUxhar/FGfgY8v8Aa2
UcjHitdKlz/LzRQQ8GcDcmw5b9+F2sJ5SVgYXZorVpgCypCrn3KcQjuuCcVPHuTnOKXrJvLnIDlU
4fKdBfnBmLQcW7eWl3r24WgxIB83TLTbrIPCJ6NNajQAoJkkyEr6HbOVMFwThcOhriR0rNJKigX/
9lkJizQi/K9cWw2nzBDkVVGU1s4D8Pdh0SCKXgRXOoX1mlS+zbZi6oiVtC7MJicbjhI6QCL/xyfR
xKwCD9YvV1Mlm3VwmJadIQXFOTcccTCGnH+Y54WxYPSWe5zLNtdUbfYaHcv3FMAdhq/gxAXP2l2e
0hFa7OlUykg7Fu6RJzZuwI+wGk0p2czdo0pZwYh8cmzPl+6cqNMIycEdgLki3xkGyuw7fApoSngA
3rNeemKww5yyXxTmef3zZTWo7S+0TP33AyZtKA/4dd/85ZV6QAfA17zZ8DzE9EsPCxyFh9pej7Eo
RxI13pKZkPgEC/tepyFF4gg+Vk2Iop7bYz08CZLanO0KpLyBZh73TKp1MoN/HVcuIYHRMqIJCRqc
ZI3QQ0MslhBVfYnX1Z4wwFElwOj94/nLHqLlF8Aq57HOHhgVTYR5RC7nrJArm6PtAt5q1E8t9nF4
ZktoVv+YkmFg5AbUkFKiz0jb9KIZrIbfv6FyO3tcW5X9jvua1l4K9LRRgk+xW7AqUNlc9pQlTCpl
bkCkrsUMLg6v9BVc8peXGxyClnODYx9VoSX/5UYHg/0D4Dzb99E82cJX/6uQ2lJZJ1qHUuDjBBDZ
e2B/DUBca8NwEesvascD7zQYxuz1tUCXTZoctl1M/GEI5Hs9fat5y94DPIGCsi8ueIZ73vQuewpJ
h/Fk/T8UccxFurV7Sr5DlW7aHHETs7DVqAo24CPEs/CQpIH2sCemqgxrw6LyXEQZQqXesDz01IKZ
bLUrkbYk18hLHlaI7+hpGSm2YKshjI8vuERZ5Y72HYqMM44TEVhdit32bdjwJfC4l4KJlZEGq9/2
JpPP/Er+s0RutZKoaktl1vvrWxpkUAeOuSQWULoigpJcr+hQI4TVLv28zRIb7f5u1seOd5GB1RtN
VbIHlrtEf6uM9Sor1yvyqbc3b32kQ6NxQ8W688ax8hw1B7OTcVkrrLpyYaRBbcBnvirTA2F2ZdzX
O03Yuw6H0U4n35c7PA2vNIz54+0dRUB9FOa/QKWiHcWjp5Kw5hIAuBZrUX6WFyxEEdLqCMFVcNno
Ulz6jtzJosX1IpWTeVzF7xAi0XEYxUyroAH3sFn7d6toRYy5SXOz8du1xNTL4BlB3Ey16foDQQfF
praX8+obZm9lIKwtiF+q0dvqxg9ejlFLIz2qIaNHuivCDv0rnAoFLsW3V4WtRogvq70B8nBa6bi0
dZBM0oLPEKgPQWfENMGKFagzwvDfeB9QANaNE9WKtxICsdSWtoulxY1Wq2XP19SiRomJIzwabqAW
UUjk640OGj/oJ9ZwOJfxEjSKyXXX9PzMGc0IP16X2hl0fgCGJe80lmtKxpzsQgECD+5NNQ295QN5
9hXk2gAi2O4qsGDYUfK7DZefBNKtEdtpmYM9S8g/Fm8e/8m95vxCXB32+R+yp9Awbx2cFdC8VIQB
SmhZkKps340l0TmvrV4mpZO0wf9MtYH9d/eidA8Yrt+rcUAoGq1Hn+zT9DQSbeBsLpP2xAtSIWHX
NA8yfdhT8w9R7o2bG/xwzdFy+I9YnMyvwukfhxqe1RyDQwGJVAFHAIJngq/FKHt1t2GAsHL5cfnl
oNpez8bkAGBT2iteo9DkqWWpp+D1xPgXmpWUSrS2HEyX4ocbv0cYeJaVWaCuZUTnIf6K/nZrmZXJ
GrOxNJPNag0ao+YGCWGyp9fPXwq9sY54ZEE0Hd3QTW88NQMHNa5gLnX89DJ00b/B7/6nTJNBoJjM
o8rgL8Gg9YiCvJHYSkvtzJJvIhDWFsiY+GWOdgu59gdgPCQFDx7U+JHV8H7usylBgX2FhlQCNSEy
BKnrZiv2wsjkd4XRvVXjT5fWbgB1pek+yJKJ79Y0bLe76x40W5TPnuBMLux0dWr8dudCR/69LleM
UQ0f9OdXjv0Th8luXXluNXe37W8VAOcVXrD949dxc9eY6DHHYzVYE4ekDLiY6s+DshShQJJLnZuS
RQgkBafc/MDy71B8lf9in/av5DxqLIgzZujGgcYSd8ge4TeGUWSnkhM8V9zHkmdfE4kPPw1YCeR/
5886atYAkOSFhMaaHQ+zRbByg6zQSyK1gcKctFa6fYQWEOkXspnv/dHNvnLT9i//liSDlIHuA/JS
L5jpfGaFda9Ikd2Axf2x98yOn3Y1qGf2ovVk8VdW0KageNZRflE/mruc6Gbn+p+Ok1vaZXrVdIxM
mNMYdSqst7RO8RPPL069AX+Zc2Prn7mpt/9tZNNnoSm7G0pidYmbXy/+ZP/58KI8wBdQ9PfUE2iD
Y9kXWbVlR9MvjmrTPu+A5c27XzQ1aoGGgtSP93vj0g2Ig37Jr66GHWVQG6HW84+AXUDskxvvcdIe
X5cjKjDOEcRRzAIexwhRR8YhKo3oXALP7bmExIwmpuL/edAiHWhqn3V5DEupOlxzvE56Vy35Nbuj
f65I9hv9qhu5+eI6MVm0laDoeUR3pPcFKmdsoJJeub5I9ifWtCLo1cCQ0waut2UEorj5NNXrqCLC
P6DYBpbJSvWJ+Sldyo5Nln7lxbeEpM03nLZBjCKh5Zo2Qo/HNTRvDoq1MEaD50y6cbR26bQ+tbNZ
fp4fxS3neunGQu0hWbY6QQGzxyzcB+NHNn2MfjwvqmiwsExwaMi+HcSmkYtziyZXRijFE2XDu5mz
ZsZzmjzxGnS5RdkwQi7BEtjPNqkfAGjRJ1dK8IvQRcS0vf2QEvWz4i2D9gzsGKGmO1Ns9Ba9m2FC
BdbBGFwPWwYbo/1IUPiZ3waEiNeRgifbq6dg5vDRbDv4DECDac81WFMKpZV2tFHa+rCSL7w9YxE/
fPS0vvOE3V2J5P27DkjX7RHWAYJdMICT4F5E0hL2Q50djER1aA6qxT9fg1f72WEmtoMD3oOQEM5s
9/uTAnLzZ5JiGwZjyUHy9sD1faqgKFUeBqmT1VxvpL/KSud9FrPflJ/+bCdtoGp6tQiaxy4JtL3Q
4eNnefTdkfep8hRoMTpEX40F1W34zay23IOyf7FkvBrEkd8VoUG0tRUrp0f7hheGX27p3WcD0dMh
PTCqr/zS/WAYd1wWMNh8dvvo9z6TxjVghjBMHbHFjvG7OMJ+C9aT2UbYoo4cdXOpPqlDSSsYyubo
Q0XZ5LCJd8REbFr52wqjDvU1Zk6PonHBamAq5on3ImlZtjLhN743ywsybL5ZfQjzkFLleE93QHMW
HONpoz7KDSa3AKkdyJ14rf99WXgjAVv1eQvJzsGtKhnv77E5Lw+ob4Iia//sTxSSPl9V+dTkwiQ8
YOwyodFz/DNaIiujLkgtgOS5Frik/Tp4RRa4YtTU5AYE0WtonShTUpUlTF1D2Fwr04Ia5MEZVG/d
1AS8fzQBcDzbiPaumEUPhoVztOTW0mxud7X4/YQtHZ9ZLFBZQ3FL3Lhbi9ityTkIIqRokQ4cl0lH
hRqHw31jFEm5tCaYps4HxWrtZG8V/jxUwl54gGonZGyRe1zMtl3F0acA0IAd/wYPZCk2/niGDg9c
AkM++HdAJPk3noJ9VKNBhV57DdTsw2nYdMdDyzCnRZpt7+yrP6YpC6NGytWBp74Frp5AFI4NSo1A
GItwtcENHYUSTKnzqtbXz2vzW7LaYa7/XOHmr0Kz/MZ0k01WJ3cumANitVMUUkhkaYAxYh3g+1wz
yGo9RbSNk/9RxBTONvtsgg410xsio0Tx/BLwBtT3et2KIPR528/QaLAkAMpxyZ8bQBsWisFi1NU0
FKRaibUDHKFjeDkScUCbkYx/gyVvhGkvoQ7YvDQmKnk95COaBROdOGS1HSqcJlMPaZhVTrLehOmB
6C6OLyRQnLG2pMUkVHnMRfiLJvvO/IJrWQG9MQvSOR9EnuParad/gbPXROuGTMgz9PQXflSbRbNT
VBvfLoR120svsh+9lUg7JnikUMhQuJJuk+E97C58HkFpJf63FVg94iqKg6CPZtzAZHXcWppk1hgk
b2xyTU8VHl3fFD7mtUn1xtwymzoe6ixfteXxb1l7S5v/OJ1cr0ImGkaRzNUCGa9ZPVtF/TzUcDE0
8vokDDHlekmSSWXMQcQcTj1MhzbEWfDMT737F338DQXOxxOaT912MFbVTK5lzjPrNc5zKI4XIlRJ
5jU4W38jWdZK4X2fI5KF0CDGf+mu69fHXYNQKDLXyWtL4xu/grTFEtCz7qpmPEtvrqOc71BiYcbJ
UOKyLYEWJMDpSXZYwlOFJbpk08zTRzSmlec8hg9FWVLhSvs+wprIXt7gMfBgRccXkyWMkt+I8mMb
a7OUvcBNe67QeJ4V/fcwlvbH6sAtW7owjNqhismYGC7oF3c8tbd4UgPPhdgCo7bNOQ672nGIcjex
K+J43Qp6GDyBW4IlixIJqJxTXSiJs2pdEPKaqZUuKHHteTNW6GJxxc/1obIOx9P1C4dx3H5IeRVk
/00Fhz+/Vks4dZPIF9MmCQ5WWUQK9enbs0eD5kOpSIjvxKN8GdwEhkbNc+ofGsDCyuEv8stgPuEO
yuhGQ/8juQHlMYs506ITLw7Ew0nabOGE7/SK1ebgxod65j6+bSx1Jul1a1dvoKiKfZoZIOBOqQiW
l1q5dmnfIcG15W/jFNwxAQzBYjiHLAOOXaQmzeR9PffOErOUJUNlWVxRLjhue2n/emLcgyPdyywW
axI+A7VCx95ZWP+gFJ9Qs5qVnOj/Z0xE9MoJ/EjMdx+7IuzzyKtOxKzwJ1ztkwDvotVoZvPE4u6j
ary3ZEOdG6Bblg2bKGt3OAYgl8YSuBLiUimcozwNcfnkMIg/C4i7J/PDQcskYw60EkLCoQqteQn8
uOgPkKoMwsTwgwPwdzTZE004Ot68Kh7/p8/vM4kxW+1tFV3xr9Jrmgz6xkRZuyg3IYr+JQgTDuu+
3DAzbBwH153LppvEPKBsPNWSeRJPWPCeNGowxUQEQRekXe8sZqd5ukv9cuQQVuRsE5zi2pPDI1Wm
v+W59cp1MsjIJK8PXMBdeHaP4Q/ruidQMhIXut6p/fTMXshWRqdHM1ifjyS7LjjApvHVI5P+GmX0
ExeKsxaekzTZUO+71aVcBUNAGdnBPKpXmx2Ao8GdU9BEJu6SOc4w3mhCrG1FmjviVPgc7VXcwz61
v3+E99Hyd8DBqkKIpQ1jWNF6ppaa5FiveIVnAcH33SvmVOdxA+avroltR6xxnXmYkBCCoWA/zIiB
2k1RgfPq8PT64tOxoEMRfkaE5HVIVvn7OGNPs3KGGWNlam7iJLh0b+rkyziO8k/RWJrUn6L+Wo9L
JzAu5vrVT4816o8KX1KzKVBQeEEmOM+p0P8omAql2DPpObFiJTLdJwHvXPlQPmdxkezsNBQp4YYy
u163ofQrpky2LNAVHdxCnjW/3Iifd9BO7ggKYUfy1RLZhAWAU56FMv2mhNMeJzL2nK/m6UKUzE5c
sL5+8rXw/BcJQ4nS6c92YdhFAIOTTW1qrxc0RO7xgc6x1mqlE3a0bneFcYHGqfkIJ7M+4yQxolwV
Kg+5TdyQZCkW2f4ar/7qlhtLn27WGuAbTjBFapn58x4IIXeI6dVS6KAutmzPGBd1WI4v8dWi5LoF
DAFUWaf5e3etTl39KZ7hIBe0GGR8e+qEsNFYNTh1Tsk2p2vg1eXJsCdZ9vvcAf4taLAog+6sbueU
IvtoOTS8UawD43saedcPH1VlHRqdQsJFm7HylCfutd5is6Luqnct2dq9bzw/2taXD39YclC4VV2u
w7U8y2p/Apafe6RHZSHE0Lkm/FvGvg8RtmD6fyWAeaZzh/4zlID28sPCZQyiCAIkaBODqZ+x/cdP
ZH1J54GwfhXePanzudgjDX/as/L5lZRl2Hn5ORGonmmSiEK7BN1CT2P7gL8U1Gju7o9A+pbeXLRB
jQ31toPSt/CI/qsn+uoQ/qFYgPJ0JQ5TLhjnEH70rHKhmy+2m/EGeUN3FCNKlrPjdsFCL9z1U+vy
XTiSjNs/9QIK4pXU67q+nwgWPNmBmeFhBjOENZY98SxqBCz6yaYX92PG5ySiR1OCEBuKbK4lg4kO
2E8/OHUgBBAY5gKSfGr9cF+WDjZKOZxcBG0WU8b2yRsAvAkjCqD0Uj/zslwve4YbSQgLN/7XICvw
3nEuvglCP3TvmliaOjmedbFfm2UVyop/QsMC+FgptkUptvdR+dSqF/aeDdtMWsxV0emQFSxShWuE
Exqi1hsSidsOfZ9QM0o55D3cGJvP+BhTFWM2TxYQ+hZaUtmSStZ1Iy107D1zHEhhiyAR1hFjJfEp
haD3igydO1eVNc14f/ZY9pudrW2tzn9HLgXutgiPRBa9zZBFeWME6gFv6OiXVK3ihvKj1bRevDG4
8e5SDoFURsDqVFYh4XC8MCFte1LEMwFQaxfHGl9tCHJ+1/ta2noCy57GyZz9mDTRLXVdHq1elkqK
sw2Tw+L/cuGmznlMQIj7lZMO3VFqs57xFt9cJV/3U+b8pKaw+KlExHVsVBO3kwc1dqP9k1BC9kjE
xY9OP8sXoITH3l9XbLD42EGIoWU1aaSNl10zQqG/W6P3eeiZG9ui4G8yFi1WkhvTJRTtt7j0Ucb+
JZPQ2HT33w1ennsI/3oMfWXqjEw4ENK+nDbwoazRMGFR/15HiPsdE19pujNkKP328VvvJeg06RIm
Rljyg/K32StRdiHSHlFI84AK4O1BLjjET8pdqHHDaMMRZMU6e29zkDXMpuGtS6kDol0PGf1A6ewN
usO0yiu8c5qdWZmiuCllvrqRpO1oykZZ6dbMFYrwdqoi0m8DtX0l31+yuJ2sPH7zxmB4TMHhjb+f
F4MNTsFsxi2cIwOVREm8kiD52HwH4IoEz6/ZKZY1c9+NQ1fjpW8l9FrpxsMaIuqhiBviuaYOeSz3
EZJbxjftZhJPtuCQ2/oWCEpwY77i9XO06KaxC5w3ZJTk1tB2va7Yrplgak15zZYnIEsDhXn9R/zx
6EaLcjTs6gUzT/a4LfNzPvicsis6A4AjLp41Ii2h4AnRKJfSzKq7gRtvIYNY+SF7TOqj0dU9RfUf
8vkvLn+NghinE2k4Pz0iN4fn5+tG+nl+Um0CEFS3sR+KYOjbkvid4AIapYa1PiAYmdx29LndVKQV
9gjLz2NIeuEgaGqjN5ITW4q/XFU8OCYbRAtylf6OX4RnGY6h7XNykL0Rg71P1f5F8lV7lC4KXMmj
UkH0u4zQjB0IMTalXdiZR0NBqy0aR+UG9VCEss57Pv8wM48vpv2qh8XWTaObm41tFypaaUm4qrqT
Jx2cLn8ZPrs75JRNQv+ZdxMq8lk4jfv4VG9Atu2o41aXe0FkR9shq5E5wZ8yj0loi1CvjS7rn3yZ
wPF0ScgZBYM2X/Vgk1oyBXjnMzyl0CcFBcjLvlnMCzu+ll+wT0OrOlgdgC9RwurR6pRfFMSX7pfA
m/M1vRXEW2sL+FW/4eSMGfabSvQjS1RrFltdfkwOlNy9vl6lV/azx224mjIXG9ly3crQkV6WhUsI
xukc/hvG84zhSSsNyaAk5XsDM3oBRL317xRQADiojPyP5r0ubFaxLZ3K1hOdcxC/GbDCSVp6kfSx
ycNUwLkwWU2FE/FbE6RenP15+kZ0EIby919GqMTRomgJ1GtjcfEWfOjMSljRJm4nEVaWEQrPrM6C
5Bp24wqARJDvC5kDTE/hM2IC+J5b+F9mFKglCScJhWgyYevz9O+9r3HQmdUNzgoMq/VC64WZUiUD
bxGJHMah1Pcah0636PmGqCPEzKpsV8uoDNbb/ea4TOu52e4ScE0Gr6gH0ZB7rUd9oeLKmOCupzYS
oDp0EMrP2/HpouLHjDl4SVk9rfc8IksZZ3XV1cuUpVsWX9ZXwq0o5Z6AWHH8UZ6GB8rA3+tUwBmu
TaOvyy9rs2Ekb1GvYLgK2gRDZti8zvPh643M0kCnrg9TIBl4m5GpUaQWZwMAbS61ioW83PaQx9p0
NRzHX+bdR2loszH+bENxXfVQqFUBgIwfezFlzT7WqlDtHU0a1AykuIq5/Q437zDaFccyK61plQvZ
r9oewDkXj+KV+4zs7jJAysriseC3miERxFwm9GeWLpGj3/vD34TID34bnefWK167fQ54fiu1ncMm
fYXRUoumoASHtiZNr6wD2yux0ru0ibxXFobKymRcvWFLkMqPhduelaj55wHN83RQGMdQyx9zFLcN
rEeVC7g8ZXcYc/CCjeWhVHvr2414zeeUNp4WkxuGud/QCkEKae/FecZsy/ed8BqEEMAB1jv/E2W8
uuI1mXHzbLRzP9+he9NePm2RRBsDHCWHyBwN+5126kqYKeTgJOBNdIHPtV0tSk3x9rbdrTs926sy
OmK9yGbh1mCuPT0Rsu9Y3q0pBWjieTeLsyi9Kkm8ugZROB+inv8aMuhOOSfCVCJLVI8nwG6c/6g1
0yW8IxT9FG/TOGeKK8ylFGehBi+mf5aOKmzjo9l/tdkor0mxP1oKQS171ZnNpW18d6Yo/4EwWYff
lh8ke9SCnS4ww4XV4CchnwkghE1fMdYdQS37ClcpQ4y3pd/qiJophDWPb8hmKEmJ+cFYGQuQ7+ll
DgqIGG7ax0dN63VUESAnTgDo6ER/iKYxqVBa5vT5FvmsdF4/ZDlHf+9xNwLeGLg0d/JaSDopwZVN
bWBLjcvvlW+LY9YZ5hjTltmfoo83qCi4Y/fodJv4Fms44djbZQjMreRWZSb1S0RS6375ORX5Vtho
0JrTiXyi9by8MLsnGV27b7eC0yPDV3FBVTegvy4xBPZ3Gpn4BX7RSVfyFiHed2NdXavxMpuvtL3T
3wNyH5llE4IG9bkgciv8hqDgAISrDpcFBxHYWnR/3krfKeKeKY3KIG9WNTfxkdcVrb0Uqk6zKRPo
xK8PqzsxBfn5hl+xuSMOmWvPLPBk9m88rnuwFKBE1Jsa9qEsRNzVHRO9jdxWcdf3IqptF1ZKSJvT
ae82lHpWUYOC5H0efpAL++Kvkvn5nYNFZiBekdmjZ6huP52QXfcmcbxQYzvDUeX/zktvW5r7uqCz
woZFgKkmkQTUQvSsQ0Z4MLhIMfRXC2q8hdKxequ6gIRTIAs4NK3yC+pyocYoDXVEVmNfERpN/gjW
C4Rzx9VqGh7b0m8aR39ecDB7jjRpOz0e14/M9BpznfIwyu9B3E89aH9iFEnINpr0VaLRu73bpQM5
cb3QDzfwfeE2rmXFth3DXqELD/R6NgTWhQGXazFQlXwhJP419h/495sv5IzQj5pXEggQLrf8N/3w
dvyxEeoLSv6MsKZRDhqMQdznQ18I1F8fLCdrAHCDQYnnY7vaV6IukCFYw6vPZTyBLPY3Aox2cC7h
B3RlO7oUzotaogWRraYB0j53k/Jg3X9Pea75x7Ga8+W4cH1fBcAcgb6aMHX0sUsIwJs6OfC0NZhd
KtMU5HEo9xI1SLjnR0sZ4sxVvSvkVnhA+eizkP8R8TCTKK26usdfvxviDF66/KhbkCKFgpBkD5N5
FmaUKQJDCkmePYu4wzgZ96AQfMlRHspTY3c7oOBaVn/J3iNFcM4y2ejuTAWxW/su8W0TzfnCT1Mb
nT9clkMHnlKRxhjhBkh2CTQvpBAgNUBlLOIQ1WYcrgeLQZxY85r4bUADZS1VwpzdIr7xJHlhLS5W
YWdWtIRxWg9yyH5xZvbWFF/hinJp7XqIzPzwJg/yimmkzYcsiinJQ6CD63szvIymXkPY4vxZe+Jo
2yrJ851kRf2fPc6D5fVFTcP0PaeF6kzoq5sRzkPhzenzCnztypBSZvYeEOf2pXVmEmQaIh3XE90V
u7wdmuEaXq+ebw79JNi3qlFgnmQn5//RiAW0l9dAGkj5U30/MVTaCHvo/ziiJcbB68gVa050rqi0
ZqdSLGoZ7zuy1kGIt4X1uZhghx+xHm8ONgAmdBSh27ahp9hsjVt8gCdzpaEVn9QEdIkCXukokXoX
xrGmUnbvTyGaOBqWI+Oww8oWxBSVxhEPj6LrdbCq+J0SXFcZ/HLBXb2zFFw+AiMAG+cbU4QnyAA0
LMdUO1PlvefTCTu1F79rHNaPvZe5qS4CCE7fO+5/v9OaRDSPO6LxL37kECHZ1aRoyZ2sJzPQgS2W
IRGe5czTpC03uuaVo94wvkrl8yJ4LO52U4TDguhh72thD2fph6Dtu+l5qtlcPm3NbKs9NgDUr7Wr
NJnU8E+8Jc9hI1nP1nekw0Vp2vegOSKbaxvylHj/UNUZOaTUbdE+UBgZWNWvIm0x4MK0LjCPs6XF
s3Jpa2ZdH/EEpNtNJc+HlMQhhPk6jD8Z7VRHMUKMdTMyj3Htiecx5ie/GI3bUTxfAeGEJxSdgpiZ
yxMFHZNHUg8TNAUexTsvnlSbn+JPTEtyPUPtT5ZX2XLow0TZbs2SvhEpwL7jEfWFKtNuadqo0n91
pwccZfN3d1FTAaSUAH8tSQlG3Ufxih/eClXLK+MqpEBRYyt+je8yAid/ZexwMjV97J6GBGwvTT7O
73bI/2XE/Dwi7DENax8S/B07mg2+VvpuC5iU0W7HkTHVswvMhQubYyoL8nWwWImO7NPjCEOGOSOW
ZDeV8gQRWBE9gsKkmvEQ+tqLZRYVv+5Ie4P2hQAOaIuBCZ3/TQa00mGSemat3Y+zFjZzH+UM1iNx
04SCa2Ecbu5C0Fi5SwwyzqCR6JdbEWd8dRnnnOXQV7u5LjwMyLoCrV5vuSJEuxs6hU32A3Q29Bzb
68Y6QNb8uGUgC4+6evG30NNOOehujG9w52Qc0hwONcPZRMN8+8szC1AjV/9y8N89xcVei4MilDkX
W47jwmvgin4KAWcz8OAgCgkVyT4UJ6kR1PwkSKlKSPmdJlymioUsDCwXG4oC4Q1kp4sNB8IlxwTe
Yww7uCX8N03NbTLq8LR8JXeov/xdmgvMFIeneNvEIi6oHKT2Zrg/TX5bmXIX58kh3Q2thMEXYxb4
gXwjY2VVvFsLeoLxkn3OishW5BxjTbgOljG7wLmOc8wJeEzV/dDHcjNndADwCvRezMyzD0ogvGyn
KFZZ0jsjwgGcnVE28Mh5v91YXBfwicfembv4mt2LNJ+KM4bO3Z3rmFQxgCevJZm06JdsoE14K+1G
+2kZUlb5+CN5RTKazncbgOg9wNKWsOGHHKkTdZmngueUHvNRgQ0lQFoWg4gUJ3sDWZwom/MasXxj
fD/WM5RiwhKdAmKM5dIim2PPnosNKMAQTJLFExqyrCyKK9d7VnBYj7cZsY5zOIyyWa4dDJRko1Tf
R8gHAHnexO9W0EU10NK6iLUe5xOl5gVpyvcoQ2Cnud7Am1oAYPncmqY+O0/EmKtgdme1eVYAqSuC
78i+5FehHs1M2kcVJBVwcWICVX7wvdpSpKTi8joZRGd2iMUK3+OGTQjqkqMi541Cdl60I2Y6IG23
u+QwpSgf6e3w5iMYcCf676uTPzfjkeMWmiaWhUNbA+YGXPjt3CDeH7S/n0zDiLaNFXO22mBWE3Qy
z+/r5BoYpfk6T8zzGAl+f766eTn52ILef/J+QetNVyHZE1F0PQiQ++ovEd/iSEYuSZVrTn7cGasW
gIz1IygD5ktCeHZj0riuJ+bz0f9bBMvEfZXQW4MgumDgjl+lrfRewfICGmnCx5ozTCm8Z+J/enly
Mfz3E+ONzN1KcNrzWRGpblqk0vg+xayaz9tA4dUdse5V4qI0sYbMoKPUWtInJE5VMu3tNvI/2WBE
AKWDFKpcO06nppRGgpJE9pk/Qiw+SJKOV5B3tUjzlFUdqB7W2hU8mxJeyBO05TiZkZD5rZYdyFku
s1SgioeSarAw3cA+HhKvy4gGFjNjdjoap4zI9fgjoHYtgIlcaR9DbpNghgaNnZByt0s7tYwGXMhI
eaJezIFdL3QxxSGOYgeR9fpD0Mrl9lx1pTkrO7rt5zC4VsBPGQuQixlRJRmsKd/SpOyP/WpI/6Ym
Eck48jkO4lOC/IcC2p1dGPYUnjtWWHkNxdSsmCH5ggmfBI7hVSsnHITXmJlBSV7gPeA2q38CcYXm
9YIDEPyVPIQebByelMspMwUO7LG7PRcrX8jq9qqZAfXEpxzHIycKz8jzLpGRIOUYd9onCqVboKT0
E/LLZx3umvSpYLKyQpNW10TgqjjtJ9C/J8YlAklNCNLwSpOteTNdxE7oriZtaad6DPyyN80AdnDp
KQCsP10FjOqiYWDp7zSDF2YHA+Z2bMfBpiQ8vt7Fm5sx4aDlgNadAMMLdbBmMr7rl3vfzYj9DYRC
+hSjTtpt2keVvlk3Vrwt4UDWCbGLh4ZTVZhVqihNwmK8PT/wytz+6/sLe2zxi5jA6wnriRIsB/WD
M5zAxnMY5s2h0WbcR9SDSe4RZQH414/6DNwqi9PxGEw0IR7xdVsNpGmnYbZNS7U4IWQvQvitF3Nc
AmcXdr0mJzcKLBYhLD/e5o2Gjd38bSfRMe8S57xVr+dPBzyWONLbFZbWK5KNAcZf5APJ5lQ4Vk5Q
x3SxSD3eczk6OkNyvrRtFtvkAvkWbNgX0ShsYzVUC1On7X9j5yuoUeekN6aZ4eSOVNiX1FqpYJXA
fTG+uNjiWeyDrqUg017F+++Shko0G/2ANZP8d4Jp35UkB3aZy4BGwpUgL7Pmgv+eWUnXFuCeHgz0
1bTnCmM6IayaE19hb54aFk7PokjyTA325SZwDAcLI4ucYmOa0YHrYKwC2+R5pVpiZ5kTeNpgS3lF
VT+vAWKH0VFhppgbgzB9It8dU2/7RnIyEz38h1DPpjVo81GyR1w5mqJ2TXRGXJHbVi9ZdQcTpScR
L9Hy9Ja7lT92BypatjXsMp0R2srloKM4IQYdSfhCNwEl4SYvHPODURn68lTjqb/J+uzTZQYTEDCb
O0XMSFrAMqE8RZaqTypLpx0gGXz9h9YlDOzOEVHzfJ6W4sDQAPsOupqic+HjfdxeeiFA8E8fL9Yv
/TJGeDP/3786zeWjK+i2ZEuFK6wzpjtJvGHsNlsW6bk2bZ+3VSVUthdy3oo1E8ZcwebX85dTzJ4e
GuvIac4rH8b/RhOSt9dXBmSqE+P5TValVSC4Gl7a2bg/GQKx0euGCZNyO8sHVnywtKsRm5cZoV9O
g6NoEo2KGxI99gZH3mgwALMpvVh94EcycV5f49dnBWJcfd9NXZ9UAmfkYH58O58U6nQN3t7NrD4i
0YbIyyXZVOc95LGFMlbZOUldYuhz6CztIsfuzbQY4kiU8lRuXFRKscjmHFFaKlqwOuQRVX2FOuTF
RjZveGo/lC6CJoOZEJEMHoFoBw2mb7/SkAVLoNc8UkGwcxkwhoUliTQxcf31MkQkxouWDDWtwjcp
5ugIZ4TCuB/shHbTspSIfVRLL/HD9G8BW2IIGSV1l+JLuXKYb3TSEI5Fwmx18ISScliH3lgJXPiM
faXtgdNPPV7Y6JqGeIdjpf/3aE+rr1skRRXFyW9cUesWJpeX2uk5L2Pia6qgcGrNxzedDeIH4rti
1C7zc6WKaSW/PXfVyjfqCWciNCUzNodc2GGrIUm8pNmD0JTph7NO66LTX40AbSqrf4qs/DcHJyIs
Ft1UI2hPqUtiuwbzu7jUzTJxXwBCedkrSmFl1cVUOsUCvAx0OpOKt2oIVlF7UqNbn21hkiZaFetF
4d8doxZFy6bgFKof/7fDeZuSKx/GW3ifb4hqul1vBBxJrdw1txQHMkSprz+Ubvay5/A18aXBH5nx
fmcLqqGljOX40bBiHXg+1RKtPq1HOscQawKaN7zFwY2eeGOv7mq58NOGshozcBpjjO9Wx4SNpilp
V3V78BRoHwAcM7K/iCtNDuGrPVUOscZhc8M9ghaBa6EcUu7oo/YywKrEgPirNoQorevvHsoZ4Bsd
X/WRaXteKMNPev9UUlEtSfxTcnXl+sIpGmqhIbh58PyPLh7pz+AQxCYOde/PKxLL+wr+hMH8qB3b
SQTQCenevYyObwxRuqcvTGG5SeZ6G+Jkj3jlocOBCmvMnUgYyvWBykHJImydZvkLBy4UvSD9nUw6
dA+PhzuRKw6ULJIeP+J/JjfxuRIxqUDdk8L/XpW6GUyzT2WHBvpRpqZmcS+UIYIDuMgRIQLzAAnA
VBv6uVkNDNCjKCK0c8TeNkGHH0tLbCVNrJSY42HPtsss3e4qdT6zDZ78KlWupFVqxxtS7Orxrf4K
DZlKZf1xehUiQRjiARJgQHXjbpGYo8kBjwTK1ulIYhCMnBewMFCxVVnu39hF219NO5LAsrB7Nnt2
YT4ZiwdFmGbBR+KiIyZoi9yFdM/lCaYsR50eWQdj0YGvW6EUGDwe7QnMySXUemNpmUnny9ZAiTff
5DwFZieCTbYhUM+b1Vkn1Kia48rR1qibKaFecaDH2Cmh+q1eIsScACZLF/V9h/2tfz3kqMJU27iY
Sfopg7lclcPV90IEA+XEt5PVLZk1sy+WAKFGogIicBW2j7p+jrVQafJvQpLg3tOsRRqAQ13be01h
2Eh5wRTMmY0OXgK6Rmsym7hmm1c0bzHaeRVwb15c2TqwYEF5hFLFx8+5mgkymVPHNHCHopW1lffM
MgpE60Ft3sCUpy0QJwAPBQOoCmLI+Y57EyHmYX4FNkWFkJdca93k+2grclc1tbyrXjgXtzwNI2ju
q2GPYphI0re59q1PgJBtRsWEZ8ccBYr96qkT+4ohv0XH4THkLkRVuvTBkOk5zuuPRLhYrVVL03II
3YnnHXnsKzuR6QCF6Pt0s0T8ofSF+qAjisxMTVgV+SgM7ub1r77S8es39AWFEoPgAAMsTlzYd0E+
NuRJ7yzKYqOmsYo4w/1lqumDWw1U6oyWuVx/S1Pb2LVWqThV1agjTcRfnz5L+rkdZndxFc11Ypgy
gaVnwtrpFNrRM4cZMxruh6RCz9v3rxgiufUMoIY+dRn7AOOiH1k9Nd9bY95HAZY5/XRmVwSJBU3Q
pDHLaGphM7W5VlKtS9tboBsJ6FGbxGDWuPZHxY518eVGagKlDdvJ9nVGKleg02vm7fezvJH/6xjj
kAcKH4b+QJ9YkShJWGBFx95b7AxVyMLy8rmB672RZmPj1sOPIsYxLjxmBRnTprLxS/RtYrTu+GID
0HC8emssJ/oQ+SFuAWSQsQfmOQNdn3dmc80JHWDHBXMPja+7wyacAtfcRXQ1+ajIh9Pa5NSPeN37
lasMQ6sD5cA/SwRcIuGYMPFGoFPpnz/ia3JCerVbh2XR3N3kTcJKF29zVNJdRl1qedETQhCd+9nQ
sDXN59ZpwsznbVpcECyMx226uKggg2OGQpx++e1nTssm2LWYNsnsaQUi+/4DuvfZzAUtKuNfqAXx
TH1OIUAE7DQaLD6COWQOnd483giIL2HOLIR8p1AvwJ/Xwz621KVOPxwFHbpe0HNBGk0PYpxX+d1q
Xz1DY7mlPLVVxjwzG9gQyOqhKI1V1up+X/hEx9bxz7bP2y0w+AvLplMyBxo6M0J8OUitGseSsvOm
XbsTqU04dzPhSkzTrRboecWyg4aLLOeApzqn2YVnioljdWFZcGeF6J/wi9WErV+0OSyzF+k5A3ti
V1CBvr6FukgwUom62AY3EcjjzwFk05dwjhqs/uxclPq+Ko8YC1EAZbOSa88IyK8YPhYMM7RkFJr2
HBRMifkWKLqeQCqGiGpnCGacyFoeaeiJ0GV/iyZFOL1i61DNsr+anFx2TwTIv+kk3mNCmuB0axGY
txJasJIRkac294GUGLJHuJFDFNDUeA43CCrljwfvcPdG4HUdvlSHzXr9UlBnbhHlDfdMxq4fCnh2
M/P0wstiFBZ3gf3jPfw67hU+lcQIyIdAI35+imUJKQuMOqEWEnpuULKIgyES8bzzHUhAzNQwN1cX
/XQbnl6iQd+QWt6gsrxHRz+DBmCkKkWqFRKEOMLQpc2CtH4XgBHpmwl1PjR0J+Q4p0RMfpC+OLdd
O5Ni95j81+utZYERm6LcSdGs+dUMwXaG0IxAhAv+Li1O9PCBFYpt6URefkQ9VLZ5CHmjgksUj9E6
NyYDbJqvvFg5uvZbtx5JrAg51zpsMqs2Rh545pjfWJ9nZxEMNyeq/juwTopGIzDdMaTV/zoSAmgy
XtDdAQOlvn2EtuUG+SF4jqqwi5awjwFkJrJRimRvS0APKI1DrW9xAuQFsbQOm9M88pmeW8NcYmYY
yEQ4v4VFWC57rd/ge9xTWNKdkFewjSYkq1/8qBthktw2rqyAy0oRYqkAKPVN/hcMGxLPnoUv6SGc
S7qAZxQajeqEm7J4GjMdKrBfkSqybDhCMPaLDtHcP08mYtY2fI8DXmliqts/A9SUCzztPEzKy2In
ENT/L+2qXYHpvGQLWyA2LHduwsxLUs9+dCilKCH0jP8xxD3PyGYsPb43pA0fdERJ3bmuPUQ8d4OJ
BIofqhf3s8qQkblmmtPdPNgaQN9BeIEVl81ou+LdcHlSJn2snZyLr98jeYZJmQFHsTNohjmC5WNe
z/JrlkkvF62osDWdiONxFYbpIsHTzbg+EfDydKiUuBT5k5cjZG8DI2iyLSISOJFC7ofEYYYtM2uQ
sC6N2JOPB9/gP2cwEovQykCLidChg8VsPD0oI5SN43zA6ySVW4XlEpaBuAs2gex/nNkv12wTSp7U
b7G5rqzsjDsXqLwciBqxaa7HONUOhelcQXCzbBk22QSdaGqG40xImRECtDqyr3uwKaZk84ZLwdEc
LXpFz4eQza0HuYhDuMMH2qp9ZAzIYzTLy/ApIvstZoOcfVA+GpjsmwWzTO24FibpvGVIejFRBEV4
ZcVS4x5nujR55ke/DM3kF5i4pAiClrtEKN+E85EZ07C3v6Z2+6YGVxEhmE8Mk9NGrSfz4NvMXiT7
ozDF3/l79QVzDQlc0nYzFjGB/7m3rAfGR5wtVsggZ6QI9vy019/MegTDI+uaBlKMWuGbCUS2rZ/h
eT01teSPx0IwREqC9w6aHjPISRgSg5mNBL96vstTj82jpexj2PtBLQEiyZ68XDyxeEh25mEXBqee
rQ6oYxP29qLvWASYnq6VGpb93W6TK7d3aMOGXi2IIksQ5Rx1MS9DyErxwU06sNMzrc6ab1kf3Lxf
sZIb8HRpWDVWOWCWv8JTQtPMPSpJaITV5+sGP7m99eVRzVQHnb22a5PArnscprHrfxbC/+yxflXi
zBFxAJwbvGiXU4uUjGfkMpXxVZTFdtVgTbVbmYzBcxMKyGKFkoVjHAh17gMcFNXpK6htvb9fLVC2
1DDt8BMzIrIlFdAWVyF/QqiE7Tql2+i740CBo7/w6dNzPi16bsI++dldSxf3VWFagq0o800FvzxU
mYpuiE5b9BjCBeQfPzTzt/B23kc3BtKqKY98nx/EH28AqVK2j2mPdVR1XNIcx3b+LZW8vlB/HVC3
uaPT80yF1vRlWkviFWbWnLkY4oPXMEH3IHELq3xgp4+Kl40gfIe9C4CxzVlde+pTeUQogN2l86b0
VQkn+qcH03Y24Fq0GKKdUpnRmd9spyI5ttLpziojD6Dqdu7YWT6V0EuNBBhs2tUw8Y1hy76ovwYU
oFjjZHakitf97/ZTZvSdb8XXSjYMRQ1wrTgk6hJKkAXx46xi2gh127x13Ye5Xn4SG24eGRHkjl99
+0dj05TiQd1a3YLMwSNpt6+GFI6Hop5R2Dt0b2egYoTKqykxO6pxZPKbAP2ZYE920XnJATwtG622
rJbTMvqPdiwxqgCE4QzZhgwTYscbnk+Pw5SkH+sd3Yi3yHt9nImfn15yJjev2iSGIkSSgBZ5ox7Q
oNkgZ9lFOppbxR8CqyV3aUHlGz9ZhxJPEYsHQ7TsnXoxa9lf1u6191yIkOXmeUkBGXUNFNpWgIgy
kMrt03RjT2GnSIYef4ruJvjT98noy+ZZecEdOX/UPUoha0MYWVXtNJDXvo1lPHI91cyTU8jgfWP9
ak+RP3f4chI8O6PHX9l1xA5UETnx7Ygjj5EU3Q9ODr8Nnjll+hyxekRIAUz3mus7v6JF2IO9yVqA
osmB9xukA8ohMbUXo9lMTQazWtGW5AVGu8UI7gT7qzP0jlmkTxJDMAHbBMJDt4ORnipszDdpd8vi
/YHGRQtY8hE1vZDwWKIspgUanohkLUBOpXr121cenul4CmjkIuxOkLpNpqkzu75HTlAnrKX7lbC3
wTidLXQKBw1uH3toKlBOBG9s2txxVpjVaos1wIMQoNp/FKHJnqJH+Qli24cb4CIl1K76n3F96OIw
mzKzr8EWQ9JphLQtRVweqVp7+9WWSa85j+2g01ZpTz0e+epfH8JSj2872X9cOuvapOlV0K8HpaEN
lDuG43WSvgNREEi571/34DiGWQbiJu12HNovf21ACNHrRcl2byuTJ1PGqA3Dtwl4zbHCPolBISi6
NRdSeOKNk/jVFQvAB7Wym7JCVUjE4zHHQCodQKVUhuUzuMVIYJWdf0SQP4o1mBlx9/P0aa3RfYq0
BdSpKsnYB/lIzbqZ5vvivGt2xtRV+TitaEwGwLKf06ixKH7iwPxC3Ym+xTq7qZnvoN12IMl+2Obm
hKvSsaNKp93JLo4PitNi8dvt1NAwPrLiqkx7+r3hMt1NsUw1Lu8777dXL2EUm6nP0uxJVE69NUNA
u5GrFnLRCi9fwjirvpMuViYV0nxVTARmgaV9GtWuBrjlz30neiGOgpsu9Daje1tw4kO1Xciw0b5o
AEXioqRrj3AaBZo2P/aOjoSiAr7bJ7YEpCKu9YH0I+Ot/Wx7F7AEc59FTBUvbzVF0beBNbZk/hZu
SkpqvCUM8GlbsK8HcC4GEvTyof078B3LEzCeL2uTrm1oWM2UX58j73ot7Yye70M3FaFELRWUnuec
tB06dUrMD/c7VfGp9kGx/VsDqxPRJ60aUPIDypVg6tFexHf30PDpwYyDoYRtBJN+mcKJYOdiJNeC
56JiDdjjCt4+Gtt2C4/xV5eCN+Tsicla4HfKg+i/KQz3pOy4KICt+bVGmeOnrveTzm5oPitNnwUx
rZZB2cbUv2atBbjN8j8a9s1eW4w4r/PZaQytPmgxAs5E0fMaR/uk6O2XBhC4ZGmBfI1Vu/U55xnx
8lyk6c53iYVe3bWUCzEkvTq798y72fhLW1gNYUXPFFJtibQ78OL8nhJ6h9D4GTzvE9w/6mtpe5VK
lLMfqMCLEIp7fDzWZogvNSELVe8J/5i7b5YWYCSkWL/hsmdLwFBRX5YWYgPlac+hhqSUAUr4FBWT
5yJhMKVVtBrx/Z9wTTtGb/aa+H0xvCqxU5s2v6fHFrU0RMKRxBpv2eMEAGf9aJRnHuT8g+Zfi+7G
Hnqwdm2ySaIYM/W99XJkJ8wJQzbA8Gi32B2NZNjCmuD+ivcv9SBWqXZSSb0bjKxg3LPnAWgOISez
kQV56S5OxBJaDGj5gbeyD+NX7nGmblw4WNnW0xxIX9GGPH+xeweB/0eX78mWBfMsioxbuZpXzUKI
QcCGG95sKhc1vswG2GOplg4HAI9I4KC/22X/Hvp6a++snzOhrwakZJBGvqNaZwzLAYMBQJnRM1CY
bWlnRtMcFLOxV+IGrJon8VGvdtOu9ljk29yYGgPp6KiR64Thrc4SxK6/AHCs6aFd+RpV4oWs2DOP
LqBBZUzYV1XPj48/U80nwI9XJXwuuNpsysa/GoCczGbcR9NFMlSK/JcpsiID3NhWx0y4WpOh92cb
XQMSLfRetbs0zg6LkAdX2ykW3mZj1TJKYsLb9AAUq1hj5ZDDCdbnT/aWGyoMZ6mHQZFPLfQIvPgK
WRX4Kil57KjMOKKb4XfFnLQsj/W8ZMwt35xVo8Uax3x5EGVuCHdXDt7QL8dhML2wFhD54rh+5L9T
ROHdznErO95//uux4lzmMWiZyv17WmxsWYxDF3aRZy8dgP3C97y04B/IC6bkKobVN2PE3QRJR4Nk
PAXed1fdjGGJANcU7qS71FoaCoOxvYvoaxCvkN/2bAruHoQRvyD2FftpvO/yxe6IiYBXRv9Q5aJr
hYS2dplxFt4QPkTO+gMA+6veAnRER78AxgGcbIsIkRKYMtrmalJq/nQ2BXeUOXbH16Yd2lZ6YbjL
Z3L69er473CvZmwQguhU5+KCbpBk/fI7oDXdz+/CLEZOGCHzK5reWXKMMX97z2MLe/1p/4Oh74r4
lIqD+931JZAiTwJMlPeJl2iv3VIzfaNKR07MV2pNEkR8ORvbeEFItjpIzGCXP2Bhw2bt0FndQYeY
ig3z/ogkC/vBvR/fH0bOg5RkdCWPwaxW74ckqRFg09wivxGzxq+ohFeAjSQctHhYZCLAOXKCa29N
mR4K6SWKFP3vEA0f8Y/nb+qu1SyHRmFExhTLSmJF114H2Bkw2dugevhT//JyAG6Xgl78vba1jzyz
dqCHuPUAD53cK6004edVP63X482DRPMhae0udkpJnA2gc3ImoO/8m2rpSM/5IHW5+LZGTNMObeyM
3ayMpgmdfjgbp3+inPfEPoORCMyzxf1sMWKmVj5N0C1uH17k4rQH8zZiBaywgtT2hK2DjHVLFHlx
WhaB5KgQVA6c7W/ndKZp9sTy1aHgOXItc390BD5FayRSDJ3XI5dTEQjJy5grfD7Uqry3UHzMsgTR
k94osuUZLvmxEjQRoZ4i5nxI7Iiu5Fuu9r/YlwwNHDRYTQLlUG3gaZKTrKsRCTvzN6kr4kbNIn6c
AQnR45XHfUv1YtRCCjZGKu6iMRgtn5Mgo7jcSa4WoTFSrZ/iVHJ60xz6YnDY0SK3P8JQwt4mtSHe
dV3Rs+IZke5ovm7OAr3ywi/wgcsFk7zkMl32Gu3vsMiz2EnFnkKUAjCZiV0epfcZyV5VrqVTJ53g
T5Bt3GY2TuvgLc47yXBbzJ8ygubYTOxx5NJrU6mvXBQNYCSQx3gbU479qY12iXqHWF2c3uW8C/Ex
zVl1bV3XNnrne8H4IxYpAzVD3wzO5ltNLqUE6IGBAnqShtzvDzsaS0S203YsEfsNqzJ1tEzIzEp9
4jFGOZtc07wsiR403P73iHS4Unps3dD8Mw66ATO73JTD0RnK2Y+5Kz+Yg6abbO3G6OqKqLvGNwlb
857r3rEf894zljtXmdKDRHRKPBbSsc3+4Ejm/zHw4aLRWRBL7u3OPZawVnvkCnNAL9vmw2b6g/XV
pbK0XYkPffLuRSmMqGxf5oofyN6kvHcnhiisWuSmNih3my+1rsk1W3jm8+HOePwNOHugVBFsmO9I
aqvPmltCafO61ZK8r3DaCV7IfKaB1JGceohhfAC1qibNX/a9LispD3WWU0S4242N7o81Lu6gsGv9
B7g8qqDqN4tSXl6Ecl/YvKqDw/WDOGvl8jdBEUa4ybsXzpD7uLknovHxovZ1fYeBqLFyvXbU451t
ZGaPRcZACTpTcXUyPcawconYVOUaTsocXeR0KEAOrwzIC0tvjOasLd4jzGKBoBNZkVEGNwDrMzMk
Lk4N3vacda7K+JqAAjEDOP8JurVLrZR2iguN3sbTb6md9vmpLNbLYYyYcnSgsSPRTA3mH3ugegu9
O+am9343qJrNy0SmVo+r4ArsmgxkadGlqvzVd1xuorhcNE5Z0UacZgCISD3Ek7npDPRUOhQN/srF
ehJBc2lh2S86NjNEo4Ov6xghM3VLVBlBCJu3358+EQDdv40ZzdeXXglJDsM2YjI6e3M2tGvOjxQH
WIqT8hmzes1IUf2SDpLZoxhE0OotWxH+onUXiA80Dgm6gh2Z1HKx4m8VDX7O+/KTE181vL0knww2
MuEevp4DfFGKrKxQYTnBAM5/hDJrtkfojqCkvLbWiQonCKJIajfFNzuN+XHPBLl1fdfP95quScAH
hU6dO6iI4blotIIm+1g89RW/2laChVEC1Pao0vJouwVXhf5vv4aXKv2CCtFLujG3FyPUMhHKz5UO
n1auM6JR6xuAiAp2ks6yPRhZrKYmwifx9ksX3vp31dez15XArE35ETJ7rAaj1+FWz0o1Dkzw8uYj
7wXjuWVNFlWgAXOUyWGwODwKBAy3+5QELRXPDoIcgXWiLbDEfM0GStnQw/hoqPcREIWjb2YVW/rF
arQUcaw0p3Wf56PsUnkXFhxAdPG4jUIOh9pzryn++wn/SXClpOeXPDJjRypELhuA6oERC/rrx5n9
QBDO08I9KrYCO57taXgJ88vGJ0GX3zgzr0gP9Nslbfq3mkX43P2yEoM+ZcYiVBFOAOQ4iTY1noW1
WPy2wOFfXWKKNR0+lduN77AULwPrJWaAuLOZ3APCs8t3MJRwD2Ji8YIAXBg2t5yhkO5ePw4wlpNq
3r3WIbTlbsD11I7F3T7/lz7xKqlQCKwhXpYWj/d7Ng+QZhKKp6ISpj1Gq7o3kh4uQFB1aCgY8sFs
T7AYGTVUhknJAuBLlLMlFbt1KaToFTmCEugfMMasoJuJk3449vOcp3ZCheYY2M6EdIc7fkxYenk2
Gt+uo/8AIigPtQexsNtdXZ3ITCYYhJ6D0CWz3//Lnb1oWRvYNiBEgjxemIlzDBoIjY/OzX97FhPe
6idlFH0b/fo7oO1xRv5N9HrWz28W6G8z0Y3G6zuqDhtlfpzVCDe5VcxwXTPQ0rMXVZEAbcN5u9EY
ySCr6eIRO/0Z5Vu7aNsj1uqBjkMoar+MEQ4sSk1nvTrfHPCRJd84JqdEGs1s/Qb93eQ4U2Mln064
wB3cqm58uHH835wNpQNnL39kqUgvGRFDzkmsx1QjyHfmE/2ZrarrnbDofTGzjwEXL+tD7SqbYn00
vwDuFuIAP1NwfixFADUpCci0q3Etb/Ka4pnzzLY+G6ZP0VmBSustQwhcxEWyYzZgCCeyNJpryQV/
nFPz0Z8zq56lUtt2yke+MxeY1cYdMMm+KsFiVtyNfWNtgtzUpJBqX+o8H9UQVcb+ILOL8KEPBYFh
wGgO7LlmnqhD+LbflopeP+WooU3xUdT+LwhnDSeTpHSOd4mctoHmdhzwrZ4BTmLzjEImtXD8sEyI
ZuVAraiVDS577jYSdzRFOPGQY/YeP5zcz7i1eS0MgRd2qafmaOxzaxRnnPHjThAOKs5BqHzDGI0+
P1fmfzim7RdWpKy2WuQXtPBQLgkWzxgUIZGBCaHxkr1asgogyJA4JkUceYbg4M3C4hgN8Z3VpMdP
hu8D6t+//aX2fYGVRvAPd2aakLgoiNAnx6lo0RWWLy2xjyuJZVp7DU2z8s2Ib5f79VbSwoq+1sY2
pGW7V1HweVun7GFmGQ2IR1b3klwzT7K9XlioxSrZp651ba1nOVjLSfS11fZ/UvemH45D+BAUusVF
2fX17onKkhkEppZttZwoHZtCx7MNc8GwYQ5b08OdoqqAM9Gq9vvpN+TkdwSBsRuMT1wSjKpCW1Uj
WcuGRZrCUUzn6D1u2ZTCqclWYNXpVNhqccPkh8ITWQ0zFLqjEDC4KTQSQ5bOTnBOJY7ZDMYvES2I
wJ0UP0FGUS1PsqtBa+xrD2KFZZlDPotIpfG6aUIhtxsvW7kWEa+Ovmv6HuWVgOqseVI9AD+6YA+2
ndYSdWMGRA6yeXkmxZALNym2FdIYvJx8d6bws94d9P1jivi2YFgv0Lc00OpvijEZS4lR9X9Wd5jl
7vSh+lP7lNqcdX8VQ6Izwj/IEKIMEe1VJUlImXCgPs1gKihJW4Fe7pU4R+Ml2Qcim26/IzGMmf/w
YjvR9GyLVUKZsbH1QZbDzXd+iE8kAYGiJAUDYvsTVpIZGTd5iPxuioKbDTqaakgDhDc7n8p8ub6R
BtY57ujBmzkCGu36mLFsozGEn1jP5gj5WIMRMbAj5OHUaiOHZLHFZZku4EZ9qwKnqrgARU7SWo6x
8bBDN2BX9ZllRM28dKjicVyK5eskFFuqZfgy4mcRK403oW1RhLNebUlXOd58uVljL0l9cqciYpgh
dkcWAsoPA7UZxYL+B4U1utqlDZS4S+KT+pW6qSaUE7HoeUYsKNgPsgwd5zpWMsTrNMsmOvNpTBWh
BU75w++NavpKluwGro4RgF5Tgo8jYMp0pvaf8I0XCzyybRbzecryeFGUCinUeIwianqlwWFlFx2s
jFtMzA0EXF4xR5moJ6pr/e59UqxU0aBHu0YN3+svfBZQF9zFJyWX9JasYqt5NA7IeN8xYK/Danoi
JTj6rIC1REVGNd9FIzEN1DLrB7y/dbXJDHhsVJ985L6I5tlkbcVTlDkmHwfFVoXaiYETz2npsGkK
rK9jD1iFlCoh/IG8S01XUJ0n+LpRNb4DvqAplRtUxym7j6E6NgQ6q9mcd+2H1SucKDb2XSsAJsm1
QG0wakDmUO0wEGeJGLZsH+Qp6iBIZGaTxNWaBLy+oPihjukj3gj0OuDo+2eJoJvbSy0cDWqTdgUO
y9DwQDcD0S4pCQ4qDRxOOmTcsrNqBZ0hN4WRDW1AOueMbhBjiUv/Dhbc73MskJEdrbdQwHSHjbAj
ywklyXuhyK0KlZv/qifNZ0e9MEbyyPc4jj3+2Y9C9c2BdTKn9zzyfWEpbShiPuMLl1I6RJ2r46wk
UHTLpV7QrmsczF2tU9IQk3HyW5XOkdgRwu/NDyjMm9CNkdib5FPxUb7BlGWZjANABjGu4JmB+DeJ
mco6w13vdpq8kSTGU8XXuWZTQAPXpisqakZWGQUX/fGwRis2yHGxkFWFnHYFwdtmVokkIT3a47Pa
e+5TtFfGP9/wk3Ac9J3eBPhv0v9ifkFc4S0AGtREOhlTh/ix3WjOOuXGUebUoZCVoFDH/OE+YS6k
5w3v1jLS/hhlZ+H6WY/AAwa9/aSzB7FyDW341FrngvDsGrLTnDu2Z4/vabSGT+vbYal6jgs//7Ei
3a4Jtmuouy4LVloFqJqMc5ZLU56mwRZCS2WfHxl91ydXzkFfeWadKbn/9OFwdQTWaZ9xL9po5osY
Uy4dtbBut0tkQYkqI2WBKO34He7vuY6TZMXGOfKtQ4RMLQh2p6AxHGlmyRZmYMnYpkMa4TUzR2+D
bCiOjwCRP9cpZgswkJo68sXnFsQQMoF+IMUCxBe/2hQkD/dK+UvV2jnC8XlGBkiFAc4ezT2Z7xVX
WAJY7adxI3fjhc4SlAPpJnmbXDpl+yNPEj2f1TAvRI8x1dC8K+Bi6Izyf9u0G7UdVWLPK7m2HMuF
50FO7g15O+1XMb1sPK43A6dKSBRwArrq1VlUxvat7HrZ3A0+g5h9k6j9PC9oEgbRsN6tO88zD/CQ
ORAjiFHSipVmlQ1V1HVG97SflJYf0hDtAsZvo7crf9utXKlYqY6lIBr74YM8rHUuRsqIUYzETr25
29IsIOR7r1QvK55rRMEKxynOmy7YB5OloPHQt3DB8bD1tkG7fgQoJe8FIhMNYGSloVLEYzT7qTXu
Fmk/5ikLGan1udPACSYrs4iM3CxGVzeCnI0aMlg7NeerGpGKPGd0926NlxvYIQul8EYYdHpmU+JM
JhInZZ1X/u5HgiwdkTP25yv3wQQPO6kxM/0FJtcRYCpSt13Rv3GK+vhJFVfjNg+0Vj6mepYV+qHF
ueRHe5PcWXB8g+j462uSshdbLixaM+nERafiuFXpZxod21RmhDL8/R16YqhePX7qCC1DK/U9DAMD
nDXciAi8dq/7tOgYGO0UWxhQKnh9lJp3z8/QhQghIXsTPbzgjfCRqXnn6yv8Wagd9r8hBit/7Sr4
L/E5bySBVrEQ61a6i8GEDe6caz9mpB5P1t4Go/1T0MeFj+RezeqMr8Nl42AhQTpdJNkZPzeNoTWT
tdXdENdPy3ObH2zVjcMgoe1zPIBqeM185UcikmmbviKBXVMnmavJ5LKBN8Ew7rwhBKHYZ0luq3R5
7z1nhpPVxtM54s99PDgNeeBWDc+V0U4PtaEzNoJVo/52q5firxdIhTR/on0HOz2uBACpBBgHZkMv
JsSEj+rUZPlC97MLz2jVPMRymiPAotPHiCJYOWXj3dJt+aHVsxGj7tq24qQHnW7Bu5yuPeNW1YkY
qY3Qg3TAflBml7Dfc54Hm7Us05RaOwjgnCdy3izcNJ9AQokwRG+HOaYlcIOAgiT2dmz3fnx7l8DI
+HzJWWM0kthL+knyPUlhTzcZl2s9L7EE8uwxbCY6H9fVdsFYfbmY+1k1G1h6YQUOPomAPihutvWP
ST9w8exw7UvPjoq7BfjLna/VRVB84cTAZ3Mam+5Spsx6UFeUH+qeWAfCnIG24PNC8TVE56i/Yvce
0+ROIaSlR04oBHIQe3FHPrY0Hw66fRAhFkyInl+P4lxKlOEfSgvCuxurDfgbhhOH9PEgvmMhShaG
XoqicdqpP9ly4KESHOsMyqAt/HasO19CotX/L2rJOBzAjSZ0VCDE1XBOVtjtaSfmIkzePJJTXXQ2
xHdQbX2DiOC+azukxyzansEymaMMrO9ANDEBQmY8dRNwHtO6A2cX38lvGi5MTQtvBLHC0U43f5nj
XkZbuUP8vO4JLmZMmB55cBnUxaqVbI3/6LQIN1LXIqE+zNn+5Wl7fE7kknf8uLy0pYHWxHFPKByb
IuBlJ8KoYjUO7jiETeAm/ahRvCXi5njFrNCv7jtYvf2lpyvJ13yzntyGMc3bhc8aBeNTn7xrpYYL
Fixr7B+ioItVu0w5xu/1goQFdxepZhY3tWkSBXvvCFUDQmzxhfsho/MfhQugmLKxdZqpfu2mfRd7
0gsH1LUdDm3FifMqyDTuacg5m67d9kTEaLbj8LyKTRcUo79JYomVdaWEdCTscAEI482xfreRt928
fs5RS+GWgYU3HzUEfivBTRYDqgL8+Huu+9BC+7pHsgUtWbdbadNDqwlh3g0e1+IxDUkLyAS4r2WO
HWYJYjFiqBQntcbGU6vyR5dqrx8XDuc6XB2Vw0fqu+1we08MEZT3X5XkVEXzyWVr/ul5IDxY2LgN
J3+I+kwgHFOgOqp9pPovwY/IP+HNsu7lT7cL5OSJukSnJ1IEqR63HulLS1G4NIG5U8adkFK/ktEo
U2CX3Krs9FqAuGzhQiUmrubSki7ZbeLc8gaQqYq8WeGaoKJ07RviFTOsTNREDlhJ13ZbefPJT3tO
c6+6LPpJimXfiUVOgcF5FHk2JApJA+/5JMj1Bc5fwr/F1Lf/Ywm/Dtof71zOD3sfUGCYPIjYxpdL
a1NG8U6m66k/+//UX8txx1T3L//S4PzPJ5xwAT0i9udYIVkKP51qQ8WNYQRn21ooRyNlD2Iw/vM/
grJj7s/3rA4MO778QxxLzNjXXkYTZbEqvs0EUcQ7dmmq00HaoriEY/yIuDK3gNO61QSt4ysZF3NB
vao4tHpzSohwo0YCzzbo+F3lbuQupQ+F0tXwUjA+/1fOOYIqFJh3JqHeWfizT9010IcXfCglSMMd
8o/CY0QzC/h7d90mzqzfyPY+oYje6s7EjLrH3Ul8e99y7OTie0UZLWEY9+ojWuWkGUzL9aZJ2F+j
dA8BIlvJM5Iymzjhy8LIpk4p/xJYg22HKelaDaZnfjYFBHXV13O4MzL+2tO3NGGGQFh7ctn3L8mQ
xexGnfKDjWPB7jWvGyj8xWJsXm3V31FqqCClD4EHsTPIpSslcKEhJYtrZL3z/qlbwyKx+H8C5EZh
sSZykKdgHlHfWg3B6nW+oUu6AVdXOukmcGg4NZOn9nODCug5vPiBRxmzjEZiqiU44mdGT3Be+Ozd
sFs0J/PUhajoMwB5yzAzx7p+a54M/SLra38wkly1a72/3gHUOjmG/Tikiqf4GG9ChH3Ay1YHP1YS
tSSkf0Cqa5ftDBuUWpCzgxt6CaZAl3vzF652XbOsTNG/qoeooQ+irkFQkRYz3in2j1V2PDYNE+wh
HH/hJ5sKhEqUfJlYQkLc0vcDYtycBCzaLo06gZcpDZSX8tlaUCSa1kl0kJFo2sAvQbxXO17iqYRM
/Vz84A9B7zcWkSlLUC+XDtSMp+4c0R2/bizjUY91YKULybQN74GokvwJc0Brga/dPQWQsxrrF89i
xtSAmm7uwh86+VlD9CcNTiYNUxEuABqz07h86AqDVlptUs/BvYt6CUUqjBgSwNcabgvMl9WKReSY
deZYwR3cX4ZdP4L6OGJb6k9VPeuj0seSGtnNpf8GCdp9OYWKBa0cRjrA8bJt64KebcvszMRpA6kn
wlEYfifrgkY5wyVmqtYwUc1zIiBwnKYtgo1PSqRS6rTADvE57gdhIjsEd3lORfNCA2Jo9sKzx0rc
6XvmZYX3ynO5uBhfCvtK07vi6A4dBZlrPLU3qNo4Fkl8wya4RmVc1GApxKDv2gbLpCXsECt4IU3F
Mr0n3wJuzv+ApSeJUkpPzPTtYwMMKDk3QA9Fhl9ZjKar6Vf9EdGNtv7B4hVzUUX1Uw+cOvW+TWbL
ACPoSXFYSFkrS1kurgcluxTxpeDtv8umy6HGfmL7Q9HtUlFQlmY91JsN5YW57TZn/HkyzbyVcozB
vv4p5a2DH975pxoCrhlV056PZD53UXPxmPR1VsYVCwQXpJ/bVjy2iU80fkLbF2kfeNTLgijm1hyX
YV84f/WsN6HwPUr8hqbE34EAfv8NU+uj4Mlab19H3e0ERAfkeqLbYeTT3NI2SGSCBrWVA8LRIPMI
U/W6MMkKTl0ZDda4Obo8wSSU0TWV0pbNFzzLJe/eTyNCHdl0bDKSttok3mSD+RTHDCVIUjckYb+b
IddyuH34MKzPnvyPaGIBswlk/dTC00/M9DBQ+MmIchZrEZ+988aUKDcCbfBFYDQ0F5VbsZDTy23q
TYRaeIdOOVSjPVQcpVqsHp7GdaKEsU6f0x2ixiEMjC/+tWkAguaObwmoH/+cD6qMRiO+lj1dQA2Z
UDMH5HSMZL53XmtkphdaaguUPTPq64fz1twyHg95Z0GQNQtoAPSw+FWfPgK3G+RgHKKfGtpSJJoN
1Ql9Y5wVGOXcUZybwIZTsbY0R2Ol7dkFawisS3ROFuC2Ksfw7L8yltv6mI76K7Y/RbbfriSPvzuC
9kSrg8ZjNnlYV2yLYLtu88QKecuVn7LsHdipj+HBTf8wCzUfai+JSJY17A9w27bOXj5NzuyBJy76
/328LmgUYHSpglzosQKBr3Cxhi0q8roXJ975c7dHV0tjvpV+a8dwJkhhoTtpk/ZiqXCvKKS4RK7f
MGxMoVDhpCSJ00dtkXXDA0BKptoI78LetJ7j/Ys+bM/NDOcUxPARBSuTPqDCOgUPXTXjeDdpYmoy
z625/pfU48lSSg9BaZP1BYZvTX779MAtjeIWVVdo40YkvZ6+IhVWZ+N3dvKixBlya/d2eXi0H0/h
IhaFOO0zZB+bcF2CD+MdhJJ81XJE6B1Rdiz3JEQnkzpzJXAymYxuLw//Xet86UUS14l8veHDpbK+
fbOKoUAfHWABP22hcCKEr1rv91ScxmxSCH1Uf2wlPci4No2m+rp0NHBIIPlAcmqn8oHCUM9HDLbn
pMTYh+MiBUEzSmxLn2d/euqCUHFntsleXj2fjqyx3JLwd5sj9iBdjFJspf6dGA8AbWAcodUBXHs1
yglZNRp0NH0hixtdG/ONc2t/p5O93xmcwpjAWjZWfTYsrZkw0axgKIbyKeoI4WsE/0T4N1HnlXGX
288BWex1lzl8djbSqsQeXaDRop8aOv6/BwtDw3wMsZQvbMdodOV5Lz2BsI074y+5glp9lsL3axLf
OzkHGLi8y/pxPrwY8SBmYTSRCOGLypOMqk5pTr9G8tOOfnUV8z73zz9Nn4XSTb/DknRJSNi6jP6j
N4vLuFsUCR/BIhOiunWqHet+yr6YduNvOEvlIxYsmmLTfSHfz0GtY054ih+QYcuBxQCC+w1KmiNV
HncB1tWF4NTEozc9Zw1KtL4JzCSj6Et0IShC6+JJge8cawPYXzvcoV2Qu5w3juEjus2JOEag039C
zE7MiML6aKukZpjmd7jlaDS8LS3tyuEgVQfRiiyv8pTXECR4Iu/9hPZeG1xz53fhCOyqcOCQDq2q
DoUbDljpPH0O5H1XzfOmXU75oqR4MHEZOGQEy+I2p4Gj8UNQd/Bf6lm5pUOB1nUpY+STaLKLkcY0
dKPuWEEk4f3KS/7BU+EqgCuF+bv9CHs1h/BLenXpwolFoiI4LUfn/KhAzVyuSB+EuKeJiMnOyxn5
vmEDDB0fwozZPYpgppizzjSnAqJ+9yXehFmi5Rmc3nVgX9pTAquTk/G3IV5Wj2GspGAe6oCqufTo
yBBhrKXtgeh+6ehiuZEY9k7UAs6ofj/lwfb/ugxH+0A31BTslGjE71fM5dJ9G7vw8T2+b02tf+sy
ElZm35q+TQtl8WXk5Q/hh/hgiWD2hVueAbfHs4mQz6r7iwfuCBdDhDtLtV3phnKEpy1W7DbRhy63
fWVZsFx6/InS5frkGq6jF5lKKI8NF4Z4PGOq6nD0hhvCk8YiFvdiLVbYbZoHRosNHfWJE8+crUvP
blbd27Go47F38/BB8qmNKOSebw/M5Gqtu93zEdtJDu9y8+Oh1nXiZCDZBhA2ngDqGMYdYHltpxAY
ojNmi8rnc5pXpySZnO535LAfsLzZlVi+pMnhQAMLkRfGiP0qMW99k9Pq84cZC5XpQxC2uYwAUX3e
tCJpheY4lozohHHfEC3etkpSAo3MAV/9Wlc8BKNf+6eSzjgICET6ScrpncC03OM/IFSpny4+eIU1
wz3TXYvZXsnz5rRYzduVvRw6D/Nv1Q2SmiSZNFLvifrYcl8Nqu6wUoVIIL64ksaAZIJwdarENkqf
Aw//uELhVhdgzNGTJjUG8NTMks99DtumveNbNtObMWbccdLw5WAym4zdPBNYO6nGulbr1QYPjLDM
Ru5TgeLwfjsOEWM1tyeGElSRzEMZK5aeIQKkio2n4mawDK2WXDk4dP1Z4gaa1rwVu8Y0AsSi2X6K
rGav6+jO/zLZ/DXTkju47MY1Q6AMh7Km+RTZ5WUdzOPp4fLpFy+nEQ0mH7NuUq8HP3r+jgpfu4ec
Et3qdSNwiarh2KZmYTLe7EA+ZM9MiJv4p0sVsvMcV481tjoc7mCg1SLmIIESwzSoTrko7JnbiISc
dDMjXQ/G3dMnYR5960WqRYpjC+BtPyjtk8b5/A7de1Dn+2eaolnq7MfIc3gb3qqv2v2tad9IpSji
7eAcvSeGXTX6dbFO1prGR9TKPom4lVP3btaNLpvkPoVnSuw0OaAsNphDFHWyIzsyx2150Yxaf0t1
QcY3IT+sv7dcS20FicIMnzexJjrsvz2F6spBKlJsPTkf1AIrPDkFbj2D0usUzb6qcGLoNQPtVnIA
zpWn4VotTZqzvmoS1QDOXC/0TfjIrlCPIvAn/08nFsRMtInmv2wuwvCjtOdtvBlB3ZYR3MKReihO
VGDhdZIMbBtqqa43UPqeDyhjkrc1Yka24CsfnwaOxpXiOkCBmjX8zBvG7e3dtZnJi7iKiUnq5McN
VqjCOh4cWlZlBbaeHm8HEUraFJet3YS1r8Traj+ncY0931bDEp/y6m3NVXRMOSf2+qyAgcptROqM
nN11qalr3IiWsQIqa1b9HxGMAl13XJDXs7Mkqmzpb75/hOBoG/9MJgkr/F1TNozxvnt5xUvP1fEK
AWXKZuKTkvnCJX1hTKd2DDK5lVKxY7B62HqVRFBzTXLKZWU/NiuC1/HNW6kXyrwhKGm7SzQs+ZCq
oDg7YGOcC69j1sjMS+GS805MktmShY0atvQNLDKhiLL6ynJK9uy3ciA8jbJ9Uz5RorSX0T+IczCA
8yX4uf2PlV1HbKco/5CNfgq9zmNkUFdnhiuOSuQy3eEaO9yqCsEJfWC2Agd0pdwXaISs4Vd+bcWs
8zRZPObTJR6hziWAeJ/7PNa3PY4cWARXYKYo9ZEFKzy8riYhSE4S94lHy7vI2bbAN2Jg13D61Cv8
zvDA7r9VR2Q9drp/g2BLbncbQjsKa8qfUxKZZzuqlL9GMp8jJhulAWH7T0SSeIMr1BJblza6pAuJ
CZB2oCUMsrJkRyBDpPbSFtIXweVJ5Gux9YovRpXMbwbeplrjq+vwUOEpHxfn8atrMrd9VXhW2hf0
YPNj9nuWu5oPwmGlK1EI1IHtmaPr2j3T3XyG1216ZJFyxroRM8KdMToNh9K4DQnRnVjqv0V1Iq2e
X/LYLDO6sbNjKrwP7u0AU4XXEWaRzqGmiqBpH+bvsWO1/YYlf3gYxBuUNKkPhkaPZLmdNAybkLgd
BVoDj8rjzCpJZ5ioKsU2msgFtL2ikUABFwpD17SuUI5MtkSHiCPhbGZ6L3G6cy4Fm88PSvc+DwYP
e7ewru874AAcCr2WPVfNo9kZPjQRdRaHIbjJqJr6vydQ5ux9HpgvB2rsZkDhEUxHt09KPIN7P3tv
ewZaPZPqR6Soth9Z2Quxd4j2Ijtv3/e62SpuHkSCPeoC3Ifr8VBWAiSUiDJm93m6dK1/7QAXXLNC
0WDsE1icZbq9R1NcyItjd4zlJByqKG3B2wRHnkMHXqpJZnr8VtK3UI0QW6mNN+98DVp6HRARQK2w
CeLWNpffhzkDm32UAYkbmKHcETMPgURv5dOC/C2Pt7f/1ffoCD5n/xvcz+/GCCP9uz/X2e4Tj2bC
pw69byiE4opl44Zhwuni9xaDZZmH9HbP+3vsVVLKVCMD2RZq/f8zy8REt5aY+xokyrrq4+G1OMrs
GB7R6sSs/jGAAOzRuMb4pua4Q4MK6K62ciHS3LiSKdbu9BZRRXJVJ2qlA1ZQtFqCUpP3QQiwqec7
2dSwylSVYE5HXHLxZBJeahOmsmgwhT/5Q123j+RfLVhcH8tmckmCecuYzo6qSxWEM6hfvrBuVMCu
p9KNJq8yR8nhxlcT2nUtujtbWGIAZbAo84UD2QbU9y3/n4nD2d6fydC5PxXRGfPORz6TCDjpX51B
sNjN2SjryCVRLR251PngpqopexdJuxJhy502YuwWPwEZXXBlkDivZz1z/rAmnoue5R2q1fW/Z8S2
cBDEJClkLNVr2SKN69kBmqiafyhULP95d3Sy0VqE7KTceX9ak9bCMvhJx5UH0pC8r6a4F7jDbTyA
NrxdLzgFr6RB6dml1EOcwIc4JiWm+6vwbasI06zC6yGTMzGS+KV65GYILTYDC8bjKaXWlYJrAGrU
xsPbqYQQrOD4w/vvVrm6lFWVZ7CUTBBbuNlVPFhW5bGSPvqQv/EamYo7jo21or2VkS4csZt/rGL/
oUQfUp14eYd5IxbKLFMje9nzvCmwwC9j6x0jLmj5lLLki6iSI53jvjJIr0m1NGfyJ67kYUeJpIyT
GFKAG4tJw+OS3TUkg/E7peO1+kI10jIdwdbdDDzEvVq5+aletrymtRr19Fjr9BwLlp1mKIkH36il
Jwtwd36VMS1ydE71biq/jHmYcU74W4ZPWqPdlHOx8rLUdCJEaJM5PSu233dbN2esRqBQL6N0VS/i
Xqu1GbRsF2okb/ks5943l3aSWHRx7NmKTk7UYiJQakCDx3Aq4wuXZsbcp3jUeDDI4jAZCN4MBCvD
+Uq892H67iN/I8ccakKPBYYdFu7Id+gjW9hLUsGbCJ9AX59lI/3ZpvYfjsUbUW+w9EAAL0g99Wl/
Erw7DIH8/sA8x0ZKpI1v3due28JM2JkB4aKSiD0wQz0bQeJryoYvf2zqnTTgqcwLcv5hJlZOkv33
V4DtTWlo8ByNJ0nAl96AAVWnbvqbtr8BwS73+80GpCLrxVdc3Ai8T6OjZIHzdy36wDh0QAbpwdgx
TcKG5ZAWxzjMIiU+1aVJknY901AQy9ouSm/vEB5AMSw3yETfzrMrg4D//gwFegbccTz9QAd9XGP/
qgNwjeB4G1QTYhxRJirGxNiJnHzqQFHwo6kE9+0k6/TpX/Q1SaRWjj2yJX2Wvl6ZT1MDcFSJdyUI
KduF0DP0xktmJctIGfYguJhngkuHDOLLeQ4Cu4g3mE0uJfbxG4oeWP7/9pBIpM3aDkdMo59Gr+bV
ghh3rVsGAUrb2NxUnImfHw78jpvhGIhbFp9RWrc68y6YIpqUHT7mdGyXlHzOxRWw128LcyJp/Nep
IZBQbyC+jusJilxVFYSqWMrEoKIuFKhP45gwqO1I5H2ZSr4Ju2j8INmr37MzayFvRdDlggslWWQ0
kZyqhyjaftiy0qLE27MZWmX1FKwJaPTE905o6VIYYCcX4EOEugk7q5kJYj1un6tKL/pYT3Cj7Qzn
J5FwWIlyOuB5ey3FacMtZqvPVLbsK2bje2l07Y6nvM9MP2wdAdlF7K6hab4jOwMJm9jpOIB52lwf
Sh/RyFJzX6sn5K4b6TexQguKFJepV8GhD72QK5A6pj2qOcr0cueL3aoRy4gq4FNqJdZq+Tx83EOz
rl8vBez4oAlGlb1Ib2tbzEHyrCQLAKCeaMK2Sb576hG66rxPgbzulVmFnovMgTA1dSOxa7AqLa1w
GRdxdnwSkI9g66+Erz7VI36KgogE419zsd/yeyIRr5tL/UVX+s5mETbxRP3Jafa/zvMZLgXyF43l
QbgHveEv2V1nA0Sw/fjqn3halmwiiwX40AUYvcRmb/229uXgRA6O1kZb0wk4vYEh9plfKJFYjifJ
gunsZ3385flMQVZivhTwBqfkDEfP5P71eu36rGMLBURShaPD7uxi2fb/UZ0AUGvphbcQny7tUDX3
KmnP5ap5r7O7VbK3iGASH0KtzeWrK/noXQFLYBEpWgQsH7tzwR2sF+a/CYrMvlTYnqL5jwQ8zJOj
g6hTZfn3apfHviI1pXrswQaqrRk+A2Ye+TPSjcYXJ1UMafttf4vmx+9nQI9t5bpKpXVEgyMFw1bi
b6qXrJKfpMYQuyfFwROEsurb5SEbwNRc0eFGvmdZfVROgwNSum93QX1ERBioVuJwJ/SUGzhDtEQT
sFVmUmQuo2DLnBLmZzYO/vnk2M56IeuP/DHVVImElHzusFIV84/V2xYF70mdRQS9Adb9Y1jeOD6m
Jy+Dj9n8Vl97V59vl76yMB6epjs7fy5VOXP1FwlnzO/0ghA3Ecxa2RY05fhnZaR/yVu6jtcYHxCa
Lhcvq1dRg+4mpaZIiiJRxVH2SnBQGCWqsqmbNG3odflxO/VsNLO9wP1nU4CNi8mhLIuFUr+c7/Wd
riXKXuYMNCL6I8PdlfNj23JT/xWBF+p0/MhWuQNwl3SXLeZ/BngpHQGifcMW2ZpYK1xo84rrwZ7q
P/9crBXFUKNjdT+1GCMpZjULIU//5ywvpyHOoQk/SQ3qWuZjfonGy2vKpdp/RRsiRcZs4fwPQghE
HeqyH3r0dUTjBJ367+qcRRMVU5+xF7SbD5dyj/AZy7oVVdVn689ei6MHPl4+zQ93FcYCuumEe00a
toA7EYmgOS2KOwHSS+MeZfWHg2d69Ebk9hfkXuM77n1mcjYz/4YZHHPNtGCXZE+3FrG22Ve7DJ97
xQem6kdlDyy+uq33Qu1GOB0BDmZKtbVH7rIPNwzrt9PIM5hNgnP54aD0wOAUQIeaBIIQS7T2Yjpz
ZNd47G4siFqR7vPq3JJNtk7ZmboQSLlcgNjAgUxWWW7NiF7fXOXpFYIPHaDAWxi6UM+zQXYztGK7
wDXMp9Vqy4l2gpbIrWNqVdxUpzyuY4ZkY2+nhlh/3ZAx7OHN7ghWyBURhuYB0VCSz7wiAgGl20+9
XaGCwnQlXA5FJUjH1Bw8S6Hd9fvZ9qFKgOJnBgUgb8Npev5N4p+DaDWMiwIEn5u9JBlYgXFjfGKg
YJvLBGL0lhqGONR8/CpmUVFSkUV1ps5KTsw4+BqQuRf8SKSc8oXtjQ5cZDJDR0+n0np1HBqWGzH1
cvfzNnv1CbAQDjkzfXd19OtAT81+71TpXlS7G//csIwqHIYmqFpjFjXNAEFm5Zxlc56UgfTxTauS
LYv0KDybDJuA3ZMB2UsQvG7zT454lurAEOp5ihNGBHGm/vUR80zHkgeH3k0o4ditgJJHyrZoctrn
C3K8Lm3AnoGboKPNYFFY2+7fF4Aht5FWPrkU+HQVMXoB214FQjZGgZoxSlFtkklcIoxI15tXUjkN
L69I49AtHl2QeoZkuL4OevkEOsJ33J8VaMysuQkJ2kEKcIRC7fJ+XtvcMzSsoBg0BhG5ZpPKqttj
S3QpQ8RWYxBb9uh6mhqUznb2ftOTP60rBfg8T5HR7EAE1+M3BRPsPboA8SkbmCW2IoqnOBuciHX6
9Jweyw+l69qwgqSoHHv/uKca7q4cXdVu2uzvN9WADf9dOYP9j2yb8fVrQl/sM6FQ7n5XDbOOVIlu
ayb6SjCXSS+yX4KEDum5b9n7FobB6Qr2Oa4rBAJAen+RmBADQaXJV+11XKdph4F23On62KQnDb1b
9rLRM8xIbUuJu2UiS8EvNPjPU5GRDbWN8O6BdRYve1uASRy4MOBKDQp8tz7NEVpw3YNLkcNzX6N1
L1rub72lO+g/sxHXbJbosDTgt3tdBOS61I/v0VIdpxrla2TAR8rzlwQ0jN7DlK4WXOxOFqzfO7Z3
pmseEF9WXlSMC5h9Mxlba5S/gXoQhACNBdjDPA8V+uJKJShKq6ecyJ+TEwSQvGNrIROLF1rnHk3A
0R8HVJSZFKCQcWpH3G5sIbfLwwYqG92B9umYuSyLngytE4sAm9btdKi+AM0znAb1/Q5bfK8tVnhT
uId6NPPfQuNbeP39X5amlXkm7jSwgHyAIEfxx7HR/Ydfl3E0fpMLLM812UJ2A64mmaDQ5KzXgEaK
lPHrNwNKKoX9BVarhp/LTMNOvnJHYtg70dYIN2UpgWYH+NjndEOctwT/e+U9XtVCk0wN854Y5A6T
CKebZzsvTimh+XNciK+TpmloQBFoyMsoZVaMOGcjwYN9pYSzyDXIY2YgYz9U7/gHwTxxXBvlece4
i7mYdUa5dHlzK4RM91KSFeGnXHHRNl6v4fHLDBWQPeFWzHl2qzocFedtWsN9zONY91SwLdeB9TDC
haPc5zFSAol79oOhDAuMBPEYMHbreQihY5dl9Gvou1kazDUQSYo0rOhWsWbBIGnuTTX2ZR/QYJv5
tsqIS/U1grD3T3FehkSAbHItCXH4XYpNmqHZFg0tFMV59n0GGe8sDZ7DjuJGPI5vce927L1Vzobw
nU3YXkXHiP6M9PAgYoHRD+6hyqJsTeAIc+6vBWanhOrX0S032K/xmNoPUlUe9BcePRRecH78njRW
2lE5GJeXsFbuEsci0N5u6AWOWuYX8gQsP5UcnAwDzwdOs0DNo0C0kIBz7OMsSo51R43HaFB9uLWF
HDY6Vg52kYNe+wXoVlgPneDfz9VsSKV6OiyqhWGbwnJM10sooK7QYXRTMQ9WJJ1hMzao0ghbRQsF
Hjya1noUDJZZaAU/jmIk7IyjJG75veM2PS7uT2oLq7ds94OJADTB3+dqznsdL7uclmLW8PyA1klI
xakIKMv328rd95T0qes1okTM3Kn9sdDOjDzIJEDHzgGz2srqYxkskNsgZ5qCNXdWL45KE4VColhN
iO6ta/Ua/KgTw9lEj9g2uCCVHYJ/5L9FPapNpMQLl5b5ZafgGhV1PTG9d4++iu7GwwOKhrAqYHRt
FQg2/1MJVceuIHhaIDvsyWo4ZVChKfX2IkkDYY6CGmTiPG3gLXvwgO3vm74GkrW249cUVnA1U3pJ
WvImqxljCtsNV28CZkiRAywBxEZQ7+deebECaKiNcRveS8sIOIZw5EjQlwokjjYp6Dz5yl1cvIlC
chH7bKW0/AuzEzEN+u/UyK978beTSXvnhTnSEQ1wVR3CCzIctLKX9VniLH7hkjupoDr9dRWWmesF
sopS73ekDvqeRwap+kQKWYZezJypXFKoMWQMFJ00y78BrxpjLoltTsnTXQc/4ac6ha0weM4AEuuB
aXNZA1Y202nN3v1rU1U6A1KXM1jA7RWaeB0UoKgBmUGVhVEp1s7RkG5jBaCAJKvlErtYV+4Hiobz
LlFFepxxuwuM5Uz7W4ZgO5hP5Dv33MO9FMLFlvkA2F3Evsmly1QPfgpd7fUEFAlHdgPRumHEALsO
yV9//L3UMrpOtZg8XhZEP/0Q0Jh6WJm3BpKNkN5inbImHbzSampV3xUJWa1Kwko0mrviDmz6GQac
/IO5v3wZLfF807ZMUwX5SMQU6cEe66vDBxcuEVwPmWFFJb4ecqOGPYh+P2GUR4nFELjRp+lAMwi3
P7WMSRotQC1Txj+1GFkYdlSfgpwoKrMye/ZM8p+jczDsPF1cezkkwhMfQZk1fa0PziV8SyV/7FJR
3dZnenSvZjhxfKapFNBAn7ZuaM4n9SmFNjpRgmeG+oTJjyp6VfFQCgexXpLl3mX30+aMHpc9cEzx
Ip+6M0X3T1BqT6f+EKaMsEKws/zv0tLWpS+tGl3sU/pJSSaC866TBitxr2pwvazL5BiikYjgjGNq
vFmXZaZW+7kuYs75FDNC5cT/GTPeXdxnM/J7y1PDhhRpBR4HZiZRr9PU5jR8pHivn1neMPFOLLFT
7PBzIMRhZIJqRBm+kErl5LE1RHIkNsqUrcrLMOwSt6TaGUQVh9nwco5WbKPSsfIVnSBVH/OHeJYY
1VdBhHWPwqT4LAjVCScBzRfKtesrZR3kTtEl4NaBBXQVZA0uZwpqrhkw+dnXtMh4kYLRSHI4mS96
XNr7ZtaRZZGDysLrMjP3QzZzpaqW95Vvdue2HVaPYR6ViEma9ar9lrG8qsqPbpmduBwzEy2W9FUd
AIVAGTOTM+BwDdcqSjeOzFOVTlPz/WvIDY+ICIJe24A+l9yXRFhqtJurX0lsBVcW2ia2shyHzHO6
Hxk94wz2EV9rfUtbZuXJucfmQU0ICYBZNpSgbRUFRZJ118UpbbUrKYhPZFnu4bUx7kKNPIXepIEN
iirkDpz/dWr262NbLWu9fRiHvYPpkR4jEn7Sn2fKyNcPuw3Z1gXO01V00ulka0I4Z4AYjyr0klZG
JEvaQLKQ/9zY59NZ+dCOB0lllVVgSBQqqVpmSBoIUc2+/ZuwbfIkWuUGzQDErWvcPMdOISe7HWbr
vxdOSIV7HflLKAZ0BUtaYF8ylfRb+UUg8Chwje9QxkwY+C0hVOjk2h5r1EpAq1tVO1hHycmedUV1
ph9QZs/5CpFrxsdG+F7h3CydbPcsTCbp6aF84giM1G95fZ0PWGo0FYaZ1UrD3o41krAfSztYdtwF
PCAEYZe7zPSlsGILxL3qfApk1nXBM5GEC6yiF/UFk9nRPswvutSQlXg7CpIT4f6A3vZqc2n1J3VP
HnHsGrrN9UBbr85YF0r8VI4VowVJzp0VGRnO+W6zEDmjMIS3gukhds8gMQXKvBELtUXQA4mVOXnB
BmV/G5gvDjKyBip2NdBZb+iz6sUeLu98i7FKO7zHBpubxoye4gNc9Rg4mYpQDFzpW6ARUUzWI0/w
Nxv+a6KIZb7b5IMYGt9pZkfRJU4WgceFIPx4z0UJvl8pwelY+zklsUgj9mhAnp1RsDkftGFsUs+k
owlBo01iq0HS/aT2VfgilU+VFla8rRGQrq/ukAWjIXi7XqOiO6rREMwyCpIn9qgZywlS6wQGjk0z
rhMfbzsKn4EiFbjroSmSKeE2w03l2WKjkHWMTTl8uDaj/q7O3sdiaUTiHXOtG2lzAC7herSJyoMk
aeXlujvE54x+WJZdf0Vt7NB/9nljQOe6HsxL5dwgtO+uS8gTfK7OD6Fw/ABNgHJahYok7x3avbFv
HcBKtrnF6arIry/a9WZA7rfnU8sSbQHRn5VPksk0svSCgbBnpf3sZENhWllXQ3nXmV1S6s0Mr0Qc
7ZxV7voH6QnGZXeZlqrLyCJGLQzHJMa9dJnYTzlh/OteFSa/7GjFh31GuxilJakGHkw1duWMQTgw
/F3AzEkSz+2n52prVqcLzIH2U3q9ug5nWeL0szfI6jAvGezHzySIiIgqsHLOOP+ile2zrzoFkjW8
vxqJRm1Geod0W1dD4umcaWHOiqblmnf6PXOlpBOpwInHFAg3rp6IvBWDpDd/icZacD+LefVq4RSd
nLpzf36/C6Z8oRebC76IuUFB5ms0lgU3pTkHp/54RBWPZ60J3UrJsqw+iw6tmN76+YARF4gARlmI
bk0XeyqeUxGG1j6kkWJRYkRHCGB9fxhRfE2fkYACIiSKbMbUJabX8EkO8J+gILhDc+d+I2wG1E7a
do4pxKXTR3lxlKQK7ZTrgGpmgaGlR52W5IoobNrLJjpzefnNxP5Wj2nAl8yE5ix1zSWUCy8MyVva
Zx5vPwk6ITL0YjuHQ61br0TbMCSMTCBL0qW7CZaqtjRpnMbtITrryYPynL5G8+K2ZJi4vNJOJ0m5
eaYUuJtskrcSj2wKoXPeGIgeg59/vyr7jzIqJcXowY/N+IsDXR+BtZRdvBSZ57QuMo7SO7IsVyj0
cDqRi9egPRYgtIGqMNeFw5cftlMtI/5GFEl2jQKOdIt06GnOsDHIJM/r/pnB1MU92Y1M5Z5Tk9He
GniprSSc7zdhH6pOsbigGirow6oUSkchGFG8SaMUgQnIF480FQ0xF0XbNgkn85gV+0cackWXpgi9
EQxYdrIiE/x+tvc4pWeiKjUEFapAhGM7t0WS/VRJOj06brjNalTtOgkB71cnpuMCZgqiF1sWHyTH
kVrJa/WqLvEmqenmZgL1ducJqK80MG7lWsfXB0W6vqBzpWPJ3mYeu/+xFbXDsPjGTlB3CPNe2fLw
E9mprkryjMHyDp7Xx6FmuMva/BSN3S39AYdX+1TnXgi0hSHtDT8apG/Nyu/GuaQylFxjrFpwtdpQ
fwawzI0wMWDzIA9qYHDAi9BwEKYkmm8zpenrqeuNKpdXxQXVuzdAa6wg3zESqyhNQDKui/koEot2
6KCoLMpO1rMitVk3OFay9Bk1aKnKuYNurZYYQHLnpDbED4B0ivHASGYG2wX0R+QcCbxgv6Dzl5Ju
TYVTeC5ay3avAB4+b94Bd75LaJR+V3KN4broiBJDLWgkz2E8UcTF38RHHIW/2fjrC3CopiKzf8wD
hFpFQugdK5yVuwoVau0eCduzTYwja+I4yHSe1D9jyCgwBUCvTtT2FREkKcvHLIGjcWWI2R/FxJWl
n4I77UMIJndDvnYKCw+s15e1CvL8+x/xmRBUAw2e9JVKbhSGTri3f2l6aGmLE7+LT7QzMG3yN99o
XQpOLdZFwrNrzX2XHuquQPxVbU0Rn2/eutDI3bWQJBlwAqSs0/luTg6X19DRuCrgZqJihbWarxfk
BfSIn00WOgJt4M6/Z91jxvk/LD3acdMNcfypUexMGNz/SECsk3+SvqZBfqtMrw3v2ZaE+s3Sd8bb
obsgT52vEMlhtAY0verg6ok7LniPnG3Nnp1zt1Eh0/hnBBaENJgmiPpadtC6/+MhfCX1etlieoC2
+cdjFMYtw8za/PuRxVIcX/OM+wEgoQ29ysPwZaYPCxcNvbdjfBLjfWWyKQvqo1VXmX6rv5uOlOQD
SroS0rHR/etQeqPtG/B8qvADt89BsxahEk8/HMKhTohsSMcizqQwB49uLp5FixhXe85/HI6n9Ah4
vO5BATyxC70fS0GJ/yDDpSNCQ3zc75dTNtdoLly+DgfSGyhLEQOrZCPKGVeInDE3HcgmGRVeO//0
FD9YzLCVOBZc9uiYF5mrip1PGI5yY3pgBxq7B/iSXbt1kuoP43h1vK4f5lktSpNMkIiXa/Si1HXP
3bc8uMxwtWYaZhxkkld3wbMgBaNOQYVJdkJqDvqVtLInq4HtMHkVBoGVcCx1oCxAMnr0IwavqNHG
pn2I9bc489CeEPQGOVXL9t0SjfhY+8vuOhxo4/hJu+vdMLQG6s3bnZaa/AfS4OY0sMMhx6n6K23e
ecPfj4yM7ZAH9qILRKDOLQDpZ6q0wT2lnsLIrkie0+CrKa5au0D091/5ujqIooW1HOtwKjJEkhMv
sABhjJosS5xVVf9krv2XKWDFICV7shhzC+RnuXQHhKRYLolyO7cuXnIU+nSJCwQq8lEK1dSz3v+T
rY9Qmg2osxT9WL3Hoj8sKIEjX0GTgOqQLh/zsVXCl5fp1s3nRt5+BHSCqB2cCVH1s6i1L8gC29tr
gzHTyWVDiPj3vcPqxyI0brFJfBQmHgXVrzRaqghG+KfqntEmg7eszTP6FtV41iATgF5Ee1sgOmRV
bTLyNMnVbceak/kKWvU6wDLDKDMnzAQ405BZdPvfiGOesHgs95K7dzzb7s/5csbDxyzFMZZxdjxC
lve1DDksvwUMNUuXVEj+GyylhAWc8Oe1oW2baklbifPgD8GsPqLg0azHQ/dsdoDljC7ojTGs5AKl
3xgaU9NTTrBwTMeEJGb+cFrSjztX7903hWKYFwC2q2Piqa540tLGSNiKZFdJIeJg/+qRGrUnblfO
yG6wzVyGnvSP4VnqIHD3km0KxTmWwvSyZMjbiK14s7c68jdZ+yig2SUNi3p02DQGJll9OOWTOuRo
RWYoIC1t4o7Sm0sAa/PfnnnaJHQ2RmfUPaIxtwXPcA8Ki+JfHEtEOPaYNNIXS4dY2N/dyYQJaFps
mJvv7PY9fLAEow6VbWwDNM7PuXuAnd5RkSVMs2uWrodQf5deV/PIT8phnYgvw+JDYAujgEnw5Hra
8yRPbkurxtRIDS739SKsrjpv/4AiG31xSP6AvnncOHECZ4TZWkp6WrHK2f9/bN0e5fKV0UI+w1jR
8RGTSL+lo4revJ1rWjJTxVPjEyQe8xuczxzUZw7eqPx/4wjHUhTn5HotNT2zfT7dw07sPUQvNSFB
/1l6xKzOUXfymp6huGJkRycS2qDhH3ms+1YIS8ud82tkeZuAR105G3QIhySaSTkOmSCxcYaUGLcx
NIjli/8ikHdDwJLNVaBEIf+Cm7NSpiOBLCCS7MHBXtR3zpnPIVJY/R15P9gVcEUHgdSXyDQiJROO
9oeWBzy102jNflvTQMBCTT8kw0Wk1DkzkkhmmPxXSo7VxBLswD5KMew06Hqu0+aUWd4S7K6UW98U
U0ZZ/JRVIc9Am8CBKCPHJxeIEescjz2jBMqDQri1f/daNB2/iXO3YLB+46UZug4nSVXjjejJgYcx
HiRJoRomwswapgE/lIQR5I7xBi+JkcTLuhGCoU/rR9aiYcod5Sn3sSxsKKkPiYeYSKm2b2lnBgRW
a+mVO42pu1NoL2oM0VoJDpAYIIwYhiP+/++FOSPARWiQIQjJv6pITV2/+9xyjha+HjBKhKlloPKX
Ae8NsLJ1IqmYMgv+20SW+wvvJF/DkGlHXi91M/h6wmwDPgD5h/PWD043rvjj5VceZy8IUBC2Figs
yrrLrMH7o3mrNczQfDCtbFjfrhYBd/TliPlAOJZ8GuPd7zUFQAQ4Yme4fZkGs/72Vd+OqnXC+2yC
JszH4UW+vHX8hHPwdOqyff7IaXBGIDAmnXXKmWYPNJ9ECD3lkvbhQrr7JNl7wJ4SyQn+bogHOt1L
pdhbPJBATlrFZB/9w8Qlhe7WuWS09VWddsqhzXwACNbRI155GdMOr1LMWl23o5pJuyrhJAvP4QsD
JobpcSpsgpfeR667sJXhqIJpX9OBzOfs7F406LUeednhIW5SBb6FHn+Abv0pA2MFOgEfinV51LSk
3z8f6aemQIeHmlytQ4SWfx380PWqoqX3fpELBy1aZ3o3vuezvJSRCY1CZrkzkQy/vJrKX51g/aqN
YDYnhPnAXWUekOyJiV0nTyjtDilPJgs69XKaHgI6/iqDvxbMiQigz8HCcWBZdJ4YfmYgxHkWQM/Q
gevPZ9esbkfs+fEvum9cF3NyTsfVjjOdgu2NUeIdmWsn45VRYNprZT7e/UWWZKv/yNC23EmsOMoX
zGdliZSkOMbqrgAR1zvja0CjTpMKPmLvR5ZPPRmpMnLCot0MyaJYJ30PEUT7xyysqTiKXGDYLiIV
hHBNosSg78yVoLickmgZyEU2rcg7/V/GasIsPZg4/zGXBTDBecYLVmLAjeQPrCZ+Eezt4m27+IP4
gPFBBVigUHo/WJqLv06DKNmW915TE+jjTSiEX1gO2e70zKlmqG6mmARAeJvctV2TbL6kEpLQ5WFZ
nD+0oCvWhzgEKzktWjzLPSC77c/QQsTwjU1VgT0+oD3ysgTqpGHcfWtaXI8Ja0b0TE4dc8sgirta
X1hwKvdPjtsUsImNKTVh0GmtLa7uGxO8mWe89Nzvnx99Ks6LDLokBDttVNNoORaT31oG/W35B7YI
kyHSNTKAq2sKUg1XkKDwR/BqOhVzwmYKwO1Zg5XPN6qJzux4R8b6WDkZhwxTqfYo3WuLstmXi+OY
7f09ZwZnCVooBHTbiH91fn9DlX5yGfTb7LOef6XcDXhfE1MrNBGXET/kG29G7HVoSZvpIQAs5m6p
A8wkMRb/9+Q8P19B7xyOtGd/bAuv/ENyGkBV1qE++U13ebU/1o8vwxR4yMRN0FTexqdjyfPC38M+
2ObTOB5RhylV7pUZlV7vFrVZvpdCRVrm3u3Dk3EX2Tq6XCIM11jI9uUsWT1RxFJQjCJk5gcTKv9O
0aMcDy/6Ei7q5W7AxLYad4gn6sZHXQ5w5dhYmZW52OmLCrRIG1J14tGH5eQfCFWsJtbNFwvHnLGJ
P1y/OvvLl5/4bmob1TvWdqD0NqddwxRq/5sYjgyK8MjiFWb2ZSxHWNnkJG5LQ3DnXkyKrXj1fSL4
8OBr6WwBDAKsaiQGUFBLA00qENr9QLxfGjfLXlsZfSle5EYSThQpuoMAX8nS6e9yPWpfQSA4ijd9
S7MNiY2CjRU9i+D9a4R/BKPiK65ZR4Uk2h9Rgo+xJ5ZjDm1LVyWFlO4odFByZzfAGk+t1hFSriDQ
aVM2dwvnnpFBu3NDvyO/Xo0EPHFPi2HSuqJfSqxdjOzQtcYamMMwb5DDtgoGdWIsm/ROZ2ocARO2
i5chsA2oEDLdrmc7UhPNr+u/SrgwjziGJ0UD+WINo0zqwQ/zTgGurrtvpa40y4uFSrPh2njtSaOL
YS+6q/tYDbEqcMEGjcCrQzmNjPyzY92t6DDcpX0J7EWFJSeCUtWbic7iO1ySue4cC0f/SqqwQDoX
hbi1EO9uuvE1DfP1A02iyQG1vlK3VRHSDLlz0jRsTw3eVTSLHGEGX8TqrwsPKnSAvumHUzXTuNo+
hM4EPwHhI36cYWYQDW015OeiLUlJqNtRNMNcUKvmQap3PcjXLsdpZCYWOJewlO6oTjrX4kYhP48U
dUdF4DGMCedMiZWETJuXQhA0spAXahZAXjapdwaMrKQgiJD5DNLkAqy3QGOG1oZ215rkH1kZpFq4
oTaE2QRY/LJFHiYTX0cZ+hv9hpY7ZK130RbhWuAzlZ8imjXw7nFhEfwRsbJTT/2VRenvf7sYaFrU
kDpru5XHOZGIPSMQMM0Yf4HK/ecpNkcaNZ7owXYEJ6zI0Dg2hTCVZBkw7sjcwhH7X/Knmfu5pVCX
J0QwrLMqSxasL7pjRGHkT/UxEFklXOI6eiX/pjBKxuR+g9AT8KWkW6hZV90wJERZydaY5Td7cJHX
55TB2Q7xarm2tt1RKHzMi4EJiIdwSUtKjUDXdDvchlJ72zqv2NfQL5VqXOY0YAXtnOsQWG0mGpEf
Aqu/yq1u3wcuzkyiRfQ+EStS789fU3ZOgAVpixJFH4jTs3g2VzSVUO1fcfOHffG6yF5ui8f2n+JV
nqoTi6oa9r79Q4spNJznWo4UvNsKxx/M0Yw91npia6tfZeDuM6kl2GVya0pj/f2HUcD/1FD/PY83
KhOPqM3MrA7qHcaYHaCRXTdAuZC9zzEFcuyH6eekV41/WRUFN/NAfmKiEuV0xHBx1bbbIsizL0pd
Y5nJtQlhpUeyuwkYaKh+Ph1579swyaBA+EB33Chdq4JhGsv8NKoo/8O2rRSIjXCUBsR6BaRafvQM
6qwlUjj3oCn2ESieT5gOUiCJ4yclnzHduhQdDFeYPvW+WdJoPVBdVWbXISrjfYTn4MXHrYhQnukG
pVXv+sdanyeeYKBqsugacn672c7Py8E4zrKKPlU5Qznb1G/9CVq1RIY1F1QUa7HgU4xqWdo6icla
2KLgTkCIM+4hrsNAA1DpaCrvGUV0c91Z6CUVMzCJg1pKVJbdPuZqIEG5/7QeGtQCpZeJcY+V4CJf
8eJdiqwjWMwihpQ87JpW2vEyztjhVCYokF4TlFLju31akiQZ6oTjrZCSD+JXThSgbg3JqFFHIfyx
lVuKzXDpx/tJJzUGHQhe3uSCaedXeKGpWtKSKeI0omUWikb8QUFbtNgs17tyY2rnE4ZcfeN3pb7Z
xKn3Ujh7o5v5DA0NauBPKH4sUwf+9zVoNhTp4BYTS3aciNkEi8mnI1HVcFz6ryEo+AQmzQJR2iWj
hv1yXq5qHFgYORaw+BeUMjPbLUnVquiuOOaVE6I9igy/HkpjYrQI4Y86oYEU9zzwLdHibe9yZ4Jf
auquCqt7gb5nHD2CCLOT54Qh5E6MeWyxFsKgBE1deya9Pc5pV1q6r1WR4KTvvWywTIbHzXUmHJ6d
2QlxiKPIGygtWWFVSQbS4nGG5ZsvB8N1VILJnfpG2NWjJdllSuwq7sEv5y4VUL0d/x2C1yXy2ckL
ezG4jix5Pmt2rVtNsQvliLTUr4QbiO90pM2nxMNUUAEwHmpF0JO6Q+pqMU02aQlxgXJbJ/+5aABj
/qI4K6DINdn0EadPxheARSxYLbTbojrbiuKE2u911xGnoEzd9sle4sqaCtJQBDHltYKOCudSgsXC
o/Mpik8VMg3ctvVv8xYB1OwqWcrTgFoCCXrrJ2kpGFBsUjrAT3uylr7pzQ45OH3VSN0kTCCGsIfs
2lWwRL3wkrsi1k9GXcgYVfsK7tUoQLc9zNJKT1vQkKmiqzLrNatvnoCSlEzORpC9SXgo1ekE4I2h
1A+4dXuMJNzknbjDrV8PuR7qRi0JBnKuLKUvaVeqYHoZCSq1qfwJAV7H/seEzxnpX91XrGY0TzrY
lDcWC+1RTHHS4Wv1UaIcxHQWm9G4biSYmLyAW+PP7c1457wAbGr4eZnGoKYBOHag6z88uk1EDdQT
kSdI2EM26EzSodEyb/AfjlWykCPYyUOFUllRYttg8oja0vfwfiANz1901Q9Xlm5tmUcg7XOXLgKQ
1PL55dZlb50y1kgMRGFR7590dGzIOh9w4Sgdq9JHOnq9DRc6rMxIfZD8M9QGjTbioNtGLXeV0iYx
gjz0qMP1ZyrDI3nMUmS/Fjpqc4XvwKpQMOXfg7WRFrc3Ib58Y88bO0f6op+mpwHOqetJDer6wgX5
Z/X2Z1bdBgD4uQeud5mEi1y2lh4YJpa759R3AJsbCI0WTdlLN34EjXvYk+bYjLH6XV8lVRlqHIJf
6zU60grqr1FJ+27YgpRPaC68ugqmW1ElRM1n17/gKhIVk1tY/kjOucBh0ejQ95ybKo5M26dD26gh
nX1mAHLVvHFCD1IRE6c64GbEywS7sK6N4CVdHR0tZnCaCyBQqK3Oh+R39PGu6ZHwGS+7Fokdb5e8
32b7OXV0QSS5oe2foah7mhbHg42fXsU/a7iaIzYSmeXf0Uj/kKMPOlNKNGLtfd8qLZNiCcw4BRd7
19shGPO7padSBSeqVTYB+keDhN9ZWTMlWUk1G0dJFliKF+HB9cewm9Y2ezme1VMwx6rLY5OJKfrv
VMAbnNYQai3xrGNXx3aTINqZpFFSLfl4DdWgYzJzzVMzfsbRf484BkgP6F91FIScGF4LGb8njm5s
5g+gSFVP3UKnd2xCrEhMeiWwMPS6pfk2FxcAwApgR8DjgRa2enXM4kLmcqoKbm/DjCLZyO3VUway
YnFAP8qlZnLFIausubQJZw8CsQIY/2B0/Fk0tD0tt6X5sT25mxauFSwvGd11DAdL4quwTLMj850H
UxGsl7UtC9lLAg17SGN2peRYLSc/LAAEFwE76zBY0dNMPfAncjgchnxTZBb2OLno7C0f+Q/u0tJv
2tGbgrtB/QYkxLdPLB+ycraTmDDjZRkeRL9T1T3yTQ5SqOecpnaHVPUxEa1X4iD+3mZPr2czG1d1
awahus1o7XPAni/KSmNtK/TooHfuHVulwYxaYqEwAPiwhM5i7RSRzYEpsvd3CF0QIfukhnZHwJnX
4GSnvjs+lCjjnXtrBN+W4b7TnwNAYSxhEkC4lJ9nQtMfjccOiF+7MHckaHCPDlK+g/hN6uvAFsS0
qP0DeTPM6DVJlr2kW+luKCdSZku0tB37bM0UHBMHz3/SqRY2tgGResJpjLKZyICQMjWYxMFZpRYV
fRb+Ich2iMa85yRi6RwAbZ7bJ97xcRjH039M5UtZt45F4qfERrYt90ahZMBDXI891wAlrFFKHlv0
AGt4eUx6sjF0RbLx9M78U18Z8I2SkE1XyFM32mf2/SEwa6cXwZCtmfvzhz4bUTDQumh9mHnwmYSI
1JnPSs2n7eNIZ6p/ez+tlyXWX2wLM7JAxKQ2bEXEffHSvrJbPT5opU6/HqDDfewVyIZyKF6TnetE
Q1CtxVEGCvz97rpoIawrflju6tsYvevONZYNakkQxbZ6CXGCrxpIRMljqwcVZ3LgVkz3xp+b+DZx
lVYwggqJxIEHEUxq+swwX75cuyRa57b0e/SC8v8qL/LHSKryQd6ciImfBcacVFO0L/4KHokCyyz/
j5X9UfM+HoZQmGIF30Z1Fmb5RwtHPlUPAZSAOMAze+3kwQXQKldZ1LzTSbyFsX8dCfb10IuaVjKm
jGg2cR+pHUI9+cTR4vDLo7rnHv27xO+JdCNwtVu8PSRhFYfnamPUasqU+nbAgOU9XRhSRp6LPRIk
2XGCRrBup7weOxx4TM7h+be8x2DPCe3emiJDK9dzPRUxW+q58O6NtsK1XvJxjw9hGwYi1afu1bD4
jiBF/GwMuZnzhj+SGJ/eiC8sDb+Rud6HgvYcA25UnZ+fZtE/GMSjQEpQVMzTtqnHRJlReOVLGZ4n
lof6aoIfnGTotVJtIwwMImQLAWB+TEc9CoilI9BGF4b0D7oDCWEVGPgGqmzR1tomXFYMAlY6IPtr
rTruYseysoE7GfARAHzusqneuDe+FuuEsmtoL5T36bgx3rhoMMsy7+pC7PvcwohMH5tOQTVQFTBm
N0TwOJwpZexNnmdfTRzSUAOjBpTlGwOopYm2FMW3yAc1zPRhGdEJ1O41wE6B5H8QtqG15EFFkbgq
HLc0Wc8YG8qb6wfawOm9b4z3VdiqLp+LVfcKz31grnOZo3KQ5yEJh0f1XLbQM6FZa8qYFs08HziF
oaK1jLZg2e2SZt09OvjNKGRYdR8BcDOWoHt0vlX6WJJQ2dFGiXYn9UjrsNNoI6xxPtDj183bU3pP
xmgJXH28FP3Ptu+nyaanaUsr2LgKpVnaH6AJsiFMC6pPvVxHG284nQIj/aY/0bMmmyb71VikPIee
hrJtCc1YoFpCp1p5ISYa8pUUHHrLkl7w9+aA0c2IOamGhqjoe5wZTAuz2Ki/vCFpvetZ2n1GaOjv
F1n3bTDsbxpH2p/af6/co3vbEnBPFAN4yRlFJoQKHhL51VcgVgCky5VXfngtgzv3A04wVx54X1El
WeaSI6/bC1Xkcw7J+9FB6g3AVvV41i/6cJB9m5Xyqw2495p38GNcjvCEEsSfSABuA5wFvzFOMWuC
lOW4pFPHbgpObiY3Y/ar3kSL+bgH2p5vAxJ8PdI7ptHLZpJZmlXnhYO8oiWNmNmnAvpsm1Wjl6Py
VZCjs77E/7NiCgE9PfqeViHPjKcc/UprHQTQTxIr0yWY9RvkdSS6FN59SO5E2KpS68evUQS0mdfc
V+kT28y7fPLy/IzhXjKR/yj1Rg9t/qpfxeku+12ZQHkIAAsmzwcUWyRQwkUxzy+1xoMSe6Z62GDR
p3pa2bm8H2uqIcjYYbBxbGPxNoJvr/q8M3NnpgJy0PlP5DVKjCN/jQWIOtXbsUvkR4Pru2rorgA6
EqRiteMwAS2xHYolVNsCYuSjmBgSKSo6Ms1va+DXNGnrdnpw/b/lLaNiBoy+rECGXZf3SpzOeAuy
fszacA8jsZtMsyELPtfJi9upv8pxPhjiHB7IwzXZuVVEQGZxmSFFrdSyKPnxnakTMhwhnu2U6+SX
3E0aXwylIiwSZg5OmBQLKxCokgWgttqMnvrVV2X2gCPzqh5ufxJ7O5ruLgeLAnJOXyLAS+j2Nj8h
KKqq7y9VDAozIRf6ns7q2KHptMPTFJLvOop8UgwbM9U+KtQRv+C88xXQY0odjxE8lfi4G41pq5Hg
5j4TkpWY0SODWweUz2frZZEdqucipyNdPYC8dTJAvZFJE+nPhbwCuIHhq5wXezvTDrjgQQnQg4zV
ufc1idNiLOIhsmFhFAWU+na+W78m0XSJBHspJcnsd8Q/o/x9e/sxR98rQjuErYCyL4mDUrNS4aVF
ginbaxaJpnK9RBKup5B/44H3lJJdPYlyeGkcSL/B2Ee7cGkdiH4/PHsfg9MoOQdHGjvuf+Q+GxJf
TgkUlnDYxoot6e8XJBYiEXtjYg8YBHO9MbOxRdEAIaTWrf0RYTMn8Jw8lzUFNZPh3+ZTw7J/BcgR
2acnSyn8M0/LQZmFo/OLLdITK2PtCRUhBLNjsRkGd2JWtAGN4F/O+2lxJ/aupFec8zF7CBu2R2sM
YaRDuPc8r2P/3OKyoIvIulEPbRrEw2zUXwqMPrr4ROHnFYEmc/QVh0h18pKsO9Ffwd8TI8bRNUGZ
GbWWXhcwIpmXiHr/pSgA4IDMefJjvFJegDo31j/lA712/YGZ1C1/FukOka+b6CpKeQzO1V829C8B
RgWrSup1TYxkNvVnAqI3JQIDH7TVjRdTlzcj0uI4DZPnfw1TfwcozJnFkBq0wryn+qhuug3G2le1
7MyP+aGPIdLsI87NmyLoB9LA7sEzaCX3i11OxFBAC0jzEYXnUt7BPuADFzgeb0bV9WpLDZs+WPy2
bu6RXkEmnVjl5QXqTWzhPVNJ60dVCVXBFIXTIARV+DQySMR4FB+XvhrYa51dWTqoSKS+g6EiM4Gi
mjDhiLPO4Xn70zxdbqJP7rathiAqmwMmQBC0JVV/UAnRJ59zAwxPaZ4GnijWGoUTo2p0SEImxh51
GhFhkUX8ILaFwqUxtDHmqXXnnn55FRXNXJGxjkbOXSd/fb4efvuvWLxCN2DcJKOz+doxNxHN+Q/G
pwM+JFtw/MLvYinu6GSqgukm8RyrU1/IjhFLScV0X4YsYvDq4JOqo/dyTCs8+Hup8mcj4idrUE4e
QyouAu063nN8EiJ70TLwrb8S57C5nbqZgfWUOdIsqzF2MigczAWhX9kuGadLUKD0075oHk3z2937
6XASeOGsDQAarrMjId0VIGcUjwBNoaiOFrO4CPeVS7UzWqlibNy/xBwtGJoYzBJeJAjo+UAtWMGJ
UpgLPbbi9QnGYtG+U/63+gRQV40qqaH4/Z1Te6wNhPzZTu8FMfP9mHIj63iGXBtMZ2mpH/N+jYG4
vbaUhFyEz1whXVXgPyGViRYhD4iplpFNmOMYcE6y0cLRKAoMclMwDjQbJnt4YxKe+53pZ0FJVGw+
TuDVe4iE80cfI0eSyCTnfhTzQjtxNQcu0TPRh7xb3umrU7XpyykMTunvfbs6JFbv2ADLNyRAgdIr
QGXKWk78jsTOX6WXp9QcYyxuDdwYaQY7EA3YIQHJUVJaRL6UNxv49YY7FsgPz9wCekUpnBqPnc6g
v4S7a0LxTNzJvn63ady/tXsk9hM+2cwTI32hZqfLBlwZdVsCVF2g9vLM1c7NKtRBS6slARgjI6L0
O3D0+i1G3Gj/BMBzWoTkwy9wqzBI3pHcZ23ODqphVHVrWo9QqPqlMmvLHofy1/8sW7a65rbGZ0gz
CpPCjyU+gYNx8DrQzKCTR972gLrn/X3OhL9oFz+6wlDuv9twR71Ns27+iX7461a0RkYERbhkPuwy
K6U7/EGR76gKH64Ii9ld6JyBDE7m9CNGJiq0rA0t7XUSkPJmChp4uAZn8XbcXXtud7lNVYkF64K0
RlKuG5S1ixM5jTewQE+tsHAGYeia3JHT4+rx5YuR8zDXDqZjqnkgXp/h9GvFbv49g7qV0Aw9EuKG
/IbuQPPtuC61ez5WP6ORSJPt6KXZ4H8Dr6yBQ6RKSBX+fGQmUa85bLBrVve803UXEYy929szFxhR
U54p4FPHMvgbBb3b6n/86W7k1H9LEDc7Dt6+UoQl2OAC3wMT+jYYP+FcVyrKvqFVMi0xzyC5VC3O
uZFIFGDlyaCBqPagGfksl5cFAYsuNvpK29IOiY9WRvnwI4xRa4jHrokPyvuvcERie7XDgtai5kXt
ZBJbhapLkYejFg5nu03MbAhev7LqmAHj9AbrX401u1m7v9Yke7PNgl+bm4zpcjnfTSWj8DtY+Azn
aNEdMZLxE20XZE5htv4Y7mHJCNq4AYjujUguCL4oWFO+WaqurvkGP0ghCt+ehx6TJoF7z24nPPVN
aw73gFVgSKFA922l/zyP4/XxMvhUfdOkM8LB8G4YHC6jku+LTo5ljLfWst/VruMNnJZ1TFlbXBpJ
4ReljUk+UAgHEeRXZHErVvPLB1DOjK/Lykjf5nehwXXDn16n0Yt1iSMPhimOyJcxP+OV9Kd+HxvZ
T6N2HIjfqDvNUiQyURMMlbnqXbkFhpdG3HMJ1dNbL/Ua0SGYPzCNOwkWV/ww3yooz9CFOke2ayae
W1DJhFzOA/LpENKy/YU4my9i4ezKQa0rRi8y8/sAVMJU/7+ti5MfhB17KSQXDQwYIUDEeqIhmCeP
SOxIIJGMgyfX3Ptc7lv3eiYPgeCHXjmwoEVXl3vU3XR9bd+l7TE6HnV852zCAdl68g6nd8ppkfDw
u4hCPJ8tn/nOpV9zPHLO7XU+gJdOY12PdReMpzjMSfRTtxLvWRtPdOoVQOTf5/f9Bh29WjC7iLt0
HJY8mmWyl2KZuFKtKmjjoEEnBBqoni3QSF5+eMgCt4dAT+3eZw7sHeFU8vOFEYphM4Y5qJlBKZBG
eb5TRuBHnG5VUaLsiNc7TmaHUrqIUUoZzRwLUOIVVopxrfZsbZyu5u1gLekasy9jX9Lpe0d6VkEk
zhciMKLzroMdEDeswz4r9uQnvCY7JPxMqnpE2jzwZ+w8oX89UqwTpHuEHdCWnFphnN8K6qoCYYRr
817x4PkMGFzfpZ2E9k/jfuleAgIRqE5uNlEq3+3Cdpl4tOizdsLlngeADNQpykfv4QmxCKiKSVe5
CdIeihADXNbOrSLAptbXz0ge5SdiYrJ3goHZJVaLCCbV8gp2AhB3WMDqpGcjXaVmjGGBgm3QPrYe
8R/HEb4o3ZTzxO0Aj/qQ8grImy3ONSpJ8tGeHzpWhchv0xitNwG9u3PHLaxBAqNrZUaWJFtyAn4D
E9KypTfCUpndF2JlMKvwyOc7x2TjY1vvDFYxPyMm8c7+s8rgPXHd7U5Z+l4xu3JzwoURhX8J08gU
T7Rx2DhoIxIuoGjvHQssivcmooCqUej9geVxQ1E2fXYCqoyZBDcAHqhMPLMxSctHeFPrw28wFpXj
/0qhdgD19i8qvy4hVD+BEHSvaKcF3hKCpNnn2djSmY1C79hNz9P8QhBIeVPYuBsq+CuZ1X9EF4lv
NgSuXFvpG7x8GVoCXz0Rqpqpb5liL0V3uTFyyvAV9ezVBODSQK6KYC07aH0vfOhBoTh/1Z8kHskP
QeN4Y2vCxPX5S14boLtT8HAyG6H6Uh71zqT2kIXClj26UvoWLRNimdLRT6sNzjpIOzSsHjVEWg7F
ktzxI9jweLomr3JxdDipoXPOz5RLFFBsU17yLbl0CvH+fTmkkiV+MfjG1vYphONjIpGRYsw6C+fP
eirdRiyg8/y3Li47s/6G4e9bnC1ndFtQp3FyDNiTtRMbmRw6Kl9Ur6SrDt74USa90GDOM9vbLRSA
yuHRGljxm133EHbQj5FBCRM31HmFIn4vJOI2V0dfj4XHLLo5VLyxLOtCfRBgZt3UOSp+wL+fh+k7
1RaCocQG1FGnkJ3P1pt2UevmnXhaP44QyFvbmHOITQmaihH76P2aJh09g1N3wzXIoL3/V0+hN5vk
XY0AT5dzbIyiYl3JBaqeql+DBXJ1+YSORAQbhWlMC9c+yjLivlAnCGS6es874H3NryjhAVkZDDbB
0cJyQ0WjQFbKYrja6+fn30WjBvMWebCGZHhBs0bx2TC6RegLoZgcHr/qY+2Rs4Ke3IWPOiVasaqr
0DkDgABG20ZgmERwA+mQ0UanL2oQK0L6hIqalQTgQZdgkFcp1B5A+xRxzsY+UGW2bQYzxD+XnWiN
MlvZNkOWAC6SEwvHEyU090o4//BxX/wIMmtbnv0Ec6LqhtfTWaPg7qp1mvz4jOsByoAYzp5+AevC
GoKN90KS6GWHsmbC7uMUVLFxYC5vJHLLxllER735LPO85EI5ahLXjK8/gdcglJtfPY3lklmmrcJY
ZKVJ9ZNxtQOwJlb2CeASJ+6VYp3mEKvmRTDdmUKkcS5YWV49nqb3CTcKHhMJVKeUW1ar0Boh2u57
Px9Tcp3+248KsgtK1+uiKUMF/fPrs0DTTuULdy4iDdFNi30vQXBj//t9fHgga0ZpDhuH88N1Sc4f
1j0xztE+GLd5C0weHnxnBg7q7UmQrE67mHvhxeM0xYsVYIwWzxq00moFZNGBi795HrgntW7h2ODC
QlcrGy9hPNOvT90nfTdXuDHbRkR0hO42X0hR4kq7ni2427kQJprUU9dmoka5AYhAPejpBMjUA6GI
Szsg+a1KA0h2wpVk17U3e1AFlJE6/tjLj1JrZRQR4uUWhYw6ypFXA/JitoTkX4DFxd3k/e3rTP7z
pEvdiV3cumG/CCHmQya0SWjhy6EAFA/R+grGOucI29NJAmEotQP4m9kMQCymP5Pyks1H0HEcjygw
1LIv5uBoMXpuIQWm4PKJ8V67mz7g5AFG3DidCkCVfRDtifIDngqZpmvVSja7+s4QhATM0aSNVi4Q
/EvTF0iMqn2MMrFvu1N2HbVe8Za3EUex3q5yezHYipn58kTQ5mEU9rgMTR6MdrJkD/tBgdAphoPU
i9d4M68coQ3XXzMgL257P73BK59BBDvF1EdQtJBI3c2naF4MtQStKdmAlckWe4v4Y9QKPbzvYQfi
YMYBFezZQkShATdTrJaJ4BPGYCkBkYZtLzhg17FwtttY+xWFJN7p4M/aE4fsDek8cTM6NF5FGJqc
Jq8tBqewo04EZLipE6JpOLwBoFn5RkeDPQtPn9b+vHtpkROw1UshBgUKE04zfA55mz2u1uZRvoLm
nSDyx+Nowvl9OUeu+hDGn0ZXGPYH4+1gDp2MQfMweVtd/5fkfzSJ4DStPt9ry5j1aj51Kx2e57aT
cW1F34zto9oh3LW/9rnveMxZKJ8bdxGW63CkhaRSZuqNb4mN11ia0aeRGQZckT99GSwZXrbhD0Am
bSy5b21vxpEMbwxTKTohHIkhjuMPU2BbRO27i5R3tv4IMyrGv1p/6DHlvzvMSr8EdF5FqbkafO05
uHjY7x5p0koHui+Z8Z/2Eyh7P6HmV5c/kxQ3GNTRWg5vuRdKZfeVXIicnIUlXUJ0vBrFHMP3PHuX
JwzckRkVWFyAmWgT3EiTJz9XkCE2rH+nrjgKXFWU0FAiM8nftXZOyZR+dN3yupDzxw6/18pD1MPt
qGgwiNQOMMH9V8jEtbt54ZBA5edn9kSyKSAN3zeQaBCNlWIZSh2CBU+cIuW2JjGxP9nXppK9f5XB
hZz2pShtlK36Kmg2vse3x7A/AFwHGEFfm6TaCpZbB89RU2Q5xMO4II0wqva0s5oZGcf2kqfviXAh
vbS4UlFIjaEOxAxaWp2rxZEe9aUrUDsWjAYQL1CVuxKKDqB/K3A8Lw8gIG6veC91IYX4ge0KfcaJ
DfxCd+5mMWi/Md+zLueO1ewnmB+NAUMdpUdLks78BMR/v3Z+zDUjvn66DMM0H5TpMCox0zvsJsnT
etfd15cmkhMHW0k8X3VlV1zvufrEvSSWK5ytCXokolFijbPGH3TcBSuTzXm6wGoq0xVJKWASrImv
tpcp4+IyLKUbHsr3N+ZUPtIQvCPzH91yItV13vqMzVZRbfmkOwbuahOTB7DGO3qQ/xjrYxW+2ywK
wbLu0oJawbN50IWQMU8R09JmmII+klS8X0sR1Z4Wm7zTvUO1kxo2NEk/PpYfx/13ZsktK4KfdS1C
l1F21muHmKPTdahqT2i1f/dSgv+0sgPjAUrKAAoMWqmaA406T4eaeyuMk3cGrnq2iicXHMfDCZqC
aZjSx4bml9Kw+DYQcO71YnPlxP/FKK8CEz4NQAoHkDybYz6+a6j/Z2YTlkYcBW/3s4L1j5nFE+Nr
ruCPAFP2v/4MY0DCqqitQjGAibEcYtICUbgp1ytzAw+2tyIR4irLu9y1Mz4SpGluBT4kdgqhm2VM
vUrtRlzyLgH/svBDRSa2l9TDI2SWW7dsPilEDw79T7mT74LtUVyAdp9BOnS4qAF3EQ5uilu+CoaG
z14flloqqmOHvAp/8a9ROQ1+9kuTxPL6shBEZDAKF6cOPPBecq/M5gnmsLAEfyEhCnKc0odVKbuL
JnQ0D5zmr0R8V1UtuZlOEhDf+IS74EPYrT3uHOpSKsttuDhMFtcfp8D4NtAeYLcmq/n4hwH8Fw6s
pDOWx9A1u9oQ4GH1DBYFzULz+xwQjnQfIYpK/JUzKLG//g3SVNQ5EbLxyTKktIxIcXY1P+VclK49
KH3JlioNzvc+IBB2J9UpxVeGOnCzuWYGUn8AfbCRPw04OjWDcqkQhWXT3OIVsjQi4TU/E/PgOSL8
NYRPGhR2vBxFVLU7gklWhW70RLRJSGkoMyEkTJ8SLI0k9HM4ImULertPodMGqpdOmrRQZIjf04EQ
rj6jd10nXGEl3ldM//GmqtJsJhSpdDM+c5f0PPXIPv07+BF+IK5gdk+j0uEYW2mFvUGesN48DreO
Z3GrhJnAHR27e9QGfmtOFTS3FN8ZrLCnznT8olGK7rqrWxo/dqvNNVw4BHBse6/yFcDrkyO5wEty
xa3QAIjvbr+8iYtqWZi84OWLVcL0QDnKa3NfeXnXwpGcEEhRrwZuNgR/DNBVWrrN8/E9Ts5yvqU3
6yEslmmZ1uoLSlxVJDAi2e9DSMyug3mj5liNaVA7AYua3yea+lijZ3FrCnE3d9hhY50qKCy7j4Hv
z9RdqnCI1SB5HRCCST3Asjf2+WC5TX08ZMcYjEG9Kmkz9O9TJjzOUc85vrWpBNKhhitAtjkCZMIp
+vLNh5tLV0FnkcLm7IaW9bKqy2DRixdc8fExFl0RwQ0sZ7IQGEqziXw4q6S6b2zBP15h7Cl8qE/v
UX+kfk6wsL3hxFl2lamvbeXKwv2c9udgvHeDc2YEud2yXOwoPNHgg7rVMW+LewW2+9BTIZd6bFyo
CeGFjIETJtE4nG12aDFpzfD6b+b6pJDBgZIbgF1Am/zsCE70JWCKlMCTlx3B67q9zN+1cTkhml2Z
umN2NoayQ2fw149JVoVCZYmgzJ3VMDBmnVwik4muguNi+sWmqMoKHDTwiWo+r7kPa/JEi28ZZoxQ
qL+EJ9v4IWFNfafdIDpoKeb8xzBQ9CNM3c0Dh2zq36k+ZZ+jrmPMoFcYLcyWre1UKFzY/Gfh+Nc9
hR3hDQ3BCi+LRWqUwW8HOvLl11baY0delXzlBGmr4C/Dtb9/aSZH0pCmUmOCfITEUsEMbFsmeYwm
YapXYbirpoWcP22TQdeidYU+XrlZ07q8FxR3NHrJPYG7XaLuxnEHLsXx4k1Hbeh9HB0theKYo4a+
OWgfxb397UtK95U9HANomQRH648QnviHg8fz5XgygyVQoIXRfu4lpnqkUvQ5+ldGWFcILNMQgbPx
nqX1Pcxy82/FcaEybfrZkZWD47ht1HByUa1F+LN/M1iYULnSHEqXfJv0voXXGa4+2G9da9Pdmgzn
vhYSh2QIw9xjF5hozGhc3Q6NGnLOKy87M0H8obeoCih0LnkNk+BpAAElpSHaJZy2Pqven2Ds+v5l
WHcbyFqwsjX0XfU0iIFjYMEKHwnwKFd210QWhay0qBSSXHZPYxAzRgKPjftHZC4LMd+WeIRiItGO
vWWdtYzyrdi67g7SeelYCpNAXxse8garmxgBTtm8tYUOg2Xwy7ZnvmHXTLTo48PqJpWxIvdu5g9f
4IAJKg7RlCX4FVjUo1x4bQpruZwLmYepRJ7n9XTs15fnPwtGm3bkbm5tQW7cpr/XQETU/XsU1IB1
VCAs4YEaFpkvFRGWy5STI/Lhpn/rZQ8NPeBgWO0NKuU56Rgr9NuNhWj456kU6TllktyMW+o7Onxq
+jfaOqGgPNOiyiV3UKjIczp59oaBHQXomGIWwaHRKY4dTfvs1o3KlfdWMOYduG4Zur/VW7TgZ5eF
YRyYnsGGhcDm4dA+M01pTOsfz0yn3CHkle/232ikkb/AL8Whk7z8ayMOqqpvzPdp72fs3bc81fqN
XZAEhuB2qejGkifQJOewMyZaGFS67IWPryBCc/rNRS39KKw/TgN2+B5r81Qs6N3u3ekd5lF6S6Zm
IL6AxaM2ys0iOtFh/uE+qbClqIGn2ykkg/JMMUm2XTQoBJSb1E8+fpDLixcLKVnswpUoAl9TSTbJ
9XwDsC3oJxVWQedpahb72ZYDLx0VZXfWVDfz+qGyqXmPccGehxjv7wbYBXBJq05mzCqMe/cr/y5n
gGr4NEXSHS94uEBdp8pdzTH9YBh7kGoxncJeMRya323T3iB3vSUD/CIRkG+s6fsWRvlbpT+GS3jU
nvsVRc74vKg3f9lyLEPy4VZhOQ0RoBUAf2pDjGj0aBSpRu6aJY7pVcrHou9mm5hXYxtWmt7saQH4
lLRI6LgoMamxI9Kq6twe8yn8Bq+GiR4LWEPWCkskIAPkO24CWLCSkLQnQVYjvX066SWqHP8lHy2M
M+Csfr0GxvR2/RYbiXjV3yUKVj7mVcuoCXtwikNdpVUcghgqV2lXBczDZCTBQ2DCZnPinkJylGiO
hDbyngMzqJDN5ro2ObVwIEWkiCPcXzZdviJrsrWT5YDiL0b5zC4r8ivd34EBthEVkxKxArhA2Xhi
KcI1GjphEhBW95Zjk3nDs+sIIDySDwvIev5L+kl7u1LYuzKAya1hYQLJ2iPoYa3fbK/PR3RkXRf2
06V5q0ixrv2eA6VgcssdAklAX6dmJEPfVAV08DZGWwJaz6miB6oUU0OkbipX27MfKrF5vRe03Y9+
8qzD8SfvouqJlMEp1sAifVFMc6CgvxL0htF+QqVlSam4aQ6g2EWUm546G3GWMWcFZhkBAQ0WxZC6
uNiZkVpXDsmf2C7SO/HieBs5JempG7Nk1H0MNZiwB7SQoDzYHhQ8wgZSvpZtfiVmbH1X6lMXzBYC
SFUQCl8Ktt8id4gCysGk77My2idHAO7ab6AYIo6fNJS5/cRaT8hbAfzq7iLAsrTItsimoJgGYLQv
heOV4uR1yQJO/dNgovRTaQifBb20iYpLeWsye6+gaNg7a95zCbXbA1M6E7gCKflFL9E7k3G+r4ec
4KhUKrjReUkSj4O4bkco4OTk5jLAWYdr6M31qxkEiaXPae15hHBDyRIRofSjzbmYS6IEj2N4rmxx
QQg0obVBCfoS/pco7LBTrsV3MqyPPpPhXQguUIWHRf1bnvBdel/m/J7Zj6p5BNsrxETVmK8xtrQa
1ve315OlsnbaK6wTQfwQWNOiXGBM/VEHpisXOXNNvWGyYDaEO8SMHJglEoh/3eARMVlLQ9YVNT/h
4qA3PhJuhwjzVZFODaC79Msvg/8tR9NdzeIpT6tUrOHsk9//YHpcEo49I5sRFdBg4tlVASXUxdk7
oEipS88fWCJd/8e6zbQXSsOXDTX1poS7N+3N2/CzM7YHUBxZOrr6wSGkoyWVM7j9t4N5Uy7HKI6X
1i2rebJtScunuPCZXBOpid/VZU22+nLUoRVNMeRfFf0Zm7bKKUfdRmXoMAQtQjEJb6phBACLQTvG
RSulf3sOZsX6FEMiaon/BBfhcyANDTkM+Yifm7g//gMCYLudCNMP9lipaWMVjpzIX9slxTYj+Cuq
66FbmA4GacxF4ClQdbXC3ql4gAArJ+898MZl/mu3vGQodWCGjqNYcyZUcI1cZtQMcaz/dkOlvDNB
eWw2fw7jLsAKGFe7OO58EDV7C7rkng4j+FZGlN+hFQkCROKY1Hy81kQXraUyAX9LlzZi9DGhSitW
MqHdwL+enpFRNq2F1UQohosIE7Qiud2UV5rGXNdbu6bNHrtmr8WvgeFi1XP1SNX+djiyra37vVl2
xg//P2xmYBIsDv0Xr32jt3lNJFYy5S/uHDXREhkLYITSQn0/7NA/NSaJX5Nc4RfY+naS1SLPuazO
FUhEN8+ZDM39hRK+rgRwqVsvC99U1MAkrADmKITasyV/lnB6W2fB3ufXhEFzxXBESLZK8hmmxvPI
NbC0VTN1ztCCM98R+d6uiHIxML/AL2q02aCgfB7nPEcvMuXfPckyYDWCOY8ublHvpOQ8pDSv9FoJ
0nisewf9fgIIELgiO51zlhXwm8E2tEa3UsPgbQCiqZg1L/WFK0OcwnYeD58P3orYBn4q8hLJT+HU
RtKiMblfyAqCQGwxUtGt9I34Una7c/yI/szVOfdulJADEqi3m2up0ASIMqOM/r9f8crRlX/mNgmZ
XImSyyLH1IethbGi6MESvWgbOQWM/UBE/ByHJZD4D36/AMqAOtuRI/OEcj/BNnrt1ToUieDRTeio
nwfWnbWGLgXYZKVfl8LYJTipRcZdDawQvU7nobDvurZwaMeSEwERRSO0+a1FZ7MEmshY2CRY9MH9
2PHXfXGOuTAClp1VxXbNLID8/UuXK93MBfV9OLtMW7YS8oIJnCX5jEmr39Gq2E9krhsCxIQl1FOt
e+e0XOGdxoWhi/5rynDhV4MovIzApALkpIv7oZGRHvz74KazDmKFv9bbDSq5BS8qO5Kp65dLbGdg
aIarbtdufX7tB43qjrbC1AlJcpBF/477GiBz2FyKqraD7NvwgEJ43Lc+RYZ6DyVhbi4LyriAw7Yd
kKtP9AUSIY+Ia7sc5O/figBJXdH+lCneV5ZPtlJ8PUQcUaLzFd/8LYuKOvhRxmTqqrTxKAPNsCTQ
OZuCXyGzfxm7lWgXoesxw5+quSi7mMmj+QXQ6BX99yNN0e1QFnI7Hh+hsisd9RqG0w8T+5ssvtxU
+F6DUKy0PHaA1VjIA4yRKA9pZ/ukTpYfL/xEk2DSTcxGYL0VwYaAv0CwmQ5+j3VIDja9xilh38vV
Dou473Bep+6Kby0laLVWHMca4Yxf+ZirucbTGA4hRzNrKfICxpgzM9A4PDCuKIlCykCyyuDcvY+h
AUtpE/oWngl6q1XsiAoS2txbONDOXxd2z89/q8peCyghwP5j361kCXL9o5NoJ9eHIyaYziRUIYqD
moBVjKXgish+exNY0twg+/3S51FHTHd5K+wiUv/P3DNgWkL+l1LFq3zcmJsUeG4ogELbxw0g/zVm
6ye2WdxUQRMtO6f+EGNwBdA8d+pJxA5BZsIHBqFPIGi3HoHzDxbVEBDTvlQx17gezA5uizuhHgGR
Xqvxy8u7PCpUDnA2vZhlIjWuXynRmNAIUqHhidMFfm8FjESfhH8EKQonDuDVHOivJXtRRTizYlcG
oWAwz3JlM60D4KXSEkMjyB5iOzL1XINxHXWuYA93w43BI9h9mbPmrTQqdvkFQjrILQGS9JavufNs
SOIkQo3CAzZkMGAmeXJsAjESc259i0HJcYrE/bQNEW8mSpKIuo/XEPxy4nFu4otjtZACPbfxmRSi
xCoytAR0ww+PXx+aalWuSaWRTCB+IE1zd2p3r2N6VQlBXyUtAGzNrTlQ00QqocrWOJ2uimgykzsw
gxWIdkoJmC2ng0tbYVn6ixSNVPJVQ+B3Y+s8tBqORf7Qurpa2bMSK80Bq7uEFnZrScxWCP46BBOk
w5ryI2f6Al90nLV7ip9EVbZTgmJdeveu4gOrnKcyJJ79UO6pVrddVlR2sCTYelB2lGoYE+Lz+GvF
BOmCOm98OjBGlmUFJ7ycia0RPkZkpP1axBFUjUkD4la80a0HBNpepR80DbVDxr1ZQZHYKOHPuTIx
+7vE5q8gp1+bf1zKIhd/LxYF17sX3YpEdoywW2p85YbjRmQ5C3KfUlA9FscKM0HUhOVIm32h9DBM
rd2wsvL40cAfwJCjEYblHaFaH/XpZ2Nsr4CFbqQrB/srjcDJRfmZILUYAQX7y1eSamsJoYMVE4wZ
wiByt0/3mQ5qIIcHbybqkhOH9NS0yRcJs+mokutaLakbQqZt/otEFwr/u9PL81oxpR+ignw0NzbF
m8rF+nAPk+bo4YwHEiCJhle2r+FWrk/aWfBigmXTnuzqJ87ATI67VdO5E/ZN8+Vt19fyKTbkFLKB
/4smRYgDKMNKMqbof7RT7NxL8PFCSzNCW++fBojk5Qr5l0yC6UIQ1pWQ1yZlb6hHMxBJtQQNHjS3
lcTwsum3/aLWvj58DJKoy9r3g62G8OS2FPpbI455zakIYtdrg9i1Bk0rgyVCKdW0ad/qyW7om7SW
Bwq8bB4n7RY0Zi+eRxRZM+DhQYBF2HQUskpb8MjQokabT81Vs268H9oBQcFB/ovEBzoJpGfMfRra
w+drLc+N+25YwiS1CF5sk6Ud7W2I0RMeryl9zspc7YFM7A1vyRD1golmnVqQS6reCCX0FAXUN9vo
3m5Gfh0QWimNvcyJd9lCd4YS5sfY6XBMhgKnTgl8RMoIA2jmIUK+0trIFR/79PmWyR8zqv+PUdb2
z4uXUo8q4oExFBsNiedbZJrl0vJezmV1Kf22Ga6ZMdSvgG/fZ4eQBoO2GfaVEK+q7ueapgfQmWUb
ddIRwAdBUMoAmzQu6b10YYtNTtcG+Go3hPpO9FRF48OtwMCcs/Y3eoFdc6P2TgUP3Oj/IpMLuXcG
W2ve6Hr6f0iPA5uBTMB62mIQ95b1Txzuuoj3bExmUxewODiRe2xbk7AJEAnR8cifnYmWJDGQsauG
InPh3ttb+q4vd0B/5c9iCwJaEuWdEEJV0hoj9zwjbNqaOaCr/hxEYFi/2Ndjw4meQN2uxwa4shvL
pdiEnpv4UVgygcBPZNxfK35oudgkdfTzSVql4ynw354vRHcefr4Elr/V8pdjcrAoQOOi80v0103K
aVGOc/yrLz/E+mPSns84m3FDPKbJCOLrRa2xKzQyomBBYIcvsWkqL08+LqfWypg7ep+Qtdsc5Kep
fkS2HyppNfrY85H7RRjHgOB8cr7WfaQNKhSke4D8R3cMf132FNQ4ifYV5NjDWinf7Be1bjPzrRgE
RfJtRa2mp8FDy0GrVO3Q/LZqP0FdU0HU1vRSYrExZLIj5Wz9csjWdj58f70rT0NDwroL0NZXHhzq
jLDDZUS/0YVZ3+8NEXSUa10FSlvXBUA8Rvs+1SzngXwoTXq000iUwuTpUb2ElrjCljJQDCmTYQJ0
oA2vemR54lECaPHkel481+ccN6SEFFOt7ywbnIoGvqFI8o5sk6RHfocEJ/fytSMPSSFmWN1CZw1W
f8uyTi2DniAfd+Nd6NFqspdOznur4m0IAMr5WeuHR49gsB9lMw+pl+ReqzVgxL3WjorLwUJazhdb
AoVvW18b/eX0d3TH/PL2liSOr7qGx14c0ZD3xru/UcpmnvoxemicH/kKdpxk/mEe/lkjuS5kVfGa
uSV5Uxye7vTQIdcPlFzYuh3DdF2WBQmxjnsNm8RZoRN8yb6mO0AR2MhzrcoKEuZL6h+JC5cu868Q
97SrQ48HfkDcU7AGHcTkQ9bd2FgySOXYoet9644TXmEfRU5hT9v74N/+UECRtcvKVFE+jblQUMoj
w/3UF4X8yby8mi2RaHHJRjzRCJG7UG0OAeRbiuQ2TrZHs1pt03t1grpTZeV6FJleAds9tD9OGWMF
X2aYXy0UTJdPKDzzF4/Q7wGD9P3w6QEHJZMQfFb/vMy8MStLSKtzYMyGIVRZK9+tQwEivp0NR02+
tG0+5k8K4Z2bzh2zQt9eosLbVPMMmvlBWsbIx4oRctWkxaNmMx3hJ4NbYv1cBqIpyDaNbK257jr7
U29jmrdH2tsBFJNpVo1RZGy6s/ih/NRz6yTDjdSlSu3vaJT7p3TQOK+qiS7tY1/Za6oVUr37IoZJ
Vmu9+6dV/IZjPpueSzQ4qoq5Tk7X9LATa7dT37Wg5a9CxvqOjtu2O1aZu1pExrkcXgQB22K003uC
R9oXw6iYruaNy47zWELXoOyz2ULUxn5fSjLkkwwUftcCcrm27pn8/0VkigAnpsqO1hdqV14Kof3p
HbKIunMSdR2q3wPhQ4+tsxqHQLW9NJWRwPB+/ZRujdybMsyC2qV/yGcE5lc7qLYbE47qOfvSRTvC
HzEG2AEnAen02nPP7L/G3mwyVhMahHGp5q3Ad0+i2wFQjPbCy7yFyyb54kWZsx2xSQ7oVr6+e6y2
5rhWFGCbg+QrBjTosp/7I9OEwHmg5PGNSo0Tz1YLa9mrvBCL+rt1PP2EaByVhi/i2es63zBboew/
cTwjCmDvKsGQpyTWbV08FjEfx4ZyKxvjTrl03/AvN8tAzVT/sln6+xEH67vNSJFRLOFPZGKxVnfp
AInjU0tBvX9ysZWHCgOzEBd6cR7pb0EHGaiiSnbnF7RNLEx0z5APhjPaI9EJf8on5v0DiaZTJhcC
+iVpGL+uaQR/EMxyYWOJECadhjbYYQjxqtVpdiUfZPZSLx5Uj9tq4NprrFas821fAE/toea13K+R
KOjy6vtCc6GvSRIR9UgfGZAEFy36RKf8Z903+nkf79MSxJ6+pbhbi9ZLedNO9or4PSJaYp6fW0bJ
Iwe1y0qNmW3LePuQird0gFh0ZBjDRbhAfoHVnLBdfQUT9803DcMR2Bo6omZyxcW7o9Qbq1z30hU2
96d/O7DM1lfnfsWJgOn52iDQ5ejq/wnvPjLdCws1TIxyXzg1Hg+j1UvOY8v5Rs5HoxGPkWoAAYaR
RZ5K+r4zOjCvG4mD43KPlLdqq+tQXbi4H0f6qUCxXhx4KXoBF3IvbaarvGc2wW7M6kLBgdHCb1Ll
qVbgLEL4j72SrKl20UZFIiYeIWoxp6Ozj1VP84LZLjrgtbfhk+hVFqYRmvoqJMA9Tufqbolh625Q
IlSr1DyPTwYqp/Dor2Z11yMz5zgxq4gH2GKugaQFTWkrcCzRPGoHBMBfFS+Qhwq+98/lp/r+WQVj
WLCa3ETWj2fShZh/WxLzIkjbW/1Jx8T+vacYYdnjZhVun3IpyDjJ9v9jUT2pvr6UUeRpMokprP2h
flp8fVcd/4kG1e/UM3XSiaP/99iH05QRooYvI9wiln0LAlX2zZKMDsClD7d/rxKk/hKdbplBiTz4
S0dlKH/UBd4VsOkt1GkUDGgKHCXRd87kYnlfTJmlOMB43RWbABlXQRmYAqPDaMaB6F/j6nsCOMPO
xYQNB1gbZEU1IvSOlCtMQrPA9AdXGXkBLcccY11kKVYj75yF9lrQ9ckhtN5gZ+Qf6Hrpf9a0qz/9
TBM/B6/R9e3VtdeQZBWs90E4hoKAdwHAs1p6i2rG1pU29AHmMTnQq0oZdZ9qSTibc9a4Jrkcyky0
H3rK4CjmKsMbeiWA2q8xQ3TdpZaAhF+VIaiWiCtE1+gm1EMBc+UQlPq7MsvchjhAATmdUFyN/fe1
7SUrm3k1aZhcLlF6MSEkbLe1K8NIJpvA2VRzzLKgiV+8uRb2NlDXA1C+jjj5WcIH2fZmC6CVT3Df
qDnAKzt2y8Tm7TOBhkFEBzw0apSdhDZNlz+O78ULY/9x0NvCWEtwIKDS0RLy/qGLlEkvlumfJ2lB
dlgYuWBy7dW3+NW881s3/NgbK2yUpnOxo2ryUmFAwL90IU+vVCklbXO3ynEpzf/MH6CrncWspxje
tWESpyLpmCwZ2bWfCu6ALyHmv9X7xWAfouyJV9cmkXF5ROtKnJ9XSQ3mJ6HBggSGOpwNKZPSqvBf
bAAWI825XsnFSiO2qUh10XZeaTT3LFOy2waxJUtJJbRYHiGweR1jwZ3RI+9TGvjGwvcMZ+2bPy8J
PVqT6+zKxnoZ5RmfdCzOJqpCkTD2N89MFI78b5iAINaZmBs2FMJYoupVqqqf04x7hxGVQMVrbucn
pmGR/dho0BohftDNoqFAjB2RB3yqF41f0gpF6kXdwqs+XFqmAAT5V/iGOXzRFkS37MFzk1eStlRT
gFpmfGhuDRVQzf/hy7D3ZT+V8lo8s36s33qtxigmFZI8J2U3VxuD9gVHEqtaA3bvlF5JGL1A+6Ve
TIdPZKHtZfAp6wx7rQG5yvWoTy6N3uWbG18BypU+PY89BNWGPkAm7Vm/8KdHAxC2frbsTSHHH3HA
3PBJ9YUD93aNb+7tqkMZknDD1MzDq/ChPZue6Yewt/b10Jl8ecuqrK6m206LVM3Mo1HwSJQjfAq0
te8XGOWgf4tbbuGu7DiRjQMa45uGABTbqoG4yeqhgIg2xBPSAj+0SlHyrD1ZWpQSUVKRliQBS6kj
aBxWw3Y+Tj0oS7aMo2SoZaeATnxJSSwKxSRHqb/IUBBZJRjuFiI9l4SMLkkM6L/xqugWhxYneAzR
nShL8AurgNqnp17lVLfmnOesdGNRiKJw//RL2n0TrMx493UAROoLimpe3kMo+YQVff33IHwkv+fY
hu/gPc1+wG6Gyi3U5+LqvxEJIvIZ+tHdsYKm9/4ntQ1TiMBbK8nuL6dWqI4Ace80949rQ60JfZl/
4bZcuU+A2+eGBJJBNOeHRboDijmep4hOsuAg4ELgnpTH8n2JNkFw1k/UqJuhYLoCA76vN/3mj+1+
JXj4MxbHTJdmj7TVfcN3fxHHCiwzM9M27zpc7zw9QJt1thKgQoXoaBvzVEYg5IVv+DB352Pth1cu
gBkj7MAT2UeDYvSkruq23FZI9igQy8QAdyT1cO1emunbbyGSQEvrUCVxV3B+O34S+lJjr5W5QuD0
edEQfDkHzo2oWjM19duul7IWqpWkm6q93jhtJYqtFHnDouLEFXK9oJrDLNXQihAOPfbPK2dHl7WY
BDCNHgU+54A3tLgEy67xdsUAeoXwjdOP3OKj00wQrDBmO/Vs918KWOLU8fAkCMVNytlceJxmtB3S
K9jCrnCyLRLjplkK1G+PCSF1W2ecUjg3En3QhHpKcTskQ6pI6Ir8NgwFBe5Xx9dvyzsXVnvZnQfO
tx8yRbcwMrQbhXoTf3/fhTggGANzP2onrby2hF1kNVo1OUj7tLQpyCr4BcBhVifBrJN5z6BGvQQk
w80M0q9b6H00JDFPOgmjmaTQk32jK6rKeAakIERCtQQ4QSJdQtEmOTdaSLTqFrKV7k969noOER7g
b5hP3UzYaPsReR4m02tjfcpNJuTQ0WEWl8beYWJmvtEUL0r8luPGHbKqEvy81Apm0ZBjZpuLz0fx
VzTbt3l+kY4Pyxi6xdrhbeZ1FxlrU9RmACO5Ej3CXpM8OITiDRZIVwa/f/RDvRn2g6QZoET4HvIP
Aa1/vPTJVyKCB2thNZFCC6v7bKtQ8RbIiue1GwfJbNuHXgoDWVj4vAhYGFWR4esEwRsBBV9qd5wg
RT+zpT8PxNGuOTJN111zPpyvh5kAuvgZinr5wMpXmW/n8ocByaCmZ0lpXyPm9oufJS+H+Ri2dw9n
+TTy+XiDLFz3enazbStJLCiGPzacrFV5sCV1EljtbUpp4/Pf0uEIxydYh7swph/oKLz2Eiebsb/Z
VEZFL74vSfkdQX5xXW3z2esSdlCBBq02BAI2ptRlXBzU3OY5RmpkO0c20HAEW0F+TmWVHe0LhHKm
4QoMxjaDW+kyrGJFwAQFl6lwUQdVNHqxnkkgCUEocWoyHPLqNnMYlEbNtJKNu3RmufCtApGAcXCK
RBg1yMlcM6ilsCRrVq+2Bwdzs7N+Rz7eBYMdO1JtDjErZHdinu1+SABjIJUBL4RROpqZDRMIXJME
OxNKCBDhp2FAxrM4cxEk+F60PaspE4gA+cB6QAv0z7Fy3F3cdgP+idMrq/RvJdTNjTwGiNEe57Bc
4/lsRKX30pJCyam9zLRCpRAGCw5FWvWGdrz4JTXdrm3KMgFuy1yOCrnhYeD+SVDYmowtfoaEz+C7
PSxLcZz0LLkn28yZb3QZMXZfA6IhAQnG56dax/sDWTCPRQ58kTNNnZCXpVZSUDC9Sp9JmXwkJq7W
MgmQ1TTiIaPvvKUJm9lDJKpLvgOH9hoS2M3GcYrywFZwZpGh3+7WHyU4jPj0u/RSXdTjmjo8YQY7
btN5ju5LigGueiM4I/5EFMHF0Gxe0eTddd0nAct8xk3ZmTGh9+/j66nAQra/ttix9NGD0YYafgRa
kifp3JYusVlGYX+VArvRdwCwRY7DD4BNEK19UDsLpCs4MOdrxxGqnEaeQRE3b4B1/Kf/gCxHTsim
dTUgSPqd2iZzHY1IE7+oucxCk1bkwTh9pCKqlQDMQXL1Uh5ZhyY1LpIx8OnLWLCNqibjEFV+Gzd1
ONVtVsedzlzIYStn2yg0V+rmO+feH2LWWW7Ogv0wYlBuMDyebKjX0CEOM1Bifnjq7SSGNqvizG+c
cMjRN+z19rOBXnxnlBi/XZg1K+hIBd9xgiuSjApKCv8GZdYThkgZASkH2AXVCRC+qYE6pEbIbjok
fzEnXQqIbVObT52ak1+21Nz7xAX6ef0RSZOLGYcNaNwj0H8p76JQCiMy7y0KO1djpyNtaJi0w3x8
NEV3Yr5WSxZeGWrpanA82ivD8Tl2LOkrwB+egPEbnWjX9mEYeD0PwP1vkOFHQE1Zo2QDYYiLdG1A
RH+Z2po4lPo4Z86w1KaadiIIV7ENncmGslQ9l5gqQoM2rlyAYc153iS7QD1yyn7bY9bIBpLBSrmq
fkQ1cKpW0YJaOncOR7RUSMF46qm7W+mzW7gnjCDtw7tKX/lZjARnH2aPKn9vNbywYKv4dIxbksMX
RfBWKVFk470ck0rYx1oDMVPbsyTvg8kcbYCitFXg14336OCrXt+UIw5tS9ZZrk/HBLXoyRiRe8MH
BsQgRHpoD/4pWJ17i619a8rAKAXfsnY1chYszipY9iyTT7SK8lYYdLrcpXYv3SO7DFHY7WBtVyzF
2nLEvocPNXDN94U9RQ/+oAHuawE+vdU1Z+IvuB6CJF/YGIM+Q3P+RsTvqSd4AgNE11BIlJKk+qBp
lYQJGtxs7igTz2Fp10oQ4qwBYZjl1WW5mElhMAGd2MIrafXNXJ77pU0bSCahL2L1+OdsF6+Hxfpp
9d/MWKYDPM7KAiY5j/tkR6ITjXkX9gJj4ZQTJ0Tck8KZNZCye3p6bbMPx0Sq2ZmHE/rhBE/8IPbY
rUdWkNq+mJR6tFJHU6tLKHj3F4nf+P9ug1IA3DD/h7EkgXwE6VgSmdzAzRVkQl3WM1rAzTG/UHuI
93t4mm0Kue/OHewFWu+ZYXLZDsRhhMpx+vyEf4K+oJWKgvSJIzccUcBDnvL/JKadCxIW7D3PhV60
bZeFWtDzP4u6neSoOK8T/n+ChowaPlIJM23+QH4/4ZwsTRlZrfVH7PEBdHUDR90T7hJYf9NQ5ZHx
pb7nQnzXXuIoALd5cHARGO2r00Tq56cno++Cs5jI33Ng4aELWieZRqe2YzZ1sw/cZxi/wfObaqHy
yZR7ZAueYc0SeZESMmbRZRX0oDLyVwkGzBYw7MmdVW/GvQshA1ALgwIKMIPo95JIt8Tn9DMpOweY
6ztsKFg9OQPxIEroIUI9jg57yF3UxGctkKr+7xHJBTQCA9mtiOB/CZqTckiPqipufnQAD6mSFfWA
dSleVY8bGA5lg4lRC8PPj7xz5E/SM/d6YpQVg080LE/NYVXxaIAExVrsUSccUGbjA3a20lXhNmae
xJc8p53Rk3UHwRfwOHomCotjd8tqdGYnQnUy9tINAQxMItI3X+eSQrreqt8LrIf8PJ2p2DZSlQ0h
8bqHyqVMZVEZvex7CAabwMV9TQk3pi/gXMbFSfDqK1umm9sSqKBj5WVJZjhmgHR2PkB5vc3vK0Wo
Uvc6AFCOd27rhsbpbD2lpMRhLLGJAA9y3pQFxPunxEpRrkmnFFWaMMkD6qbVpJ7VvpIGMef3a8JM
wn2Jl0HOVGXPUTuHSrl7Pq/KUHreREZ8KSHLEiWFbFJFokeMroaH1bn8PZmY0dYiAPrMJcM/WwlM
YxOUXkaIQOw+Dqdb8hSQ+9L2GtYlZ83VMor55Hyo6J3Ehy71JovkKK0pSFipZ40CVmUareQkHspe
UaC0Km0hYpnSCqZyiX6MrkEREuiLR+Qiz8SSR/m3imoNdSfnxK4qIXILbH+jYfKcY1teR3YajrC6
1Lh5C38LArR8hDXBjBkU/Fg9aHkltY3gzWOLqY9ixOPO42cxLpifrZLwpaY5ZzBKKjLTst0qm9Bh
9yV+GdeIeCxxunuIu8QEeti0DibUamEXfXbRHbJWvguYC6QzBRwBt6yutfiANHMeajOzb+Iif5y9
8dnS57j16UMBvK5fmGvjsf38F8Ui4Q2hmpbbWnjY5Sw68OoLGZ1HgIzbHhqfyUWAMdtg7S4DWWS9
x8ibiGE2l6Qq8XqPmzv16WyRXG/nnj09qa/iizyhq3NnZkMkDK/GH+2k4kpZRpCkufE8JOiX2Cgi
cIY00phJHedS9wNe0byYELSMbq1KMiFelMF+vvtMmkIXCCGDYVPzdO9k7+r+vDYu+fOOfWVh+erq
6tiAflUoZyGcoweN+1YhAfTCWdMBXrg4RXdmj9tl39v0+xeDxYv8vn+TH1QZbwMQVqZuOgQ9vUt6
XNOIzEFu73OeJ3/slTpe9TZRa6PweNsKqo7yeFmClRsM/1tce1J2qQyrXH1R5N+G0Pz9QA3HQN57
50oPs9Yw/Bu96ZGjLwglUWnqAiz23NwzHXwkVAneVG7mUnaJ+Khc5+QcqNjbOIDCmyjxCnyGxaIc
pxKHxeEX0arATxnIGp+Nh0L4j2LXrqXi2w7khYt3Gs4yU6/C3pzSFDp9IescEXNlu8U6Iv6NtsRp
/8NgMu8H7iI9HOn1wvAUjmgvJscGl7zzlAz6fwrJx1Mls2WaOzGBwhyIy1HUAeaCpCGoETwJUhov
It60Q6JQM7UjwdGUJt0OWwMe7yukBlc9YZy0ngrVeGOVsiuKBZzno6RupMb2r7xHEQH/y/yJeaLg
YHbx1TNuqIfJjG2XPfHqNH6rXXDyAA2KdJYWi7elnnbuDtZ0WlNtthM9I7hrIiLvoxrFhA8VI102
B/bVUBx2pUX276CzYWFONx5RXROsgS4Jq9V9JpQ7T3lTRNlhch3+LEBDNCzacq+8LR6FbsH2Ft7O
aVkSmmQbFUXqhsECIEfUih4O3NnkG7kJwfvAznYVJTl9SnVKmUd9+mxnfT7dMSXC8x6J1ZsmPORu
xrxn/DBsgrJ6BJRce/Ly0s9p+dlmpwPAvWXswBVKMui23ySf4UWSrkEzDW/x5kAoByNXAaM+M3Yo
Hpqe1Yjqrq6BQ46b5wNeI0I1gywQICI+ZwYevpA9JWxgf4dKmAMUlWFkPElMqgOyH7sRH7lORrgO
S2xIgmWJdLc+Qp01E9ABEci0SmARnxiiDpie8x3lWsIkgBAQO+nDGti/C39MXwYpHV2fWS5N+dW0
bcczcM+D+P8HZ4jaU8k5SbDNEjAWEx5i7ZFR/wxDepkgDXvfP7V1VQkgQTVbUtJNFvK3TSPJcvWp
qk2QPyn4+fQcewwDvIHbrHwaPB9zaOvoLPiLm+5OHIbuG40YuwLohSaRddX4FPWo37S9jhdYhIs0
LwfKL4P+DeV+jzXbNWno6BOb1pMjZEI4IALXZCn6eeTQnivu2ia+YLD3qj1RE8nN8R328+h2yJOd
ssUkLLsb4CR49oe0vdtOgNhLwS+QnPukBui/w61a4Ejy6dw+vz+TVXw+ESeoq5KNmGydXJ55aWYZ
Zcz4qEr2/jYqUT73GArZFdru7f38xcp6b6A0y6YJqanxhX+liTt9hJzEeFK+PqFLkuAXzuDyaDe1
7S/ALUaU+1D3z7ctpzSFsHbL4euB5duKgxeJ5cIY3ntgYzXNhnaNa2y1khR2yyN917WvM+0px3LU
qpDRw4Up6jWJtF0Jlu94nnbxC7W5l0VwMJxCraXWietYIVX38eRXL6BogwYvR7ihSHDqozspTbhE
/UBsM4PIbzTxRG/tKgfPeijPbD5Qoh4yvSpSXsy25E7SiAhwalRww87UjN1V/GWzsR3bSAf4nHZo
12050YNL+Zm5K2zkSO0xC1yebg/ky2AS/0KUlGUp+UGR2Y6Gls9KXJCE2BWniylxwd4Vi0HLoOVG
ksKqCVzSJeB86I1ZQjDrK06qCPH6XXLgi4oKx7LMEfsZTPqmyWoJX/xnNGDEK/TEU/jvmyiX/uyA
lDQIOdEtL2AnRBQfD+lCY3FAn5AnCvCAyAa96DTn1NVQvg/37EFHGnTaibBbKViBW66L+2Zbqs9S
wzJjdm/MbHSu8ZOwZv4PMMRpFzBM6/eQdS5ofBwNy7SKnGpodCLIQGJquW3PinHv+wJA+YeDD7+i
9pqQAq1jbQ6e0sfLVmaW+TPkH2dyDc/vdzQLgQ9h/V5383O8cRIOczDCCc0I4xE8UniemfLp8l/k
C/QVhMKKOiP8aYqPT7XOap3PLG1CxODQ8wDQYrEovVcjjyKfr4mJg9GIiabchvtL0PI+SRTPYvea
XfwE0aZLrqBXWugU2PpGgPMyN55O5bkl5ml9Sk3ygBIauCWtqSpfhwgiJ3P34yTJv16Q4KEMhfLT
dGsyji7xf4TjEw+0Y0WX757k/Z1sYaQQR5shJZjboxzVfNt/+qZDHlDvKRF0kyjjQPn7YM7F8Pm5
b5vX/oOod+rYI86tF4A/5UnqDATeT7WMQHtpy33dD3lT1Scvut3Ksk7Wd+Dkflpm+Ydzrc1zOuGl
kywZFnq7C+Cqf3+5FsyLFZdbAB1vE4STRrRij54H/0wTejPr0Yj5G+YUjysNvCrLNsI7dXH2F0im
BSC3I3ia33yb9bwx6Gb2gSCmTDzcz5fv3QuvtixylBjrUS1mTDAFuis3ihZ44TcS+jNmAP4Vnu2x
yQEPCRAWhx/q4xPgJvTVGHIMWPLizajD3NfAqNL7pt4gUZfZk+s5lBoqRUajkTUTH/k9yibWMHQq
E5kOxB9fsrYaceb9qjAxdzmUTR2WITDbqT+1BAYTa9EHvsC7Ipui57m2Om22A2C35ykIFztrmH+B
uU296KSiXlEKaXT2COYptfSmMFOtrtmXu9yrVGuGMifA2RZN2TOqx1Jjbf9KZSWn73u4PBmRC/2C
z/GVVn91F+7aJIHyr1VnYa+E7yzTMu/vJa9kOvy9fdTlCs+7xIM7gyHj9UXkO4I+2EXK+INEivvB
Wos4djFJy9STjb4v3Z6kgNfoIspitS1R+7OvSkd5ljTe1Uu0P7/qvWtvTrWR2SdLS9lmTAyibvNE
Hi0IFdBbbDXgKSCS5U0d2x8cgtpkL6IL3R5hn6PpY/4pp0GO6o/xCOzuGOXkJWlpi6fkxqavoudl
hBtgdciURsEr3H784PRmpZ0D8UupfoVn5NHrPLXZqki6vAua4YlKjtCAzpTCRKiqb4W9kJFuMneN
hICmtUR8n+RxOOdfFkojMGvBuQY3qTylmMgYFihv25nzYgOqvjGrs8VR1cKBts5AGqj4sjvphmoi
65CfoGQzDK/mIP14MU0m+QYM/IuesP2PupoESc/ZhF25fX8tPIlMQX9SxvOgohQv1s01FtF/3ts5
2yvaGQYmapmHQiW6OyZNswGPBVrcmvPmwK73puVTFUZQZiWoKjnP5a5rOJnCAXIA5+bNHQgXe8Fa
UUGs/1mAZdB1iKcy5wu+c1gibJYW9fyEh8qYsqNDw65mF6Y4c5D2zIdGrUyfffGykOevntD8N21L
Ylqwd5rn8ryMmP1cgxZsfHSexTp+p0uPyZOp5runSMHsX6WneLPnQgQSv+DzhD2G2m2vI6SxaAVz
d6sQzsGJqEF809jzpKtb2CzAgRZ5LNu9bkhtTqq3Gs2akkYx/R7Gut5CG4oc5661vsx0pU4TBSZJ
BYv1qXgx4vucuvUCQzp1KJlR10gZXjhMi7t0MvBsmp3cmaH3a/XtFGGnNj5So6u6rqGil8KqLHiB
pxlv0mzK1z0q07o1NxXgMyDmfYVe+vODNQIjo2rcd4j/L/LYkgTaIXysHr7AHrZTpDh2Zh1W94cs
KrgCfnsJspdsJmFnTd8kGPJbqNYymm23eZfFnRAS/rqBPrgsxbWDsu6+vKuYmiO46rbhot7VYT40
PohEYCk6OZM1aTwZnuT/keC2nmWBO39zcwp36ifEqdpmLOVz+hwUGG8nvWI4nEHLiX4/ri3NmCKj
vGc0dw0dp+wfzRkljS50ZvJfB1DGiRiUBKggrlqtywELCr81cd0vLIZ7fQxON+xtEGyi1v5kaks5
KHCi5HJWiEifZXY/xXhVyiMclSJvndsSqhsH8kfMlr4u9Y7jziIUTlr3zl3ovfDlTtl8afvNIG5A
wJxXbW8mBP1tqOrl53n14aAlnbtqGJuA8Or11IstB5RXmssAU+HNWZQW+10lspxiGGWUMIDO+hGX
FlIzbIkRO5/qRp2pa7xNigX3C9GC9rQE5RPVkVOkhcRlYazOEKhjI+wPSrOa/fa9+UcbKv1MQJHn
IFSogpacwSs3cey1G1956OfyC4a9bPmypnOqOgLNuOuvAvc6w9u/R2WJ4RwyQwGgFBoHq9fohoxQ
qtw7M33dPYovEEGUzCqnYlAANq2CbSqj6als4jE0jIPJekNK7h/RxjZ8RbzT0p6bXOsWmmTMCHw1
h4557fPpmkrEl3PXvHkGMzvmZNmbOCN3iG1rgT2ZEtsFA9cZ6qKbPWcpVCW5kMED4/8CAWrY8ejJ
Yhgx514J5SJbv5COIVOKTV+SLAriyt9o4vFDc0nF9bdEL71YmgBXDK/rgGhRQRastp92BX2J8WHa
k+XTlR8MBuw3PmnFN2GhOOQYU77iGWVZKDlFyNduSIWwGoVkMdTEqlIQwlo6nOB3ZuKYVO7Y5wQR
THN4AnnFmkaYxqfjvFRF6aKDwRjQK6CgFnHrFluw3a+H2yw1zIapAJ17dJzVGfp+cEOGvMMCsXGc
vkmlFMesCk+a/7F4Sgar5alPCR8htauyAUAmvMQgHOqI/aSq3dzgVOWZJdWvfx6OE7wCBFg+w7ju
1rzDM3PrI+gOimGhb2CoLurZE8F4p7T37t5tNhiHBr6jEtRroi/LQKSaJk0fyJwDcc6kJarYVYor
Bq3wxeEFJrXey6/vbVkEYJBizrCkeJEOKiGpoB499Mo7UXEARk7XtPxDFMNwGEOLoxLLQPfE2RIY
y+BfbO5cj0yU3X6X7nacku/o1MxtDwW4DTt8LTRNp4//x6ZBrnVtQBciItqJQVkWL/DXo88fRG0k
Sunpa4G5BOqssSyAetffLCe6iZHYg0C6CkEoprXdkaluRHLbQ1W46dB5tHvKU1Dxn4nCly9usiM0
MNfVv7OW74MP5eY5iy3c/2YKQvL947eSVUu9HnhKB9ZaaWJ6oLTbM/YGzkZrCUDquhQzwj7UNXL1
2X7r+hOniifnf7zpl+bvqFHvC4UDZ8CkwJDwMgqkya7dbrGFyj+gLrAW/T0IOyK/IXZsIzd7DjR3
sKD5LkFiM3/IcE9mCJ32Za/sf8pequJg2MysrgQ8JzKW09thy8zL2JRwBMKn8LwvxMXSMuxUp3EB
/l1L1NP2FlYpNaxBTeh05ME7aTq/qjWgpDgP4DJ24WIVWGqD957bHL+hnpJj3KwvkXcl3DU6bjSp
uA3X3gpemYtTYL7MZazAOVPQrpWZfqvOltkjT4v+OSzCLO0bve1Qtp8K7HRZoRUlIZzlnkRMdsIi
PZn0Q6a9QqyTJ0w6SHHdFiMCELLXF5gaUOORzUET43ew8aN0rEL42yxmIYhuL55gtXxp3Z4miZMv
TlR6bLG68rZTXlcA7C0Axg4Ktwmx/bnUj8+IoUAPSPtw+zEQ0663dSPfEHRZbUpoXFLizyKf+oAe
KWDJTxJSglITUtn0Xq/at+dPmTwlRECv5J1uz1YhCbwwJzDSS6fqKptVi85EwcXg43Ed6y1EScUc
ZIAe8rEpH3cOO2FAkXODsgsnLKybsWXlSSXsCSHFNku/i6vLPTP5ZVEHmuDwQv2AUUJBRIxysxGt
GiDkxuj83ZKTFIyXZISsYKTDuHmZqAqUbcqQM/yTDJyZJz7HtWV5R+/rNxSZGs96quXUYtgoKLfy
sckX04UHRHHiuKb6NOhmelY7oZXhJuXTihdaSfh6RU3UkY3Zqy3FNu17XORgam/g5wuHHMCI7fEM
KNT6UuLbwFs50QP1xqNcBNAxIWwcxHADTRR1qylHpZa5hRGcrGHgtpXwd28EMqla6KpYPlxJXLNn
ps9PdEI++oq8zVfHj6qob+3UUWXIdVKZe0pBqOqqbpBE3+Ldz4O+GwgkJvqxbAZnSj0z58hvYY0z
2NT1gWFdQ/IP51wfZpdr0ozQIcOm5EAfM6qKSMZpR2cval7YuBouhHv32myL32MlwewO8B9FjffU
eHb1FBwTb9kdq6WZu7uFIVdj2yU+ReGYU6HJZeTEIswXYxmBChFWtQ9n0Uou02Mg/9RU4rMzZ7mo
mfgcOThLfqOug2vRPq0GHYxnlkrYvhWGyEWrQRcgJeUo5Cm5EGKJZouPkY1ax+dpaCKRVhiSE8w9
7buC6QKE8IIf78Lnw1f6lPXf9LRp1yBd4cZkuAcVyiC34vFd/Bfjk+62PyPRBwSj0qrWlA1AxPQL
4lsuG+8TSyLgczYvEiUWgH4nIDuu5geMoZMhuq45Tja+6UIf+Sob/d7BhioeBDv5KlNhizt/I+25
ju2dfdeAETTIqo55BgYnMQ511NqlqJ9jTxe5uWSEU0dVs0wFIVGa8rjOWkgG1lDxm4DNYhKAqe5N
CBOXvYnSHzu9vzpTH8uy53h4Nbd5eykBHJQmklqn1P5Mv/eOo6jKkhozGLbpECF9GyZpC80mUh0j
Abo+j6h0Q6mbzIuWzPjL6ioEiaMCdPxdaXMG92bdYmq+WhS7ZrW0QNSBM9PwX93rdfNNbHXIGrhi
XKl22+1J8I9ni93YcmttuGlRHdSnDw5Cp/tWUgKiaFWDHlgR1kfNdONMPaXcDSdzqyRDkyMqmZMU
LziucPyBYmcukc/LVguxv3vXgvG+Uf8PHjgTVwI0tADHmwfimcqXOwYvUK+OCjoLetaHFuVbHNEe
ELulE+NSAMGZtJpPRNdrEuFb+JQPe3B2iPlMTcvfMCJUHL5a0MFXs//hPggRkd30pEElt/dUiyZ8
6vmpsUiIuEUOgUU+OYIau+6KMsSvwyJoYTeeFp+sMrz1VwOWcIaNlloIR5iY4v3Lm1rPsnQVUwgi
HqU5eHmStb1sbHM/TMRz2ZCXbOhvBU8QBWRomskA7RdIPL0r4T2YI14e7VNTdum/9OOtVjGZUmwn
50INNVL/V52FyUDS2vJ1BVUH4KgzPQO5rynvneXyAOtb+p1nn6k0jL/naT3e1l0cR/sDBR4vraJW
Ywp2/YQi5Kx9In8/UkDjxiwWoAt00en62fo/p5kzwKunelHd9XVk4ZVJYqFTtO4wpaEzqeEwIzij
m3RqzGuTCwYvyV5GRsJNTr5nC6TC0P61XUNtEUGKEOMNn0Nt6wN3b2mkVIW1eeZg7aEj1xcUgz1F
yygbHU1KCEUJqnU/qNn2/YyaH1c5io/5i3scuYJ1mW1S1IxIkfcuPf+41Xb1eInkuCrBTvsTquWP
ihU6V+pqhyK7VeLL5yoZCggLLL+4ljDVTeTxQYZtNY7oloK85ZhQgJ6H6P/g3kBgrFmNOW2oO082
pj1eJhApfSzgfaUSQQAClq+dR6wPNyGCAAGMKaL1X4qvwTG9KelBZ8FnmYeWmQelxmhYN16c6HKy
gspD59f8gH5Yy8HZfJ8byn2bJPnQUS66ti9u43/ZXh2Wey1V+i8eSv9vYsFNA2nWpEjhy94wqPQO
ITAljwqLIcJpIjiU99SsNSu2eH5h29TMDTrLIEHnsPnEet8ZCDP04FBGo/ud8jZW/TgvtKKdsN33
J6ICpdcjFWNt6KGBEn2extghx/AF/D/BooUQfQmJMUczlmPZee1NfR7XZ3lQAV9F4Iu1Y/yBdXnm
CYBFmXFVuP0v1DOXw0OaUNiPOZ6owhGOR4TNOnW9w9prmLJw5tQuXsORyP+bilo95XwJP41YBuT4
Ao5py/9D/uGURyVBrn/GSrmKWojMkC+uh+ICZ4a6zoCKIXRyPvksYoCLV0/bD84gXhzKdNV9VU3/
2rnbGBGFwtpVK3LL1zNMiZ7ZR0t38H/PtDXVvNa9NSeR2wweTARgXqMqvj88WLiQWnc69wRBIQAs
d1q2yFjBPhJ7Cd5W+ZkweBWE43/kWGkdATyB7jzPhSBlowU3IcTxxyxlW/wTzAZu+DkdoIzbAKO4
c5tCGOzpgUSk6RKf+vGY3gqijL5D+/RpC3MiA2kRB+fsTUK91zB50CWiz8SButhTQBYMhdm1r8by
No79CQsAGHUe+R/xFgF+aLAmBpSMNTvLwGOR1s/ABEMIM9hy7H/+BIDWTJS14uS5cEAE9U1YfTrK
19uZTA7Xxp9OP/MAez1f69B8N1x/Ni3Zt4wHhL51fdtK6IgvCOONvKcN1yum/MFBadie8YSN6oF7
maMDYEr/+CAae4n9ZsT124Vb3RJZSY6/zL5gKRSjV5Tun2pF+oSoKqhg5E+QTwsjWoNZuI1x0Lnd
9g+dZfBrkr3XBia6vjKWkHcKa3J/19r3lHI7rVPa+4Za/cYJmkLaINXWz6aRBmdD/ciZqF3NeOPD
JCbC3QONEQ10bfzkKiuREUWXKt5o76QiWeGmNRPA4J2yhG6FmKm2NOUvy8IJzJnNchXL2MadBIeY
4PxbunyrUNq78eBsioGk55XleoWVoiuAsqAtVlksc4uyeaECQnwLHWYXq97k2WtUK4Wvh44/eVKw
iRD0JM9Da3M3cgSqurwM604wKzGaXwUao9tHC5ilk7frn4pNkFlaaZeSz/aOEnVQKjwLnHbkPVrn
t3++RTTu1KKdSSbt0bANXVC//fTMW05+iujX1ulwb47mWH78CKeuF0/XoqQ+MRImlbXCwB3j3te1
aQZRyivD1TN6lxdT/rZH07MQyz9SWVwidmXJ+PRmuKCpSUrKYL9GZfubwTuKqw/Un5RarlEN6kQv
rMEkQ3vKCPJ2T74q0jBMjKoV6W1sb7zbmXJg6u1Ts90tHl3oJl8WRran1eCSubLI7OVWKhrcuCnq
7d+BBBW5YL0RkZdAU/Subq6D+Rq8IWMDIJx8UWqXkzZyoo9Y4tLDFhaVQ+xDmc7MNCs+qRJY8ofo
cpJgLWaRivGhajJ3gf3qx69qh7RpO8tsULvIkXFMqtkPMHvNHb+iGyrG6GAoTG6AO5dSSdg0Z4OF
CoIlnGSDcBkizeF0pNX+2z1xoQvbhKgHGakNNAoUxPFB+EzisFQxgi7ovsJzaZ82smXUbQFdYCAw
xCbvB4qPJaLQzje+hlceug05wjmE9DR9fjjcIhUZ3pr6xsSCzbkWJh76LaHMbyYaEaYDO07GXlOP
LxmDTCTFuKluZpNOAoA6yDaWuf2Z5ebKa5NqsQC+uS8aB1QxW8iOl6nGdlgdgr3xZZTth1E3Puts
sYsYNmPX4sL91QpZMNnhiCyqvDjr7XCEMg+YFB8Id0oYjuigCS/MbTBDk/aN/xzdA0DQzHr2d4W+
TiRibDtKziT5VrgsIAstjfC7cn8dqeekNnb4FuRwf5AKUg83ZP81sCQW0p/dnDiCdOvLF0a8ldHb
oDFFJLwiYo0GBQlIGhg9pXliRWAOkkUTRn+OBk9dEq/S8HTr5fBXUXz5bE6blrqqF9F+qXUD8I/7
FlMqfuVNzNy+UmcJI+ULfO3q7P7Fkd4FyoqtQf441XmZDKMaGrjsh8HTsBrnBxmZ+VLsHpW1eVUt
D7gV/uPFN6no7dIUFW7YdOidlHpKYIKq5XrNQZLcBu1DRAPcJB+MnBi8Me6hng1L2JpOD9M8NYRf
e5MYBO0G+P3tpRZGeekcgXU4W71JGexpYJo0VgCzwgRwJweVLI8xr836tHC01jXJqKjPaaKOl4ow
pcx6oBGYd7OvrxRLW2wRXgooGQttzGf7XbedNgL/EYpSc92sRWyjUlGS9595e7+L8ZBD27ll+rKE
qLH6S6WLMce/1h5OfGgEZnmwW2aaZA48opasS8WqNpuhMnZuQTBsUaWYzJUUF+Tix7g+Uqlk8tZg
QSSZJjScv76eBrCmD8QNj6OVErI1jV8j+F2TM1rDL8FoMKXgjW24bB8Kp/KvfBwYptV2nQZ5o0P7
NKwVDKZy/s7tWFE8W8M8HcFgNicoKXNd2La51TQdf9PZ/RLMlbGvwebFnrHEO3L37H/Ssj/qKdJ7
+OTHJIqlfi6KK5THj6pFa46yuu3GjBvcQiN6g0APJxdYVP4o8ZHgeaIOweCEFRUaK/amxEMQojgQ
yNzzzbgbWptnqdJ8jdTdABoL2tDA2bKaaF8AIskKP8UODqr5vCNfoDdG5/Db7Ch4peR4y8FAVi0+
mXX5mIYRmC930hg4s3izJUS+tRP1kU9a4JmtTKU9kTM8dXGEUS6eA5qoE1T0lNK/ingUClC7bPCO
tdpidoeCStI0l7nfyS9KEkFZYP+BdC9TrC0igQ3+pxNx2r2BR/jxQ1ymlzjlTxretUtSURT8KzLO
qEsflMmOOzsM1SXdH4YbeAulHG4mVcnAQeqXy0GTWFz+0YnxP/xxXCBDryJa/JjiUQHY+dwWRdLv
TcndG/G060Bx5SH5wbcN0RJrVHlsP5PRVl1mfa82yPPN/4c9PV66It9xx8TpOKzBCNazckxwzAgf
HqXEptor2DyCYatMeaIt825y4+e3uyoLsPD0j1zRVKpiRFCuzfDqDgFFTp4ss6t0iKP44EcVnYgU
JX2DSuozL7SEWmiJq84BMRLTW0qYBtF2oS4nbIERvY1/uwUmI7jQwDFod5jPAYVASKMKkig0wKOU
qSipGVdu8GERL7ti+vWdoqs3r98mg1eeWX/Mj6+gUnWF2wgszQgnb5vpBPnQKM/vW3Zvk6DXFnBl
t6WlEpv21Gw3Hdf1M/W1u7DTOJoBfqm1sugXbUis0XVAZnPA5fixyqL0/zjZgUzj6fkUwX072mRr
iCy9mkCrkR70DJdFsuq0zsfEgY19oGyneC7/9LBvUjah7PqFGHMXIDNzdzgXWZOi3+DYbZQC1Y4S
rkMsnSP1GWv0Ei1kF0yogaXfuleg5kBGeMz0cCOnz/DpUXpn3ct1Ua43SHCpNOaO/Heh2VxSc03d
zR0WeFhpqxQaJrVZgF5rlwyOE9y7Zpd/BCL0pWGhCXW5YOVBflOfeQSNiU1qhgKSRDKLS6ETcX7C
fIBa3HuyEXZ/x4lIn3pJiAHpeDxeeYXy6nfIhCuYSljy5ksGYdnN0zEMRglhkvBGBCIyIqEzB4JM
0z60UHQZltsWJuESMVUYkuR+nwxkICmQkbiHC5nSHw3mTGLe2rcqnVkpW3ZgvFZkPk6S4IAKsIgY
4i9J2caxwc6LP878COBTAR+NXNwvrG4rGpDmk9h1hpTeg9d8Hioa+HER5HObZwy2O3CXFgIyvCNc
swvEK94b/xDibGiyNgg8JlGZAzpsxFJDFf+jLlOyAmZEbpZuG4GriEpDJGZpKroYkgKpiPZJDUoM
7C/9NrhCNUJD4cx3bBzhgNb+x1Ret8j38OWhTB34Si5YkRHFcUg8EDjlwG7BqF3SVk7Pvbk0U4eg
8qTN98sKEmRMmA8wxbrjC+JykUnuBrBrwandXRyL5AJYoMu/aHzQkjdlF6Xc5jN/+nz5gGAUT3QA
+Ua3m/xJgJFbIO7WVkkgYBF/cH05HWmI+SD9A/qFUiDe4QJ0IYdIfCuvvOcivI5oYv9rlX+H4sUy
ADJsnBmKkRt710xSmAG7XPLAMsz4jRKRKhGztXDvBMjL7nNRmwQxVbOnYVxw8JTOuG+R3NL45Z2J
YcP6/4oMEu9h62XUAxykqnOop5oAENIKgUGVIhnpYPRy9Xmdik0U1m671pHYskx8Rf2amP31V0nS
q7wMBNdYenbBLEUkWYlNLY7i50uE1vcev61VBugI4WRjiXJPGVySj2OYaY+Vu5DtZFarvJcl/CuM
K13AHT9AwJ5CnsIzIJhO6Co0Kk6wJ2NSWiPW/b6Rw3k/4cee1DaSNxdAnO7rJgCAggOAEcH/HeJj
rwfTZ9D7l5QNarTdlpOFV7nuXRmNpU62MQkZR/+/0RFI1DULUyXeykciRvekqElNIB18dYiYaQtr
Trtibu0u+CJtPUYLnc0oVOtX+n2UaitmbPvKjPy4uWDCx5NCwy87cyE1wmy37jtdQS8A4Y5N8PY1
L+cf+Oj4TugnPSRnjDj91+Evmf/RF+ynidXpH7Z2E+NPvP8rXeO8nSAPk6Frkzh5OopmcldvvpWF
A26+MHnenLBvgoFxjXod1c0AUSEY1N2eFwxIg8Q9ZHIoJelCcYIlofi6Tu0CiW9PSbGf69Onn+bO
4ggCzNJNcy8PUqwQFxhEPC1I2SYQu85V6BV/stle9hvjKp8dN0mj5Xglr+mrFPjrncNh2vak0PRw
0X04W5gpO99VqDi5OG4VaRyujYcYXIzVtFpnOGIisFLNGy7+QwpK9Bl3N3kUrUjz5OcRUFl3tbmr
gOMlgCOhK39p2GgGh++fC701EevmJGn8IaZdLkmIPtRkH17qLg93YqdtKFCjLL9yK8llAp3e5T8U
un1THVcbUXlo6S38ajLNH6hh6IuY1upCPzKAGk+s4J1pMGOWShRW9B68OnaXwAJORyijNKHwasUd
HNfNZsVDNVDl3/L86YTlr+62WX+z7pC05GDRE7dWpMRitE0CFXzZlWdCGum8pTKedU0lw1JcNHr5
COSqK1Z0PWRrJM5V28iqIZqfBDVB02aPZEkLoezXUrdLxVWpL1mDK3m6uh05FbFZAcxiKg4MuOmz
70uWT0MGZ5UPhU5gNeB4iE6nV7tXlZVC6lLyvQStKVw5m9AMga9KLnisrXnURSMFz3Nx3HGlV2Ha
d7yF8f4+zpPBvM3eh0KgiSe5p5VgQFTc9YpWVs2VADvwCHIQ2G/GoQ7CvyX177otF1YbwGB8ToF5
MQXQ6xt6ibvfADD/xGhcghMhw7FnMJu2ymsvb8Txu8Aha+zaeTE3UhicP8pkWBlIXKy4Ho7n3wTk
otadAUnm+6+PumbOgCKfI5f5V4Kgybu+A6tCZkeU8nWpozX1FgwLdkPt8dTgYFRfvovsMZRL/iOC
gVIgoVXypaIbvBje+FDpgBOUFN1Ji4uDX/89a5WhfiPrax4UPHBR2pszTvm25ZZXbRl/V5+cdKAQ
+40qGjW7SHBEsbHNmlDCvzvs+wnOU8HgMQyAh+YjIJ/kPiIUR2R0VbV7URLmZCyDTXgMBWoyPPsT
vzWiFFwZ/7Q1FaOcH7DGV7pdvwdwBjEo29qlTzYYHLVoSMx7gNqa4gPN51wW9Ur80eQZAnjVJLFT
TRSQc7kZ6DgcSDfhWzEae4mk1kC1d+CV5gLwQPlcse6WZFMVgpsuTk7HDbo16BPX/h1NaTS4AoDX
o6mKAdW5ZcSb1g16SDNxPyB2PRAH1mQaQOoInbnrMBZRJoNa0YAHnAPT8T5EHAzXT9xwNK9zaDVX
V1ftVs4cAzpQ3qCZt4LjR/K/lG92oCWCqIUqNCUZoLmzNIdOTQCEAePyG2CifBt0MLFi/2kMxlCS
FcZdUjlJ2829d+e9CiDiVq6bpLvyF33r6uod3lXhQoY3cRQO3PR5EtDJUgqTh7ctQO+PoFox/Ado
wIHa/BXrAEUdAgVZnvFAzxA8pN9KjJKabmxK2kZIZlCBIkEieDq30BEL65q7wx2vWhuUg17xDJ2q
sF2EfBbWiw268YbN0EDCLL4KTm/7Ic6O1fv46IY4CTC2N9w3iHWoY2hDn1YuGrcAvSljvnwzMV7h
YQDqzpeoG3KW5pEDvBlR9SVH8p3bf2rwAs/8wPJtO/IzCRWrOrXOy8yHLd9Wljs+wPETGWU05Xwi
g2l7psxxCnwHD92GZeMuXhlZoyVxU18m3835lTddG60oF4uwMEWlNUmui7whRJEzNtMic0eBr3fI
j4bOrdQZ+M4dLVzbZZi0wG6Nbvp4QAfMmJWDMvTNBZtJVurM9exszW0d8kramS1D2vC2l3+0mxkP
L3q2777QWu+v4jDXIXkENz0Q2gHXadM2HKW/csvY5j1I79Oxs1eTz+8sVdsbA/aG6EkNjr/fS/x4
ZZwVhMcgInjwhjdpvrkvT91AB+tNfm/3Ks07PuAAR4EUc45jynOiCIEdNQ4jyFpdhhTxmyKkwnMA
/Z3BawqVX5P+zpZDhZ/U9S0anU1nLSMBougs3prqEV1sLjnpsNJFKwiJuaD+2hVr8RNEl2yk1Hxm
/bGdfhu0lnpHAXsZhshkeifZO1MAfS8KeDSE+bQ9XkVMj/y4rLHeZrN3z+dZkVHeAkz0ael/gnm2
pwqByRADurhqp4Ia+9XcemN/vUPWOBYWfkXulF+9m84DkmDNPk0UmN3+rkWkfgxDxsKzAeINsT6u
PI7gymQRjZLVWp8FtkXmn2X3cEj1+QzFu0b7IAGtkBn6GUygaDNs4zjTmAfcplvEakYqwnRZu2M0
8ThU3S5XSKLVYMnAjvwVqYmdX7cY6ga9Laq4Ghn9YJnt33wMepqbAlegEJhOHU5OTAzlRO4HQWqz
9JMvoVHlgViyvtDzq7sAF1yuOZVft/Q/8AnnhALUppxJ9QfP3Gqwbqaw3dCDpH9ZaYMknGxR8/MW
8tHe75Y0QkqHwqzuTi1WxEyGSXwweHk7tgIV4yTnbzwhXB2fh+J0Du8/228Z6jRVm+130ayLODZg
lo8w1jXDsAW0Um5n3TGkkjrjAmwmy9LyDyV7BogKitIawPa9P90y04uTsAM9aNzzAWguMWUZvBaO
zdOQG7F3+5vrUOGvManR00hSPAMTIWnCOEH6wA7Q/2psBWVWKBMlYj34tH6nuUMVMRrayrVpWQHT
+zbpzErhiE1rpdPH57llHeMRKpP8CWME/VPVRpzOOHIb3rjaOd1K+Gs0m8WJ7yO+1w2P4jSYax60
a5XScAh1mYLOnE4M4cdhN/e/yYRpt20eIF1OpK55pED23VMSMTCM6ic+9C2opnbE21CtkII/04PS
zWEAjYnHwWRrVu2jNsaF+SaLSKyVntZ226T0X73Loo2NSQ68Rn3VVtL75XA559fjnxd7AG1v5/o5
+QQIuh3yFZS9QKA0tANG6BTvgBiw1np6Gx1t/JRrGBPmHJQoS5VBwsCTwlq6F1kGJGlCcJHsDaVJ
1tUHNrFSJzLj4RRCJPiG+QzFwLydJJtDmM0hQhVQnveobuCtbjlBBI1NICNxbpIk+0nVzyO8rjIu
qhKlj+Q3tJ1xk33VMbjcKQjcdp/TjCwixd0D/5dce1uMeSvsiIfYe0MZ6H1bgx60pXqza/W3N5IW
S4dvhgq9T+9bGanVcvkCYKS3r0ae7O15VbU8+uvWTxZrpQ5s9Uk/EQ3X2OPtITxwuvmkHnVfzilr
4m9QpfPzHf4svquf60wnNC/9mctxq7LKDMdeTNUvnLSoQq1bTeT4kRoBT/vQumQd8nQHoFXr7Bx8
yd+iL35/BmS07Wr145wc41YAyidG1GXXIaHtYAIIV3L1il+GxkSloQJgMTCJTiH64N5Mr2mIShOo
GcB5VCRS8jcA7r1RJT36FliSV7PgOvzqyHKUYgH8BNDkYXyQTl2rfhN4QUgbfRNqrcZFGXQTjTey
ISMmGqNSgcspEAnvDCdqsAPdEfqFBfUNx2a6SzvYzuKmZsfShWvE2VNlnGaujkWTF8SCWHFnJ86k
6vviqdOKp7Kljo0hILtmrCjp8dabbxHKG+4sLleYHU3yMq0S/2Evi/Jm6YsVgxwCkUZxXMp024r+
P3pSoVX6R8q5PArgIPzIJemHodFXAFZebryneGmU6pVeYR92kvpn805ebIVqt0IHcjR6v6OKs+kq
bD7ZhPXel4fGXv3XlZxW+YVdQbrYc1zyrX6g5/sKnhAwa+DkEjgOfd912EeOEHylwjDxFMRcL6wv
c7lVFMqJ8a3pi7tjC6vZgtdl2dVF3PsuKo3eFSHprnR1NzclIxj567mSQirYXfoAFGDbhgysU7rd
69hxKk1WTvhnLl4IHdJ+yoVjTwkYDuQoE2KTw0/Po7JkbHZ3QYHLcaB4bTXWd2TJjmBU/te3rO9a
jjPJyfUdAdDrcX27T7vDx1H8cpM339GLRUrDy3Fp51GFInqDN4QW4FFOimbj2+XYhjAlR9LI47EU
7k3QWZcDGE9Cb1VvEwSH0RKUiaqQHNOQLTGYfBQLXrueRbqzCYqAVtp8fsna0Nn7mrgvAXCdTJ3J
E13jORoI5wajHLJi6JybN0NZrD+yBIm5vR8+uk+yNxoSwt94K/sO8E7fqeAFTR7eHUmR3daG26+o
ov7P/ZPd60ztmQYMzuOvtmIlT7Uzi1MP6+l382cS/nveNJnINHFO6dFJxCyRI4wPqymELU8X38Uj
jIYYmrKkbmFSuMsHwC/tnxV6+1yHef2MHtwBfXd78+xz95TDAjwc2WXRxwmABzOAcefY36dyBX8e
kInw+xjXvd3MGuAyHDgqvS89UTntmpGXwK2Cn6TaRbZ8Yowp9Ie3umWYUdkJ7wg22LMiCJtYTXMp
7mFFjTNIQnajMB0l0MgSlhiRsdLZ4SkmukHiYzHIqWlq9+0pj/84/At7Zfc81FI9WdUeWN0EeXV9
ro3o+q5ruPa0x7jl21dwnrs47Zs8tvlUXVzwDPxFefim+0h9tY3RoutNrIO9ml9blmHiI20dXyFe
M5QreuD1Avgbbyw7g0tE1F+13uJCOyOwB9abN9dF4kWEqagSISQ0KMaySNMAma0UrBSlj6F2lHy8
a2aQPC2dY6cDHaWvOfVGWS3SwulBNoBupX/rCyUueca18YxyLND9jJG2GoQphf1ea7g2pxk14wvt
b4bre62Q9bgHPg8D3sKvzp6CFeAeydhD991VfPzHYRfpII43Y56jLFkYrYsEEXu/m60atFm+vLO0
gZdBfidPbcNVE/+m92Qkln2oYYaQhKaoj8gj3+tBc7QfHy9HoWt9e3dZ8B1uSPyeL3kSWVzrELJl
l+3n6noJNhX8S5PSG4rzOFfDBvUEifuc6S6kYiZJCbq0BdDKMcSvg+kxhbpbltmC0/evpXgkABWq
zuwo8Fwun9zRZQW6M1bkDzXsjVrcleeD1YbDGB/MrAi50X+0jEzPzoat7Ajx/Z4XOwC/WnlpJLob
2KWPjL2XCGhQRpIWUoJBgbRDpC87SwBSbtSwgGjrwxtVb/c8Cn3ArUAbk1Cp3V2gs9DR2oMaJuE+
q0Npn5tOrDOvWMGSq1TLubjwtmc7WGx0MJGkFwiiRf7hNv33jX9qA/RsWPPQNJ0Uqe8Fnh2N8NsB
0b0T9yCqQKA88vpIO2RoTGiSmBybEFksUVexrQl0ApaMpgkn0nWjuZrDo+brdauNW7OkDPti3gAh
ePioovuBToJTIE92ffcKA/GCxz0xEyVMfD/ex4Q2k4DtowDhYO2JUTvvtoMOVEG9GAam3Qz5QXKu
2XGUzB+0X5bGhSdohOafQFop2G8y24/Zq3fUnNTWETiE+ImE8HvFfpI2ZHVWj1TGjS3iAlyOTc13
FjSPH5g6AuRAwoySxbW1+gYzfbPdWdzUbQVyM3JrbYaN5FnnbfMN2JCYQK9juBB8B97zsw6RUy3f
F/jVgsbw8aByZcQc33+VNc2wbQQbBq9Gl1Ti0EU/uoOLjLmDkdiaOg9p8FoULOu8a25k9jDJjV2K
0+eCRtx/mE8Wec7PyJ5FMY5tkZ+7ZIizZ6UbEflNx8GLp9kKWUzcPuTpla1jFUolfaSafuDmBPcJ
vQ7Qfd9NoJMjlkOGwf3Cu7ZUivAQxE6V4MN0Yek9o9a9dgDBDYsMovS6I856UDg0FpUOY3zGmTv2
E+I0dmUhOrBMb9/ggZ9Rq8w/75bDln2guROL92PiLnv1n1mn5oNB+mMndMzoVWPKD5HvgPxXYFI3
ZPb7NazGT/C7sgQs0/HV4Nmuby1d8RoLKpVVvwXe0zw1XHxdL9ei/7ZTdfeMUH7505/PEzr4LqCn
IwNj5xDmcJygLSWW2rUY2XioB24u/bRNE54v+afYmJ73ZlcC/z7VikXl09lLqTEaNv02RKsuigrI
3zxD5Fo765OusUzORJVWH55v1tyR6oTL30Kk2eoBgc36fH52aAULGFJR0aZkokT7pzHx6PvA47z9
t1H7ApOB2ygea/pQSnSB9cNnCoU8raD6e4pObKu0tVZsUrfEmlLrvT9COCKyiMkX0zQQjEYQ3FDx
txkb0GoDRfpan1lpS07uKSi7rimbeVhFpnQm11H6S+mpIRQhJQi1clf66jHyc4gIrUbzi37/IPxg
x6nNy+b0928Aq1tgBmYHqtoEG89SCEXNEZgvHHaShbsSaWzKnenV6GP732ae5GGYOLB/TI0DTM4L
H5lvCUeHJO/ljejjMg7rIfB6eA18llN7WPsDeRjaTcuXaSxYHvJut3uCZnKVgC0TdNhQ7E31YiyO
a/XTuhTZtZx2yJT757nhA8F7xr2HUs/dw+rm7tFT8D6ldF5EZ1+Ir6exsanP5apWs0S1dtkqmJ0C
KaKYuan7glMylYN20DP7FnFt5tjFkFzGzB+YDwsdRwYJ8CgoH5OtlA2IFAMQj1c93Z1dFIOdGE+O
r2TC58YpdUO1ZBqtHKbnpH09uAp5KzKkhYEzKjkvSoq/+JSo39XslXqlpgRpl0rX00/W0/b/MDo8
A/jnQjn/IOwgn2YSBP+yAwYU/UwPFr+bgDJ0vXgHb0J0LiO0CQ+jm94AZqFiiZgSMUOWe5EoGOIt
YwS78oX0Yymhpz8JqbQiEuCH3DF+hIyl+PhNwRZCL7h50OAw8acTZe6eq0+DPboZJstfHsmRFGR/
q0UYBrgmEUZdjMrKfo6gmt4dcR0kjNWiuUh7iZhMqDSTXxN1dQxbzLU0GCSGyqc5nl+yXUv1oPay
t4TC+jNXbk2WvgaaJ+0I6a3YpfAQG2QxKxNFSoBv7NoDWBfng7x4PU9xyZWEgxWWBXMlNDWz4Rcf
cPHnFKedUCY+HU3ycy0pRsMj0QrpKhRXTIm/6ZylcM/InRb/DDMSZKjh7PJ9CNgEPm03+G2cmUn3
IBhFpiX0wxJIKgKV7YX2vT03jpIPzuhapjtwP/QvjZrh3T4uPIEeM2mmefkKuB0t33VR9BAg9z38
wOmuTYWCJ/8gRyYD7IDVbENI0ccKNaELHZYeyvXrYAVKICqQf/J76Y5n3dMu4f5eHQUqsCnjIWJS
5DUgXkzpv8SgTVWHvxYF6M+a1/d3RkqGrDtK++BMJMY73MLOvswjbd+0hiaU+YHKm9cxf0L26d21
F7dRBWrA3bRsguE/kssf0HhYPYj28cytu+hl6C3g+r9BiRaTXbMae4ZQ6+px6LE1yfwv078hasbh
+AX9DS6DRPbhujtTLeyK57+MaHz3Gf6BcEfyfd8+QvxnrGVJYUoG94iXHP1Lh/i8b/GmY0eCJlBB
9qdb7d+DU/naEQKv2TgYuZ6CFZYMTb6Cb1OFTlEm8BGRt6SVLNG29urTOX/bzmp2AVkeUQYXHzNd
65njlGXJtEZLeusFCHrZM3xlyy5A/PVwTkc9bfVHh1hUAnCvggZ8G/9+jY8j39XjWctQEMzY2P/c
mqHhEbrO5cpWjfr3SVcMzarhBFNmMUCEnDcqzM5dF89KkuKkSIaED1tmeYhWa5GnWsCvPW96AasR
llIA1/3BKrr7OzGHsjs4g7vUWIIvdGU8R7mupj+5Vjt3v/G0opDuKijkBMHav0xn4AH9QwaGRQJ7
0jKb/5IGclCbO+t+Cn5RNVwD4OvSlRc4FJ9Cfa/efXp+y05JZCvtGHYOJcUh5g139rOhB/dkKg0m
04A0t5vOihJFOxQ2+B/j+/oKqjqN2CYe1NEU+5o7QEmEsQPrgsjp8NUiSJt65kUXcTlqyW/lXs1j
fInOccaRmhJcdlwxnHklGdR2gKBxrcV6dQj8t8aT2vlChl3FdNUByYVZHlfCMjdX6MiblMbTHUBN
BaF33zPz4LnhXSN1u0IcHLCXF7B8wHxJ4aa4FEGygHYrxTlkaZwV9QwiqivgdXBhoDYe0J89aPgn
3W0VEXNd+DaS2cPZcW0qXOOuzzj4wfJd0v/Gjz+giubYJUoaSFSd+RiHwvqqq06Q5ZOZvYYJOtmm
Gt0e/SYMVCR45dtu1RJqS5D+xsghmDc4RHIR4yW+EkfyMLyx1QCOUp1z19i+NGfLVZxj2xbYomcs
PqjPGz2nnZrPoMFj0uJKDFiZqxfn44w2w++Sl0w65WAgP26R33dzJozSpQ2Upx59t/jBUOCtu7Hr
QtZ0211k9QJ7HICxSIqPkn/mgCy9SP/XuuR4/9uWm9Y0lnUp4Ez9u+wkR8kO8bQHD8lQh7Z6IuUp
5QwozbUg0p/SooIomaopiKo+bJV6st2BNo2Q5hTrJ98mI/9s/V/vlwKVBU7tOdWpecvUhi+yrXxS
HkK4E1XaaEioOmE+713LxE4sTSN5E/6nNFSt+tFs1+dJaKjx68ka7EC5bqQG6NPIUwPqe5cJShKd
7gjPixGH62FAUQPOUx6g7pN80zeHp+LrXJkIee14/5PxoVqYr4WPv7mk77xL9xOY72suHXkRin4o
N/I75Lq6r81pPgDbUOQllVLBwQ/7EQAPhhQpDjG2Xfac0zzLwtvxLrYPeoe/g09rAu1qVgVesIhk
N8ev4B9L/jWtkAMi/Ipr0elrlovN+tjv+mZ1W6bFtrypRU2z6uK5hqVGMf9caJDuAvB0eLZi/kEi
4Tp1ha3yQmjWon7oGX4ch/OUdQ9OAg6vBjI/b/0CxWrOhZLSbsXXGlvhKxRTOUMEh9Q1e4Qb+gqZ
3Qj8or6uywnr35u9QuYIeIPx5tVQICVDuAesWMDinYNguWvXpARZmiT9Cf3awqg+NHrPm8SV3Ijy
MLqhJ1Mj6zwFOMQOKlng10BWX4tZuXLjEJ0a7iYwNHqxX+ZHDOU7HNzrHGPGzvVI72FFCPl2uQNM
1Mp+LTiDquY4kGAnCWAmLO8njdfkh5OFgRBasR8QpQvI6a26r9QJ7kubHs8iCH5m3v5qksG3Om4b
T2RS/jxQp8HdzaZKLJnSEq/h6Y8zdfDjnYKoENXpJpjpeNAAmGDSj5d8MQ+922O5bi0UDTq5josq
6EuxRUuQNTu4Kcs2mk6j1FXSUSIh5lYnJBoY0SZGgq8VOkOE70QBCWWYXYhUEGWAPyoXcRHttlgc
hZL9rDK2a6y6mcN/FrZyxOyeJD7O++qM6mpqYW8TlhGqKBvuIZMTNUgpBPXJXs6SJpbDsgjjVuTa
qYxGHhoZ4xErfE8vohZffhZLWC4SPBxR+J4Ny/yC8//NHg9DH87bEm+N2KbX43kcp/FvxR0cj0Xb
CatHZ/IKezy3ik9wH/g6PitdqaXst5wOBefgTW+VsGxsxtdg1U4QrcDHIeM+VRTOXkFfzTyxepcS
W/b3YuWx6sLxpJlYAkn8g/ekzx9LidIeoJAXi27BI7YLq0FU7cwZ7QVDCPJVkE0zUH47CHm23Jvi
BvHaT7NXPIf/Y1tyRJRwD0SkalBi78RQkOqIS5VHLOMaPMUJGKDa3en7/Ek5Yannsgk3HoVHTM3u
mn4i19WIfpR5vOb1X3sUL/Ml3gzauwnQ8q5ulzNnyUccjv9sHZPtIvLvmJyMtUU1Sc8rmnQpsN0W
ER7LHup3hyJWCqmBgSc4aG2zNff0zl+N3BtjrnRD0aDqao3U/HPSgonjLY1JIgwkrfgTLjAK2ZhN
wmm/wRISbkcLpuH34lIpx1TxKvXMHVkI2N49O3OAgmf9e7jZVWAXNWNVb13Kmhz9zOmoh5uaCbpX
529L4fTNIFUaq2L/X4k0HLXgMOJ1bNFcgENvPrx5FBjRdHoeVliYeeTaT4ok6DIYzxg5r+zccKCA
SyFo2pKrFZWnnG3eImsUW+Bp6e7V1TUBE/inaMO5oioI4E6hTPt/tEbQ9kAZFN2/MaNMkoJbx7fv
VtNLRLbmMGQngnABcbVCZ5jQhB0+V1hKBWVWO9tkf9Aw6CIZKJTyS6xPBWr2oEknFBtvYXschZL6
+K9wwVTpts8bkfGv22JeiPaNgRNEikNx6T0nVl3AH0Ut2nyiwclDiOp58HXL7fipy2LFZc0NEBYK
GgAe0dt/HiH9FCVJFkK3XxVNRLQdC/LTDUZaY06RJx7d/B+WebHxublQWtYS3EyRhGkt41cF1wn3
nGHkzNFO6ytqL94CiW/K8twOWwzgRGjK+jjXexziRveMdgSTRdqn7zT3ss/KpFQjD7s1ZcF4g5CN
HsRyCz6AKvYd35RU50af8vMgqHll8b/ZY7cGYWoW9/x7/joJOc0YW3soxgHOrLSdC2dTEUMqVSDv
L6ph6NSyK9DRZaLY3dpFHDHcduHU7/2pt0sbvxw/qgPWb0QmSnF7d9f5FUne6kGK4eM2NVbPT0Rc
I09VM2NQXKe+NOpvOgo8Fh199j23Cmar3fbCElAAE8epcRucnu2gmO15v2XNfM820q8445G5wV4l
fLz9VlFuE4dMLbp3jcOpUC5XCqJjqkmmLlNB5RK2ZWo7ruopWEPwqQWnnZ/MC9Cv+q5FQrXCrmHJ
cwTisganvepcMULd4rP5mHj1HCkt0VnthkuaVXBMwLQiWxiGc0WIzxpbkB6hIvl96VMRVlDIVE9M
7AJUykE3Fxyy0R9VmfsMpi96RTxbVLcSAghNfi7jNj47Tyj3jF5puNzxiosRMKqxoZ+4T7IHgEMm
Txnz9LqMesFgnAzr6BklSRiMOgl0LmY18C4ED41HeV5iP5Yl7RqMTx9DFWc9o+yhzg1vAwVaYvGN
TnoiKawiyDw2bs2EjWxIxQ0x56z5UzABSs/8wsFKsGTbvp3npiblN9TQrse24Qxfz1s3bKcPqC3L
k7zn5uPjl9DYah2XBqBFDA8FgD4Bq3qLxYVhc5KFXBchG64r3uq74Hb7nKbrG2HupA4gQIrzpf8q
I/3nMTjQ0vHJaaWRYOl/HfEQFoOXAxVXy984NGjSdkd6Cq/t9gCfgrEWsb2IsRbMW+dNsZlC5yGF
7ljjbOD3WsVjNCJAhgMRMLQL+jXdWZGSdMRVGmwz5FdIpny2xGBrt6RGWa4rE5/4Vqkp1uUGuRlX
MDRtH5LpuW+ETDcHMv3LDDJZqTGRdphtcM2mS1q6E6yZmRWCiLpFGVBsF6Y3Or1S5fZlIHFCebJP
RUlnZDWW/jj8Cxzukq+6T2GiKgfEp+v84fflP9c8wPhanzHL4JZonueDofLMGX6xcS0ubDymV+Qm
wYbyo/mye0NpQdvM4cxLWv57cV32A0Zmc+FE7eKbilqXnHQtJS4sCAE8Bg/jh6tN+rp3ClzmF5kd
3VNBCGoZ42vM6WKXU2zzaX3LmcpybY2dSbzns8DNjDvFa7jH8kILWLAll2il0LaAoP5Thj4aR/zA
61kHwpWL3oOfaW2jmuIODY0JizZWJEqneRZAICk/2gAQ34FYAUmC1dxXYDw+feMdf6FTKp/fnSct
2F6/05qH8qs7KWu5aYCX0nDBlX3mYkLYhTbzHAi/g6+V03dKTj/AtakCBItgvsODG3m9T5O/kK6g
zC0LX5wR9FafwB11lP7mGS3qBulYZz/3ML6+xRbhh/+0wLP1b5hI52NmCloFNpVJclLjXCCogROa
TgtKzd4P6R41gyqgxlspj30p4zwU+ui4zIVEp5i6bXCuEdWN4VsC5rhRiSTNrw8wwf9QyOguOROA
FlYoKD7+conPY7x9qs028hg1K/DxC6lExJZkXptkzt9S6tB4EFDx6NDMoWGV4odqzYHM4vyDJ5P2
aXmDda0Klfb1j/UsB9XAZ6dC9UsrfAF+x5HeIog97oK41dSpsrq3DQYrurpyDFEvybSnIMB1ip5A
iw5ZQ21uKH04bojcpbXKMqAXtnVnYYzSTFQmUl8gQQZhCo/Glnctr8RHOcmDgsKHU5g9J0E6asPF
lcgl/GIYhKu3eqWuLfIK2MIucGaLiF7sfJnEnAebkaAVs23ewWbsjkvlvtTjMHHvfYVwxiJhUIjR
IJWeMlXXMJv0NgF7U9H7GN0mKX5HpZCcUhXSxRwWZpF/J1s7JxXeIcnhtKxaf4sBeQVV3H+45KDe
KLqyUfljTQo7apprB/0hpHdiSCIwGqY2GqOMxWXXFDMLQRmzbKUNjwG7+JaZTEzEJBE83k1f6cUl
fNtBbEBBphfTNE12q+bTUGpl70rULjxjsa1uF9j5x/ARxW5ge50wQQg1PI/x/SP+IxV5sybFU5Tn
5K1+TGnecrpsUExZ1Qe2i3LsymMym6WkvrNAOLeq24pvdJ3nruAwEZFbOf8SgueX0G07R8eQOvT4
32t76aPGhvLZ/xz5kwo0II4XJ/ehuZMBqZQEKfC/B7BekIyPW7RmZV8XF7nk9oKgbDcZSvajR6+1
98DlzZNGM4tYCdUzI4k9evzCqjtFfYXJDKulprRrUPb61C0HqB4ozmEFDr2moOIipKf4rPaqJChb
QaDtcGvmM8zBLbfuhRoQSjw6CdnsS4UFE2wqxW8O5POIGbCuGiwIT1UDysO1oz1rvSyrH2UgmcVs
VAXw1gjLXBnMoLWTGdFVb7ojVQNLxkjQUBj+AMnIAl4GmwiwcaT31mJAs2hmHNGU58ajdUBDxEwd
K+Frrjn4+k63ixbzMV0g29nxGDKQZ0exa6kjzQxEa+0Q0ww0w/oSw0JDnV1R8HxId1KlAajtN7/O
nPUtHMTpg7h6c+C09XliqW8FqaVlhcnNZjgp6H2UoHlx0fQ1V0z1zZNs2OLjEKCEUq+xSNyDPuoJ
g8B3DAawSiiGpgHW8UlzOOuwWKW5Hin3Rex5PwRAjFWvAjJruW4qc61ywJuXwZiQZsXIpZIrdFi+
CmxTk0DaLQOqCC+8l9hhwZW9saEyINcKYAw8X7Q5MXaL9tE+k4f1c1aIf3cRfJ5rkuwo3yPCuwqT
l0bS8UVJMjRDB2nh/Jz1XrzzQUP9qF1WLAtDzsCgyO5qDKQhRdn+LTCBWAQDjvFJWZqJt1IzlrnS
9qkA2lUuGucLORAk1lJxIXqf+6SYNCdgfdnLUAofM4R4+PF905BDcPS5RGc4CSog4G9TqQghfLuY
hpb1+U/PYyPGxU7k+wqbbqj6JtiZY1r6po494tEXSqPxEgYFDDwv1LP96X9LxOshn3GFTiU3Qztq
qV9iPklPkx7vl57o2f4nfcmkGyu+1XDgSjvlGyI1wUgAQgiwr/Ev7OS22Jk6kyj4SZAhn1fmvGbv
0EMpY95bzSEowEuX3WemQ6aHoVtRrlOO0nnNyU6dauftxkMNzmz1w5B9DrJBN/Rdf7sGARNrNTfg
5DWQnD+D/c2M8v8sLufW5keldJ4L+AToB48BrBijiBfTSmb5b5S9IOvUbl9ZI2tcjRs1UA1Hgxzg
d4Sc9jNRQQot6UMPVnx7R5jaFIWwXYTM0bb4dQBLUJMvGJD116Mo5CLq7+tGZGwJJ6Wiss9IoIZS
vrfds9IZYjqwl852ikSU6IAfe9jXP3oJd8T0MGJovpWlblYvpQP2odsgGStoxYfqh81iygc2PhmT
rOS53oMsl0SwhwkTNm+Qw42qmVlgAtnCPHHXghpxzXCsWkCz3hDR5vbdWQzWvv46gtyt4BwjndAo
7nAU6YnOLNF/Vwg5CaWDmsnPlyuLoDLLv5SfVWs2eCkYAC5Ivt8fA3G3vnpZKi3jJ0mi0Qm0BvkX
ztzTpKFdxM5cytFQCdfZrHziY0pCeBcrDgeU7NVPX4avm2xhuZJzQpnlKykSJwr213fiZs5psyvD
1C6q6RElFoLOMU28QHVImihUEzioEZdBXaCA5Sf0FMHxjhawI2FunW5F8kOL1dnylyvY1Xd2mN4F
MmsasOvM9MQs1iLCPlX+lyimXLoqCnBMVSY7GjvbLTdezuRNESiM+EhppPta8lXQ9E6Yrv9yf6sJ
1ead00AY/1YtQKW+ZrUxwDruAWbG8FeG3HnfozScUqVHV+byp+/V7JutxmFsqFDGAzrgJspYp+Fx
YYSQYYYzPzBxK04ThWXUaeq6mbYDERq9IgjmSpOW6UlT9CyDOpeihm+8FcQsrOjXLfvN6kHkkXta
EjOCMlZSU+OcCVzf/W7xs4934mnqPa8Yuo/WbbEf0RVyNMRxrjYbPHxt+Jlnr0QEfkM8yLPvWqtf
nXM4CXr5IkJwKgp6IJCgQkEp5nmpf4E7Kg0IL+5/zk0XIwNMdxEjLetiFae/WAdXxnrnTllp7Lhs
7KYiDdi8KavrYd+lwJFN6erCQpTkVXVDu++YnKhObx2kkDWFF48clCPLE5DA4aF4+O7H9ydhxbFo
UnI9YUZLybdMBXN3qgN6iVcwksjObQqWE/T2bcocKkkp2bP5Jh6CZB2KqnCbiFbhHlTaHtrRFoQh
u2qD3Xc5FPH9bvz0b6F5qf1r+wKFgUWYtnHtnRX+BbwnVsSaQuex4USIU1kOiSvRF/5DqQOilfaN
0yMgJfffzjycJ0DZkw1lvypDBNcvd+5Sqq+IT67ob9cjcMlKjCUvUOJM6obSMLw9ycQ4ixQH5d2v
Z3UFJY3tTwk0n2oFqWckuFpEXdMUx9TpiV8H42tILPVIV1i6u+aWF8RjunoC94Z+VPkaICWClqL8
cdGXSlBa9ABRyJFE9JyzsUCPKRtg90AzWTEnbHcQBUHfhykRaYzkk4vwrtDnxh5J5CW/UiESj4R/
9eYYoZzTpd5HKNPnjU5tyUKsIYzRcnWGWBeX3O+ee4O49iSwNiOpBrQf0ZG0VUS2EFAd7iLKQLiK
qugSV2F4fDOdzz20HcB5t3SluaJJY9Q7PhJkAR7PuLnAIBrJQOVimZ3u2XiVI47fQ7CzCISGZySa
RZURy14dC5PawMuubow55+HxzIZEBtyy5TMpcOP9FGsZHleaqQbK51h1aIkh2oOLRGYjLy/aD6aL
Z/53vHEgjZXJn/LNRPc9uKYvHtEPOYGLWlGI416Ly2qWAiknqOil6hjSka/NftjmdTX9IkgRtStj
JouF1SPiuXi3O/Qrdn67UQ4nxMeKHot17hmro2xe/sfUdc6Jynplv5t941b2GeTOzfjZesvGNfjy
7GRZAvHfCnQFDnHcohahJGMZ7j4+Q34gVfJoAUy6Kb/NrBPgN6+eMCRKReeuJsQX2nDpN8lgLFmJ
6Fhp0mJFLKzgg4A7m1ddat69bJbi/NarQ2oaz6yK7ksYyWJXJ03GR7M3ZzyJbbbgIveyFK4Ab8oe
1CghvevVFVFtRyIgkVQWMQYqcR+hvi/GFlPbxL6nx0RPzjhzD9tvmqmkGkKuHoJLWIzv0prYM2Fl
Ld5+YW59FmO49tSf8WPAEBpaIN3PO0ej5vQ7LCbTqAN9peSR7ZhJiFbYiL5/PLoVW7FRwdSBQLEL
dxMvD0vmSB65iN196vAG00Ie2uTDpnMQHXC1onPgjspKHTHUUB/UdrT4TUGz/k7V+Nhi5NVOo9iM
005/O36dpu6mpndVKXRhH9huIMiZ9hOCtFsMwVQIIGYrN1OOw6+ja9jtEmw7mJMm4QrIdCjYEcnC
Panhva1vmHPg++pp1UMAlVrgs6KzPMgNyxcVmSQWULMMWJJHLgL7EwqchKSQJrI0YqP+DQxWwqwN
Wv5yvExNfbD7TGymeQNxJnisCsAmTmSJwtyOpePMf1rAYoMZX3PpjLZ+HObn17UiOB5GnG2+s7cd
pwQzvA/AOpQQkg2V6lx7pJbA9Y8LbVM7yOzh82aNg3t05J+dJVvyFfhcDfrs8YkSNYvwt//Ni+cP
q/Fbap25yZK0I2NidejHhSOhtaNzCPq6APcdhOen7hlEkW+TJTxnRRGR+czvL2jmwEu2UuejX0Fa
vmSlt6cwfJ0FY7TrU5Eb0zoHE2vJ/LJMQ5cYFH2u0YPlhnTvB8RCabzzM4qowhu9bcP3JOmpnwqX
pXRx8P4Y3oC7lSxMdvYW4S1xRtt5rJ9ih//DFWL7ZdmHtuHgWGtAJfeNIbwccKvMTy2gPccNHPao
6X+v4PbGUYnFhDtjk2OwM/tt9Jiue9KfdcShoxiTDNXE4mreh6bnNahj5n1/bxuAYMaNhdwtLyvB
kGq/lZMSHR1Igwm4jKYR8HEvy9yT66xMiILf5iqvUHSmin1WvBLfNi6HgesMldDWAB5KF3KAYNVb
48lmni/f1rhuYvO+n1PMov8iVzNVreoQXJWnCQo3txgtgpQOE9M+fBgrwwDppzfhMdgAPo7HUX4v
NTAK+5Z+Trv6fdmoZeGulX4iALGLMsVRhMA57qyY3lh1BI8wD7R71kQRLqRx+o4kdKN+qFiS40s5
fbxMlw6oSTjWytKboddSWhVCq8YamA2byujQ7Bi8J7Qia9DsjYv6d/UeeFSVhVdfgx5pV6LQGEFJ
Tge8yUa1toTHI+2C1EAXvIUepFlLtNQPR9st5mPgfpy1VbNMMf/kczTXjtDyzh90jl8rxE48atqr
vI234+uwKVo3C90Ce2JBO5hzET4zZbSkzu/ZwgyfgoJlXvKNGjCBOmlr591BcbTOeroeIdJ/C2hV
fUL+ot4mM1HEsaGvbeN6GmJvC9jv614nkURJidoIIFAWk2nulQsAFJ6oynf7u/PnDxM6pxV8kciP
rGkRDa7ljdM5dLK47X6tH0h2ibFsEeBU3iZKakqkmj/hIjTAA2tjQjVRpV0rk8r7Y+lesMiwiug7
3lCpHXTEutSQT40XtC9b2rZ10FbuWZQx5+Yv4XTGJFoouLflyJTJshfq+9KW8yBjGn2OlQs7DHOe
ugjezKLUYBJYCOHPCipjLrqJCDwmXs3UxERJ/k/dP4FjJnoHMtV2WbWiYY4nV8QMNw4WlSsrg9Ay
5VmQaFW482j8sFSLm0fYukVGEjHCjwhxicrXoTSNzB2Uwkp1uZUhroR30DQBjvG8btibZCH8cXJ2
jjr4+gSKsEC4gD+Nbxc8QzqNbufcRBe0hpReEVhVlKGRbmyoDE/strVJh0rganpbIMzxRLZJlNKR
zEifO989dCbTnCPS/jccvY2JAqV2sdCZ1ZU6Bu/KPh5OaIAGFF9/A+nzRrUOpd26SvPLFfTxHtIu
kVnPlw2KOGDNDd0INNQD9FcqwincWxCRUh1OwUu6H8PRbZ/evNFfOGKSaquSQlcSf0sMUsSC7n/t
RmdAMl/u4kNInBt1D5ytMbEdqOz7lzaJjwOEIMgMqOX9dp61mCId3KfCNyRtXNpOXqTOjFJEMUE1
8XRLWR+ZOIHuD7VObtj+pXeamcBbEJYAcjHWsX7cCKlJShT4G4jBwAR3fPe09wOrfhvrWNWE/qxR
Ly+EfyaDf84mWdCdQdr+niEh8GpT14BSv0tq4XMR5rRS4zrsVZVe7uEQXiJxgNK4zHp2ymAJN7gT
ZaEqyMfjmEySwSyn0iL5tzyLOKgCQRhlyz7JOb6v2VTZcfFKC0PBCroDHAnJfJxd9P7q+8EsKbgN
8d0ggChpBiHl+ZwP+Y9Ui0uvekJRsPyBDdfp/p3IosB9euzWvRS3g0nojrqmONXaBt5ze4YN/D3h
mwpAk017PqzN40sNr2qJv3Mw40ZWW7D+tPkKKQ57GaZiPZByl9LCZtrUl1tHkyQqYC5jFNP8HP+d
EcpcNC1B758xD/asa07/6qimFUeD7rfmfBv2X7Igk9IoOekHkX+3muY+Zae/7yubup4lPfsr8IGU
TAdN21EGxXsfRhLwbhg43vyqaRAcMTnxUycS/MMouJpbm60IcwrBY+cFORa1QNsjedKkFyxfzMhx
S31kTaWUdfm53AWrxq3elgG6aMYTQIyRfibZPutbqItT4URUuD7DiU1dixE2JGPOiwm4qn5TRCh4
4DCAT2Pe3BPShh5P0v0yjDOcPn8VwIXIoY41a6LQ3mTKt7XODrg0bPoHxBI5dTIAxyjxnjIR9/5A
MahjAskUzw0qkJFSqODYr0YmZ1HnmonQZyKke53qJi5pduf+COj1i1pLjCGtEyl2mFWAUtoonFdt
QE0wecsboF/U9qkVnHVb3+NjKXzvIUnso2FGHLaW9Yzy570+hyMefy6QAu7mwVP5N6ZojUotX7IA
NN/h7b4Z4pQpFX+9jTAvKmLYHSrlyRSbh49SGXwoCXnqlXAjzTt6K9nFimiO5gljLDnoWRN9t5Gb
wPbtDZEitQwEwRiizv4yzS8qRb81XPJyoss2MpvcsRqchg6e2Quh5DUxiJWNg4k+T1WwKKdYYYFE
PQtMJ9dCYgVXosJk4VbeG7jhHzFiFr9+N61weF7Ig3tswhDUz7D2pKZwEkcFrpH4TQydAG+5WXoX
quO0qkcSysRiojvd0VykBBV4uSuJ4vQ/jXKt1CKe+57kM8N5JwoyvnyheEcnRP/5/6FYelWbLuDE
m8CdcQL/UrG9Yb7E8Kp3PHeIGCyw0RJULQI6Vuk8f4wJxGJZAGMjU7fTSwR9Vp0Nfd68n2QxPQ9p
aSzRB/EvO3U8w8ywT+ZJPtsVhfEjl44XPUKKhIbBAQof4xI4tEbLJ6gIKTt0SNkvZvdKMy2yPX9R
m6sLjxTNav9xQjKRey2SJ7D+Bakzy+VLKK1p2nXCeSGykR1aKyKWF0bIhaSBgDH//HHfKCkF++m4
Ncgb4MOl+V10VxN16mt7GSeDFwT6POSB1fEva2yluL2kgo/9gLLdT7WEB3/IWUXq3Sp9ToD0NwjX
JDIKyQLLncpPPcVNpjraw9+T6Xwe4KoV65NsPOSnVuq0a/H6WxajaWugbtjP3+RckGbCnfuUqHFZ
4JtQrlnYO22tz41NbOlxUo0hSNoda+4yM8TRv+SBdI+5HQ8NQ/y5N6LWuJfWeQ/12LnUPzJSB3aU
z8Ek/te2JJO1RzqFyduB4ikJDN3uxA+xhLs5G5Fc0hgQFIcQ/ZBhq71ewzzaHSRuN8pNMBFJMGdC
1cYSPGQtWRbbjqgVwenO2Sx5GvTn3O5LpwK1D/gmQo/OfU3dPmme049232HtLCgodSu2byvcGdnz
wunY7fIs4bSDKZJJVL6qDO5+OC5wu+BYAIE2bk5hylXZnnfS1WqfmWWPKvczudQsI0YtqxZGCoPK
hu2F3YpohD4Nt8u/op/QTsEcZoo0iBGOuHqzCOjMecKN/SwnmW1zlNq9eXW2BCU08UAIM8HdUO8z
yfyO4aX2jXxnL909GC5Bx42gZaiWPfHEP8BtG+LUm6ejwfWraoShtGVPEZLnhjDVFrl9ZvMcqto2
GLqooRyXYK68NsKCfuFh/vOf615Czwo5jUprTqMJjDgbDSXQjxFx63nyyg4MGR21w/6FciFJ7rK6
OJ/Dft4admQizPx4NaSP+pBwRsshDCnYDsx2y4euyOMuCsK3wncl+NECY5GAwJUvN9DC6sLPycqS
RZs3nuhe7a2LC3QrKH20gWxDPCv1AKUU948MLoCoVVnKgJzMtznISRy1erflnLWImldexb27hNZW
7yL/EUDJFcOpg9juMTNzdL6PgyIyiculJfgvMBu3GwqQeu8yTKaPeE1BVnCcrQ75wZUEhpDIW6Lw
qlc5VQkbqWHbMrkNkMup4Mp0FvkNT0U3+2WNKs7OZIyV+ot82SMC92x0reykJVSYRV6XQPCMj7Tq
s0YsGXmhlvuZLegx729wOFVQM1eKGVEXWM3I8F4UzPxp184ePdR3FieiL5bB3bEgT9l7xkYAnJcI
U6hy+GLWx9JUHJbIpL7Dsx2fSWer2FgXKwi2kJ0KtAfFa5o25yKoJSb6+2EIM/MW35WCZk/UPrfu
4gvA+lKOuuOtG0Ba8fdq9PCaQkDTmTm3FRhInYbOf4iyCikNd0qnjeMitqxyUMnNA0oauqnQbw0G
8S+iCmmvL3TxBjtF+652iTjXpn//nlk8jZOhXe21+p4r/AxhgCXeAI39Am8Tk8lHV9T9fYamsoKg
Jpf5MiVrkEpVvW9F3IyoS4TO8Beb2qHgHoKce3MeuarXptEk+WDuUPPHJ3cheGPQRlSPFr+Zm2bx
13Dr9wjBKNurSffVVD3sxbU3NjRqeIAhyHWsNCf/28Ap2ZcksNhpC7iqcB4I/upvj7bdWTayyvMW
T+l5SPbzwdZmB5QVKzFiAIxqEBDfmTG+MkAb4cltpl+q+KOtiFY9/BGCfCglq7URxn8qaJhzx2Fv
iC0CRdTHI7BxKIy5icLgCIQM+phA4ku+CYiZoU9Ht7DmiYrGh8mGA8yFPi4Jtz7Jvl8AuEyAFa9w
ukRO8MP/oY5b5eGIWooZdvBWZQmp05b8BRyRB2r56SFQ6cvuAUZXxxlTOMB6mLdPfnb54S0W881M
g+V3w741ZCmjhv9aecERgV9/8iwE1CUiuJPBVgJ/wOLSjVS0OJwoNw87nPFeQWuuxA4QB2U+A2nh
JJQBhYpAILh4MD8tg8vJpT3EnzGRisOdoRAF3T+1uxa4hhQuhzky3GORoySkSQsHX8u1X+ROT5mw
39y0Z/nJSLQ9y155VE8upZo1Aiun8YXkxvxc6MilC+v846kQWo9M0GAnhRwJSfSdK2vO9m+22zxe
uaADjP71yCnaKjc2iY6NVEUn7HHUAwGqPZvAEpe1lH/hS/G2mbm9YPmRCk/UN4G6PzYnXILB8+k/
C3SirWsocN7fJ7d0KRmYYhdHuKzyva4cdd37UHXhbhGZM51eePsIZFSBiHbVWBzjyvQCx8VumvgX
/m10NUl+Hs6buiHJmNSxgVRkeL6oNgJNy+LMkXIxKCZrQc83OXoGbwqk8QmBajIpG7dC0BE5PcPC
DshB27aTEN2io7Jy3yCFOZK0HjkHisT0pVY67ONbPGopVO9WtzHklIqhJJ6dNRUQtS/WisaCoKiv
/w40A27N+asgOjdyI/rjINWLD7j2Q4bTxHmOhiiNyuo0J0P4EcbTCGS65Hawh/OrAbpkX29FK/2d
3tSPyDOpXdePzpC0NqSfoDPV3Gdcsy080htpTDxdhuPHqPlZmjsqB6RaMYRMMUsHqwiesxVzxzWQ
tJ/WdRoRhsu7P6fD1m8FX0nSan8Nmx41EZPlZc1pH6DnLX8RGqq57/u/o4J3qcO1mxyycoVg/Lpb
BkkU+McNUGH412srNdlKmYML6eNtR/dX0mJdASesuVbdX+QO8qh/Rviek31vb5kGkUvYdLi26Gg4
/N7i272zaOb20Isv/M+sTXxumbMZqgRvd1o70q00zgfoqUoHAOAv7Ho8hx0IIECw4qIfSV1JHpRy
oe9dEmegfPaNgNa8fJcFFk2SC3zQ//pXcgaQHcokkq7heDcHzLZQwnicEqjxgCwQOIiDU8V1sj10
E69TbCT97m+s12Fsd9b6D6VN8/F/v2+ZsGXAlH6q7dIAkyQY7xljYw9UtSIAJ874CMfqpbrvc94E
BDTnHCi5Qvghaa8LTDVypaFLGZccY7JtyFebW3EDGWLTOq1yCbF7PtioXPRDYTFp2qVDqiA3b1U6
r9VdlsZO4upe680/ySbdLcFzxQTioSh6VGcjrhMhPxmpU0/g6/YTHk7uYzLxtg6cxSrsEwfkT85i
UdALivQDCQzVgTv4KKn8bS5mV3zLZeIfg1R7mYW976UxFvWg242n8XZ8X/JgknwkLZXniRV/qF7A
1AnuTvrKpte0neqNlK6duVtly/mZ9fDd8PSdXux12wylf/gk1TujV6T4uyCLWxECWNYUzPNPlEQI
S/smREBpsV9iZ5MeoSFmTgjpZz0amytCHoD6lU+Cvd0xih5keHF4rqw/TCvViBTR/oHEci480FNj
2+ZV+mlxRy9Tf4Dea7oKdThbSccX+e89s1mSGlSW4qhDtiMxyywy8F3svrca+7NYKakqLuXwkOdo
gQigCoLsjtWnY+M92TsGyPskP8YB0xP8/3rKsTorz6ow9uSaHP80GyZGUHUIrYuUeIRhSGSbGzO/
dgsb6S5CJwJAJ+Ag2c1niY8Ibqeb2Tslt6rCiCHFYflMpLpDhIf+X73v7Wmr1KFomQUn3kOyGDXc
FABTJ13lDdVr22Hg1GdKcj0vAu9cUdSs0lYfo89zhYvSJ62G0CvR8xUT8OSgYtIpTnRlrd/NVZVY
LzkqJpnvEKQpzQbOj9t5FBAlzQK37qewsEr6phq5QAMHQh2xtfJfcgy9RGDmHgs9y6+8gEoNDrEj
ZI9xqHi182S9XkPCf8XZtNU+mREw1C2YeiHDLshwoP7pwsCqKzNTogBCzDTCMRgCMWgEvs27GuMu
Tnx6BSDHYwWg2pgHGzkTC1XxNU9FQLq25AvqwC6cSPuL2fydJrDmGQHSbZAi9snrnVbktyshsfPy
1VZRnAs54wHixBCBqh47gojEenyJ+TEuXCUCybYhPFrJHW4BcGquN7BQCwqfyO4Rx6+3ftAwi9Zg
2b+7BneSOrE9fx9rfJPUeC3GTuiy5h4/f6tLWDI5bdqwF099CbinT+cLsLwNjLn1Q2gt2vw61kBd
UR/RErlBXS+ICs/BYRx+W3LdU6ZowQi04xQCM1LDtSloe3Fjn0/IQmx7xSSz4t0JxS9VzzYDcpT+
FRhPXEUUOuUvN1zZLOgDbin1WTx/K4v2qO1xItmpA1ttXHCGIa0e/e596Yu0TFk47eK6NIH1HKRD
aOu/Il5syIiBoqFrnt2eS6g5CUzMgo+tHS8gQ4LKLZYx0zDCUBo8FmxOSaFbZwm4zpOHIK878U1K
/Uj+3s3Xcn6NfoUUWW5uh/vI9K5pU5yHZevCzRBYLYz+wP4lQYxdwRSVlKgyS8Ze6DeF3HSAQFJB
FaIpIqHQV8FEcauvR+1PAenJAXTlsZo9WbYmAlfC00+eUZO1bZdbk5WQ0MAytPh6zkPWIYuTVSCD
Dd6QwIqCcGXaKDZ8xAehsgngMbB+2Q1csxG4A1W8mW1FcxboiG/o3sdK1gMljJ+6E/IpwQsAhV6w
JntoabBjxnxsrVGDBrvhPfBKOagHJ0ZmANjvJJHk8qlAVeTIfpORAypyo8u6OX7Ci3XWGHBm6YNy
p8gnUOT+zonQKb73wZBebA6mhJdrv+QTQyg9GdgxVg6rT04jCs2qcMm7x4jzq75gZSp1MyxpkWmc
ILIcB2Khx3JpOqWWldhGYjqOmegg/gOOoRcfPT/a6K0u1hdwfco4yvWpHfAiPHCTuocWrsRjN59d
k3K5W3vzX3j/oDD9PzTFtmytAYipGPESzV21tjmSUaRKTaUqanmcynXM8Rs1fHP5d3o8QKwsMFCS
M4YOflQV7Cbp6n1lW3EHf9gGru8Yo3axS+maKSrP99QSdEc0LlRQRxhnNjMiIG83+6uDztJiW47s
e4s3LQNCS4xti0jbMGqiemjzAAUlLFGwzj+zYZIqWAIlqCFLUeNm0u0aM59KXLSpGFEPJNGZ6YPe
Z8pngi0TgD7GoZat2iMXLeZrJi85kjk2JGS0BvkngZt8g4HtFAemeSwg0gMRqxYkJ8tA3H13UoW4
qKOz54vkRoeBpyBxPDD0xCpDS06VLmTo3IkHGivKT21wMzGtOakjKPa1FGZ9WuLeTiSmxgZS6S9A
QsNRqBlgHMeXkeyv1YsdiQjWLFzOEVDSRkwzhT6EAVNU0myioyMXc3cdpe/yARQjLtU5yjftzyv5
2c4olPN8McHbFfcFC/gMJKTiimEB2bnHxwniUV4wqgoDXQFLr1aEtxBfmE6mMSNHboOwPGaYOxSW
pAIyGiM4Tn8gNhcvUBwxlwkS2CxQSBD71G2dGGR1r8VSrcL4yfW8PhDlCBe8/5VJPfUNjjE0dvfD
U6YsNBtrevMFr5ZSVzLLpzQCVAsZGZlmsxIml/FWnmdcxeJsLeMfeIEtaQYRV+CFR8X37VB0pSkD
fdbpJAeKBYZGWIURvy6dIiA8l3skAF/3CTVzsAQJlzrEj1ELlbLZBIM4IjVo6nzXj8X8DXiYctF8
cHcFSDKK+J5ukimB5QZtsYpL61QiwdPDscogykwqdh1CYbkD+JHoJjL4i6Ycr3JnrW4r0vf4uFq9
vfO36beoxn7pDlZZ28OshCcMErxLNsA/DPq2SQ8R+4uCcQbMrVpJLJgCJMJgKOG2/JwPca5rBYKF
zjl7KFBv7CysabyRqpk+SE7Okp0cBvaCGbgi7SM5JwT7b+VeYW3ZqYel8GzS217wmk6OwrLuGMGf
Jl+52KrcszqT13nDFQvsiUSBX28CQPLv1tiK8YYvuTYtTPha1pALr+3O1boN1WJ83jI6ScqtthRR
IrjM3tWxNIJMayWXsqCNOJt86chn6z4y51L9BP+1Ohp+uXPmhQ4DA18pupZ9OU55yOR/DwM650Pd
GsnomNUyxDHmY44f6Mpgsy+JhdYi+cqy1BTO2m0q9+WjF1kR+wl74KZjpfEcV5QHtmBAQXGhw/jc
sJWQdVlXIUnuLDf9mfG3cb2mFsCgdepSkjHuFKT6FHSiV9mLOSjzfq1x1Y1XocZQ3uqgcSa9yEAb
SRjItBj+OER7Xy/kQmHWA4ldwBWTlVC94/T4UbfB9YhHOBaqu72WVE2o7A3fRli+OczvD48MPcWu
jxFpT/cMYJlmR3OsOxB4qvMAHrvjDZv/MtEdb7iMzzBP+rpO5UL3BJdZU04K7h8fA264m4z2MOuw
gc0cRzQgJcsEXDc/aD/vDhuhEooSiz/wKK6kp4Mv/rFLAp2vvQLl2KzLNAbhV58OZmUnZQAhWwUg
EmijmywjOnB3ZwLCaTqf0qj+ywE38cItVpE9fmTiMFjx/JrDsLlCWQMuXY3Eywf1hjQdd9TJwf8w
rphBmERmv6ilGG2rZ9ptR1h2kxsIHGIghUxBgsAayxI+t7a9rC+r6KMCikkVOtC1GrnBpP/ta+iG
HH+seExkWYCuzvRmH6j9d24qjqtog+OV5wv8EWFbwuwSt775PO3CqjztICaP9Ek+67wkteWtppW2
riZ6YTh7I+pbQ23sT7ZONn5930VQGt859Sk3z4+BE+1XfIBg6648nNldij8WfpSBeAglom9uttov
4WJrBgeABS7rXF6Tjp+4ib5R5NI4UtKCR/Q6nVqF9NpGH8x7BJzS/4wWtawtD9rWA60VGpvHk7If
wdckFtQRXySJsD/k6LN25yY+YMp2xZLTvaLrLkePdovLxqeq+vIosFms4sYgChVNM0qen15OnU9P
qpNm8aoEsIqwunAcGDMWTLHSyjOQI/78VvHXo5MRTS/vkR6BI7I9zVcQIw52cGpRcKsJ2+QQzMq3
/QHkesgeH07KC1xu3ejI8Oqq/MQ7wcV18b+MRG4l7vrMyh037Fejo+CTmbi/4nq2NoLc5c1CNArT
VcpxzZnOrm4duLbAA7HYiuujP91YB9lQrhblzxhD7jV1mTmXBHvXQrNtzqbQG1pEZaWTdN2P8Wjx
QAft5ALHDf3r8aAtP4OMf5T6I7iEDAhpAOfK7NhNyUB1hYvWN9Em2b4Vyy9y3FHXO/XbR5IRdYK+
1HYYuRtD3wf+PGJaT9zmRwZAdwgieGUSOXyXmAw1naxjC7b0o3ezqyF/soPeO/SYsUQjO7IdStVc
IGTW/kfPlNTdACFRZfmbt5vVNCDmaDBIrR72IO+RG6oMZuP6t9b58oxn83zKOVV5KZSOnhP1w7oA
XC3I1b4Da2fWgqV0UQReBwo955n6SykIN0czgPUTaZzRI7aTw48swpR7oiF4qDopBn01MpeCc7hH
/vqo37EO9a0b4FlWq5e0rG6wMItvOD8/P40t9IqQ2rB9qvz4gEW1Zu7zpkZxjSVyrmzlz3+/AnjU
WvsQAkBO1KnJRe8dco2bQdnjQ5rRoM8s/+K/WzNbKgK6/nr2OPCJ2epMKtaWIT5VI1R9kP/wKjP2
dMmLQtrDn6Neu7MNPH0+Dd0S+jR9M+MaRVAXIQnh1vD85ggv3tkqAvsN7t4+ON3KEwtTXaHDIwTk
+szSWiecLKVr45vRvdQgPzLU+PFnu9qVrJj+TQOfvD5rtzZXzzJB2V/IxPyOalestcev/vuKlKyG
hkQ5Dc22mB928K4pdNUjZ98mMkDXpfCF25epkjaOJpeu1hvyrIMGvKlb9FAqWkM0jlkOhxr4B4+7
OCbwB8aUHmiZbIJvVbiknLuJVCcYz5We9VjPsMaGO7g0nf3zKYOK0vy3itw6iweZu2eycX40r6Ik
R1cmud0qTksqdghY6b9IQ64FniuG6yuXXXGtA5OUPDItCMNZKRN1inHztdGjZja9gNU1iwyhd16D
RnV+TCscXumT0hyuPO/3UUJ5lsN+Hmwo6GdRN6h7yIxQ9rT+3eEgerhHjP86PJU4xPdDBIf+QACQ
mvg+LJFiSQ0NCRGBESrGvJ/41HUlyCEnsIHtss995Oij7uXge1jaK3fNtnyB68b8ROAZ5sD5qXXU
DL9j7HY16HAiWf6mwsWb+4K6IxYMtdQlsGV8P7dk0o68sONZex4Ukw/Gsvz6ouDMVf5PZ/pVa2jv
3qrvuRQvJ2NiUYClSQ5PLkdx98eCjipDwJK05AhRidQaShcQJHqSFJgLmS0AQc3VaI+vNhMKGmSj
VinHI+zUh7U7dJUkSohdfJYuveS0g91fWshYblAOYDZb8Uy78+yzPV7urkMAY6Inc7HPeCQGelr8
O5lGvFBl4rfUFqg3xMlQay8/joakTEFK+p6KK4HfyigMODAijwU9eWconmDUtGnvArKoufJ2dVuG
ognAkCn/mJrsPUx/2NG0+3VoOzsq7giY1fAd+uWIeU+SIfQdl2+38B4aB/IXTkLn26rvfIBP2ge4
EQBVUaatQVFGHIR5+rfAfMRPNn7yLayCXTgh0ndiWkO1RLPikH0hMtfhfbSKlIXG7Fha9SxFc2M3
AfHHnh56OYrHHTH5ZJj/EzUyUKfTI3GRIq5sy6agAQB1TsnlJummEP6MqM1tb5V6VGZOka3iXbfA
7F642GzDJKgs3z9Zj7QZ+/57Q+19nrhrwPbX77TYhLc48FzNSF1pGNkQvaXk7EHh1Ep7MrP3sPn6
Ha7O5YUU5/giSqFuHj2v00ZfIhsVwAI4aw2WDBBgL2chHchP7fPHIFKVRzayrHysKGkXVBitkUq0
ulWNrSkKLdJjki3kX1+zB8e7BhzfZnQOhM2Fw8MkBiFBBqTwyUis9GqHEkGPAd9uPJqTFjxaZLuO
YXFAgqtxNrBioEMbM+QUQaQamgkyuY4c308Jm/cz3uU8qjxTqV3/28TK7ZE6Dwz9CGKmpROtY5Ch
S3UrTWuKdWEaJXGE0X4K/hBroa7aKWD2lwRGNfLtlcTJMhxe0DQXWd39UDayIK/1vhaetQTfXe1G
k+6EWBWdE4s25uOboSZEXPx52Oe0W6v/nbknjh/Vz5zGWw45tnJe/s59QbvbjUPTK9C3nZJCkZNl
vDuxHaIDp0S+r4QmHBb5hc1E5sIHspFbVMs9SLsSSyXvoAotI2kLRt3lpvYZjEBTD2O6uIubvSHz
Z1JoYx9hM7mYhnmdrH/yscQJgboyP3S/TH9ch4h8UhpKYfs39EMLHOcGXa10TftydSDETi3fs7pl
Ew8o2CiUuZ5lXMLy9lCIJXlLFbcQD/jX7BkuHMUCDTexJIl512bAKNM/g+ZRpWm7n8t4Lr4m/aiM
v6BKmv+cmadbN95htsoA/szbO1OPEawzBQgHaj+clUXKMqrlL4KE7Xvq3v3K0GhlMHuqrzafW5/L
WnZkPInnWdmdEbF2eYcQpESVuk/+2hHj7r8vOVVGH8qGA1orbDI3+wyMdYwPOTWTJCWVdRBlR5qe
j0qe8zlSqQsJWsG8/IIt1WxUxtVTpGLDhkAi2+4+LUpiZ5GhSLyah8zMNYQX9TJuCzAbfHKufRuz
qh4+j/4KkSQ6639jhb0nhVXgPSoBWyn+fNx03v04skw6h6wrAz8a9C7LQq9PyZc5tytd9yghHJbE
eAPfkQtJ9ohXse7eo4VGCSJFl5r+j0DkdD2aT2SMTB7KXGgz6jOTrBBdwx+7BZCPTCnXlohFtrHj
jvLgLaq9/Wf7hXeMQ45nFbGTtSrt7kantOvd/6SJtXtuCjY5+vyVhgMpO6030TNZi4IORZQKk+aq
JwfToDyq3wRYlzXjbUCMe9KSRCLm0lV+RIpEqCP2/y8fbJJi0PqsmaWjac5OW7GWrjaJDQR4q2sJ
C0ItJl8foVaPN35kF5mLD53INz6DYkapVSn7S3Wq7Adeci20pvZGEbeTWOVLuNbCmoFYgZX/JFdW
ylKFJ8UNkUIWIE3M4B0mTIKnbhZ50J+h2fIbL8biPlmt7sV6o4hBqyGS+WWTxLMyy5ILKcA6xhko
HiBHx9Ec3gn+NBB0KDhnjOH2IQeLJWLooQrlog+AYxl5cHwiKfTdGxQGOAB+OTPZZUp0d1o0EqsD
v8Rtyhgb49whhNwd1PzrbxeZvQGA9v04m7yOA/iRS20TcNNJBwt4CA2R4PxgcjYsNXUFjdogMoVH
uOxIfwPt1gKuX21GQE3RgqhYm39um3RAdpeZyQ2mZyv9ckaWIGbczaLe5s/lGWKQd/MRmCsr0IPL
i1xu1QAq3n/emP8plbrh4tblPpUisFlfQD6lbWgxqrqjGjyH5SaZDlZBcHWM6fIEfs++vFo7XCEs
/0yfSN7ekikXCZwl9piifNYSnB8mC1hvCsZeZA8XiNfH7b3t0EJz0siY9B2SGo6e7GdcoJp0Iu3S
BCzNZxaLY0eLgNzWLk5hxvU36EO8rcpEQSxvYgbQKEvv/Vd3YpjEDehAeVyCEO03h6cLqxSxSMSw
9OWmmLs9oGoFyFeBCEP2rzE+hFRh1cdphCnLadd5HrxikVeQ9dfhjRMbsvyl+4amQLA78BYl44Rm
MYrGcxcpFmWVOA9X8EUy7niokgYkRgu0zj3/cF+X+xJtwvyJ5qYsk1u5GMT38smuHFIkJ/zhITAW
VY0hAz4/G4UHjJ7A48/f81zJQoSslTwOHJyehy5hM1D8Rju2hSYS9hy4Hk03D9nvI+cv1zXrXG9P
KzTvdkpMSqxT6rDRCNyy8BV4IoxNX63pCvot9BAH5Fp5NLHwwSKhEd5QRcxu+3C5DAl/PbMgQap9
vnRQTR7RPaQIgQWxyIE9mFM2kFprXvVpaA7vPSCIps8EIb2X1/fTdYtXj7kKgtdMrkaq4KOKplqJ
UHne0e01gg/gPVhDGE1sLjcrbED5Vu/cdXJsj1Mgwr64pE28swXDltJPuwY1FykaP0GlMllXY4lt
7VMCesh2ZdP8KsHgOAnoKO2JNleqSGbu6iOfLgOKmH1pq+L08sErjRNR/cNKffjrtxo5Rh8RtWKE
4cJRyC50MmNo7hJdscQVDsDS2YYB2ikG1DXGSnIqxBUAsDPhA/+B1UwHGZ6/fj0PYP4ab/mcBc4F
PE7OAI41OScisN3OhQqy+CngqMtj1YnLwgpfu1UjdqHhdzaeSYmUsNrvydQ3qamu4KW3SnGJ/TMQ
Sxgjx2gVLkhWTgYdciOMV9mi4DplWRfiGLrVqyNNEdeEWJ3VkkiiupuKMYWimO4n8xtUdEW5h/9a
MJt6FCCZyJ592H2dzZJaZ2IzbzX2TWgexf2TuKxjhY6ZeVvWW3DCiv3WPRSGZOt+FjYkJPsrhRyE
piG5Tj56H7DCrRkCJY/g29aMbGMTrQV4VEoHobU1IOKdykqWGfLkYTIbxcNqDSnUQl8fGqa13b/c
64vCVf52sq1pBzJZO0IVQ8xwkqn6AFwuAGHKD1q9AXEALuZ9xV0ic8GqnjhPT1f+ebjajy7D79wA
lbzvcyzyji+ByP5ZiLljKiKJ/IcumUkeUOtgabRVrw4l6M3eGqdCjaPAPeM1tqCbxCgP+hoTtQAT
5dApBC1/Qgh0PfFtJhCr9SgcWpS5obajT52+W+cLmRwVi/sr4QediWNoNf8s1VH0buHz601v0IK5
qFBrYUiW9PYPPDNpdJSri4es0+aiDLgE2U4ggvnRlcMJv8Nod/UVOPeilDCOnoyF1pqfLemUhVcl
hatS7NGlIK9/LvveNqeB8pnbAgkH6hIKBbm0j8oN+DT9mIDRgK1QcD0V7837eIIaOXm8bDWv+nly
+hlWFO5LGotzgZWirfbs36z8uyZYbp4o0E2EPLg1zEaQXtji5IJoAIbegGgFoNTYE2H+E/vgaeKY
OqSdsB+as+ADoUBp3F0MS/Gw7CCVTnehfw5zXyfEX2/ccf1ogi0hwKNJe0hSDRhdQGuaHQTZUKcY
Rs/nnGo+5StJs3rKNXYdbxagXSMVTtji7QzwNLYJeZ6MXqWncVC0DLGTNPdNdFdY81xejE+DKD5F
t6ngXEeiIjf0dBEEXqL+XqIL8w4CA4sgbvDyIxpZWsrzAoSlt/mT8vtJDJ2FkHuq/BygsdMCIl7A
N6Dkrt2LGk3pnEaO1uQ+HBNZ8WgRyWsYvS3JYgq3pRjL9gkZfZLwNl0sJCbCerhv7XM/UklF9mqR
2eueKAhG5omIls1hbZdThIEU95sDyyTApVvY6aC1O4zbeLirbQekh3+GoU7BB1v9LEpP0iB8bPa8
CjP+e53gv/qsy6xNVH3qe5LC5muIUbtv0Gry5moxexhLQF22lPNt9EiOqCv1/5t7/eRid5SOV9IX
IhLHlpQuybxIfXyEMKj7g+dpnjB77h93FRGei+O/LBwj1uDWAZRnYLnFt3zK1wkp2tiSDDuTnXVh
ZBgzF12z+DCz5yCAJJ1R7Fsl54yShGzMo394wHV1g9rd2aw4Eux8WRyGZePSCIx+VCtn4I9gR35W
7lJByRvgwi+S1nqLoGQZVazvZJn8kTxkbpPBQBW9PUOrQnN/wCNBhGURpOb2L6h1M1wzxBvcHZ0G
tvy+5rg2ZC5FQ8r+GDrEjwcGCK2omLMs78k7cYsFwSi+xUM5sEu/EzFJy+Lx46xZg+FHKKGw+V2l
sZpX5qyCaz+3yCS8yRxBr64r0IyAgKUGPfBXa1dm6iPPF0e4n8xKmh/sHuntNGiATqG72Gvetot5
pDhGK1sN6HmA412pntIOc5Wde9tVFDJEa51UIiBayWyksKB0goXCiVMFTh2nu+5QL4hq4uSXeNSZ
+dJ5pZSMaCX2p2P5CwyiCWw6F4iTUH3v9shgK9IMKas04RtTbTsvcNnUOWf3vehIkIVWynKAiPL+
/YYCryxK7IfjmDzBr3fBLOn+GDaN2AAjtJaUiHDL7zpZ3ZJpQ+cdrKnYp1xxt+fo57v99DLciUOr
7NDYCqEC/letDlzSIW+VAMRVCnDCziXc8a+jhCVGIknzCw0Itpz1yBFI8KkPu0scXz2Zbu0fQnR3
Ogg6Ll7yP6Vhh8u++FcGpls/D+oSKkIzOmH0j9R9PM1kNEAadZsWI10TYIKi787Bq/3ToSq7aes/
Chh8/i3p3vKjXDPBAS9PrJQ7UPxzWc5G2wC/J3IH3X2nGdJ0tdMn73kElYBpkJ/EsA/FnheqwrDt
Z0n7ySb72btoUEdQTDNKkVPj9mQzbMutKjwFYxr3amzc8U4YqVBc7kd41bO2yi+2Y7ildPDPU1Bs
MqVj9aKu14449mjG0suk5UuBDyO53dlm2yyHWBlHUv9YEClK+3mvCWIfjxGaoVx2I9jpWH8M1yXO
KuXLbt7MtAQFEmJGcspsahS8QMrp0Lg/z4nNUYLum56stqmXfxNk3BySS2KGXvLF8Q+ysEzPD+i2
4gQmCzGWRYiBUyu1K/vJi7I6xFr7PRhRODAQBf6CrPikpnuepnggjWhUXsjhZwUFdzmKnBpJGX4V
ZDPnw+eKTRAsMrdGehmNSeIIjGVYiWv9amwB/VLlt7/iiQsdPEs/27hFXGhZratrkdCXGsAspYG+
XzcXQaAnoWNs0+ecm5wjZnZM7JzhdQrmMlly3NDZ6QtBkA55mStF9tzWCtFkg/wLHRZoQMhUwaR0
oh63NXGfXe2IICS0pb22Vpadt3KGZXzy/J9Ck3T+XfMiJkxxyzyuDYSYQp9QMj/A7WsdTLuh8f+k
j58xjqxAJoZbh6KlNXgT5ZB5FUhBCLWO4QAVJaIIVRyi7KeAxAm2Bc0ccmhXuf5UtyD8wU9gBKPh
XHzqGWTgIYDK5+JbRWlovF1XDcJtP3BVsl/As7+pSXQX8zCJQ6Xzto+QJL4GJTgIxBv4+4zkS4SS
jh8EWVz7WOKu4e3oTRVrvGson8P0PIasQYGV7kUcWMAn9TZFw+a1fWUHAVn/M+H3kD6aGo3a2FtC
O5+4KOCTRrVbUTh1YIAvikmYJZiwSMOKt29NxnXoU1rwYHNHxAUTt8gACDVgT2wFtRCSvZSvfp6J
QaGyj8CtpB3gPTwlpx7gIxTf5Vt+w9OMjFO8ENYolavyYChXbgpUgwQq1vkdA2SHHcE7phPebjm+
l0UqvcyXsJ1mKT5JJuPzhuTpUblmwP4u7gOmGGMFfJ9FYzRqKEHNp7JHv2hz448LS8ju+eo8+tiC
jjXEHzBUpSgpJuZFTqXr3ZTN3U1YggLfaU0WRq88GNWL02RKy9digHzPD3Rp3l7BSzz1bQp0EXar
WSORs+r5Zbq5Y/KVwmo5lBaR9rAJW0v76WvAUwHbe/20iov59Hx1E+8dDUntQapb2m+AR2vfbCDX
ez8/fGe4TgazXQN517nLscvDUJy3EoAywP3mE6Z+XN1ZIXyDTG2av7xRCSmb1A+HI2qpNYa+lPXz
Vw0bC+Ynvh9evhAM5tPhGEhOH2j1I+fUiWsSimWz1PrIpzxFlmhZeIqxPZ7BML7g81YjN72sH8V1
q4sxLqa0jka8AZktxoz4uKzDNC5p0rkq4TjUZJ7C8ZgqmzX642i8qCqOOPJapaKHQEXAMuyy0oF8
LuIH1YUC7IX/8si60WWiATm6gHmjOKRtIlPIqZEm7kCCWQBHaAVvYSnGatcuABvf5496/IArR/nl
to4im18AGSEyLdUZUOYmlHHV4P7GSjanAP2Q/b3ts5T5g4XG1U0V+3CJeIql4sQDC7JUHs62ghZi
oAeyy4cQ10uVsiNIuGT6HgtHXT8h7jG04iprPCqsRsd7HSclMZ5CMqShRmCcRZhb4IDFfXV4R3yB
w4c0DUq98Qgr5K09NyW7SPdpEvW/I3obifh3pbkGs7VqwOvEteXWstpVS2EAlFm7bK0QnPc2ihR6
dpgujcRpaQkfHNu0XFAFWLi5uF1DTzNoxvKC66Q9VDikkMjsrPcWvsKvLAvBjjguQK6dYexbxnQp
6YI6+MMtQ02ECDWCO1xZLThGcLdRgNwGqT+a82fiKhkutDaMY1gLUrBzFYz8imCADphutxpTRUY8
On4WW3JmaJ5vPgdb6ANY34cWe+2hqYtaweW1STQE4u9T3um8YfEfyvlnwePBVDtfxYxh/YF63PBD
j/Q9mb6gEjLL7TFDnmc69Nc6eT17X/oiG0oy6mLZj2HdI0kD/O0xSmzDXBlF34BCCkl01IQWXnQH
u6X3x70Y4YTE97bjJy6hv/Cj3U8Dx0lrISxFGzTok3+KWzsHez9tvOlaxUqkh6275wofztrzn+kW
u2Ddax1TpwH7G7jhpD4b+llpq2s8nSjvZWQoo3s73V5x0n+UqTf+8rsYB/yvVa0zCBqdoT9cOftp
g7htEIXjtFXDs6GV5QJb2Bnsljk8MzhN5LcqQyUi0kTkWNKfzxGmWjnNCi1jrXXQhanr8OgaLEJI
/jw6MTh5WTr3sTPqcM0zRHyotlpTKCiih21aACS5o0BzEY49Syvq6rUZMJm4ETVPUC3StxMKcB/9
M6vnzda7wxuTW7CJJW0bNrvXHABFN+wkjUW1hcal8TFmwCKydmEz3wyo5IO7d8V6Ph9Mx8ukIF3M
c7uIO7U9cNZzTytgke0f/XLTY9GAtkvj2aho/jYLOtyFW/2Xgj1SgjEvtZVO/0gr/TQBYF2u8UaC
VQVM2zoMQYcjCzcl/Og305rKQzozaIgsTVfCzmIq+QMgowppWcZpm5mwGYTUQlkpNfApq60lH6Xk
RlZc3Ju3YouncgQGbECfP8MvnkERZ+O5iG/+H8WLO0vRFquviS/Cmns49DCKB8sbmQlB+fHlTu4c
MMkwmMLYYb71/cSq92IXDtC09S9lPsvQVqO2u2nxaGdJwiW7VPreGyBq3+3/aKt1M5kzQKjvRkV7
ClZEWZwgK+PYAFN03a5DJAwn0G1D2ntg0IDh8glJVJigtVPzCzZ0RmJabqMbRPZkFK/biALexmtI
U41wtkd2f0Ak9R7D8F08d3pQj+2uYM4tfXWvaVukMN3AseUrOXW7gqCecrO8ZXsnCJTkau2NemBB
Hxz43Tib8fUVc7sWhVEPIDIGs8PlTSw/aEkXS0Af2lO4Cd3eC5u4w3X1IznN3nhVBjnY1oH8sbc+
r8RsEbTd29JS0JzajRvLdFquaQaZnesx6VEF5AxzGbunKYGg1zviM6zHWVuzQmdcZt396QaW9byU
IAi1UnsW0e029Y7au5RyhOnoN7avMjA7MLNeCZzIRtrW96xC7QwwNtWAkTIuACF8Ef1bgTk8odJD
fOM2j4ePP22N4uwC6LphXubJ4BkY9p6L4odt1BRULxd1IoQa+MF1M4C5WDMs95qVhZVKlO0wR4rf
bVyN6hFCxefQItbfDT/S6+LD5nUFicGF5TtIkX1rn43AkdnPvExuOk6pgdebt5lGX60WBGwgj90K
Uc90dLfowwd+DewIgfYhFy5llFj6eaf5C/M/dSSYZHaWUxq2vX+6Ozr7vVRnPIFfTWGgyPvL4UT1
8vlrFcUtaiKLW0UMfOZ2oI+6PKajLuM7XZNamfmYWfYmjjXdRPVvN7VJf849qhQexA6jHLlrLnJW
PMbqJw34O6pnjXhHeU+TP7ckd/TKl7XzKK/90sxXUTpLOVIm6nDgmdXasWT4UR/hAacuw/zSRw7s
hqOF7B6emq0M1Mp2HWZtxn7ICpEhA7ycBV1u1CQvJwjZwfk1Ldc+LInf5BWWn9G/a8otigjyy8yh
QwjBjwG0QMwqdAB7X6TKEB18AKx08l6H1VH3AfPBV4T5s29JIQMUK9ZEMs3jOtRlWA7SS91acU41
78UNvVLd7AB56o1uFfJlw5VR10e4fLlK83H6SjSEVzcYW7bJQ1E4/ZrxcqZvuXRIlTcTBhNIarEh
HbyPzb5Wdf2lNItBMeP2PJGfdSBF2D4WPjbYKBI5tvBIOaCgoZhC5n7m4PaI0xoms1Y+ROnZUi0h
83QE+h61HvFTePeJLTZuefkgbbuud9bajS+HlmLTCJM7yuoWQk2f11m8glxGeCRk1/DBDhmg/YGe
KaARaGaKLAPcuaIfch+PSKfNpOUFH8E1MjDT9WB3DLrX1HqVc242HxLo6yJChuhfRTLHaawGoz8U
IbovEwjkpmtz2EUd5OOjYe/0S0yIinyTwT+ks296+OA9uR89nbUevI6K/slBSBCVcajykPfENkXj
uss10RYB5c//PIwDL6w5Nniq3RgLCtgSjtTELmCpFvIl9g9o9HD4xEgHYflYc0ijqMFPZu22ewfo
HbAZgTU/sYu/Cw+ruySRiBLy64ulMxbXjWPgoyA8yTxs4sAjxCPyKjJCrTkvuZdh0PK6tV20O1Op
g0jtQLnc0p3GItnaMBXxDwFEYFQv4SKVJeD6V3uNAljy72/EHZTdQeH844hrH79/NA1fKl+jiof9
e73lmTTjyY/RkP0DnQcBnYnj7PaLearp320gxTmhZkleMvbTHe/tQOZWTv9+oyjjWshOduqyV0Kd
UhmadVcvvhutTyU5d+5jwFmqm3CMoAMfNNFnXH4bcy1+aiUzZFb1RxV0PwakQHmFOjq5n4GZX1vS
w3Jjng/lmfslpBFh9Rb4EOoSsOByxCHJgfP6CIFfleBluouwXPZbPtOfJB9sVCKQzoDALsg4fZX1
gkOU/7e6QrC5dVI+FXwNBt/f20cvIHZwduLy9m7Rf6pE2M53OR9VLgeBsUGwdlBaQoukAMwJWLpi
r3TVXEXEq15PXh0wD8nKTf3RedF0JLPxXMjoVMOcbnu107w+N3syqGMzeNPtGOcxi+qDZ+Iv0Kip
qjjo6r1m1Ly1PgEUIQq5yrVrCENCb8TRNWwXe0CktPFOrvYL+uz2XOM9CNaXzEbvoOWUsHgiVSai
H+owcDctwoGfFtJ4gYWnRYpQlzfm+21jgN2MXadGvt2pRd+C3tNAl1ymsIyhcVJqzM9kOf7BIp6s
cPyEaA1Ea7boK2IhIFL5gs7Kuw9IrdjzSgki+FlI7OgVd2L7fsXVUubkCngFcqJ4H15ZuIlggZii
zeiGpwlL0wbM7/OpiRTIMcKVIWeJB0EouuqEnphiTEOTd0G49MxUv/xKtpLLveZLCxfY3WbwqaIC
ELYkVLezzTxpyj5EAJMkOacRxHwQjW5rO1RyMRR+h5BthUNd7+Dgikg6rnFUo1sGpJGRUGcd4P0c
lc1iWwJ4pALR3ohMLzALJhOUxNufNj8a+Vdr4oOUCg3TMPpO4ax71k2/pNX8dagRZFCdnwOxWbOv
Py/1xhv0XaoMwbD7nJ0bPQrmxdZpK6zOYB8A0Vwu1XT50mlviJifh05daA/xxK9mBdIDHL8m5wlb
e/Ijlb7v9vQWyBLPR/iA4yaQNBj2SW8EFG55VBxhFD+uN75g4Zu3hNkY2YLOhpFcy8iTt3Q+KZhb
sY29GDp6VezjIk+0lVAjF2WizYaLRLnBF5m33k9eHOhlP9HtMiIROsMJ+cHVF6MeDf5/EcxV1tm4
CZ1AKx/2VVjXgnDxuNq9g7TyhTEo6zVYPQ4oJ00RN3+dJWnHgiAUG7VVTScHhR8H4vKQLij0rjVS
/IewHPnU0/VgDYAF9TbUlkxhVO+jfoWQx4/VauvCAcFgY/RZ+HMdwjXmFcGDR8WdQriDOS8kwiCe
SQAoB31h/fHxUeF7YpcEHYUISftSuwUVHWhGd6nQeni+Y/c4RrU9FXX9o+UI2/3eNX6SiGd2Jk6X
0LDNx3A9RhWivYOF42sp9XyK4U0qNOl4Fs33pVQ1qERWhQ+6aAyITeCrVA8FCEo2Yl9dA8OMIaJX
Hx93ULai+ZPUNi/GCDGzRqYF9EDoW42A0ZQOQMsNgf/s2tP/XnBD73s0YDuCowRR3+aTt3iVD3iy
EdBPFSkULfo7MHDRjwmzvESQ2HQVuHkW/eDmZYl7OT6mWS1o8sfKpgUQS415zw1on/4O2RoM49G6
xATdHQ3yIq4SuX6Q1JQhGN9dJZdO4RhqLC5ccL+F3RG2Xb9lZUHD1WrgKmg6Izbnto/haVc3QARQ
vU8La+J0q2f4LIiBOUecAHqGGtxNvpxWIQoh0E6GF8a3gfZAUKOqk2JvWUgmuHNaoclcHhE7ysm8
sxyQGKOkC++SEvjDULPwoa3T5elKWiyVcx89+oYSkA1x73lFKiT/xFF+I98BPRj02hXG+UZovro4
3E2FULIJpNImBXKDNMpD1TUKbiZj2WpnmA/RO5VYLMXp0X6SqTB2/XrDCNNAqr7MzqZo50yoGf8y
eTWVl3zeZFR3EdwbiQ3qEsyvRDe0MasWHRG2VLmSPzhdl10RwTMVB+SHBvcjipgnxXamkyTaO78l
uEGFdLl7p5vRkqzXal0WK16FcqnWUCqZL0fbINTPOssN/ZN7lZ6iZRADVgx+iN+PmVPgV85//0cR
OeuN15TgWcob/AKxLsGT6W1327DHjTQ8hAnr+yhl0MiYoYFn6e3DuvshEAI0O9VVPTQ9jh+qwSqN
eidNqTFeV8+09mhcsCCESCmfj9siEyhAPeW7bhFcF/2iIFur2umT8PGmmcM0tdTtH/kpQL1x7ezO
OmTzRUA7ju/A+meRa4rGNHcKFyKTdFg3dAyuQw8GGo8KA+yZY46pamBPmCCSEvbNNJnPx59UDcAb
0zuGJMJYL7AiwpHJgeiltXSOvX72UvYFHrxG2g7dJbBi+m7Lop56KKEawKP02GnkYWensDePPKib
xCYxT9ZlhsSXGLMpa/EB9sI3+qDj/cGk6+RtwH5sc77anEXTgo0RAPUAPCpN9GPyBnQpzxF/mWoQ
QNt36QywmtXCYyty0bupZWyNz1Gm7h/htL+psaCfIn5skzBRsFPL3KGa5CJhOuq6TWvLJZ5oQVAG
ex0O4G7jwrgtiyd0fY7jUbcRdM5FHsWt9nllwGZp+6Cbq9I+4VpFkWhFarxkwSCcMOxc1CJ3o78H
KpUTmEZsvyuxQ1boAXsqMuFI4lYRXy7AL/6PvExEoKwN5C7rfNNz8rOA8MWm1DeqaQbgYW+HU+cr
uG3LPKMHrTlo81CLs8TcqpipfgoFipszLJSJAsyw15wVcq/ip+uzF36uF25sRgtvLfX8WTcCzJrV
xigj+OeM+wvghw0Ye/2SOrNV351apUqBTjDYRB9Hmlw1KnPxNZvGERWgFs9euRTfF+IFDQt6GcBC
pFXhc2uU97KEJ0QJZdAllB2oWC2XHLk23Xrq0wE2LgpXAB979qTPutEqAfu1JrwTgzq15c0XrkvK
ONKGK5S5vU+7xc4UTnumjphiUoKLh/GSBsssQxwIt1VMujfZSHTZVfXyzQSfz4jq5aIU3osYL2jO
kBubOwpyNu+EPMypuhhMIC3o9sQa3ft9fXY2JZd5W4jUY4tDpmp/a7TmPrTb/+NX+ZEdehEGx7+T
7V+oads6+940BtUSqXTXcW3t+yya0ETRZl5bI6NQ9+6jn1tfzE8+EroH8n2CaOkxymnv9YgwH8yo
plVhPxSgjErgJzRzvykQg8fN3FJMeDKMsHkFS5W7cudrzp1j8pPxcaQhjV9xaLncjzcq4dxd0DRP
njMUyPsdAj/OpsQxwRs6sIjz92E7VNQTLO0WmyskJsWprvx9QVtCL6LCazCTa+2CdIpJZ1/SGIEd
sYzkWZoPatASUq/oc0Auplaom02K2W6QDtapM53+rApXgOqEuBBF1sWv0IwuXXpzuqeU89XVEMlN
Obxx6k+1vgVNNpf1EHen6a4xnT/G3X99ZJpiEuM8eU7tyCK+ldgmkHZMAKXr9czP1vbXtrGRNOgc
5rufS/lwLUIgMklRx7ppdcKPqrLMU4axoJrBQkbAILgliKgjkGw1UgYtG0FbIQoC7HNo/aV++uNd
T3jV8tVmBgHqC7goERRX29SIMH2O0QQ/sXaeXFUOIPsXZOWt0lM5eWDvhpG4HasSpoDcjzmHRoCq
gdU3UbWaTOAXaayiWzNCE9amPa/6ZB634/hhCVMeWYgsEJeMJn+odkmGZHLfhIJLe+YMjmX+pW3X
PHoNkUFiybOL7irdEo4QbssFl0TVvEV0CeudFTmxjvaSQn+dSopPOa5Nnqj17pBXbk51BDsh/Mqk
UOpb386qcqWdH+p5iLdaP0xIZJboN2uJBIU6p1lnsccNk+nY/B9l+gh4o/Spa415nK+5Fin15L0B
dcj0MODsg87AJmD6V0OwGkJU0GpCx0qBD62eWfspQOeqoUBM2X0Eh87eu3ZEN11a0KbdNGKthNyn
UolyKUWXjvuizFTZnSbO2Iewuw+CuqkaCn/xVKIGcP7W8pHNfya4ASfQHXxCUtkcALJlmeQiGJar
6WVFJhgssJhr/khmDm5arJMQqfx8URYQj8KtU6Gn5Uk1Y9hS5fFZND7sQZvunQM+jUPEGLCI8sfD
OnCJ/i2SLrT5mXYtGfdqnUOyrfKbThkYb5UN+0c1akRP7+x70l9zX1+8z7vfQXfOG8PXDYzjx8G0
URLqjmMcO6br+jRZGtuby64FiqS/hEKTXP6xCj4h1+Lg4vWNvFeQM+uw5QGv9wFjAqc7i+XmLbKE
pCUC/HE0OY2fdDgk5AXzocK37h3nrg/fBcfcOLSdBJSDHpUzf4fGnuAkkhT2Is1BHco9c72Lg++G
If5NPmtSHYtpZvj+tDUPP5i/RjoWOy2cNYAqAH9UqnmgBu79GINGPU5FDJJRnTe+wkmwg7Bl6LBa
FtxTFQjflIyknTcLVknAh8P3snb+KLASfs+pQvWVl0ejstnTl861iHf5lbWhykZnPT/VbGj0rT4M
jeyUZA/kecQR1Il3mCbAfwxZedzzLF2ql+pPXT0VCE4PrEZbFVnpSIDhd8u3jO/fH2/4002rgpl6
gShTMgsL7KcY7iZDWFu4Da5xY9w5Dba2SjFnpWv9XIcP5V8XTC0zN2+v7L96EtB6//N1jm2qJdGO
AgIBmkjx4peXCKcOwcGBMgKghig1pSEISZlLxmCpGF9ouuCEjVozczaYQ1/b5Hoixh5t77+mcw65
c6SsU7msUVNFt6gpg5mBh96B0WF5ZWHhZjhDzkxIhUp3rjuhGIcdX0AqtVO8DhiU0FU22N3W5KrR
9UmRLgPasEy1gd/hnz0pK3a/Z63CJsMWAn8xdMPycQARteIJ/Lcy4wNxfZGB0j+cQv22ZIY9Bt+F
+WVig/ZBaMcYdhaNdZivt1aKlq/advJDa0oh8WVSJszO+bqwV9BvLLvbzzQGh9skvG1Wkb3kuszA
l7UMqpkNYbSMoBpxsUbJ/7XsXnNrZihYcTDwduXCuxRMaXEMPqyaHCvNu0b/q1O9mpuJvztiTAbh
jNe4CABx9K1zcJQEZcF0oEZb6wRHBQosrznxlQxD/MpBh6UDuDIlIfg5ocAzjprHWg4yuWWDR+qm
vR+jYmTAlPs5C8GRGFsNHBg+K64LTQo8Wq8cjIh4OkAaSjgWGGYlx9kmX67yfdnZ+cqQEQmF9x/n
QAuUGyCf7g8ZKJRaVORRF29cRnwX0mpgSojgsfZ1DpwIf0pg/p/ABJ+owUFi4DQOwsUyQj2rJDbd
oeoTVB0GCs/J8by4QQpgpRszY2mUhsjAC0M7c4JuG2qKNpYmKpoD+OXA9VuPKb7ZtbWC7u3QmY67
TqpQcQqQyEtPPUVWkcqLH51wKXPLrQiBpXIv/8jDLsNfwFdKCQ3tE+FVBnZ0hBsNzfaqx1uDnnVO
e+tZb8sQQVSoWRAzdXl1XyNCRKy6zgIw+LaYahyT4kERUUDp12cCycc+eKBMfA4X1/TvkMBBdXIg
0uUmkEWkexR/gJyzN4GvzBfW/4MGJKlFen7EWUvvxwupvs8T+5db7T9YmABgVLQnCASj3Ow4k4if
X86GLjDWJSyl2AdIIHJUh53gyIlCCejBEp4586xITSBmmr8ncyPY8Xrti8pYKFtm524hO7wiJWB3
Q/yKF86+jKDlU/dq/33Ood8J3LIPbQ03UMFDzTa7J3PvlqgHWrDvT9nnfn22MM9O/1G/qti0Wgo5
1mQ7ncj88IiMPuXdY8jzqMZONyENzrpQcSo+C3Rz6QauEAiIs2z70t5Twn65gzhC+P7ru4cuW3C8
r+pXFL8yyw4ihUptq/Gmje60jds1zwsk7RV1GtRHrymfEVM3xEm557eyjavTBjtav0wdDYR3Htib
GWkR1svGHc71Q3WBSbyp3L6JPREwU3UmP+cvhe+Ll4jYcrTUUmMMZYjysU6sPaPKe/9tNAbkkdBn
Cq/PydzAdVdbaC6ttZPi4Xurs9LEj3Y/qpp6HIU64f1qQosAS2aNDX/ulSqckj8NcuB20gwfKU9A
VLNDZ+Eoman3EWmhYICzc5vSzxqL5Y+nbQtnXCfHrz7vGfwogiK7yQgsg008jdMWmT5b8WWa4maB
YjMbS+D1nTSniX+/AzuwDt4fiTWuCU2V+sP0oiTy4P5OBYwqE5PLZLdfSvtMAzy1LgbBz1eTFqiI
LToVdZ3ziSEoxSa8x5QTM+ApWWvAApxojLTmrr9kBViLfnXyG0WAh1ygUfqSWBUAIiOiS0IljgMN
x6zauwq86kyg73nyhLccoH4Ce9z5Z0aPLTSe5H95Kt5nwgVTJ1okvykFHOGIWijBagRtPkE/w5fc
m0cO7EMdfq1CSuXLcPd6DrH1GFGiBPe2USDYEGErlMk6046hNN8DtFQWk8YSQ+IMGgcbheQ7+aRM
YE263GZKHyT6x01jWyAaGvDJwMFMCyKLo06+kxYGVWqLBGyGaAqlfNMaFWLH/cy1qKkXyum+u+Me
AiOvm2oRJAZGJUzZJ67PaUZuzcNwyojPlAmcFkaygKLxuccOGYWPlmsKB29Vdby0gTxpbIZlNVc5
a2daPsrWJJQTt43p5tMBixmXJBbuDVleqcj6MRU1LrGWyXQFhVsqMMaiDgwUUcOunZa8/49NO4LB
g9076KUpts33HFmlYSrV/o828oHIVB7HCnKNB2SYRvvG4ZgO1JVZOwHnKTZc7/x0nfjqtEoK92V7
bhxVMhArw7tSTTi6RhZ8SIOe3DNyJL0Fqz+r1tQZLFr/OvOJaBrobMKtgFx9/OitutChROWTUmxL
HZCGw053h603uVyFfurLoAq/NJ8nFnNk2W1pXTop42wUYB1XvgRiZ2THXvlpSJp3RRcNihJQMb5e
Js42qJOqsUvEjnbjT9l7447f7zSgx6sepDXeheLF+uK5fqWszWHfD9PDxYrdhYaEt2J5WvIk5VCX
AsV1QsmVbvDA3hiI43ExVfytpUENnafa31iPBzTLCSxxRX3TpuGQgVW6t/t2OfBE44cLruf4j/dq
nyrUU4Uv31tq//FM7D6XTm6fUY2tqtUfN5MBYcQ8y5wqreOh6UULINaTkyUzPiS51FFcGwJHrlOm
9i6U5OX/Bxlzi4MdnaYmxHpaxFA9Unoc4lZXbsTxpUsTmKV9mtQiKae1vCZ5wYk0JsPufToJeicx
utfPbwNt+hvyWzmhpYPHqbX24Os2NpLf00fZZpa/mE2019nO/dlGT/Y0THWT25LntGCBGJ67YQji
k0kElIq+vW3N3RU3VoWDv0jeCRQF7Gb5LnU1ilRc9V89q6t/f8wT1QP0Y7QISrbul/m7V14BuYIE
mXDz/e9TE73XX+EIxavFMoKWJFQhDMDLxv5e3dA19cEFxJkudJK61d8KS3tyUOAn5YsuJSRaHEXx
CjymMCAqYwNdV2FpJhh4ofFDndTyBPv9tD0dLgjwXKIexvt4PCY1v/6/G9yRzUznHFRz+LGUCkyf
6vh9oKtQxZFtuugXs8Ude+9+aku0aDNdaCdRTfQU4O00UMAKyyWs+i4PZWjv8V4ciyW0/0iLlXSg
HY2CR/KaG2cOAjRJz0k0jldoEIGdc0OtN3hxKcaKO3qUzKl6ZIHMCPtOaS0ujT5QiBCb3Lj5c08q
djRGQ8m0a2Ty6cOsRUehjrvETMAOiYG1X5yPgHPg0Qvp7ORFhdPM5HrmnXfWVkEuiH+M6LqrpOJ9
ouRr/RpmeTWNEHC/YYK9jrpS8iO7JLseCg/eQluYVwRMRvnw7TAylxBpIZ9DKn9mHgA7nc6yvnmF
0gpq21Wj+zBvarFBzXArEx3+7XVUxMk07HNKjd4PdWBV5tOTFpzrr9jL3jOFddRcGXQkFcmGnzNW
ohl/7DiovUYajcPW2Q9en0OzVNmfDDLkG8GdAVQvA0g4kw/q/LT8L/AezY3W/3DdDhYWRRPDZSHT
gGD/4/GuxzOgKJIXbHZCb0DhHqSP/GjIAbIY9MxBCrgOH45wZQJlsI+D2cRaLepeQ3JslBphajKV
02V7UEXScw6sL1S9JPZd61MziPtvxW6jQ0JCY3h8ogoY1Vt8G0tBd0PhfnhBIWgX2lYDiljq5HXS
tNXjRkofYwl/dltVPZzDunLUP4sJO9q0wA2cWHOK7JPsIqIqEpabnKGdMkTUPpzOl9fMhkzT/d45
klKpKEvJud2JTGBR5PoApuQcT6nkwXfrEwQe4LhKeaF0/4U6wETX1M8KAg7fviadYY/bNAlzuCEH
8U4IPeFbuxdKQr3lNa2HsRlG/Vnn2bNq3RxYlmiqdX7lyN3BRrXUXg8rd93JoMioz4oe9mgg5boy
EIqVLz/qMrMQoAQbfnOoHJuadOVHFlLJfaMyPH9yEIPtsplrPiB2Jupx14QlnlXWsvgEa9kmBrLS
Xx/BlgFQFWA6+1TkfxyrxsV0r5kgcq+WL/um/e1YFd+CuWU4VnyZfO7epTPrKkl3ciZfV+JM1X3I
1AtM0lENKoy+cnDjgsg8sOSuuBYZDQbxchjlKHhGoRgU7tCHi3whww7x/TzPinzgmE6r5zhXtEKZ
HAE3ROBtAwTdRWTUgtyvK3EK2AOzAhJcoQm+mWNgjejqRidE42hrKi8ET5JVxVwxJu37TfGjuiRi
zXDws+L9M2zspBOcXCkjfYY26opf0DniS+FNLwenPyOFgoljpoqHHfMAdfY1RnXnc9gvP0dWg6jw
TsyqFLOYFd+5XNQrxgjna26KCiF4DglkPjy4riG/niCY6s5VV0T/lYS5qVrsIHH6R4K/BmTU6Lsm
ajSiJHNkfnQwBZ+L+a42Sl0i6oKDRDqgf5MsyJEK3uz7CDft6w6vpTbDNSUc/k50yuAgCTUIfhxq
NG6D48Do+wZt35Irdir/2dknC6/xNBl1jwkXMUF4lZHngGQTUpv6G9+jYxPz01z8Hde5tQ+a1nwR
xCdWi15rDyF7pqCRNxlCUa+UOIaXg6+u2fP8WnxXGi1vghXcQ62uYGC16eszuxG125kD0Y2Es930
vLYwdTTbA4AfFSlFwBe/dG9sA3zy9vVo6ggF2Uzy6Rz5vUFRwUjsspxVvoeG8Tm9HVUJrIZ6KzH3
L7G3+to6qVmJpOpaWcEDgYlhTsG4g73oo78eyBQHEha+BPoVwR4JAzShWTGccWNA/W3zirCaoa+e
1M3gBYE/zje8SQU9u0tan0qEr2FIcWs7d7+3XssI5RHUCpjXXt7yY6wwwxNf99hFzU7Iq5lq54pO
eOgggHKmrMgKrFMfum+Iqxe0wI1/KmExWtCNjrteaZinmnCDLWcjbYoWtnNuHA1roUU/4JG7s5fD
l3BrNtJhe55/xQXlak3l1PzJTzDkCsx5a2Qp/uyNzBUfFmIYY8mMc4XMGLV5D4o8LbRvAdtC53MO
wo6MLQRPljPJmrRi1B8a1UDCUYaYW0TBldjubsDTxRbIzXHWX1PAHmb0vvCanVexQXk7y+zDZi+Y
MdCc83GSHfiu0IrP8DIAGaY7jJcMIMUMwfluhER1YvCP9D7aRpCF+88TvsxRwCYi0CkskED1eayO
DXMxdyxuONgNjg/6ZYsqDN9vmFbHtGZD5crYy5B8iBlhPKGN4MzVaw080SZxzUNIvQ2xCjxxYkrQ
kCpOjUj3+42ThKO+2vvkCUjQu7XkUtoYWABqvpim0eH7eiHENCGoK4LiNe1+ZF607dFggN83OsBk
eEmego5+34NfkSoE1kHaa5oOmXov/Cug5p7WQPvbHbM07xeeFwmSzj+jE78bITfXDkCVkPJrnZs6
Db7shaw6zfKAhZIT3U1G37gU0z2efJ+Y8htl740XFs+YMxulNM9qqwfgdWHYb1BzSCukWZ92FY+c
vjTKcxlWF9iunW7a65O6c0G7C2uULfEtCFnuDqgQg/vrh2E3ugu1NR8WQxzMeScWClPFu/+QswVK
/fUm0U8R9YtNRGKF9J1bdcLrOghDOkG2s1PXnOfFB59s8jiTxOYTlol2bWdHkwlrwq8i+gBi5tM8
ReJ9omXOvIF/pQhynRzwxC2nD0kcO2rO7P6x9P0y23ykdS0AuVn0YaUHqS0x9aWgHzZPul2xUPuF
/+gfblpLAfkfKmNMU5kKhV5t59qCKaNj9u7HWEpAdidHgX/fhyrXh9eqof5+LoS/LfiA5JAhRmJz
Zs6LuiW7TZKUVQFKIao5h/VU8QP3oh8uSBLiaeWU6nxaH/TGiThQFqdw1pNFZADH1SeKA1MkqNA/
3ExhUwAAfdfrRnTwLw9m2rcywrPJ0yc7H63GcDUtuDuVHXqy3xZMOCfrB8UcXngB63t4VF5bFn81
ru+ZRaq34V4Dx+j9NgP30uo7kWbyR/787/4jWqwra75koSnIZy4YIKAj/83kFGhSxRmf3P7YltN/
ejPiPlLRMN8Tv4mt0heIh9x5JmY9W5jZEavtDlNewDrs+E6KXO/lhejJ5PprFYnLL9zT+r6Yc9Y/
K9mmoAYLnEIrNWinb5IxcFAszyvLVJqQG9vPccSe5E6RyQCF2hgMpEf0U/CcB2cbYuH561N1xAw7
T1JBpPnKgT7qHn4WAUzrb6ASRwsMw7rC+OOMVGt3Ak5iJqazpptVijvvOk/u1ja6oeVIs0vxR6Fr
q1CygbWAdtjj0CFy37KfGbB6ttmxQiGZRGeSe2D5w3UYpQuD/kgmBFBHIC8AraUQw43YmAAWt+8W
KICIUE7phnkcrZir1MHU0KKzJVdTdkTMUbWTqbqxdX8HMSj5ywZKReWpV2VHxn3+rvyalaE95I5P
3Cx8WTlUCIu3K+24B1c9Wdy1qEZhPOgtIN6MfgzQVYIhuS5NrLMSCmNkzr1Zd1paJx25zCgpnUmL
7TLhGJv9o86Uuw/2KOyJN0LV+pgdCk6buh4DbWHvFNoCSqal6xwxMlveLQ0O68tJQb9RcLQg5LJ0
gY6JcT+efykB+encvOGb3uEtsogmF3CcPGUg87dZEsLk5L4i9j94jX9vjJMAmfLoxvwsuM9qPwE1
H2jgVShF4Ucn27dufjetencxT3/7MzzJWjwCvIGMSEuGBoXupsvfF9yUmei4Wc9WCkW2Z4e4KNvM
u8TY3vkqYcKFaj1zWSRkYyS1uK6IjIDj/9xkeH6mxReE2mFQJZAyfJqI8Is6uHxQKQw3/g3wVPT6
3y6kvGhP8z4wlndcsBB++pJsbDGxQnFPiY7mxcfj+0DQlSuK46RSv5OKvcK8g8/2J9Qej8eOTkbc
aOKi0anSysy0NmK6rGQJDzICJvCpMQqdG/zsFUIAHyzouAfpVtqW7C9ye9lb+pfr3ydP+Inn11QC
69qLIkt1+OooBEbKvYsJmOXc2H55Vof8mL/7yx1SLpukJmKbW9YiqII2wZ8bJpHq3bpaTHehQ9c2
hz/enbmyGsC52oxiRCWNPrumaIQmHEe6eR0h1oaEQTSWkCuqA/gUcy0A4Pi7V2RexDNYutjCmWzq
uCsh1X+2Aq7rswX17Xicl5mxgWQwA2fXk+qZdDMLUcYheICEMp/3VmRpRcNq5BkN2X7aNeRlUnd0
l3+MJ6uQLEGGf/VHUz2qYnc6mLnL7mxnWJHmKBXpzJ+aq/g4PT9hiSGxTSnJbydpjxzYeYeWowpc
gctVfA2H5LML2CCAKgka0cteRhW9he/3EiWzuJGhCTn1y2FDoUcoarff3iEvtAgdZthvtViQlQNn
LncZ8cgUWAKCc/jMxCillPmkfoW1zqiaMeEMeNp1x+dOhVCofzu6AZZe0EfBB9zyP+MZ9gtlTc+C
bgwJbHSOz6Xue5u41QMsV15NxO13FfvA5l5VsRJIGg7PF/5sTIABcAAatJCIWcHyigvM3UUPw+li
ku2R8AgdhRnpbGejJ4YGWTbBfVIPTupS/8SAO9Ao4WLp/IiWpB0QkFGMTShzr3mA5wUIiWFCNQCD
kI2bWusZ3fUvSgG3ZuhVJql9CWSZWrqgSzwNqa6TLlksNC9ENTvOBorupJBXBDRh/MQjiwVuhtEK
tKka5itQ9dgYba6aF4sIssAUhjft9mAMWJ4n3UcwOxEjAtVZb6CdOI/wizBx1DAH26jDHg/1Wqlk
rvKJZLlrSal8UB0JRqi9gWkXlV07/EA4UgSWYAAU69z2UeHxqAm2lcRbZ48D+LAt8oYYQGxHnMVz
KxEORt/PraRerp9ty6MJ0ujY1XIvGj6qY2R7wua0/qI8xD2Zp7L3AajqGZu26l87fJcgG2Yl4IKX
wCRHEudZQ1nnummVC+SegE0eaNOQwmPDdkmF8WMljcZtVEYOXNQyJWwSy7N3NKT4XIb8H1CMibro
hLVUMO0ZGg/tcLdvFcQ9MXdQNsHHj3gqTl8Wz3WkDZDvjs69ZGNcYsKBev/Zo+kSe4Bs6xZ6/WzT
MZ3VwQl99Z7TLrGXVevYt/gJ9+XE+Q/J7kyYX7ugip94eYlMrpDwm+lE6e9E04Dx3CofIyj7Lr2d
+vevsVWrGMDU7F+3B5niHdcP/76vIRN/vgUSGWraLTOKeFWMioZBHbkebMgwNAvskddK13vlaYHA
ytuAZyP/5XoYM+/KMbSwH08ANG2EwYJXlE8fXTQVaX7c/nptYTaxPZhdRxXu3+B3lz0ygnELbVDg
7mIGH7q93LmqD6KnVkywLNkJd2P2KduzdFEiUjmtqNdhwTM3W+JLaTrvSh+swWB3eYu4qEXz/Fbs
mhd+EobcpH8hUcE65/NHusK1GmhWxgXQ/eUGSoq75SHYTIkRofUix+oUMa6pVjggWu8nyi7gOg8G
ApQi7HdOujE7JxrBBLpWQB7mttY1N95sb8J0OOLhD98JHAq85SY8GMgBc+JKIVCXLT5LNkQyA/Ul
c864L2OorYtwp2HmmeUd2q3hMuwNs+S7mWe+ZmwtkMweL/Gk3Usvhe06x+ygZzqyNI2N9Or7hk5e
a/rpCCsXz1iGdAJ+GJHYgSGR4hbew9BQ3ooTB3690Gkvjiy+aS40wVYtMKBXpyScLy0gPp4aGNkq
Cr1K2eaQ0bWMUSNddAXdqZXve4e+koRXt16PgWtnhJPVz0ePnei7PrQarLh5Gv9QLJaCs+ls4lN6
/OLS9emmdIXBV8LvwE+eGO8UUu5bOWbnUzNrdIbOUDARMNQ7G2MEnTox8wAdJEH6VPUCWmCmdhuF
JAo+oR8R/BZWuCOgNi8jHKYxsqUTLxy966KhlCyA1GQIig2SFnrdd5oXUR0k5FE7izg6QWU67Tlf
PBJuqRtxvvOJau17vINs7ta+WFoI5jtWstZPDU0bFHglsIycM3dufe6jQb739hBFTekNVeyI9SkU
wB9zWenB7pSNgYXYR+a2fVFjk0EnkABaVhJfGi/PAduuaB03jmuAPkgwh1pj65/4S1pFeZl58c54
OH1JiVeAyiQ6ymzH3hs+0Zao8YYc3N/x+o5Z9J2EuZZrnteIiYwqPcl6Mk8Jl0HamfV/nLjv0nFQ
g+lS8Yjjsog9znffuE7idLyt2cjBrtTDgclICdcWASRjilQuKKQiytgPJaf1vRxB4qeCgsXI20/Y
Nq57hXhVjTu1mkHvfNG4zVs/vHb8G0Zk7kHlOuCZzIFVSrBnbtbfa1EoR9o6Jf64JO202ho1mVx3
Ot5wEqA+3BU5O69j64egdsbjhSe4ce+8sCFAZBUkluc8L2L0rMPOfUCokUgvrK9li5sdrojW6YZD
tUUQYEQLolUc+ZKdB5EqTf0GCocnoaOQc1YgitzQCVoBWsg68YSom8NTODikYvyKpcoskRr8d+KT
Ik6Q6zVHGTnJGPKUspmDs+T51g4FnXV6Gfpt3W/P9lfTIQ5CjrOyDVAevjvR1eU4bbktC8dYdTr8
NLPwzZAlEip50AcyPZabFi5Qj4buX6eOg1pZJcz7edW1o4ayrAfLTQ9XyOiNuKPMiIIWPbz+dkVN
6W+C/lB8g/S8HEfrBdShYfquAeyzsKmABU/ND0c9Ev6yoVEYbLWcedc1nY82Cj6wMbLnRjDcnQBy
CUwSxTSRCNAAhaeEeNkX2G2ARWpcSmptdEwIoQRYw5aYThUt//GQrPZiezJJIxwOkrX7TAX5Apyi
wDUQy01+75P++YV09+Cnq90zBlD1S4ySTfZ9fMPO6HWwgzMy0PTJ6elhpbuLHvV1wQKRh4u5KnXk
sXAn9EzF0jNzTiD+IMn00o33V5gYBBk1M+me56Y7IUzmtoFvw7OoxcJZm1u42EMONxO2cBR4F/Zz
g9pNA24hsFwqpnPulSNGS47VRmCSEdKBtZ/oXQvO69x4cxwLTNCvht4S8ljIrTMLQ4eSUAuCCgUu
eLUhsZMi1CZbC/QZoQHe3jTVL/+lcaOi3GYXVRkmX9se7GBrHHz3+UIlaiR/7B5GKadZW6DzPkYf
Si4JrcBDFnfyWdrlhwqrgq5ziETZUdcLkXZ45IE6KLbw40vV8RYReC5cKHKKcm/tujECYtb+g01E
lUYyeG5RfIfQtoE2eP/JsBlSBzxSAO8E1zNJe5jKXqOqmsqGzRKUAdm7OlpdlPIPnlc+DVp6cDRM
jHv82xSP2bsREkmHJF3kddyOJINeUAwlNcOrNXtKJjo+xsNGoon74tSvkyMbNYcQrc56Pi/37rdL
3zbC4FLqw9iKsUcCd+FBND2tQsMR1+lq4C8mm/q4LKPRRv0NWlLNo8JEUUjHJziOGZEoFEvFfM3O
mD7Nf7a+DOtqx1RsGO66K7u1bMueZG6H8rh7kq0ve2TQryZ0lSsO8oH5jOBkICWdsxDu6BuV0fUr
Xi41KwAK9kBVi33xX5+Yatg5zkSTZu4Ee8BIMn5RU5k7pxlJlzX1j5KjBvlMZbii4yEvCvQe82YC
wyYYBM4eQsIiSxlXqIHjudlcNyVEAGnfw9ZPOqahQOtDeDOzsNhFLEItCd6vRenjzgZc9RM1xEdK
BHhq5gmEO6gLDgLupkJuFdyp46bak9hv+x7wJxuc/RQ5CY3BcpC7Y4LrhnIz4Y0kgxDV+ZYndFhD
/ach4C9sKqg8meZLuEphQwppFs88z7JARKvr513jvctQo61GhNAkKYpyIWFWuTSqsMW+UzvGW+QR
W2jwuDML5Ul+FPcTBWj70tg8JP3/RqjaMX8QTHtxR8pIvea+bGTGeB67+5hA5r8ZtSQfxE9iPWBM
+e6hWaj7YGMiadMt6VoFXR5d5LGIYdWosK7urff4rLZBA8vjTJn3X2Aw2zlhrVP+4Al8z0REuX7o
dDNZj60pfH5isE6GaXo3czP0ZyCHOEuALHOK6QQOCH6p1tyMyZg3NdxFzRnIxXS2PE8XjdZdoGcG
Rtm/7HfP2Krn+AdrR2TtRqYTYqDKiLVchT6em/WwaEYeOYOGPYxjvSwVUdbE01LOAQ78KnEFHmK5
/M9vDOgFREtOpSoQDSKoQwuY7aYdl+a5zKn0mjkc1YkB4QHUNNGIHs5gQ1s/a+xuW05TtQINo8fa
P6Sdk/Vvs2jpPOVN1KZ01ZpDAgOVyrB4SfgAONCli0WfERsmcjxrgRX2YCQIBlnRxVFrdlj52y08
+OPeKFHoT/LqdkCmIap87jshp+zaes0mj+NRBUZyOqwPgqSWqeXE6eYIS0YFjaKxfmsqOQLolVuJ
Elgsp54SP+mpVAd5ETrcME9ePpNH8/anpvfTKR0jurIVP1iLwCk76hD4+mfF1Zay9+O2qH/q6fCB
YwTMOJACPQ+kT7qj9nHx/pHs/6a1EALZ4bjqtdfW5TMaHxz9r1i3qNY5DzEDK16qDgpHVQFIfL7N
LxqIWm9D/zFlzdCFbuSgRZzDf7Rc8PvanVdsMy8btFZ/s1ofzLN/mPiITmB2b/Wxx6Rra+oAl1Qi
4D7eps2TcRM6AUhhNJlgv/3d1uHM2ag2M7H8WI12K8vlV786yX3Pe1V/QNByVtDSNE1zTlLqkY6z
pm+VW8DGEtT43s/J0pXbxsCPjuXdLmE2qLDvx1/jLEia5zjvXJj6phaW0vAnpgMwQL6u2hF4KnT3
ubDUm11x0Bv/fZDq+It0TL+DvFgp/WexjKkb6H9pKp+03tYG7OwJ99fv4QCLKVeEehGckggTIPhv
SNcSvgIsfKM4V2jaEkmGjDcD/v1ebHaktE5FDf9JyPye8dP1gKu8bx4bXjklRIY2FT2pjewtSudD
aQHL5kwh4A97M4KOo4UjaLLbhY9IgYgESmr6/JqGX7+EFxZK69lSEFF+7FoOw+PsW0rYnLWJwYAn
xQcbo4uCp2QDnBZdYgluGwM629e/l93vU/lUmmi4uGqvILfLDG14ZKlSzfZ1ijSU9W8UJSCzhJH6
bcJWk23L7rFY6JPV4rRcMRBDk2Gv/h+k+D69q/k02RHNYjTgj/pQ7Sb/+13FD/kIQHnKnz/V1Cxb
cy+pR5IOszaCh7g4daVAa6p8VFw74gnXNfk8bSJr20PIw6vJlKGH17lWUhrV3ELUTkEtenZ9mHkv
Slnvhi0rnoejtQpjc6cKD3Y+4gUpU5lgEYPptX5IvIONKqPJa4piEHYlXbLoRMPFvFD7XUzoipB4
3Q9M4f7kXFomZJnC3Ev33tqbZ11EmEW47rCoZNdS1aaQm0LYCKEFg9SSNhJdM1n64ZxegOSj+Qr7
qdq7lal8ojtEbil6SCfuomdkoMCjCPUck1ze87ZuJDEeZ0rljq+1DLX5JysaCgrkw6mgCRgSvv/m
5R5KjrZ0HQUvYA5HbhnQ3xcZoyjvED9Pvz3kO4Sx+uc0VrsApB8KugMMS+vplKWqNyq0OgQ4YCxf
jd41mSnWitBfZ3ySAXU4Umhw9cnOALOIus6dCFSu7SPduAoOHzM5+ouIvXyFmFjE/YuxUycnSECf
1nVQA+XBkC5/24eQZ2pFkp+KBn31v4mFQUGO3RwZ3BVdKBgCc7U/8FPp2nlCgmzRuWY+XI1IwYjk
nRWukhIMoArVqKid1+urHSF6TLfiFqIFTeECfEFVaI2CefnOx/AfWa0lpemF/J4D4lun60ZgYqoe
IjfcS5Fe07igI/RX5IscGnJFV9Qwz+EJ1/ylEftnZhkIabeJIHaztrHRr0J6k3ytj722tkJC4Pqn
VJqbXNrKm1QrRW4k2nFZOIlngUd9BN7TgIYpP/AqlrUGVpzE2pzcr9GR8ceMK7FNOER5gNzQmjvJ
aqspudcj5Nb6PuOSrU6f/j5cyXlv2s7yet4kBDi7yQJoETft+Potz4XvXpuHU3TH4Z9DSmacluB1
7MpcjAdUtchTOKqZxt9imgVIw3oB8HNslsTbbXoA22ruezjpekEAbB4KxXHq3pFXF8O7Wpl9XOKV
9nhIDI8PA1MNVbZpo2wY410cwJ/n9LlD921ZrnTBBR5XYNWhOaRBTi4qYvXGO5CY8+LfzrGvtESI
iexfIDzrKR3NAy+2/taMpMAv+STSyf5cVt0WdEeJMidQigz+4USrbF4Zocg4RfF4BQM7t+KyA3P8
4yYaINvSeyJ2/CM+3uEmM/YLW0ZVZrSvyKAlFgpDlrhNM2mZ5iQQVhl8zg3YEJ3VizNpFZ7eMABR
EmUG6v76PnB/xQsRhk+1s53mAJ14ihQK5Z973sPlos83+ymAE3eNAaGXg8U49A3T0s6H79o7pV30
T87hygdLU3JDxETkrNwHvp5J5lWtvZAvdvs/AHYf2IDEpaeM34K8ER5FCqfZ8PzG60CxwkGJXWAW
q3+NYA8ZpfgigGz0JeCv2NzxpCmJenL5ROH7HxTkEaOmtIkkdOrRsR/VwE+6wJiuFTtK5w4P8wx0
ba6eKq0eodkrqede9886EIPwEHwusxxOlrlZQ5MPdkc1bPXKZ9TbBFZRBUetTQWkF4lXzAtBh+xv
wj+1giTGJDI2Yshzv5YecV5nwVgQZw8W1RUEz/FGhpIKvWYz2lDq+9J5tLR1P5ey2cdh7zojZTH3
I29G7CT1v0XlkHfsy4L1Nbn7hgmcfwOQj1AqeudmXm1MNEB1ILtU5gZCrNoaecKP97CRlVycyZ9a
1kGopVVJXeHKG/fxbPAUooBvv0rkGVJDdijyyK2zBh9XO725jGwMpuMXp8/bWO8zjXH8Lgc0btpv
MHcTG9yBRAwRVk3kw+0tJ84bMWr/XWTKoEhrBHYJg7AUUDQ8rTpZ8OYuiNMnyWWpvGXy/lgeS1KI
f090ss4cDpu3LfK0GMETOH5kecVS+bruVTepuL44kUSGw6rKMyKLtrJYr5e5Qhs0SWGlwVzL6kOj
/EFECD3ct1jTzOuS4J4AYNwAUCobBcwFVrCmefsSRxqd4PVCwkkUTnOkDsSJxJ0Yf7ptFfyoY27A
cguOl1Mk4lRK+rQaHaqXrv+fDV61a7x/lFjmS716CuSVtXolW5MEOXevakBuecfFMi0R2pd0dh4t
lYfLinhWaAYNoMo9eWXiG73r67FHe4Ad/h/8Um6EnayPy4YSYsWec4zt2z8zgcdFrZnOb+iZV66z
7XkL+iRRAKDz9FramyDbwVsccj01kMFuJl2YjOaM1mh7EHdl1Ro6ynoCWQqXSEzHcQOn8Wn0Gfaj
ZO17gOEavhW1tnpzmYEeQu7F5ZwMKAlK24VStx/fn8jBtnvFscBp/midvIlmw8ngLcpgY+O+rmj1
GBtDaqFJcMWeJJ/0TYNNsQA3RpPLHhLrxjb818OBzXIdyUzQ3oZ7bDbJocAqH6mjiheopkbWwqNh
t10rHLVOE2X2XviAOPwMEK1X4vuNqjBImy4sdto1l9oF27lAtsGRFEyIjdtV+5NMea/oRF0ZCr32
wt0evsOSBUV+Elov6mHJoejyvC0evQce2RFCEWKT+dBBNgxKe/aLhHzPqJnu0urCV5h+YAPVbUMI
81N0w3kB4DCD02RrEWmcIEbBklvqXwvvRs4ItqHyHjDBw3RJlf3yqZnCDpin5AgXUNjI4Rm3AXxV
PAhjNAuJWEFEsCQgjIRTG9raErc1D+93c8u+D5FJvC/wq+NBKB38iLcoRY3aaSUFMcgZWI+wb7vZ
j1W/TeZSO76Cj4qsaaYkK9Dd7NZ7xWpNIE9ViL8ZLH3MneoVKF56Kluq9cekCqtjxXknNYmhPRzn
7Ni+EMfZfyVfN79qqujHV1iJinyoPaAjgEQjaTEjg9AOGt6Avq3KjehIb1m6U8UYPadiQWp8nAjq
zYpeu097C1/SXps8JzNmKzmZVUQn5BAgNRAQyWMntL/qP0w3wuu4lzqOl2ZQu4/mXCvq85NXnrBi
WZDwDF3jtFxga71XimnjjhdeqGBRUbdyZwtQsDjKSUaPm4EvONF8DqoQVbmWuWaZFw9AFvrAbajr
OLcrOJUM0mxQZHuMcsYWAwv9gsZEuQPdmVtXENQlePTNEsCy4bfuekx0V9QIX8uPimLs1Vn+AlXB
Yzdk+7lQZnOT3wfP1YjNJAE5vrLPlDXSasdsMvKs9D19aUQwRVUlDH/PIoE8V3m2k0KmG0ccQjod
zMJdN5OtjomE8BHEctFU66icW19dvxnOPsfFw7ojbgii6E+Tgm2F2CcQP2nnqOXPKAYrT/65PX6d
FMCs7sVpiWT8/zCdE0UnX/yHwbjaZwCsbNDGt5H92IIp0vvG2H8Ut2PjE4zXkTU6Z0aO8d7r7k2R
mhpCP/ZhtLwGmBw4SbGRPLQwIRqyDNsrhI1BEVlNcAsOFT9g3lpweLQERSTgENuZysKH0DOd/gGA
1IK1vckPxlcpnolSjAr478OtYqdZX/uAsITaMMJohC5aMzuQuO/y3HEuyVRvlxpCHZ61ZQI3HqLh
khNCpFzmtW8uPVd3q6ienCgjeGrH6MJQdUcdBMfuyDEr1srMZAtsXH86LXQIJB5+1+q9aAufrck6
x8uKyteP22+JWExPv3B248p78FPdFXyHB4ybMShofK9wtfhKJNYqxBKxS8iyMC3sfWnoxTsyQNeC
Esy+2tc0YmLS+cBO8ocH/dMnaK9HOS2NeznxvPCc4nhWWOXNDDcYMcRTJljF+11aQDVJ/W5xJiTV
aqC7nY6Wl1P1EDRhY1b2MIMoPpxcpMf5ncUVgG7DNbWB7XBSg6Ap846lCR7I9j63K/adK5pUnDC7
c9xnt5eZFP/glz5eSrhHR0AYK3cO6o5JphwAvG3DIWnG3jfTxr5frQIranHqu+ehVhaaNuekgybG
/0oagvN3Pj1v8Ig6sTT3rqdXHtsdrFxrLDnW8vcdRsFfIXA3O2fq3Y2MWHyFSEAN7WPR0jYORFQn
o+93KZZwCxDjvcwBZkUuc43KwqdN1jojg9MujzyR69OTqVsHPTG9w21QsvsIMmqAf+WL3osmOq1i
g9pjk69Ve7ozeVCwwFFqt3nB+Yo3QZOOgsPAWeoWzT7AY6MrmBtpjssdqFwVUBG3Qpkup7nhKIFb
eMIfn7maCrr9ZDJDXlynWNIuN/mMxmTfcAKgggwFkkmh0yQBgX5AZsazOJA8wiScRDZPxmRpKJrf
6kxJZ/LeJQdayUNNuJEnp3cj7OzeoDSvSlexmquV5a//QJYWRTECVnTbUGelfHQBn+m7wahNKiUt
d0YRFPrurkPeVi1b5oI3eSpuigWDkSDwRSbxJLh+oWA8rtiRNm3T+EEzoHfI8jfiU82YYD96V4QY
6hm1D4GzBxXSY1E172HjZ5wPKLttx4HnjpjyKyhzO7XprMvYCV5uie6/zNvJ+DHRLJzJf8UM+zzk
Xmrrl1tFg3setrrvv6WIrZddiuSoTsxUYKN4ROLc7zUWL1Q+7hxIuiNAiBVRvLnHmkGE4tFvblvy
OQcn+LNuUInc9/IfvJbNpnwe4pXINzC9n6VrTQrXvUQvlpAIVWeb9YcO2yHTkQSRKZSU+Magw/ck
N8A0sIhBpMNmmRUdIMEqBtFB36ZoEzhBsD93o2V6gHp/cvkNvRtT3ljROUm230MQS38btT3+alsI
3VcUpleM5NAKI1Zvu+NthYquhW28EWhB/SFxNznaPXeQ/TiXyEeiBfRksZkVXiWS60UtkOwFK523
W9D+KyLFLmqiF6CTkdKoQAS+e5OziPKIUCVBYtojIqAXx7xcew5JJNlXkvPMOFUTNJF3mHI1288P
XPAb59nrlMOzVJR7LNCw3K3dyicvqdLY4SE/l5NBmWL3mx1Lx61ZK0kDbl66bUXCJD7Ulk2fLeiP
KfVqv82MCzaQxNqZtel1uMIxA8CdxZNvUZ2gIR5JNivgMbkZLuHnfTUv+43yZK0KtfYTWs78eSKV
C4tihrlM7AbhGLa7aihDsw8kvhVLc32M9EMflGkkL+WzelAG1BCOEZx331M2+LkBQ9ZFe3Gqv8r2
iRPP1jaMHDqnp9On4FK/z1QqylfNMNTdo5H/bRSX7HRsPiMInqn+JegBPkJVYhS884VnLK7yLEYj
wROYcBRPbTj/HMoAJXticcOIvuqTs0xwhTxbkMO58o0wXnkmi5l2naImoRktpUfesksLXcaw0tQ1
qi14Z1VHhj/5sedUASnhormWuE7kkM5s/tET0jssFGMmiSoEJj5u+A1lZPgRVX734gn2d1X+dNDf
r3mJJRw8x/PszwNqbOnp81fV+LbVdw0YWdMJhYCdQfakvjyCCnwO6qPFzYZazUDWBNBihDct1emk
yTqGNi0KsfjalAKZPPcvXKxFu+lfwjG8eZhaFL4Hv8YQ148x42/vr18Qcme/sylaqnwYDsXXXkUh
SOF3uVG+jLy2JO5B3d1CrLEe9lK7WpMksw5STegrwCGZNprP6IbiLPdSHnE1RIRWdfhahDIpThvd
V5OwJLkb/Nk1rduVHQ0MkkaWwff/KKAs0tDAlQYole56tttBOSsh+h5z0ZTvlIHg2bfBbfqUIy4W
faMBWfXu9xa3QOTCipsIhmW+qrKpSTpqXkJvkd7ebLbjPN7efR4mYdHGXz6Xz1GPaDPKjXtHnK+D
Y/oWtWrwVgjgcyrv57A6o4k3bE2h0tdYpHvcrkgmG9mT0WSwPI+29NxmC8lLkYSFo4/Kp3dh7gwI
kikQdQTV64opUlC5FBigxJD0DX6D/Yzfk8WeY6vw59JNjpyI2O8YLa7mT2nd/bKBo8VUK2DD9Qfe
JLpjDQsI71yGfKjDcKVRIhPx/DfoInjeE4YR8y2tVT5tcVwKNl/PTcsGabLx7IjyigBvtd9NVgDM
bfzVN5LTDtoQFLqcA1t8eeXVYYPL3bPyi6F1X67G80GSj0EYfn+ah0fvmrNV76ZrUFLN/V8q8hSN
E2FgGZV42mA1hFt/QqakxYGqWk39A3XDzYKpEBp3nh6+T13dWqgh+ZlM2U3xmHzzOSdi29/O2ECu
oewgapxjKRAUqJqP0D2xTueR7twx6UrqKefNSTvhFQf4HKTihyRPOa+s++pPOmw6CjQ9XBHoaJ45
2i++QvXAyEJz1w77b+GpswsdAZqHWGew7bhDjbQxKU0zmEgEfgM6DIVglqojfsQ4Y8SkyWYJFPP3
IIRZLBtFsMQK8IL4JMmpyutJ12YWa6bS+zFkxYgZBC3zuzk07WvtAG7nMHda7osjuAUcr0SQnztV
9qeZFsUwHrpmd2NfoMd/EHB0Q58uaIuiDLCs/VydRmKuxLsHXrC4bnNjiHv1BRNxOShnsWl0vpEU
kxzGhCRsdb1Nrw0vY6e3WXFX2D92t1Z917WVNPxNYeXUInuD6glpiQtJrFyOlHMsAp64P29LWS7U
xRFl8WrhdN+pPLXqb2eaqump/UjBedbScpk6xFPdLMN+kmdAHXAakGpgwGjraRDHdR9As/CaGkcq
pxETae3AYe1dCQGL4r0MQsCeyGhg1Pbw5cwQGvE5mpCLlAV8BgyulecjS4kWzTB9wjGfrfwV+3l3
KAk7rNbR3aO0y52gM19XOklj5cXcOerLaH9vkmqXmfgyp2rzNh0PkgUwmL7XfsAo5t1AXDqj7ogt
Qd/bT9+xoLc0MD8IlnQnIuHxtHc6Kn8empAMXcL/uUITjhEpTOL1WSNn4HVDiXeQ3yGmos2CRrQU
UG2SiK81fZyNMsNpw+HSJTUrEtR88lK/z7kkRxTqFyJRzqmk/7n20fkwfZfpkLkVvn0WnFHQKr9H
TDxHFz1sM1pGiDYm6jSf/vwxhIg/QOBadoRBnOmK70J6WJy8nGfQnSdge14iLnTysyE7WBD931B9
KJFEErGyJtvTmW30QDTXVwPw6hJCT33a/9Ax+hzN0mIMZQjwd1Nn8V3IHlZrhtkxD4Z0+vjiKjJB
OTBiu/if3zZ/upgaEW8boX2/eB1SeNhzoMWQ9ndUd6yMej3GIUZSgbl2hELe1COcDBzFUfkJUwrL
oVUMZC2rK+3Y75bSL7VdofENQbr9wc/tcHkmIJs4rpS73IYOXwZf4kI9Iku2qWWwvx4OIWODO+l7
p1W9B75tEVAVgZeAO7GQlClwbmtY4wgn8TpQM8meuImDC2SOU6dOrxYJXepPb/pjPVAg/dabN/n8
cpwuIwlMdRH4mNk5XPozQL8V59CW4fH/jk9ycQ/ttrzh3us3PsrTyFsjZXYryKCFNPSPXOUSXvXz
jvbij8AAIgyb4ZQYb9EbqPo8Awjw2RP1nEnwMOMyKoUmFO+ZLjbrdJrEgM+vrQ7OKNbnOEZ5Kiuu
dhel9Z8KbUeLaZEsBck8d7bHxwwmiFpV2tBh8j4Euxp2hKrS0oD+yCn7Hzu74Z2lYrjx223OtLmq
gORj6J8i0MLVeSmcOAzeXUV1ZFjMWue5bKNOprFATU69dSIbAVRl4ZB1FM255iPG55dQ1QeKZzDR
pdk6MXNjUhx7OBaLu20Kz/0Grs6e3TyvEFeCAuGLUZINHxH4PkTI0EqfUIJLXtJIMdGndjwlCDLC
GGjtxZvyxuFMD3nf8xSeYAUjyOlnBvJppnEvTkJU652FEbvX88w/KFRWTHCQcM5MQURj2kngUulI
pNy43rbGwhehWOU00qykfgFV67IEEpDYWEr4CisaYzYHIlD+9AmP5GiQxpjYZ9/E1VQAtqqbl6WP
fS83Ic4yKIAdRaX1FbLsUsHpaN7+HJetWN+89+R23JnesEfh/2B4j5jmEZ/oyJk+7ZpVMdGswFS0
Xech1KtOF22fFGKOVvumRzNu3zdu5ZcoyJOP207hnT1+kQzGHr6t5WQsdaNDNuYDvzx87tbggYvF
X8oZyIWMG5ZnTF+DkfqF6OnH1GQIcRc7X14HZXz+OvoLLu0vyGtnfmZN1OMBTtb8kNL4LFaU+4EE
a3/tnDsJldY8I8GTrnSD/jSF6a0RKXEj1J4n7DEt6TMiwP1AcCvONdVTsdJkecTSoVjo6q/w9ocV
yxvdoVQuTVonsJPpEMPgVr5mdExEzuG6SR1/2K1ZE9nTpDn/LhhSe34xDFd6+FxYrP3b4cA9tTvP
qBL078OBnYWB0M2d/Mi5pFbNeek1dGBjaZ0oEgQn423hJ/HNm9jvIdW3NRF59BhPU1KAhhrfXS9A
QfhRWImONRzGd7jz4YllT2rrXXxebCWnfwoiBQ0B7qajzbnOWPvh6W4GW1EQAI+b5dXRbhSEYGZV
W73+CBfimZW8khQtVL9h5kVGLkCOBtesm80emsyDV85cw7HBAmyjpTHn9EkG3sXmqsI/GYovVYyF
3KJkZlEBjAujZjqOWfeGB8a9dcwmt45NSaz76njGF7jDWNQCHwGnmazInVJ8cZZaiJxLCZJGFufd
DaTuS6eLfSPUgcU4B+q6JjhTyYSCAvrRda5zET1aP5xYXbtBxC3hD7BaYHhzQAUtdBvCFfEtYs81
YBzPtGl1dgo++9gE6hDFc7OjLKhQ6q1+ohFxMkxv7GRn3bkFOcz17x3WlWjMPJCS4NcypU1LlwuB
S31Z6tO2swFbpHDjDDZEcFpHWrF00ZHF3Yd95EDfE9lp5O8KtE5yZS8dWWyUDoxNhkzO0ENqHShN
DBlmaMdKqYfZZbKGsOnx61BQvibHQ41Sjoydg1jQt74E2UX7b3n9z/hU19rjp3+pdluYIX0OV0yV
OIGRz7VTt3Vm53zGTzgCIAg3B9RQcn+ArGwzRu5kkOhCxDuFDhetr14tBAsNlIjFBiV1YVM6N7rQ
UWFX2mhgZVWL80mmxA9C+Vy9yvyGNvRtmc9uAx48j1bn7aiz1NpEZst/Qg+0DHCMsntnsDeAwkbT
JGwJwxZadWQ9vDx6C1L/OeOh/NsKH/sin0s7DnQZoRjcsfN21ylgRilSqx9r9OwQuGGxpiIs+4zC
kV8uA3zc26a9L5G0qDJLSV+l9zDeG9MNMPeSjTVT1SKLZWDggMkTp6iizT4pwwFDs0SbPdlSSwex
LqOwRG/fvT7eaGJpdMXDsT4AOcRSxJtB9grDQMCHq5SMyzqUTaSV6+gXsgkBYY1ggUKIxVwrPGB5
+nfILI2F0umS2BBPvYOtk/JaznVHp2NNjGWYGxK3ZbFqkL+k1CZ4UOs9p6SSpdilesgLP9yrg7m/
qs2G344U2B2CIRL5ImcDJgEwRE++If7c9fjnSx95Rq6BUmRFkVHGy7wzD0TGU6BKqaJFJmkLK0bH
/WeVIio8CQMvGKTiSN+S71U5iSq5ZzxwlVPz2ykCVRNLWPnvQ9ty0gXHXOcgEvMyCHXafSf6/HqZ
KhtIjkd/zyoSNbvYvWNhyLMOo5FU97tZ9vOWa7AhUtgguIaaS8C2yOESaZuCcUnvt24ZCcLtAsUT
mUxQ6t6qpPRf0I3htXT7ykS/eBJSU7ZxYqW9m4OzB79i+DX0rcsTHRvNmSGuSm87knA+T8042lub
FGBKLc8873Hx9NeUMLucFsb4XUwa5wljm/bSGeV/79SxxiYr8EtVpNlFje+TzlHdpB8Ruma+5E7b
RB0TzN4Tsptn2HFHKNyHitADUYM8f2w9/aKmdAgjF9bajH4tK6fWIWxludo/5z2HfB2GByeqo6fx
OtDSSBv5AFLQr8G3Tk5dsIhw4/7VqgeQHTldvkldHD3yy6082TyQqWcT/GgzCp3jSEJpOGUzM+5J
XJC8A9UPiLBe5ubiue1wiyZIIrbB0Zx9kHlNp8sEgvq+iz5qjbeE1chLHOrcy++uN8rUcba1uxWJ
xTdrfzVVU5hBoXUeidZzi/xgUjkx6M2mpf3JyXtFX6dpY+IbS4OaIVQwNT7slB/LyNldCQwQQ4OR
mceTKMB3RQUE6CpSWm/JWMSZfQ6SykNNr76DceyJcDSfZS+WS/21aXEWCF0m+wcVlmAB9YSFElwH
qeRDG9yDHyp2YXbBp3+wE3Nu6FTnDPjny16Gzo0GWY/zfdb8wwP9mKSUBh/bC3+o4az0huZkdTOi
KI8cJPKoa09QiSII+4s981tlHHzkgLX+oJJk8fvZ/ta08BPeKPvOyusZMS6L0fjqrI7dqRqAX0/g
n/lmspDo/KvP9kWvSgb94e554tLE0wtceIKSKI7RldU+m393Fn47oTiVyapX6TRHdWyxrTl73H1P
GlGyk0loqwU5wbPltjJdduZ0QXyCcDkTMQpNtsXx1nCmwbDIiH1GiKIDpAo1ZDo23CTeKygpPMAs
sSWQ1z8A/Y2yHGnI90b3PGC2zIROvKw0UnWvef0ffk9keZZ8Xe0e3UgGUAU3bCOfBN1dsJznsnO6
FpzkEG1VUqFkvqj+tI1c9YLvLCWQ13E/cKwE3mCYYU7HsmvShBR6vo70rPH1XSl8ggYJbX5ETv2U
rJAntEH1swm1EVFu3IRt9VvEzKy75b7gszqCEdr+IFuFHWr6fxSbHseI4p2AqKQgNppCQImM09oy
K+ftHXhr2HgsXmXRCHov6PPC9VQ3GYQJEawz31kET2xLyG7h5KHUzW4KPgVc30/Ap1URaNGLX1EN
AREsQSceWESjWSPvZPu9oNxW9lZKCeru5b77L4aQoezLQzoX+0ZLMAFCwVjTJGyvluEHwhXvVyBz
qdLzeHgzw25+pg1scWDBFxVqWg3ls3TIEb/p94sA2BNbrP7n87svCRCd8ZJJoZWl0cFb/DHic0x0
Op/Ce4SiiYUyJUWDaztpscBbHAApmSsgWQa6rP4ZDLG1HjKAnFU40a1RwmMMvQMhhCW+9JbvJqo5
HJEUSyabJuF4NS5fHrwIUJRbmrp7+5ESgmlfMs611xxYqk9vensDYqvBfsVSpHQfOSxAOYYhCImK
czP9gh2bfZSIMftWJ49RpkVR54pZdC0go44aYNS1cAqOzE+Bm0JyFjJMX6K5rclgaYrELuP/c0A/
IPdMJOn0upcbfxqs/7J5ThD45Cii+Vdgzz5rPv4aMAgTgbKAM4CMh7rZWIHOmcjMA0tfBjReFuko
eRlO1HY5egkcXX/LhEZbzc/G1dRwGqUZVtHhIo58LMqC/9ZOhALSigMBhdjRa7huSrkd39WGs4WN
652hXWme/+0abU+V+AH0OtZ+ve1Gb40p3xfT6ei2fgazR2HKpMDevpntYJ0Rnb4tpps4/jNudjik
L1wXEFCqicGDeA14mBXMSkH+8ilEVFWIVxPPkQAZ8FQmF9DPVr+9uoh1YLtghVOn8AGlx4xhhIuB
W+dFOVy09GFfn+jVmokTBwWQv/Z9edOrg3luzkoD4kSNaQU+i3iouB+DHkDoEv36aik9QLcvEp/o
6dVmZ26pAXqRyeGfDEe4OYfn++kiZiDESy7Fk0iKe2veH5JXX1YvbX0g+fu+GGSYdwmbWYcGCKKA
AKqnMEbE1o/pMthb0nTvluAfzcHUX5//ZFpc99Ter8dhcqIPhQAdoT5bVib1ZzAs2DOTH/F+EBtc
ia3bLSURod9Gt9UNjvKTWtP9FKcm7JItc+th54fQaOqEtb3jIfBF0EXLe2YKGAxn1GNrK5H3EbHX
A/4/ABwVuwQIvmX+tK9y4BAdMDUF3KN/RmcaSZx88jgapHbnUcJe1EC/DwUEcIocSzpm82OLTgu1
40EjW/c4QGsWIFOG2aS/CKRWsW2S92WoORRW/4aqn3+UN00gDmMYSyxLh1TSDvvuRniM4oj+NN0V
H2X44noTMWUaF+6P7J5kxqieOP9QUFiqcuYVnrLgmRsLSmdx0At+UG2sYgwSRJJsYqwMlX+/+CcL
iySSze3YvwMz6wX2KBYx10jMSQhm2rmdJzRsGj8c9QxnRymDcbLuY6/LX1R5vLPslI8KTIH0qjX1
dJZSvXqoPS8eMh/xgc5X4EyR+gCQGsayhgnsopTxrd2SSzm6JugJzkmHXrwVB1MUomTWTRW561DO
Q6dMVGG/a+h8qC4jGkczpPrZn4By05k1C86vEzMmxWEkRS4Xs6SyOWbx3Atx9Wd79WLhCn5+6Ruh
/LVa2zV6fTGQ96Ulya7qxJII7mRnledVfmGdfnxRnWSZq0TM3i91s9XEQ8R8H15xZ26jN31DVkfk
VGic8Bw1WF43BbORqbijVJAs6t2pf8GlrkJ3vrg29mmHSpgOq/E3pzgYlzC/BFe88vQhzvgmWJXw
04Dsq3dFBROGdPpgAYvISCWU/GyfP6n9qQe5dTDG8v2rgQ4VsbWbSBNfMjwM8y8rdRW+IxLxD1AP
OFjJa1kBSzTC6XzW/zPyglW5+9ldVo+Ch/88EVfR9HISDjML8JURZ8neVk0wBrDGfabY7yquvhB4
aygnOBQawfsJiNQfROy/HSHOAFXMiBJFdethJUvNOeKgibmOdguqYRqKTKqRVk6wTqMpzkJ+Hv1D
gLhCToKixlmSfoWZj6lGRsSfh6IhF4bXbUTr9oAd3xcK3N/D71004+xGFaTQBColo00rt9wWuS62
mi0XfdB5l8lhHrNOKQVGylghJgwNu/HEnTlxjCcBdjECezpAELtI9ZxUmuVvb6fY45c9l2xALM5B
iE5ge/5rTgUj8j/0dWWyJfYghxKoPvyzN+hrKq2i7KHueTHH8YovsJ7ZuX8G4vFgSnTBr7vKWCZ5
WH7B5ajz44wenh+LhwXpzUAnb0bzbTaQ93fWP49EBJ5fW/EClXi/MkBpa/R1SCJ0b77bQM/+cRF0
ALPUXoqmCm9piucoR4H27CnXaqFrJY7bQ82IQia1F2Yc4fLUL43Sx5d4pFNTPNa6ctyn7cyPVoeq
vEH63PnNV6xGbrY/jtIq2vo2qiCkqkq/adrxHTqqR0tp5BC8qs+6ywIzxFSQR8Za3SUU9u8TbH9V
kl7CWujmYzLoOmyWyx6HvVfnFOosR+Rl/fgd3T/QWZwxwJEK1YqtJoCW9pHspo+r9mnSaUu/yB+n
9x0sGv5+T43LQVe5zBdPP0j9QwbR3wcxXRf4UZYOQMasJsBOgt/xo3JA4kQfSyL/4T3HYBSlyEqv
d8QFkxypqL/5yANLBln3mzJ7deSNwkB1G0ngbo8URy76Z28aq/WO0X7OKTpJOsae8un6+thpjL1x
F/9ZndltI1M9esCOVagIqgbfDrCcdENgXi3ujLZGaICox8XTrc2Uf0hgdi92eiWt0tWoWr8iflWd
/Z0ANWndUdSP168FS0arLzPm4ZMptKTO8QXO72J2tQcjaQKy+Z5xs2+UFZ2EI5JcMHX5VBepZcgA
t5IerPKzZbshia68Fe7RWryq/fs+QTi3FctQ9fOKHwMJ7xPHTewpU0EgBR3ZP/ABzK+bPEfAqBg+
dM6Ek1KTRKHYC9Rqkd+OsDmQO5Zw/3frNPK4FmR/cyhWERCv1vOw6DXUr6x5orazvBLCAP1Ey5hd
6hA4InrgI7+ZIptubd4hGslDRzXcvOoXzDzPrAME7lyBvvmhZavlX9jz5QeqJZTuFzPVUfO9h1L+
hASrVRii9E1XNxJXG6LxhL+nfR6s8NEtvPUN2lZnukr9DvIfoE38m/jhdxhyyZy3qcLFRxeplmJA
qbGfvOqdyky/T2eD1ezEvMRfGhB3/cNpjxLyabmcU5zwjcevuXJSAyLxSAiOmYjGhjVRDeGRqVLq
G/71BYRuIuclZaPrSgxaYRI4H+Jafqir5GM+K1TobXbVr246Pc4pqjCZsWa4nttVPkHgLDFbV6ki
L2W820tIs829EsIUxkcjFFe4B22f+f3ry8vBXKd1HKSEQGRQdFlSanomcoC/PqKWXbbTvHj7s4P7
6BkOVrzLmPQEHUY/E8mI/Shj5+G6PYcH117DdogeBIiNt21oUgHL9QGD2Bc1lq9lfufpNy6i3F4A
H3ZQl6OpjE2YM0SxcXMjq7VoJJU45XjuhTdOgkr//ISkxmtgAlTL9JSntfUqWxjmQ6dZ8ZvMeS7y
t8BFvmdAHjreRYW7et/UE23pogRxM0E6WZZdTkEy7osF3VpOYLmibMgxvhS4pPzpGVcHNdZIJ+TQ
QWY+BMHcR8zW4LGWKlCqZ3NcIDxiTxhLo1wYlaUh9IzPXQ+LW7gmKDRi1LmZXFj7pXQnEgJzvGtK
WbzrwqFy0eX3cqUNng8t6e/BEo+JAafCEziBGpuGH7mGSj+A24hlzLzUvoohTucLh6g+Kn/Q7wuY
UIupulnV+JXrP+dI2XXoOBbHFH6LBTwzMm8j3JKt2ceXLRhuQSaYIIDuZyP++PtGEfkRur4K26vK
+7HGJWnYojl9vtV89t7WlD210TQYwU8nVOHRUPT2sjJXSSSAYRbaFKXUDIwJi8/KYgiOeiA28G2Y
wQrXXn1o1nS9SqrJi7jyLljqt4jz8YcycnMTTMvxvvCSWBZE2GxO7J6+Gpte845+GxvcdIqhusrV
vHz1Sh473DSWBlnl+Mkpna8t9D8xkePDuD3PDiBQnNRCkBYjT3lmI3StfBhqewyWTBSTbeDdr1Di
57syB8/nYowLg1G2kZwtsnF8TjkCX28Qd826fqRgT9y2QMUwyliayisa7U+upDqXZvKPBUTO5bKP
sklNFBUupEESNGAEGH6Ok2NIXdPsxNXw3zPQKRkqxvnTXXIOQY61m3tqCCnMxyywBdQCb4GJr3fD
ikbbSOgUi7soRRVFM0sAAeC+ugIrmA45flQ8CW1TvblXlXagkP+19qtJOJ5hRP4jPKOH3v2OpB+L
4PsL9ZI+aeW5SLvFfkVruJmCHT+yjzCEEdIDHhBWvvoVAL4X0tY/Tm2xkjwKZY38TXNr1AreOof2
MZdpwQmIe8otEPETV3b3S0qiefM4JFIuDuTwK21S7BCI4a2p90jXaX5Dbwad3lDoHtW75nBxprCV
hdv7tnVB/stU57KCZqVEEkYwkFwai2eTXNoMVSfY2Ysu5Hi+1qLUBXVkL2VkBaHE8B9h92E1d5/w
Sun/z4YpQU2gKeR9lBckkAoe3wYHt/MtMpx/FNVF8FmIiBIQgQfsR2aUyA3GMlisd+8Up7rZDWFY
rrd9m3z6Z/C28dp9tI3i4gzil6JIZl0h79yIRTGfkEdas/0M2vCpE2DR4o8rm4h9rFzCM/ZH77TT
xj6/+M5FcrX+k5gOg/8mZ/IlgVjzf1Zr5smijSHoRlSBf37sQNZ1QZUepxvwocbslCV/NS0B5SoJ
0tHmhSoE9/qgUXSjQMdCwE5apHbMcOIxjJ0qhOh4FQQJ3W4U61cVlOsrpyjvKp0dp4I94WVBJSOJ
lh0vf9VejNbr5uaCQ015LFdykrwwHHrfpRMpsBg6lZwGfZ4jhle62xcH2baElf5iwokNRwARqBbX
NalmnYDcdyCw+uShkbB4OphWtHKFT9HphjeBE98YgVSWjPb/rCBnpuiUPnstxXRrKUEftYYij+Tw
ikox1FUpk4IGKobaVH6yIQtM0npuon/exK8TspZ7vNBW34Ke9JPhF6CqEw1joD3Ldk32+sZx4z/7
0RRzN0O8ryr+YT37eAETB8McR2ysPWB1SUl+P4r5D29k9bhcjN6PCR/KYS7IUHdts7Jg105xWS41
glRRrQ707W9RcvXD9BR/55zhTjrQiPMmbXS9yMOKAlvey/G4y0nt7WUpX3d1cOVkeKJyX3xo7FN7
xRT6QRKzPPdt2EXUgMvBE+fX3u7AB9OjDIQWdmDcvn/s3iGbaGIDT4BDmPY3DBybjUf7pugyMW7V
9nwfqyXu3ICgJPsinm5SuvOSv+1tfFb++dHDklgwzUV3Vr/wIAIybonH7AoJGDUH0IxdQUSPEz4X
2lErGborFGn+nrTrcBIw0nUiv/EbMX17PyYH252pRTautDKYTjDCUCgi/sjjaYfDyycb4jO81raJ
Z1zam3mI8x5LJ+0zTaRWuOy2AdXMZ74Dng/zy+3KCgbjjuCAUJR0bY3MLAKD2321OvJSRDLGGFgW
XXRzto6mFtXCVVVy99AcAOwalBcdmJhjrDax9tlp7rMp64XyXuHw0XlJNdN9wv0QLFQPtQXUESVT
4VoS+EiQRZyVglB/T+aDqYN9YfMhwMg3sU3rVKs4TqBnPgjstVDCDYjdldxNCsj8Wy9KYpnyGJdN
ioMg2jLh9hc5xSDHc+YkxgNcke11cJG1xxQd/EQDdrAcoOsau9knSDM0Eb/wFWoLhainthpif1ks
DLf37gOfXidxEfyMyeMai7jwWeo9a+IkdKeYnvel8NCKhxkSel5V1E9BPmFDSzsSgqzlBny4CqjX
YEX7hTzVMo3v/RJX4gnIeVIZ0coMuH2pUTdB9XtJcNClAWAlXQVUWTl4ikULODS3HjLRwwG4DadX
BsUELxQqj/u7rc1dISr2htqbzbIEL8XT85iAgNtxwSpCSSM5v5ZZnzMp6IX8b14syA/K5GKJ5Qoc
JtMGmp1dWGGoP41VrHclrarmvISHhwHiXLut2dh4ZlJTgHqX1iCkxoGHIPQ2iwJwbqfsfjsr7oD/
kvQT4GeehgNP5DIPfkHAddXMluxlTLUH0+4Mr03feysblxvAmE4vr/+8wkxSJMQlwhPHY/ZcG9sG
T8OAQnNpWDnit3eQajcfUuxfggq9iGLu8cdQMMQdvUqy8EBxrJHPpussf7G/Vjo2WAeZjIZLh2SP
JU1YmLwo2x5pavyUzGlnjV5c6GgmTiHXcYfLNo2DKyNtywVY2wXFdNXgGnagO7OOZba82n0DvccP
3oR0vUXK8UIbI73rkcYDrUdAA/iVYfkxmWrVahUaCSJ2x0iHBOJtNRG+BtF58IlYhlfetWlC4P5t
+VLvxDlfk/rdcZ08d99esnWo5fQm/5JqAshulTcopAHSDg7hXB9OGxkqmq+7VfJfjBED/ILiLskO
W98JB37Yt1VWlVffe/QQe9qbrghDI1sdRqUzP0GkZq7fRPWCY1rWgubvf/faY+YIGm/UPUVBefgj
b0Yaz2NbxLWxWmhRs34SBmahjA0Mx2M3ZpZVEKds7IOkcptpei0zJCBaRXq68JnQ6At994aUSRPj
Rc1tEKpBttoJuWR70o6tSHhAf+nO0EYprjhE/lvhkOEs5/eQepZi0dLeDXZE7pbLtstdeqJl5J1l
bDjZUmyajbZd72nODChkrzDxJi3mpG+gYY2W0fJe+O0nQx74qo/DggxXJBlHb70auLSZkDi0zgiw
JXArMYJQJMbu1c5CBIUPT0Eu+R1spYcVmxVY94S93njVvU2541c7+Uejr1/WuiZQrIr55n9Z6ghX
oZLV5vGElwoJShyz3fBjnOTS7oTnkv9Ip8byfsACsj74Ul7Q8Hbtkt/5/GVVjdhA1a4RWJtSFm7H
EN2Ns6wAfF/s7V4cWBjyKqzf45ypUpto9fKaQXTd85Q4E/SO4FHnMWQROSPleylw+7FukV0G6Ize
5osgkUCkj1qWa4+aQas2K8aJbcASJNPxqeYHenMzKxNQP+x2bmUozC41qpkW/AK/DY2mp0WXanGa
46B0gl+K8+yxGR+bs1HwG6GkNKzmj44EMXMcXdEMdNNCaKQ2PemSTSKh9LjWwTCX1iLOKqM4n/UX
8/f+YQ/So0kE2xgICj6HvHbdeWShaJZ5SCDv0XTfzIejtvnv2ARwUtfEv+vCRVc6d0Xv9C85Hd7z
xXsOMP0j4wIEaJhMhHlqHIprrULVW8UFtuuTYmq1vAwUXwmCXQWmA5SxYdO5fQLiCgy+eLg3vwxf
UhnR6PvVrDVtQ+rnYN898tMq31HGDwcvwDOOO9C+4GNo9YVRHB6E0ONIzONYm41drhFI+BjaogM1
+HShHUWRqum9CZSrdEV2RpNsSju/f14NxxzX9u2X4PhRMLFLsid0wBrnoCE2f4OMsx/KQQFFmEJR
RUNq4dxKPoe5Oarqf+MVqpL6TgGMWiDgJu7oiROaB5nb3M5DaUuwwfQ9WBvfb0Q5rH3tNQW0D142
+eAvl2fdpfHrTlR5YLz2q8U75NGO47y99aoeOYxszHGf+8LJ9a7j8iRyMEOmk6uJgd8YhqHqdPb6
RMGAEWjPRiV42yCzhk2k8hNJuIbUiHqI0q1EUvQ/ibbBhMsZZ7u6ycEUtzwYdKyx1k6Iv4jNWLX8
LBc58H5T8aBDjMn+A2RBr8xczeIPu2njMkRM26JIMItsX0+s/DqXG6mUzcKalRDRRxp4GbnqRqAg
uIfMJys9/Po9mvJxNoC/81za3GvEX3VZL2SAPUR+DA6167Ek3s1EnitOsHAudS96zCPeKsBsE7wn
x9xABLRG2NFIHgkcfP1zulxCywWHerPVu+iB82Qfs9pffB5L/Gi7+BOZxGDBneYIqh2AKm7WVOEC
Rzxww6HqfMIN7NRL9Y1VQn/fvoJ1qY4GyV1I5CGz9chffwvJ8XoshEtrdNjpNDuKdwxJ81JL/62N
LJhrTXR5uIT/51T1vA6bsp61hfZcHcjwcU21k6MsLAA3/sjrmfsDZWOlbf7QexLHowMQKEI3IZxE
bjmks0m6HMEszv/w+MiBK+rJSIeTfNFsgjOT8fUmhbB+iF9BXMG6j8RPPcPNIFXWkDS9MQHM2uVH
UdVER1eiPpM89gHJnfXlxZsG0FrOxCUWP0URVi214tgIbpqzgO3aEUezXdC/v3O8CyjSy05LTHZ+
T6Vl4N9OZUD2LIvEkNIs4h2bY3B8esjn3i199zf8F26HpJDczxrteHmmuifP+ueJvluN7HHgXBH0
szQCi+hXpGlPTWXx9BSSBN+jqKO9TR3/Ca6UTZNjGZNNYJRn0HTckIZ7s4k0a/D4rqhg0AvxPb/y
f0Jl+LEFV0YrfXO3vL0FMEWQOz1QZqExX9mG6qI/5ckOB03w+hcleAVSNbAo/gcmnpY3BY8Hd1Ms
eDhZJgxxzffuz4Bnw9dedycr7f/wCrikviNHRzCxE7ypqQA0FZIuZNRD1osNdqgMwM8VYqVFWs8t
vase/o4WQTSZ0i+GmyaO7wbyiHF7sKZfffD1Jsa4/TbUSr7NHoZd+CLGw4qgh1jot0AhtQILbelq
WpaRiY8olXQAuHuK+f6CKaVzPceLrRHCDY6qtx0KQcXxsaP2kGAHEXd5Y5uB8hWZEv/7aCoujOvQ
xGzPy6ix4uK50jqFWvKIYPRFdbDOWTe5F8C51lPMjUDpqEkFISowpzlChawy+YPgxzZEdCEI195f
qd3grAkcOQhRTHCV1u6ouL73NP15/KBq3qidbcGsXMtw2EEzLD6UOnW/1BOQZsxUmC8MM9EiouKF
CmgVr6P31otjkUrIYXTBjwqNFDiMAJPuqUuoe2JrWFbGBJkZkk2X4pDIrGZma6rZBNkIcUOX0ynO
UC4ARYhdwlMxokM2GUZl6WJaX946Gg1Xh1XJVobdRGEEtoNQOPo0R0IzoV7ymL1AZE7WtVUYQtWP
IgYv5vATfKb8jRHW4Uf+/I8YHRPE0w3kbU2XU2mBIAPY+XK06wIT1RvkrzhyZXeE3xS4oZi5ph6y
Y4SV7GpNOne26JdRFcAXYCxksOraGkMTmKwTWWdVf71Y+ea9cJnRooG8lI7abNMV+F3EM16F44AN
yM8JACMkw28qWdOIm4ajAf2/Qxu7nplJ7otzHceLxSyVcjRD8WtBRG9CfaqP61xBqDmFGYvkZ19o
pDozBr6CxJxc4wAAzfyEnelX93GyBuZNZy+QZuHPyiDKcyr2mHq8aB6uQq8839jAmuwBFGgWvlgl
8GALQralJYpqsp4eOCr92N9u6J5Yl7vjT2hpdkXu5IjIV3YmKeJGXjYGH9M6gryjZ3DxRjlPc9UY
wH/i1DVUBe3rA0n1smftmSBCf3atEBAc/na320l4hmG9g7VEmSazc4KikxOnpY7I+kU9HVQsnrW3
X2CCVc/Ft2aPOybxQyasrBGATHlPe6hOSFbb9oef/cl2M+ya7xsyFQjIWJgPAvSBOkWcAJ4EDT2d
R6rcNa2lRBZZSYxM9fyLzaBWk6QUPuq1cNkn8p3ySyWa5fxQhhC1v+10uGLJ04XQ6kijhd5e4MD9
0+RKtgwlv/7S2TFa+RDRr02oKFf8gHtsfNhqYd1A2t5Ac0dhPbTIxX6Nop8mf3otAespXIaAgO6X
iSfpR8MvV6Y4PbuhjKAkAejzEtHT8Mq44j3kddqlyIpcdS1cig+/SBLtTDcNjQVnQcI5yASrDpPv
pAafVdtgutYDllHvJwVtOM0Qo9nZKS4n2hovITO/aAoHFivx2KeqR/vk9NZWuqaGReX2/MPNt0ku
pXNa7rfWoPFHzKhkiQ4VxDg5jfe+MrO0w62zjmRcDiDL8D6fAfCW3vS7Agz5C9JfVb+KfXoU1V+b
a3G1DBfK8SsMOfcl8P6vQvIWDsJGhp0buWYszO6LbG5GL5qvpmSUTqD0Sbc9iiFK02Il0S/r/+rt
TUnTzTjT13Xa295NOdz/M+CUhWuNKo+sEyGRJ+fZOXWGCHxKzzLXxwsDJp6fegrV1nT0xL7rq0cx
cy1HrbWJaqdzHfN30kxjz406i/r8jx4T5hC30Dm94EBCmGVTH5gRYJUUShS5Y4VLSoSJc5cglPUq
TXDcRQHO9q3xmRSh4zJI5aYsaZ13OxNvD+tu78nTGpWUMmNyw/aFEpZvkDDhQNS7SSzyquyGu3bx
r0pyZKi8WuJ/ahwUIOtXYSmhpc+Ny2doPSdvnw2FWhivlgu7gnWG3mBVAr/rd6JTKDczheMxXZ6s
5ODKo5asMxQ/trcrq482e2bdC0tjaL3qk2RtyDHngiIL84I9WQmCcyIRMewHeZqGPiWy8WujDAAs
x0N/QyrgC+pUlKUqdxkTd8ZVhWmM+y55GYsbL1Zk0TE9oN7A24tNpidQivot/vr7qoqT4+SUi8i6
RLfKscxwBnHqO/evG+GGZ9Fgrk6BW6cReJ7wetsUtXg9yvcT2FO1Mb3jcHUeaKUJzASQ0iDN7qTE
wdyVew1RZQIsha/GOhZSHpJHPOyiw2j7O4sLE+JsTsZja/X8G7dUfw6KgvI/jBg0Y7OZ3dTxhfcm
vwftzw4D/fbgkxOs8aEVWZMlGcyt59J0bgr99NEVISnlkKFHoEaQzfVPLNaCbZml252HowgUICT0
qsguvAh+0WekjStR7wxno+ZDNUcSx0GClrueaoPSA7qrwBy48EO8gZdNSbRcpcmarw1KtiGoUHXu
0aeqDmVk9XXUrUCp8A8/eIFbZ0upF4NhlO1VBBGyUOEnfncy3JQCuG1s8uMX6KLFnZbdCBKmA+Hj
e4XZIJY9b6R2P4QSoD+NBattJIE+NZU9TtZ+JGtRpRIYwgatwy+4qB5qeEELdM23AHuTqSZsrNNq
ctAXMAf+ljYEDALW7ISNlSbMfgIOlonOoLil18tSnu/Md82GxI0GA8bsNS1PrrEnFIsB3IAxlqdY
McrWeX+FYf7VMyr3O+gELCVbGoFmSJIEWQ4rE2M1mqlLk6LjLhgTBk/QOsJvbwb+L5YfkavXBpzw
mCEE5T289FISx331sp9UCw+OqA6OEYfJJRGXCg11QiQkZ7kckEOZUJX9fUoi4Svb4kHtgmHjuXs4
51xOvProW+pfOeJIoQA3v7slZUDt1Nc458OFSjZhkcagw8TPZdF0Y0ROKpoKY8K+y5ARL3NgcdlM
TJBUFX8JcCL/MFxE2FXXbdep+QHWZlmpU38PABgvK6HmkrynYrRfwaanSKDYHE1r4cYd1ZfZM5Xe
uiYhM7D9Ye7RADB96/jXwsRCTSfg8/C3pkYJ8dOBbbZRuYG9OTB0ZDICOj2CYp0/olxgOy+SYB4c
fuOZhyxex9HciipXPslM35TXI0uzYQlm35cSLWQVQHXPlt3KRvaeSZiqATy4kRipakoBz8C3rZR7
6oYEEWA0rVfGFNygluW9GBlZjhbvXvFQgXMES1B/PY5c1+PeVVKXDrNpwUGxpknSXuHCEw0WY6I9
Z6nGPpwbOosu3WOdaqo9nYESFHcOrT//E6Jop3UIeoIRzI7KyswFhmI8CMqrC/GHYJB2LAfufmMs
R0L4WTXoqPBuB7nspP5KhBxvC6KH67svxdR5r25li1qqbsGmncXyiB3AbMUuemSdTr50Qje1EpWC
hclKsHacSFs836Jz4HQta1H1qgSRbK0pnR4B6hJAJFZcR1uTPwPQ2DtxHmyC2REANzsLrxNI1In4
ATJm/AArDEuK3gIdSYkdwLtdXTQrDLSIN0cjqBfvlx+Ilz3fW+3VoZschkssLm8zBaW0jcOqLftF
WWRfQQMWB4xkoQ0lcjL/WmipLAF+3sXwCByr2fUyKnziTJd9XaAM2szbCxVbEFxA9mr4ksjj9Ulw
UNJDCVL6QrZDO65XKgNMw9iCdlambHmI8vjrLNMFwJv6KRAQecNpqAb0y3cp/+ES6n/R3tDEBGVp
Rb7PzZCMmCVFHPbD0ha8lkq+RBe5Z4Zz7XJyfUo2Y9fa1bvW0mU1m1dnDRh6gp3g3b1XAr5tihE9
QmRLkFQEecI21dee0VSuBZrh5fQbNiTuJnVo0p4Mm3SP21EKHAtoWAyEe/8iYZ82JGXJBZi4L9T5
cUeWNQJsDEEESpV9rYxbyHUyPoBo78+237oznEOdu1lpIWxNbtm2Q5EfTpCFypKKm/Qvd1j5TsEy
qiYJM+5O4Vprw3wsFIXzNmgrtHDxXrN7AUUEg76MWlPKE5nBIbryg1xdoDOkf7xjCL1YNT0rdOaF
8U7wTtv/qJDCp0j34ASwSt2IVA/TJs9zv4uxB0hrfAY0jkxPN+UEmNqdvlk+lcXxlsV19KxHV4/3
yGwkLBbmmBMhIinzktLl2O7OFcrsOhuzL/cyutMU09bZeXvqYI34ylIzINWO/v+REF8xamP+cwxc
9TYMO+u0rHHNV/10ApPW9lGE66NXdVK+0UvnW18G9mPQeqVOW72fw7f5KOyZZqFsbrm7DfPWWeQP
xydg9vMoYnl+uDzunbRz94TtuacCqWaFvJps7wF4vIf/IA6+WIquP7zukDUCAiyDQ9w1E1IhE7pc
oUDXjhVyjOtOkCG44v+3aYVvt4dqxj/7UUm0edcMMR3Tn1P8DkkdynKDSRjnOezX77z4btmQl+gF
aVVBWiTjoqerXSu2z2CkkZa3yZetH/M6A8xYJ+t+22CFp4khjhDaN2sULJahMq9Sd8kbL895SXOp
NxkGOZNOWpNgO0g7YGgLus9B7vb9UbuYbwz4Aep1nLTI4nzqTPkHuf5Gk+tENzi3UtQCiDx/q7Xb
tC5kf5rgxGiyMZNkJ2qJ9zNX+JdcPK9HmRF+3NnvK6iukJXCxZdvnHvCdujPtpARTZxxFIJlAkJX
8o3PnnJOugdn57yrlkJ8vYH/WraF1wbnp29+FxynJcKDTUqHaovqJD/+Lnz6APbo3R9RoY13XnVj
5VQPpfMZHS/MCZ9I7e2zpH52fas73/IOoEZ53W0QgU2B9+Gun9jkDTFgY2gf4XzopHDg2dtLbEPR
DeUkIG+/W4VvVPDK39rqzM2UCUowK2SL5xheblhUMHNBmZOeZtcuy90TaQy8c8g77unrnTzyoo2i
IkMB7ouPhk5Pk9wiGo00LyEjrjVbjuz5zD3rxx5/F0SUyR71kOblIStvYWPXr4JR6aHA4myV7hhm
z+mQkGoBVAW8I3loNve0C6sURUmVlVe+u4QkYXUI6xtc/2aeTY5555x+26QyLcpvQmc9DnaVhn0H
T6Y53hdhmgV7+bR/ZCEpu47eQoAhKA7yPUU/fp01ANSA5iGZ0iYiN78BJu0D9ROk7jt7U+z1NN3/
h4S9JanJ+2zQ7ymbgVMwUZlJ4Uf9KBdL4mybQ/015G4YqBdpIJnq0QR2rEIyNc4blWteo9V/UOSZ
5IoPf4Ki3jlkRdqAs0lWGFJaXDhJZ1YKRy2YZ9s4iK3wdwtSoJ72kIm/44mG+LfHkvu4tT13xnhl
0VDkCHc4YijXxFEwqg6HdXpOu5GhoaVMM9maDJlpEcKBKcPUj8djXjtI6/lWWicl1KILKr73SVr6
LzKJuC1xwcK3eeddtP2A4OcIZigHQZe1gMh2+H3/6MNKfF1dOwt4/u9ukHbaMxQrUemATXkC/Sou
6nh6Ntn9O8obQ5K8Axjfwq7ANgeHk5xrUgu7rQete0Ij5v82RP0VXWtbC8pHy+LsDRt31QXdGkIw
U/pOO0NP2Ftpag3wdWSTKp9Ewevzi1grNrit2fvfbQcbHyq4EqhV6ugnOjxQt80kDhHcR9nkzoam
YiOjEloau5iS9m9eXpCRUtLC0LBsbnNUSjZhOl5W2bK90QTp+xfY67K0NMMKko9WwV5X8PUn9pLR
cKsX/TpyO079yB2FzhD1EZm1FrxQDGJra1zpgHolPDRziB5HOfZjF7+ck/QCynh4XkkRitWA9vaq
6EMxzeawXn/QFbc0VzLV1bSBPdWZAC3MJmN9c+bQo4cgXaRmUTPtvs0rJjfGAK6oQUIdWiKMo5J0
PmCx4VD/aIPHKrlpCKixI6spDe1euKf8P4t9/oPxTTN2cvaKGA3iIN/Zv6TfpwYZaumoLVfomRV9
cIi7eH4xXwAV+fuhoIS/zNEpqHiX2A6OkmSfiFaeUEBHXq2qkv/um1x9Pv7kopFHzQRLDxqDngOz
vJgA0kkdBnvkYS+2NYfM5fyLTGlZs+6Asae/vCWwiQpWP2dCfpmDaDVTaxx+kHQu5fmPMNAC19QT
S8y9XmNDOkgL/s97mK8hpYDwIEGDCz0awoweJwnPkgrEIVYs5HTDekECW5fuXgUJKNnH7mnNlWoV
pnsGAmUEbFIkE4yhQNaaEP+u9uaafQRqFeaMaQjc7/s7VyCvK9Ivqy+CkSvesQONFbVnHkiq+yzv
h4Izj04VbirSLrI9bITo7g5xGO7PoD4+R8RFAj4mMZa1ZK/F8ixaioJfDw+D6VlxQwJMCHCgOM8v
lDQujTboad/FBdGtCujG9POm01uVq4qupodZFcug7yYFi788HDmryJx34mgsPXQIHKH6em60Alac
Czqo/k3mHMJpfBRAsfc9bxGu1bRDg+5u0WFYdJjNKaWKWvIFlSxrMQrk3k9hEHRmvx6qP5ebyZua
qjoGcv2gUeUTMWOCjTEO9JF46z8Oh67FD3VQyTtOJv9DPeqKtVX98Z+RmjhWZostVPqXbrdTL4Ke
yk0di5+pWKUVr1R2+eaSZK+u6VTaHyqoeDxacnE0ElDbEAfXQfwnLmKYlDArS6xCL79MSuZEJ7w6
pOWcBfYATZ8k4SgWIGzQYXQQrZ2jwI9JFV7kWSgcwMyuhZXxWO9iiGuat6Y6aoqLAgND/Ui9zfq+
6GL7B3Eh7DKoT+puMaqLJMBLVEoZ5dxBK4FXtdUOVOEOyOlvIlz6NOfNC2QlduCH8cuQlLMAkwUE
9TRe7JP1J8boNyGSNh6szZSM1/0DbmOEbUvg7ORioXDO5sVrhR8nCXqKdz3Qpq2n641X/Vcq4AA/
BoQHqOCJ7rl3irn7OWJnxT4q9qj9yP17o4rvkpXDT4UlWS/XtJVjqp0o5DXTXtd2poDliftQsT6R
/mu7BSaeYto9HOYDu5Tw7jpECN6SybB9E8zNx279MzdEzbzCOHNNO+4fJw7uBdPNyPPuXQ3kqsHw
ZxctgvwxzIpIzYXS0vfPbUdj+yfhh+to4wGyUA3ggK445t46NCojUyEusHHBk0QWe0i5AZHAlmWW
W8wZLyL4cD8WO0/hB+NUFYxjO16EyvnEXRRzatuY9rMK9WkbeWz2EkuF7zsAKb27Q10ZkEFvqO9v
l1cqAfsG7XvMMuw/XF1Q4qKZa2Bp907V8G5Oxsd1W5mAGLgmk6zY6G1pFIzvhwdJZEQoBlzRhkXH
+WX1G9+7MsTL9VXjtAHk7Ur7BZpca8of0xC2QnOimSQES9ItsnwLOE5BiRWbDuNDgdz39h17EyQe
jy8z842pgpazHSnz/m3WaKdMh1Cbs/mJrndII5gRkikxaMNl2xIEwZ2ilBKq71Ezi+t3C30JC/Iz
IKhWz2BofHUTN4IqqGvNOnOTuN4lVFJ7YJu741VHGSXZfejwqOK/aa6j/icLY7E+i80Seb1vbUeH
ZQ0U2JX3Ggyzox+Mo1VpzINY1m+T6eekAeaK+/5M9rAAK0cQxIobB9LmGcbB/l4tb6kP7MYGHs4v
StfD/2cH9ST4P6Kr+Q+VIofVGWzpcc4uRU4Mo1c875b0vM8uHS/PaRyQQp4WBS7t856g+Wl1Jeob
LYOZB6hhBw0g347HJgQO+c6eozhmWXKdwwf6w6IOlQL9kvJCfzfWVaCcNVgGS/KT9fGhnJQ42KCr
eAyjY7DNGmQgF+cVTUF0Cg5r/mQpCVLFy42p36nmeD1/PIpukDX83pvrVNSV8vnNNKMa2wnfM31S
kyKjkHJ7mhG6gRdi5dH14XwYiA1rd94hPQr6PO86kfUrqTrzVm97zRxq1mHk7Bt/d+P6vLHOdtCs
QPnDs7kyHSLwnfqvjHjkZrxS/zsHhJuFAlupmK1zYKjtO6sTX+xrY+8KhSiSDW8lylvrkRli2/1C
hdkFqjbcjaz/fJI2OgZcgU/jt20z+VRQlkX89BGGb7jPJSfgK0HNTrFBoSLL9fbQ1Gd99sk3h6iy
MPf0fq0vc8jWLz0TPNGpQmbXpfvYJZsid2cXBxXoxwmUi0Qr4XpFz4H8tW5cu8p5Gh7iQzfWFrmU
LWy6b9WPnYRGE2MHTFWnpz+3PBq8kRUFAkDbWzBCyjDdmDAJsVSB6PQlCoELC2niRG6GVxo0WOXu
ha8taLLk61Sfu0YrxkVW9G8hHQRVdE1Zl3tZID8L0KI8Il5BfSdZGc4fCpZw8P007OhDu2v9Wa2D
dTdDcf+CPzJWvCXggMQBKpTc/OCJZhL3toWwNvx9NuHxJGe0W0jL1fbGxRAgZHp1xn2FV6uB0E8K
da/VX40iY6W4QYo5vr9O7FdBAlJZFTAtmVWABEnUCbKIoN5vc+wnUIQ123oSZUfaS1mSmDQdKIda
J6n2j/Qi2Do6T8T9nHmgVw3ApYVDjYRjABkEYmI4wEjUF+TP1QEFTQP359gl8H5DQ4RCU7b9mZiS
UexGhPtYZarBia5Iz45u0Ipt3zng9DDYq9aNwp68RadxY1ELKSLJQTfB4tbr7L+UuHVzLRmaLyEw
Vucdos3l68yFvSYyM++q77K57BH7Vb2sJJUMfyqKgSuKNft5I8LiGW+FCfUvQqcnMrG7CZQr0TKr
5JtQjJzC5I6LsbEttUSobSJSwqOJ+g6+scO6/+AaYgKEr+rY8cR0orOh1UH8tFL/p/zK7ZEGGJFm
iqBUX4/4hT79AO9/77W1eOHL00lN9RoOgLQOt4Dboxr5hnzFNnYCFzo895KuLwG6jPUoeGrE/APv
AgfyqkXYE/adbcFq4JMXErqeJfG28zxNZ7k5PD7GQRiMaLqisR4ZI48UlvqfMGCOR8m9iWeAMsVx
P1MQUS521cxlIwcmtR6Y46/9OImlgfrgONLeYL4nbhVgorXLfaKPDnhDv7pvhWFb8jpT9oGdHC3Z
724AoJ1EcBhPir1w8iGch6R0yZlE+ieLnJKue3A0SC2hd1JJmlyU5HD2VrT+2W/6jN/0A7fFo+NE
SECtvBGeAf5Oj7RCmh/Cw23RgSPytvCbfZ4dPfvnzlCwu+au00eD6DKlnlFNSdeceAikztM1yjeE
JtB0098qt6CZiDiN3+drC9PbFWVZLYOnT4qZ7juVbSK3eqhnnm9mGCVofwong5tQsys4NXWhHm8W
1W0K19i+0G6MyF15e/kfZ8e6V3+rDT2IDgPKK67+2/d0YidlTTtALAZrRPpyf8Gwhe86SJfhnMB1
QWDnU+VbTrL7pSFdf3vNK/Qs21caxgtAOE+w0WIE8dZckamq5005oyVo6PkYKBcueRh+Eyrmo8Iw
2dKGKyUDkjDQfVazPen47x4SzUGKaDSRNf/Q/mq32galDar44PP3CadmBeoL7F8G+CRcf+d6aSTA
H1KJ8AlpxI1hQHxC8xxaK3b3BjbSjs0C59cMxuZE24OhwQvI4nbVDss1qEYr9HYq/P4PuJHLdSPE
xgfKO+jAReG7Ovrjc4aZpuB9/KA/aRIvqCeCR9nHdgwbMSaybNGt8Ui0XW7QhqAGxWtqVOxcfEk+
9qVpmor/Ar53X57RnBtIzGO5N7UTVQJ1JHg9kWlwifeiHBbzHhdthgyt7cjtVg0jT+LyBEff7yd0
V4TrVAHZS/u+yUvYSy4Ry8SMf2UGHGnn627EkRtrvEvPd2id1nggbH1DQGIS/Z3bqpiQ/Bx6tlxF
B0KiopWusAQQpXodBWvj2arO0TYCoDsk92QjvG40xCuB28kZZouDkL2FreL7LLW9szIlJbCC7nZV
Ib0QsSGvPhppiJ20enRg12JYkzzdpEtesRCJ58lwnm51n8HJraSOlMo434DILz7lcRdzFZ9oIPm6
FaFpKJ/AoCYu7Qs8xtF1WLZ5omzXY4LbxiZRTopwm4u8BDv3/tFYiycgdrUD6i/dSID4Lkju8rGL
t/iG5zrk4J/yKIRq1E3D5FyKXiUpnp5/EFpX34zXFy40/8NqB+GVqHzxhGz6uEhEA233wKDWnX8N
RZj0p5Ehh9DOBUaOeAYSX9pJY/7j6eksmXL62m7OuiNlwu2mp72/3TlcN21AMy/HxfHQBtTDlGIT
HFr5pSYSYhh82Ngjrsl4IT3tHDgbJKgililwwMxCaGdWUvJIHqjuYxL9s+s3qDu2rxtle5OHNCkO
L9LKKYLv8aKHtHZxEGWjZ47dJhIxLAtR1tQlhT73jvJvNwffLY9NuOl56/2jxCwfrg/FHlK+Gv+D
a9PskXUpwifYQC5FRfUgFpWa/K6Uz9XbfuiUsHEZ7EOcgwFVpmMUbnExemyiLcjWqU3vvi+RNDmP
HpyOrwlQTKIlNTgtXkxPOWENsI1OtUbA66JD68cthoGbYvP/fw4lVMG5d3jrbE5htRayrniyo/FW
kSGugzfMxJFuHekod9UG+DAtQUlO5ltny8IC8MvMMuRL/gNFuXckmlty2WcqlR446MKykVHAsCre
tDnGJi12dFDvV+AiObbMa1JZkj3xdTyqUukuz+mglW5mfTPKwQNKQ466iSmV75AAVd7TMn40nwjU
OIEYpMkeJaCe/SbFveek9bTk4gxXtLv3hlLIimXHibtm9GNp//+j9kzGGB0+PUO0nO5QM8i/dJbI
TEtaZWbvF+lfV6/K6WIc9ErypBn/gBfhTrnKsAF6AkU1zppAIz0Lq9eB2eEPzMqHNm06c7MXcHo1
Jnsb6xO6N0X1vbutkxpW8UHwJGzlxKLSOmAPPGz2EDTbl+MBBqkv2Kl9u/bDfPYoc1SpUdv+20CX
LLBpjVlRN6fzyXWVoOhuWkLbhJwQrt3lz2lLZ+uKk5UzvJF1P98TaD7+Q8El89MTWlOQnmmPecvc
3MBhbdOWYlEGzbqsT1+AxtjA2zbYECF+0kMITqY6mf87NiiyxI3CVbIT55ZbXvjprpasIJue0qWz
f53HYhpZAxC2QeYdlzJ0fnERMeWqNoxJ9GS/GXNpE+8hEAyeQhlebNQmtUqN8PpZCM1gUBMEv+zI
NwmxIQ/E18FHnLcB9LQ1AYu7wToWj509JzHzHtiHsYRL2rCpzs3Rn7FepEVrXdDblsM3CNiqvazH
pi07wRvLlIUZcsSxEoAHI032JEnjrQ9us8THvKYNFQ0gG9SQd7l3rCI42F1wdjvfDWjVtDCyoV1k
fvSGmbE+hlVFZUXlg8w3cl9OBykUUaDFG6F1mW87vM+Z6UipIaNNuWqsiBRNQ/dtJugSup5kHSxZ
2NBp3odKj26LZtpU7e4DqWYs0+5cRSi21OUZFdszx+ufFURbxZXbqyApMMMC02oC0RUOTAA+H1X7
VMsqasx9BN28XGE/iuvjOvj7Ycqmr7QBEWJTXxx9wo1f9+PvxdR7KUYfiZz5JBH8yk/JlEBUWiIC
hkqXqTp5ntVOOatXmfHT2U2REPbTNqVshPH8Pk6GYcpjWGb2x7v4MLHDbh3kJQ8QufdOyk6MeAf0
sovJ/PHXfLPS+uyTbq5XwnkEr5jB0TKOJmzHruDLPBY5uNbgEE2uclpQIdifPo6fb9pleH8EJk/w
tYnX4pBXrd8pVKdKFYy6q2h9CKO9EA0coOyJycdwwlG6MmpJFvpu9PDBqYxxnpkr9mIoGUs6BFrL
0sqihxt6VtQZM7TYNQ3pmcJX0h307izzYKWdFJZq/m9CcOVi888ITaAAKYrB+Wn69QA+QHUUkuUN
iOC7dCPddRnIMDbNu4/P/3nZ5EhALoU7/pmsWD5RYCHouTJk7I7HzGEUCVBA5iiOK0o4DQNaO5+4
oGl9uxJXgQUmAekgC43JhQYM4xU7infyMqQmuuvOvrJMKLmMIW+/fbdMMUHvcZEXbIOHgOJ1eXgj
4ePqK6rEiYJe37iW0jc3wvUKwygcJ8JktUNVloMzfz/Oub1PAP3Q6uS/p+mAwM+GZNdql5thNxd7
E3YdVoN9N0QZbE3ZbEVokR7xGCw2LA4IemEHDHgzyqAIidx6G7n+vhh40Js10fzy9xm+Y+ACpmRw
SUqEL12Fr/kJGVNZnJaB+XKLXBwhs4PrfQvwLo3nl9jRrFCKSJUrbtu727I7CeaTms0eeJVFb959
h1ukAtxH4tcf/b6yR+y5Ve215waK0hAZFcFx6ueK08RpxooFTd1eGWUbW4azsGAq922NhAiI+wyh
wY969/2xRQF0eAIhpeQtbXdFPJKPpBCwDNpF6WDOBlpxX4G3IGCavNUsTmng4NthYgG2vSXdEsT3
/GkvcEvappeTMgxZ9q1XvcLQX/p82AekN9EYtUv0k6HxJrHHwi/5paWOWEJgF2EUl92t6TPPJ+KS
X3XnvVluxQ4fMWkOGuxr9V0y0yVAer2LquXkUMnd1L8aJqP9xu0RYEKXou2A8rTGhvUaNunl5362
WVtKDNay1L20ml/3gprsu6a6538Kvj3zMtOWhEfWuTxgcXs7XDmCM3UxA5KLJ/TSWTcn2uNXo16L
Ur8V45Hi8I6CKcdYlVlqx7bMiYflrp+FPMxjTs1lKBdCzLt2sxEVT7QzR/Ba4V0meW3VNlUrW8Ia
XTq+gzL09aj70rNNp5rr2I29ZzjG6wsnjlMQTJ/XNsupMb9vFdSHlQjDK1D5JkrL2XflArxYnzby
BW/q4UVHFgfR0TsApOR4ZRzWd21Nia3m59T0hNLQKAsyHs+xce870yqwHnuoBdxvRhqtmduI35+C
Q6tObINIKJF98sIekGvlaDV1yD6Trhhj2byt/UXRwJUPtFxDVRjFQ0FatZeJ8EwlMEBdCmou3DCb
5xvdAT4NqqeRDhGu+Hy2HRTGHufKcBEG38SCMmHEnwhdhdOjBi9ZWJzVOuztM3DoamdRc6hQKJPQ
KwNFUNypFTHdFIQqKSg+iqC5efiY6/JCXGviTnX2pVOAUtfmf8iActiUrc8oo7XxUHoFLE3dZGKf
SsgrPc/LBpG23hjQCN1+2OuT0G32qkj47DdEmQuQGmZBBsgcb1B8M+gDH+TnIP6GYvN5iL83iZUj
Kf90ET8f5YeeCMKasizuvrok169jzakRhktu10Nosp3SiB99KcX8ClHaKGmzRvk8lR4IvzLZiHsw
wcd2fvTGZvFrcnrx6GvmYMcX+IYn/sz/rw1bQr4cLLE6VffGMP6BB/GhsQIPiMGRdNJ4ZzgNxYWe
axPCIs/dldbp/rmlJK8YirbHrXTW7uxen91CQsIrWhtNQzRv9LRUpfLemxXuXAHYW0LHrbVbSve2
Yn61VwyRVa4Qv76HuL9fGtoUVuOIhhmTTpXAq1PYcqzNBYdPr2gcV/+aLGr4hIH3IIyv3G6nqKTU
Xqc43Ntcz5fMKfPTLWaLAgwzP0WCVEtZPibF4H5y6QfIKQ/Jx0MjdDfPMm7bkk4B8ZNYD+MmgWJm
Da4UOnxR2E3F+8iUehuoiqNP51jOybOC9vpmqZ/VlabmRHnoDUcB+Dicjc38DbNZsXh4YnNZhUgR
x8wfmwh3rVPEntUbSgAjyfadbU2PwPJGZahCNNEs08xSwPtLXO0rgy69e99FXuHexmnTaLlTzldH
8I3inSws3f9QkKqZ4PoCI32GOcFrwlY2sTCTlKtWUoMy5IsDBECcRRGp+tmxjJJ+qM7InYgVqBhu
Fn7eJ2GKAdR4IxyGviGrNqd0yHCzDJhaW9GuvD1rKpyMT7IefGX0Z45QgZRTNPkQ/LWD0EOs3NRf
Zf2owA4jOTacdItTXrb78yg1UdJ3xMz4HL1EaISQ8TEN39afL4aVauZEXxRIa5LUMBXWmURTrWvq
BHfF+HcH+AbwL//PZTAkmakO9I4xCznIFV42Iv1LPSkfv/btPV2OuiUzhC/7WLpfu4n4jLfK2w3V
6lv2GzG8H0aXHtWxNDdbw2vsiZUoE1dNQfHfh4xsKSEBQEcgDHhzc46XD0Dg2Ml8e8JCb09AJQ+/
0Z09t7DsikH0FKZCXrEEoqL8sE2N1fladIx9y0kiojhZ9KvgcPvfgiXKGh6w0cI/PkXtAbEpThvc
K2KRu9BrGOIlUSRiktGDwQ8MKnolPVFQam/cVjLLKZOsQFaXDp41ZljDY3NX9MPYFuDBYls+4ADX
CGV+5RZClLmL7iJdNQsdrn1brixElfs+PZqjlrGLYqptDjUOVpmU3izRZJOFM4EW3p9y9EFSRCrl
a3dcXw6dHVa2AhCOMJM70QotjAqtXvmXhgsVxQwBIDECh4heEXJpIXmp+E/66d/iT84bzaMRdZN5
0akgHaUzRsrmGMBfVCo4MRoQltvGwKwFxh695Frx99e3T56nDIRoSpgunEH2MyjHmlW1b10xxktg
jXsmVdLppuhnkowpWar+lOZTVuhSUaKmXeFq2N637NDNm2Q2B1PhNrerBI3SlkBWXelmKE3fNfNr
V0NHMu7KwhgEymoMOwcv/j30sKMamWIpSgKFYgL7z347WGarB45STkjLRF/oCJ7MdGAS3RGHAKGV
AFc3Ktbw0Mv+HeXIyn2QTrqMfMQVAXfuDiY1+4LdXZvU8129h+dmNoOyvlMb26m/qOKvJs5z05/8
LAVEQyoOl+LwMuzk4yr5RGV8WPfCzWLGgcTdJU7LcQemv0KHMIMmKGrUdHdusOejr9iDIKzX+e80
lfjjKn4+m2QsF0VbUPbx+bs74nE/AUiNx3Aae9ut7fjjjnzHrwnd0vvcDoYSnMC3/V2ugDtB1iwQ
VSPWSr4YZnXzxzqQg/P1HQeAz6auNZwDptjuUVywify892htWCOXELDRUTL+4jD0ro8K+pP96Gve
JZMOUzXcLktvdYFjGMvnXRHIdS1v6r9dvvdSIpDDhgNbkwbgZ6R8GrYo2gkucTQeLROTYg3Ub+ra
R48eMh1s7hevsdMhiKDeMQ3qMIFGHKeGkz67V1D6Tgn/gxuPFv9o7s/ps2IYSgxLMyH1o4g89Hkk
zzINCRc0wcObBvY/cb99ShkWGHosOUoUSmZx9KsVJLCUUUYyNtK91vnuf8lYfkzA8BJhwIudZNsa
hF8uiP4oyNolp2h/EOj8lQUkh5RkqQQHXirzB+ymbG8Ji5BXKlm7uyNh53Nw/uNepV4Tps0ndxqN
BS81+P0wJsvURrlL7SSup49vEY65FluOBom0jdfP8yiB5T4138MX2ZhQckLenXGeJeO5w7Skeis0
+L4nV/QiSmbkZhyjaBank3ct51qplc6brzFIWqrEHs4pMCT6o6rDZTLh/07AH8yFxMVvf9yeTxH+
A2x5ue2CHz62ZSTd+NmrlwVlVc/Vnp2SlMKthE/+pGI42yCKbxGRxh3WCXaDSZkotyecvhwq2iFM
06/wF6N97UxIF2FCb/np3Tv/PkMuCHjFZb1/HwiYOhUJuSHHZbJXhkriDsGvPe3U4BOgrG+oSP/k
MR/Kdl9/VRjH/IqbpVx7DFKMc8gjMoFe8eR9fZ45qi7hDZ4zouPdLEhLx7wnm/BZFZkW1HwNjlAH
Uyc8p4vDgD5rnLjbXA2D/TilqrrOm/5pxO3HD0dIQjDq31XZApknroZydxJRRCo4LeEtThN4POvB
JE9teGB53NiEgWr2Pmbn9qgw0A9DNnak7OhO0CjlqWYO7lAiGN9WugLI72kxTYVHEW+rGOZAp9Fs
XlCB9/Ytm/cidnwcJ3Zh4vSFeDTXQgV4kjafA5tRAAW+wX0754J5XaYi+K+sGBbXr/osfj1WgUev
g7y4ew2gZkKIVV4bGyYFbhG5471NbunJnkM7iYi5W2ur36Xsm9WqO1HzfWz/9qBm9cAbd3u1al6N
f+Z9r/JCnqUfLACjv+jHt2iiNwrvGYRiBsLSl4Gjzb84D0gpJrmcY+WfALYB9YH55PIGZKwMv4SI
aAeHhrpMe/LkAbBxE+Rex0LMsGPtcI5kjwBsLqpgmTps0Z2Zu92CFyQKRpBQNFDIKtdbsPk+A7r+
hzDgg5w0WlpNBVkC3Zxb8OgAiVf6oqLIDUSRQNOMqJ/xm+OJN589Vou4hLgGXqdlQ0eF3LF1qq01
+BneELt1NW/QgOPxIINGGJgTb/3xlozONtBCiPKtFP6XjFxCoHiAXJcgUtsTR8YUPHWNWjNDB4Tm
OMirpiFSlQ225pMOqGLLZc0/3spj7MeSm/k0bVVNucNoZF6T9Eg+R9O4P7QZNYFDJYowcIL4KO8j
7SSP68OhBptHdbOjcUuGXrJTZnYN4ATG9TMSajwU5ji+lZ0mTT7TYYWdrxjMJ9/9GnJM5uulREMn
rHw42iH/TDrSK3l0ekFSedSTy+I4tqdRNO0a2eRG88pBQvwOJjFj96bK6PP00IKxFBe6RUQWuiYf
HfmjsaUcT8IM8nZbqoCiQ+ahsjXa1w3s5fu13yqByYvqbq7S3Hs90O/0tRRgXd9I9FvRVsqtQIuH
VorKYbXDIuMg50COvFSCae2QLgfMONI2Rq1y9BaIjRowyDD6jhRpDhNuBSQmtbsnTO07rATrw4JT
7nEtBN0bs05E6DjLCgLSlGcYy/20ylM4DXg/I3qH+/FJdwTVuCguhSTVn+BNBksZSx+IfRrQ14Rq
s7ZgJsRO/tJl3Q6h7OMe/fDYiJS+idV98FTz/QbSJfoKO8F0xQfsxnSHbzAulCaDQOTlTKrKnIyJ
EHC5r3RhczFx5ef6gAqsGuMKT5fqmJlHOPTnVL3tVE+3fUgihxERY9VrQwdDBchL6h4yScvnj7AT
3BLdQSOc2rPU7aGEEZuk1jMoEwIv5JMNc1vtGFSiGwwzuPwARcfm11VZXA18E+YarO/SDQa6FzPm
xpLlRz3W6nd8kZYwefmPmdgv0tNaXJ61ZuocnP/By79aofMh6OtERprPvAYKVnI9M/qW4GtOCQa9
0xRmKW4Fz1sxYEr7xFDGE+CvVoq/wC40pn/I8VAJC1fAwGfjUMx+Cio/wIclgOPnZbKfqd7HIw/g
1qxggJj2hnH/OSNdXj2C8dabMmB3hk/EBA+O47Zegc2Yp6OT4C2Df2LKMaZFoiepzzJQkfiiWXh6
wZbSHCJEfWlJ9QL4OzL3nInSkftHRXbU/x1wSZpBDbmm0JrHnZzjSnnL+8Pmn6p4ofUvgIcWt2Ns
02XkPi35mRiyTipWRg1krJRI9TKySDg+PYbpu2iG76AkSdQTEQ7urJoUZEgn3050UClbxjlV80Fe
j9KwLbi9YAhpXuMYN3JR4c8xLP8tGi8dnl0w8t0WSrZES11oZeUz2qRLynUs6/OCryH4bKKDVTO/
VQIvn8G6N8oVCrNXy9/iKwxvyx0U9LzfgUvvtHC70AWz8r7cvCqu7Jv9kQ9Kxvu7zm3XPh/RQzdL
d/WLhlHBc0XQ0LzxW5+ONGtCurSYxoN8OvoTp4IDKGXfQhuwpyPI7JjLMkHPPtBTUj3O+mO1PuTT
6FHVzK8dbgAmCoQiE/H1TWTy4+OR7gwnLHpYmmOsfcs9NgTpnkz/aOnPIzSpYFqnZvhb4q8U2d/v
ZQPA02RJ5T/RFyMlx3oSlTOlRoynOixaVr3v2WMgzM4ZyZYn3u0n4A0yYdiGTfLYNrLvtPckNE75
OOVKknodY51fB4bv9ywKbD2LoAogcY1JUdWBkWYI/+fgQ7O6f3IFtJvjUjAV6JJw8yUbUWOOYMOc
jbzvKedi4SGWkBauajpFVbuZO2eKs7TYzqq7gt1w21vG9G2l/VuAPa38zBslGSYORFp1jT1pXMFo
8EX/xU/rplbXbbBCXykkhTw4A5Zr2BCQViEVRSQM3/5aWy6jst7OpZmQ+xcULVrtA3Zj8pK15O3h
AZ5SqfTE86/IrxjEAozwIrE/MZur6baDrRXUe1iOFU82wHqavLtYDLbHbSXfozo2NrtAMx4xf6FC
kIaYW4WI5bx+cBdXPq7hK4y/xXYSWeUSLhNFb4Z2Rl4DIdckgs3Tor/qzPfX9cf7w3eLo1acaNxr
kdVs2p41UHi70ElH+Os6LPh/ni48rNpA4mwyK4zrzRSXuxR3LMp70PMTl2420TzAHh/EowDKhyyp
tRuWoXvEPxI1LDchm5fyf9Tt+Lv0knLLRdwAIIs5dRsv1nOHT0dow5CzLSD0kLmqwwySP6c8eNNS
LH8P3ynNx6fpDkU91Xah+v6k39aDKAiGY8RuIwoXZOKpUH4LRMly4H4AuAUDvp/skh6GUuzOAV44
VkyZ2Dy0KtQ4mDgimmtcAIKSFVhKBvRfkso3QmBUDtHNWdVqIvIrpBlUKqxRBHoOaQWr9ZHLvMZx
zJMy6yp7k3g471bGOsOvbfLzSZzZfMTTWwuWNAhlQoe3p4IxKR5UJoTHd3Lv7ZO6QT4vIIyGPmxI
X4n4hawcXqXx+uQ9f87NhanK0Ow4VythZ28jFXNTwBYQ8dDhRayAcJjpWZ/ckYYrkVogEbdxR1du
nMEv5INBPnte/1Xk0CTVvYhDKa9AxFjDkmlH4fuLCt4ySYT8v3Xhbh+vnKOLWBpOoczPZ6VpTkfJ
z7qzjBAmf2ph8FMfHDakRlwZlOpgFXdXUQNVjt5kEcg995Pid13eHEUvcY78MfmCfou0biczA7/k
FKlPvZRU5e0ju94imMlYM3UoMSTuH4fkdlsSg9TsMLC8x2buoFoDUeuoJjbkArK7qVq/Mxx9N2P8
tWb38mB8HV0rrF1YPqHt6zEez0p2ehcEI46+nisNIpNboYn2K+HRuyQehI/NzfFrwcQlDvKxmXiv
br91iepc0XNWiZWCRZYdYFgCSLv25RTjHykdc5VdNB00KfIOgQ/gGn8V7yv4IUiPgUxv9aZ+HBgG
XqG32KzfK4+8SwgBUSHrkKqR2KCqcrI+L1jlc6+li+NTnqQPz+exbYLYGss4JfXHsrg9qT+kIU1F
OVPtU/QCio2+pOr7qY8sFmpsmyocJx35/eee/ebHNCGHrln51SPnKAy+v9HFcEkfZUhkdINUMiEn
REx/4wAEWe8RkwEvzFmyHnIJdrAR/S5Njb6+wkqEVD471hBS3a6U4KCoLYTFBnhX4ffyDo2cIMq0
FlceurKZDvQqHq1056gMsWivIgkkHR3oqxPkFSvu6mtml9D4c5QPRXxJF8co9BxbMguercXxu4yE
tDnJH1FeGNUqvEHh03wQfZPwxxSqiFXZjx7F+aEcUm4tTZZVi08Fdp0GBrl4nF+ylr0AH6Y2A928
iHCpRFiMo2T6Vxk0Z9PsmMMjtyFYW9En5vsWWnsQEdlCV79jQIuoy548ocm2SDCOSzHL86EQFf4j
A+S5QV/CPcYpz7UO6XdsJXY4QpV0Thfdiu/sZwKdZSDs5hGo5WOYzgmbbH7WjbDxzQEfPtIpG6qx
IEZFwAcelIKCT2tR8v7qoCZENCRYLp34bQlXcoclrtPrejtVnmlgV41dNZrRpiTwL6HZj/UHQ2Lx
jGY1cl41vNQgk4XAKq6JsbL5W41x2+lE27VMUYgtxmdCnE1nfPPeh/JoLJYq5CRCZEBRAmzXKeSQ
U0eQpBgzqN9iCBRTspDXDPacRQkkN/PYs+iIrlVksJ7CNMD0mkpX5timU7VoK+IuvHm/llTafDQu
19BuXoFjeexFsERzKY3TgzraNFj+kmw6FUruDgH38c+nbUl9J7maft/BsYvPwoQV6mWWc8MCBmBH
BC6qZQX3Soe2y08wG1i8EtL6uS9EL5rAwCSvHsani9jYBnO/x7j949xJ50i2R1iJtdvXm75KQAmp
XZHYOLj7lwB7+udcUd+f+i1HsMZrpu+SUeCWS8+hYGommuwPhBVX3kEiHcLwhJwiTbtaH0L+TpNj
FFWsPiFHO5mkx1tcQXjRAe8Ai48TlrgRCT7e5B7XzH7x2MTScvRFO53IonfpUEAoZD8XkEG3Y3is
8cI87Dna1MODlHL2O0hirNwZFZlkwvhj7ifWaY1E7jlAc4fiHg3eReSgbe7z1yXh1wF69I/rMb3y
pAHUDBC8/c+6RG1hx7RRQAVpuZ5+6oIpp4zThfGfrcO/YILgGYtRwZ7o42+LCsFug5M2qbQxBvkQ
WkKXBpAtFcSZ66yqTj822YNWJLAhaz7LPmLnQXHQVN5SuElU8i3gVr3ofkCXmP+pbRoUoxlGBw5n
vXahouHcmZMMvC0Vdwvt5qsV9asjH+f6Mv4GuuxGcu95fVXhiNk7Ezege+jVYbSOs4LXeAzV7cmh
wn6MV9o5YqixZZp6Z21PcT7STNXIQ3ZYriOaUkNN1WsEJ5txyx9/RvkMTj2vPsv+IgXbGS9z4QjP
6GLETtzk+m8LXm215j6PhZwsRcVwpFnx6DBh1I5rRu41vXXcvMjWkmS9dgg62vwRFPP1gCxW0a8C
Htvsp7etyV0nfa8cEG8O7s+p1effDAmEPys9cY4rvT3Tt2cRVSIPTDn8EC3q3mNdzt4kA/tTJilQ
KdydOYmxfLdaSSlPFMog/nysvIq7H7fdO2amaE3yp5CWVX1SxZoBYr8mzzNVaUYedouDnUI369iB
SR3454R/p+u3kf0Dp1Xths8hBX3AsMbewMr4JHk4EsyXpsKtQEH6lvS2GgY5G31LFhr4KGjMjJxx
1Tolpz9dCSKTGxKIu+wMdHQ7UfSB2G50ZEQVKKvbuLNHXW5RJygJEYp907GxRWcU9LzuFu5GKE7U
QJvQdzU32xPpHh7CgUYAnhzt/BJCRq1I5ahkFfT/IJpUQisSPcIDZcdy0/pAVRpeQHTaTHgNqETM
AMqEMjyDBN1F0+Vkl6pgKHPCii+zmDN2viOAWLlkTzz6cqDR28bYX6jx9v4r+NagtidQMNMGLKPV
DzoF9VFZfFmxk/A3l+96DqjyDjuWEXRq0UooD9TDdDhPopvG06s6lcQnOrxDDEavrwmI1wqdgKcX
sVekjsJ82N3RcuxwpVeI1iveDbY4amR/2DYNyYlP++weQ/9hKZqiQDXBSnEyVPKX28PeF1pdA20a
NpPiAeYAA84Vlq0PEtfQBER8hf31IUmMFuJD6eXwLYBJtBXFSv5rtm3avvexJj/8K7vtaA2iErks
XszvyZIiSGLzqXFl0hvMDp0hMTY6uKAlq3/c21B2q5srgH5rx4tbZFLig8tahAripXhH2MIUEM5q
5mGQPM6atRMrfvqTavkvCTr9hyiRy84gVy34RgeK+TNP+jTecHbTsBcB3B4EjW2VaAT2BYODlv+H
g7hssToDbE9lMzm1M3pYUCXcw/+YqB7S/7uxJXJJtsIrz10mUA7PG+4LGIN71jIDcQ6jaBRiPvp2
EQ+9lck4Cs4ZUf2kd+pUfmodQBPHkEL1/Fi2RB46KORJGwOhAWGLadu9f475BpKlUrNKwMa7pYCh
IPPyhK9QP16OHJHsoFG24qQQhAC7dbhNVIw4XLL+6gJzDTbW8NXbyphC/IEiqC4x5TZfepK4eIBM
Igb0UrzzSK74aGYpuYqim1GyXzrd2qaSnUhg/x3Ib0QKJbAjXpR4rLpWgxYV6Dw4yeOq49gcVc+B
3LaRFhFHDlBZFaceb1VgSs57URdxKO9V2R85epeCHiW0CyTrp5ZrBG9QAUC7mY0CpFMtfZ/SPQHU
C2GVgBphb1bCQV4zjUR6GpNU0uGLe8iPXONSwiPtrN26gvxc1C57+tV8v6bUKuk+ng4KaDMaBmqt
u5PK/QSHVdGCol1SjVJzdhp50DZ1eUPwUCtePap0FxklZ8Meoyy/Zafap/Aj7bxAeaw6oy4zcqg4
UjI7bj77JsWSWnpAwwIaqjyCXXcNdLAuplcUIHMVPhiROmvlUTmGPerOn6AjRPYd2E8R6Ty05uxq
rjxX4qIk4BWQyWtEdKGXqHXACGp/Hk6apqud3hFMJi1gHYoiBdmZSKiVEkQkU+7HeC/oasmYNOfR
fBCNXFvEEzTqXoCcOg0CLdDvgsWrHZ83MMSLlQ7n7erQ9vaSi9ydB2HhMG1cEOK2OZ96i+shk20T
E2uLw1o2AxJpAPoJtdlnh2VkxsoL3Xu/u752ABcHhpFERkBEi3wnV3PDdM6cGtCqAkLfFrJdZ+Od
18M+dMwBUsq68CVCODVPpCidP/DWpryjHlB3pOjQEWGBlYKqtEF9rZhR6ziXBUG49Ko+OrFqNMCK
qhL+qFur2/bh+O1QM+xorPHuPWTk/FUNf89FJuNkmapJER61NXyWyC8x6qK/VwyieiWVDpPLCYeU
MYthF/HqOU6zv/h4JiftUwVyKCgQySrSfwa0yEu8n3Cvr0wO6gzpeBuGz8fezajb4BuzgoMADAxw
uLwMJjxzlycJyYsYcqxZpC7x3AeaxulFJQRPEHeATEK0UKYqzImCr8aKpancUfy9WtIPUmKUYC3/
Mdk1IWP0AzrqZioCPMSebkujk31v8PgfkXEwBRQHO1RpRK3Z/cZoDOdxE+9IMwGfa6QoSj1ngTw4
YrA+fDLzsSJPP+SQ/D6ajbdLhmk5hTKaU9W+pKlsD+YA5qsVYAwb558VG7l9gU36p5ePs93LeK5G
aQRz/dyQxWoXQ+9/NHQ7VhWglx6pO48QyhdwZH7x8b5dRwg6d1+1VznuqxBXUSVO2TolAbT43sl5
KJ6Pg93FsAM5P+8Ju0v6AClEQW43UAxL1TLBxLw6j6CLdjpYOfYDxow0PUbB8Ly06YUz3L1V371D
9b/6l5t+IYnR/sbgm6LJlfOzd57YLRqdSpLwQFIyzPxRUsBZs+ZA1cVRMMa5Puan/2u1wlCqFFuk
33+rQcnXBedHoJBjSCqdNQ0km2P6GAASktmE8rycNA6h5Hw0vLQ+M4RqiUmV4NSWNaRfBiQp1DZ3
VnoghLn6AyRzuzQ0Q1/vgHiAUzsCl9/sQh724EWAKQhRKmbPZR/FsVy1Q8ZHFbN1tw145OueonSy
CiKFr4VH6IbkUhrJAH+8A35qdsGAw34sxxOTFRagE2OzOchXqZjSbYWe85JG1qYtwW/VAjY13U/i
3my5gtuoE28Xaj+h3qlj2pDAZ2oXgEiyVqa1Ug/k+LO7X2E19NfEgSwtFTvrKM66at/1rEaqGCNV
nkfRnzLJ1H0Pj1iAnk95YO6ygRd5N+7BBwYzI1KYxsNXGZufpxpaplPootIpDojKVS9LXLUdUpUl
VxIBrFs+3xbwCqFToedGHD5LKXn8YHPdQ/Wn7ly0DbgYj3YoHFYuKs7onomPnQc2lbtFB1ADFEqw
FkryUCO0EjJ+wWx/lbXAMNVD0KnCMy6YsFbV+jYHUGLzRSvXxc7O/+PEOdEJjiSun1BMzwjWw2L2
hUogjTsDHMXbIxIsaSaNty+wxqgOGJtDNiAZmnmn8vUdIrGuJhHlwkLicwFPp5J24MEfzHdc5ykt
ZoPD/b9hw9+dITJJqVB2CjHCXG7ZrpU0DXfYq/vKEXE4ZhBoo1Xk2uICBIqNtTUez67KUnSlo7Fp
Ar7RFDjmH1kW+wsbXHY6HvAHnkBkN6C+hwZbn6M/4NXQojp67brX9UrAp0mZNnTdRtkq8DzsYHtM
oQQg6oE5B4/pOGqhOTVh6ExS+eGQ5AUkgMPu1RrdKjRbpN8RKYBy1eymywZfGEX24dMVnjvYFxsw
StNOFyNGgk3n6C5DNuD7AcWOHH3CN6OaxydJOKzdjPegnRIvpcTZD17JYnV+wVcudfEw3Xm/pmJq
+ygCA1UwCxh97hhv+nVogZlGIqTvbi9QfVsseY6394P4nlnwT43Js9MtkUmcM+11Nj5HEm6dfrZ6
/ald4KoODuHzvvniDFIzyHNsHItNvxXLjpbE5/kW5COFXWuWipR6lLrVXy9L8yHPI+nAhJwhVfjJ
e6FYI3ctZy5E0iExAwOU5x1A7OQFZrIqJfFasecS+mxgIxUdTuFgYsGzu2uxBsvA0fEe8W9U0X4z
ZyIH3hOAxqDcQYi/msrlXUO6hBEvV7Nm1AIhjqwob3t+Iwcj92jh+GFZ/PeBtZ92g/Eee/cuhwar
QSTo9vMHTWPZgSmm/g7ypbSrxGEVxn+R3SZvoyP6e9w14gPKW/AgnUldQFk0S54iuT9MMzYYekTW
T3pSeWP2STtGCsji3FqV+JGISFUMqADS+QuuZOf10ZZ7/vZspmfksW55hoIchZgezcR1fxPd7hej
sx+QIyjD7zyG9K1RgZtrY51Ei/9LU1qmKWb98Enm1Brbt1ZES4kguL0AFPIlK1xa0JTdfh8x2ILr
BL0znpgLUIjQrCURypBIAQb3OPig07eMEEii3oZbaahYx5EGVXRdeVwl1R/gre9qXpH4ylFN6zcn
lYI2eCqyT5Y4OD2bzBk8ExFl5rOyWlfQDxNtMYldp7XtcCNaTW6sb2pjM67lemwinFEXACCaQwcP
lMQ+zg7nfqeCUd4/XUu9nmC6irp1gn0rwHtJqUimdRijV+kd0jhckJzrSQ4gqkh+sV5FcF8WfXPK
igkZYaZQ8zLLF/CLYt4XeTcsaP5t0Csug+wRj76RKjcKG0P8EnMNEwDw+wYTHuiroT2F+PgQZIZS
1ys8B3KXVltJKwzAhRoPuuQ64s6otG7w8RToA/5DlJxhcC1LkSUYd/u70K0tXoPAdA/uNebE7wnr
iMPEjdN2zxz3M5jmflCIJkpXYK4zDyymo5/UpOwvOTaD6ysLIk5D1FC4eBkeW1T0YrfQYeAXInd1
TeFPobAUPECGmQpFnbZfojSlLRbp74UDIFWqbfX9HmhQRN9V1+fvcq/nqTI6Th03/M2uAk0naw/Y
3vu9h/e2r5y13gNJibBUVBKsraOkLo8ArgGel8WfvIcXprTaSFn9e2a7ke6YN43DmC8YpikYAmc+
R9ZqkZ3NXrHK+uS7O4ysvmiisD3nyYUItKcYZTtNlzIHQO1VAeVHlLwl1FOOaWY2T7/jxVJVjK7K
69ohQzQ7MCoup0+g9JeIEcOfA8G9L2ErIySqr3UJDgH11b1YXX0GoSB5hRyID9KKTrjdcn7gbfmS
dr3BURDmy0Dub9SinWafayLaG8rlLw5FiQdVgMXAuglD4Rl8Ur9D2mz4e7gAsZ1pode6GHjSJ7tJ
ENlnxS2Nr7QPXhn9JQlfcgQ333qZsWqOHJ1YpzGtorNjDJ//Ps7BP5YPX+yWFc50wxUn1It2tjnE
iSTCSDDhdZhlLuhfzqU3sEOVXsqW8XtBDLPc6/oqEvZmwC7Q8zU8ULMlW9IHiNGo6V195XUnanJR
TpJmQkBSlvc/6wS4exTWbQhocjGTCTCwyD+t4e7OK8MFHg+ujSKPH2eI3z6apWBBPk/D09elpmRs
U8KHvdqboXrsNSTSdkV05uoC4S8u6BmGAYLRXG/v80EvHxBi68FbYqn6zq56wbP7lpWJAohY8LH8
/S3s2jOoEYELn6+4XVjDldQlxOGLFX5zWLRSHFcZTiRkNvllpOwjLNIZ0OwSQQcHWigpnOFI8c6f
AwZor/6/KcBfBalyMet1yY+Yw8rYSy/OKtWtE3/jmpBdNQkDyaMWQVbedDqPNr/yqEB5v/9gyxfq
ntJj49tHb/0if8kjJMH/oZ25Qd6cqmA20f1oJ5QJw8daHUqQ48nveqYvR7WFljhaA6ajPjFPB7/H
XWS0srUUmaOsLGNiOHpvWJLd+zt+kQL4rp5zJfe/F6Sx2uf7poXsn9dVkPQItAWk5M0ETsP7QWSn
FqQzBQRnxR3Z26/QuNjz1+JeEPtlOhYOakkesy0zed7EKdl6829edXfoBA/O86InFAnJ/n5017CH
nHTkX5LxqBueoo9W764n3eOcJVpcuD3yhf9DMoC5OoNVlD3wM0wtwg2YbbF3fP77kXXPhWZR5lT/
c9Z8qvCWxvKnsr6QO2eqb9KFRSKsNeMyTnC4JH/AAomFjzTHa6X/4M3aXMjasvk9UIuikcE2t48T
euiisQhdrCtplEUj0I8Xw2b4eUE5ITnJ5eQ07UY/VhI2wAtaAEtScH1UdkLZzoVYYxwPP7zkeYQr
6IcThMwP5QCu2dKIXleOGBciyPaVAatHXlsxblX9Y4H/X/yVoEWtRln69UG84/uYEbfNgIHoLzGA
2dn+IC4wvQ1RQqzIrzc+ChKtGspbPr2fJ52qfYV7PXXMOSnYvQYXkp8plegivHxg2sSVjbWhLBQa
oCDwjCRQe8Lw3FA4UHAOnQfskK2PXSipZQPfxTdBeDQx0Rg0ozpb/K9Oi2StFTgIS88PhFG1ZgGe
jjDg4qmTuTfdXwcf6Z8F+jjvsL7hkgKzxtOtrIliEATScviigsAqDacKFHOMcpviiH0ZkvyvlLCT
6HsLHm69jZHMDGx55DGgDFqbQQfECjzOUp93tcGu95AiiaVcZNYhpRR6fvM3qW8pV9Lb1IAq142e
rq/H6Gla3OxMZqncia//2r0CjVBWOI+q6Nu7TS9bhq7sb/MNSmw1KmKiWNDOw3k91lB77Nfqnrse
YycC7gYjME2AQ7Uq2EVaXj5prxpf+MLZIwkOMFyYUh0ld6PXXYEndC2va8PTH/oij+0zhAktzNa5
EuGeQtUk1HGSRzyo4HnqPXSBe+cifz7vq6Fxh8+X3BfN5rnYV5hAKTLX+czrjQKWoGp1du4KCJ1/
6EMNZFAQwbACCRSdn3s4Nt5Qw5DaAoc6WC712nRHst7mAvWrFS43Zx/brZJ4391KC8CVy7+6WVM5
WjzGghyLSmu/+elrv6OE0uVZOaVHLMLAAZdNYA+l7TiXO14tKLyZ7p04+9R/QmFQP6c3wWH564Ox
1osbbPleLt9nNUB/kXJTBThLltBye+wibj1b4aiL0BNWiKg7TEm9MQAG7K4wPyVr7OJFq8GLAv0D
tvC0qlQXyAGp8P3YDzArNKPVHCMIq5IZEMWAJsV/lS+IOJ6Fk+Hrsun2sObJ8qLrDH+EqD8QuOO5
OmEGhugLvvV9HzPmAFipFRZ+U20LFvj0TDt2cbhHAPb3cFdmAEAdPoSIzscONoLVM+tztwBLTcW9
P3M1l7gxxLeVnEfGxM/bvluslBl+YRwiqKsTHcGSNY1udYwTdcVSbOt6WiIUaefYSHguEp8MMKND
JEYGE0MDtVpdcKn4RRESKMauINbo9tt+6kxBOmeYWMI+9+aAcjhejPfPchDYN8A8Hn55mc48AJcz
Nu9uJHhGKgBG3ydNwFXNF+DdIiqdnTCG8PZybzWzIHqqg0LkmT0D9Xn6CByyWOLFpI9ArEUxwQ9l
PVMLCkBIFYRnLkVXlIelgU9nnZqbXIhKU9ANc1ELL+HjgyycfPUrmqfnY9PgyQH6FtlyGgzTtDwt
S5xm77E4K5MFurGuld2odx3vn+EwD1RmUnyb2VewAzKreDfitdUtkCFM799YiwaG5++rYxIaAbZ2
fZgfiF+4kQW7Ca3+KABdNaxDuGWF3zE3BcU9luxkX72vbDU54tiynunYmf/FUASsnnkMBRdrqsp6
46nO0khjQ2+yKZZCwr4lu1HMSx6M4qgs55HkUO20MsxmM4XNzLAUKQYDoNcqgdNdTnnIETJZevAP
t/At/DfnBtYG/oxPzqYy1e0Ny9B3J3POA3InwlbJf7mudR7JxyjvaddiL4wth+1eBo6qFLUMhC5Y
ew37SH/XtXDtfWhNpyN1jo64632HOZkG45OajNAu6PSfSWmu3i1vnz/bdOTiq+X2DKdpjVzmYV3A
DLrP2fLVznv2bOJznEBu+2NYZN5PCtnPP0QoUDs8yIo4B3hajbkdPxpFy53II3a7AyTji1HF37l0
nW4ZT9X4EzVuG97qwwgSQR93lZtdkIZqjHIVVo95IizxoGJBYTJrS6A5UcGPjOwzflTMzTGPyglM
9+GbZHVg9pjQ5SRM66B2hscG7nkPphIKnhrDw0VQcoZF3L5WN9ccss1I/cXsmMiW8XKb1FToKVkI
IEjqUvteELTTM1FQxGqJMwoipNHZWB90+2sJ3fi1by4Au4NwfZmToobILWBtBmT2Zg5TYCo7kO2V
fQT0BlCVWoHkZ1E075fjDIY+EUB5j4qtpE3yILQo9BxhtG0EtRqE7j69BM7Isxdjs+hpQpajwFec
7TnJjHEvE9OvzC9WoRGlLT+iI609C5kKtOHUM17xdoxVtaKtoyuyDP7tsameMDyRZrmPfs0n0LyX
idKDdhLIPeTAJjs2H7pAqapQTaFBd0BrH0W1LXpaWntIucnn9VAJnoDiuQFPSHYOr4CT5X9+ATpf
THdaNUTkc3hnO+tLjvK2QPcDvGB4DW0nQ6QIyrioCkBJ/dm7CbDzRkoCEon3hqXpzypjeM3yXegr
/6vxZ1nXbBK3Q1Kswywz9pWXmsf2xOXxoj1sT8aVyfJdS/vb2uKei6u5aD848z6lKnWkz/Wepacr
Zm2esm6Aqb1jL7c0ZjZbEJAT4+0zx9WJMgJxOXzRhUyoJHPNXLfnqdaghjDuwi1LViPkrmv6yjmG
J0A3Osr4HpS6Mj64OETJEaNADhQ9Jh3qETZaD8oPpnfI23a850VkT9bqv4BCCDLId51aE8S3NLOt
wBU8hupBvOcWKFd1bNeF2LdRiGhCHKUdgr/D9xiUd282c0ppydP8vKYfssX0dtbJdnNOR3IBHE8e
BjLUzkABtBrckrgoGqCX7yVBs0rnZIGWM61NNEnQlsqDPdp19AAy9qLHhli98mzMiGbzc380A8T9
Ep32XBm7VvHogHDycMR0oL/Pt6xYO0pIwAY1jmQkkh3HtHl7pAKxJiV/s4wQTrWZsXbVaIhMYrY4
xrNSb7VZHG9ao6ryB94UGW+b6L/3XosrFJAJneGeLZnHnNxIoyLhMzMjXrYG/nQeHd2VF1YiF5es
UFl3gLgp8nlVu3ObVYrsj2QVP40nQALyh4NICtLWIU4A/WDKYjMKCT8NC79WUSO71knzgdC26+oB
P56DaZCBn6b2j4ftU4b4mSkcN9Lww7vHya7g3srXwvs8acu85c/9kRgAf2NxJYM2GQOZsf65YSc6
QA1oZT1fKPVMVu7iqfurFa03YT1OROOD7dowKHMa4k8g6S9hBPji2RYrQ2rV+GwK48Ggq0RbbcIK
k4kdo40ptVKGRgfMvuei8d+uzqmZ/jOGBI3yJG9Xnld685DVqfanpKUshHv4WGFeYT8Np689lr4G
oAVNcG4CWhVSPGtmOHlmFx9Zv32LDoCKnQpbwETLSL/1aQ7S0loE6zqJ/ucMWhzlslZNW1uzn7T0
Qq9DMMOhN/aTa9nYc4WS47cbYb+9jGUuO1kKFble9CgedMG6Wfe4dPaTMPYK1kxJkBKFAAJmP6yw
bgos0+ZAruPplj4isbuQ7Sfl3ukdKKD6Z+toZLVqRvAfRLLgDSxyxB+WQi69uzkpomAIt6YqQ9aE
rCUwE24HOemNbr5m672Gow93qotuyyjT8+s0iogPP79vctw81a5VdSN0jsiY6owClxYTrySdzGkK
bB01POoS6vKMCw/cEtcxSYZZ/8oszldRBW/XmhKIu2AnnOpH5t4MJ4+j7gF2gjpQQKDZ77095XRJ
IxbHHggYKPLsHv/8VJFBi6Ki4UbPJ/YsYRaNUKE/WjYBl/s88HCtJFdxc8dr3ME7Xk/uAaqfzfNG
tpReQvLQng3a3UaI1PDW+EhkQWE2i91nTYeIkAFrryK6jGJPQpjWUlsU/2zxWaFGx0T8B6P3jFE9
BkZVRQ6BfCB9BdnoanNkzFywNoyC1x0Svet4ta74wjwpwWQ9NJSffULoD9xmp+yfScAtz8eXLP/S
AzZzXvo5Vlful0cc+cDDB9TD6TSgEqPA8xhEawPl1kyeWZ3RFWn8O41mkD/qzAr9NvfsSAo/8e75
r5oG1SqeME/KiwI4SICzCSu76zuSq23FDV9+x0pMXeCXYw0FAKg3Ogm0t/x2c/xf5tjRF35aVqTe
G0OW4wrWDMsYbrJTQM5UnLBn7d+fqQDU+qVB3E2Fmf3HN0Menso59RxPzLkGDweSt7YruO10bdhR
FONTz3nrtWLmKI/TN6lZX1E3+AoGGQjU0ad+WGi3f24RWesHeBdTFeEcicbb/57zz1snxxlAlFst
xM/kKpal/DThSsxiwQ/abluk/Wv6mMMr4BimMgSvM36M1+8p63Nd1NgP3x9d4dIBAm99fq9S41WD
sxW18odHR81jxGjsH6Dz88jwvDqpibmlZ5szIKV1/fKN5W/q939pltuVFgPsgnnlD5cGBjiQakdU
HcQFpf7/OcbXB29VwC1qTZD1S04j0oOEPjFlHFqW/xzgeDL/ED9Sx7+PfzGNU3xQjdo5iaWrlpah
dCT576TRQvC3l8etq8N17Ud2S7lfXGVr1XUWY6AgbXbH9PhVR8dwcVNYo33RXsco14dLCYuPYf1R
sOhSSods1JBBRhbTPVJqCm+5S5LqI8XM9kkEad0IgzmziNpCFDKb/pvdB+4L6yzJYL45Yb2g6kBo
KNEddxu/vqX1ffMZt9qO8Ut79nBuayOGBWXDWTqjeIMYgJMJHRAhvo8AAyN1iFCF+XK+KhlUsN2b
zrMuTwEOJH+tlM2UeHcGuVn/PmXV0kLlb8mzeZ7S+VHsOqEbF+kNenPp177EObB1VEgyoKX/ZZvJ
CmyNZqOcsWJ5FqABvkQP41l29nDWkSvPhYnmh5aY85gH9sPaJVFjrnxlRsydlofm9yhtgcBUNlHT
nlk6Fcw4P2eQM8U5CtUwV6QB1eulbQ0yx/+TjngrilgPFUlDsK6z+M409W0xzOoo12Rsy16nP7WN
vpq8tMR7gxJn4S5XiU360tw1weFLi5vfVGOSKcOvw0sQKP2nJ6cUSBW/Vnkmb3WI6thowwJLYwh0
Mx/7/8+qQQsiD7Q3QiZ3gGSweJN+jCqu49XgTUA+KVscb9l/7/uQbQuOVzFVgbNJEosfxGeUhJDM
OxTUjda68WuNNAkoTVVaU9JYiwSDPZ5B8cXzqCkSMBORpvvgcQQT90bMenEk9Ffpv8tPJMZOJAay
TUtrrnnBIXbCG4BLw6WEMF7H6q1E4u9BBVDa18whJsG90xqp703kwh3J9gxT05PvqGkHw70XwErQ
Gdf+35a7Golp73aswu7BLPLkqcB6Tprsx9WitNPFDr2qYZ+wOobAZm4DfiS8g4KLeLNlN7X83Ce2
Uwr3CvgI6fCsBlxujE+1X4I3YY+vg1A3k4Qk2sfrPF7PeEhwT/4TRjoH5lb8xZ2U+WaDBNBhAwX5
FFSzxNbqKhvIiF0xpB8pJTg1XKjyPQSObl0vyPxzzOfWcqMPCsYNcZ9vOMFEQ5KGlrsfmIZMzxZB
JPBcFWXoQMZR2eYYA1y/uXufhXWf5Z7P9lXUtZIQIn7LPznwrq25njqKE+OfhayUJ4iJH6Rc3BxN
6RR5Y38Xie+yjaSjMVUBWnxSPnMFv1qL8SerwxWblgH6t3Y+4wqX+UlS1ThYCFQK4tnV+fGxtL15
FyBADIfQsWyiB//ImD/o58d2nKQ7DT82/ENjkK1TCifu0ycWLBHho/eM4/+ekoN5KKKValVIIW6F
1mwcmZrjMlXtnw6e6fLLbiCkR8RLPk3h9k7flZdDJRYF3dAeSZF7kQr6HH4/f6Zcuoy2+MGIyUoR
2zMNmRCLHNYV676GSjzavNUqM6LYzVBNV86VNrktcPxMvaaA0RdqcXj17PxelA5/onh47h6amCiK
WF3QsHgT5H4UjCriRhWq14HCOF6DMWk/npubMLSrWL6/iUAxXcUL5I+gqVJEQjpnDi49tYuLKXug
1icOcr8a5cEQffj3su6ccUjDhEwKabkoJH6UMapLvbhxSgyXOVjHkTcJ67tU3azsOekA9/FJ0oGa
+76sfnXx/OJ2DdgBOyiaPTBJ+ij1RvhYMHxGVoiCW7FBpvqBlIRY0DlG2kqzG+LXi+FeaH3nfJRW
XtH5+2YAAgyoPRpQX9aWRBhrSxWD1Eq8a4QS3J2vlK0N05XvktT/rzBTPbGmqhBAmnfQwSwKxlOs
Z7KemYkTdC+hzxWi65jCcf+Jx3yXi7Drru7EOXHJmG6X+hiJeogXZ/UQFmUk+NPP0gCB5Zr4DZsT
+WDWxz0yztPWQoRimLokvPSraFhNqJgOJUxJq+4NdSrnC66SsPhwvMuRQONGzcyrue2UPFCvNoWt
0KXs5in7TknYN0sapgcFhsgd0Wa5yyrxHBtNPde9JdZfdjSjemIjut0xfYyN+0qoBDkTHpwSU0KG
BbcZ6JV9TFE16jvNn67BuYXDqIHS6BuwTv9Hya0z6Q7NKjfoZ8onDIOu1etWu8daApdF5Pv3UQDr
/TP4GR84e2a1zftv5cmbTzeVXzyttDpnZzUAkhaHu/9aOh6HuZk4HPArWTutfEqTRmvVchBr322c
Qq1hoM5QakhQ6lBwZNljpYmlCuWuHOlP4FYHWcP/m5deTeJyG9HOKxgJpASTMBpOn+aoPZMTt+uc
pE9O5vS/Kdo6JI6/Hxg/sMRKsFmBBKCBjer5Q1QFFwEVnqpJZfbupXq19PiOB18biDydutK8JlqD
1xPbI+sdvJkaZE8jmN7wFHqT0xSf913LdM46QQqPHndiQQHnE4YVlFwRXT6knbcH2bH03ch2kqbq
KfbIk6dbQXp04Ln2r5NP1ypOTF5esczOMF63qGiIekzSxIeS6/dWk0dW/fmzO2nkjYbWZMF7N7bF
80IQCwNJq1iueJpz1b1k6dDPbGB9WQ1/Vl3P168Omka0HXE4BR9ZQ8BmIx8QFh4e7nDC80k6HB5X
J/alIBdQQHE79xWGO5+pDs7esNqTfDqqa95xd75TpWn+Nww0LlBabiBA0tGyiwMQBxgP1gUbxQ4X
X+pNeisP6kBdssCXo31BiUExX+EywGy285dE7YK26UbjouTZAg2nF/DGiB6l1K/FS0SK54KLGgpv
gxUnusKpUfjNl0gZo3932fZzT0eA2OhWi2mFOqjwYElNTzUpOlnS2M3FcQs30LYIDtNBojeKG7SA
X4hmUaDoJiC8H6CGIMfFqV6z/2huktaAHGrtwceWasLpQQtkNWFTpSY+0Bn1Ley4dIPz96kspWI2
KL4Dfl0IEAcbn11DkJFaDomVWE5aqSOUPspXbRiMfZ6mDlaoY+c0HMsgUxu75Yk550wfaee76yxr
r2H1jr1/KWp6FAuv4PekPs4AAWGteDkONt4UTtVCetNa2NSL55m25FkJGB7L0ZefhEofPCWksp/y
eqLDgnhkSE6XcDfj79jb2FzmQoZaSbWlXkRwQnMvB5i8FJVF/oTzNIghlVO4+gUdek4wYBY9r+31
XJfetyG/csGcv0UUx0dfm6mOljB1LXWaKRsV8/mqo9rqkq6jrv3h8vRixBYbpRIRrYf6MoG7tixH
Y75ykv5cOUaccAaRv40pWkhXphi0uHtckYqvFTomvfFUwZ9rxn9ZWReWiYOS6DQnIzySC4mbpLj+
iOQXJARJCLLTZRwllHhhEGvOq+uFp255ToFy1V1bTenmKXUKZ2PpD1VbuZ6xDd8fmhyBNeXDd0f3
yIGii1qEMxlcJXljt5d10cND/bpjxm3wBgDHlFcjlngRRzwGT1Q+x6ywxwlrsaQSJ5ypkhcyTRJQ
ig+pI649gfjGIjtLpRUiM4Wh7PbU8siaQ+v9DA87Ck4aM7Bm8al/tAmP6KcsnkFxjHiuJnWm5y0l
tYvgqwq6dW+mleeNv+WjNeQHxtKeu4gw4LXObVl+CgoqwWQROZP7ehGPIAlsVDOO+3zr02arK7Kv
MUXq9PHEtg66BJLiU1a7mJejRrmB6wGyUQUWZDujcmoDlk/pioF2T/zGIOAiSeLD/8ab16WSJ7pk
ItsT/blI3txtqWTgzC74fwrWdAxQ6PCRUvfRW/WmDhg6/ZwhYuxiBRm9kSgE/1Eumip3MYfzyjv3
DSxVFl/7BlOhjzmpFfSV0y9aUs1FiK4z0GAxlkOql7W5xJP6f9f8SXhoWvwwW2nfRdulUT7JvL3A
zlCMrz+wuOvAk7g50cuc8w48KYFpxkVdGP2l34RFSZgbNRkfIHvTRAG9by4BiN1P/O/+nR5lLLnM
CC4mr7cabpH3T5ZJ22tf3ngIKppYZODyz/h7ZP0n/otLlAujFH6XAkp+3loVhiXY5CJzNtNOr3kL
hevZNTEYlq+3kL3sYTXjcqd/+zPeybjHFQVLbes/6OpqGAQytm9vGl2gwWLBRjMFLkEqb/k1kdif
QM2PvgmBRO15bg7h5obTMpBf+l26mxqwF25nyMs2dEuBA7/23A5PepmBQKFXn2qEBQxg0cfNZTtq
fpbom8xbgPiXqi3d6KuAaWCeILM97OXvhJcvWR8qzAI1j2GcabfkcK+JBMLcybEfBF0X8wBEgU8i
istC847qLNqey+v3Bj2/YgT6Xsn5HzAWlGi7dKyB7zlYNSRU/5cP8QRW+hZ/2wqYl68o7Bv1Y9FH
Qz6mqI1P9zsyiH0hKuhBHcYM5NhhdwgvyNQumM/KABK7qsSCdzmgZUG6eqNAEFE5IthBp/XYZMKh
2L1mNr2Orhyk5bSnjxgu+jH3rDxk7HJ3v9QEOHzEAmCT52gxUnVsofjcq4FUHTPp3h1IU9xaZ19F
BDVzNdnl5qfPX6YhhDX9w0Gv8OgK9Zlomg4MIS3gAboqkNnncN7PDyyLgUW55ml8ay2/uA7Way1f
a6ti7DoNCsfG/K8V8d0r+6iffZI6q4OzQ1VeYvcnmbcf3myQYdTRcUFT/XLtVrwcfHDhhr8Y/yOu
k3CJx65dDT2vdHH8O6CSsH/kcijc7NWqItehgLFovOV3v88VdeAK8HNt3/nNdfSMuQhYCsiyNXAL
DVs2uYL0ND+TXdL77D3SUMtZosxaW8J4qd3KTXVw8JbqacAsDQlhyqfIyMXOkS3FQqVlDtSMWN8X
8sgs6XY2e73qgAXnQYno/ouf0I/O4jGJ/fabAQlytz7P0PM1ckhxguWf1u5HpmgwJb/sWyUxuaSQ
Ha6tjS6+U3Wv+2+o3BWDKpwRZoeneWkU+x8dPGsSM3eVEaJCKDDSHBqDa+xqP44AuB+rbR6iCBdJ
fpUpflo555NKCxQY9zwz4ckQQlGwi96/iGMGxd8XZbVag08pcXr+0CtQKNCNg/JlLTM7frhTJ5ls
yMQKbu1MjwIvlbBNDrbuvgzgQQJY8Ygm2XiEkIE9uTAppYDHj8Z+GTAChJ5aKEP6dqny67NVFvLH
7iq3xcWkXkeM+lTTRydBdORBdMk0yFRU5pwOl10PkVzx9Q/19MkxXwMYhU1nmvrHD2gUTp7tn0+d
sfvMZ+mn39mwqCJqGLihjo912cNIn2OKuwYEqr5xBTlPHjjdtdD3kz3SU3gkEuWe2b0qJD6T9GgV
G2AG7wZKt/X1aI+m6h1mJa7xHo0FsgGzoEKVLjnZ2Txq8fLewdOWH7JJMrZao+fX/o9HvGhYAq4B
2pbD0UgbHG31Q3rq5CJws0q5gifExFt6xswFzq2A6Ghjf4aB452RU2SuP1e4vYl1Q/YEuSoYyjm7
EmK2b0KXjmGwe0LzxgT7p4IkvzSGuuiTZ2NmW+K4k18aBmIFTwO0gLyxOS0rvRjdvx1hHTlzzZM3
HRCmZT+UHJSlNCoBmNTeGZ8rmeHms+pVScSBcRpcDDXmjvDZeHP7yQxH1tc6vND0q+rjmTNKZnMY
/R+mxn4j/6Q5zk5cr3XHQ8TLCL3UhJNlDXgzYEGB7bOZLCRAsZFJFdi8wp6/KDv8vPWF5YFoMZ7j
/KxVsyPuRy1v82Cuo6/+9a5iMt1HPKOhwQ4dTPu6878qT12itZ3Kvp45ndMfV4D970jWZdxbT/85
2VmqPYw1Iw0Kc1wYYCsmLUuy9Qwl1Os55B9AExTUik2nC/0nB0zaurPsNxWC68NfLbn3ieFoyPb/
cL/T+k9ut5kQcNvgJ6DCoe5N7abN0hmupsJBmw9aRi/OwkE9cWpM/OWrPPey65ei+of4m8pIwoBs
J0xylhd/asR8S0HSUMVHctIctkooDbRpAGcG23wWyz8uWIGzmZAfROnDZxPzHj7ZiW3e+wsTeUt8
9fppCG0dyvbZDF11kBTs3EUFLROHOKLLX3TAT1UyGAPRLEaLad0Qfr3Id/bsNVD7opzPVuhS8UkN
eEUx0UXvtppdFtaQU6N6Gqtgoc0E/tXViUo3+ratABZXI36IVWlM7Nqwi6Vlzf/43+2gMmshA64a
lsznZLohtcPuT2EBsy0t/naCZtRQAdcrvsbWb2jBXos/Kxnyb3yVanR/DAXiJVqFs0nDWo+mE/Rb
MTfJAkHtny9UCjya2QQ/Mn93nJC1EmKw+5GtGhsVTIjYLtSU6ICp3bww8od8AZdErRinh8GorONL
zgpUoZAoIyGX5PmygcuVKClZB9b6Z3bGgbaeJgxAAkrCWlCHbHKfR087fll01I/XHK+roPLWTfWR
654Y2lVD6eBqc5HoqfSUEHCPfjlFuYGghPucDSzwBsO6tMQ/JQaWU4QL46yJ57TqT+biPKRLv+ty
EiWXecopqcC9ahyMirvv6kvTta6JrIjV6mwRKB5zgXy4S5dkcj6gWHEFjIdwhgtDvpdzNtsmyJQ4
M0m7R0W9qSoW4fHAU3JF3/SVUjYDdvsOOFoioJhEZC+jLuK2g3w7d4zQ34XNJdxD61C0aL8A1ad2
j2fMZZo9fhSJ+Wu+giDNgNyYj0bJcBCx6lekE2v7ftoN5032PYbxgWOJ+793Hnn+egDDKx4xikkS
MPzKrk+HhGRIjiJrThyTthHnT1sFwByVVY0IDq4Yw9A+LPIt6h0UwtMNdvMjYON/2yDeHvhaEqg4
hHXb6x+HlTsrCooWQMqcUbyXZ3MEvi7lQjrezuzB6V1Hwhq4CdrugzAGZ9FCaGJ/uuMZlP6oJ70D
UoiUb9/McwqAzWv70CODa54BeMNZpLUwEROhxCWtv9S8MKwNqteq1XR26Z8cDCw7lOZhqY0iDWdA
307LBtC65nSgH22IIHC5otUihtX/bXEcJk/GhdBlmYbMeWPBF5DTPtcLss9nWhWAkj0vVdyNMRdr
WxuQrVpX7N61WqW0/IRP0ATqyGICCqqVpGGTMEhVVqVdRLNFJOBr5DDW6RnEbK4GQtnaz9wkM+Q3
ATnOCx4jg4nnVDkjO5trm6OUd4gFzvzZu0qTHawlO2If5DLzvXGXIOyXgOEKEJ29sbVNvViwJvq2
Fc5CrczOxsUHKdOgTJwpktlH8IHyO3N/V0enXr/AB8UYgoYI3Xg/c0e7/yiwX7ccU+aYIY9B/BCT
ruCiOoneuhUOWWLt0uwnJG6H2fyLbiGCDiOnB19R+Y6nAA28KZKSq4oXqRDuhg0A4gDdEYVoFZyq
5JWdIXG+JPHwH+x8aEUkzB9VgK5Os2XHRdH3U04cGrdXYlXkCQ5nd+w7UsPxIcWj3CdJE270kZF4
2fjHmtiXM5mMXkbQ2r7SUxxhUfAFmonKxhrOBX7HDIHsQMFUR0rtGDXuQEDLlS4nVLh2DPs/eMCa
w7fENZWv95B+sVajYuC9caoEWDmV5ce3f2IFHZA3Qnf8EW4OVAL6huqyIFqdYxDvIbtUmQgTtpvK
xEGGCwlWGAybGfKxgRziuU9JlT3DDkE5F0x86lh8Egzzgg1bGkKhvJtQ2XgYCIQ9jvnWSUX/Jyxm
wooMivlRkYolpA8zBAE9MTKDwXR5Js1Br81CuyiHTKBBpYvJur6ZynqL4Kpg+iLsaX4uiHkAQeFl
txpCCozUYhxsZO3rcK1bdesBNcEXsDA/32KvmEFw+97oCHcoK2dixlDluvA9dRJN3ckX16KGAp4a
/oGdGctul3WAaOrluMh5KOMPh469s7WNOaY7LArgryitJm3S6U/9lvzgkwE3ohu51v+qs7uwycx2
961aZlVUP5F7vloA340ob490cZzD6MAzG72VuXcHmQbIY90ReOQz28fClF+z3BxWdSwNgcUAflG4
dCoN0EmnnkkeyUV/hiIAd93W3IuN7WryCru7WYDQfhz20SrfU8dMxTW7MZ9IsVnBiQz4uBHIizdk
u7A94QOYKMEynOGidgC+IkdQBJkWapTXb3GTRh15B75ixpXF3rahlsY7KOu2Rhj/AmOY6e4zusuQ
dZtDo9XWK4bag+FNJq/Vp8oRZlRy6gkruYJ86eaEWw/5fCXTSJm1Sx5kD+bsMklRY6kECYA+ogB2
d0V0OuZS0tM5P70K/kRyNYpixX/TKvNgC+n2dRSxhdv7d+peCtfLCgvpJizvCkTcQk7AomDA/R7a
kC6X7t+Xxh91vlmYdE1hIYOgJoAMkjrVVcxy0EG9qF7LcwhPOtnou+eju54mPUB6HgoIWAzegiT5
k0gsZKQnAUvCRMU7lGu9ZuMInE2kvcGByLnjp+smsNudCSA+OuvAgjhDYd0YkSI5gCUNeq3H34DM
tCHdqQySwB4WV+ilKAzCcIMj2N1I6tvJIQZrZ3mQx/ic/R5f3P7SiwEe9Mblq9sOhXHziHilWYpG
U+RDZ/urI+Pbwim+7gBkPa6wRk3DTCp8x1W4VU2AnksNiGyA5RceIlsxyXlIs8AN7AKxSzRdiAfm
jmMyYy9fYt5oVa7gOM0eInHUssptbgsBzNOCA0h3N7j+8y0w+0Ls6Th241NXkxrfPfQ0kHxSrhDM
qS5EzdRNIckQ8cpRoLjtuzRA079F5GbALHWkwcBZzbzDxC8ZBVrRo51qdKkUiYnfHNYiI7nA3Yl3
cwirA2VGbRJtcgNzaym94vwhy/4F0xFrUQYVAvXDRZabHRxHDpS4ASPjqoX/0GRQgFXKLzLPTaQt
S2A2KqBPiU2etBZCOR1gkx7QScFu6RLNd2EP3WoSPu8lYh5/6YJThzrh2TqRKN/EMmMHRkfP1OxE
dC6sSOAq1Xu/Mp38L2jXvr2+o6/p3YXVA9CbmFb1zjI1553Xqb9k92z8H6Pwcr22ODZ0i2ztvT0e
CltNkjmxAPqMcxzejMcaPr7llsMs8emWmesJK+/LorvVEWjsrRF2Uw28VHjCoYhop/CCi2JdEX72
qA+LezlONLlBAilWDRZND9u+w+a1+ur2Cq+DoY/dNNv2Yb/+rJIjcE4BU5dlhAQXWIjqG5tx7O5i
LQwRx7QfJCTli7GtbMiPJXtLAh/Twcv6UMC10T7Sy4dTHkqC/doW+OYrw8ZoviqUvP7P9vRvsxtV
i5K3KEA29G1SbCQhf5x3WOdidR3u1OYBUUofdslJpMsFj3QTMqCOUMIlDw6xvslQfDms2R/QBaXE
EiNoTvh4z6cB5B4dSk0NDEJdUIP/9uFh/81vk+ZY/BZjrDMjORSXcE1kzMEejheppCix0NpHQOP7
Wq41BFX6c30hXxeLxHGTsEthotyXAAkmGOqprOBHXJ/Hl0JcEDyuM6zPiDYBGug4MNgeQhCrButC
cOdC4RhkJ4scMU/G0O9SmAG8NfRRDmKOsbGP661420CI+EdxMvZFd4e379hsCtKrMdO8hPgzAhYr
2rDWIk6e/kxKbynb+SsTxyYJmXQFvXJ3/SPyMjbOgGQNs/Eb6JNpGBC/Rt6E8ndsMTQBSshnV1ds
iXXpjXSpGOaa041pXK+AtkBCWc/nCJH1Avyfhc2Q2asJB+KgeEV7oWQxGs2gvOCyEMLl7Zngh/Gl
HaGLrXfoqxwhADZ02s2ao0bnOopCMhdUHpPGebAPDgRUN8cGEXvIcqKRcnd3NHIHFfj8eBhzepFE
wa9W1H8ESaD83wb7PesJwxM7pP3HjHA2qfaSfIE7JYpdIwLd0g1QqA8KuvBuRB3dYpxvcjvp6B35
+60V2szA98ouMIzLx5HFlixHoMoZEunzeOPmDWw2xup2ADNTUlOTPrBxTOXr9WNANOqLLLTWM0FQ
LF+fmxy+kfppAldTsKNdF8HBG/lurv6BFph78F5UJs2cgvrxBjgcEt9aL92f/tjKWPZZ92zy8cjW
eoRza0xymlptJZphQyx09Gq5slSL9phnY/RKwhyDzuy5sDRoLGzvTn/0s64XvWDCUZxBllhX1hsC
aWYdoJHZsJ+dl4Kf6ZP81dslCFruVAeLI7xQ90u16cU6BY0EKQKvyIXawa07CVuTAWP+09B/mKCQ
O7CNUn+UyWiCsmr4OBvj/XCfNULV0Kdq0t0ANBFrlgEl5q2xGAMWo96Q0SMZf1u+s3Zxs+xEzQFJ
vHkWd2+nmiDzrQdxg4PKi0jejdaVs0AH19tuwjbkIQVWDP/WsIGD6PraV+yqFN6nXan7Cw+EkyjI
hwa2c7JcQOz9KTG5ZAsMDX5Cu2zb6ZoG0qcH2nARvv/BDeMgPLQa0ePXultYO/DJQjjqtIOqGH//
OB7xY+UPrB+phGcGxQ8R00/m/Jeiq4dED5rFexAJMDy8r9GqjSfRORhJ5WXgGkqPz5tk+qRRikZ8
jPzuCEQq3Az4jBkKJq6WtGjRBSS6cVniDbCZN6Dgl5okgJQUn4p/o9Q/WyldQRCeQlHXImgGFqya
Z0pvp/NfV9SvZr1h8Pu5EuZNsHb4YslxfiD+pr4rK9EqPY3lTgUILmuDXdxiKxib4Q25X4O6ouqt
vtXg4X7DlaPOD9zIGTXLyeapJrP6SJ5LaaFUN0DXsrhR428XhqtyNTk7NS5EjqstxHsB4UkiFQp1
ybXklPXCqVZ99mc9PtXdZZ3jC/cAAuQC9RMfoK6D3xU9N/Z5eBvsbBxU6qTOac/Ir9iPPWOHH3h1
84UV704NHEtF4kXJTbdc69WM37WHyMngXdJ4qzfjjLiapfzVky+Q1E7zTwIp5FExf00oqn+bjhmB
docddiyxeRvxVyISmeM3iersnAiIv8yABNwqri63rU20JQKBeMEQGmOL5Gs8VvZQsZlf7ocs8/kt
5Juh2zlOtwz43Zzg/H0IWTypCPsus/v8F2En964/sozxXBxs2+yKkAttk51TVWkZ8n0OJwwEB9Pe
gQykRPlQVwROpuYL1P8gHNwsEEJKGZRfUy9aDIupcK8kg4Uhiw37dI2wHLRZx6hfJEWdiUUMowaH
5BJTKK0yHNHjRVN+YMzGUVGbRbIJxJWo10AQTr7rk13XPQEKpQV4vPuk4HaX0G8KvrhFBFrclLaX
fwKKuMW5UhF/OTcYJRRyoi+RP1GwW8zq6NdYm1XcQKNkhlZq/un9Qxor+57StNdDSJA3X64xnUbV
FlrsyLVEgXdKKyRMwFOoI1JOxntbewXIOIfs5XPl65eGX/bg7pZRoINNrxKcCilJn6bKenzQYT4T
/DfKbfKA0jl1s+8uvltfW/RuSy8sKtfIk/K9TV46ch9Liu7lT5BlxVv6jyayRTFUat1vYU6SU0Fu
rMcjpeY94nHVWHkiCMzIdKdcFzIdijjETYzBgR0UbmtajR9P/ggCu9OwCAyyaFU4dlUOMR54xyNu
CDes5Of8ChXI6E0hSP3hHhM0DrbXGvBxvFO9iOtMBaqdAE26cmRngl4+PSqNQG9cymwSZlCWD9z1
OhSrb6C1HRWxnrY15U/w6wrm3aePlb663USKrltUVE7qxurPj6hLLI3uZ8MWcT5vjUIBc3avUs7p
xfomHk2wESUlk6iNALkWcdHLSaEJw5dqSX179TPMKY/91VAXGN231+8lnZ/OooJ92fBs14UUeWr9
hfUcCpgzMuoOeOCNuaWneT5Gzx+R/FuuUxuDU1/c8BWIyIx8lgpLhAgDK0+QiC1Am0svx4epg9MU
mAk2hIHW/EeR6CGwi71avHrD1SXV70x7ySmTcE7yA/VP9c7aPVDMswWIlqnnX7r7o/SAI0oMwbSD
cHjlQkR111GwvkVRAkuL6r5MkU6SqFdKxLbc8DWrz1gH3++5b45FFAdtzDyBuyS7457lWrvcUSjo
OSl+tQkFkaCPl5XAjVnhyPVyKD0ODUQmpjTft0CWrNyCiCb1mUIv/+ak0EvVCKF2gz8BKwtXPXtA
QtAkUnqoJvB+Z4tdVRrIvEXYPd2f6cPG2FcfQBGponU2D8MsiEkwYSCJ6M59mlE/GgXGeXBMFf9U
4M3koGDATy0yKwmEdRSxgh4I7um4p/b9xXEQdVBwkqyYMij56dgevE86fY7Im3slLU/rV3GdT2sP
ftbnm5lKANZOi+JrlBXODMMDiKf17PeXcWLA18DwxGtKChF+Q2IMlqeNzKY7C+N86/+6noKFzgmz
6e920yYhpidkDHMw0PiMAPtg0oEdSMDXWKRfzp8qBNpzQtL3AYmrZgUeSOoGCvZ5CsO72vT29XSP
yy3qgbPiwTXm26ZuuOX0KporZ9oQIpVEO0utcqMP4Ds2jX7rNazwILAnIkDpXFZVedUOaF1gPfeh
KMnBXxTVLixih8RVPk9EXR+0XkzKYhfABV+5qI7ZM3m/XrKbNxMSazsEXnDzp92O9SV2WrBBgGf4
mWgs1lF0VGKGXSQ/j0UjcPY4yHyBLpqMS34XMsPz/QtR+dra6nWR7KgOxEk+APlTJqzz/QjZ10N8
h0M9HvMZY1XI90PaJKYQohZoYu6h9ynlC2Sr91nUgycdGBuBjuniSfSsiavVWEIDKitnCQ69QIgu
+2QdTz8rglETAx1qSDYRckMQU+GecYGsFPcgL5YF8ME0BEC8+cLKEuMFWAUZXjNJVUmUW5dLo/P2
dQbT4nNYVFSYgeYNsR3Ea52UGFUUE0UVq/3Q7YS5a+xJRc9fQ54kmLGVBZhCaNUVGPZlxsLBQHRK
G/WWMEQbRB0vEhcB1c4OzBew6vwrQCh5LNHLqkW9M/Z4j6h7LNd5LWadfj5sWltcNPdQlHQBqOo2
4jSfrH942EOLb14ho80lOFFHSw9orRW5Wrd9Giqfg1UM47xokzytzDJ4rMzoAfCumsGPYdXShoqF
NMm7dJbOGSWC9tFfOiE6t9CHNxbQgblH9KAf1ssNW4tdVioJmmLTT5FMxDYBwucerh8QePRrCQs9
LGcJqjhsZ/9gR1X1j5L+KWgoLmsLR+jD31kYSXvLLeIemB31megbDxhoHNDiwU6BrmsCDDcc9T25
T3DQUIZ1dYwS8P8xo5VUbZ5Bi9MeI0LPsUMQ2A9O7aWRjWh54T8RhJ9t+I6bpiQnsQmUl8Zd5acY
1jAQ8gT6XnOmM9XSNwIeXPU3XTOya05ik/wfzfUUfgofmCqkvdedKso9+ge94zTBRcOSW3bPwbI8
KE1yBre0Cgz0zAy1jFiZmnwPLuVvf11I4JQyc8t+BLZ0ACQ1ynUmS62Ae83lV8HT7BSB4Sct9MJp
VD3tmp7wodaYjyfAOqLkMBTq+UHYOQg2RmJELqXrJfFySjPeEwIptq9Vx0rmctjGiukyEYYpicCf
sdKl0RDKDR4BzPgYoagV8IA+eIK4lAWYHVFloUATndRQfw12O+DyctyGhE3obzaauhbGTM59xSpY
8bEm08iWAalNKRnZoYDAmCRbMrn05JPL8tTN39pazsUF6mNaWTG4u5//FuiRXUOh1gX6Zrr/GVp2
yt9PX+FXtSfDpMcX13ci+LmzjstCQawwMxA1+Lcpon7x4UL+5YicHhJ4sF6R+Ftq+KRNe9JIJ7xz
XJu3UbOR1fsFqj7bRmW4uiWW+5S3BCuTKA5NNa6NM+hMuJOggwSMWqjq81B1H4dG+g3UH+g+5OAV
LCSoEbp61P+zAWEgArQFiDcKENu6b5u0qpDgQYxBYLG5+vFVPtDmAFAnkU3RuxDT3p4E3G+C+9jE
1lfnU6SCuEbculo3AivU3+Ckbhj/xgLsc30Gpe7ZiWtpAO1P+EOlqx0j+42OqZv4XYmkcCu6OlX/
d9ldZvQvoR549IdqsW7zD1f2cBlHe8ROuOTkuasulv0x8wsELmn/ihlfFLozp7tF7TcFEpc8yh+g
LRIbMFVCtQzUhlmugOoWzsAVmfOGsyFiEcrLcIx15bfiqiDRnf8hGBZqTYLgHOv3AD4cl3Wj45pR
rBWz/yi5Y5ozkFZpXTwhWmudLAgFykrxeAt6npvV0yPa7guIuujJWIUwpvb+aVtajUEGrF1Ycb4W
DHfcjsEoQ/eyi9RYbXS1/rLbJGhH4v+cHO7Y1dMvXhpnizp8IBomp2r8wIRuhfirhGk7pBeow2Wk
UrevKIVCOMVjp3RzeBzCBjpgREoO51vU4+8vgl5sxLq8/EQknvl0UKq0kax8U+CuuHNuN/I8uGhO
FN88lsSWETMKXjXzdRS3Y9E2oPn1DbqPGuuZxHZx0qWJzzltUnyiZZFWqRwZ3Nnb9o1ntjEF0Jvp
Gl0lRFqYUeNtSUtZOQnrredi7+DlLyWYyOstutDy9ctaDkLgw03k4eiVR5vs0wZEdDN9A65hx8uI
l+GhAD6ni/X0872VtznTk/ztJvVpceEH34c96j1gt77DBVgIdBPAYyj5flAIxcWYrOv8/ntI2lEN
ig2CjKmEUSBzbmAZqIYQJUAQC5WVr50otRg9nlOzLAViyfW7NQr8brGi7GrBlwJPOeFH56qcLKhX
zgOp8bFOvd3fendKAsvRQJDCUTC4WwmP/GiocnojECYe7lu88yj42if0lVFpP/3rmHAdd0brCMGq
9PjatdsFm2hJo5fH564bPRn8U+RhxA2lcyYzFcs+lZKGMOAb7LHUdizcsC/ZFABLDuTffGWxNstc
QnEAKa2z6PjTLj5XUEhIrc+V3uEBj0TsibG/H9yr1KesI+vvIFAu8TLu9TZXtRexHJg+9Mv5WT+m
i7SSMiJjmpYKV+t7gnd23s0Z7k5jlBVG4QyFoA/03tbMwvJSUOFqaPFy/4EjgBbDz7MJN6QaJDsu
dGWFWDoYPSHWwYE983WFbHx93c7pMhLSbFuuqrQOW30Dpb1T5ZQGKVX9IhDu7S18I3NOErytMSdN
sXDO1Bi9GqydSC+bIjCzQVljrb1tWow8u5RyoaGgcb/VBpRHuSeXNARR/1B0w1IG/ktM0jf4CrjL
gFf52Awca4nuEMSCBm4eyNsYfEUNNOYs2b9p7hp6Qo6BCyTzYZkFHIgqi3WtOZmiX5rlMvJOicfJ
mAWfmxuvza7RSRb/HPtxP6z5UeIBP7wpvwzEjqWPtJDYyqefxekYEpgfxc//Nt/7WNJ3pXJHPLPv
vmZwyfxf+wTVadGlLjotLXEKK7HweINc8eWB3Akl94vzh2HGqRs8SlRurz+VRNDJV6oAIzoUexV0
kDJTULfNiuWwkvHOjhxgrabBhWHx/cpjOIiooqbGkHzk9azKntwLbcuiTzf2UpqgCzMggJXrTdLs
RQJA3uPste8X8jfzvur/HD8bFAcmD2uKflWEUrtpPEsEnpRsbq8eQzPK1k+ogzWN7B1+krBJ33Dt
mZ/mfEIYQQxPJiS4Qa4kmM6af2f0++qJgtUfZeJh/gYZTsI2Jf5JdHNYfIt6nzdChXREVlTUZgSM
oQqn17PofWMbtnkUqDleeq6octTz7pbvJlCUbew4fNyeSmK57RBYjhPJJYijqbGpvO/uPR4mfQZz
l8pH7HlJdBObrW4hw5aGv69e5gXkU8dqz4G6uUaYv/T5h64QQjLiP0N2hwlT1gpTaIDO2GXqJQnB
ObNivlCzkbqVgt+Erexiqx+bEk7zmMUNg2JWXx6XBXFUmPqnFTUFb/RLeezkEzU7Is41pNzSwzzy
jH7VmVNQ57HCQrmdzEbiIsdiC00EgDM4IKqBQ4wMfurahLtdJ7JBeWAQ3aVE0GwwlT+MRE9QlrEz
d9y+en0d0kwR5ZcSLa2FVjppMROc9kTaVU7LNP/yBDQC3kgrFTa5anVLZx98lQwy8SgV5gWganqU
/rvwtEfiEqx32vZjlXpRRHaYjYd4cOt9m7CVqBX32/6eFjvFjO4uxAxcDmTRnSQYHPCch4ALgND4
n8VPUBj1KBDs+o4/07d/MoDWsbDBeoFCXEpe+dTmltA1OCJ5y5W7sbZLJbYktDKy/aclm5SZY909
44wD/6R0FirNlb3eC1hg0mhO/UDHq8KGMoPzBp/SBkaxaNT7fv/ryj3JiKynRVROvsxUulHZFPz1
wFDwZSprCXgi1BLxETqOhJwNVDtDTmqI/ZN7ZKZcMzzFghiZ8Zdejt0CmG/iF4iRRqSqwz/aAjcB
Ohdp1ksxt/t2txAGSj2M0V0j0izLGASk/PxhZhHCW98y6aQ+I+pct5sAyhUmGiP+Bpa45JeWFBM2
9kLyV/YboG8YbQpKEvToau6qtqMoodufFyJGCupPLWYus4iYARkO5nOp8+i0ByJpeI0tpU+AcK29
EzMKl1xZ3YQzyrWaUoXJYJADIFFzpUcrOGvurWaILD6jZPdrOR+AyZ2TsvNBkykaTUefOD/UUG/s
wNFp4CITfMnVbWRnRmYXJeZedu1ANoXvgH0PSiCEbighImblJMFhekgmkLSAwLF1FeF12kksSyuV
EyeLs1CfSyHkHtDLSj1KbC54ytmo+4r6MiBLE/nPKZdReuzoP+QUer5KacJgfmhGeMktdMSxqusq
8XQw247Pxufo9zzuYioG3WkdGekn+9IExUnBzwX9D5ZtE+HAaTOyNfNla96rIm6z8ELTtwgd7c0B
4Ib3rXoATbK9/F6Noz4s82urZUEDY+bSx4UC1cReaIuT6yKQ5pNBvhnL+O1cthBu+E7vkAaJfQQr
g68CWSVBKIERCpY8CoShpWyTpk9nxkJMJx0kCOoi7QIkOybmznBtxUzprJT/fkXmTf1ypbVomAog
d7SzRmH7vD15F8tP+60tZtU6p3CWm1WpXzAehV1nTMxLOSwDCMelQoz3nJCAUGaUm5YcrJ8hGMa9
vc8hYjUBeu70fYugBPxIHYVBqqcX/TqNdUvhqWmuLdrD+1QZIK24p7j9NZ+beybBiA42+lSKV4xu
0OX4QUihJY2n0aOldpDTQpWxHXT4fhtUnp+jVLERBrDc+sDTfKod4ZqfLE+YtVqqru1aqRc7lAFl
/SQKXyr+fwl/xJvpIs+C7Tvao+a1fGtzlUnerfzLJ8r7OMIKyP6BCnO1lsHxu+7JxpejXhzw4epv
xdDt7GBxQgw6Srm2MRb6AjJLZuoGxCoS67+sOErBSN7WlP6uz13khavPQRHtsQ/53zMBJmcu/GrW
CjTUBfKlsc98YsfW+1JmQO8HBL98NUbaP1ec+yEN31pgItRxeFlDTFYmFlMyKNV0zQjh7Snd0VI+
gt8VDfmL2GKRl9s9T11Ki3rQcbZmBJGlDtLXdSkgxcDa5sEe4eHXTM1vFNN0r2fvTQgBzj5b5XQn
gmRt4UlJfU5A7VwcJVT7qvvsxq+URfSSzI8mAB/RO832E0t30XUu5Xx85shkTFBxF6K5oz1pqCHV
uOqktUwsWLuDudDntiiOjMKHwz3Tc3G/pzIcGGAFYT7fjVgvG2jdNmGMORcpAi8QO8IhTPW4R5MR
vpoEjVbbJeORMMunYLs0knqzVC2uucOY7unGqRcov1yIgpI7lxQle1gnKL4oK4Myfiw5F6YsNtxF
/2RuFdReUPNjw8WnsAOkvUzzSchOkHVBc9CgkLmyORnPHS91Mf+o5bHsPUtJeLT15kNVrhHMu1cX
qZBRwpJLfpR4Jp6vwATMJHp7q8HjKYAfDqHpVXHgUJwNNke6TjiQJMVCaQQoy8dKMEH3tcfis1R8
v3U24mgCst6/gDgNhs8CRIegGKgg7Dy4DFeW0BPrsmue6l29eLU7CJMPKE4AxbyVg0rczT5i1chq
9GZA7E2myRbSH8Qg5tH3aHtu56jLN8499RoWKs0obWa9ueiZd2OMKTkJE7GOw0S+Fpx1xJh9SYuG
9NB/lPlZ5knOB5iJq9kyyoZ5wf1TPCpQLFbLtcLOlbiQqu+ZTQSBgrCen8oyH9xuycQw9jY551FE
WqCphXoRWuxZGwAbR505bbpj5qNia4l/Mo15v0IWFpd8jEibLYMaeZoMN9l0WSFB8Cfp4rXfUx6b
MSz1NRm8EQIQS/Djy196U1Jogv0oytdllBA8OCZVeWPj27XyP4cab5tfupUX630LsBzLh13UmHhB
lGwQe9iTEJkTr5OAF5S6wGRCE/FHoyc2yY9wi0SmhF4fx0J0bjZpEUIkV8UqQ/AU7Tdi6DKpu1QC
kiF6wEMnWY7v9t+p4y+oLWxXK0OGF98B1ZlLuIqr4wU3ytsdpZJdpBHKR5K4rXV2kPKHa6m6jXlM
Bj4D3gvIwNA39Zamzskz5CAecoAGVJsJrM5cwsBleKYpD4+2Uy+64gCy0InCgfoWehfglN5fU7+1
9toaNVapWL4zlCqXa5/JDcPXxv/llZt/jwOdnu1SUwGM8qEecLty48F239Xc7qq7ToyASha+tbcE
DR9FKaRAaCeCkGZ+mgtYZ6bElQ1joTF2rSBlOxBarQY03/g+O141xMtddQTWgaEtiJBMwmUMHOTN
XnH3DRICMVkK+0b1CD0FdQWN5QUyg8hLyQqzG4xEcju5KZRx/NzR1RLbfP+u+R3k8dqNmmB3vOwO
MjTWvcczMRS/vshz/raVWJyVQPR846409MgveD0YrNth5Ww4+crvLLwy63iOFTexG+w4rNf9najV
aSu3zvQhpxA3kZOANObRR05afgbCZlrkyxEPDnGKH/jCozgk87VOdLza9wq5fskHuYx/NIvcECpP
O5vs8vAGDC6Up8QnieWztMwElzJUxnoCkukdR/+lim/AoFxZFQ+/yJEtP8pNqCoKDxOAUNDfdF2E
Day4ENgj22fYzlQ5ttaTB5QJZ8pFXrbi9BQ9hal+yCSI6RRSNFFpN3JppIe6nhpLkaOxkq80Kr7z
RlCcloEmy6sUvfNd28lCfaoGmqupgNSYIqEgFZyyWIyh03WebEKdD9kjpbUyUcTeCeiVmj/ao43D
QK/xg+tQD4lqGAuXwgFGv/hvVLhjfeBPMe3pOe7kAnJn40sgteeuU7XvFuTZh0pUm2sSe7Jwvt3R
yHbUzI9fDLoPqndXeOUt6k3wDZhF1cBsKUhBzKqvWptdmqoVhqn5tYGVmEtpZbEeW/t7LbdkOqgF
VmWVlpb+lPaxU6rXoqHv6NBPrklfd1Hn99tHJkkoiErlpJw14Js6U2EJgqtjpDtHUHp+oSc+8FtT
5c44smN7NCVwLaMkRuJbiptkKzh9oR0iLI3o2STZLxlyQvM8wxqy84sL+ApiW+qIsIosRwVqosLh
i6s5Z5x4RiEPW26PlFjvFpJUgbdIdBhIZfet4ULm8Cc/X5y60xEQJlUURSARSETACNeuqxQKe/zU
7MyRQzFJ7QZEeNAXr1MBzgJKUqIsmmcr1o2TmfsUh9XtPB/FLqc4lzMvgUT1h3LPWXTO1F1iFe8Z
upkkx60X+WVKiyMygDe50S/3Ie+4nE6kVN++petAuvga75PVsTJvEcADk3udel4ZYc7KKFsg0O+F
7IURBW548DhxJsDUlmzbGD6bX8jUxsV5ix0gxIc+OBunm6zShHV1mcrLCOOYNmd1014tuMW1Qy0r
sDKgCU1tnVhMY731DxfIUqkkHWN4+PAjkNy8tOw8+ww/ToWwp0rm+o7SVrySjUrUb5Rg4a+nY70O
5pL3z+ZujH1CnYQAKOd6YbQ91z1OX3/gCQN355A8QaSmtbAyeEMLy4oL/4eZZpvScCYyfWFlBE1h
NWRzuS+ah5cbGXCKGjiLoS7uO1xwWzJzr5PPY/qVSWmx12CYGNL1YFpdxpq6AwDxUGB39R/mlnOS
YyECokZ7PhSY+TMMkuweQt5KbbH+jVPOy4yXEi66NdqzvI9wJMLtPmU8jSq6Qb5lEiGnhbPxV3+x
gbtRvywM9q+Au0MVODLjh15yVtTCtZWdmsch0BQJVBgVfnD943Mx3k6g6NZJStlRk+cvUSf7pI1L
4e5D9GOENy4VXp+1+cLSE8DOh/upQlfTIvcHF0VykdcfDETh9KCkGcBlwnCjcMw2SerX5GLzXsJD
VSSFCYA8XTOVPtAESzZor61MuxEAKAM6b2BKUHmilmXMjggH3lZQ6oA+Q6Mlabhh2ZK58x+in3Pe
UGhQEd7ahGIckSYE/mWGzXLu5vKzdN5D+v6n8e2Se5veS+Nr8S0UYDrvv1CdnhgNlptXzfepwUAL
nZHupX0JAU5+QAaVwKOjjTX/GdB7eenCBg5ui3Upv1X2nozwBOe1ZUBEbIJtlzjvFpbzfzhqYsJW
j7P5VwGEOWPeigkV7FSPxQMhos7XZ/VDN8UJiIMryx76+tO1w+yWFA3sRm2FXaIRO521AYzUryna
IyBb7EkQyRjwqi4ciAd3funDuOKDj0WpYbs6ssYNVNxMKQluVujmWsxGJLHotV/36hxG2snKGVWm
AzkN/JFs9Ean5oKzo8kpB1W+opzKejXY00kFfurVgVKom8bRAGgtRwzu8VfATZTXoeZijIX7RalZ
Ze9md/P/Sn7WhLzjLidY+teRxngNmta2IFCPr66/pVnh1RAkck/d/8ppRfQKlHhAZX7nIKUqUOoy
oBHYyfkb6ORUtMlJJU6sBYGMu6StvvUPZHPZ713C91dQrwkIz1G4LTdF6nAVQcN8rVX85KyYkieo
D8J7YJG5QJn65Kw9UCpU7oFdrSJ9p0Vkc2yGu5WXAwj3R25mn1VzYMQICO9Ip6rzz9TJzLfl5dFi
Rl48VGMXmbWOIHkBvl4bjp4ZMpV0UKXUGKx3HL1AQn+rZ3gxPyTq2rRYZUWGflZan9/ND3eBo+6a
kGRiIg/4uKgK9mAx/Dikh185jLSje/+fBUw5xNnZYpFV2lALZ1o7zh8QbX+MMhbYOXMd3xSXh5kC
1LGyd7wSZmyvXW1/VL/BdqQcE3P5J3bicsTb6PUavdhM4UwuLw6Q5UfX8ly2W3HKTFI35605HQPR
1DTGCpu3HAK5vnncP5NiCRCRZn7sUYRL014+wjMCi4BQMlvud8tGL9E7o/kaUyWFG3Mgxo8pq1xP
2YrR9nIj/o4tk9MjstB3UqyeSST3eT9ZQvi1B+9Ge3D0LOmxMHzfTKG0pRCvJIB9QUParty8xza2
dyK1u3EGZhf7dPqXMYlk056l7gNCg87aZYhtjwi9IINyFcJvEJ7cuUFOUgPvWkUXphDmzggeZN1o
4cJh9sI86tAgZ4sFV4//tXRjofHrcvH6p0fHQOW/VYt8XTgC/UuxbBMpjKWk5lNvw8ZhCEKnKoTL
0Ri8kYRYXE1gWw1W21sggKxUIWXpGGMtofIKtGeaSe/FIsYEjQfGmo9Ums9OczsrMtfB6W6psWaQ
jwhIW94uEmk3iiRTx78zF7R1wVSnyLhLezCUK4loyydMo9pu4IJJaMIRrtoq+P0A6SpFsSG1HD+T
hH4RtMUqzsqGlLbtDcr5LkcwArlX76UPp3YzKF2XppRlkF8LjA74ZzJR939eLsOnzOjhCqhySheP
R1KWnjh/r2+kRwjre/kIcfA920vgdA+V/ggrk3DcPtzQnt62DdWT5JjdYF52vVIKPH1ciNV7iCzR
Hgx+dmJdX+THeMuSd+SJQ6v+EZyYlrJs3js9sk/nL15BfCy8+0s1eMyFU8/LGHremLG9lk2x5VRY
eJSLSKXpUl8q2rP4XsgtmW6VllZc/Bm+/ui30x5WIosMdQyIr/QlNwggwxzyNCgWQZRCz2Sq/S94
x/Jjclr6m2ANPotYcendpYxPIvn6/CEmax+POqnWUWiCixg3/m1+6v+6Mb7BDhBXejRU4o4s5egc
Senn9RcTLItdLSLLheX+P6CudmleACwpvaXxVvXnOm9PeAje9emKS7GDCqmGWMZXLACjjLqWBt0x
diH4RH+WqCMZHPzzNCcoPa8b6l34ZVV9qusLX7HyOmCPGIT1B412V4//cTr2EkX78GUXyVLEVpxQ
TpGoolEpzahpe6AFd9S2dR5rsB7dT//lcc3rQEwGF45bPcZrjv4DIAPRQdWOjVv3dvObj4+aGTF5
brrlZxrbsy6vytGmuwUAOeYvHL9khbPaGRubfqQpRWT/cg3QOlhQMgvQ6wew4kNQ2gaFS6SvZit1
wSdjr+D2RRK6x7rMQI00ChFrKnja8zgjZfIol7eUqFuXplZt+dbm+P2ckEOcHpoW0CPHhrLQ4Kf3
a6+wOfcE7rMyp4wunGSsvo02wajMD+zqugu8NjEfKQXCWkSZCECt3NJbBw7iRlCPlrG/zXDrLvCp
PEEkJslyg00RYzub5ooNR7wOJeL2bFpL94gtAtkrcOD5LnO7Jc1JROr/ttKbDo1FTVMzGXO+rPLm
sAWZ2ChRW6qnGApoKylj/3cackgwZGXvkjyUGuR/mvnCHfInegFMMDWVozXrGHf+lho/JC+jeXxJ
xpFP0tD7iayhYrE8J0fvrMv4faMkkQutDUxflWH880FCxy17OIQWjjgCpMEAFfvbmxLjQ0mit0ew
Tm+9O5Qh6q69Zw4xPYURpZIGAgITl+iTTK+QjsosJeX1Qxmj3nThSkID72UdGebfIUawbuXiI+4b
RRNhI095t4Qywl2HRspRFXn9+QgYrrH+REOlL/5R2urZTBzzaQOFn9Ch0WnkT7r+qAfcMooKbdvI
qGQLOxVuazYD431EP4c0DcC92mrf9Y9DQ9NMhM9yJQmwgsVrgg/bqj1bZKhx1BGAGpMdJW34e09s
E7L+xDxziEMMc9ho9dXenxO2o24yQt24WH9hHk4r6i5gvN6bSAx3RowlZl+2j7RTrQAiEYmY0UYG
E0UZYjmQKdYi6lYqyHn1U1MkoLPCJhdMe6iYk8Va1WEzFLdMK832YeRDBeVc3I6B26QtmmJ3kDky
IfcWkczvUGFiUM9fJfzGR36KljXYA1zSFu4K4M1RRME/GlRHf94wYJP/tZMLSJLdVqLv+H9zdNT5
OnxNmaPATaEUhqo/NLwAxNAb11SI+jhn+KoypgRX4Vdo8Y37y+QE3EXmhy36x5iPLzcxIzo6Nd25
izbQy0Y5RT42POI4xZRcVhA33WmIXNMsZaF/4LRNuceGkic1k5jNCLL0qRnaXHpbLy2cUWsO1P1k
9bKs0tjtcDFGdbsbI+MzMyuDne3wrVPQmwj3Y01DJnEhrFDb46bcDl/Rq14Ak0byeD2IvEQTFCcy
edfLFN0eOtGOawWMuhB6kmDCmj97dkEa+KYufhKdnkK36J51H3jrwVZU69ru9d81rDCY3ApErZhw
z9GE2Wt5x153/9i9+nkkjjxdvmKxeUkcXGFfVNR41C02QnyXdYipOELubyxAaD0bEKtUiQQbHsOy
YeJlIlC/NzC8pYM7ZVAKrog5zfJYUr3uCMgsuH2SkTBDm/2CUBoOLi8lgBHmyrjs7+p6RGPJcyhk
e8ggCDnb2Ps4vJkG/E5eHbJdevaUhcklpqazfxJPbE9FuuJQK8I93CppBlt/2RrbU5xjKAD4codW
EIZ2DvUbBNjCa2FF0qCYdhw06FzMIBQLvojnShUNXjPX79o15KfVuiYQOsQjrg+KgjWrlonz6cTk
jnLcdy/I3ABquVhmLKpsp5u4ygU18IPl9J/gRzqIZd6M3f4FaE96OZFJ2yy+TSYUcBWvsuX2x8/s
2rJjxCl+LudbiuI3K2i43zwEb0qXFOHvxfMQXk2NDBUYuNGgkGGxHm0bwM4PUbTJtPppwW4OUTUI
rh010ymfJDiMk2QzVwHurgVOkcROIs4UQR/4UYn65F/w9uz4+hl+ljbUphHxY/rSdWB3A69jVvaI
aRoTuFlaFbB7dJq+qBErb96DIewWpm/QC47EO70bAt9RLs+61zALi+hr4yHEcZ4LO4t7lk87TP/9
ZagmP6tFEff50g7SZ4t5lBWYgBLWv0VyWhnopHQEBVxSSHBBQDpYXqfoC1T2seYMupt1BYy+Io2K
04KbDrTLNn+Ue3sVm9OIuCgs+1G2ZawVKvlpwln+xlo5iRbj8l+lp278UINA8rw+6D+5C7yZ8TDc
itI0b5PatUb8Of0+6cMtqnX73P5LFXKI4bB8mIEdEklTUZhoA+2I5BxU9px06nvYdJa1eFtCZKe/
HC4QFCzCyyVBh4EZfF51XEz8W4a35DV2+2w9Dy5Fo3wMl7UxTDXxIYuWltX7I3ooVh/t4H0kw/9C
fFhSgyhIPn2CcGvg0s0SfJHnfUnbjkq0Mbp5WRbRE2lhebXQV9WX+VzTqZqolAq9nhk0l5sbGcog
ldvTZEE5J7tTGRCo4SYlyP1kDRPltE/Bk2Za3lDSSk+21I64T5tZHpFcwUt+/DUGG9wm0QjdTZUf
r9n83GEezLTmvPOB2A5nj7RVu7JG3sLFtJijdJIjzXYjo65uGMuwe3bxAAkTjPReFgeOQ6sBYduH
WWQpO65VBiUHcZiFWjF2gBdm4uoOxORa7UQPUQvKXy7MM1FGGy7EBBHpHi60zYPeIMPiPGpoBXio
2kNra++7H25dgBuC0DZLM8R0J6zKdPCSaYKJdiOwugxesLBY165ORwlEGYWredWSM/iBk+J7tn7T
f9tGqOuV68VyxjhPqTLs5Nl05fZ8VzITDlaWJhu2YqQf5BNnIIWR6Z8wdRPMMxjVjSdVIKtXDzHI
xXXZGnnzk2lexIcbLrMg+/0Dijj6pjZVo8yJmSqPu4HiYClIteK4GRvgq/AjjLyuLbI3bkWcVecs
KWmhRS0ySXPlUvqUk9d3aRY0v/wrm30mr8JVOs5RGTxqAEaJt2E4XijIj2DAsRYYMJree9U9qOpq
tIsaDN5s7qRdvSVvpgKkaxbPScA2ox+hHXyUZjAZ77qcTImlcgyWdy7Wb74zVj6t+QaL47VSMbMy
whOfoOgZoUlUja4KP2/b9ruOh6ykpPiSa/KNDZIYVzHARzhsuGL1trPTYv3RD34WlzTlm3Ii/9mx
B6aS4xEyGjR1+7xLGWvWZIV/34h6INpAS+Vq99vzeN2meGRjHY9QQY4tM6rPR4CrBeon+kxP9tRb
2By70/UPmjd2VamJ9dr9Tid1QHUwsQtloYOzhnmU96MoHjJWViz6AG8C05hLhdP4ypS2vI8dg2mR
YkTmm61tLFIkYDQ/2FGu1KR976ECR67LdhxysmiAfzkgyT7mnPxtIkM7b7nNvM5xN5boZP/EFhx6
uaDvvMQulEIxOacBi5+rIJWKwPoI7bWqnMnNCfu/QjpnGvSAKSjB6OpLzP866VWA2FX+KPDmJbei
Bhfd3TNNCwuQSx4mZt+/rF9RDfuIXkfh6S/adUHf4Nb0jpW1XUDpEqjhh3pUwpvaASV3Tm/Dyhbe
zNwtTp7lV8rNq0CkOGAgtVChqAAPnKXEjiQLB8ysgsfdjKoJuT5LGYvPJqrlIq3Wx2RcEcWoa6kZ
XFCTulywQ3lflRhqkg18zjXQWCugn1neN77EmFozY0v+BfhrXey5S2W+4AStbsTrdCQICt39WEYM
ijV6lT2ctpz0RV100nV9VJRBwRYbYTzpYU+v/H70zD3ORVsH0fr0wrGOKMLfa4h7lOi+J+iJdhEj
uva2owtNasWJa6pd2QKL+79fvGi/GVjmwWmIOTVP8piPGyjcUy5YBpIoCJ1X8eTiUx1A0iNDyRYd
2X7lhz2zIEJ1aXVN82xC/BpEryRkdlvdM56ih14bpmrBMvLoVCkNJ/nrNSsPcb0u+fEhr1RL/XPK
mFa0PTMTX7R/R+JaZk7pScBUElrAYVXZ5k5Fd41PNB575rFUwDIT4oDbb9zg7uTI56E5+ohBzR07
NUorFN6aYERLna7+tQy4sSlkA+pSaTilmZEgAoGouD7mqrjPEvDARdYAUDHZoydqLVfmBfrlRjs9
mRMDwESAFi/m7T7aPoPQYebpFKJbZ0ua0eSa2520TGjtlaB02zP2MxxhU8wppDPoabE9GZ9dwTw5
w3ceVDFdnH6UAjWEvQUzugQLmffzPx8ILu8kzuhGdm6c/F3FuaaTj4gY/0ESlklhMz+zM7hVBhZ9
QlCvVFieodlBxjLBIUn6UWX9ft9Go6P6zF2Jb+0pj5y6BI4cnpb4fqdWy93cVaqKlfcfU2ywl847
oMNbxx7EVt+Pd10IWmLzsan3HM8CMOEKBRFS1TBb26vZ4pEw64+r5nSyg+ODNmHiXYu0SvBC7qQf
A33xK5f1P+hBKwOz/hTNDheCwumT7/AXW4aRP7HKRH7K8XrzSpoRl2x+rif2hJpTYLZgTR9n/XvK
W35OGFZ2WvLn+GwAIEB9oZ6XEoZTyTW44sEKnbTr66uCxA0yJSFSJco/XMOn76FsdmEQ2nJvAP4S
DEXOXxCA3Dmy4JetsUW2pNXLo+15OE/pM3JHcx0QbQC+w4arkdI/va71/Zj/2e6DSzwumAQfoCao
p5clrEg8nV9TroTxe0YJWt6FGJn5SCoDd/sVncUZpfFY9oCERlXB9OOLvBUlarKGCyX4t9d2dA6U
kKUHKiJvXmd//Aeq3FvHKm6duU1cXaOQymItCaVTpgW/3Yp2ftIPxA98coRLfy+cIzvyWj3iPI15
77dW+hMHlycQy0dBBPWj8DrI+jxDuaq+cel8zmE39Xtht5JSYYOPy17HZfOA2uNxjcmVm/HDigmr
n/m16igdGElpaMUijvn7qpBLCFBjjU2Fy2zyQk28pCkpMXZMyrEly3mOR62JaGa5oMfRexkbOj1E
cTz0XQBQGqzhOd6QdaqsrcLl0Zue+OBntXKRGAB5dDpEkNpA0qOM28oSIdGRI9Q/f+0hmeCh73Wh
XfMloH7NBrX+zIZ7uh1hjB4teChJQ14uegKomuNz/ub/KVm6+7OkcuUzAWErXBdTgMBnIR80Agle
MltLHUTmnciLkPRiIiQ4jTgT6qFokQxDmcpI9j/nXj8P2mYKq9uhM49QeEMyYrNGYQwoEIcfp1Au
1bWS6I3FhxOSAKQ3hDJuD5G45ouQENr6CBqdT4rPdZiBvLlQXl/x3kAfY9CRTkNV7bQvQGCf+i23
v4mL8w8RNPCnY6qFJhXQWdrmYvweWKOfABlQnsFEvnPrdXWESfzY0z5uuK3RQRSUguUXAuPaaS4C
d9TMJvw185iNeKGu9VOtjbhRAohtj9r5hRA6Viw3c/tPQs9eZNUdhk4Lz6dososHq05RUa0pIHUp
e7pzoI7GmFpboT0lXuKsvPdmg02JYmsV/eq2dIrGMD8Qv3PK77R9wduxB3I0WOjnIi1UEBBEQVYL
uazx8oeE9Sz56YmZWaBqEXnoLQRAwEJzlq7FEs3otmvaNkz7AxYP1ANV09D7f3Wq5Vx/JFXjkSSc
xCUna45pc10u0WBtYztCK8LVIMHwSb1QjvFMfylKhRwMt9t/xLYhwwkHDShcVnYAmbS1K1S5Ff7h
U+VlYklL0Nz+OdstT8QKgbg9o8xj8RnCp6QbvEjn1xZgnYi+wT3qki2tmdLAHjJBi2Dcis4KKXOn
O1KTNyCn3TNRquTUbm1qbm4yl00/AkPQRIiLlHRpFmBcNbu56Jc4hprjhkuPEBuqToNejgI3+Rsx
X28G/IZ4QK14OuYI/DZKYEae2+V3F9+4bl/WbffNnDOQhyhU1GKVrR4I+tm1/ScN8ZelFo/wHIdF
Z4RK7K2F9t4APeIhxzoewnuej/j/kLQPpkPs+riid50nRyFXU2hqYzBr8N5cv9C7gFUGzGrCsUUx
JOIRy8b0p4IKmoxdizUUAq+hDW6maAJschxPacYovIJ9MTASFAieTtZSekDmvrTWIcxiOd/WSVl6
GXjeUIL2UpOiE9LOrs9hA2sTI0ciS9B+xBx2nxLJBuN2b4EleKSTEVsiB6rgvkugm5AALsGBoaIL
z6z15n544sCdJltE1t+bQWU7uVIkq9S9sJT64ql5PMjzEDd1JvBIdR4EwYCjkxSgVw6TwlVx0lqi
7gUMY1N43mV/wOyoohBufyAMN91Vp7yGmQUI4vhSBqttEn54FLSM1F6NRvbeUTQPCS6MBUTlwcJo
WqCHsn51Vkk5u6tHMKxWjmuX5XKGW7DtkUVvg2R6vTdun3wnA9oy1h2yswURgVwr4n/tjsjctKtJ
mfD4mr1j7ys7e4ffylOLHhVehbhAxI6i25Hi3Gvs1r03ZqN0wLyD8/ZCmj1JYVURr7SCooxaZzJq
/czTupQ9XF/3bZbu3m82qGt791g6f28Zkzx1dINwJJ5IOPtnnJu8KikiFuQ1efZ7OxDg8+DBTMTx
kGz5Uj0xOkroxldGmyXCwmTDvm+/+Q6m235OScV9yNIFg8GtyxllxQLzVuP1JuVGmY9rfHIge+ax
iy8SXQWyyZeI0OqluVF7dkHQTwYuqye4NV36Lz/I0R5V6VaXUk5vrFvfknVUraAtjX8MbqVaE4tR
qRpm7n+/7zWRSB6AvP9OsX/41Xs4MS3gKBKZj5v0OKfi9KdgEsUDChP6m5w1QqVfEPz4pk03cdCt
HC2auG9SyPQLRB0Jtgd2vlclzIxoaFaQiYeIwpFo4YmsvgAzaEpOQwbx8n5yLKTMtDpEgIZJy94m
ltwyUrpyaPblfY+0AF+aGsJWq6LVgdH9t/8k9G1U0fw9edkf5FhJGexTfiLFla8uLV5U5o4gH57Z
4UBhCoy8Af/oXbPPqi20ee+fnuT/NWYRJC2svFDWPsO0RR7wpfu4HUmx0qLidDjGqP7fsLCmZ5Jj
La69lHzcZJGRN3RPq+nxEuNga3RHzdPCG1pzZ0s4kY+WxTlTxBLqeQ4nMqxU24AEZ76fMUGRCOLC
4ZId6r8nEY5jJUajhBVudi71ehDpqxN7f1BTKz4qiSBT9BoPIbUYkFeasFO3BxiVZIZfTYTspAYy
PobvjzBU9fABU8aJEtoR1l5P1rfLGXZfid8qnPm2HQTGonbIxso3UnVniJ8pxJdCMPlsHaWaoEnG
18KjL2QSLW+AZ0I55GpVs992eIlHZG147DGJpwcaur2YRaequ9VPMhfjmYisemx0LlUoLo9fY7jU
KJIhAQ3WahopUiIRYTCR3WiTCAmI4kSzIAD1ZHjq2h50adIgbLlfo/aeldmKQpTwFsfrRCF1W0Ui
o2c0A5EcdbbHNrnKHyEfL3NoSKLvh6f7hOqsoWddHuoJ9F/F+nSc47f1m3yrxIp3p0GD7r66RS4I
I1AZ6fbyad2BeqRl+nPCsw4rVU5ioncn0f6vK0nb9VHsxovtkfY5mZ8xXg1wvMA7SZyuXCFVZOFM
AJXfluiyYlsirlqJyGL0rHVGSyjBz46QfCx3lMDo1j57jOrC0hEW76tfOFkCOiLY5vib2XuL8RsB
BGlXCjvw3pcNbS/Sh6LAqIsOFNj4JTrcHQjFow63jZtkdyJKH6AIwHkHYHHKwPBuFwVQBqtT3Kdv
t+FD3zc3pqDdQm54QlxDtSp5woh+mTwYymcZ4g4qDV3srVBDppQgwwJ4R36zQ1l406AxkIi/0yxQ
91aT4jByPwAHHd4PUBy+4YOJnlvX0ftu/ifqSbvUubQm+m9m5OQ4w+onvm8y+TtIGVbZClUVyIxF
ZHMkQ0QgptNnmNvInXObtvN58xY3T6NnP6PGNVunY8ddwSwFl+eD8ZDYrIEAq5qWOVqt4/7zOvfz
B+FxVRmYFZEGbTlc7w/wC+eENBzYKjuac1ZQ3kvvGRzLzg0O2OkkTsrjeMGHuSUVULByqgTXJfhD
yycyc/UHbCBUaECSNu0q3KnAetFMLx7TCUr4EFQita12XskBWSPA2QwDUQ9lT40iFdKtlK64KCEJ
SOhBSLAOrQAykbk+YMP07XW84VOMczBLvD0qM7XLgRnqlOYaMVXINftjDY6/d6F9qaScjm3ARlI6
wHkOe/kSZBw0Ep7y4ugrg6rZ96wuVsnuhHG4mVjVtZW0NTpTf5G/YTnia2NMMrPadskTismNamwe
nuyRbsqFYO/RaWutCbAA9NNjhv5D1chiWN18hGHroTJZvDE9RXTbVsDJMokjnGuiN1BQSKZ9rJyq
9i/ouGdpiokjGbKT24N1leTEZf6Bfx1TSkgfUqb/q9By90emTG2xpDevLAJI9f1rGYeVNu2H6BE2
HHmS0/xNvcmXzUGnc4tUnwcwTUw3lHsUYoj4EozsyVhN/XHSJLUV6hHYE/+1yWwMoGUcUw2NIzut
C8dVWf6We4tndplZUz1CptGAwWXqNw9H9FgFjJz+0ndKnPT2b7KyRIgSsZzj0y587ek1fHKkqfAc
Im75LOUN5u++6brWJ+UBQ0DYX4XBebuJbiu+o8gJzp9mfTkNFokTgU8gCPBp9J1kFHR+QrI3Ybkx
zOGBgFkR7ar1VnbqG+7i4QTXgD68naqjYCalRsCK2d8Ms9VF6YqSZi70zflzftooT+Sa7gqKli0R
spuyoEJ+jA5/qq2E4pBOUQWFIQZmgJdimtejpCaU4fbUeH2D/Vk33xMhsGSrneFSVD0F7c4mtx2L
6O5+Lb/jf6XLtb9gMaR1FuDGLy0Gfu2v2RxGGhSlZXY+el2qr2tGBBO6kxqyOxdheb39ZG2z1AQr
ZCF0HtL44GnxTnJoVjtljMZEisB0OiaJga2kxSGWy7DlIXmGz/wYu60BEu0EMwcEN9DGFBoc7SXV
rXxdsYw40YFMC6VCLUHpB8ilHeHDIcW10tPxtVZvpmjET/AXsXvEgxfP69zzSGjdGegcKGG43KjS
Dgui2iKfauth2y+mvh2SWju40vOKiJBFCtsjv3WmRt60kcicKryOOQkLpf1OuMWiYUVZUun+9OUD
e5pfjvq+NoIDDlMmljU01caO2V48fiTwNHtF+f0dlcQKZ5Djr0halwyPOUXeWYrmB7CBV2wZq19s
eqend6PWniRaa//hPgqouvl9EK2bApBnwbBY0aCd9yLAvrpQ5Tp6v3jY/chcpohnp2EAmVQKI3rh
odV10UW/KnWmrglS/jqE0uV4TIByYxKZ2ohFDu5Bx3dKAFyTlHSQZ7sZvdhzUKeITugWNTwEMCDg
MjPTDzKyJcn6xYoMyNy5QMO/M/LgYBS/Dkb3EyHUq9u3G/aR+vZkiEv9tYysS8EUSk8OB9WrAW8R
m0qwGvN6+o3RWCpLM7iSsb1s/pScFIueMHzEtRjaxXCZ6zOJ6vP6+T6fZh9+5baEUfWs/bul3pu1
1BftZg9/d6Gm6HjQhavf+lvwAzRybovxDTfEjRNYc1/dGUKDIAfAWmACAT6k1n7DwoZ+4hFr74gT
Z21XCQGlNqKArDHAxVlt+zm5pIPCtkLphifKeVbcDmG+4XVY/3f6xbjNd3HFu5rNLzltFm3H4j2T
MsyDwXpRr2xJjPPioDbzi3tHbMXvDxhTxSLI1dAbUwhO5dqpcP757+XECUTO1drYEkwwGzJ1r2I2
tDkaexyRCT0FEKPdIl9UoLcVQ47NDmeWEKP+S6sIPEBxOT2HyhqjYQrTVC0Hpg+zYduKVf+Nx429
S75o8w5xkccGqdh+e+HpXirVN5M5OyPdoppsrr8br+O8R6gtKMHREtGCISVR8ZvciFk3pLq9rlBF
43/IC47sL4bTGR9+0lvx1x2DfH25ai0I5lm760Shejp7g9YOjrW9iyt0Kw+igMGcbT/Ojm/oIwzB
qQvIqcJ6RObx95EkQL0eYh82VJb5SQMA1/9mlOmg120gKKkCqUAAUIfa2fAdyjC2Li5HEHo2qEvd
hBdA/Sj6rh4h/4PbhgoAFkFR4ROCIeWZ2qF7UQr3i6kzSKNpkl3ZCzCwHYtgSHvFE2elUQ3p0onP
ER+Ev2Lt4HJuThIPP8uQJPll7UHrezF4hTeUAK3JrfFclZItBkCqI5xJzeTNDTCHloP7rty486p8
qaHjfOmm+wEr7Bi18BhTmMc6I96bSZsEnAilOviqzar3AnjtyCo266N5QLw70PIW6j3RTAWBt9zb
vamcSfL7CYR1KbY4DK0BEUmxq+lFh2dhbhA4cWEonuF6S0IKsZE4i7JonBLlg2/vEhhUSsJb+mTp
O0syn2m4W68yx+E6N3fBiY6d2s0bXYjy1M4gfAfo2JZNnvL63AyiZXEDE/sTBTSBekfhqz3LJmLE
a2vHlp2DA5nouMArJSEs1Wz2HNqjrEl4PmaruYKqKuQEfpHG6tro/w7Veo7W4O17HZX3S6c3Redt
f+EFhA6S2LnZiONtuA/4yNvolyXbQlFKLDIx21PT+QVgIYBLUL5P9QcgZiNC+wLp0Kg/86myUZOk
lcC6m/stCRqkS+yJAmOS7ztMnnyMG6DXvADCXE7lOeEqU4pq/8tJBk+3s7DucYwrGxLQUpcrVOTk
S0b2TJTX1ZJt/z9LbQ5EvumwSmTLDV3nozHi/0Fi258kukXruBv9ZNYr1AaEoq8M5kumpKVEdRZZ
5eniMfLAdgOZ6/qJ501parn5ArfB1/7f50IYBbi5AfIFvFmo2SHViptKfxd2uEdGMzSZDjMHK8ws
ehDoSZAcAeaXw0EMqM40iBUQ+QBVnm3FWbKTTdtSMxaBAN+aIqJd0TbtxnAnTRb0/nRk0iI1CEc/
b4J2TmKKd8eVF1Wai6tFF9pi3OhePHP6isdbMSTbK8zUt2+ORhQxWRfM2CU7uR4xrkzRZkU/YEGY
S0zu/XXpvsZZY+2Qiapa8y2hd9uFnAxaLU3gYrDICA0CLMqXgEXZUmUGLh7f9ojWiO97Vjr6hwEZ
JCtlbIZjd0VdyoZEGk7GzFpMK2zXCQmjIC4kTzwIFu1slKbF1M6cnwmp8F7vvbChJY4UUKDNEK5h
kpjh1WEBpg5Uh5mMmolrtshHJeq+/Rno5+arBhX6DLXvvJkDWMP34n9OE7cyxR7/S35wqNQDTyGm
tN+3q92ltwmTXuDwCh4nNWY4GM1P/KfNikKiosZhJUzSHnhZBcwQFj6Xw2urd2DpUP6xeNO5m8O1
sgTs0V7s4XuLufNZDl1cfWubDhExXi1wKfF+1erjoW2GXiP+J4WRBm4YwGYY27tZo0YjaGxNxm/P
cVWiC+AncZNc+kGWhHMW+Xwq/X3rS1SP3/AGdolSntYk3aR5Ht4li2p6QNFZks0WkAF8zPMb/HQ0
DO2jLfa8Xx81AIaPuR686Ww5c6BUsQG6YSQ9KW0E1z0RNeGm9mOPkH7BbMiyC/1e8D38p1nMhkHE
vValAnfzdjLnlye5FqX3k9JQX1CYNS+Bo9sAHrVdWqixj5RQ56MSM9vOz4Rx1jjqavsoWopv2ZBl
xIYOCwv3Zqw3R7UBFqHXF04AolgtB7fKHFRftIfGZXYP8mOLeRLI/639wXPMhC9aZlMPrqVfCdvZ
Dyl1Fw0b5Vkx+1SlOEGBGr+Cn3x/B/PUHxoF/qCoHvEEb/XxMHFdVsdtpskxnXPrw7uKXe9HoCfp
64VLdJUFMjLj41IH/M2ceEi0jQcadhzbCEst5Y9hlx6i1UywLhx6W0PiElrJ1KsYyzhZmqLwMPAe
HpLqbxSHbL7OEMTe5fGd9WmYs3j88f9Abvi0eseZIv90vWXm6aPAAOYiZu8WgdC/A8PpIf5rZ8Dd
TRQ0LOFfakkKLBd/F7qmUzOkN83oAE1JMlIlPJLkv5wqNap1OifbR7KBT5EgHpEZTdZyXKjbS2j+
5CzjoxmtiNn3eGBRKqRq4V/6KOXplFZCLTcvvJ9DKHVxCaZ9iOmZ8Ma3KGz2/+YngMjawJddJeyb
0qteHiTK7rNynVeVhBxu0oWjOf3i1Wx5xYoWzX/JOX2sykTTY97wwtxrWG9c2YiRvoelZOJfj4qN
yTv7lnKNVUbmW129KlrPnDvHCIB9JrEawbrXV9WxtvSEe+p7sZw2LI2G9U4Z06LV/TmGYR++pyN7
KLbp6QpSTgS2dy32qWcEKdFXwRNm1Ebmb5R3MqOX2/D9AjyqFiF/25hU7c9a8KbqOJrlSMcLnQTc
CoxDz4i8cdw4fmaiEXeomUcxucW/hJCrl6UtWGLXpWbe7eX5zU+n7VinxDbOIZWeKn08fSwo4TqO
0/U7A3RB+FkvKCLR+KCptWMu+iZMgG0wIQ/kB0SKihxVpQ1i7165ev5ZRpCjR/xdR5JNfcvUb9gx
WCbUwC9DR4eTPiW067xChSo60YRed2rR8rGGkm2sB8sLwcTS7bkjYXz/y1moTXcSXhAaX0jheAUP
0lrnrVibt1JyP6BzpROQFfcvSfhOu8EcRZ0gQFS5nFtLu11UpIqU/eNFJdr5v99j6H+MR/7GoIPm
nJkHUJ/VW/lDgj/kQzVOcRgy6ka/caRj+iOv6RRORRQkIBfijRI7Kj0Z6D8ze7jUnI4KmHZm6no0
0TAAKaVePkWdVVJe7UFtJQsSSIgYW3t/mMTCURNJuzRvnkj+FQWOvH419Mlt3A13h7wwdY66Iji8
//wte6jW4lvkKbTuaZX2KtmTnfJUbAiAlMhqeMe0Oa6NPQL64mKi/Drf3sfhO8/Joqq2D0iI/pJ1
r7BVEpl5JrcgpogDWA16yJ05XzMVbnQicRJ2Z1dJVchXgBHiqX5Gxv+nJRiZENg5qBzrBJfibms2
EA5zY8zZcn0+VMx1C1AOHGCaH2Pi7dHsGijp5oMieM2oaGEPVyZ8WH99ZbWjIlLJHIjHXl/y3IqB
IGvaFRKmEk0rZQoDNp7aCpheO9GfR1uu3C0ljLV1bjumdBYDe+UAz3jWTvZOHNNYC9vqbaSdIV4+
iO6tDt9VDEZ1aEJrzb0fm9bqHSAOTpIsHVAECpryxhm0bmCJ5Rcwvho/15TBbvoJaKEEybWkC1hQ
VMmis1IgMk8edloWCFxX0Lt/B9sC67iHkwOMLPgCkRCxtg5gVZOyIEwrfO7HqpzZw36yvrlM59wq
k5yoKcRd8on9H+YYbKnlO0DjuDZezqUXIGkag76pGs2ytv2/Z/7r84ft9+Y5R2oYoCcKGZlqK5zk
M38E2lmw4uo4ZXYV9NPBtxtPpr3ovJlohyj4rWHTkA5tUmoTUncm4xHMnJduu/jvYtJIbGsKNWoI
6i4v5jC9oL51IQJP91nDDpxiMHqJkegAlD1Gf0wFGDdT9qaDuBDwUS+V1PvfC+WLimK2GjJ32YJY
zNA4hxg1DXY9l+W+sFa+TnOssZT86INGJP9kA37lXrEOcnNM0uc7QSBV/CHG0gz3e3SebwQTeX7s
jDL0ho0r9rLyyv20rdmuGqzn9vA9dHEGdEk+23QLNwauaBS8fb2l/3jq/RO3RZwXqefxNPI9cYTV
D4CSbIM27HrIR04bInlkqJZtjdF3HOKzw+Jcie0wzOp5JILOTVolA5y3QKLZYjY7DRwkgwWq4J9h
rJ+e8KGUlZBcRGGPAdf9eNW+REDhh2BiLvMd8k+UY5z8pQc/n6KTbgSRpb7qqWQ96BMOIKZuAN++
QRepyN6zd17TJ+DYbwTsw2ePJv7AYMMAUQzFNRmHTla1NfMFfsVHALArxz4lgqfqipvgCtP25t2n
1EAFuD7S9ptaY+nINk1aRW32aNczAabUd9DkEKdhmsLKO/xM50982vmZbDik+5lfGCwSoqcZutrT
i4z+SDwnn8gq2la1VUe/ZOyAkFceDscyV9/m/zhdTmLy5q48kET6dz8yeCrVbmuIkL7CFZB3zblh
i3jZd47w+r4VJvOBSw64E5onXcS/TYanzwOFomGovE+DJ1owiYLMea270b69ejc5mxdIMMzz3MYA
G2VH+PGc2xpU0wj/ZCyvYmYdcXJ/aovPAaqrG5N0OpdNKpgqh7Ieu1SQlBoXuGyrMFUPINveIGOw
SbemjALdsF4jATXzPRmsBK4gq98b9Rv7Y9Xaic227T4wOq6DrHEqiX2jOa1fV2ehpo82q9gI+KY2
/DY4qTUmM5UyGxMfTlwqftxKOfedFGl7Q6QcUEMY+cojKW+mwaWSGnOZXzQSiwqfEgGcN/LUtVcK
63PZnRzUPOLdaVIUxWmSQRgl8Kr2JoH3y5fqFi0NT2BnTe1GGXB5Fm3godVT80v+gp+QELTTehV3
ALA8tRH0yWxS/M+0sUsKGFYDJ0FDfmHg4KT3hyrnt2oef+BxZOjv3F3preBKYn20pxqUSNCxOzz9
LKvoOH+9c/PvO5ddlfOIUUOcui03D/tYlQ3C6y84+KEPvjnyQeQoaoQEMdPN0SBbT7eGjcogSwTy
Ar0KHODwp+Jr6jy14IiisQHCfFUDOpODmBPX0AAPWu1ameg0tLjL5mbH12Y2n1thQTRxpgNAbGOa
H+tQWqFGuJghsZ/XvFOCkXY6n4da3JsyjKUx4KNZaO+GnVkZgeCmejxPZs8yfk1HgbzJjj37a5ld
ekZsV7eHT3o8h2bZRc8Ov9yoaV//NSFcQyJjc0fFsGLPrhGlWIDEzYv91pdn5UcV8VjqEdld7YYw
0sBNa3jetjBUD0rz38NUqJOu6yuIafjhbw60eRl5Cb3bresseVwTRyFIZimN9uPOkVInEjvskGEY
NKWNqIje5rUwZ7UdJTG4clJeOF6/2yu72qSf/fQvn0BsF/QlF3bPoOCSEzL6M3RCM8cKaohngZFl
RFcNroYR50YYmjkUZtwdKiQ5M0rFdm8RQNmpW9vBWBW92+CfQpWD4T5FOL8CUyEutB2dEi/GBGpS
RFg1rbuoE7OawVzb2ExB9Ccbw/o/qn1ueZaGQD/Eo7cc65LjLPpl9TLgUX3kz8uwD4F4oR2ziSfl
WfxQMUKJREPzXpYjgQDdaRAArjd/5EBX7uRV02pml3tQ9Suj5z7MGiUsOgr3XRHa4Tbot99qCWMh
h5ZECNf7P5SxxGc/28LJbVA2hnzxj4jhDJavA9VoPrpJ/OS/w7WG+qzPFacq6qxTU3k3Jrho7bWx
E4q27nUtq5EQGXv0Cu6qpF0nEJUkCMWAHMMcoqq/nHqERIYqN6FtB6SXeDm0Xa+N/gakapMrMdvo
R50a1bXQy0oJTfhr0QA4mBbr6OvGyFDV7w66iqhnD3ilNsEXT5TkB3G6rLL3faWETeQvsXzh5dTg
2Lq8cyhoY6rRAftvRfWfoYHPpdI8rjuVdMURpO13neaKKXo3s/MRohOcBi1haa+hIH5GG5w/q/t1
xej1fJKDS5yxzXnFO+1IJsq6Y6chhi28pFQnwn3wDo+eZdM0wI3vhEGDGbPDYEZjCh7n3YHkel6y
S+0uZRGl844CmiSg0s+n8ulAnyIfloPOuzEsxNY32sJQUs+lxBYt86VSbsPHzrCnw0fUL3zt+Uru
b5mxYpZUSH4bJ3JgurJrNkEGrlnk/9qJBeHeLQZOikASuwSpS9WOqA8C/2aqI0ecSVRD0PZOKhd4
QzCsOxMrihS/ZHhZSOsWkNaTsyWPzzXVcC1bFGynZ03m7y9SsptEEIid4uW/V4yGdPLQsBV4pd2i
0wnLw3TBoovCrHfC/x1M7Qsmdks6ARuGa0PqvYRCU3gnb/LZOYgpzQ7TMGZHrf4pDBeZjngAHfx8
+QNGJhhdTgWGt3qfuNOqDo6+vf8MaHtTAyksjlJ2GxWnyitv9oV+B8tBUV945HIeunCupZLytkrv
35D4RaKRX/sF77ZXiv1gCVCiIaLQgoz4kCgS8drp2QapCam4F7+qiHgTKzSxe2sjkWNiphFsNFUI
8tTxIRH9gPzuzZYZT+UFbuPZjqNErUHHdzNKfxSTGZtT6VsnplnJ6mxycdp4cB+iX6wVVPisCIKd
dK7MbplRW0tcwLj/c2i7l+eeqIkF9sTUt1k0hx//v9CFCXNT9ntcXelwJzg3N4YnbXVHKUbt/4GL
r1ckZxXtXtVHVwGjc7TxF6fDe4MjBkj289iymZzISXjKYhs+Xx+a2Fst4d7tpEJoNe8Qiri1l/0i
a1Vb8VseiGvqbV3MDfSuCw8RXdkK8AErjyh+PM9JUSwuMyWKH6edQC/jab0yr8kOjK1y+0A7cYzG
ijNJKkH/NI/k29GUcwRo8jTaWfVPqXux4l/mzYWOak3CaaJ0bs2hWyVJDi07A2rtQAoWaDiP+tKR
9HwfDs2MSuriXjD4h05qqa16WSS8NFTABVP2QmPaIMFqROe+IM0m9M0jU7QvJ+xtuoJ5qerjO8KQ
9v7wG0FNLYyWvy7sIcI7rkcbw5MTLJvrA9zWhCXcgLYpxDnH8yVdb5rzgCdrKzRckBI6huDxkreu
fzIhFftCc7TV6SGm0ey7QRiaXxMqMMyMdbNI+wjQ89l19EiuyqJ0eOILsnMc65SMNuJKbMK43DLH
cxBwKP1CJ7IRu0vAkdN6LQsLJI4ek3LDVcG1AQ/cdGrkt3yjOCcXmqWfs2EYKn/k66HVjcG/yc5/
blfCcdJFwT2irE/UWqsscjheSWaEuB8lxmccXSeBPgtwVK26BUf21FrzdA5JWL2wC/qtIGC2xBiT
Qb6l05L702jd0TEN5ZHjfh9b3wCISLqDXxhRIvCYijYy5xx+t3s7r1jmYqqqY1WhzKmhs2g0R9PF
RSbMREHpkSEHSlweKAVS8jyAuci3eCjCRJfXObGJYatvglEixsEAYTdiavQq3VrMJYbIrYoNV9lr
W9rjvFJSjtWqxz1VhTbY/dbpSjEmRsB5fW3Hbel72KrpCRxARedd6tYqKWXa+5dlqqVnCcB8QZif
jgM+3SRAkCgh6Io1kc+Wo25YrsTZ9jb6tsyLc7TQdQD/SdeKlB9fRI1fEHwrM4bfST8xGDJcGZ5W
ODu9NtBdD6EQWW+bEiGijFCkRSRZ5cs6O6i6zKd98BABAD2pJAS5YkExAF24N6HYg7uEd3XipOdm
ylXrcTkMhhcEWOd3vBuvcRpqUSmUR7kIFdsMzsJ5tE5KLEcoxfSQi5c2MDidjBiz9vQcL7SiXFp5
5b2FljGq66m2147S2i/E1VMkhGW0R8FgM+X+lKDPSrnheY/xO+YN2Fq5QqiPalG8x+38YI1YJdD6
jz6vrff4OiH2ktHdct2l4YtQmEXCGyzWKmfV5nV5vE6PdtcXoNYd29KDpJdwjydIdpAsePqA+255
dWucOrZQMS1bWxYQUK/WApGZNfQWVIaJArhuWNrlEGN7vPLtO/0gyVIHUlsetlshHCLio1QhWPgf
3zsCrhHn+Hylnx0vSkICz1RdQq/yrS6IeWQZcyTuLzbSWeISGvrqShLffugfgD8MLTMU2us8wEoq
eRrfBHNxD0lZGmbr5g130/WRSUSXnnGVr/OZxJTBPUV8EdNAjp8XXRVYlSrlJnmY104Cgx9Femwb
hVfGTUM/t0y3+UozLUR2p1Zp/uNB5ptAJor3cjf8UL73YoMwGQ7FhwXZNZfufGbcupHOeOlCTmvb
yVrSzk3MXDSd239ihoJTPbz7j1C6zxOEK2MEKXdZEyBW3cLUEXmbfKCqwd7r/4Jc+TKjbmT1k4b2
wZIv/kKS2E/EkCZeMhnqtdC/+dBx/EBsdgkvf1D6zEAzC0hykSO2ybECAGYBJwMri4ROQaiGOxgX
UL/a525tPboGneEkOEbwzYDNvDlkvPUqJJtvKjgZ0NI45w66ioVmgF9b9Twp6guX2Ep7TaO/EYAo
vH47Ao1oe/pvOJX9C2cSWubqryYx+8Cp3joXgoxGIauIt2BcKejbvjOWvjKS9e8hHsBArctQPJyG
g+7AanTOhWALDdCHjQ1N4jCgzt/9mVmC4CvxPr0HszUrUXuLqaKBzq4ngG60rE2kS+BV1y9xjtj0
yadJgIUZmo5wiTfFU2nvOugnKiY8wn9Hb03QIaLcIChnxGBIEonXFKhzO2GvwC7fdAiVXoE8jiav
bogtRKvnxJdx4yfXfurMm/MCCCKNn9UKq+MZi1XIHbUHiTImx0tohWuLdQhDLtX5mfSIRB03NTrB
qEbpdh+Fdh3HyxFjdQzXQbaGu03dJcjQ0VNfFAzOBUcr9TD+6/jjgNnUraotOZDiCaZamhVdl9HA
b2tR8wyq0VqgcHEh4/NcltkGlDREflVAbZslGZWvzG/SDaSFmld2MQnucVKRNShixMsA33OsF47W
rI6vLYf/2u5i1dOKra5dRxtQwxb43tZJ68/MvGEqAaCHVhQmSalovF1zVq6rGA7XyEXY/iWAoVzQ
dM2nGgDnwKvOFYqqmxTsyWbaSPkLmMHoFul+OZeZ0aZwxwdSaJo7hoJurUqIs7pEZrkVZndVb/KX
uHqXZ3tiuNUFYTOCLQ/5SYho/K5OfzLMA8lKA+5bJqX3eI4KXYQv3J8Dxq1MeRr5okIFEz395DUA
IExHXyiS9INwbMbr5JG9GXFVo26ZRvW2r0nrBjHBXGPAkjVfJJUa/GMTmVyxEOJ9xWFlVinyrLnO
7tHghagyz8wIDVDmSjzOpM0fuQQt7lfADhfBFeanfqlrblnCd7UYWAsAmJeWDz8VAylKmIqLheXK
MVq04loWx90RqUlRYJV9nRnvimlB0Y+8VoIFCUx+N/49cR6ukjE/SSXaLtTx87atnPoiTMeVXnHi
aVXpJF44S2epQ5rducNlJKTMiyF9M4Egg//jPV2HA0jU4eYPYsFtlBziihQWUsAkJodDMErLlEE7
Ov8N/ARRzJraz92ue+SrIlQQUN+p+Mjq2c87LGO+Pjecl3c7FI8zexZu68N9CalNRoEK94Cg8gyJ
/xWcMgMDcR/UAch2ZAc21OLF5rUA7/4ky4mcZfSHuTspljbpsH+mqm/mLqu+wH/FBFgSHhb6tzVl
4/mFDP3UNkwbRAN+BL2q46pGm+QqnCmFVKyyOzXKx8Q3p79+05pUxTV+T03UHh6Pc3lxuAmE6V9E
1vRjZofg8W3sCX/3buKsE4kH1r9jXV2eVmYdIhZrNAG15CZNHSFaThEp/6mnwbn0PnSHIXTa0Nly
SxvdiLjUrFw36Kf3+ddB2cuNu7t4veLpFQS9IeYcnQPDk8wpskaOUtofJ0KVlNZVEaCNfAzHaSio
wnkhba+MB8Nqii2ba0BOmTEKZKnxbatgvLaa5uidQbfNJT5Qvqi17aEk0YJ6R1gKyPfVJ7DQ4Xzn
aN5sukbu6RcvBZhZsZNCiaE04O+uYpgJHRZZw/QpIW2IJ4MK0iKdhb0ihTqGX++15VgFQgP851aX
/bBBZzfZ/k7TvhqcRBtlUiVyOzjUKqpXzRyYyfhu2TJ1EgBUSZm3Qz3Uq0VV/f0pnOgdOyx5OPGv
4BiurN9soQgyj/FANMbGoLYqrjHjZpzxs1dpiv7DXQb8L8sQcB8M6hpJvNOqbhxFYYS/ZHDTH5IS
mztx9ZeBs9HF/QDsYoZBDxY6XGNfCV0FaYLEmJCdfIYclOGGcUvJQeOsYREpCOg2sVrJs+5DJInD
eNsMgbFVZszwjRrR9F0H8ylNomZi7aJnXFPjGEk9Jv+RYxsMXvIn2rbNRc+gkuV+bFuXjHP9ejTi
/meLyw0wf8BgWWg+/lpMYxAcizotdoLZn/lWe/x2amn1QZKGEVuJychWDxiF4Y/ePch9XzddaZh2
ri25qcHk8hVHasJN6suy8bKK+JmWKO7M9Q4xoy+l1ae3nMCkxxTde03hGNygG9FXgYeAP8W4wC9C
cafNtsTntthiniI98T+7G62/WPWHzRJ1rotjnICAMWfulSFlMZVqqX4/SUn4Pmns3Tts6hs4Unel
xk/Em8H5L3skb2xR+EMbAvLw0dp5h51xtNt19GJ4YPw0FOfkfM/ZJ+fOYCkFqePMxe4r/e3ia5jP
MGQDfTuWxQxxiDNd4qIbkMS10EFd7OGKlBUBZB13rDsEvQ8dSN9sKAf1i365B+Z0ykmyuZt0ZZ35
hCpG8YuNL9/QJPIBhLAS6cn4QTV1w55H0woen2ghG36BgkLoG8rl+qOwtSn11cbzGASQr6sSAHRg
NzW+SgiD1AbUZzFswgVxXrHgtb+Ej9Rd9v1IQWUi2XeYssZCATGsTCQOwtHVXAcXIMwpkOT9adJ8
Oy3B9/RGVzGdtVTkWCWONFXK/yt5hgdShEFIZb77R74ieqLd4wVBZ5gV3bV28/Sy2jqcZxutA5/O
mkS3jdEgB3QqYJSXKivmCpWVkVpWwSwH1tB8UUK+wcCwF4vR/xdXJ7LDT1H2IvLslW2HMP7HCSbf
2PYiDWFp9xYnJDHbuWgeTXJMQ+6yxbKFCDoZmjNAPqfraIgsYEi5tmsTzMe767S0zIaqRGottxn1
Ce2Ibb5uYwpGffO/pP42IVwcjnDGlMlPE38tNQYlYj5YHYIqtd8cLAUJY/3/9QAl2aH0WJI9lmWG
9y1jZkLvCC0jxsV0ab/9s4dXXB/L1/UE4VlbkiqiUswSDSLYsbGYVUksTXHt1TR65QjoIMiGJE+C
Y3I0p/7WpPsQ7W5JCS+mnYLK+s/kw46BAT0BPdZlBqp4E2O3rHi06vfdL1BoaKfPBLAr3M2nLGdz
ION3zjz3nU8G7dK0ZfG0/E83BL4pE6DKb95v6gzbbhzYh9POZezQJ64nLVx1PG8HbnnW71za9jnq
PGJf18EYCNgHzJW1eWO1nNoDgrAhgE2Yvm2x0kHZab58PpwwYIs1jbfhWOuOjS8Sm98Tlj9ECKG/
mtZogNA3I46SyHTwLj8wQ7tEDzEKip63TTMrNOO1Bt7Bs5+GGGjJpHYOT2cJw4NA7UYtsfKoCDiG
pl5lv+NUW5PH0o4ORAX6z/SciCM8Y68n/qHfipqjqo60pL5TnWpzn8aS4zMKKlqAMEwLZXalVB62
9xyPv9mXIhMHUh5sm7Em0CDI11NPboW2K4LQJ/TW3TwyZWotyY2mfbe3Co9+xsh5Yhdta8FUuUmk
kCQAHRa2DSQB1XDVnUgfpuKqksowNoEdFUG3y79zZwO4OMWr79MxzbAK+O8bF/zpZydBPpBoOqTR
jNfIR8y3lyU7cOHByVlt7bpAOg6jp3r7+Hq6ZTWQkgOdx5GrorLPz90jFGEeUlFUa9UWQbOVMkMh
SBteqQi6q0aUcfqu0XU8p1ee1C3cIsSQv0fd8Kc2IIGAJ/M0yG/ne1DwQNoCpLjOsWHnLZ6h4ekc
v5DHfvb/UXqOAGlqJDw+pbHxHZ8t24ouseDxxLjMrZWkOZ7CoJU34NaUagBWen2D8rBVkgnm6703
4c+Jpex0hvujvjh1b2t3nPsC61xFYAXaCnOPeCEQljyUd09YOOvuKkKkNobdrsIuJzJPA9ZR5FL9
rzLO3X2YH1JqJpKC2IR+C3IjffAqkP/3qMfhHTYZIKZQylH0CtSk4PD8w297ofDZAlt4rzG1Bk+n
+63Hcl7rgK+hrE6fpAQMqXIHz2+LrpsC9xTOno608qbwvdynHEw9l8B5nenJ4UExT6vDzD/HaWvl
T/5JpXVLxN4zPGf4tnSWHmW/yHpsYSosow79+M6kqLvt10r5zU169wTwuSvXePXlQ1vOxfNVQlP8
3s04PeL7vXSZ8CucoGx+lrnuA+0Kj9utPlWCmz4H/CJumQPCOCe7OkCbWMyX18w3ohRf1kKCJHjO
GzPNraWOCIsqT/qdwPAh4gBQNnRLqY6x9VcFdUfvpNGyOMDbgT6C9k8tOgUTPNh4fwZ8YLMItvRh
vrxnmkzLeU2hXXXiD4QWJqX41oXHiQbsifg63qPFB7C8bPn//PL7ML0jAbmLRHRmWH70glLdyu3V
OEq6owzNjKOc0N6OVgkFYEE2sJ5Ne/osnY/k0mgzbXKMRGf5ijYrXR3sIyvsDci87NjNUQb+C96J
I4nKyyHvq0GrfN4wJWlHGPjhKhe2gVeOX999Y3/JIyiSLAGf+m6bcfvruv2uaV5ZjmSoq7DQE1NW
iSuoYYFncZXufJCaxjuj6w7q38lly6g7Gb8UfacpSC2fjG1TxV12IoqOn2/2+keNRSDQ5MF6NKKJ
P3gD/vpjQ1kBG0KZmbdzCJ6AKtOF9I3LEdFKdXVctYCVxYVsQ12uxLxZyqPnwhzLUoAZQjc3dvW2
xlg+i/0l/A3cY0NhQXCiMzvlzJ+nUGUGyqCiZbpfEbQsw7W8zyUd0EkefnaXhl6wjXOC8Vcv8gnR
TS1AjN5qKb3TIPxmNBuXRHkMyz7q0z+cNT+LWPkbAKNI1N+69lNRn4oDbiMNRmILjO360H8IBdZw
3uudk5yCgp1+N37/Voh9sHqP4jjvtFJqiGdKhoCFWofy8R2Ftfw3yhU8GLL76+MCy9Vl/EzP/tsG
NvIrD++z+2JRUHVF5YlfSSp5q4SMouVEnIYHAimPS1XxzFvlmIo3ASej1ElO8bEgnMATn6gZlH89
KXzAkf03wxeKBsHPDAMMl+qvcalpOQ1Bf2oO3ZtAnnFUfPuRxTY8r+gZr/XOQ1IjpBpZiEOdUx20
vLMGf83RUrmxO0X0D3Os30XUi25MhwZbvYugRzx4aU92B+umnsQJfxM2RsHCdiR7wBeJ1p8mIkaE
94/9m3AdwyzFnbaNfMoKucbxHBhinJHAOdpfHOw5+UN1dV+kEPgVV62Q1QJEHQ8OExUW/Zxbckn4
dmkKdfwFWf2nRnOIGE1j+4LPGPNglnSNjB/PfENkSTQnowOy1UEwLGWPm94HygzVHdbhQaZP10zV
Bmpv6L1kPm7f0rddumcpuFddXrh3SF+MTwUNgz7Smnwb9exIxmyBERHcGl2IfhTpvLJle/SOsDBp
tUmnhAVo3erGunKYOIN2sXnloirIwfK5rxozuGdf7zJLxglNnyIUufSdSqz9heYGRzeDLnLrjYHZ
TXxBeIZfukMhf0YZLpSTZCDzEjIDgTMVxsnuFLFNLWcB6vVqCJfU/snZEsWbVl2VYZYj0Wq2lM6G
gAtVVsRWEAOHrWVUVh7SKhTEnwIrNK9MxkIdkH+qf87OevcN12dHrEf9Xzap6kOHLQLKIpzi5JJF
r7glIbcTVXgOxagYnA0RSIdhoKlsMH7LsayDZRC3UHxk9cLlJrjt/ECmKfoMODe/DfhM5N/jG3X5
ut36XqhegmZEPcw7oPpkd13U74gJBTxtDjRlvP2oztoC8MWCAEqHBKXPErfLueBx4wAzyydOBCXS
qYpyCKE4mDJJy1aOp4UE3RmYWcYL2mRKkpnBPHr/OUbfiS5FGsqsKvAT64TS2aj2eH0jkRlded2T
gVo2vdcbhW1J20swLOe/G/juzQGRqK1VW7FBEDKV+RHoq2OYC527qohdK31GOgmGZ1Ki9WT0mLJa
B+0Od1Cov/BVES12W1N3wNwV6qngapCm8IWXTAMFlgfct3xnkR0wJcy8X9ZBw3a1lkeFZj0lg/cG
+xtG2/0vsP000pIs1iFqljjjLBdk0hJP4Q9vGJgXYYYRbUML+/OLToFiL2BQLeDMr+yFDqupN4DV
Ko38DoryXe7bSU9yZGi/e+ro8DXQoTF5RufsjRkVjzkbOibiyTF6iJYQZVzNBuHvIFWc3dOaOf5i
nWFZcjeRX8aZ7DqVFr3oI0wD3cqNxs7BKYKGBOxb+EzzXsSDc0XGeNk9C3hyQ3qu52P2uzanEGYi
PzxauP1O72Kg56nczYjwF9papwDrrC91ttR4gAmYPvcrTJl8Wqm82URiD42AtuntUFmbFlhUeVeh
/i+8+UOU1Txr7flTu6C1dobwi2cjLbSLFZmUgwWtP+n0jfdmIxyYoP8I60T2UIudaBs0r2/HPadm
we5who+t0F3hcXWZOVVImGlXp+iqZlc5kTyw7j01N67kHCRlrWWDWF4XBezePDgKlzoU3yfoQVgJ
dP8GzNen/9ugZwa9ZctRpZRZw22a0oHDDfdneS4ymj4GmegQTX1F78BrAqUywaa33YeLtE9J8CQF
f5Q19T2orLI1IQ/HO9/udAINyArQqueiGQelqNFwM40/1WiD0hyWq4kWXyin1XeJKmIbvNjB+8dF
GRkW+kOw1CWL8SPSc4IDZkUjUnhG6qWZ3ZZ0g5rSyE+pVm0G3LAkum1xeNkzHW0EiussdiJBHdgu
8eUWvTqL65Qcabh9Z1Gnz4JU59XsFusd6P0r4Eprg+Gka7nZ30zvDX1lkAEVGzktrdYcJJ8fPrjx
0SOkpZ+gAeOFFjuyIYsuZIraOZMU4KOXSc1wie9rQNdNqk7XJqQWH5lI1qkDRu37Toh0bgCC6dKv
fAtuaaj7SKwvjQbRQtc1IH+jZztLojABuE0dGz42zGAdQCXJE+Ha8HrDXtcw9VUnjTqSJLYaZwZm
Ee2ISdozhuxWoQLNDaUAT0OkTuiaYcTi53Ge0pjWegSbAEq0ueoTIiEZZnx60gZU6PRkGAVLeHwh
NoRh7Nnyi96imFPGO6hYC80NOSX3uL0VKV7Q0lHpwH4b7AtIyC9z9W1zFXvjOBNcOJ2cgUuHBvtv
MPnIc79Io1fG/BOsGz3lmjOqBUVt6J9gZFlvi0/tFTgz3d7CzoXId9Evk6rfbBu8CGzoAAGQK4WR
FbH+re+iVwCGyyIAKa2k5/Ak3C6HdEO2JtcEXV2ZiheEY8xAZ8Ic4qEFMgkqpGMRWlRKac2bOYnK
4A1nRdbO/7PEF+TtLBC8a/Y4XlxNyzHNMTI1S5zXyQThj5RU38+bPmpHkgnp4vwuhA+FWZFCBtzb
JsT+S8YIm5G74czcjHjXe6n2R+qnsgE2tj6JZ1SGADnADE8ZgK0Hz08C9yryRRMNy6ZqkUHeutrI
t/ZUiMa63YdfRaysl0qSFUpG3zSzghdr28watmjnrn2RQ2ym4O4dGol7vRhfPXDs1YydxmDUpIjf
2r3aKGfu+R1jKZpCJsX95mb4IRxPQsZgv/wbC+ZljhSSB91Itvlb42xzA1BGJC1DICV698CmslAc
FKZdrj+j+zx4MuVV1xKUqX4cEi+Yzmsvc6MXImXWzvxIWucOwdVChcpJrRyIk21Oz5YmWDGBZz2h
u4LrfZSZY8iryL/JIbhieGsfsn6ywhfnn8OVKe1zVB26Ui8y4k+AC7Lynlcz8kFcBwgOZ3BYxDpm
sCTw/3+X5glTUTqShoK5pe2gjDn0i/VZG35OKLEEPlSyn0zPJAx1wTouyHZUoJZAaTzxNemLW49J
ImH2tvrLIU5NyIJKv1b7Ob+TCg9fSpMx6L542twbmqeP73thPpyIGEIzIgp+AXO3j7p8TLwPAAOL
XF2MxnhBRQZG5zsj/dP+ZTx6S+S8JortZ8GyaEeRFqJ+SALcHSy/DHrVM7Vesm/vB3XweQHvd0IQ
LB4Is5l1idRRZ9N3wcvZSCPxfyejUhpndzA7wc1xxC7IwwF78ih6OIrHU6xQYdOVVKRu1zQXEOr/
/H6lEvWNzq/LwNVZHc019jhvDtaVG8IG4of9EOWe/CBSemf9x8GEGN8Wifq78+LCK2E4TtM29p6W
7zX76p+UuDI8iyIaPAtGeaEyCS8ENk/CC3P2VfO8nQlrZc/IiTHhNyLrh1MzZYByBkZ3Y8/8Xwc6
AX0hoUuLoypDigOJaMG4D6xJoyfaKMZOnOybzTqHULhvv0wJ62sXriY58Zdcfvm/QZvkGbw8R+XP
y5QyOCVqrJgFkH6iBPQO9k7B08j3D8EpV06W/rfyD7Pc2V+vnMPWshq0JOe1UO8hUOEw2ko0Hwr+
ZWKi0Aa4Ci0y0C+a91bvOG/hnA/saYGHTUHPOQHYeQh7O4sqCEJxhbnP3tGfyVxs6s8t/8noDeU6
wYatnsmD6cbpguk4CkRUFPBNl4aYexQLpIfvP+qCkDzmBG44LKwGnsZZKYTWiu7ibDlrGy5sBYaI
aAyzolYkx/l1fK89TrAQzz9XD9emIwsB4pycVPkSVbCgIPQpw9h3x4ZaolKeCnXmMPJh0itxpVZh
87vlY7rQZGNkaidtovy9n2tV3IjuIGL/hmI/xrV8sanQ2O6cz/mrxtl9NsSE/CVwKOWU8uSXrEWd
8HMxRcBw+H5yT1kNU5u7IUVKNWz0z92ZaAPpIkfWg4Rf9/v6K+MKNgUKIBmaTa6V1n1/r14JARVy
gR7qAM8Fod6N9HNNVv8T1ytrsPig4/JbpHkHtbExTWjqMIia4jmIMQFRzFfyZ2A2RJeeaBXUURfd
d/ADTJ9UESA363OUd6vvAycGZ3gn3sUeWsdMO4rfPihKm8/E9PYgMO7yFad/r+iF3M1BXXaiTo0m
H9V/fk1EZHQXrSai+KrfGUFztP363fIEgI0yU+Wq7ckd7lcyHFnIvFTeRoz2MO6atxjjxdwni6nf
DCbmk4dAoi6HHKBlOVMly3Ray25eyS43nPxweTSDNdkXsViPQ1ZNQhfDhtf9eTYBsilCRqvJDudN
O9d4uwwubHkZqPXPWOCCsKkhJV6ulvvsJ1Yz4gMy0fkHZW/PyT2bLQxqqlzFRxrRensSlM7JyHYE
Yuf6dagneR8zX+PN5xaqhVZq3g7HXTMO4Sdu3dCUz/BaYtfkMcp5zfIit1RziiSc8//lb7RdcgEe
fSL2MOGCCG7SjB627AGptgjUxFDW4WkN21x1LzTXNxqLEf62W8JEf9EE/La2eLlGpEdR/sC8iQ+m
Wsq2JFCy5ZwntqjV2DNpQDFxSluYvfcwty8jlUJQVDPBBNwu4wHckS5ZPJa+CSI15n2zOX6OTQw4
XaLRsOorWldEsluoKu0ClE7JaQYma2Jqf64j83zgNFzCsh+CYXc3sAr2rsI+8LT10Lp44MfhdpxG
WOKcuMR+UfxNDNFNkNdun37DLOnx6Q+g2B/IIjBlMLQopwR5snB5X+nVjHLCavWPog7ISFN/lASp
EPwqZ1hR/zwoDoNdOJHyG266lQyQ1jy8keOBvfbyhv1W9l2wK+RBfM1vUw7D/JaOq5i/2/Otr9I/
eJa4iVZEbuHFGz7lL7HCfH1DL0hL3P/m1uvaO2NTDpFh1z+OPeOYqmG9iuy+VueFm1gQnVbK9u04
GU+7r5fvohgHAPk1/peGogxRIbXHpUuLQB2KMM3ohwOzYvrt+nE5u9zuirOCUBvU1qLjBCooqFmV
mXogBpZi1IZ/LGvdvkOB5vtur47I8SsYF/wicM6k6AGGiVc8s3IxRxNuqkbzdCsDDvvAa/0oTSK3
myC3jhkn4FWMMM+QModb3Jw+UMYHL8TqgilzU2NgqeSVuNr00yVibFC9MlKqliJcQv9RPzYaNXR4
dWUFd+50EJPBm7iHA0tIs2QCrkR8eSAeFf5W/O4C4/cL4aTJqPr/IhhTRQmkCOuOoimgFMWN8tkd
h9wgJh76jE4Qpc5cKVJln51mt/JHVM0sQTB0hWNswDM3D/1Pe3zHhigRiwMHmcA1yH+lvBCQ25wQ
TcbX6qPV+teDaQFn/aH8rDVB+44tCXI5YQ5cp34s7KpNmWtHjOBtbvFi6s2y/PJnuWCBoNLyNG4M
/roKZBsQhSLDgy2rYIr4XVCyM9EHKttjWw13cLbaao1D0MaVj7PSPEVJpYxhuoxdRG2AsI1zWu7j
lviqRymlN3WUko8fePbi5ygIo6JK711yKfSPB5BvT46MWf8Xrqa7pIeM54HHMJcXwl62KwTMO8M7
HJzR9nXE1ri9YvGnlPpWaFJPdijOilVmJ1+gfgLhSb6PmQxwHRbSV3PU4UDDTzEqJgbKWsObZRSh
Rqj3j7Z337Kr82unuvduahuxcmx6x/PK+pDvZceA7Bg69scGtIO29BFNRwmO+Sa3ugagWgx7L7P5
6NI6rOoOdFdIT44JQ0BAhvkgILDKik3Tq/ezG3Ru5WgAzikDn0ZMTgBVPR8BLznK8P0enmlxPDvH
fh9cLHBdFyzzaUzEpBnJa52HXgjM4kozSXL8qXpvfxZzNlMuiINx5Fr9vSDlUwIVyUfgdZxb/JXc
6VhzDTpDBATe2HescNXzFPBe+c4ZE4X5pkISD3Xam55G602niNBfKUzxDiNcQ/cnVOYRPJHtRtU3
03IOjCSEOVXD1tliuYvHbXwdiItU6vSCCjcyhGL8bpL99ABt2K1H9ljYWkA2NmR7JFIbAaU05mJz
l7jPvjCCveDLnUg2U7W3NJaoNpISIYpk0BI3i5snnGMhb5sGD0x6mPuh601TLcoNSBe0dj2q6euC
416hZ7xqMaOfcn3vWAqCrYj2lx+6TNSgnDCDiUCgv3B7VcCEE+CDaFWjvlQZu1w5AdDer+KwScXj
kXetJ69OS2lRefVjvSFWs8XLjQgkl9HD62SMcL8dmTHlVx7TefaPiZKsu4EUnZJh/u+R5ZYeKVjq
5NE4pS10p2CVUY+mgjL8aL6vm9yd9ABP4+J5wbbs+LgznSqZM0T2uMJzhEmBYUI5pEnuUt5vO8tg
2Wy1UrszcUqBR4oWvcipWqmxye/WOzaT/sNxZsldzF+mmBdiIZ0I10bX13ilRRkt6iVALDAsJZSo
u0LcQjnA6bith4rCqdCm4b0X8ipECmJYph9mev4QjI0ivpf7zUrQbmdq1ziX+S78QAZtJiIbRuPU
1lY7RDPtCM0ScZHI7BBIO2vhEZr5uZhKRLozjW9p/RFirylx0MS+JsSZJz3kKipgLDWNgdu5Q52L
f8G1tpnErtHdJp+r1ccUjtk2qF+kwgllAGgS7gOV+KOZHBQ3BXyHV8ivDiooF4oiNLHothlW8Dfi
6huHdUKqgLZ137/VErTP+gxjsZ4/a/iTucQlSHH3wfHCB3BmTGhEj4rJeMYRfRfJ9TlYdoMPob9a
tZHZVP9rWobFhEWH3lp30Hy5mYTWqy+qL1zvtrTk7d3nVmvxltuBe8j9IYQX1Afd9zD+Q+xZny58
+3vYA8jImyPVf8gTNiW9+jhmXmatatBkZaoi4gIZo+uX6hzJzJfuy8tr/lfsRy8LU9RZ0qJ/HKDQ
Yv3FvtYEyWS6Z2JOvTdXf+CMeUmBXYHXqO0MkLBRwk55VOMVLkeVqEH/PqnL+Ii7w2QHtYt6fX8I
Xcbseqhk3foTS06O8CLbYb62aHDUYBT26JZ3OuDfQJq1OkS7NZ7TNPZ6Ei01dr4lxzMYSgP6+C5I
lM3OzwNc0hAKV8PswtFrMZchAqX5hE5sxvy65wHJu86A+LqpbPSm4CXSNejcb1I/ZdinDETgJ9a3
fJ3RwB9QBF43NQYd/Jm8aEEwZcNfdTTmpk9pFm6Vtjumsp7NNPfeHyQP8uuR6eVsNI9vmhF2UwBd
DhT+tUyH0cm+v5b5973nWWwFXdP+Rh9y0DyR4klkMJq6eRiwWtCcHAYBT9T3ajwwBgde6DFGenZ9
+ChRnCi9CYY4aIANZs1C+10/3qbOkCtzv+MPnbooggKl3XNKpHRsRznn5oH7nkdXr1/7xcAOAcig
mWyWH3UYNkjDBh7YK5umro1yqpdWQqsxCmYxyNlGUAECm9A+59u3Rra36fJo+Ztq3TArRAXyyulz
SOLKH/0eryzUaD4esGxwRX0V4kfGgEfzGAd3DbHLoa96YqMM5E/hi3ZeFdhtvdsMERdw18cAgLEu
fNk31Qa3EjiKkMcMEReR7Tn3pMKKhoXAgHq/+YNvbdJkryK8dy4qv5ZHa5WY1kPM2X8WvhBaHQVW
7QhMeAiK7rfbJga5TEoZqpqyJ1jvsBiMNSF7orV4mK6bseGxu5Xt3EXyZAg6GU0PeDpAyJSIUmMy
sRkEy3fGOI4LHNBL+XTYW4UIYnBSS6t61utUF6xZ4D/P+mVL+CKIb5MsoRMP04Nv8OrXvymj76JX
IfS4G4eel6MvnXyWQZchlfOsN6SIrmdKI9mOn8UY1b4e4/0Flj7gUF3wFo2+4LGk+hdCmwRp0e77
jFL6Jwj7nULbaGHIQfSW8qrGMpnDtyQGnFdMpZCKvhs6k4zbqm72XGquD7v6+Yh0LD8Ev894I6ji
hRB2X7WfTeBJ0q7V35fdTNBQNW66Tt7rZcOhmWB8zYoHImRp8aQDpfOnsGvE8Z9vS1A6ZPVswyDe
jaBVLzxPaGTuFpxDUn8e9YXAl0doaR5ikGwfuxkKREduWQVmzEn8lJbko/sOruF1Nbk2RTFA/6O7
Z50BeWD9OeIC8wq2tEXPLAukE9/c5RzA4SaCRcKpRiK3468jamK57Z2zN9WXYWtHh0wX3gt/pgJH
RGIincSmKi+lYzwn+XzjyQQpJK7A+fBmYifUgCfndXUITyLjI61gfsHkm+VGZdWnkDbDhn6ez4Y2
KNkQ9+FSoyqyxIKMnm49alPmfy3qcAGQmAjGXQ5a7LqyAHTw0sPZX0obDpOnvLaPXJyO2gYmNK37
4E8BrPNPqdYQ9RVtGYgcvlptLhYtTQmQ3K/iDUrVjIla82/7/+W5O5QSnFwSujoDfS7wTCbP/gAe
pEb3XUCOUbD7AjyVhRkS8+aQmQvOwjUmmxh5wVfzaKczvxmu45Oj9fijyoMNQWEoIszYJdqXzLKn
o0o+d0Leo10zzHnpMtoZujV+R9u4QhGQwnThsUB0icZesarIV4oSRiAwMP461tgHohtEPw9+44rl
fnl9tsGv0JB7NBPSrYSNt15fcOQC0htjk4NHZ1pZ2FD6VeC8zN6aYfMvcmmSXk5foQ4vaWHKYkCz
dpyWu3fIQAXS4u3YytaqD2y4KHFsq4IZEn1ZLRsVqedff6GfpTJIKAKZ2g6AimL0aIi7mpM7Mykk
JT/sL9BDHXffmID+0LEE3Wr91Oku7lu75hQjGpJpj3ST9N9EN6I09/ZAgc0XGx47clgzPuGdUrB9
Jl9bhdaOx+TEFuB3ucmPiddqcUXgCYNukYWvtIYC6wJLkkRu4zedY1uUq3TcpfG3v/L1+T87XyFV
aFTkt//FQFGrR/jjA4InxLMC9Fz3xzXbtnfaHR+hVMKYE/t0nxxFc1iK49mp52nOCLHR8e/tDUY2
7A3VciKw8K31MkjpDABU78XzglJuKn4eeLR9eBsh958ktWxy1bumuDVCnOWOlYgSeTvtf3IXLBmh
TxErBhElCNkdoEoByktLHX1YaxZLGPmWpQC7htQ9eXBNO7tQWDARe2D1KQDZKWpSUjSV+cx3v9JO
p75MlUs8aedLnjGORYKn5doQdBG+XGnSAdiiarnI1kQ+XbK5EQXW0BORTtR9hnuCfRrkWgJvsFhX
DNiYvQmXIwcc2UlxomNZ/w3Qp/kaOXEux6hdGFNlD61QIXPWKa404Sxg5vRBYMs77Xm5pk4RYbao
E4YyjPE2BFwwW5cuD7yLZ57c2KMMTWKCfvln30NVWrSEwwz0fm5bPCtur/n6FcdcJVFMXzaW3IEF
NwqydRMeAPPhoqyjTOJFzxanp+8/N126KtZeSFM5irO4R9O3YeKc9P1NGyS8PM9ON5dIatIT3bZH
s+uQt1qk++9HEMqEs6On8XSTph25rZQnFNTMFbXXu8qsu5NKaSpyDuz3YaMV6abRh2CXU+a/6FJC
mzQ4V+Y7NBOM4oaMHDskiO+zAsboZY52kLnZU1ZearueaUWTlo6kALLsDQPsTBcCtNpQ2byTx9iP
+cL5kEkTPlhiwm7CVQA5KcYf7UnKGltj3D5stgSjrhuxs2M1K0PTaM27hquqhnAAw+7qgs2DBd4W
7m18Hh07IscEPvQ9tdAqBEEpyGncfA3yDxnmrQdUcU469tVpZcnDFRPr7F2alhK4Rw96IMftInH5
6DHdLyEb1WOsJKFeKnh+1/G7QpgWcmEUuMgAwlYBymMjNy1wOF/oy6WOA7uYBTiahEZyELjqq0dT
nwlB/rxIhnmlRtXFCDT5sOsQC21P6gUjMpsrXuX6bOMwMbYN+9/JbLKJtcVmyqeW4wT1noUTUggE
8J9zlqKoGVwFUuQrf6AlZnY6IWIzMqpD/WObcWM552XT0OFvtGHrShrKvQssWRsqwIsqaB1MjZcG
g1KHq9n6PGItIT9rqJPZCUcj4wiCiDD5zaZCLKUFxfkXLZyGlub2b2k9gfWDNlpKacznEzloV5FW
x7c5+nTRl/uTEoMx4NkVR6ekdaBGsXE7JiQyABVm+mNJGLPtCBFhiIF4AJBbTcb6uvz12oNVTNrf
7AMpVEp1CiBq5FsiA//DdI6pjbbg0mvYstrzwiHj9tMtN+3v/65Ot9Pxo8CIe1zRqTNOR98GFB5P
rdRC3Hn5SDaxgoLcY8Gid/TRDp6An+Z2JPe4k3DKfNUNyGal6uPKRmTwIw4jkHkG+f6JHHXenum0
4YaM+F2movIy4jNv88RTXEIn7SJ5EJStwvhh3nyed6H7idD3eSd93dnfFzukuMwx+hIAovfqyOZT
7k9j6epSq+WKxnPrTOLfCem/Mz2BhJnwSomaL3j1j5/l9Xb/Sd+34Dt66dKkmuq9TkDdDrwynPZj
ZEDGSshKglYD3K2qLxTg8nsWjY+9J0ATmyENJ2/8LsLTtuM5hhghuR0Cjhy4S8joTs95gKveG7Yk
aaD/Ww1Z3NXpQO1zZ0PEV3nGP5+RctasGpw4dt3shGJDqL3p1L7SZ/KkvA4FT5WqAfUx8l75Mxpu
ptE+5qOsPgovg2kG+2jkhsKY8JJVCa71kyH+gHxnnlR6VwzPcy8j9G96wjFeGt5Ow/uyc+CFl+yN
/4VVDMUwUB0t8JKZ7uX03oJLg1hO7EeYw1lHzpGJQqkuoYsmYhJ/azxunfhfCH6++rGd2aG4woM3
EWu5KHRu/qz5A4LK7zHv5aZsPV+qXgOB2oxriFkFUtU6Jm2RuRV9yMBRMblWbzDEftvtJNO8ehCH
izZmpOJ1EaAUEJFASxuz5ky1XM80a6rR7Nh0PFRViozmCW7fsOudzsuOFTEfQOEWLUiZ2LXNR74v
s97tAbJTydA/fwylJe0SedRzY/qjoJgwieDVN+GoOcwakM1zF7LKKRkgYowCm4TtT0kmPwYs67NH
taIJGQi0ReTlOYkPu+FoNhmMHG7yDORbosOwcfgAF2RPXaacRsjSaszbhTUddVPalDvHUGEFb4K3
K8R631KSMsNcUOLWamIa4YElMe5AY1+o9oqmNKzpswnh14ndUSK3k82KOQoJvbkfOKAp2W9zDhI4
8S+gT3d4UjA9bLc2Cd985Alm5B+D+tuJ8/K6ktwEjhjHO2AvwS/IXrV2ZL6WbVGcMDGJvkY5EEra
NdpyMZ6+Y6e6RRBdDD55xv9W/fkmVhwABXtfTFGUiR+cMIe+GU2GPfnFcxAyM1ZLJvUSRIsULr8z
efxJNbxHD2mlBJlHoitKIcM+14YNkAXKy+0QfcEQtb/2hOxy28Fgd+HNMh4V+yq32DvtwQJ4kA3r
ITvXb016PGwn6wOzFiaHgyESbyzeL3XlrE/0GB6yEPembwSVdt8Q4u24uqgzTdHf/I5CIQD9zQl/
5M2GcVdG65uRVlZ8PLujuSB4g8qJUFws7BlL1NMxq7xmbcHIxGDLu7iMxf27k1lTPEZn91xkn1dt
jp9rFvcx4pcO0SyEfxfAbHFFjCJwzK7nXoA/31CTU6slOQqgm2rziwo+lRe2eQR0LbyXthftoTVU
+AkRVXDmZIW9ovEfzNKLZwi4ikny/lVZtdvEM+Y4FIvviaO6oOR98TXeHKppsl+BBF2emGgKqZ7n
py978yDqgY5kpjUmaZ87QWAGoikfqRiHMb1Zt0Q/Yxb7S0whVA4CFHN1uOBX1Tybg2ANulRt/Dh9
GuklprIhb+fPR78CuJ4oyJ0AFVN/n1y3yU1jFmhI+ElUBj+/pWu4fYJiyh3nocf1OjTnIAKJNhwn
XBAGS8WtrGXttuGdG4FTFSeE7fjY/3JcCRrKGeBxVMhDdJh6NM+vK1GvS3h91Rt43DqQY2vnrnNX
wmW4SP4ZfGMPYLv3eWG9Jrxjgt5u/6m7fJ2oa0Q2LR54lnpta0TtvUrT8xF8V2I3VEtdpwRt9r9j
mV6xbk3xvBtSB06Yk3sTGWUDsO360oqIs2dHNyVX257oFSaVzaML9o/nPz96b9fBlsuH/pTBnwrQ
HXag3ldfdeI+wSZ2NNqMOKtnlwe1XNSp6/LF1/pES0v8dW6MC07jz+WhMbQeuKWgeD7xCiOTl/mL
osn63dBG2NAbKUXXHsabermLllnHXcfcSbrzZvfdWmo/BWSHFHj0YYoInCVAzVC4u43oz9YTXJlE
YFrNd6dUWPaGGbFWFhyUBZBmZkWxJxugzyalKNqU4Sb6xF5NDCMdtSXiOfof3cunSjyAw2DRjPv+
luXv6uwujn3P+r08+Zo/trTThIaZBCBn0XZ1MHig7WPMAeMuLQecXd4wTW3U1uje9w/s6y0HfkDa
ga3tDCwM5d53rK015FGqEMKUr99pAy34EmGM3YL56jKkDcV2RRMm8hI3IcCalYrEvv4cDvSD3ZBK
9WFRw8fZq9wW6FSE92SAaQVu7pEBx3bWPI9B15Z7zx0TghHRuPmK3GcEXXd4I+VGQJpes8h5imYj
e3frTRE7drNMxyzXMgxcTaENKRGTgFhBTImVFWT5aJprFDL6rtdt0oU3fJ05G2bm7Xu0iqfFo58b
pvHOu1y6o+FJUq4+BeduO/CBdtDn63IaKkH6QI92gZqfaxFGapQXxnqXAPouGTr2tcQ1yvG+Q5dL
Tb52snMeUo/8WBh5w5x229PYCYcLzJ8Vz29Kp3skbVQd8sAUfxCXZnSL+u0cBx+7wVKv0oEhBlrS
1esUrXmpfDvmEK5Fo/RfDbK+P1ljMkzfROSv6paFygLWxaHFbuPVbmMKO0ZHqUjChFGhWXhsfJmk
IlFwaHRGscYIGhV27kUpZMrlwVbRG7VUFlsB/0ZjdDWQdyAfvHgiGx+cZM3kIHiW6lRKv5LIjW/A
OBZGzkRY/2jUcI1nBm4APi7AoMNJMr+dEiwWAR6wZbWnJJs02ZP2tsXETC5IqwPOLEBJa2SnLRc1
wFgWq8/87omhCo/PLn88WQcdkoCRzw9lfx6lepkBrmSBRKKaGAhU7zSyu02f6k0zr1ZVx7QFcTPN
x/cJ3KZq/tqfaclg9zian7S996i43eK7PRKF9pGBhWOekm2epHgYexiFulwNkIBKrwylopFj3NmR
Kfo+nH69D1dhmFJ7Sk96936sUdJLxXYIoji5pQxCBUFf2GkUhimlEAHVAeqmAod8o9mu9bWHoawV
/xVJYl4P4+67jKiy2oTOfEa+/QMrYTFlsBEURmhROETzt20LMDqLR/w0kVKx7iQ3Wsj8Jvp3wqMg
YmZzB08W6jygKj+SQVeSZh11Y6vFxXeo+6RrCzPZ1rzeed+l7b26TeY2fEQIxiGEjQfkaDwYk4fg
0ahWq92r/ADB9RH23vpccDdUU960TIM9x98oKzhYMu+Ikxp0kIc0leh8Wj7X8YTxloWV3s7u6D4v
X/JMxeHmUq3UsYwXgbm8MHd7lrm7I7DEUvbz3GtmFgJBvfQ3grialhZOZ0kun2C2DYlsuplCrTjv
fQAKrVnCll66Z29O+GSMPAL+8qEVLCBWsJ2w03g3JNSFtdncpNp1fVJHUfA2tf6FN3Ulkf8UUgr0
PVYzovKAtHC4HxfWD128Y84p1z7NUeSHgXs3BTZf82OYZcp5AzmDQwhz6a7qtHPM/Hr5nF1kXW5h
jjW7/oa3W+/vMg4AJRMqKv0w/l5w+zwbqAMrYexKc6Vws+6tHCA6G8zelm/lqhrFJm1mdDk1UzYe
gtnbxZv8Ag7vLesoBevevfp/IK/bWHNs6JcAOdhlBe4K084IrMYbiG/mOtU6skrJL1A9M+UPsaYA
hZ56DWbWM+XGPfM7OaBC3f1jCETKllUWT0sKF1PWxkv0dbkz+2Ttjlv2lpwHwItIKBrSuEWn9Uog
KlVF5X/oPUCH9OmveHP00UQyT+wPxrbz7Qf3XjzrEdFXLwAp5Ix1dkUSQL31sSJ9125IGNHyM65+
r1EDcphq/pUUrQ6037Y1FbwiVSkYAq+F63DFL+JL8O8rtBzH7arN1HUS3uyT3PnBnW4mBLGqM0+X
knf8oNEWXiAix9GsIB8nZOzvViLEa6mEhBPueUv33/fDOuaEkid5Ox+J6oJACU03VLcTv5nJXL9o
lHQxC0qZa9IKLkcU/O58MadySeQUOjL+HzJQTAwsCOnwj/Mo0NgCWnL5fYVztPqOwsXAY8Ia4mf7
WXvTRVTo7dBkwtJdVgqBexdZdoWRp0TBy61M7pHCMCULsfb3MTsowPSqr/CTHZUK2J5+uUTXLLSS
ezUEmyMJGUkFhnuj6e3OvlYmthVRg0CdPBnKJIV8SeEu1IeOcHjY81gwgeXmSYdOdAESfL4TA14c
eG/msRYR2C5IPsE2SsvC3HLWqbZ1tFM8oj2TJzoaUMJiTR+ILgKGquydHybqEbF5gHSPv3t2ZeTb
EA4iXpXz27BMH7al804oz5aBK92boHtcxgpQrHqKn3NzwKn+gJlrqXeZ/KzWKDKEFgHE+eu8HHh2
NhMLcKI3tnJ0Ru8x1r19opfT2gfrIdTsK/asJv31fDcgX7c01bmezDmrkiQUdiy7D0nk/sekJCgi
UvZX3KKuvUvUHRjSjjeDI4gbkwZN+bGMqTdIicjm33fZjB+L3xrxiqH/+uGbh08zydPodl1l6V/V
uwUomtxUUPjP8COJ+8bjGtgBh9dbkH+RAMU3Yxi+ivlBIjVnKtCiuBvnQIEO97oy89XvxWgoEuD/
qo5Uwa0gHqjNtooIAjxsYpWFZg4DwyRy0dg5N0AAD2jn+veIWWLH56kabBafGd+sdXDwlHdtXr+n
ZvEPQ9f9TUCxyVp3OEhiyUK8UIA+L+O3em6oZRPgOKgmejidGk6U1ZqUQxKeheLDcXPdw/frU1sN
1T2smX/euNFpm8yHxSFRKPD7Awb0yNnQ2qiAVrWZw19CQd/xXVl69puEyWUv9oJyS1Z2yGBpUTNH
LIcm2pS77y38ThpJ6lSebJnYYqn4JcsEdxEhZQSG50lTdD5QpWJW5C4z/2ucdiTEyye+TzWEsfFS
jS2C86F4L1XHWM30875p6IvkH3UiLBJ/VexVlZu/iBj62ZuXl7AoPbCkdPFskyG7G5A4JJATPuAZ
FY1VE1d6+IjwDYuN4Wogw3Cu/oQrvua3DM9Gyf5OfikMkjlQjqyX/BfgALnOU/wgduBM6e6pCZ9V
H5MOIt6nAY3zRPEdBORv6pB2JoIBKPIy9N5qx3I+t9ropIhpNy0ZUSYgboDWpFl+rLKenO/TV+gt
RZY3ooaffOSk35YbHtiwnWiw5HWqU8MXfYzb3lax/9YvgVVnyVyttnHihtyiYYRdmyZ+b2RVFQrp
G+QPvLeaqW5jsPhg0/19uGdqEC09rKgw3B1a1roOcfEc4AJm7XHom/DjG651Ux7+59IXre3LDi7I
MMbx6BuJsRoaVYv39xdiSQvM4pQr9r70Upcz1rdQQ4sEeX3JIOxifAx8X01CRSJqmizKLqy7F5pM
coQOygJCfpLxeXbhtd1LnxXBf2J14UUHN6VxfDm/Iu6oMJs5t0dlTChbdhrhnFPx7+EAnEqbhN/h
3otY51dtR1cWX6HyC8gXlSinLwYruTWfpZU/XQumf0qK15+0I59OV/aTs+Ddo8KmZGbUi+yNehjw
DTSGkarUXnOkowkWyV/VeZcMXZ4zKf+mgPQlBA4k7o+1NFy6Q4mHWr8GwgstmUyZo9VDmKV6q+IY
Lt0o96E20DqiL7MFAKl+84lUWUuW/foCha9oK2Mjllwl0EI2cg6MuFw7LEF2zb2qaK0ecIk0sG4U
vTpbQ0gjaNUUQ204s02+4SLrQ6mKNCPz2sWviUSIZWlveONDDtiCDEXMRj0oW2Ypur80aLMqYAfg
3ZZBkYgCOH02uAOMiRfZ5WZbojWpSWa68FOPfACgEbTKd8NFzapYA3ZIlExyU0plPN8T8qP4O5xg
Cu3dYC0R0PmTA+4PEVEWQD06NRs/jYlhbn1J4SY4N9KWqQfQG4tNG/0Ks08p+XvHIF6Wz/BqwN9k
+Aqei5vHEUMvyig769Ubgn18x6ZHMkPcQh1NJHxFVIpxQvf4D68M80mksP/pNVWo8hI+49MCG1oN
+TPELDxjwyP2EkF+0NhrPbRTmt7sTp3Zak7P/YyX2oDp1Iq7utAh7h5AUdVbz/FwSShb1cAIpFZa
ldbx1TMQrbUuxk12zWR24/2xfV2ZLxFm7WSw5Pbka7DgkXsReZ0nnS3L1E4bEgPVqCKkXdw0UxqO
ITyKbqiupdfyQConBFO8/pbWc9DiPdkJfTx5ATUzv2wm4lyNI0W/oPxe+ecceJ9HaErqxSvfBCRn
JRyZ/uBRV78s2SxyE73lJCVg2gxGkCPN1UMus09SVYh3OyMLnCY0On+hUPiuIVObAPD7O5XYj7a/
j5Z7AtAX421DjAe1AQcTs053Ed9tGmypsje+0HC2I8kOluKgaatF+abq9dUx+pTBhyy6ZyUgGqov
BjCmAB5yzp2WuFIWhwXYei9jZIwJZdMOVbF9ELH/iAyyeDUIS9ESd6SckQdhoM/TpVIMZUxQMUEB
mZ8A8/qGxN6X/zux4N924vgFFes1AxW0k1+JlMG/6w/QVoRh4FcQW+5fLn4xMCR8LFnkwn97Xc7o
1FhJLL+L1xxlmpSF9c215iSrQHA9rHjjmuipp07oSt+y+pTWWva3nmkb4GT1/jUAFwrOiZVBck6J
NBhrGUia3VbcUL4IyI3Laf1RGFBAF5fuZbqVC8YbDg4f6k2gXRV9kCal/ponSU5804iGecSEy4US
eKueaS9j+WZBqrWXDTddI3cjJnCVaR87wgOQsK0bWpWSgL/09pD5XMIIK8KjPbw6P66n6GfxhrBt
bK2qngSVUhhgJxLdnaPNt3Pe7kHdqmSgmy4lwar+Tavf9qcu5iHnCrwT0RfKZLjPcAkZXE66wCF4
qmQ0hLbfngCtwPdoXi38wvShkeHXghW0Uomiqg9ggGibOAoW4Fu4g2lOjNOEnIL+S/PgHmjhlAvF
xP71+3gFBlwVqe56lzQxUhiJDE/LneG6iVSYuLfF5PSCV7BNLOQ+IMk1+PEgxX/vQZp/S5c24pUJ
+xFcdR6Wa8pZ5pkz5jPczDFoDkSbW9y2HHtbasAG+jBJ9F5u/chTHqGTE6r3pYxPEYK+T9Ats5Is
+5j2GmT5UC4aO2gGze9gUzoDFKxDOEy0V+Mz6GF3uLspP+NFJ9OaOkGEOtQZ+aqX0u1E59efeXYB
ipMkXJqoND142VqRvgZdr1XgHkFwXBIdTYA5L2SI134bnwjw5VYmv+6DOXw7uwHMvnWdfJNkkyz4
D6eYayigvFxgchzBC3bGDdSXsNXbc7pdZDMU9ycHrjEGPpE83t4psT5ghslikbcnNIfF3qVy92aM
V5h+M2Jccpn4HrkSe7TlkV3ezferWIbnK8D1wXfqH3K2Nw48MPY9ArhzbqZfWSvxfDFBvOxzOSc7
QuIbYeu/setfccwkVKXrirIPo3SyG76rGyW2m2sK7gbnQpD27URKyHS0XflRSWEjH2FnOM8lxZle
lX+B35k18hmwSOx8RdMqj8C2+XC9y4pY1mwSYWOyPnpRoSfepurdwRAQ2EANTJ93cV827T3R5DM2
eE8DaawfUxSzgwOdxnh4TVA75+UvgsBMM1vcy55K4bh6FIQTzR9gQFe8+1PIh2ffnZ3ngvi+04XE
ekqlNw8m5y29TqEDCeawNe/Q8GGI+rpB0jcOwHVVwrfNc2MfPBzEHQadOPS/xBjsMuCG6yFyQCMf
hoKZSu6NdNcvanyk2IvUQk5VgRtxQYubO98Mx4eKoL951HEuhiWwN4RnB2upRpxlXuEg4vgYC33V
5xN91PNn/uNOHEDOiMTiiloGw1GHyXQ82RJg0201nWG45NL0PQlQpdrti7yXYu8DW7RT1zBAMAK+
FJXkhSGQD6hrR8O1FRjJzOPVEe/3cpaTdXjkWc8Fd2mFeCsIlpCuyJgk2aQYNu01S7S7xEnePOuk
S7Vup/BRvyN0tMfYegdpa63IUCONZMhBh6fk22xoqDyPU7J/FiaC1YgrlJZXs0+lEu+24fR4hwV6
MAtBhxKzuJfJyFsmsRKQ0MBKJfv8SWxLXTLNOc0e4oZt6NU4RtJ+hk2EaPj5NLZHF04lgQeu/vB8
8ZBoNfmHVYo9JmQofxxZus/jwtxs17sxn8eRjpI9+iUnNBVRUyyAIS8gu0Y7ZBQqR24U8U6VLwtF
v3kFxDdJ9A7+883YE7Y2+HVFbn6iadib44XC27l/q0jgV+6iaDmoW6ixgmqpmljVKlllJtGxD/O/
rUtYeapJOlsT29o1ngXL13aLDoo7fU4jpo3+cHNaNMxrGbTt7ukkC9PsAr6o3/pwcUddkk+5Kw6Q
s3+7Ac7mpWwk8e9Tk+GDe4t4j5KzTax/bOqt5DPivYiIh+Yp2PIajBKlxU39WQhjs4c0ZYksiHP+
icZdFjYXLuoftHo0XnvUWdTg6jYYAqMnx1YpVKSWiXc9pl3kHZyd2GeB9s+1EVy3/uVdkTgstR8g
66ElzVJw61ZIugV7uQ+bCNswskGl8uhuyrUHbj0hzGdhNkAWpVd+OejgsYS9ZXGdeIQ5wbhyo9Bo
qngD3buHWatOYcyl3M/3v01+fH6EXK/lvcJHAIjjXCiy84HU2eU3QyY0uUNbwAeeNbmlFErHiKNv
mK9cm+NeFGR8juo9BzDmoTDNbFhBIWb0+DuOEAlizy21fUl4/zrWhPAYcXcVPqY/3VKVCQH6BJ/4
SIgghxkyYZ/iThtH+QPrCOyPhQK/CdGfHX4sJrtSiTC8zf6gp6euac3Vz4c6uvqcGBf42bJpQeCh
BhauVIygjZIcAhl0FqypPkK9cr9v+u63Ruuzpp6tMtLm+DxyznAVShDxjk36kiKCpohmjx2T+9Yx
dCmmlqN1FbBcxldzMVetcGXkzORjHeMKZF+3aBIABJUBt+8YYDlFA/AoOxuSDH8EDjODSC0Z1LoX
0S0WGKjSFuv9GgM6u977gDTTYJ0pZdWfTEn/1rqrgSFbDVFfrz6CDnR7XFATZYtKQyTPQEU5rtNS
xy3yVqtM5viBEHpu1XNriNxotfqdYo4eVsGgarohBZ0vtdahctZzaQEVZsvx/CWr8zbPkxkq+Zdi
+R/ZJDUnF66l3qzURPEvSP7xXxKKW1XOTWP+Z7+vX8Ra/MSiQjWf+8s+NR/VYXZbkYgioGGUvE5H
7P1LsEBeAu86eXnVdb97q2atfBT6XyicYyb1MCQP/RzdH0mri5hxMqvO5kNsYL6PIZxbJnzFjxYX
HIKutXW/Yur2dCIN4kZUd7zqkmZKWnj3mMIdnf9Q+M2A59PSKqK5WYaB+iQExYlfckqbxbB5T2ks
Q8gmIjMFeRV7pI9BQJ+HcaxlGhymH9ixWQOqYxl0KBX4iNE8L/0v0CO7a0sylhYcUhIeSubpsAri
Mno6Uewy4dtasJldx8wqfiry89RTwkZto5Yck5Ja1Ipa0O32lTF6iUPUnehSZJ3yWWIX5rrsTeYr
EvGG55UGV+3T13zRewi9xOWjfghDAF5Q9JENarA0Vs5ylxp9k5I9Hyn9yf23vyZAb7yy1v6cHOrO
wc+GTuh/bytvRmwF1PQL58O4TnoBCPhwAILoYwdAuww++QC8kBhb28cprCrcPonoFzlsIQAr2IyE
e5EnILjuQX8NJ8TSuXdHoAzmbi6ouB6fm5/GfecHyfGveppr0E5adBhJ8aQVkvnfZIWF0EwVrPHX
Lbcv0tAkymHJFfFjDGN7IcJXA4DQpTgcLykmUu+i4Jf0Pij664ScOw5o2w86eOLxtBWBDUCBjv7W
5d+q9rfiHo6bLhP3XxP5Ti1Pgner1qgA3Y9U+TLF0G2iCZ5lwevo5Vnf41xTWAt6LhtQs7WWzMZd
Qgsx8NB0FFfyxKpjdHpvXsiBGfUZThTf0SIiESjl6Bd1J3ukRXu7RQr11qC6DSm5jZo25yhzWyZA
AWYBmtjOwueKxl7qdIso1nt+RmaSEVFwlqZp7jeqmitk5eVo+GAC2UsEvJwgS6HDRkcheGmOWdd/
c0CkIMG5z1JtqlZ/k75O2qK4BP53utdu5xK5DMQwbSXfuNc8LZbgDGg58Ks4je5j2RdOIJ6atben
YWSJPRdUcGimpcmL6mU3SwGV5W+dYKMAiMsvWHiApOFQbxlmQRprSKCqiDA5Q1sCzoYIXnhBXQBg
nkPrfWoaqQl2TtD4Bigd1Q7KwJY0U8XK4aFUqhIcHn8xMgBnrk8tPJ8xgjTuR4dbYpJigxLq7Cy9
W1Qxda0jTeZvFEiMr75YUwR+O6NDnxb+T4vydJ5fGamVvFzkfO7OYA4oIX7ZN9+3EPyjklGAHbBs
wkbRX5d+v553CAKxJOzyeTwb/Y8SJE6ynIPLe5e4WV8OxzqGV+7QJGvd3LbypyN8ulD3LD4mSk0F
zDQU8Q9Z941f1CximLCngvJSuLsQzaXlYm/BWJOOnL2E1bcEMZC751sOMC5IUo+8kmEqU75+u/GX
Qu8WkyumRrXrjWM9hKgVeP7CRXSPLzoMcEcfcdHIQ+oiO0hI8C6idQ33vV8GLMRSNA1QTc8ET3F9
aVQDc0daSH9yXH5Ek3wasiywv4e3hSR/yMEpfCpTX5s0EPjxito1utixB1zjU0YvNjkcwfAv9YCK
A9ajRC1N1KYHD3rLn5bamyciwLO9nNeB4SV82+X5i+pDE7Ns6W+d+zzVo4n80OK8vWptVuk1LWrv
PiT6JALo5CFud0vFkDcBLbMXU5v6sO07xr9+ksLchiFqeB1CXcdjfTgBigYKzX9vry735bgyev6Y
hahsaCCRFFucRu2s4d9s00YfsMHnygSFHKvoQ9tUPDTSqdyzC+tAbFiSx3b8ODJLzmST2/sewtuv
SKddcIidWJ/1PORGP5coRdIxLMKgQh+GWp9OTIQt1+r3TbDrBMgavI5qKwG+mhLfpG0bs7aDTrvy
hb1CWTS/l4FNzPK8aiOkuyke/O6XysThwUqpsxBaRdk2U0VjnJDxpjz//2WjLXzpm4xw5WWFv2C4
bs01B/Sfkhh4DFNvQhWgObphg2wBVAigX5IrIwy8sMx5KBWbO23zTTiHyRgHfVcSOom9G/4kS7A0
pGQgAqX9wqdmrrFvJ3Oio+A4maGmHwOsy49EYAI6SRn5Dhmp3xl2iGege9afgXgzATmTqMD0xlQY
kmr8NF0fMNYgXfNgp9fAhPddna/M8Bo76lw/Jq4uBE0wash9iALUE372bKM960OTV+y+U11Txbxs
7p+NCeatJHqq+Qe8VfcpNK1Ag2AE86N4E6hU7hIQ0Ta9C4m1ghNH4VGHMwUX1msOrnth21KSS5X9
+tJSmGj7qdNPodW7t4d7tgp1Z1gM8/creqZB4W71ZXZ3suFiEsygF8Rta6cP6c3hHLX7OqW6apG7
CTy+/Of08fwlbKmTaFb/dA8GT9vMR6mbsvHmnD65RNKSAS1QJsMbVj8pSd7PcU3AyuPPbCwX6WdF
3tSjXtxnMB+7/TBzcAkxwEbOLXaVeNxqYRGuG/7Am/MvH2/aoJoSr0DWf96TYPcw/J3swiv+UW+R
Vk1GJGu2ii0AI93oN+8QmuR+f6YzVu9LIfDkcYl1N8fRkGaA188DomaJjRT0qn9LaldRKo197Wv4
ePPtoXepYjywBHULQw3PIPH8g6QYH+a35olrcMyd3L5dziETs+2JT8ZoM/snqZQ/9Wf79L7uJ5C9
W/ca3cQ80bhZSClVQ7Lul5DYhQB4x030Pi8AhS6sP8D93b0abAbJvf+iSDPsqtsJByeXvD0hpNDV
gUtgRpuAIWHUZezvIQUcQLp0OGQOJqQjwLpS1blxgZafT4tGWlYePBxNxNcUWMYvm2jnfrGpGDtQ
yh/FJ9Q2jgN34laQDo6VBCNM3xhthB3eevDpyoaBvjmUf7Kkof/R9vCWxjV9+VcYYIPIEtG4X6wC
kdl1rPaG0cliNFS3YuA6Wt1mAciPpO/38Oql0hCn0kWFVr5PhktoUDqxNaV0BZxaomYxTIGsgeuh
QUumv85YuLdaCEXWMzxKjZnkBTLrpiQA4as40/GG0e7pBSuDy2TC++oGrsVSiKJS1Mk5VbQVbgwi
6Lus0vL6oc12S1V+5UetqkFR0JBXvwrUlMFJFPNWck/qANVvlAYSkP1HulcHGSb0A6yziVX5mUHF
4NxFLxtgWY9erpNjDqnBhExQdPtcC6C8o8chOZABj0i4IAr0nwhkQBhzwA3F7qT96zdiEhqQlQEu
kGdCUM47yzzyBq0FVM6CZ+STrko7MF4trldBRW3lccx8BdjfEvGvu58GQf0xmSoAuz4rPmXMAtAE
rCpN2N+KHuBGgomshFCeKv0RovCRj3VVmP7rHFsuzYMu+2lwemkScfZX6v+FEGLaic9iuYOp2kiJ
1Hc0hMLDEbTculeLOqtJaIitHaIU7AzNbKKkEGJ4hv7hzWigxwZMUVoAzVWbVtMRNb7iSqFNfuYH
7IEwnOYR02MynfQhIka1AX0RWhqBqMxDCaPL75out5jZMD9ueRPQuwkMazPVB3a1jPlT/ss3Rij1
3ygF1RG1oN6yLnwOpnxGWcmo1Ee9OLNwavPUWi4lGuan6LKEI6bgPzzVxN/paCQe0B0YCRg3M+S/
WG0V4E9ItskCjyDDfldE1vJiQTXPUJFquYnjRmqzrXZPYa8IBBdnwyVBuXxr4ZfH3JitWZ56BP0X
qgCJqQ7VjaW6Eb2NY4vyxLE198xA7uOHHn2HmsoukCR9Uzs/54epQ8sSA4JDBNiBUrjR4zrAmptz
YLlPdiQwgGljSHux9zzt5CJmNQfJw66B7ov96GdSkfPKuMcibim72jcB5RvsSMNUDMF7gbLIApK/
Rr5+OiJSetz6XFfQe0+O2TCak5s2I5q4X/lu32BFF7BSxWXNiPKtAqFoisi0WKiEWXIY82zNypf+
MGfUfvY5kzHK68xx39B56IjWa2QWaFBc2ZDhaHhWT57I02ivatsb1n/7qLsUahIGdswI5DVMuYDn
XdnVwOIKFHiOMJH0lh6Vu8p/ehXjbbZ0xw/pTCbYhYnqVcmLehZz5EjaZR2+pJllwG9bX6ZEk4uS
Z/5vfzAmGBuGmDPaup2oBHI/1noM+XuUtmEuyxnL0xeptoX4UZDKeROOklNRZErEYKnegBimXMpu
mT2rvGuhyAsGPIYUrNpF5iHwOHK7IxxrSLeEUFahfcnoRgsXSva3XLtnS/KZ0qQ9z9Ygh2hSynJ2
lAeECHC1vsPxTjgB2i2kF+Ln7QX5yxQQieA/Gk8rsHfnKtao1QFKNAazCjQe5t9ofLR8tFbdSiY3
jJVlYUlTF1ZZdJ9/mmnFJFPJZQO33ge13ta3x09h/H845pG1oFfdauHZHFrnLVe73fonWlq+mKkx
KOXsPJQPKrZ/OwLDYIvelF+vm/8NlC3was4IBIa/t8JajQBlX4U1CcfHP3fX1Fc49mqKwlz7JAj/
vDwo9QUZzrVSjS7PanUVovYmsT6lPn300YhnedQYiYYH3OeoouWhvSFoZaWPkhtC0gv7w/Iyu9b/
zsIJ5Hk3ZLZWnQ7l2OISDgR6+WVd5bgKpq+QrAui9dUOsS0j7ZaemghOFZiwFcUZkqC+HrbCYEo5
Uz4zByZOnww0+KaYOV/g3UYIlBCXDvKx7tOGjXuQg0JCAmDuqpKSDZDXoy50e7WLDWnuzVf6pitQ
wIBs0zX8KVvYgiF+z0pS1GnDC/KBAy9vaaE7gJIN8PQgSx1q0B5UYvQBpQLBlKsbPQexxNjdktYL
/PdQWYu4ABvdLf2MXVQzoAweLdeGnr2dAsVvHZylPiZN0se8IM43q/rzzS2/jW8WcnEgeOAsuqXo
5cCZJciP6V7lohSI9fGSi8hNrVSeHIxi+dG/Epg8FfBAwZsBUWkOPRPegoTd6qjKgDNDI+KOwinl
XO+fseOflxiOw/1ZZtkBKLWqUUOp3rtVl/05meNYMLkyPoIo/llqPcIo+ySHKsb9H+XV6a0HNg1s
J6Eifn/3OQ4lPIphFGCk5/8hLF6cEugZc9wx5kC4DKp3zqkHLyjciaw6pLD78zFObgKQp4WVzdmN
h2FJKonaKGHvN2Dh+RObTUnlw1jRa/bIRedA5s3HrMC1AGKnt0j1H5ze7jKwW1J3rg2yMe2N1IY0
GCbIgrlpjGZjJzcniJqwbRW4m199Rkmx/gCe9CW7bjAgfCu+soFhcvPB0OT0rnIho4ULkheOhC4W
njAoVEIweD7dDoKW999vh4vylwmSXXujappr+dtTsxUZFSdAPO5lJNFkbOTq+5dy9jFMfV2pg7Cs
GIl6bonaLKulxBsycGgyk7HAVBG2Ry0OLBDwNXyTYN7HOirM0fsOLdM8mtU73BCUU5lmr57xzIRP
KCJGNsqwNgqyvmVOoCQAgNUdAzQ0Df7iwN1CX7MSXlWWXt6IbAL5ibA8EJyiTuv0oVz0AbOIs5mk
W11P0rOcJjv4022vCDFdqc709yGTs1CxdHBtTdemSCgAS7ZFXg97qcoBvURQTK7fT2SDcRe+to3j
W3OLgZWTvzs1B6Mym2UemeAvtA/TToX4ZYHXYCZ70P0Bxx/4WLJOv4gdG5FWyPcnmdUmoVj/cQMS
CTePKhdzDZnDrB/tStPn2DnsGYPggZZ7N1qZ2RGOLLqMezO4NgycM5HQp/e7NFWru1vsojXonzEa
x+TPMDX6bQb+LrCiN3w6g32I0lonuTJRe6W4zUGqUCtjwZGzQrbzoCxtFXEBaP5+Gvo6dfCC0qW3
C1IONWvJGnmRT1JUEG4r0KKwLVePrNGWfi6NLxbXtZYo35SWvsKk44Xux0uUxctRTSPwO1+z3JEH
+21zLgzy1LzBCcJ9C4ioQovHARBNdsy5xiUO+IwI66KWVXDmb6Ce59vLpDvKfCt8b7MimXYIdYZB
t47VeVtQboeVBg3UDPbJ3OJn27ZLmrZyn/DBxI3MHO63r4SmCE5nzgUNAjX2XoAXehYeffBhgzc2
t9DRNVpMwyQD6YYwf5lqPaf+eyFyl4qkIa9GJhaw+hNjb+QBR//1wtbg3Bai3uVpizXn+M0rhd2Z
eAOljSoc5FQyXBwyJdUstAtBft020yp0HB88VV92jiY62GHpfsRC+j0X1DaFwXBGmDCYUroFEjuW
3sKXuz9XMG/f2aA7lPLryhLJYF4lLcwwWrvLHjxG+9U2Yr0Q0v2/sh0P29x0r7+8rdkhNtnV2koG
ObZje7nwMNJ56yjPIPyHcvpm73+iYBuBbROAWtF/eliIXQD3BknckYkLzkePsteDT/cWqkf0fqgY
urJGo3+UkXpirm3JRBhIslw8SqujrH4Rus87zwWALfL4o11vL7QQfi8lJbX6SHThRNWxLsFki9bq
4xKgyvSMwqkfhmit4PEhxuLmI4lEOFsUWR+6D1CegmRu0OA1kMe9o2+s3uyKBPhLqsOZliXPEajm
xiLRaHYGW9J1L7rxl6B/YmEov5ekUNcg9y2lm97XT8azK9BpnM7+DOapOq9DslpSo36OnGRCteds
PiYbqxdHe0uPjwjcgVFMK0BO6NW6IFEhNJ2K8QzjeLHR5CAgXaG+LKPDLeH+aLJPuUe8xrdSrOu5
mPkEgq8oyfaUXHiOREK9G6at4T+fVTcYJTU5nJDx7TteUN3Iso73szzZAFkFs5ghvgjsorYgNLCR
D+OSzY+LH2f8p8AkaWUTVKergnysOOtAbaI++I8VdjJE09bWjeYjYIUt14N80d+rl0sq397HgJwb
qXTD5uD0hxcsUxwY9ev7b0bxHKvo0kpi6AvoimvJSFdjSB4H7wGBff2eUfEndbIbe6dZTFrJ/TFN
/L1LKarjhrCHNdsX7qhdcVpNQ5VD2hEWNPV6n92R7V5iYYUK+LHt+pZV2q23ZWtzlnBm5E/myIC5
6uFcmcTWMp1T+YPCtyJxI3ONGllJfRQQIwixdmDcGMMVVVIdBtlDTmVY3ssvWvpnlJEmMX/vwGzC
gYd67k/VzF1/RGH/b+jfUuYe7Feh3riYJrcWU5tbnHVoVa/iPFTndhiqyYCmqsC74spwpzTM5obr
EZLs5c7vV0cd9Md73aGkqYDbT5wVLuvZLIvO1eGwKEo9uHLYTJxz3ZrEAIZvfkXt0tJDwLhyj/JM
AKKf8sj+fPJqrGvH6vg4bvpES73ZV5rStdytZaRY73aBgS1Pfx0l11OQgzetooj0j8lv4htwIAL+
TCxq2IhBGSvBafkCieEu7h3SJx4ZApOMdXkPSLVgnpd1r176ODcpMRxPMeyCbdR+dK52ei0zUjqg
Koye7ABe8rVfRg3jpFetqaOxyk84lK1iaC6rRaLYoi2iKbEHGmkYKvs+N1QuOVXaqmTp9yTJo6d8
nexaZ2qyfuIeDl7wj6i/a/+MxxhGPgIiGbkAPenq/NvBP0Tunsi6ffLzPQL14yKIgfIjWtt0IM4c
NQEPyUM7e2JvM9ENt9s5pX/y9NnkvAcPdzdnjQSe937IANXAPjnSNO7NlW208CQ7YiUCryigf+gM
rEvPbRkKsozxA+YeqjXDkC+Wwe2hlaLX4A4d779TuqyYfDtJHyt/YDqaVaG1D+TdjLR3z0EE04Bh
4Zb1vTWwLZesxVeFul3FLITezLp5ZyDYRMdArSz4HBEgB1iRQF0nItxChVQ3IhEUbuli/HwA/XcO
1iZXRGrmkxYc6Xm1Pd5H4KbDxcSr9dFSTTnB1Rmj82yhNPp2KDK1//lBzC71LM6mEcEz+dv6/sj1
quv0W9dGoOk0fveoFpa8R0cUduj47CJcqE32IjZ1wSpr+D8Bpb8JpOFbSk/0zti2rW+Lv/M6bCT3
fbAGSFcaLqrU1HQrXBJZtLlWslImyJzt9fVttpln7xwmlpqlwE9Fih4SboZso0qct/hUEt1JTtMG
GxZ4HDlThmMgYMKI9KSwJiSF0ULfG4AeDdXdXm388FkQpPsFK3/Pij9uTFlTgfCshX91PWp7G5Fz
irFP++dS3h2a1joER62YZNlBeWOps8V6R4AQqR0/Crrap+X+iKVJNEdx17q9pR6TUweLFSrkvZBr
xBmm8iy4ns1KrF9g0gSYbuEYRKuMm+xd/CcINH9yQ1hUtF1guBe/QcgTAIW+pAE1f6kAILwQ2vL2
9TSRjzMeIOYkpiswCy8IQnIJRiCD8d3qozzEI4qkzqMEPo7RsOkGU+gX/0m6XXhintSndBTKNPbF
VPu3TwPQIA1c0IO18qCXCv+zxVMdSA68yfOM8ef/wULKXKImB79z1ErNOAEn09GbCzBCNK7lRnBa
zUJ6ZajkcaG0dkXTfQcqVgYRr72BVmDM3I7S9X53M1BULwjS0wmkZExprF86xlP8uvpd7NTalwa5
E6dEIYGegYnQ9Pku4+uV2oyXvwtzRjwpQ671ruDfup/zEp3YzjIDmntqXbr+pXv0APTo/N/ElPP0
xhcGdzoApLfnbQ7yaMI8TFBFXUU20nx9dVG6Gab9bDdbukyZZu7NwVAUxly0TslUghXFC3z5zYJg
D++W5mARKLYivAieMUX23bSCSIrKeF2jWE1G3b3IgbzYXRll4QWFHkUR6wpHuKDysdDyLyBhxbo+
Bx1V4+aV+sawZJsoV+JtvdPLiFvlH98ZvMFu5A5dht1T9lDm/Vm+O75IyVSjKXa9hYGfJA8SeHOI
PrilXYlctgun0GOXMsVMo/+oCsgVO1ieBVyvW9VsnAdI9XdKr9ardLsoPn5U57eppYUrqGquSW9g
zWqGw1rQWCapoX7lHMhnYgD6DGyiFo5+RRHOvDECbXoYlsKfrMbguaRB7VvR/6zpXEllOzOdysHo
iyn/Twb7vhYNVY7Gu1RdvYPVUfjlMwZ8cJ9kjcUAe4F93fZe+RDF3LuDEQ3WaKwYipiqbmE0xxuC
HoQH5O2XjjRfBvgOjk/qytQ6AjBDFO78lDWQBEF+5CEZNy4yI4ZOWZIMaRGHA7rcHVk2afvqecXc
IjH7BHZqbURGBjlAFWCUunmOoC4xiD/5zUKKSSIRyDkRm52b/6V1Cz6DobD5x0AZ81htxfkt1f9Q
1wWJWlyFjWYHxca/lAnhjbs2FGcM5B97YQxCsv9hRyUIaXQYCRw55FfoPr+JzRF59kJiwhCmwmNW
Sj6Ab+55bQtSLqhS+YuJnDiNbRy6/ufYcvcElHl4VriCrUD5K5JA/Hy31rAwGDS0NYaVNztRE9JJ
4730vuKYqmJSR+W5Wc7mUn8FkmoT6xSDRLdKjSvBOwTBPDArAj6A0JRuaEU8SktyL/NWTnt7oh8t
DVa0W35PiCMAIsrIV2C44N8yHHgEmhTp/16npvfwcQ/WkrtTrrUMLNhV24QuhjUPuhXlP9s/4u8D
OP7USNUam464eX7HvgA1Eow74Q8dRw85cTWrhaJWhSTCfimz7tdABBcwf4770NwImSWlVfMrPtmk
I/pJnwVBKHti7TeXvwFetgAafxVbmahbLcjjqVrbYUrvvdoGmzf5k1FlpdkJdn9ByGFEMDFoC5py
r1uT8ockZRBtk4GdyS6JOLclH1Y1LYIY/GLXM9rJr5irhPmN8asrpfsZQc6vQI9f744LzxEqxoVR
DWAwhegrmMrXnN4jlDyFm+2dGckKAJk4kwJ5Xf+CM0fbPnTKzPa1kKmjAiD+l7SrMzYb8WSnc3oB
/abvYxU1AiqN508is5Y4gqpIH/Wn3rDXirr84waG/EQ+z0AsoS2Gq0Re5HMQSsb1WugyEtI7N4kw
J0tEnawzWCGThGHuYDl3voFCNIEh9/4rEFd3M+hr0AlGPqb6N10fvmTYDUWDWK0hZeVYxs3oaIwb
28/HrrKeg5CMde4ta2pP4fpqCBoupjfDCx7sfHpDqVJduXcc9d3VHbbbrdHUa47BHQHqaxFK7php
voCGLgW0vpUHv3NIeSlgjlQmLaRX0h+6JcX28FiyXJTRpQ6Pfp+PG2PH+VM6n+nUeicfB7D2HFG4
2k/HN+HC9Fn1AuKlEQY6zNxWvYY6xOL6Ubsnf5mccQpOC8+bV5PT/AeSZNR4aT1VR9wBKPmp5aYS
NMVzQNKumc9GN8zWHw7Jfo/7aO3HFqhk5bBvjqcAitl3No2GPhARXK91H+3C+5MMhJPWsr/xjeJk
eTaCqa+O+ceJkvQO+TcecwK3Eo1E4dg6a55lUAGhTQ4M6wpuoB/Jk24PQNg+i7EtqyTbf4h8wSXj
grITFdljMxVbhTy5cE6wix8IsQZlldMz5V9nFA4I9pch7NtS1ZWrlWTz5Fs57IASi8vay7VaemEZ
fryWtykvF0J2lQj+hKiVQ1NQqRyRYofVzw46D1vAeC/9ypSCrJewfhf2Ju9jJnZd1+nlVXGidYeP
97j4xBKLagiz+hftsSpTLaZ+eex+geiufvJ/ADL31JsUeBo0eJkU6B7IYdj9Vn9QuGjFCsKv64Fz
zi3AiKPeu+SfTVbwOOhrloXmhluL/3LjFaLaRcc5LxeQDXgst2/YeRzw/aHRuOh4dtxU6aRPZPJ6
BXiR1uAca2HERv6Jn3eLm7I1RkjQMyS1RUsY9x8scqyqReROI1VEmp8CF2Udzz3A6MaS7doFODf6
PH4PhdsSgmYMQWuv0aYl36XFthv1hB7PEJugvLNWkG0EPnJ1JWrE3D8/GYS54JSEZIGl+0uehMkg
0ceM4gwa2sngLRBwqQ8XRsqNyqlLlpqSimlYqfJJwbj7IB7dKO/EYNfvu0xbhUJeBA8TxZpF8dlK
lFNqXw8NVC9W5zpGV0aO6gl7YsIdIIXoh/76mTXvsDV5os0nvvH3NA4Cia4xWjjqOmFIHGpTFWDI
+rxicQ05n7HVQyUjCDUvDGWh1+7ZnTohs708TgX9fXARZXzx73ZGPPtdabndxeLRHvJ6QfGYQ1M1
3eR/DTqliF5SIDHkwIrVNQNnHzWowgfKEDQW9ojUhp9qlTtr3mmEj/LaxVyJUTtqhXDzzJR7++g2
HQrnlWp7LxzijHVnd9sOx958yP761R1ospGxZ73kNTq1mc+AjJHaCxVEK7iJaItiEXhevIZeavaT
Bl2pM31Kz8Y6vKGBeEIUyhMqapij9NKuICfCkZLBxTRNuIlyzrJxCDPsTYTyWPRi60Q77IOa7D94
I+w1AOXtITICojfdToY66c+oamtdTGVkdI4noigIPMPT9bCdM/UWPR5rIM7ZkFFYOYtXs4BikmnW
yoLbwnKTvsbtOjIRKSCpdpLWo1R2pgN5FYNt/76W+5uRo9U7+UV5MDRBXwKJdt1zwyberAfh3F2w
kFnDoSHc6rZw5LlkvXtuGjiCqbswSmhJBPVSqN61MPJLzcbSrpC2k1Jq75Rk+i8OKbqgsn/RiHDT
690EAfEXXXxfL2x5hn9wm0j2+NSBQfLHxGW84j4G1Z7khz+PbmgT7d9F1Qb/ejr7C15FWVtJR2DS
AI2w+lqdYWKH1yYeu7l2sHU+fb5PeafrItWZdJ7WeZ5O8y+KQJE48E9RcAeAXZLous6eTQzg3Iwq
RRwFGqJHTgMfQbXPju0PCNdDk5+WkctaO1wesTfUPZ69iUfAUhEdyCbXj8x1h1XWLrZ0gQ2fCn+D
CYiiHwVQFjzyjDDSS/iKEouJG9BC8iUKjoKDPyAASB7O5IqriHXpUl+Ij+/hh+XsbjMeUFz8f8Wi
Oshum4CBCQ5nJXGW/INgSGQcB12KiWzzVV6Nr/SLxg39jCsCRZqIOdBg27g3Co3s4JX0qJAUHhmm
jbLkvQMHRAs/YX57AEPUygpNiwxkdDqCDPRZFm1y6qoCAepTHr58WhqKxhsNIWI1yqezW4No1upP
clJp8TAnqGhQYvyE5b8mibb02cehsrahlG5nWfXZjeE0jH9aeuxB4hf50vx5eX1zP+vTHFpaWGuD
2//MGgd4t0KQf0GMsi30SUztGH8CDRILS7KUsadAv0VA0jdO+rGyvVWDMFMQxvn6gBDQ17Niw8Ib
SWjt8lvK1EgdXHY3VZsOJC5OWCQIhEE8PAg5LGlOAyEwyrTBS9epYUfuQgyBQo5wUg+R06ULCurz
XarS+U4b3nNiPZVihfAH5wk+1W06kx8pB2X/x5fX1Yj7gqM9AUuyEyeel3dOfQnGGFBxsJ+k2wIJ
okDg7ebhQNicqxNzv7wRu6dKdfTkfDzvnZjt2heeTc/wod59Om1VWIQEIETLR7MWia6Assrb0CvG
EMeMGqUJU9ZFxrWZHDfcucdff7BsPGzHVqCSw7H7Opa9eS1t/kTG1zNHMTtfSDIFDmoNUySV7crD
hirm8/C+d8hE7jUvLkE/ZAfXyo77Zyzs2WFfO2nBce95xJBgMeUY3cHm9Q450LL0Pd4LawzjQd57
a16j+DDxQ3UBCMxvreeDzXPtpi2lu18P061QYqo5K3lAhAWhflLZxM8Vsm6xlxef8KxasYsZcomI
Hwy8dIgO+6jsPYcxnSqMXkqJaLkW2jd6EsdjdJKLZ9h1xJ+Fz1/w1J5lXsTD07U++hFpKRg+u+H8
xEjYsqpWUsmSjPGLjArTUsgyi0IRK7AVFA/5oH6ATZs4nuAfz7L2EkhATXQTMBPlS1zwa4i3Ax2E
v2AEkYnqBV+pcdRf721MAnw4lH+8Pf4q86PCOlVBTPAL5yQWppZDsxRKPV3ivitV64T4q5A6JNhI
KazuxFC/oI+XcmMcAPaTUgkInutLXoAZfWVHB7XBSVfzVDhui+/e2TwSYf1BM0qtylHxW/M28VcP
MHxl35GiXomTixmHxplnWfzCTpewOMa4Oa7JuJLGK0EyL1eKrMeZ4evttrYvRvO8Vdjlska7ea/W
kDGfFtm/Rb2ZWZ+xlvtV4TNuX5GrLaM/7K7i7TUHpfpbMpiXNmRYy1wsY/Tg+TwqDp1D2zGoWwgv
aOGLm66R4r9sGKw/VpYEJTNTNmCSYAz58WVUAR+SHHW3NU3196WLv8wdIsUGMvwddWqvmbHOuD6B
F4/Cy+uf3j5Bgs5xDgmZ/WzeChzqoAX6P1M31bqto0gaqY13xF6ArUW00AMmJwWODVOfZFjeeBho
IByDcwggEhCjuuV28fC45vn7dz457FcFD8a4bzPi3y3LXrcUlPjvMsH0bzj21ydvE5VhRdtDyeDl
anOuUnwCK6VF+gCqxBD+nqp2QzLgb2aLgA6JiaUF0gGxozLEegmnGcFLd80wr1hzQrqbPGrcqnUM
XTLSr50bM7OVWF9v6ytBOM7a04ehRqp/I8KiA8mvfC6u6dATPeRfWwYxb5yV1vzFIiHcDUYQNXd7
R2FKZ6tBhHPmC7G7pyS0dGUR9Gw0Q5DCv8/2Di9UdsMwsce98QB7AijRHadsAYlidXj7LhfTxZ8X
k240/MLaoPdwsM5j3xIHfMcgpz+hKKPM8j58dFXX5Cl5EZ3A2fGcAueJjmtgBUdDQ4pmbqkHofZt
RQUTZlXG0qE0DBBk5YOsIUkCCQAXzGNGxwcrqpAn9aE36GHfuq4xkyi62KZ4pVgQw2v9vgBd1Kuq
QMI2DCz6SdW9YdHIfAyCRgr6y06slpzHi4HnX5QspihfVcB6RSm88nMK/++Hu1RC2ODkVT7se/kQ
knZhn4vkwHZByDtgNFUTi/+KMQpZCbzSnDERm7V5KQBYAJHmmEPHsIeO5WXk0bNnveuhiQRUb2/P
HBN1r7qM/DJT55FBfWViDZbadBqmQXBqBoKL+I1eHc7Y6Isaeg8RkGtafG3MhKDVbiCBcMMF3o5L
Es3dOhSnrp0jVaozoR5Gvdv0ndLVtoM3PxSiqC9mcxcgCyVW3v8tDuvJbuQmvH8fyptnjrqDVXp6
4IdYCei5miUNDYEYa5JrrP0qqjkrGy4xZayZXFKMRX9EaSB2KlSJbFw/bw+rfpdytarQIcscqBdT
3fd2iMQmgBBI0j2lmK+/JHNDca2qxRyv0m/Ex1TaPKRY6LKH7RqQZrNif6P7MZfKEKC4Jd9IaFCm
JfWeofcTnbqcIQjgkixujN+nwhKbgC3y5tj52tszg5JOZGHm9SSm/kJw0OjRhVSw41zGRecB+KsF
xLhDhLQEiOhExjFBXE7lQfUAO1TZBZ9Bfp/dFOM8AXAhUQ7437k0pVVsnWpegRX4C+3g4vFBKigo
56CiqYc/QJDgTXpO5D3ASIvtQBJloqVnGNI8nC9gQ/K8+mRsqtfZ/oytPe4f5moj93lRE4VlXm8w
sJUk9FXJ3mvOyn/ph/U0xiQ4CEMei9QUbHtpga9TSHBeXxzKaedtBLMxRvDml/e+q80MiLRfQVXQ
1vxzzAVkvvGglu5F3fo5HsyHpBvDVpyHcJ0/+J8RM9PRhKCCG4zI8WqN2BQN+jfW3WgvdxM4L7ca
3C7YMJevcO/uqLy+vQIPGg1qjFw5/cnNBSGA1o1GtM5UgJrB843N7nbwetF93mM8l2VvwhhnLV9P
dwBslz+qPeF2fbJWvEJDUAz+YGezlUKYLsJ+73E5Itqc78nAhgsQC7u5NIL82CUNDsek4OSw1gIM
AD0TrKo3FvKRk5umWYkKtsg1+Zs2mEaJu5lrDnSf1tLfklJeVf2YtUJaY3T5VebD/zR332UobOOa
aB+1qyngSOvvq2ybphQVAerfywzBuhwRojrag2MOx5yXhGvqna5mfbeK1I6ecSASnwe5AvDsdKAB
UsvgjRhgiC1SQfJoPLk8ywgn2peBb/Lf90rK7bGt99l/GBNxWWjOn1q+6Yk7naHs6wz0675g90la
Gnjc1RpIRCmYRvFChDAGRFHyWA1c4r9p0M6CaPUOCwSdkvoIqjEzZag8s72o7/1SDVb/C+lgKRlH
UU5PpcmlJ6+JqVYjSdlqnbaJjXRHkaeqUHGokt82FweO9y8XqKa45UcVSLLxRD+HcBDIgisagoat
FnTvoYWtVh2WkFBLbkWowfOFwBvOaALSmUkBFLAeR62fIIeDgxmo04ILwBZetDjeuJ11yZB3CLKT
9cKOCOtaRVTxf5uiRx9YVul7ejHohHQcgdr+If68ku4/lenfusqTwsQ37RVSDEABfVdOu/7A/RZA
WAMzMyqC748tJO19A8ln3VALrOSVdvEniNTIDjAsv5pLWT605XsKeIRw+36s0V3w4A5frgHjQ8nX
jlNW+ocgi4U6Uj52Ugsj6SDZePj4DXUecedXiqsJLdmG7gLfWu2gSs/XgZXTjKoQJPTrRY4ilFPo
7iFuoAtWFcXlMqLrdsjBq5ybF2aFwxmK7pnsMNmipLhwPR25MX0Siqq94QJVgDomEiAS9a21OguN
wZKi+UG8BkdaIxaHTEHtokMTdU5Qgm8QCB+eEtBwHF2Gj4COJeMnHdRQ++ZlzZHOehJiWY1t5fox
0jUXDxKQwmG9iebsAQoDFeFYzY+los2eJaO1lxaxMja/puR9TDOhhLwFvVO52e4onodmDWBzYOil
jbjJ72sCqsWZQcrlonfcoDsq8/8ToAYbjcQAeYEu4bX/LntxWmsBbaqKDryWTIEa1l3jJaAEcH8M
t8fNCx3LWBlue6crsxmAF6eXHpWrYy5gU0nYJE/PmJNBJq2UhdtZuvSk6cLDuGTiK20LZhE/JgT0
csm8cV+nA/CjLpxws1KC5KACn0zCCuNHPi4m1XKIfkTgEYS4E72QTYm2twAZmLW3A1b2UwVRg67K
Lff93XXOcLqTH6v2WBSQnrhryCveSGReuOkl4xQAIHaZiNjQUlSR1iP0qt0nlw9oaxzb5fk0JeeG
srC27963q6VX5BF3cWcuKhZVkdYWXZaDkPBbiGSRseA+gbncdLjuVLIvefGjRNCF0dt4Eb6ff1Cb
mGv0uIOvDP0/A20axScZ+50E54QVXHoEZhoHFX+WnkkRAjOcr/yK46tOG/DBh4zU7QjwQLTAjRe6
xcS3hR0EvZos32x2lS3WctBbWnpWxkj9fNVmrXyWtwM12kYgcfwWYo11XGHXQG2oziRp0CltCROO
ArEfzyVkq62s4G9qrC8izvbAkadr53RF2PcBPVCFITNj/kdM5apanXr6H4BWaTf1TXtIlHU4pBEb
abmwLwnNNGlKND40wtCBl6MzP8SwJFOPZplrDmBLqqJkx1qhrs/EM/JFQmIQHiluLVLNKyuS2Dsp
Ep/6RAgEI9dtaeV9AouSTz8IY9KG6RZB/Oz04vJyl3yWqCgAZbcguAINRDrPkEhWi/QyAHFyp6UC
Yw+kmoEkddBhb1InbYT9A7Mlt+3uMgSA0vmbGGUp9HvTEXWEJzFMK2IdRI95j5i0SQtDjsUpW2xk
GCEkJmNKptvCWuFtoDjQFzoSylyjfzWPV0igps/NXr18atwvXRelM892Or/X+5xnjImqvJnwI1DF
e9VUQG4Tl7kfppxTe4SJTaDWuFJgbIDmB6SCgkha6vI9gyCu7ZxWowjc2M+pgk2EJLDCrTOca8Sq
Yy2pKXaUgtLmDg5v9RN5gLAvCpr3XmvEYS6nhUh66YFH+BvnpZcGYheMhdPxiBtlA2PiqOIjLvD5
TKawiWQC/30C+b5ixdslum7r2XnP439mIiQlXX1R+HJ/ItVwTJYi3ij5/KgU4txhS/0nNAzVNhGe
lIQOP16dymr7x9CUue/OoMErOhum+/NNY4ml5hpb8Epq5wimYLDN2+jKkDeBSQ01UlGWi/77nfr4
BotxLviIwdIVfZIqD75M3mFYdunTkbT8/el0c2QHXqPIiNMbfKK65+T4gddyP+ga2QJYAg2A6U2h
KKZEZmf9qcvQQD89cBRMYEXGV56kcg0q8yT/y2gGpYjGHZCmG9oJrrZabyIJryZFGyGruWB1N4w+
Y0iOQR8gH5g+0Gc4Zx+AFo2m/T+InpwnYgtWtvyH+yG1WyiSTX5sBbgGlq3oq9wMoxKiZjW6qU8I
S/MqlK4oHuwzso+yiJPnSRNtERGvccWSNiUu4pPYQbdt9KQ2eRAUed6COLQ8YPbvhVCht3bz8i3H
vCx3Z9d0srYxLS6/doVgLNoXLleLafxPS/hPNlCHhqWP/JpTCZSwzlN5obC5GXJM8NzeN6se6qb9
q7ZS9jAYs7BJD2Ijdm83VoKz7b+nEVQ248ks/yG64uj4vFmYh/wfaHCJPpqCBGQHR5QEBQePRV/0
FH7OMjSkad3ZWVmTdOWQBwAJAGxJPDMWRdUFUQFNvDl7On5nC9q7PvCXi51g1SV/Oul7NjxRZSuo
ZApz2LgJwLaLsdp3x6/y3clZDZVody/RCw6SDEZN6bPWonLfkxjFLNRjOe9Xj82RS71dQ3pW9UN1
JGMGVMSlRquZozcORyzA7U8fSuHQ+/g4lg91Q8VLm0p9u57qaeN1hLwsnil5CGqwBCCPGBcWMBql
MInY4H6yoO6j3xoQZXQ+M0PKcZqE8NQQPcHF1sJGC0/QScFX0zH8xOGf+LBo74APEDxE5HfEHHDE
DTCc5Mej+8cMGS/A6jm2QcNxu0WYeZ9P7AKzA4MZptRigYJ3dxXp1+9I03j9BMNs+WF/BKTrJxvu
UtEHFWQnzK2iK+gqT4OIC4ZfeUpeCOFsbxtdy6sjGI2Cl4tLTdG8XksXX9jZP7aTSjzY4Q1y3aC7
yqZwlbAR6iOQ6tiK6+7GhKKvaK1eDr2jrNZxiJZY/xr4Oyf8YpXHdO1F51QiaY4gnYZX8Z0Temhf
08mBYDMx12BTiM2CucyVmVkcobIEhLDlvxxV50agkP2bRvVQ5faXNteKKzzHUvtqXgcVFvu1qFiF
xenjuJCvNPJ4I4vVMCWYllK2biqjWYLiA5GD5Zy5xu8MttCudgyEL0ln7D3JyRMT33BGindiZP8l
5NHkfOjyW+p/Mlum/gPckewjq3S+V6614d2oLlQ6vBLMXzNXREXM66TEugK5kbuGaNHvDnXnR9wy
eccGk+JPBYBlvdThHDs86GVQVJFwVppUxKf1TELgxFmeBPH9Fblti2ontZlmWmoV/o6DgPEB9yYp
hMlHUqlw6X6TWrtYgxvcrNWj69XVMP/b4t22uzQsXtD9JeQPEPsJ/0Vgl29xvdPQk64DQqfbrgPD
GI/3OxE+zCFiyQXoOoXkKRJabmnpxITWZuqtDjk2V7CSdhZLHesalxH18OPmNHOVDU6EkBxB2h1f
q26e83ykofWmjvFLSsAgIKJIXSxJbmAX4iRIibFdWPZDLgoovnr3jMd/PcJiI/9adjRNobznLuQG
/984WvLo1dlemHRnLe3hJAxFb+UPSEiYELWekgxrbFAngGrnImXd5vm+EaK5jGperZa2ASftcHvk
qIW4kHD+06+BLGUR26NrasAsPKnbiHMftLDCQrTzyh4kFfTAbOWG8j5sVMLd49isWtYA0lpR40YY
pD5TKSG17FIIZ7EU6hruCC4OIR+d0opaxmaLD44UoP4e51NPplEMi/Jd1pjahZkInfALSoztOq+l
yKgW3g2/NJj5D+SK2kprmy6WDgPCyJYrfhmBkbfk/1thGZlD6Z/YI+urA3Bo+zcCeVFhYUkMkfIk
135yR5bjAE4PBF303ygJ7tWTyFKtuxmtCOiFsQhG3DnbRYW1ScrudIIz0CGp1lpHOdfGpLHhzJqm
NjP6Tbg+3MeEwDeTmzydFhV8mLB2GlUH0ezr8ym+PeLMxmv/cmKBUFsEu3CnFoSH4gEtLYsnQY0c
s4/FLqA1e/M7mmfnzZiu/s8f1CYzLOSNg0MmFs6DSMxZ1IfIBhPCqDpH4Kc+mhFctaHDkK7sEfua
8xFjulrJZrwX2mCmkb7E7z734KOueeZqpDCkX7j353zGZGcLi145zHC5WKbAcALNzuMEX2iHiXgN
zi0puZ980YEja3TTIjj2KCKd+3UUFNpSD8uVbYEJRRHWsJ1IqNymzA4JX+2wDcVrxxdRFP2U8SNe
mjPvPf9kfXflIPO3ZSJ8hYc+RKhjbmGJtenhMOCnEbStf7eRdH/myYHVCM7p+OBiN9eFMssiWaQX
DasOnDc6t3PGq7EoXyaCYI2fA3s6BlFjE4A1OiaqOuAFr2z131e920QJXHMyAOKltHn1qGC0vpyr
BV34qqvaNfjt4MXFCYDLV80UUbW0VW9vn1o5rlPpLgXFHTDXXQCBf7ZWLRu/EpzhY9pEg3L+knBs
OxlJV2qcXeH3WfFby9RPEPmdtMVfqgmCJzB/2OK4stJdH25NZTRdkkTp/+jZzf/YBfDxqphegM12
jRzXvucUUS7b0j0SBYTUAscnH3p4Lsxz6GoeWEGTfzF1WiflzbBUg1DLotYM2dNKwO7l8t8dfBkj
tGlalf7jQnr/63FPpLVe9334e1g6v8J+A2zWDVSePPIQQIEM6vri1fVqGs3i5iM2HzpJ/iCYwt9h
I/08GPqGuSR6nJ9z4S9Y6OOYkVzj5bu7O0OPd7twmLPtgOkYcAHUROaKlfIkXmyXkkpifNGFMzPR
kznqnFmHqvR9AVpNMoiB4yogWisO66Mp41pr86x+RI0fwznnSRgG3dQPZqYV280x3KRcOrWqCJRP
Hx6d5T3VFIM1kU+o70Xq2Pn6pKyD3qiOh6e78mKbCFdWYQODJ8OSVkshLShmX6mEKfezb8N4VDHW
YmUx5vdVLGFMeszLivFYT/zi5z5DEfJZbhhpC8X38AN0V3uYi2En/Q1N1+DQqdm7JmqpIkr5s5iv
31MethUqPgk+D3gobBUyQXs4G7ZumYJsubnA5Ek8FRlwLwJfUQ7lLeSdEK66s8osNF6foyrEUw9s
Qv7fJAnqYq1f0zbYp22aERixjHkOLeD0AbeU/2AzNKYqD/oRD0N41VUigd9Kn8xVnO4ed2nYzOfV
oVdDot0Om3M912+CnLirtbbHHNGirzvhniapQvWVzdBFvJNl7nsYHK9RwReuIe4f3ZOm63DlfSFh
kzKptU2yG0yiOZg2qfk6D4upRwwxDjfbQptJq1NrgCWERgNJzYc+XQ1jgmWsaULJr81LN94ar3sf
OvFufQgLwN8eFX1ig3cyZiqb7Mg6PM3rldnbIHEhZg+l2D/v3tty2OEVFvoowBfjXJ5zKQi8bFV8
gTdy7Cz/u2dkLgb9lJ91JEaY/w1uChaUUxSXfwqR0zYiOTZm7JHLWUjxIe/gSwmxfSYCl423Bemy
TpecRxzs721phM9/1kyDoFq4kfLuUiINchOF+pl9dHuMQSwSxeEn4g6Nou4FCExbxESqR0QbbI99
KIRQuZyhVXnCEGuwwXtG55nUP0pKOXXYstV5PzU2x0hn/VBoorq1tgDnqtqk6y0T9TpDBrdPZtag
Oc9Hc3EzY8ZJSXPXFKGuQEN4ZLFOY2iuvZfEVIqHRbocKP6ToItq3QWTZySNUHsC3o/iVRJk4EzE
INZnt2LykdrkfK738rxmbGkxpUc/mUaVATEDGA4kWb4BsPzz3hzrq0IxwQ/EEPb3qYRqm1dtehXz
/ta0xGO2BR1D+IqMLiB6ZSk4J/YOaS8xtvl8/0cI3TFTFzFzjjex4MQrQzPcC5htozF6CGhTAMLz
Umr0NVa1Gph2/S3b5eAz5frGJY11o54ZqqDDjedOdmu8QkOoE+zo0kHG04hzHMvRlRvomdp2943g
eJoZk4jS+SRhItmRXKodUPHZqurNOt36TpnCnswOwRCFNXe6NNxozE+uIRfKx9kzFgM+0HpxK6lz
kJGQIt3Wav1Pfz+Zqs4GhikcWp+VLkIg9K6DO+cf6ziHiqf03H00t18chE15Uwn3Ly9D73qq90PV
VtgAPb3h9wCps7vdpUoRgk4n7dGoToFZfa6Ed3hF9w7dbykp59iNvd2/cuEkLFAD495GWp0MpCOj
ZJS57/0KiW2l1pC8ECqaMN/atz8e+ooQVznDxP912Fj9kG/I7Fdl91EBWrgFbSGQ29WWHSayhd8O
1otnWjize+VARDB2TQ2HrjKuKJ4qXN9BW50jr8pHh2geKMkCQgMoLUQxULLFmFbPeSrZKg19vgbO
DPQ7+n2Wbix+onffKXhwe2dWaFkZGmLT0bfF6yPA0y4OK7DVYz10Ma8U16rox/TP3S4L697McDFd
BpjsQgn7gHQTabJ19Xbb/KDmQqPbJGRS9BvnOaijCmi6skQLWCeWWFBkXOob4u4Ai0GUcStOUu9b
2XE2E5/Kivz8le+QjBZ/G637qxxzaKt5r/xHkFkjrtXW0dxjyFUH31VtDVmByKDcbMnw4AWvBr7k
0BbRC23y3yjxMyqe2Cdp5o2pCsYGvXBswpuNde63sWPskqupUcU9QRL35zUADuXO0xoR+sxVMmIf
tTwasufRYudcWANNNKpRhqpNuMaivg7GeryEfFIGfY7WGVLmhzXJwCpSVAqOboutFTiPLyiwuuE7
aS75oZqap2F1mUh5u4jDf6YuNNUnF2Qm38MWnY3TncXkfInZxO0ErnsWBb4xFp/xNdPG3mwfGFDF
R7oC/iiyr7RX4lXn9+usz+xEqAh6uoXMcUnAU+CpYUK6UuNIkZcw6oqS3NQmi28gS4No5/G7CkrX
0rrTKe1fBm7Ukpefow4G65wBrndW+lX1XtwDd+AaQrTzr+KEDQRPPSF5crji8dNf/x9lBrOuavYc
ed0ciQ7R9GRK3oq62MoiI2HCjrpWHqGdzixBbkO8mCTu3tI+MbVo4kLvkBSIaH/ZDB51/m7dnyis
TyIKoZFIpKu7AoHdpOZoK4VLklzQaF1cBdMaZ+q0lctw5Y2HXSltG087bU0nDi1nAekPl9IVXD9V
zwtCERBypvKjtZ69eAcpxiY/xfs8HPLyUbtvi4aTbUIQfeWg6OkSYQ3AGYh8Job8+Kr6zhWcWt48
XzQnIMhvFexv/i62CK7+OD8FMxTAF7TfhP7O+Xx4fGjTl5eiI9POyQVBYbuhVSj4O4iEMgR+zHDK
N46mxBSd96oQvuWCaHj+71DmytRr1fKebiChcHSyHXZMTixaRRnGbGzKjxYCUHjIQJQwGDcRnUP0
ipZDG5X9ux1c2+sWVnpXLCgqI/mMMNK5WzZdHqJebfi+YMTULH4AadS4Utw2I2l79lnGsQR2B2D2
7sMi3NwXMIaUU1xxZox3VeVOIrX9yOQxvfh0B5UfXyQcSwWuMGd34hHiS40+2BkUf7pjStJ9Fp8v
zhzQcBudmxAdesgEIYTJbrLyEv8laAynVpbH+oeVUv/Y47MW7ytsDH4gVOMt+KVKZLaN8f78jOGu
fXILowD/P5c0UuLKjRYcFC8yVsEea/mV1ZpJ+92iEPzIgUc91aqNVdzHf5SgICGoQdRHUnG13Ak6
fyufkVvJP5g6H2mSzFPdkDJNxruhZbNa4bBCF9xvK5oQ0cIP1f08wj9wHdHl/2C8ukWGUk8iVxxu
aJskg4KS166aJSp64gAA1UBjjXPS3W8H42hyJJpfNyR5TyjYdhVO8pkbngVNlD4RFXNhqMH0iyvd
WBwlXbSqDeEegSv+pZ4Ge3z3YbkIKBawdA8wCGyDQpYUkMZos3WZs3INA76a+R5hxEUGC1uQGC1Y
Os9YQQBRIqOp2RINT6NqsHIM/Bk9tb8O4HGa6duPHhTgDvVmuDYEcpw03AxGEk9ZUeCBeQjTg8UM
7aC7Wqa78pZv6guAY6We9eHgV6atbTdWzMSKozJrC/2XyczhHlvTEjGe9FQnG4GYPWdOsp6IHvsw
5qTRLjKNJKGM7BqRLSRR8D8zzLXwGO0JD/v8A21scCHzbp6bnKWTL1em3oC9UKU/I18jh3MfRABR
JY+ecdV7sljTYZ7Bf11TDBu4ooA6bPkAdKSSkd5/5bb5wHu4KGj5mD7s9ng0wII4fhP23XNtaeRA
GPwC22nD8WwJBDxYWjWvoFB82dvbs4Nf/JqioVZSX7j0lwRFfHIpHsj1UPGJSOutE89VoX/9OTFq
Ps83MQGRYH4IXQ07mvJLBcb6S4RoylAUBeDaC2WBbsyEHJWnMOgAlEWvLm2gm2992NxVlyYzjJNA
R+W8wcjtABvG9i5FbaqDJnZAc8GQVeYIJ4wcf/qwC7XuIfzYIORORv0YScKh6YqTY/G+7l1LYoNr
ZW2H0OAr8B+JStPedDMHi/VNTe7lDZJY6u4F27oNwygfB+gGjmf7pJf/YncB950aVNRiaQpUgH6M
0qnlXdLishdtzbcEIgn3exgZ9Am19jACb7IScIX4mOY2unyaWpKEwm7yhUJyNYFL3i+TeeNFd8dV
bExgr0EwN+0nOGXWtHcCGvO+RU1UDobh6ljegCh3nPIkwsphDHIjFL1wmEUAnrgwSoYrtrn6DIDx
AANYQAFBVt0lTHpz94UU0wZnbtyIlL3r+V25k8YEGJtok6kcLgigJbprR8ZgpS0iCJUlp8oXEgC2
lUzoFPQE2X34D5ZA/0sa4+LIc8mrVCXrtuoeEbO1IjH/mGI0WKm4MsRmLv0/exJ04rwqfyYJDU3I
Xly25QSJujTRaRhR5uRruFjofRNADBpIEDRn/vm+kjqztTAaQt9RGvY0j6tH+62LdTBVPX/z/6f1
8cgV46CpF17snmZWkJcdW2NA0H/F5rCmNhlNzmAg3CWtErZmf4IRwT1fH5gJXAgSuhzG0uy/5dU1
tSM1haeAytM+OzZqKaFgBRURtQXIiBcF49XM5smPxBWXPxY5n6V892JswayArE61XiU+W450BxhV
h/pnMZ/o1JYRnmAsPGjoTHxhppC0bzlcl2oiUiMJwQrfplnnaYgiAhFNXXE3boHn07eieWZ4pkJS
beRaGkyrHx0jir/zWrpTKl95aIUiOj8yvHo0oj1iiu5zW6TZgjco+8MKb7hhXX58k5LJ1nVdeFBt
SueXdelTOwNDgkkpX+QCCMTmn7MLZOXLhjOzvcW8KnNzJEbBKN7F18GeQeFVdUV51YkN3Dot3bvB
GT9T7Iqka+I8Np4+ukUHtiFGKOkO1fGKkydlOwgnFgZ5CeHsfUVhF/S5DvxWiYEyeYKZeyytfSuA
v0XT1qo9a+kkOcWUMv7ZcPnzlw67dyvERkRxfwM9jpD+Jq/0selMSvqA0avVVdGF9Ck3Hc0PqWax
PUQvPH1KxdPGkmFEboAPck5bICnaqBvQL/+i/dipnWYrt4jDgypCj7UO740SWLCWQ/YnwkPHs1+y
bfAw0O9YRZLWlM2Ei65swrEqdMkjqG4W0PeTnAGjDUreCBn11K1NcIBJEt9dxXAvN8Jx75sl5ioM
+g9AovqcvZPUzIe+8MYV5t4dN3xtLSB+EQkZZ0ISRK8vnQgXSLcX/XL11kThioa9ay7marNmL6yD
pRUKiD1u9b5yJH56nJlq9Gm8uP3X2aZhUjm9S9VHzttxl+d7+DCIRmfJXIXJRm+CcA+V5XWFCPeC
NBTBvnzHzFrHABPgmIn+EhO4ni7wKf2+Bya0uXzwhmFX7LqhydIHhTVmnTIPDCkHhTB3mYqjrReM
P6/xfsfthQN5m7zJyN45v6ek3/UsP0shUWJ0ArFBLzGl4FfZbRRHr0Ips8pU+KgVDLGkV8qLJy8T
ausODJuUcXRZN1qBB4AKQ0dTm2QnvRCFSwnpR1tcYECwff5PQFCUhdLjDffTCbe8mWW1Cjy0I0Um
wGuVhq9T4gSIxUBwxotnjLLUlVL7ga68TyeHVE4/blv0rsvfiyc/4vFX7B8Ko0GqTeLyh7J7C3m7
QoG6tub0Fa1DCOM1DG9dwSLtFYzvbi2z/nLVaKOEMSyEpMZ9RAO5sA00hQWUssYLJcn6c9psC5ZC
rAMaa5G0Xtif3MrsnISwJ+dc1MbTD0QQiF7uj3Pm8OOi4unfQB37dGxIagHQKzJhCBlirWLyDRTN
jNlfQ8o/9n58cYADf2bB/aIDqugOlVne2J8BRCKgFagLxTsTQXgdmFSALa6BTEU71D1I1r9gwx1d
HDqYgkR78DxJM2Li4WxMHCDbabqY2IsAy3vEB1k4BlMWQIJ4OZWlGqha3eFKR/FtifZoLLc2rFaz
7zjcLHdRWtciN1GHf5zSzgEbuk2Ss5Py+XDEHAXtnO/+84kh/AOETd2vEj6mOmxnw/fm8RtTag/B
ta39moBhkTNNQ7LCrIiciIdlaDt9DxE6Vpxfikn06dQwc4dzLD6DMBL3EakP17FDRMoBWX/qLAvQ
EjqKng/3C5vgbkJXCpVSOUkMmcMeqFtM1SZwE6j1WzkJh4DDtR14FDavKsWObWB6f0ygjZvkBzBu
lh5zxiSqQZdLZX4yEQrVAwgGnvN2OA6O+YJfb3VQB3fa0lLuUcYZvCx896/Yv6qA9aO3gy4YMPSI
8e6cmyahfa7NDvRlpZlVZlMFxs9Sta+dHjfe5134++dTQPUunddHJsRD1MGnNOeYDenqRCzg00U0
N+4EiWPpDUd2HxhlAxC7ZbIeuaFWur12aI/dn6FiQmZegMmf6i/yLNPBzCX9c8ZGU9xBMw8ZTwvz
GmSYC2emhygPD5dpaBAcWj4pYWtP1eLUE3Gb0Y+fBScxb5FLcvctltrzOJJfmHg375bBIQjiJTXI
2ffvLWj81D2YctCMEkx62huxeS6Pn1msXr0vmbfxUd/xOPtQrdlTyxBfTcnCOmtE0nI/QGZCC0L3
PPi1UQftGE0G1GYMbCjzfTDhgUIfjMWd2zvT4pS9Y+D8ikD02OIqIzF3awNfJM/ozgYlZTUgsj+T
I1QX9+8wFrBb9ZFmdphNcI+QVPG+9qisPLXZrtnqqxhWd0EB1bC5WkfRpnCH4L6/1b7FCZcJmnJB
5vPBV+4UJ9a5aN0AfCP0HcMwj0GUWESZRTb25DaXeOZzviHVXnx6rR7mHwa6A4NxyMZLy1+Ahz3b
oj1SLTgfHGNy5WYiSctOd0LtSplqY45jjTjVWSpm8jkYPhQk4RqLSxKAMShnjxJtDtLT8T8uxYOI
ot1bS4Y5wnXHSOBOP0nj08y11LqFtgD0wZT/mt5cOsqsyJiJKgXsZ6Q+8UKvQp8wxHeYCpGSQEOv
aVzZUYcN8CScCEQvMZ/CO7MjsWHNnp7yHjdx1omUk+Fnv1sC0Wkt0ROPPU0eaG3Cv//fJ0RtKlZz
cs3j0+rplNvX4JP0HT0RF6CkCKTqHQcz4GYceCcy+42Y9wlKcVWQjmKhUF0mLShXn4H+i9gtbhGR
BO3dbi1+l/nx6XNL0PqfyMnMys7psuBr86/k1QQX1cwO7RS36R6pCq6N8FTbqsHxGfumai/e65T3
9xqCkILIFcDSC9y0mXS1mxLNcx8wwLo3L7G0eai0ir4/o8835aHckDx/bsrs+83LlXHmWwWvujxe
rxX5Fo9JS5wNRyEevlU+70O3frxxdXFqe4QzobK+d7nSKHcAImqOqktrHXN84r6fLSOPePSeDxXc
0fw+qWZ+j18DP69hlOyBFL9ynxm8x7wwxniNDFYki3XN2UMLR8On9sSsfx5sQ+AUnEkKy+t297dk
diuQYGmmeeo8Ug972KMMBy4LxKOWoMKg67Cncq9wO3nWTZkd9DUfCtsubnGTXyHLzI83PZ9UUniv
HcZp4JFEdMjMx+2/FpD9tcO7pVR1NOMznXQ89bTmhPu2sg+5PCwDfxHDHZVVpOJWb/ExY0mihg+o
oq3KpCl8KX9RN7OObhHn9diqG5hxCRcD5GX6ccdDpaj4fOaty9pEynuUsIG1oOtquMO3rr5bdpl2
ItrK7abgSLgi4JKWubwqKlC+P3NF3UEskq2v0QB5zBVqxKr2ZLHdi8JBcFeQYNME21TaPz5OMbOS
AcVlLds0SI/rTWJYYo2nRVwj3vFUzmjFhXqKPTrBqJ4w51h+mx/SdFUQHbga5kA+SxyOh76HrSTg
mnNKdV4xWnNkYJS/GTlzoz4kf24TEUxMQfGa2xi5gFUYtTxBfns9N5whrSCg116NhlFzLbnVzGHT
bjdXfF5aoaFdCAoO7fVmvusw5Ib0WcK77jf/JnGEoywYHNMCq/85OCyk3dyMOMLePcZBkxBvFTdX
3v7GypD1sny96I7QXXAkrObWhkiGqJizDGMx4bGQY3KiruiuNPZTJuWxOTUswOT3xykJAHC5PvgV
cr3+Wn+QPMIPNrTZ9DcXCKvmEKiE2eWImeOJcfO6N4celd0eTFzIvE9atMssmF+5u3FIXOS2u5/p
xcO8dH7lsK03M2Le6rW93ewJgTmenj8iwx6FhGxK+aaCIF+O/0zsmxnii9gqscnzsUK7/lJk5LDp
rT45ouXwjtAcnYix2DqcJZ2lN74vbNotfh9n51vp4fkyH9dyHmOkOXS/rquLDJ4fhFAQvdfn7KGX
PZsXOpMET+cw2aQPh/lCQtb8bEuTbFuxbjiEEEpxiAMSF3BgHK+cBCV32VQ2Fw18d4dwHqss/lyD
EWUOBrfq4E5Kf9Gno0JVtfqTWKTvvCCA5Gj155eXGIUlLzWfF0xWJzaeeQf8Wp96GmOKb2oD4nI2
q7ZjHsyTdLKvej+voy3Dagtn6Wype+VwXBznttF07rNF3LNDgqybYz7aAugGHS7eu/UAAH689lYB
N5FyZGG+D7SHFrK+NM9l8Np+Ph2duWYjhEzEvwRM9lBjS5mkTxh5MakHnDo4gwC/oyGtYhc0MtZl
80eTYaSwggqGeN+Ezlk/9CjQ0zjg9z7aJGPC/asPLQTQGjVZm+2NguwlCnwJ8cSjGV8WR+z6Np2W
rXpvCYTZMRfE8w6/fppU1twc1WLAil1sGOciwZN1VNJFYRnpt+IB70R7qyVPERkpoZhXWxwV4jTO
zuHDoOrRh4h0+tHDorZbZ2UAbaAcc3Bx5/bHeGNmsy19eMmzslCiwzZ+2qvAmSZmoagSmmOmmmM2
eukXbJV1SLaCrfsW6GEb13ORWmD5dazAdlqGemNQdUsNkXxZmGFfUgfYB6ceRP4d2xn+meC1JC1K
zkoJBFjVlK+cpLJDqTw1H/w1tI0yWuKhTQo+fPHiyC7xjTU4akkBEO+6iZedApYNnNN5l9+NtVAP
/WGzbESrGBv6YeX91GiDcT+99uCKUQbfHdSBOB8EwoEtB9+UBLPqLt3hQ5ehW7IeNr2WmYhgEeCR
TY7p5sWWM+ICx9PHtWtZtwJKOMO6NgcCurkxpfCXG3tznu6so1W2vQ7KOUwX8xttMMZce3c7x2WU
3OwCK0bkLaVcgQ6qoARpkCKC76pX0o5KaTHgtgp5tVFO+8eYCFmwPdIfUG5Cfu7kISolbcgOF9K5
A/bCwiUfURv2CyRD3GCc7a+h+/XerA6K7J3vMLcxilVPCTi3tTfty8lMoPh5p0EG2m9F1MoNGqpU
AXAgjv081m+cdjlD01XRd+d3cpj6uBAnTLxR0mal/RycZHCAmrmL6AG3n7CDGOr1D8yWuqWUhStT
IqYJivR9fNRDzaePto/AngW6ysXDG8cPB8XxRa0ALydfNQcsg2cyyxHRmpqsH0QaBHTCPGxKCIWR
roaq7oHTjlXJj6htgEtTT0wjGVWUDngq8mF6EkNt8YSIPf09lx9dn3Vts4MWuqCBE30SB0VcoWqa
sJntz1pdcWqWAEV417w2TBOKL/3gPt2NqkCAwiSQHTt+Ps6hYpnbnGUNJOhZgjnTBNu4jYcse4Iu
vDWVkxzJy3jhPXUXAvxkB65J1KOZbdg1sdMT98xafvtY3+8ocSfbybjkgAyMCwFv1FmgEeqd0aW4
Ni+xzAZ7NuC/p5WSr/CW/8R5zwhUsJg8IV/NmnBOGH/d45XKOfbEnWtHl8N6Fql3Lof1F+CsUdt8
+BqEul4WyDoHIZtw7Y3F4mNTCSK3GRt+U/UaSckACzXWOYKxOBRhDyoYQeFulrHSz+Bsd07gHuL5
zzGNbjnRR1oTnoUS5tAGPpxhqueHaZ459c4cOrNCuMau8dA0x+oY09SSuMdvOCYqgjtJcbPCI9kE
0cB6Cmb13IScvBVpgupo1aq7809dNPBRLp0stsjXqqeaxl8YLYhRhsO4ESJiXaAZsigxpfycX+K3
5xN/frzEEEPWREn9uXSlhlJ0k2/qRgkdpej86s1Y/zcqymS8lFhS45EGiie0deCLt0I/ASuRs+BD
e9Hyjbb+zeyv/akWurfUvdjTmoEmi5azi792g1xVzQkRPXF9e8RpsMW/5+d1ddC5S5KkmyGP9549
RzNWKsT1RbOAGPpmPWW1qntfWN9Vo54cda1/CtA9ZnRmkrpubFj8MgAxMNZQ4KF75PMzJgEHZtNR
VJzNuAKPu1eUTQqUnAutrLE55iNlJ/92aZZVMXNRK8UxRFafLJYybmmY2jrNi9sUyBXEuOO9jeGJ
Oj7P55m6RdiEMS2h8s0P7AJySfy+bfcwN4140cj6RbP0xAKWMzVfayvgdd17b1pGL603XaEZKqEw
lGKPxncDyvmew+vjxbRIqXKj51wIWXCUUuWylho4ehLKHBP9RjMYQ3RV8s0ocG3WZFufvXV2kNsR
ezaKuU/a/h7TzVEo/zVRkOp82+ML2GSyFItKMMSOms1MnbHG1F06ekh7Avz6dX39uYwjIhszMZQr
YXhh4gedLhwiAvAxkycDWJHNK8nlla4dyN/uShgrMia3DgEJgC2BOjyT0y89SKNhvGEF3TgoMCqb
xVMkRu9jRFi03OMhSLv+PH5lNfaT6Ld9kEGq6oWwmvGuy9yKC8n9Hq0u4oywIn3BW59AECVrF+5v
fqotLoLk8Vrpr7Wd3DOpDtfSG4UTO4MfxhUlpODSfkrJHNJte7Uszw/Ik4OUC4JxIJtBWVZqGX2Z
NE74do/yJoaWLOFtcaQQfgpNrjqPpnXbS8KnSrfBptiJ5LAG/fXbqQi2I8N3tkoDLnm13jVKWlL0
lRSP+xpy1dMg+PYSg4NMFDrgxAiHW+MXFsm3w3IiQeBa+wHfzj6k4Ti/BVNfCLOkHAREsIetedgw
JowcU/D4VLGfXcOseiO3W4tuReD6sMp0sKSxwdWANav/Ftm5LlayEs8/4K53YYCfFbdYg9TPGWLF
JW2ACujuCtWTsK5Ap/41+SLsdisW/6vkD4PRdiiKuaFKoy6pVzUccw7iDnMiEwFoAVFKcTv+55FG
hTFmVAYlYULaoJpaz3mEQJp3QDUpSYfoQppgjb/+nv8u27lt+0uRcLCwQ14h2Wxo4p4YV6Zsq1wA
thlcAAVwP1rVNXAje97uoBd6H9U4Er01tPgpBQP3jjDk0Kan/nmbKCSttaunRRumQz1KxXoGm7gK
8Ipe/I/yk6vPJu/7Tkh4GNcjeAiO2Y6QnQrxNJMD/Fr5H/iNvT7f0pH0lof0HQBgrED4ENMyt6vy
VYZQUZaRKiNgVXo6IX1fI4VqunkR5LbELlNZQX33V9bNwCE7KH2MdoC1atjSjM1jF36eW/k/+3XZ
AGYNLqRLPBcYvFUz4trnRFJ2itXfWWb4qjC52YlnvyNvwvWoggBhERExTTDbFzLPKF4u2XNCj9So
jLBnIsP5m+kZcoUQBUPrGDQNFcqMv1UK8HBpz8gJaKOxFLu4FQxqW9wvLHcn5uyKpDIQt46wrv2T
Oaz9EeepEq73vXoS5dhyScYcoNSefThMPZaSKFR20b6g5W+vjwjLygBD/yP41YDEtfxLfL1RTyJm
bGCUk/vjC44WUxCQs0MiDNpCG2UyP8z9lNGaVEb4uJOBh9AgLAKswZxzhyIL0N84L8Pe1C5a3yoM
Kx1+10tmVytKKUGuDiSdS9VEl7z4xCOyi3aTq17uOdB3bXVIusIZEJ3zcnGTcwtvwCgw8vvRQom+
fPZOBFEyavDSbJrl+gckr6dASXKhKb5Jjg3Y7OiVG9jJAlF31/O3/ect9jtwH2BfIvTCmbQ8eeDz
X4NMpmVA0od2BNx3dsQ8Ubr91fnFhLMbAhUp3/PQzHcZ4m3VlisY+v+4ue3AQskzbsnHbtojl/5N
HxUGK1kfYRam15zokN81ctX4DzjcwrcN8EaHiOy0UQTqk21Up1NIRubcN+4AVlRtUeKlKfWFqlH7
iliMaRv0gSH/TySQHioWxF5GxzcvuYcy97/112goO8CpP00hmrvcSHI5mHdIVW0x/ZuIdAa5Sso3
ycd+V31uOC7pGQkyAPsY/Xr3xi9nwtVPRkqXHwYIQN74GZiGstoBxzl4ZyVAHD/Kq/B13ofhhTWv
Kooj+jFl+ePRXh4E+6tGU5gRyQw6rbGpw3HqXgs0NzwCeu5yl0ivM5d9Egi1lVpJGH3sVVQwJXgR
pbaWeCNg2ArNZ/eeqFOuT32zgLlD3CMgGtfBeOWHcwULxUyhgZnWhrQvg8P2rONZjR3JHjRPm+pe
d3h+5c5KBDV71KR08EUhbIY5+jepqRD2dv2xDyKiiINyj/qDbaz46MWeEhNxth1mwkBpRJfpKGcB
mMo5+1GCSpTDtCJxcR5FlPr+gXLzT/Wi4x2GfBFoxef9HnW2k5m2roxR118BhxFJid6iisbRWx9n
5I+VG/YVjSyT2RRxjgv6z/eWS1ChANOeGWqGxg2gMbrM8BPsXxsDymVT+hD2kyUO9WwGL0WAScLK
44R+IPytCZB+n9IaBIK04OSZ0fOROgZB2IZShT0ZSUw9FrbbwNdo7dm9eIPSzGAcXM5nA5r9qGC3
4SYyvIBxQgvR6EERXNzZIoBADjbq3SBzKWJoMvGfrtA16B1VZejZ9J74JHjsetwaXbDSAiSYpPVd
GlAWqjKcTudt84z9dr2q0TIBkoZpvJbRZLP3IlobESAw787dxVAnccFGUfLqNPfVcO574nleA0UK
9P7eMxXHi7samxDUQ0+X7y2/nVCq+UdI3NGQ2sddZAf5aSQauDa4KNjmEFT/zg/8YOFya1YSGItA
rx8Na940w81GmjBhsB59vfoW2WY/jdeA52jiei9sMAbxuew0vT2U4+CMxOSKK/i2NL14/E4jfXIo
upKXz3PPKXLqV/CwV0NFfsblskiHcjYXSPBCC0j7f8jeqX6QMZolqUv8c3lJ7CmhkGJzKMmwqK0l
c4tvfLVMNLaRNGhGtlk0De691E0S43XLTkpBBpTAtc6iDqVQzQhwbgWWBvAeIr1N85JKadi2K2ag
vVlHFOVKwPcLT6N2ny1Ntts7jRgU1PMGLGjp/pxs+VgyPJ4lbk+HZOQoBV/tkEqfFGWRNZ5+mcdZ
KAOUf2ec7Otvm5L8Qjr1NfoCwYb8QUPnIu38Z1bMOePGvoE29nksIv2be6c7WYtHNwH0FxDEXExU
IkUrQossWj/V+H0nh407aTxOaQliKZ618rIDy19Yauczv/uH0u6+9/1YS1PrPfYrMj0bEvvBj2Vo
UbYXntGx5vaKI57ECrGc0Xe0wiaAkKHRUnCYY68/5RVlz/AN29QTk8kiQAV6geZQtKsP7x9Dj93M
TXf9IyQlxHlwpyy+6xheD3co4uuZUXRKp+Bh5Hz9wwUGp8ynrxVd8Xt4ndOof7apQEztPDJVjfOX
9XHtzIeKGX61dr+STaoYB5oOKDLUfDT3DD0ARO1A3HQmuAAmVGham+wQCizhskNI2X8G0hiOtCN/
0NXVGjyK9BEXT0yVt63VKPXSaCdFRbiqUp78HjtfaJFHDTFcQzuM7DjoPksdCGoHpzBd673f7spn
/9GO+qqsxKdGpFVQB3AmtELKTd6pDLXGguGSKrqcBCQ0AtSWwRdrSV5Qj3h9Um/k3cKBfKjgAw6j
1FFn2XalOOo4oSliVVS4ljPwHl/bwqBlC/lmU+TSv1nX3UutKcFQXiAHQ9sLKhUNQSVV3QFS2Z+m
H9ChEN5PRd/QOfgl1djcgLlRO0Dzn4aRQNxH2fS7OoRuuePtyWv8M3Lt1S1IX0v/sCcecvRFtveQ
JGQjWkBwimZCJxDPSbvt7CMdibAQJW0+M+UZUngYL0lwv1C1vGgpeqhYt5qCt2U7iixnxnhhukrJ
kmvCYA43JNsbjjQb3TnDq5mSqgnlUAB1BQAWAxdKvKzo47swb/pvLOfvtZDFxWa3iAGz2cSmPWHM
jMBEjD/EbRoR00Xf/JakURDlDIhcoA8b+zRxWPUBxDoHet/jt/qPe1glrVxS/Xf+N+vEY+wHM8Rv
282QkV2sp5oQaCm/vbNxvkPQK7f0hplgG31pp5fz6DE4+lKQP0MYBsUUWpHS94M97kXj7ZUu3LzR
w0LzCfDyAGMSu2Bx39SnxiTyt6IutCRmuaC2t6UQEkURTBK2kuTkO7SRUoWzfuZqsw20Afje79gQ
upFcKCOnhKLvR2+AxV3rGYgbYkENoIY4d1MlXA3H5p/omzIxaVg08+VipmQFFu9/Jw7aD1YTqIxD
1akUfumBGV/3lyQvvm8J74mMWyo1oDS3vx283PH3ijpkhDOZys8po1cPM19Qa8iysrNedhdBYB8F
FYRBCvg6dNOrHInF7Z2EiBonTYjEY8EwnnkEE1nnMrgYgSL8ljSJT4PjggJzs0+0WtpYAlxpduoA
U7fhlUx9qNr6kF7rACyccmMo/4CzuZpp1mpKApysbzzJanIaloX7IjUMZkz4UMLlAgEogG4yHtQ2
K6yA8N5mNYzhbiHwkZ4rxptfInMeNjStMaTiDgxfTZk/1UC4QzCk4gCsJGSCSYpHnE8SsquVaC+u
b8qVoygor1b906jgcGNKdeJSu3k0FCPqudenLa3VrHA/YCw2gd9OQ4YUizUtQSI0xi1EAVdeUuj/
NasiigoK/c/rMTXUDfvIy9TcIGxmyc+cSE3VyQ74A86eBtaXxwuObtohxrV9iqetS+swZf8FeFUK
BU7kSKnBEmU0YoBgaNjg8Xs1sDkqTS1/Uu1XBvva9vjvPkSNMS6H/A5K3E63tUTFx+BzRMpy/YXC
d58xnDTJyiUuGK8PNPf4ehyYFho2YDj8T6vj2wJFihWy61ENLmxnmYs8CBT4VuAlyGcB+e9O56qk
4Z9nVGN8UGAc44bJuATBHbQp0I56TqOQSIlJcO1KEqOv5gNMg8qpd/5QDA7A5oTlyIYGoixj8nYZ
9x1nw8/OTW/f0ED/+1ArblRbG7GXcVGZVxIflIeYHPSK+kqmpeSfcc9FwigTq7OfSGXebLKBL5yo
f4nQxov2/T/XLzOip24tSnleiJVq0W2EDSTOtCHbTNJCX2lKOZHrZ2CqKiY2OTi+NTrQWmaPqWth
l5ZYwU0cubViC3X1PqRo4MPv6+zhgt3bbPyGWNTHZnj4FLo0SuIhBcAFsPpdfIZKXAssklVMjsSO
rqC6LNJJZlI8RAZhpVQh2kVbHnUS9k9bJHMiuWlVrixVfYiWPjbVBMiJrD+JGMqk/Bo2ulE8C0i+
H4jeu5lUNL9cjS5g7bQsECsTPlnE0GQ/9bobfvPvYBuruji0ZDZIhwBpua13hcy9CQScfdhJ9mMj
aITpHYFcPBBd/2pPdQVlS4ZoWLvnAZtSrBomqwRutgwfFifLqp5bhjuIYQW13EXLjTobKWuhWSow
L3/K380r1+pbsKAvL/HT2jQRZbemOrc8cKqPtXcGb4xi75W8S/5KT+S5nhuQZx2BIP5BMljjG7my
P8Y+ths7brZ2ZG3vVwsXB/VuSwwTmx6qNksyphgMwsAi/MY6so8PX4DVVbjMlR+/dCCmaGZmksaz
jiP+lSMM2ttgn3AnUMqDPVycayRSWVfhyKtaQeexu9yo81IF5Uyycu3ASVTuEDERcffGfIC7Zwtz
FgxTRUO/BfwHp5k2LVPxoQO4ltNHHGp6wnmnFjPfgegu2Vk8YN1dXtIYBYY86ALbe/BaPNWXlyHm
zEJLYKQs3aTZp60HgeTHQf02kRDXdXgR0FugapIYTEEE26L5K+Jxs27D6j58MXHJqpyQL6lQJQzu
SyOX+lL+KoFTSSCIOQSUjYHfnVST807QqNwaqBwJJNN3xZ6HJydo/5SLxKnxUfjaHc6s28hKE325
FqdC86cF//5RprvjkIFB0nZKiOF5fQlNh5wowiHQ7GKbFcF0/txEE+nyQrVuky37P59CnSZYv+ji
kWvRjDxdF7CGIC+OpZb03y4NGsctOa3VlmWeq7X3Xisqr4Kd0nA2p9/WOZ3RBNJfNCWr0BI+7qFz
2hV317G/HWRQ/pZng3qAJSdj8IY9MDWxFHwTLh3q26rX12iySq+JpoENGsou7v7jyK5+uHQpuFMK
t53l+BR0rvHu9A+EwGhXk0c3EfXYChPzq5q+omSSejFvR24fo98vOBre2Z12nVJyuK9HbIah7QJr
Zt9PZ1QGzIRqPtVOEfn3t5VF+rM2/xXq4Y6nsvWCe9BiVN0rug3lYpQK8Cbg5WNd2BYjxoX2I6G8
uHBefNYalgr4xoSPTiY7X6BqGG4PN3Cms5jcemHeUIuqi9BTJYXho+PNnI5ukV2r/Vi4nwuRXUUR
JcFNVBDrS/vBI3P/vJVCPO0dejI9FQZ8IhNiI09g6zwneoyyPUdMrBix5QPHOYNSAHbzmBAD8lyL
i4JMg/c4GhR49FzcxFk+2fKkEz7rDSD2g7bLnf+g+CTTuh9trzj9yUTDMFcU1P0Si7AZvgJW43H8
6Q4PF39wJRNEheJcPKW7JpnoHLoMrgtpU0Cormpe8Ns65S0eAVB4887FVB7lh1iQrVtVvtVIVRkR
gMsIzkIP9XvdxQvOE+e8zQFx2VVDaoKl8pU26vlE8DbO4qQ+auB69YWXKHLOeiKORSlX/QQu0CfU
nnW0g5mjcsrAVRD2KtqFZrTfz+s7StyWMAhNPivqd81J/1cjzY8o/tkY/PhVvj6O9hTjfz8Ml9d+
8zegMCS6GbfNEFcrBFDNxptZDg41Y9+1Ap1nxI4xlosYUhGfkYkiC23nvbc2M1LwOFool3nSuD+t
UeC7XvgeRBpfgCLZoaPD5zJugK8lF5Y0WrQ5l+goxY6yGa9oT+CcTL2RaqP/sW+B6bwr6p3hZyXn
IyGelLPyj4HUiQMdwVwBKmqhSVJDm9ultDVUhzwHLTkRmCSaJhQ0zeyy0ohAwV3Lr5dN8SJWnSwW
T/WAM3vp5jxdSPUAm5rbZOwhdR6E/p4+2boJ1HF30Wcub806/SMhqLy41VJGG72UVs8CtEta7/Cq
pqsKVRtM0DurVJVkoENVgKWQGP4ImNrHhnIQ4+OXz1mzUuXMzddfWzy7OIW49WKoCch2dCMQkJsF
ZBxvJ2MrvdNkt3eU2/v17BIIaRhJ6AEjMRpuDpECHZsG3i6c6v8MuDI28nX79AWcCEJ/hMDnB3oJ
jie3jlSIl4JmIM8D7VrPbxZbaLeiC4Z376kZmv4Ka70nM89pDBFOqevloLrvU+qaKFTKvQPRFTyk
xzjk6lgA3f4DPmduG1yFEDgBKO85y1eN9e1xPqP0adu82MQ+eOUvA1Oo96MQOa9qC1Pbj8k2MAC2
xz+9E2/MXy7FBE9l8vyTsY2A2K6farqtIrmJmQavDENH+OWMgWscO/FbwxYs1uhz+2hxm8tpqvAK
qDAMtYtu20AVQ9dYHaF6U95kJKxKJfk46UMVnLsby/bxv3hWEQGx4onmqE7mcNBps8FNzweDpaQ5
Y9qtxB0xMJgluQ9f2D0maS0uSJDiL1jjr5SVXr9S0+2Mhgb6xgC2+0K0k98J/7nJtG1Ss1vbywxZ
6+18cQ7o/W1nIsqF+2gQhw9o91pNxdO+UovEiaZhKvjROvlbwQoxHZHpb/LJQJpy6hv9IdcMCaiA
lgMKzkIICVWUgxqcsaCObZO1boMgGmV3QBplEEFFPJVY4URp/ehngETDqNKY8IBvSAVQP79Qwybe
euNsM9wpvk7tYqNJ4xV3Jl5H8LKzJA8DYGieMW5SOiOb5iKjGmjEZu1iHBTh6EM4pBkRbhBak5Jz
NG+8J3rwzSZR+W0nrfLc8H56rZxrTuO1HwGFz6dEEzhLL7QitTMSvXbttuRVVzbP8Bbood0okhk3
XHk2rsK4VWifNQMrcBXR5A8aWrnItQQQv2Wn48QMq2b9y4l/dx5V8pgWR0WHj3oXxNMbDR2L1uDT
9Zk+mFdqilmjujF0cXsPXyqEuZ9dbx5zM/EAzhaArc5Xdrohyy0RHADeQ6b4APpcZl559zQzXW70
LhkT+RVR3DYs2rXywznMF2uX9xGMvkxSszcfm8hZVHE2zPK82DFi+rZndjlv37G3RDOa2HEqxBgc
oF1VwT8BiDiZglNVRotVQHDH8EOtIO7Zs5uO2xLoXhazfu8uhP9VlT0JUt+6l8+s/US+BnlzG7PP
BbM99gIIKsxHlAGus/0b58HyOOpLkKOLisAZHG9F9/habozWv+wGLzsG2YQkBzNGaCR/tCyItGLA
yemq1VUd1fZeG/B5rZi+FLIj9ndQZPYXWos2lBE5KKEzcRjJm+Mif28izzk6FyBgUKdeMol8KARD
CXGTkAUmOkr/MzcCBcvD91/tCUISjUMPUH38zbvSA1mSDwegq6RO1L/bE/5xxsy1tQSpRgWuDgx0
vaMleSEL7p7/dtryqhR6wSYILAntjFnBtzTKdwpTF4pvcVTHNq6JwXTKWIWet2AqjMm83EXjORjJ
oMKK/PKpsVpD9W7RgQqz9pyTrVKGI5NKqbg4sivCavEE0l8paVOIpq2ZlLxgV7zKhxhxU4W5X3dE
vs5VND8noz8HnoWiKSf8vfE1IiZOb9fWFJBgC7wPPBNj6BQf101dI6YWIbpk9LH1lebLwYcMOfwB
nAeW/Ls4yrbs8S+t7Bl1egkdaxarupK3bz7OXMyOCpIeae9OF4CAZ8VLwfkcPuULjI10XmOkVXgw
0L94UxN067pOliheegd9R7Y06B7yg6WWmcd+w5PzN+0lKnTCweKy0CW9cxokYLVa/IPLiNzPD042
fzDrRyOmpjlHwA/fnSDYCQyFSbb5ia8XhjrehoH+AgDBQmzDwrAQ2FvS0xzr4es5GT7sdTT+j/xR
tYSk2iNXP58dC4QHtWuflqWTUUfEsC6TSBCTjLuZzR+0AW2L/Vs3PYfyfjzdGgIh5lrEpvZyFT4D
VUnho+7j7/JDj39V3nG3xkU802rC5991KsKwJtVo05xhwothPyogCEuxmYjJjW82ywBMgVi4IHku
Ja3vH6is1wvvra5qcEU7V8xDJbfXMOPe5Z/SuWmBU0td8Wwtay0FgeByLI+/V9cj7ILjnhKI2FxQ
Q0MIT1fxBoxXyFTeMnHET8pcdW2ARJXQSRen+IRm9ycKVkn+8SOWzrUMFqS5+i5UjJLuofe9uJbl
hFhHsJTpPsJdZb7Mi1ufwpcYBYRVjECtUSaTIjawKxSrToGps+I9N4qQhFMaprCE/D8l6KOMnJxd
i3L+LLrPRLmBstwf2q5UovbJWVzkq34Bocugy35emjI12/FboJbobX/mtIDq769+wcpWvZYdr9Ye
7iJdT5ZRzbktGBb+4rjGOHTyhBppibyPGPP/mCq40mW7tkZ1QSLBuOnYNiin2rPldR3uoBu8ND7W
9MZk/EguZVloIu427ObUiti+v24+t9JRsQAPAfHqHme0rOcvFviXOowilwZ9VNeXGZWqgP2E2x+h
HjWDntxeNV5fvv/crsBIjnTzFfIzZXVskIWtXb0Rwa3/UqYLlWv22gAWFWyJ9Kd9n5agaxr8TDRt
azy2nsArcPrthIoGLGenmLzOA4aQjGDw1vLBPZCFvGaWfyKyBztGKlP8RQ5dXEEMX3RU6XURqZRZ
2aY8br8XSlR/JpSaJ2nLG2DEedVsBYy2m8fKFnWeID4m8wNyxUqlptA8hF6H+mcSvMrekQcGc6Ff
Rp8nWDSlsQ7kSZ7hECzPOyfKXVRxgss/AXRufSd4Xf6+dDHgvRr+gPZAZ/jsVzB56HmPGM4DcyMB
hk7icUa1hN+TWAc9pNwPVHtYxiUyJqY3tN6jVJG+YKEEm0XvXYhhF/xKYhbRcN/uUFLxFH7VehX+
mojxdOQk0uRtFJ7XHH5+ek049Y7ZrFOzTJjX/04rjLyBhhVCTJt0W2sSGjT8OmtQiO1kBB7Eh9rP
0EXZkIocdGbyG1eLZ2eHgTRMO8eCGB6OeJxCqwM5HO3HjFg8WKSoQAM+v1IXmHSOZzSV+Y7ig0sq
HUij05Y6i2X3q++i4R4ZYW9chg7wwEOXXgKcEX5jTfaf04OKEmljAQ9489pfk3cZhJmJxjHonk9e
g332HYuJrdGnv5kdSjSq15cNeVFQfvUxjxusLLDcg/0nCrdgLBFpDocSspYD+Tk4mI/1bMN1lOI7
rz6PCvdtEt57BxDKSNv2rayuCdUTZW4ziwBmTHH6SZmFIhyNwRRT9ebrgi84wef0Wne34tlpEbpL
vHM4wWdIMEvUk3kZqhpsWaE4ykCckf31vGDohf7q/4uoiVlvG7ZCtF762j03dA2VbP4zbxdudJz6
Ds7YmitD1A8tDvaNqpYyQ/ENHRJ8azbJpmxIFBrwT3TV6/cspJXwT/x+t/SaORuArimgA2U63qhl
I16+sC7e+gE4rileNLiM4VwmcXMGB45NPLoYCD+Euw/TdEljctzNoPsD7AsnnVHYWY7t5qCzkxru
MhLM49tkbAGI+fTkKONj1NwZFWyfVj0neuiYuDOlKFChGSZ6PoPIj+ufPlH50go7zNuKmyxiBThO
MpnVNUJTvg7Ijnw+ZPIc1HCkN4ZLYvH8d7/sXkzEp0ZrWudFw8Xwd4NXLVQZJ12x0A2mtuYwsaiL
s9SjD4iRYPOczcHiVoqs7P+oXiZDt/f2uZgx/lH2m4cvewIIe707NY/RXkcNSw6VKqPDalJCV9F/
GVtDDbDcJicDGZkHOhWexvvOXixTNcNdQekkbL8Bp35JYfVGSnBbCbSazFvkAnIQzyatCOhR3J0i
9cJQbYG6nwk7LQAkyglLfuT4OhN44sm+NQVlWkA0tC1Ejg2EJ7st5oNT/q9/S9TowBOtRJADH/qp
EsiJ7G1k0BfR6TCD04LHCafsnAgYeGAAsYAxL+RGs11QhdXGK02pWtUFMcpHEtjta25aGupaci8m
XoJBBnVm2ALru76FGHAthAlGKzwUNmx4Wd9vl0VkoEqgx3cRa+mQfmcwN5K21Qp6a8HE1Ij6VwdH
7l9W7QpTdtqM4vPkEqNrBQvaIxYNeNwoiCFG7Cbcc8106RA5VFivEj4l55NJaPVyls8xywP6T04X
AbtQSdn2tovvoRcIES9zqvZuBQZFaclk0wlHuLv5BQ7haBdNAy3PpuVKsukTR6YFyPxUyU+Tno39
ITndVuVhmm1tna7kdZzBuvl/MVODVryZC9Psa8SwQj/prQD0r6tQY4N0tlS2pan5zp2aTmTwKTrD
+R6Z0dIjkM7Dasp7Ip+yyKpXQJAy8MCG2f0gVQ7P4/R3ny3s33YD/q7VMHSP7q2Kgt8hKd8BgT3M
d6NUU+5hEMysifGf49K20Q8u4OCpjpLRY2LUdWXi3716YA/IA+rYHMzfhENfjdmKu9PtzSsl4eW6
UsQa9vC1h5nZFyXCoL4kDH4Iny/rMPJgDWget8buF1BnaJay2Vqihr1nZpMrAXlzGgvmIJmrFH0c
5FNa+Kr3XRRRZX55iB059/wdWn/G2WkXAcsri9bNLlOWUrnBDNSxugFrRNp/jbPtYXrwiGhxOjaN
5NLGmDEQ9DMJcbj3HpH/XLEx+PKUvHc31R1V1ULlQUsM5wUo1COAgEQurAhculj5uAzehY7Qn4zK
/xPc5eVdGxgU2FfchGEVRw0Hjif149096TNNwM5iE3k8kQLRHjM+rajM6Zz74TkWZwF5I/DiQeQ4
VoqDYJ80jK4dJ+tgWQBa5t9bQ4T/SNwXxgLvhpajBGQYLYExAJ9SQUMUGeUTYlhDcVUOfa8sHR00
vG1nbCVu2jeJVgEzOxKhf6OaxczWsxdWMCFeyUiqCCC/Qj7RFkpr02ArSVx5oRBv+OqTNF8TZIRS
/vWl6V4HSY4Z2KWkvJV0WcsICb6SxUqLmWsp8EUUxGJQ0KWV9IBrlYlrgB7TQDnuV5BjHLsR/ACX
oGKOwUrSoaKntkTpwmOLiTK9BMBYqoW/gUfoybY2E0ujC92Fg9YKz8+h9TpEisVGIdVrSq//XRmc
E3+XMrgebc0Qxus2zPB9zEhaigKybXIHqAZprEicjbuKj25Zc2HdWbvHTYSoAT9Swmt0LV32eBOo
kXyTgbpJbbjGeNieBZ2X6WyvSKCf98vsCv8ueOTRtRvmzcgNUVu9bc1ID6eKBZtebvbPNee38VzU
ADKIjzUoV5D5GiOEjpxCmSJgtLpRnUeh5JQvA5CkByy36FkPN621yYK7KBHcCP9bx/XSd65ZDoM0
YErDsJYkfMCZE9VeS5eFCgZYTnqOP/g+/VgLrdOiTCW+gTXGwjQBIX0EtQ2Ioijek3uX7sXheVIT
qn2j2VCy2GcU5eniVJQiEySiunatul5UGaLd0fJuKCM1+rFlbHFMlxz4bNRrE7OPSvtV/dS73LtS
xK/Z+z00vpl/EK1ZYHhiJjMF+mHAfTFhO+iNtQNBWh54a7WXn/zzu2a/b1Jcz7v+jFXkZSWFpuMy
chYPZxsXkMR2C3+x8lfVijQh/ceX131ZG3oVf2j3GjxPsXvKbuEp+WXZny6G+xnnsWx67eMdU76D
CrtQA6ie2C64E1b7LuL7vMSVbCD7I8rnJsFAWAQuAcIctJ/X7COCqVp2T2ayXtYTMhCLVe9M/Zcn
pTWZpLKaZtP41oLVBRfY+KxQnNkhxbW9U1GaZAvp8DYDeXpUAgOSGr7WLVQGejzS8FLsG6DqyoGy
qMASMIV5To5vrNa87jaSBgyl311Jlwn4MHKk8dAkZHFnSn3YY4ol6Umssc9cnltL2/XGu3Tcufeo
MjuTqqbSiSeYYuYctRCrVWqJiZ4FEYhWRTd+ID3JBOv3aupIE7iAwYSslERs7Rgs5SKDJpr6/ogU
GOMbefU12SX5JVFAyrrEL2RqsGdG0SEUBDNexBTquSRNHbi1Q2TdUKxsCFne/LH/Iw4t9qQvWwhc
rzVozeG21aY2KXNaIFge5en3TC9tMKWZ2u1Gsdmz3a4atbSbx31oDt0x7UOzgMJ8ce4b0Vc36ycA
fSBl9lgx1YZB/yWK3vbh2tyVM5HzwMwmtonELBSAcozPmDyVm47xE95rXmMgmMy0VF0XPSjzrnGY
NAVMdmbR6MK4pk43DT6Rbw3Yl7xaVj32zQ9OKlNQ9XXA3FuIzonuv5qomIkn131oXPwv+3Zr4aFQ
1Ty83cGiqsHi+9cnDxKtuZA58E0wPKGFya8zvOZQB9kcl/E3abSr/ZOWpGp0nAI2kR+IMA4o35HR
UfVDvNm0p6xRnCWUrFmF+Srl93PTC3oLmNMIYF68JTzsLe2LgGbUyd/Ypb5ZR/G/tqSki+bFNaiD
O700lkqEqq9sMI33AO2sIwACHm26AoI4d1iSekI7vcJtQTw0jf3J41HwaakyoZr87TawcWSxePXB
0DZM72+5y3hoVSrqLWD4isoeup0ErcbLlREI9GphLMtYHgS2yc8riWQ4/gaGzhiKQANKkExZ+tI/
vkK7m02qn5/785OMqpY1w0A0H2QB6NMea+aWDsktgDGCRFwOhEg4GcM0svmjWrlrzaefj47NR9wf
hr/Rv9syU626renDxINqtHnvcEHGBHwoZav+GL3W3o0+b1jDS+cYJLpHoltzoX+xcbHKRvCNkaWh
ik0r5BNKtn3FltLOePWXy5OHfpSiKSXYByDjrRmp4slCkhLM+cKfHdOeyfAp+N13APmF5U/Q55SD
P01dm2Yl9u2tOh/reJrEY32XBuiFgq4UPxw9W36ed4KxKzu1aZ0Fs63FPB2WoYZNpy3HtOa5scN+
BWUgifzbuHM+LNQXpzqtrObTF6N5/8pU8dvJXMcEL0gpTQnecjP4ZzIMTskc7eeqapjyIqzCdaI1
h2c2RLPzG5r0xyZ8OaQ/AY8HH9oBv8SpbWJDDruzTK90QTvmb4c1VzXl5E6IRrFxQfg5nIDaq5bj
UBgKRP1q9pzb4EH3rQz5mU4Pf4LKt2g/OCGdtAwjUBdoV0e1mD7SksJN7BqB9IXIazwI64xLOIU3
oF335v5qBywOJIEdwAYZSMNdTc9tmSCxlPCWkLmZW9UGSTHjec4PLDYcB9hy9igXKR/nLoq+9FZK
Lp9gSwvBeWrx/BhWJ7kDXvr97mm5wqmVR6QkCnDVRg9B+3fGBzmUZ5QMgBVYxP76ApyXWvoKj5DF
Z2mIJXpXHhmqgjG52D1OXPA+672I4bFmYcxl6EQ6zwRcir9pwk01IPUdfOb+xCc+X40dQvVvZqtg
PHgWKqQuKWdJg6jX/09p3G4MyUSRME/pTwLUpBh4XgCt/PqGa31vLDXm71Py9UcQsMbd1aEWSgSz
m/KQEmVDQm/7O4dfDMSJmCUv/B0xZAM+MRHcch1h36h7XbsUUR3SNrr4U5RMykqO8MDVhxEdjiER
fSFMePECCb1etpLuSYLu2Fntgb+bWYpzCU4STbgebazdMEapPz35T0b4B5bSyT83Tx05b/nMrQtK
taGw7g7RyLVBFBTGLiSmkMNh3uN7gmx5cFrUKfnMkHZ8ys+ovYAA5+7foabauxa25L5l3BOTl/mF
oJVO1pI3JusM4bdXl+TFnXBbEZcSVknoXKBKCJk5mlj5PXkbCXaJFL56bYma6DPMqy3DhYvzZ+7A
BXmwZzIXYkrPssOxnAcs/+xRd5qQjQfiw6PHGvnEC/20uJZXt7YC2HBIf8ovA3ukcR31sYGg0nZ0
rmAc0CPd3YwteANi2Wyh0YZCgv5SgVT+jivAkt47I/S7Hj/OIexAmwIXxyaISVHSMu3sFfwSxf0q
zPINqX71B0KkMQ+8UVU3z60RMk3Weeg5ROpO5qkCDdS2aSx4OASKFophIOxNam0zrsdoTzhtxN65
wBdA8vZHtvgJlbfMbj7foOSfUleyY5+1mNvbW34+WD62pRwc0H90QNIAuEpTwPlimlNc7LH+fW2P
7MKiF6D5X+LNY1e48y1R4PI85tvEenxkmQ//0qO0O7WHrzuVRlE7wF4pRtUpJ/VT1nrt3peK4ySw
bleQIPsmUwJRoRBq8qlFJMFnyBoIDSPJ+lZi9JPn5tT+Yx+O7Yq1qLDwRFdnBUxdKVwIfRo8eNC+
ifOZjYCbzL+vsk447Tni/TANWwEDh8zmlTRDV106a2w2bV6H0ZhAiDyHFGWxQAF+ZqZQ45ve7Vxm
YpkCbgx2bT6keV57d0ZtFh4pXzabQXnWrVYrPsMZzUqkgrKjWDv09e1wlsadJwU3IXRZU6jfUtdi
IDhocbSPs0Vb8LHtovzYt+SGNRlAbFhKELUu7YueDJCCRJleTm1NEPy3P2zIfHLe5OunmPHgfOro
XtwGDXbyl0IJcmTWDhKiw8lx3OejVM6zyt0fOdfbgxdlW2wXRqgQRod66bOyjXW6VsVRQNTp7/aa
rSKuI4BtmWBNVVG8dtXvk266u2r7KONBdJtmVRxeq0rcNkEJEO5nW7mufH+lOPtzEaQam33PojnC
7UBDb1lWevnUmZAYpJYpYOnZr44vv66/aOgA1Noxlo5K5wBoXc3ywnJk/VnWpOMu5q0CVSBMvx98
yBDTBqy9Wxr9U+NPhBUqBvvEUaWuyP01bhKsbkjQF8IBKh1R9qtQM37VefsEoQMNt484Ge8SLQIj
JP+w3y9l7XeRL5auyEDYm28RsLdTCqCMUsdIDUuw18O+bAj86pMcJ+wWM9D/NQP/7Kt+F/gOyWRI
HUV+rsPBHGXeo5B13+643LFruxK8A4FsImYMTFDP7M0YSEhcs3s23OoJzoq7LuQNP7Qtl3wWTHZe
dgb67WHvTPE6Ig7hVEndwgeNAIoM2+rE6eNSM6P62muhcdMis1o2/NfNH0tmqYeNzeh++JG/vcSJ
jjHgpsIfDNNMqPAzTXB6y8T4ZdKuuyliB3VKVwyzXAXAZ9ty+9VLGvisr7mmQV37QiNcDGVtiEuk
7DltEEHB9WoSPR4+lbeSTI/HiI0R9Yg5z3LnhEsK26IXFMtAEU5H11d8DzbD2btBOyIKJmzYASYF
oNa7E+eAo8MJ0bsaLfzb2WIS+lvg9R7zWcMYh0EMDpwW63RucGmAInClputPEisO7WTkgnGV6qGu
wc5bvWu72+CfMwAM36qEhHy5m8WH/CjwJmY7EMUsf+H9DXZtcCambpVCchvF7M0xrVJRBXELmc25
UIeDzIMAlr5Oc1X6+sqXIBLhJNFM/Osk7XFUsXmeQUuwSg9n60p9Nsgo4NEIESnHWDd/236BGmUo
u9QaSj/D9pg1KigaIF1U8ms7M47G6FH2BYmJg5qIt4o6373gstl3CH3StsKFJax7fRGc4Ae+B19F
cjZr2vqUc8OyuE95UV7z2NkDJDxqGMSK4t065u3y5MfapEfInDDI3qa0bd0kCEy/i9F6qZ20PR7X
pcKObd4hiRRzWwtg56/Al7fJG46yTU8gUM0fC1Pmkm9H8gV8rHQBk4bgvTV/UeIQpFVLKSOeNnxq
az70112doWUKQ8N2Em27oVDMfOEEAekTPVmgAGC9ag3hyvyWBULLnVEYxpeSHTDQv+dNs40YBq/o
k9DMmP95xhmJXOqRHa6k3IPQXWR/nKY+cgHYF+xWpYRGnOnBb3jgljd+6YJfn7tpX2DNQFKuKx9c
YyyujN7KT3/VxSvQpMDpGOseHY258L56WEilkM5rMur68vDr4JJ6HhiRPN/CsxMsspmUkjK0tgbf
ddQQAJvvCCYXMVKBN3cOKYL0bTA3edkLCx01+woM4q+JIIrcM+klHWE5xhjxorETcoTwiz16JeRN
FhnkeUpWX4Hby2RONuGX5nfmfMKXEuPJmJU75YKFL8MC4+gMa70TlAmKnlGRAyvapOZvEvw2mY+z
vDrzJjEokxP/0oQkcrIFVeMwjA+z4SOI5+he48ukyC3mNlqyif7Snz7nWz8Dkkl4E19+dkh7Df++
QqYygMsBFpSSDTU7zl2gCiocLCZ9BdBpncsba9++kK8iiFjC9uMKtktarT0oC68o6cnXkUOC+mAg
xkv2pgtBwC8V7XzVwrxfLZ8h3QmtXbfE5eJfJUiO1u1O9y7cINkFVUkTe0W/UVzZQRwsst4d3+AN
0zxj8+Q2C+Bz1mHEWr0lnClKvBgEn2mzYko4v2pSnPaaOqUJHqmDoTxvXMqVTbLpQ2djx1Fxc6n9
txxvrlsxsopnxbDEX4tSoQ/9VDvM8cUYMjLQCLpHg6bxZu6q2DHF0/L4CzbKgSZIkzL8jT6LtrgX
G/pnNJHimvYxvZVvhSDFL/jiIsiu5+Z0wCWxrN6SjHbmYgLupwvbXaAgeiT6SuZMBxZ1vuFS06kJ
KMiOwbrkcOA/YmWypVZo+qlOQ7M7Z5gl3R/s6gW0xJdIdnpYfohajDSCC2eLgFbE599CiINyZjSZ
2CxufXIbzumLMMQbPRuLyb4FAxcxUzzh/P0fiVrht15PoQe2dL2Ww2b+hbOcyFmR+Y1W8pczUczL
Qv6xZUk1OZGHQn9hC/fk6SP5F4GwQ85fC5MYWcslQOYNf4XHU9hHFNI9yvadojs2q2Sg/D52NLzY
+HNaabfVG+tkvv5fpoajtnJVIvuXayakMF518baBK1IXyihy14PB37A9JQg/hha2hzx8Zk9T/NAJ
BcvP4wR8LEcHqM1TMUveLcUv1JNKmsrwlebQ59e9yhiXmEBkkP8YgRaboK+jPDRRS7s7rknnA3Ol
Uj+Dcae9KeJIbd1qClqOLEd+xcochlkxaJORaAYT5YzOxE8sokX3ZzeFh9IseVrdy8ikwsPjzq3U
K2R3ItvpjyclPvtMdXGuLI7wFrZL22f3eoiq/J6vZArXNTCKKIX4XpwvjfM30KXXBpxheWJiWSfD
Vdc8glHvv5hPizw/rcZYu0PUbT92ogcz7C0rhSnZREc6xT1SdpMtQDv1wiXbo4W89htcEodDp8vs
f9ewhT6mJ+kqV0JrEtJf1acnFaIWt/DuVtiAhaJnyxpXNX819obDGWQjczvQkNfCQmnS0STdRoz+
Ys6gRHGlQMFIFRIpeW90YwGkAu7dgV0x8qhb44usVKK3Z1xa9bSWh6bUgpuAhTRC3A692QiYMp+b
HNho2AZkPU0wMNiDg6A0xutFgijvDIYLkNHr4tyGuO/P4NYNHnzgeQcnJFMQuUYHO6oFN1g0d7Nt
mQhaCvnOHpXuEDc0JEXmN59Y8lvJkFArEkn7aZVjWljGmvA9u6VuBqROYRmysmN+V724aUBbh7C5
16nOvSwFP1/sTThUy16urzCqfs8Xnxt5N/B6cVUFGgJVTla1qWK788ctrLCytwQUKU0GgTjmBVeW
YnXoRZaNaqOnyyjNc+BL/TglpOaA5sPmxHcZjECW0T+2OQfM7nqBADyAuynUnGOaV8jsiqXqUs4W
TX2CSLtP4ZrpA26l0AB4BKbVNE4iR4PuaA+6Ql2sXc/64zeq14OLp9SerCmhTopZ0uL9hY1Cgpoa
2/jj11mnm71jNIP5VzdCdSpC/NusovTMWA9raK1e/m7I261C/VkM8o+i4xepqngyfTs39vOlGaGs
1zjiTnIfWM8L0vbz6JmXQcG5aWAVuO+wjwClkBTh5HEsLaEvtw24Ikt2gCd5ASS64pdh1zPyW+A7
dAwgqsV3IXQNTzhVPBzBupRFMXuEvVtn7ZBVCeTo3x6XRXHDCdCM3kqrvFT3LQEM1xnHS8TKAo9C
Oyam1YsIDsJt3usyruNoeOWRAqnTWFrQVGiulkkBssHLm2gg299jBeAH9ezEmjqtNemylw14m5ks
7pft+eJtnikuLU0BPrZYmDFftgFql6gSv/4WeUkvQ/dVWSe1D60F6V9BDV1xvHI4KrG1Y/WKbJ6J
weLEshYOALxlasxpLbSiTrIihZYtKh89V5m9I1MU5ZGB3E3Zbg9Nq4zBeK2xL6DaLvnoNgx9hBKE
nMjPqigFbhFQDZr6S2O67c0r+prGzgUgOJ+YRTG2ilL9C5/ykdeh+f7zkDN4Sr836v/lfSt9yCV5
R6gGcQAER16CaVn1BBs/YyjbnTuixGc7CeyA0HZSvXw1k2Nl5f/61HW7pto9uKBnpLtSEahooSKV
c+Bicx1gVUWC2iPyagQ3NU8HF0yNYVmW3p5yD2EErA7VAnJuQjUEYqIc6wtPgOxi1+SoJ4wGmxoQ
GIhhWYnp/Duuxi8S7yjluWbj8RajbDx2Fh4vN1nJKZrEI8eEIJTcRNKDO3Ggqq9uRPM6txa8RjNr
5e1SLZCpfsxpSsFeUHCbkXwaBQHQGJ4pf7EzCeK6g+oKnwiXRtn1v5tPUrNQ+ZG5hXM3n6vRkoh1
34kVfbAnVrYF9nWZAzSfTdLWn9RUxR8X+os0IkaB0Xl9xL8qc1rHpLFtDHWgTgTauRg33N16CWGE
3txrSOqlR9614ADGKNMktyxp63f/+G6yMGsfFKNLFh6LhV5tg6YTadjenjpU9UECN07gwRcXAD9b
SfChYSsxA0EuihV8qYejqhIJPPZX0DS1Qh4N+Wz0p/XhOUd20BI8Hyk9c/txU7FH4H0WSRxanBLx
YWnKK2/HvFAc9KFjq1rjvGDupqLbjkDTK6nSg2SemRk/DZwp0eR4keRl/0g/3pUfY6YHONTGC8hx
zy/0Swvg9OhbzEapUlE9ZPktIsw1iQNuQ9ZIHSb91/BV+pGTYhuibCt+6KKx8Du4bQhHV+5nSNh/
QngfQCXGpzyZG5lT/tSLXmLKmCa7tezI3Qc7urjWPu55fEWVr11fTlsUyWI0Gmc8YQHyedQagPIA
suBVefbcqYIovr5lxLVD/0fwFTi4fQDTd6uQ0j2s1a3ssYklF0yJKi3PUtZFJZON/sOuLJv0vuZd
hwbKZAVl+yf7O4kZzM84WzjotFDfTjz22U2E7RZ6KMiWkg1/oYR7t435mrZs0fkGFyexWSlzNFIh
WWTqMHkMQk8aLyEk7I8SFu/IzNDleek0AyNJgyMuLgi1m6jG7R19L3yAq1bnsieaf0/EowoR2cxW
yh3tWYPEMpB89lHAgkDrEGyoyUgh6RezgKP8IzB5/Kt0CwhyJgaWHkFdhmj1fIEkJbxZishvOwQI
W+/uWmiekB59kqgSXjRIrvQ1v0kmMlZpoqA/FSGE8xnFJ5I7cB+CwRshqqi1TYB6M8hSK2jjsXP1
YXHZUMnNm8eP3H+CAcKdr5H3rHV8J+KSKFFF487LXeLR9kr7w9AO8yGRoMk7QnE0VAHcvHW1oL3H
3sA5cXa0/dV76EfK0j1W9hIN7JTql3HhjfIyRvOQjeuW5dRYE6J9WmnohLRaFiR/Lv/GwTlhBcF5
CkrORsZxfIV7GXsVg9ZfL7dLVJJgdbEiiYVkJjlQ4+5YFD0b7KWjG6cHVm8j6+GkG72jnCt8M6+c
8Bf5Im9R3/EttZS8+BGYUKOgzmpSQbn9P8kpaA7sGA7g2JX8Gvwrqsr+eURbFZJnFemCkcAhh9+M
lAJg9Y34QtnUx9akRXur8rFvAbOLXLZu7F0m5row7BmfyiCP85vLHgw8WfFugMXmdagsl1jbBEA0
IylY8U5DegAvIutEGYzh86kLC9m/iHmLRr3dDtc8l8jHqbTH/oNCebbD/D9Qn1KO0sKS9+qlZuru
buf42uAFml/16KU4YmJS5vQUD4/IrXopv+5AkKZ+OshQKupXPrq7FqGwc3FndphfaD+gl0wKKnEy
qjGma8Mtm2jRy7v8phtw9eWAgoL3dp5aBZqMdF51BVWFLXCd74XYFAKAZ3uHLlpWcrMhEAUGwkIm
OfDPEl3DhJrWbtKUx4Fu+Z+qJMRvjXnHAGyzvRgagqZyz9hBjJLnCgNb42n2nHnm2miKTacXDicR
7k8Q8XGf4dDtZy5Gy8/EOzFI8jcTz4L7iTPoqG00Kcn37NaVoVNbCWO8EkmqvvNXsbCVdlrFPO2t
ZQqaOYd2BQnR+E6k+amdQx+dLzBX9kRDDHUbr8AekrebYFZ81fGmPpIiW29VGiM94tlG6elvAJZT
kkdLScz6Xu0MZGw9hOiD7gqK+kXe8WQl0FlaR54N66bs8HHU5zmmueSXJcDlPpUhnfXSNOI9BxCx
Y9A3WhyChvRYmx8cbkUatK7c+n/f9nn04RjAaZQ4nVQ7fblCyBc3Xxg2bmzH3R0aWU7nXQ0/aMxK
hL0bZkL6E3u8HOBwFCoavy9SHIoTKp+WufCMxRDGWDPGBmwFxlPODodaL120pP3ZF+0HH1WBCt1l
UJ79y+TNS03SEdQbCo1TCA/x5IOSZ9T2nhecEicdlHPSFhOKKxXRiOjx+lydVRfzAiMTwoueRXZA
VREU54zXas0hee8CUN8s62axlcvCr571K41OMKqmX+p9PU9B5CIsHEO68eYAaNywtExAUTZvrfv8
lMhi1T3YQaWSRLAcLkNx9Yt4wpylSoewe5/Y2Rkju3LBhKzNIAMc4QfCw2H28EDJ9/H7gGL6gH8C
BuSj/GxH9xTl4IZ+B9+LjmKvtb9ZElHemZ14eZ3uUAhD4aRXj63dhuZbXkmx+fudM4cj826Z3YS4
usb/PrwzfO97+0hYglT5ERX5LSOb8yFHlZA3j4iNOrDMiUY0PnoAxc8C/oU+etp4qR5/LY0YtCOb
ZOefUtUVVv9EU5smE39GUmUlsKkZri4P37GHQbkNkw1wvR8Jc42Aot22tqbz54ywGPv5DMRytFci
4+OK3px6A8bEibH82KaH7ULJiVc7Jjkv/DvlWV+3VgERKvkvSGiDEFRutBIma8Gl7VPkB/J/iouO
jpi/j9SSsX8bm8S1YRxuyVyWpHJ5nhYnTSpYA2D6Z/3XHykJiqVDjNuhY8OFdq2jlpLX7BuwoR49
ezzuuz1Qtzs1byG5RqX80HE7nc/o4RBCJsctQq1DJLOp5OlojDlOC1sMkrLoU4AqZW+/U0o1t/b4
4eAGtXW7soRtmWAECpdL+r1krOojPyPEmJ5vetvPmG1puk8APFcQnfk+G87OO16px+k54AEmrwtf
SJkf2gdBLgh4Sah4bPLMJLkFMaGb8oYsMONVo/LXeU72vkhTTeo3I9TpkxrE9HTBdbxEjXp192RA
Uy8jE5rODuVqglFIad0Xq5AnY98Yc5jSUJBd4Gh8HP3BBbICqfTQZxgEX52AU06AWQL5mq2SC7zY
lazzQXQHrESCemYtQF6fRxK0A04I+y5jxpSxsIIE+qypqDaKC0GHpiYAbclM8HmihtFyP7WKenW1
zOJi0B86nzNQQRI6qLZbGFHiFM+GLEc7j66zBULvZXUJ0lPwQAss5zBx5TWLc/XOBwYlGqfBEZpe
9jd/wvSLgtTHp8oXvqB/IzxOJI/p2fcXEnMAebeB5dnYfQ0NVJiVunVFA6AIMRiq/3X4PUH47dij
mK7qGyaZi5ZWpARwCFJRTKErWtoY7VVX2yHkFouyRJli7/p8B1NnGPpXMAtchKe7O2lF/EcKslPL
Gf2TaSvZN1wlSgHIFFXq+x79Wjv78Rkf7nQW8ZyNmFizCBvi3Qo/ZWjC0BGFMkKUhRl2DG0+1IYk
JqAeg/yRomYQrKYRP+SQUT1TNW3fh7GdF3HIa1EaFrpsUxlDSpwN+AV6dxJsMo4vjbvsr3gWYyMd
s0hrXQ5dXfBIFOF7xJQfE2pnt4+EezqDeaWH2fzOazjatMWheU5iOaVldnNKN4O0Nkz8LOdbfSCj
spRvuPyNkt+oIhYIxegpDWp6oiTAYVP5260Gu/7yGxZcSdKWnoZDElltFlVaRfAgEodhJ+D2EEM4
muTM4mVpcTlWb4kJBGWhnXte0XC9MjzoiXh3S970zV1ZMtM+wLRvTodkw03Fx1OCI0pzvlqyEunv
6855kj32bHOnK+gvAiWFutBu1a+8kAEyFQNIpulxJ3J1KBuYJcCxa/uY5L9WdgkHfuCuXlAo3JXZ
zOcMnUBHxdqrQl4GknhS+v0+0rx6FPFoYDZivWZj+v1MSZUfrr1XJtg3I8k6z4CJspVh52e6DOXO
bz4D75sISpWgL2B0Awg6BM9XN43zrLHbH889mBg/j6Pbz5voafgK08zAEJUvtAaHVgEfdZqbh5A6
vH8CxYs/b/vjCoJV46fQkyynB8QNyO+MNLfXVSg1NqeYtcDP+wtpDdRiVta8R3msLOlzRVpVsCko
U8J02UUiduvoJZWRgdk3Hda4sR4glFnMeVdCbVXiPo+oJry/pjiW04HdKxhBHLWuG5QdFby3RtTc
IouCsPAcVBDUA7Ga+I6HWuBy0+U6NsHqTWUiqGGfnOsKZzAMolZvOsap+bseH/nHQP/I3RJMBf3G
MS8xnNG4sawu5MRyYWojIs3n6dQlO4M38MaoqPMF16391rlWxf+d6uNtxjhEqsnfM7D6GiRDozGy
DPF6S9P96riGPlU0PnjD2g7mQjKe8qHKsSbyVOOaIQV95mc/ajHU8KRTcW7oiJhxlLTvKm0l18E8
xztEwf27Ff6jMgIC7WGenET9sKmPk1JepRGcN5eCJMDMHPumsQ8VT40wfwI3uU/w2Qbc7pKHeInw
OBtlM7CErJjxzyeso5lviDxIj8StpxQjbzTJep7eOpJQfqFV0mXh9E8LiBDXkikgS5V1l6mINuVj
EjlY0o9RdkEmYsXaCi/NI+4rEqyrGoLK9UxZ2hzY9MP3tpOZzFXNyMFQO7B53s3wh/2g7yEWSQMF
h9+B//4BlX0k5SbGnOr8Ry135OTI7tXeg/IatOmlivuQoyITYC+ap8K/AFc0fKb0EJqwgOkTIOuU
5t2dMyJyF/+VJGIrzh6atBTDpyAgwuOTikzedELVfwW9O3Ox1c2x/PUT4WCF2K4eRzOiLeC2pSur
MhJ/8EUQiqny1esU22NOi7zNiR+HvmotvUkWJf9zi0DSgVKD+VnZvm5w3XzPgmCr/NQV/qiNVoPd
ErNfAGPGQDNfcQXvCVXY6x9T6JrRU66/f5zodWKjPTBihqIWgogWetSYO54xu5mr/27MqLqweqCg
i9+d3JnkCb8jXmJd/xBRuCY747XluQvOGerI3U/dhHslXAeZRgo+4Okp5ZX8dp++t9ZSFl4eMGaP
wDWtAgbgsNYfsYLgNweuXygOyCtsuXA+TGurLAinqwW1n3Y7d6RM9Xf8T8+MnlkZwWLlAetcnIvx
mcR/pdGFDu5J3wUTd4OXQA5QXTlOTfoURDZiu/Etcy1WWKWNOv36Ng3FKWClfwGOuayrDf7Pp7c6
zDkv6eitKi+NWeafbo9JF/915/aZGKS4jWOSb9U7ad15RcrIXo6ivdzl+dcPZmRKHu8mDFs38zwE
bP7fgoGH15KAB8CEY4x9n9JXjApoXbaCdL02xa7kFzr0GA86DEbqP4oi86iHR8RQsX5UwpvND3Qf
7c8/rGO3l12wPRVc3Buzq/HrBujQaqGZJnXlkVueVZCENGXhGrb6sttUhIb92RfgFH9AvOXOJuQn
L9l2uOpNFdhm23Pwts8Ap63tJAbrsfBs3ENS6y6CeAnxiNC4Bwk7O6hqffehyXH9IM5gXMLQhssP
29l8QZICeeWISTIFslHGsCciAFpbRhqvqau3INr5y77wdygmpQgauDl60XVihmV4IcTx1FAmH+iJ
KX9QaJ4cx0gPidgViZD488GFmxa3pbRLAtFe3Q2aTOmxdhucHxqaTjkaoqTkiFeCGGuqt9QX7sY+
bRuHcD9hNZhDgH0OJEXb3AdQr712lAILWUhhRIlu6pOJNwstArTM/eJdLLCV0ox3EgtDkuem9fsM
o9WOhSaawdjPTWcBklDrq4S5SKzSOmKM6KNYByMGZzHaXGfkPesZTN0k9e8KVKuRFPuuhVHcJUvd
2Y96476zCgnULfvkV5Arn3ZPl20grirXRyF8vXJu/SyIx4VHZXEnpzl1/ojqsmG69cmbi3LuIBLj
QICYGQ/Xd/eTHr8eReepeZ+3d847L/chs1/Kt2yexGtlLCtZCWhGaGoXcc+sKNy50TtvmwPVH8tB
4AYMtz6uQgNAzIsFtqQQi6lldezY5ZveHFKf23AQys5CLqH6E1ffWJbGuApEmdIQmeQe9bqMVjue
3unhMSfrvZjBurLnbWcG+uC8fKI9BnVJHQ3XjJi3QaAUmS2TyRuRP9QtCJvtWPLUPaZlx4T9aYcL
lXjYgk/A9EAhhwGXEVATZb55EbzUSLFllg5/scCIP9ibonDwXA2p/icqDHxQZq63vcl1kqjBRSEi
YUKjEOsukdJaXN83w21SeL58b5oxC5eJ+hlIwrGm0MfOyhMeyOLR6td1bnucHFNvqSyy0h6N2YIi
n6i2TI7g+qhqiUkJH9/RxKyfV74hUUIHVlOfqw3JZlYHm6IaZTQwz6+i4KGS7sRmV/KKtBlGnG1K
RIX14jWSsONaTUAb0IKcqW8G850sSn47ty4SPsgt4Qv4q9+I7DEWfLf9VExTbsyiD67CJ05NuUDk
LT/gfMp+VDpQpHHXld3URODsmn7V5Y/6/AZzK7B8Wt+U4jsD9P4aTP/fubv3Z93yoiV+FhsdvJFp
tqp/YOf+esXx1pQA68/TrtldzJV3Y7eAFU8s3CkzjfKSDYXEPUEQG0pqQkNmC/LxsckDLbFgv69x
ydBmdUAjANSCrXPRnEftwEppH1H/GAM1sO2T5ew2siefc2G3VhnYeLtmL6DAj1Mk3cR5zxBz/Nsn
3xdO+fZZVfu6hAdJZyI6V+IrxsjjASLxrUW60UjaLrIad3ZYFrPUn1lJBQE+w44d+RzIXv37AKT1
1RzOzv3ftj889JvcggZXHWQzaMuFWbVgF9hHIwm9+BWaZ4eloJLJYSvrxKw2KNkOaJwo6nqF6pM0
D+0c1fzMo+W6GZ4tDreyifxqJSd6vgm01IB8LokPWFSuaVoBWMcGNK9KtVY0dJXLWrFuNuVdyxNR
fcnt9io99Ey8FT7c3/vF86irA/gR2BRm3k0Z9l0VGh1e3rsGQ/ABW0zG/NkoclaFUhIW72bLPZ70
C1MIFMeUTTI6gmLiBKxtTCZ0/ebH2WgKFfq+x+VhXo58MfbwcNKjGds783sIhLH2Gh5rWnFNbWZA
Tm6CG7iHAlqRBUmRSM1PPSz4T8jvw5XLOplfXGl1yO8OVBwbC5sngFbR62dHj+ZXVb//Wq8/DzkN
RzQVBGXK9qKsFv9ndZ+QyqI9Pu1tKUiRKq2mNdqeOtPo/CnnhP8Ddu+9eU0G9F7EIaMUhW2fhUz+
gbwbfoSyzoIw9dJU2tDSyr2fi5a4IlgH7SLTCLA3IfteLlBv9Evq69sPWobu0bf12DtE2AZiEaI4
H084FMGAt+USTtsRsnEX04fBbHtxaqsWGnnDuSvYbP+tBTrysaOH4VeHFkRLcaGeZsDX5IvQNYAN
m4z+3gCc4qbS90FJzO+kvKaCh8/udqiLeYwkacjs3TIvzQR44rpYOSGZrCeRCGq/iL/gHc524N5E
/rwjuFB5VUYGt7/9zSAc5qYTFkutgAL+sufzygHUW0gtCFAtJeLzX63+xYqjJ37hGv/MU5dQ5qLs
c1tf4AeGHHdqEfBJXOYqT2QXW+hUOghOr2QohCoubkkahxhB8+DP4UXTDaMJVcn8v72+SiYhYqzp
koEHA9O/80yRrJnLinBz7b9weHoBeMKp9qENvw0aLSxVB+NwdFBaNNJdBAPNdZ1oJB9pNcdkJhLX
7uNkKWruDWEm0xSzGLsfsSuHRHazo8hvAAKfT4P5NWr4KUvw3nCF1bP+Q868AjfX+EeJ6tNbPE8Q
bclOZmylauTxbukyBarWbxLJNnNn/8TDUUGRUVoCPdODxO7xYyrAur3HhSp/rjMyGcMA9TPp2Cbl
8MYqkYhHTlmu+uFyTfPXFDRRtKlJPLjXLTud3BQuc6VzB7AOQs2H+AOf8Ie04ZhZZTfc/1Tv975F
ofQmi4sV/N1PAt7OxgULqwLo3ysnWvoO3OPoCw97rPVib9Te7+rHsWU3U274rOr5jooEJyigcbCU
5+Zfyn29AUi4/ykS2YQvqX98IpoBbi49WWtpCqi2eCLjYMi3aVwZVD8Zy8lQni/bBeeTiLqVjjhV
MIEHiVjfR52DQpz8fv7NpMt6meJaZveUce+W+fVDLs2LmJvW90wf2OrFEr8o0WXyo9skbKMk5Csq
osn2QZSpLl9zgql5XAIsVr6Uh0x04EvtDNVkf+LW8o9ciCo1J6UFVhZ2LFINW2yrn+s0JmU8xICI
Oo/fS1sGvmpFK/vH2hriQjJK61nS1EU8vXzBn4jeYGZ+rM5ktXPVSm6vs3Z/vfPe5rXTKusezx4r
ohVY3169yDss9xLZAsCeEbOSKlqrdwAzFTggddUow9rpsEhkYO+JGNSAv7sqYmUcTtRiqSa0IKAB
IsE7rHMP5ZbN+mnT6zL+D4usqQOI1eyfISDVn0EpeyZDSagf3kk7PsvMz9Rw9oehTS8yfn42EXft
FSPFghEH8aBjw0W7P64PpM6B6tpCfiHzyQqvhLqAb/y/GH/2vS8zeFBIHEaWEI/re+G5xIkos24X
4o6wNNwTVY5dbdjVRQA+xoYN9WJlYA+pGxD1MY/hxPbXhrUGIEplitSKd3qAzX8gOSXMETqKJ+a4
l70s3lpnfEC190WNw9RqnMsO6kDD+1yTLvoJayhftdpY4BwvNM5DoUkwrq5ednC/3WPtOtehQvwf
zpuG3e32pc6cggdon++ZwO3wJHXUfs5yQGwVIxveUWgf20tYC8I0SC3gaOwZSOPAUJKnOGHQavT6
OJcaDTafiGdx0Fn+amZRhG9gyasYlp5sPUE3WSmYqJ+vWyxzfn/B2FoSHfGSmkOJyvOy2KylFDbt
Q6E7rcazocm7AoR9zSk7xqHzN9vqG7HS4E37Yv0LxZ/whCsJ+1AagS7dnZ3XRD+1P+rv4o7Uokl4
nuUg0SypCz06BtXuv5TclMNQ8aBhVBHvvthzYQTUl4u6nciWCYLzcFiLa6oYXjHoZuV25W2yQvbh
ZbTVOUXzOjtRuVBFF4XYLoyTvm+nO74CJ+2KRa/XT4hjWHM+uuoSqn5hytmRixP/ltRP4NEVJuPZ
YR8X1tMK3IZTyucq7ghv6/t8ppdu4cG6yPuBIF4hTEeS0T4QpCRAw5pB4ACK5Exce53MC/QR3ZLp
S3tcIvMaQR2z1E2rDGyYHYkwtpADekgYAuQTQJK6mlq+m0fZteMgohudDgeXUnUbey2m4j30Zo5k
zVyCHPUYoTnabxbfyc3M3f2RkC5PUbMylofFnKsKnUJjZTUtdaBpkqDhxizlEOfVTd/6ijWjNhM1
PTj3GTxFWidyyhmRlnI4jmpmyFfHhqXO4S/4ELZjrDnSeYUjIxTVqeI5zfT2g9uyNC79cPe+BYUN
UhK00EiTGaztzmV0aCQ9CWBl53p1+BqIr7KNBZbUOG6dBo0bCAE36YJQD6/GS1UUQgY0IZa0ucQV
SV8Sl0c3OVE4jMx97nJRIPKHbYFQH4Btl8nAdFHSVpx27Tub9e20dAXzk3v4AeWt+gI6VBxD6v10
iEysqLkHQB9NyGhvO4K2suDeEossO3Mva3P2Cx6LnFla4Ggni9ow7JYnCFNPGrD6c9hv+vy9BISn
Nn2A3ibyZnz7mhf+UwasJ6Rbbe6j9NKo3fvRsseGEsiutxlICLwa0lYANKm79HcewvGXPm6RHaZj
7ic0FRy2xJ/5mQp/81wxtlazMI5s9IWAj7nsJ/4Xp/6R7mVSVcU9GVkkDqGs/GwOvOd/ajuXqhft
sOAM8hZHy327fubYrvBC4ftYKjI9a+yuyxKARdbU3UfTKxr9bH2pZGkSikdyBvtC4NayWH0qvGU+
gcyAsqG+SfstPfGNT/66zJlO7zot9kh2s8ivjwxWpnDCYK8IctBSq3Cd8bBLaENCaPUSanoMf8Cc
onbCPtDRtdRzliDTR4QITqPhoMOWLPeNiHJKkLjQFdztiOkE1oZFwcmymBA7wt9IEneb4+V7VKf0
F9nQ8crMoGDCTVcx2vfY+m2qOm4QBNKDg7ld8y0Dn4M5EZXNn5refeIzYRSwYwlMev759SKj3iMq
uE7TUzG0z8iQAZ1b1vjZqas2LcbIPKlxvVGg9NT0sHFdwMDWbV5ad7pIq3pBAOPNts3tm7OSHy4Y
RSxMKeCj3TKI7zVuYiaEiiJCq/Z3axmEohYEs++lbKHC7LrK25eSZ6ZFZmabaqxO0ZY4mnnQCJel
PUYUFPDt0xZIkFPb7L+7QDA3xNRRH22+TCgap7BDGSFfgPg1jrOma4icbn615J5Co4cpBSS5iiAU
U0GB+1sTPTuFqVN11t+KQVefQR6WfBCMNtaUL6IpeWNeA4cosRnLZsl6RneV2bX+edofCQ5Mb9Qf
P3VZzQx2auXU7r7nvhNdYelveOcUL6589wiSPyhGZW0A9gPsHpOmQug4bD+MJToIZlwykjsosOgv
SNIoX4hZFF+5r59VTbqJhzrJ9fPVumtZ8lMnX3xdUW1cq66UBfFGZkOtVQ0nNbCm7gg8LUELAmtv
mv9Or/osmNy2tAUwTZ19UGwf2xXXEGcqsGPqgWjZ7n0J9/8xhm5WbB+e2YVc0BDQ7uIHKuXNUzXh
lAPkpl0jLUei0MvDFG329fIONPUmRQqCNGEC4NoUzZk8EWVWsg+p6fn/I98UNSukx3KSEvZNeraR
1XBKYnd6cK4EbpIeiHSX++u+M2warouD7z6N3+RPBk98dcVElTOvEzmGu07elqtyCHf/h/MqedSb
BWo0coDcci7H5CwpuU5uhvuNM7NDC+4YppkimWM4jkcr11eYX/clkpw62R8NlC/P0lHEh1ak4+U8
/XEaTPdcUelBvMnGVhYyUojYRVHDmvlS2Kr5IuQIpHCzPRBkGyJ90r+5YuqICpHxwYGpbsX7kjIG
+afVdaQ+y2I0RffqgYDfYsc+PeCOE0CtK1QHtmu2YuX61L5omlV9bKiHUo0JPVg9vQh8ArLzvHxg
HGMg5t7j/s3tw3d7owjuZb3vELSvhWRwVn1tK89hUmYd7yooMoBjvFM8A+ywq0jOcDltIqV2kf6v
wL8l/Quun8pgRhQfax4EhJbk7XSatxvQ2JkjeBWHBB20lHvmqkGQAUSPyAsqn6Q4IUKMyn+H3dsP
O8IY0vHOfL1lI1OosAuCATF25bKga0VZOGE6rypM8ODuBmGW6BCkCEaY4l/Wvxu3pjsL78PFhngd
QoQb3AUa8B0sE8Uj5oMQTFQsXN5OyVTcYYVeKY64K4nC2EFRgwIkNWmfESxEw3v9hISU0Oorea42
cq5B4kfiJRZpPuviWU2Dh6x2KqlOONXzC5zCOOxQkteDlF8IJgRHpGMtUV6qf4cpq+1jBo/QVscE
ZqMIKn/A8QItzNtwhj+jUFReCipIzG5WpwZJqrCc8NX8asXMpz9wP3aKS1JM5sBz2GD6Xs4+u/+H
9NtOvm5dLd2J8o23USk11RnkiYE37KjBunxbcTyaRxt4Zm0mGOMFKHEtmje30NlSxitFnnF9OaHt
X+CJ4h3MjV8m7hfdMq49DUYlvKD7fufRuvl1LIOjXBrNwgaupeb0BYIYVyUXaIZFQsn2ORXXDvIO
U7+XFedy/NfU9HolPx96KQZ0TCh9j6VpxugFIJNiV4z8klbhVNZ5FFDWiMmi5ESZfDVadcnJI2fL
C63XrEKWXrAv9JsdlNYE5KqRKdLnUK4IybjWW/wAlyRTLZf4kBsiSDbiWv24yQft9p2Kx2Ae6lhq
jgmLbGDDzqaCgagRXCx7JOrsp/4i0+JBC59bvapzBAdxkt6m4ZSHsQ26c7JJM2WMSarkjdaEVxhE
ikQlqkKk8v5bjqO2/LcRgGvMG4t7t/zOLREdMdUx4knBFFPomZZzyjhavO655VdrRFZBlFGidXN4
KkPQ8lurulErHdJvgLIM20TvXq8l2qBXkAOagyMzblj7d2kANRjjfYdK0++yy7zBH9N1Fj14Ue1y
uCOe+8RFR0ZH7mVvwY+2bhbnDaFK9JzQvFBcq+yi1RvlyeKEPe6vE5V2Ma/ORlWKtt5I6pa5CObC
Y9ccKKyGeejDllLIA7NBqgP4VC+Y6IgQFViIf4Wn22itWrXSA/y5x8BI5vOqbHI9yX2W0zJaNFEp
92Y3Sq3LqhMExXaORhiTmX08zqHXte5+RcY+259WReOUKhyMQhkElL6ueVyWgyx4L+zt/5I1uXli
izTSC9wncyqpIXYxUZnuQ6pdy8jxRDGSPiECWYW5srRkoV7cyDpZNcj1c1c6gysTz2AxRnTB3Wtl
taEBjYSoW1FBzKY9kzIybWTuzUfDIDMDBZF5VLVT0xsU+73y3e6Zpx2aNAstvY5Ikykqlkc23IN5
0Y4osTlucPlhu/F+7Xu+2qdQK5wEOUNrhAJS9Og2b+SN7T4clajaI00X5eRyB8xXe4hZmX0vTvgV
XqQcQtVW9TCH8iBRj+xFTwZKLV+aBLlOw9DA695Fgbc1uuZZH3ZWTHU5xw7TuEvzRD9QE5BXIf+7
miEURBxjrUuKjGNbOvjCZfb2dMl5Rr9uC/Kmy4WrwkxNbtEsVTwPatHNbN05qLV+yXysv+d9ZsSh
IQHrNq8JJat7FFbRDYAmv24bhvMCdGpe0hGiPn0sGa4sDmPRJM7M1Xg7pDpXVJRkOXiZB90PMc20
tJfoqNHIodoSDXt0KIHgdN3t4SPtRpGOxoJ2utNB8koYsur3WCw/0ZVKosF5JG6O+axkOqdMJETp
tySHvlg2nA/NnRXrS7/qAP+BwSCnIrFy2zNhwKSveKSSs2Hc1WrKdOKHthm2QpLlMFbYSsUVamZY
6frim/QLhlXrSbHHe7i9m3aS1RbNyQsdFERIhhPLfgkwIi6YTEzcQk0+CfjzJ96GB8k1JUGyZYfH
qa1y4RrshAzrCc4EOYHZrBaZC+wPmcUJKZy3spe92X37SMIbT88hTLCAP5A8Mumz9DI+Xzx5ntoe
BzY9D7ZfsxTeQmX9sSU8tRI2tONB1Agd6AQKnirTS+XY6RksPrPxC3i/BaVVzPEDJmRjrgBb/mtj
nMOlq5BdFi2QoM7IRxaPrq1fgDhh7eerdowRHsBV2l5/w225qhcI+tzrllyhDBOmnghgldXnzOxj
QnwHQbcOfUQ7rKhs7fMs217j1ghQz5zKo3mMiroR3a6gWGEs/MM9VDmJFYI+0HqefCXCgLapvk05
0fvU27+blyZtsCkWwBEUjDKC8343X1+VcAYf+Zns94eoECpJrJpg70UOc2KPoaSh4/Dvt+dXaSjm
E94xxlQp6UPdcx0hxgncHDXT5efuXml5eQFElVf9EcI8x693aDg59w29gvbA4BQIKc3igL1goExq
MwnCFxgkCSGo4je7pnzBwA5r/xqmq1mU4nbwlFaCvCpHrLOmRIfRKmBv/iGH6ifJ4KD8zTpOSdzi
MKowYEy6McQ2Uu3eiPGgPSJDnFq6DjbtPi2ielORPHlnpWPAv+/0yfK8YzghDalTMkhkomOWZTy9
kV43JC45YFBGjYBt+df2yrqp57AOHgb5aJSApiWoVC2sjNGpRyfpcFpFZGprM0KxbTsvke/hsRv2
OQmKtvROueVnQH10Ce9u2eNZOl9+7xsJ6yelpHmqbNwOfztJWBPzStn+sqYnSA5kkWusn7xTjCw4
58fiwvM9tPsdJzaUR0kfNy/Wm09QJJ1WKDZ2ccXncfDMEX7yAwM80Ky3o0G12/cxu0OaUMVabfha
3pt1cvt39ig4s7khlcBOEBhy8MYF8XytcNiowzUgSa+aRq/o1djpEzLxjXZVZ29273+PLI5exNF9
H+AxZCKTUKnhATZgXPOwnyN35Atk8daXrZoPkThiKpf4oe82BiMhS5By5t5B+rih66xs3aV8twnF
KhAxmx7SSNcvnMxP37tpwUoZeBLco9zRDJlZlV+Zn8UeWHg0MBy+Sa7Hf6nejNTC54uv3ZvktTPM
5cPgjKBsF72fvdfMR4bJ1RdMPJeiOHpDd4ksKtNfRs75gKRnBehm42YC+xQPHhP9xc0v+wOFWrbC
036R7hIPTgz9+GPRVfLtJ2tpWAQu/C2L0HKomCY48R3FIK+35QktGG50Fp7XCBcagS8n2jljJkfz
PV7wccwZzUxycnBQXrCHorpsVnXZoH29igTWq2jiNtUqNhixLfE54I4SNeWYkgnpOnfRgnjGh+A6
+l0GbatiyyBYOKHKeziXGKZPANyAVxy5MHBQbyK1cd6K5gIyioi4/lV8ClmgzBbnRK5l4984kI+r
ZaUQegpdPQqWpJEiPkGBxZ9TJy9C+Jy5MWptBVwrD9wzEfOTdxhMzJV1JMtrBlEGRvy6eKDxew1W
84V6aVSXy6Q/hMVzubNXJTI/nTIH3X2nLTtmUwdv374VCectX6woE40Y+HJH7cBKkQJLzlcMd2/q
UbS9tMp1OEZ6itfBfh3RX+0ktwiGS/W++6oqoPeuUjvs63YnEAuo/BJ4O7kyRNy3XX2pyfRNA8eA
mC1xk4hw6qRSdghi/n+UfYxgz8pLw/C9INJUoLXzkWvUoUirOp/La32a8/P/hJkZT1gPgUiaUb9v
RgJ829E2JAAyPmax/yeRz8wyZnQvQwbLmeIOh/hCUkyJzbps+S3ys6rSdB2NvH4YBRqndxGUkDWc
djpQbQxJO9oEqXmwx/vWbrBSUavgv5kdV9OkRMySxEt1H/oAqrNQq33DYLzGaIcUC7YpyphFealx
5KEvl2mWU4K+e2kt6cAEi/P2eRjcIJgbPL9LmYJ59LY4Hv+t9rToKE2lwJlBT+/dtM0q9OC2rOz9
Yq0dzJ2oc8Z3gV9TVAD9CZxWi2F7BCyB6nes4u8eQ19XXlph/SPtes0HcxKZa0UASE0DEg5ztEFg
3aLEu4H9ahwcYvCt52U/xNwaDgXem3sZyOzsiEcvrAjrXarj9NzuxO+zDg4cVY7yoGUEjs/0Ultj
QledCvfV4rv+/7rLAfjvkNM4VpC2+y9eKuWJEM8lhsB7Ox2jNF+jcNKMXN2PN30BOunBgK1MVLuL
GeDbV0t376fQdklU8O8rx31nuTqUe/8E/V2taai2Vls89Rt30bFnJLAtGJptwnG3hD0hBS+XkZb9
CvrIs6btTum/De5Pprf/Oounru83poM8HJ31pHmk1Xo9aoBFhfh/JaGGTqGw6eIigZQhBmpQ73A6
fm53Bdc+V+h/qrQBtFwbWChwIgww26ybRKvPiPHXisM14iqz36fFMrFm46V8+Ahdix/Jr74q4Gqj
vB1WVru/+nb0QumROftudxDTb50Y3CODwSZOTkgEmOrrrW5x+B7aZ7NHdTXXLnPmKK0EWtWTp56o
ZsIbcBpm24amPZWS053suSplwJ2HUeQWcoCFBXJS2yPev3L9d5Z8jvp1gw2Alu122LY6p4ZShJjn
ihQQvN/LvLbfDewDKCSiJtwdhqim1q+lMQFj56vMlXp3weYd+wVH8LLKaPu45vZIAZJBKaonrrq1
6nFRArrDEfbNHl3p8P/ceQGmSW1+FBtMr4e37V2mWOT4C/gyym71EQfNy2gQP26OliV9WUuoA/Wv
+ZqoGLdGKaGQ4S7Sj7A9bh9bGsfH3UyJh9NMt1lnX24yXaquixcYCi/WQU7ziHK/FW2Up8YIrOoT
2Ny2gDgjz0Rx7lg7Kzzpb5o1cqa4o/XFEJFPywDSpYN8setiEw/YCvQQ4xNlaH9M+eiMN7v6ffAt
RS0Z8fa0f9ydlrX2tttGd8xKxaS/mOY6Y2dS7hEzpvpUMViUhKLKtwu0+B46IRkEb+lEDzNDTowV
UF+ca9mJjCzb1CTZB6s6Ujanqipy7VGJGauDBgIAO28CZ+RIJCYmdm26/cILjLgVY7VubvurRb4H
jBrY64YMrEE04rdd4nlCQValccAo4PttLu/FjYXCdT7xETJK61EPLQkURaMrKXpnaLJFYaHlMa6m
JGXAJyhGT/WJeN8srYRHOYEhRk/Nz+XyPNOmgZ1gn6+/V6y/NOa1W2zqX7yRfFnfIHtm4tiDgtAM
eUbFeK27aJ51Wz7UbXjhHIRXg1vEFE4GCO9UDQnAe6ZDDOYCeXut5WPJ2aKQi/zhKk6wrnxrwRvN
uLZv/Ey754q/LaCJo5h5ih2tKVRzp2GtdwT3ZQDOhnKw71yvStmrL2CHPVfImy9Bv8yge7RDe+Ia
Z3f5VNls14YA/g10NB/q4DlX1z17eD1YGxP0jATI0sM/k1N+eLfzniwZ1heTUTiDEAYSHUDwJOm5
Qzv09rgGhB5cvnsdIqvZriVsQb9B+k+lwfPs/Vzl7MsauG7bbyXs/MKTqeoe7KOP8RM7J9zpgDa2
I2J13MNFh+irrltzBG+nV0SmYnxshtBuke1ifLUkZoKb10dULCIjG9Xp/bBnjAzU0SPr/DeXlh+Y
hw/l6sJwPGfprFJQI3VJOaumGWm/ZaJkFKLrb9JPPfbnpMntb2wN2gWWEwLmSsqYY+LiEuiIDFSa
2hlZM3w8qDII2e6Zx6qsPd/JpxVr804tNGR76NmbY5LCXAtJ4MWwFd17m5KDMTLKBe4DYkqeXQOJ
YLCfV4xfBPUhOeBR2FRVsqiPcBTpJox679MQ5yInFGpET8T1BTKoa0+4HkYFAqsxh6mldhVLu9HE
nUmCtGnuB5dSI4DdEFEZlXkLke2EK7D/NPlj2uzlhkoPt+KXaZZyTar24c/+RcUpaHyo4NkKAkh5
5HKt0oXoLVCYqxbi6ZP7MqdrEsGcWLPDTzLfrSF0RkDBY1AGdKzjU2+7VuBEb3lig+AHTPJzyE2b
88EDxGTDkOR/4S+stOamQYdyo+zFx1h3lLDnjGMJqNw/CPdipw+SL4vhT3kmKhr4tRvfk+WhENEY
VyOHrsNbSFriDpJpZ7cx4YI5ZKI7kP7cQl6x0qCO9aiU1M8jCoqU9DIbk4rwr1h8FS532BbYVoec
lcwiSmR4hwa8d6gv3ZELzVDm19dNdyMgr4AyVW4PO1xpHlkyqH37SzNZyeZdkv+2RDBEsJ9yPTN/
7l7j+7q2D1EAFfCWherEWAs6g6QbWRrhqAYGCY/F7avdnb9zE1n7OKBRApYHyuxHQdNSd8/Y3QnO
eR9ZvxVWB4lADfyr1RewfO3HW88OBiyHPmSOpdhUoLV5WvAUpOFqvvaMnEsjEZoBtmTbwddkrzZp
MThBTyjJhP2DGElnAcpUM9cFOfftSZeCm7vidVMEuU+ua8oatZNZAkLmW4ORPonIslQfnHR9AjgM
GVL2UEBo21NuE6hNtFXLwfkCnA69vlWTOxwLd2b9PnJWN8mTF2PzrZyIGjl9qF7RdCxQpTqLbJN+
sYqRaghbJ3vExX9D8ajzrmOT1BuY5Dm8Cq3GMd6pwt7HlKwxUeru5bLH3CT3uIDeyhdIaKwl5Q8U
ctLQGqpiqt9sARswUdNCiK6jwcRWK7r2EIkly/X06bdErigAxjScT12ca21WEmbjVjJ0CJ1sKebj
sjS8MZwuGvO017oAGTARQhwcC6oZ/J40caXCFlc/1yOThTnJKKKZTH2dFFr7vvOI+dk439y8dlZh
Bb0v33wN/HN2QM7bN964WGB3jsnq/y3UzHr0F6nxSITfxCSp37rj0e2eNmQXYdvGMEiUvHZ7nS93
hV+5+H/seEsXPj9NuzZbgKtYiRlfeT3MMZGf6TErKNt9Lzt0rb9VirJdMI9h6jQirUDl/gcr6FKe
SJ4uKPOynQtkvjYqcVlmjErO3cfnSu7eaGRY3LsZ+O6xXaW7ZS1t5gttxwNZVDSfNDhM1U07LZ9z
xUtOzNhTiNlzhCiGEZhBZHdGjxE0rCSIhoMe3dVBZ2rLXq1HF/O+HyXnaL8r8MqTxn7/WcsWdf3Z
vTAvpDduvBCBahHqJaRxteEQUq4gK6JKH41jvkAqjbC9ChRoZ1HmmJPfmtM3vYp210RXc8vJLgm9
52t3maC5a5lQ9PwOXPGTb9me54vgFDSAkwVLcRChJNwFLSjHle+0F+0PMiL11Lr4THf60GDevqP4
yEhaR5IvyVnHMZG649KRFvxSeY9bTJfuLoh6clRFDoj+eMxjpbGYdhAtL5XfDEizXDG7vmEajjP/
pJiR8QRhlzc6kP+EDr+ooQ3Tj0QPph7BPSC1kwQGCmIyrbsMX7JYQBaSia8YIiCbZBS+EZpCDngM
uiIDorUj8qSwf5TJuLFB+pqP+ewelIqP6xusc+vfl0COOxh6DvBMmR8tYBfDT4/cO9/n5Gxl6jMa
YM2sZXqbJDYWthk5MABCw+ol2TjK5LVtgdlUlDwdLGfGBQnthbDjvykDqZUnGbV3QG8GxtGKP5oV
r/CEka4nBPi3eEjkoyLn0tEIG2Q1C7B6ugdrfEzZVIVYiaE2W88u0XvGadYXQiAsWgXDjAKCBtEj
v1aGwlqWYdbquipY+tS3Iuz+1ZcEUHUxndgrlXnfGP7001pruELIWeBAb50E0eLfsueapmAi3mNQ
DlA5CoPSxIePAr6US0xy7eMv5Ibmf+rO8tAiahUduVIjDURIkGIksv3VWaz5IZe2C+B7PXIZ76Xb
l9u6GJ7Mka8kD4UjUrLVwW02fYrydyGpY4zxWMg3fawrmA+tV90DAiqBuLLzmtVxEeYEVR45OIFO
sGlrmODEV7TwtBHWRYQY5xIh6FSye8aZLGrcjyXE+Eg3QVJyRoDnE3OvZqm61FQ+zIud9+FSJ4Nh
RcABsNC7EubVvSk3GQpMRfi03F1fbEUvO8tEnGbbepDSSClMAYpq0SlpFfgw1NcyCYpW1AxB5tFr
QXV0dDdqSJBK/vbmQV6ySzHfUwHtOS2SsyBt3iwZQGJJQE64ohRCV8U97waa4RY0B654wDXKObcB
jvN19ZozQIqN/dNOzTB8MU+E+M/tuwf5yY2FFEYfgZL3dYUnJZ2UPE3HMWiCwQjGOm2wZbz3DWlN
h089cI9CQqJ+b7fNckDSOW2gSlQEM3ZwP+lbt6XuMnlIvPjYUW/hpJv8s0F/AmRIhCPPW6VoYtqM
N6hJ/Qqs+uXLEwPCP9yqAuLRJEmhzdXZ4C4xLTUfJEl4k6fUzpGWlvbwDyqlfp4BnWgjWuub1yCW
4VSW+5+EvJCVG1FmivVg7r5rmWQ6HK9/Iqoqmot5gkdAs6nb10Z01hkjNvruwAeBWFLecR8RGIcB
8LDT6ASr8ruIA1b+iFUdJxMLTHQw4tURO7+cHLDyra/l3Vh9YDalpuGlJQrT5LPKq80+gAFEQDLF
2or1MIr1AsQeJ+MC1FhTc3SQ7rzogR7spZsFX/JrUeRS24ZVhkqJWohPI8pnEtLFLbevcQnVuRIG
Pwuj042nj0VRxd9V46NSTo/401djlfCJjwvY0ME0S5pr/jbboSeZIHh6GJU8sgFhnV45LLcqKK0t
S2wHSlVle96UxGVY7K3eJyndUxbWjIIEiVatkodi1dwD8uvt1eXKDRAw6TU44rwJgJ9WcT5CPMYM
0mU8E+AAyheVPwZH0rSBkIJHCxHgf9qhBATIBnG8c3DOyQBqmVPcWVH22ibffAG19jVa7I6BFmKG
4g1UrcG1BmpRf/7NMeYSWDjTSzaSnk67rcxZzwIuqCl/Dph8anyiolVBxRyjRNtE+DpEJ7elkrt2
o2m/WwJ4xRSCozgPpIWfTJGebCMNPOMSwdxhvX3rQt2w3WCf0oIVUghBF2/1kGFdRkkf2/FL/AvV
qwV6DylxUQPWBAEgEPW+LXgR/VuQ32rmFDEcC3k00loYIFxVfocuPQ8BGXx7akGTUQ6VZ5jCiqpP
QbuSHBPyJXqQStBeUWj78MmVhSN3zYcTl7jWvNz+9t7XBhVsKRJnIbDRiz4D9eLekPO107/sMzzA
r/e13UEeifqttTfhaC8q2EJmMUTsHcNN+BfTjrRvZeiKJELD3P+tIcxYj6nM9Poev1yHt0+fwUmb
HlXfHYpl7K8wwZ2BLB0oyzZIPfjaSUl4vRFO9mmqgAlGv65ce+0fPQ7XTyFbaYbFZ64kUuFW3uqR
zHfsxbL/W4C2uKoYjDlSdJClZ9sZw+NfgZGK7+8Hc9cwl6ygtAdffHIKMt86tpYH0ZTOtsLSb0uL
dNlqUH2amUknoX0x2ivNwAC5KBGKxdCMpn0GfgDP0Suhb/uZE0MRp7onzyvtJt9uUpifK9qMVkxI
QTfwLziAKNRRf1FAI6KsrHs0/gmAZ7iTTxYI4Q7KYWCZehaALwgLhRZYtnakTyFrt++3VSfcjqOe
DBJC/FYlkYpc6PqOTzLXk5JAmRWyz5y5isYR4MhTetounxXht8asqUHlorEMT2TI9DBpTnc079l0
SXsgJ4Tw20a1Je8idOQ/jC1Vy8vnzZ20+cP6BPpm1WoohueSzgu3Is672ppzOsKcKrF8ukh33pox
UDJNOcgdhN8A5Gtiw4Z7zIfUnP/+Quqf0wAtaRhEj+6NsyF4cuW4kA9lCKD/hDQJwjwghyMeEQig
s3zDyLqCCihxgc2mKoRjameJyHJzq3p16LRVJ+iSl+GYglZAERR3CwnUnKgtgrKDIrKsN6+6q2FX
BiDpefn6gdSCngZc+eOJ3OmmxEF/SmLrS92I/CpcpF6T2VW26q8bHGWCtEObuohpmM0b2cx+JnDb
SSIccbW5gbfs/xrOTnn8pPoW0GxWh/uxCM4C+QlsA6kZyQJvKreRtWrf5QB1P3RPR70fJrN5C89B
RObPLdg/yMNsXGxQHVRf0/Buetfd3tVV8eg1wZ+cUOmQEkd0KRHJoz1cfo/NFMlpmnouT8kbnTrd
dveDqn/yCzjsXL4qXwzUMsJ4uUOyFx9fiiigCppcHo7Kp9mL2z2QDZ5nkhR632gE+5BwnqOml0p9
dRpafC1dP5ypKMrM/dbm6H7O39U6GYMWyqN5oJa8SFoun85fcL8psDRu6CRk5/uPZO0DVZI0/fq+
3abs8lxEZTGUGYqW0XnTrIv0YCcIFefZJTnDtw6ei7bVVoT3dkcq84glMyipNweD2jhMWATDu+3T
lcPie5KRYUGscDy80rDbi5RbBVqiFhh44bSLKBgB70z06bL3G0620sz7MjtLhHWwMIVVXjGqPp5U
uOY8m5ESZcg4lCwlmHMp1j6SxS3qhjfHtFVbRjQUpuFkU8ApVwOMPxxvi3OYnxsBx79GIoXLGRnb
e+1EororWKyKBJGruGl3DkPlRNk9KNbrI0ACheRhUnwKyfaRdNlj9dDDJEVRYPrQIhaPwcL4NBxh
fpuLSkbBhJujQsjPrC+4ZqTGlmlHBbAEEnd6gPAFvADIJEAyAIvWi4LMgmi6md4BEfpjVBhh2/8u
FRqATrCVZ2y7wDlcbfkQ8ptWFMzoMb6nCz5tgOBJSSJAukeROKiHvZ70ch2DLYJOM1LQMKoopp7L
CutEWYTs5xYRCAI+OBs9wuCyi29evcqqTcm4o38qIFb5ZwDLh3zkCB5aKpX+78sVpXiegH8da7aR
NI1ZU0iiaoaKo/B9mX4Z1UqxuL+AdgNARHAEx2qMfVgrFW5hZTBo7pNUUpdNIsY/HZ1s4TtVmPM2
0j460vZiv8Rwy2aOVoY00AnvAdRYSCXU0hinMqakWNWfdlt6ac1Z/Ko3SX/RzT7bClAHDBtDPZP0
ahelHJLq1nudiZVj1yZspWaHcbi9evYDJIIVBiD4c/I67DLIPVupgN+9UtWNsEZP39UUrVB7HOsz
/iZl3wvAxOz5LDXJ51t/CjBkvo4qKl9dLl7+YLjY46Sl5GvH+NC47uCGIQO2ElUED53iFS8P2a65
B5iRyY8m17js1Hcdz7hx9i6U/jIHjRYkKrCShF2zuwdTpU46Gm4wBFpCoRDG7ya2OEfLlEsy9LyC
5lGMnkpCB7T42ECeQqORI6qJTY/4XXySCU+dqS17/5cyzz8h8s/jVm1cGA5QXcO9N8EYOrhhbSu2
vxns5+bSldbuUNUYKaK1sMS3HkcNOPcPen2VCSXHHDbVKJ7zZMaliTUr1aGCFn10nKSkkCoS+Z5p
eaFbVMDr5XT9gVce9bgmKZ7v8CjvcGYGF4q6hDGuTBtCIq07JRR4e5kGVoI7dZ8Ts2fpPkecXpc/
n7/SwXQ+TFWcS/pbjM/8PQKM4FCksLPryjfR6JjrdpasX9ULictzQf+sefoPKMVMwWju/qquUdbc
MD5xIPumnQlGI8JFFzpwCcG3BrWiWQq8H9GXf4Kh3ppxLnXCU6ORB1cSO8runUQNw1t4fJCN1lVG
mOVsJWC7/KLB+gXn1xK2tqmD2fAxUqztqz0jy3Zsw6nKR4jgqd9yOOqP+nlZwux1/EsT95fXjQ7T
97SopxUc3PH1D32cj/dc49mWP8tMr7934KUP4J0vlk83+i8qTs0gK3VNnDzE5x5xcSkHu4zc8i+e
0eFmX6WYiNAO15dlm4i3ojfelQo7PwCLQMAd68qpLBy6VWMPdP0eqbFobTrI0onV0doYsezuhr49
j7YwdZbNJCInoTPl9YcPFWEfw5kzfnO6pkCF1IDPE3QoyKlwfWi2CfWO0fTUD+KrbQuNkKqBb8j4
/a0eaY0AjWiAGmpFDDM2WbOqa25yiQ0uc0TFlcAHTzFe/W0EB/NFcq3vWn+R8Y0Wcl4CRzJLRa3k
b3lZvlVqZCyL9ZUPlOAhCiK6iCo8W6vXKk7++kzZMX/YjlPjo38dexPO2lomzO4sskBoNvYyRBwC
l4PkxwFEHKr2NtXKPiBTFKM0ngjfjv+4gEyU79NlRla/M+Of+iKuhPvHa6dQUqFTJQqjrCUs/SoA
YIcHbjGPMKInrmbsKQOaL3SWjwnuh5DI5OYP4sRaGvNrxo7/XKffXpj+AuNjmOKNr0jI1LNGQVEf
HEw7eAFGA1i/lKAtJ+4lay9cw1nbYLxayXumRT37J+u+JD7R8Bc6h9RlGk2JS4A680WOv5Hf0y85
yl61ci9+xnVuR5PV5+el9zWrhQge3j0gF79Kx00Wi4kwCIhOFvIuWsFPqEa8hweIjvaMKh+54jUT
xPWnfE/QCa8FVEvvmyqEFy/B3Yv9ceRwEMU0AcdZRwAysztk0UveHlUf1ljPA/Fvtz57kfNECwXn
YLsoC6o5MT0pN6UpL0NncRcUt61myBfo30T7NZAxj1lc4JCZtXy50kFc0U+BCV4dZ7IZmZoHCJ4G
Y47to92AEHEmHAtALutiTPgq8YK2bp+M6i7XQsyNuiJaptKLH1d8ZWDoZaUkP17U3KFZVJpGBpeZ
VG7JZpSFHXO+DVozJez8zJK+gnriavvaYXtSJKuJmWmu62ZA8/3Ck8MS7qK8pzs0W8opfjdo9Lgx
7L1HXtT4+8fv+5lCNkVAOBPOMIu0L0pP5JcoL6W1vxJRfVo0f47GIbnd/fs7JJdmvyDelg7x1KId
qbYLVLe4QiZP0EVHEPD8jdPy7Q/i3ZelF1+HOlFoGRR8xLAnyauS4rPayfs3aSuaBPn/lDcNx4Vk
MjtoxJ4YMmVUc4OyQH1wjL8gJWQl1qLuVmuS9mNkEogdvUeiTKJckLSLMKfKeMxqd809m0JCQ+22
QM9y+SDGlD3Tg7ALkViISHiP5T65DAw/KZeGQ7azx9UnUFK5w7mjqcq/AAzC3QHXZrraxseYBm23
tkl6GRMJArg+hv93QJO/tB3PBA8uVwZKbEco8tjYGdMRrH5O+Rdy1XA5JHrt0z+43FPtXZLiVRF0
KImknA9bZCPm6Y6W5EE0EYkR2Uduud4U1szRlYUalc13NocRMxIdioz5eqWD54nzxE+sw2SJ0Z9U
0CbWH70Lk43DO59ndkarVhXlv5aJLOodQFsOX6sa8cfbRUFu35Mdqt3plBSyuTG+b1WA5IUDoy3E
CRdfvioHwIs1TsjEtAL3EvKifZx1Iv8N1F4SmTMjoIlNcZyDvE4gIFG44n8Cr43J3nqyC/4rzu/F
tpZWwbIufhpfgucZrUsAEb7unIbxZjaxDcZZeKst/05PyeexnqL0DcWvd27wKstRqCQU7h/a4FKg
bMUjm+z4xqXOk6UesXkWHnmnZB8pnFKzEvVdIN/KEN5/1Zuph1oRY9bGne6Wte4do6FY8WnKUdAc
jZj3W3TDFRdEEpw/QXCIQ/J8NFPumDOUEf/H5Ie2CWE6e6qDDZfT673OF9GkyQMBIEX8mOeetQ9x
WHt5e6iaPzFvxuloGs20Bd5Mas93uY8FpbxRSNFpAW+hiNV+htCaLZ7VrIGNJjtkp3a85mSl141c
SMFlAY/YVqxe7EHqRoFSt9XbHVpQQv9KCgHHd1vRiQIbjuGqPWIys6k3VXEVONP8SwmRa1y7/UNH
oSnUlXUJYGMUCvH8W62w2wxwHFYxWxGk05JYLoRhh8SCGK99Nu0eqyh5WVUOhZCGRrExHS0dvunV
ycUrHvmcL6wJ+JJBgjulS4knHia511mpWpwsqE/yxHPZ2i2ARoWgJEliwQ02Lb26/4+ZyRFki7m8
7iD36+wmBIxXUuklWUA5Zu2o/xCTF+zWsNLaICsCKk6lPUTi9aGNUaNMIEcR22QlYkDm4CyYeWxD
WBTRpwF4DIYJ5XLr9nigJyanFI0SoIud6LUlmyr3UFDRRuZxUZjVY2O3cPJnfBsVc3Nj0EhLNaXZ
6fhBn0jdhbwmfhBpk2P8iC0QIaTDNeyDDGQwVviE7J5uwD7RHJuC1IyiPk6U7hn2d8hMjlUyQxX2
t/G90KKIk9J4r1Fi7pX6NVylVpdAuvWf7G9/kF8s98x1/Lsjgzo0tVpTB8e/2gD2VKswnCgeHQgX
pLclSBYzi3bVYXNUNG+WkImE51FNc+uULGPzeuUdCJ0bUYHLfYsD7Kxh6H6VnDk1QUGJ9+T5KsRp
sPcLs1XOldNJS2KSkAW9VLhRELaWj32UZPHR9PP0o4GN7omzWJ7b8ZVDTkqsDEqMAZM05wIqfbX8
Hb6ZXQhnCsG5vMSSoaQaL09z2Yh293DZUShjVGvtDTB3fbz7ri6QhYGDd0KWjrfNAiW4fZq3Fk/i
gp8Prc/H8jXKwpsrmJA3duDYYWRLvczq/tx4y2s53p5Lze56UYjNJ6/8L+M7YJV7l6NQhN8mywlg
aeMsQ2RypVDDPdJnm7QdIbAqQLT1DRF4KrD5js1pSrgwenfj/0S6+32aqu3eSvcFB1BwRLDMJuzv
3gKO2+fVeLLYxKGMyYsqL/YtNnUHyuIj7BQKx/87hRdwxPX79cOOLuc+kLzuir+0a82XVgqAGOeP
OCDLEZ5xZYhAno20BBxPthl7FnM0BuZdkTIK4Or0cH1nGEYKHmlvJFCFPJ5NIgZq3e41r93EGmji
K3NEdEVxnOez7LHqQ4L39A3RtKBq0/zaofdbWHElrOwTSi/K+VicCTJahFHw6gnrAv4ywOx7r+MT
eOmxDogEFG/YOlkV5y/I3pSlY63//5e88dJrYwo8KNOJO7hMz3wswERnA0aS93nfGSc3wkpmA/tC
pLwpvrWLT9XMcCgB0d2F4DUH5kL/uNdnyQlV/Htw39+87+yfyQziMGsvTRpJkp32YNGVq0swRRpf
W6LLCsUTtKG7cIV/6SMKXFWbOGTzrITfegtESIjhWHbfXFfmyUJWI7Uy8tCaEQ9KZeXwwa/bUkap
YFpSSSiA3BrnJMnWww6CMXtH9FGjl68lpX9CPBe36nUXnHiR+rIwDL9Sagv9RJoP8sUu/0nmj9qU
CvFG/JYEVp4k4OVeirL/fDk79QSy53qZESbl9T8OfbwQQcUnCUrMmg9J5cCKFlHr+mHgeh9IEF5z
gG3ZyVk4HYNRGfIzbDYGcu7xtN6Kxs6lTtXZnfQ+NIVJH5/Ui2KYAc+qKRqptR8j5CtrhExKYk7N
O1nR9qlc7svVyMcymwQOl64ENMDFoZ9xvaJJi/LMJBj+rPte6o2wcFES5FROrq+eTvvTal9nSUR9
dHTkHxk9jerJqsaOzpNbsCFhGH7EWEU+5U1l0IDR3W+Pw7U3ncuzF+P3NV0ed2asFFDMcfdYTkPW
rsyXXEXNSQXIPzhX2riBjylYWZc7fs/dlfKlcyo2Tw5HI1VldaDFvJJLZBdFmPAMNEeUs+k1GArj
oVgTsNBtxL8VLxW5Pt0M2Awe9D4VcGRaMPzII2lgZCzS8Kjf1odArMMWwYTnDzwFqs4XjniqNKUK
bRbJk5L94BvhlRkka+hu0/dkPE/dMX0ff2WqrrWGWEiDY+DPXSf0M0RxF9Hyi7snZHF5+jv3wpls
ROMiGr4CrFukw3s4M8Gla9Gniet/pPWR4rVXFeEIPWflm9V0jyBqOjTA5YX163E/tl1MGYhD1P7+
u165cGesNW4YyObpO84YRhJnKIQyhbBhT8Qpa2HRzbQtTIu5Uxz9E75mW89QlBcZvddl9LkEvgcB
kTyGdR1BrYvc8OCVMM1oKHTRNvOQjj7cJDOIFcRz1AzeFJHgW7hPakrzXaUfy6zzvzU407BFrKhX
zzhS6kH9MsV9VsKGUTAsQsKoYscw6XLy3M5u7tQlVNyw2kuebk7vBCbxMsZ3h7o8ImHUOqxloky4
I7A8NfNIaD/z2fzHTuKA45GI4AFsn6SyrnV3KEY5oUW2itwIO4Nc6URGeZK9FU9w2F/lMW58PYmz
9zuXSoKB2lC6anTJOWWymvLx1R/szkN0fFUgHys4H5xQEUdKmoHtUxMl0DqG9pNJinqYxMUmfPuM
mSJp9x6WFL5OMFWFTG2KJhcfzTh5drn8egvnyco75glLnisTNcHdPL8s2BuW++cSjVD3yTX4wqAU
2sAdkU+ilLsHfXXIz48cYxL/XWH/jOTHrsTyfP7/I0jmWb6ls9Y2MCk37aYhB3TtZz7yFOfQ1BUu
xFwpJXHrtjO4zJFwTntADvUz+xeJSlvZYPbQQRAIy5wOgAFXapclKo0ciVSaZqMgKh/oayt+ThUJ
ndHj52wCxd8wQhuNAFqKh0IqVylftj4tWOHyO4pWLjtvdY6S95HlHQp8LnWA3B6BXibpUIGV9xs3
ts1EwdV21eFftJdcerjhEITx1/EYekoE3hfa88yaYs9S4le91Wv3qfYOkOmcjZpV5JNeTK7b6S6a
Tm1ewApu2oflNkD83Z3/uIDz/a7qxrTUfdE8f7BVPidK93DCZqYCKZHXgpEZBq3xPTsvPYSZ+nsV
7OB0ljJ0h1LjXB50ciLsD2B6eSaHfeIT4cLPwbg0A5Xb1YNZBh8KAC5DTTMrWOplayQLgHSGP69h
VM13KtLk/OvR+nmt18B+CMSigWKsZVfd8KA1AZk8fbSr4pEfUlRbZdHHMOxW9GTQTytTVIcMHzjr
kNqymmS3tp/F1yq0yqBw5kpUuD70Zm2fILpDbujDdJEIVZhonIOkJCLZ9QYn2cCODxeUi83IWJDv
OKh0092ayD7pVlztqocHOjYRMbYnOfdyUow634E/+eFNrLBphKDfKTHE87BEpPd6q/F2LFZbX9vv
X+4FLss7qfIOAkxzNwXxCIwXlShzJwYCLr1WUvriJZIJeZftgaKK+X4XTCBQ7bKHY92+QrxqRaZP
iUvgRwx440nKxmqmgdKlTp0ZfiYExnRNRj6YAV3DLojbc5pAzptJJ8A3zZ/opWcks8emhANDkozD
7sDOBIhW/ywsuqrDtdsbC1wC6KGmPhVEYDYuAwEHucEsL6mq9fMGpageWI4BJloEjyvL1fPXKtcV
MGv25MLeFlGAElvo8MuNad7OVGv7UfeASlWWtO7D+7a5WYWa1P2dWjXLm7tAx5z2O+Rr1QP3Nns0
crHxN95gukqoEZZkitEvlVri6OaRZPI617cS2m/k7rAKUF002I6hC9htNj5B1e4HG83R+csFUONr
H3Ab1fMrMETMuZdzowwdqS4wW+1dOnDV0FLQVL4DPzHn3ieAXxTSNyQ47RTCh9merN2GQRVgeHr7
bi0ebCjoTfBmdN2jGemh71Ie7O9kfmGEO1Y4EKD/U8pEZzu2xZJ/Elr69iT9XiJ2bWEtcAQeJR/T
MvqcO6NpNHFPNHAIQ7NoYX/Pp5M6aX5TiJzCBcsqf371R+LaWDXf/dLepmTnmUlEs2bkWrhoqBiO
cdk+721Y9azB/y1gwj6lVPoyWFnmgnZe+wF1eqFSwR4EBHf6siitcP7u1yxR49MA1MF02IwzDpRC
882VUw0AtompmVWJpHTAeCDAhDMmYe8VJn5sGMUsxj1j7le2IrOqaMTsF4AgHnU2bZFHELWKHG+g
p2SCbDVkGZ2x3egCwK/h2KzhNKiK3SJa9enhR5VQaECMCHB3d/s8H0XnuBuE3NqP6863Y1bqQp2Z
Cz1uyB/nDYEgIdtCqnN6uds8bjsStsjqDmz8C3cRqNGn1QYzselCWdMk3sHrUP+QsTvAluyhijjx
N7v8/V3BaYCitaN4IP1Z2ZEYkVPdMrNJZaMOb9EFArsybrKmXpuHy+qoWtPJKdz0RUekTEsoq7WS
Jmg8ZYr9ABJf6+fY0vBy3dFsPZo6Exfv7xS2VtcdrRz2p9d8Y2UabZ8TeKAlmXEi/M1PZivo0+8t
N2DLqv5UraefZfUv/8HwwllEPLHV4uHo6DnQYLEzvjZFvyrl7Pxm2tyyWdfQc43ufAmxx52VpXBS
KmqQZpPrwhhyF9Ik5J3zVQe3k1k+abyuxHfJQn/LWnque1dNxgPEXOEeQxPxEOPCq3bNk23rL7oH
kXQ/kajM0Lt4roGWieAV3SC88KLK2mQci1X3Bd782zGhzMSj/OoAPiGP/yaKK6OrVzUn3fsIjj01
7rkIq/a6zW5wD/wd3Uf2AWs42T+FAlRKATb8SCPZiy1mV/zXWKZCrOQOQ+xFbwC+PVk2SzABzCoz
S95H/mPsK5gJjqi6uRdHeGFL3ds2ZFHiNsCxL8s8qD57CM5os0s9Bfl4K+g7vMvvIme69XqB6P5B
/PED3zQvYrFZkCIJxA8V5/EqGyeAxVzy7PqnciUE8gCZV2YcxzhS4QEGoXTE11KrEqZ89VACLEvS
S7csufZaTiYB1l0YUFHWReYClVV+8XMPE/oHWbwvUYLgTYNfUpJH2RdM3EvXUpJi62pCLUdXnPe0
OhoJC2D/Kdrb0Txe/s3ug3aMso5xKzS/3z5eyxVT6NWs+8CJzaa8eigp7S/Ouriv8Clyv7H/pZrH
gSsB2XAEhXAG2H/jTeld1pkYVjA1Y2Qndez6+WBbumIB1/566KPFBs4ktpNtpz6fEPOIC31qabcn
jM9zYzUs7JZfeq3/hAM3bpSO2KgjCu3ZVaconB5NnQDowEmYPEPnYeVUFmq7E3CN7PlGd8c1KXOk
amNp50Bl1vtr9Mxd3SyFa5W9Ia88dvjsAr9gMopA+OkV4VijJgf9hZCaGDE42j2RD0rhgroQND0U
pW4G82uDkgbiS56N8GuIbuj1WLCaBCvmaxRKdpSBGM9Ggewtwg7h5phTgPvtqs3imgdyOnr8L+4a
oTU0BOieIE705D8/Z38RXuyZeHiohVLg/Z4ban2RS7MvHGkPky5XBfnh5d0ZbO20FClu05ocXNy5
VXWbx0B8yvjn8/b/lbjHzI2gxb8LtxC1P3yHtTbPzX4m41JwFCUsC5ySkXH2h+SMNCoF0jqj7iv2
uV1VJKK/SbbKHDCjQw1VX7YzRahuCTltL8BPEm9vL2qtworbY7PMzrJKyLItJnOv8K8NnyEjh+W0
40vxj87Vf89Oo+i33fhqRQ2s/0BQeA84t3M3gr/mkfftuNxKqeTZd9w+mtiZw3H4bzNdf3JQbmOl
ZSV16L8qg4zVIHF+7FX1/MYycKCaJAb/ezW8MhkLqIDJCeEcCfDKFdLxQ580+QhvlQ3EtmySxvY+
nQ9m9+0S/A9xFpnuIiHDeeOjkSZbgDdgKdHMRKjYhpiG/hTdxJCnBWcSs1gysbzTKKtAh+uRJc6Z
K7A4ARlO7nSxjAIpzjWySZn+lOUY4QZfIBKMGItBdtGLBBNeCzalFPYxzwuGL32XnY8mj/Z7QdVB
kR37yxDiJOyjaZoyMkJd78CKfebw1mXDM6qj2McgndrIZCWDK2eLetRrwwPdn7ZnjR1c+ZeoNIMV
E0xg+C8as6jkAl1Ptd5YdX4UM0Uxgi+ED8/FPg6yxplOj0fWb5/DN1w+Uu2JaozpsNB4rVFyTTci
YI7JEjE4Jh7BecHdXdZ+Sd/DreEQuowHzbux6GPUWX2fwlhWMtLCOdrhvRkoZaL852OWrRgagitr
IMelGLHma7wkxf6hx5FE7OTC+KaksfSoO20PsrahQr+1azyV0ZeSZJKZCVmmXPlLxONQJ/5/j/5y
ZkQQGgARq0do6t9Ky/+s46Qo44xNtnwUKueOmLQfWWa88YjNCOpu/wveuAJzVRbN8U94z4qWLJq5
YOkJNzbQvlAO/Fod0/k453J1VLEGeOWLQhjMglrKeMHgj4mSxTHDhcYDU1l7wceI6sVqe7OcFmS7
dDf78ijLsQoE4/yWehip64vqxRsKNzXDV3vAqH/REdr07MMvpxZ43skrF+AlB5UmGLO6KR7/nLiz
fSPK16CYLhaZK1lPyT4FALSkk+xfH70uRN3ykFrCEbfEI82j7t2yTKQrDzSWsbMzDf/o13BNqEH2
riogsHLtuQr+hC496RyvhdfXLDYoqs8a7Rrt3mxsjeTzjtQG5eg/BSaF7rXDzjz5VQyJsucFDSnd
iSDnKBzcPAk3ftviygxgC7e9J04cZoGcQItYqCECsPZAEZZhp1o1T5AE2G5IaPjQoDcTdcpPvSrF
0wjDqI4qGkRKQpMZYUgzOqxgEvYz1RWmmWez5eaWmiPCLWcR5tihnzQgFpXRyqPagjc0fy7GRjWl
ShDFlzLg//KWXepC5dkLWccVV3kbSX9AMBjnmZCTDdniJlXCUjHSCNVe5j1DQpKA2w3gpNxo50IW
azKLmLhiheFHoO8iv0C/Kjvf7ZQkBw5BLKgYU6mYXpFMtydPX5uRWQkZ5Dg+yeKHv3g2cpMriu05
sU7CRA1INwovnjoGYODS8lhMTfTFEwwFMWVk0dwEe6DVO/rMjU+KgtyfgLL0w85UMo7r9c0fyHRN
OmuoiVC7WId9nJi0sihHkHODlTm808/0GT4djY22XKq+M7qyhGx/dIahpVnrvFGQEya2U+h9HeNL
lsAJLuP40kt7T+VHayQPxYL+IBiXva9Q+ogvgqjTi3LsHllpsByu5nRMQd2db4XVSmPQ+ASic7td
vSPhNrx0CWn7WupNdDS4SYxnqt3W5AVatAKVMQDKLHczhwbUn2xSXf92YhLpAJvsTjxNev+SMeXT
hu8i0rWHwftjdnUSv5XhdFnQnks67fkzH/VY/Hm0gW0kyviChQvkBaPvxIIXXBmeoHCfOcKx3idR
W0xgFGRSpGICX7f6fP6yxDBHhBirobaC8G/1cCHCo/Ien0Zccg2+z+x299Q6D1J6Q5IqzcLeoKOH
w8EQ/vQK0wrqcsP8RtKa8eSVvgLC9R6POdfVpxztt77oTQSxvEE+h1JaUF3n6GHh6q+GMx0dCyHK
EXIrXLwINkbqQARxjiHAf9a0sk5bLZI6+pjVnUJsYcNtGGbPKwCZCRnTuVyv5RZJQhv8uej/TYRX
rJFAV5/H+vZ4v6+woMAXJAEwSTGIOZ1xvcTLjpo4kVLCg31pPwOMU9Pz/uyayQ2Xls9f/N9wEHwS
gvu5dK7NE4mQku5ySpEuZ8V3AS+ql54uF1caSsJEVeu/9DkSre5N4OuMm4UxI27N24VU7c65M/Aq
PSkl/Zqo+6NkOqfCUPv4QBSToX3PuWqun7T7e7GRt0kyTb2i7eITJE3WeaiqRF7UlXEvTAErdxQq
jvg5zW6YRuFacYwyrXdBOKPbJjBGron8BH+EaRVkbV1OH9O3mLM0ARQ3NWS8fZwh3RPMQxYb66hA
DJl4uOWJFZfsXNv9XPIcg2pyOvRXaNB7I5jlR1/jnhL891fsrl24Z8Hyk0zpo6nDT70FyZu3Brcc
bJHiUYRMCQN5r4ciJeItBX6lTdvUIk5MNzQsgs520k3AP68Jo6yS6aof8rtQINmr+Anp6m7B7uzz
ldCXrRb7jjWjtihzBkAPEAHSo7yQ7A8eqhBnRXDEsr+BQY1KjC2AFzNZlz55XNQgdTUJfIqQ2MEd
GYIf3+9AectsOGxUsdEfpNFUO32J8E4t1VtUhrOjbYDOV1K3Qzi+8t1jt2q3wzog8J9JgHiplamP
3SR78dnSbJbv8aV+U7W4SBTQ4Jppzvc+YIMkuWHUTgWWLAx4SweLMzRt6GJCbJdJ3xO/oO/JQCO/
3lns14BVI8nISWWnRwKsbhT3JtK7IxdTvzsmr9BKLN6M+JgMLAT1JWdexBlyZyAWhw6ti5cFflO1
2PcR1c1+vUXUAVNEtfDtXGAuLMBOiQstueFBgr3RI5snGyfPpbbQmPYsfsqVnNjZYWVLITBC1OcM
NRTNkN21opF6rrnlvtdEhAatNtRTdX+/Plo+wevB982vsos3ZBwWsYaEgL8B6wz/mbjjCKOgVAbJ
IvGJwQtaB/nhCktfRro+61rEWwr9vPIByhYrJ/+lXPIJ1NTuedZHKY3AiHcBeAvJdW9v+uA9tUrm
pNdRcpAs+i0KTkkdSWhpaHaRYmXeUgT0IhfGGs2uSJmmLLPvEdH/tmIcXQ+P131U3T/024YHjGHR
8PY4KoFp6SZ2W2Qz92hCcee8JFsuvvpCzKkkhUKgtfmvSSCHXPUhddi7LnyodzegpmqXrwuKUZuM
Pn13PsSLhdo63nsdb776RFHvCPJUWbLicfl1uAtawDzEt+V1bBJiSM4ZnWlybttozRsY61kUcFug
1R2Z+98/Fs/fKHm6Mx1YX2brk3Uf8h5szL+FcGdB7wJ8/9h4iCnwWJie67p3HG86YxGvHGN0kPsF
j5VPnvtaZ3hgadV2rVOTMRndrHF8hyMFZ+MR0kHqPBa7Nh/braxt4pHTYkRxWdgCF1IJqI6P512J
kZISgbSIwSNCXa3N2qf2NKHQgwy5CWhBDU5UVp2ojCxSytVpiSUVtQG3PYgo2GZuQ4SNPet0iYjd
FTSk7ieWkOUrbZa29O6/ZWEc7XBL6wEW9DYyWd8DLafHvbcuN3GL+F3SXCulf5QW3/C9V2FYxpDw
oDy849k1UlLP72q5hvBvTafDzgGqb5y8jYiac1c+vNKnGziyDFLbv5PDU+yDNgmcCtr9Jhx5hl+Z
e4BRYOpRgqfShg2AGK+8c+elbdPpjItBM/6+wLqEpZHcR7gFxW7NhA48/JEp0IdeU1+eBnCIlu/c
rdZTtS61JK/8wjjOoOPeCUFsWiiKhJZOW+Bms4Ps8351ebiWCiiKpWOhmfMTxS/mj0c0zUuPXK2M
TCPRSRf//maYVbpo/83+rkE8ObcEuuvMOWCO8ukPN4wWB1ZWJj6/ZWn4Fnun75IzmPD2O+9IO7OQ
/TzN4R/0XrzruSbVnNhx1NwwYdp/mkQLgOVY42VuvZB0Cip5X4AvljZJF90zyfC9p9NG5+X/uLpW
Gg1NmLoM+U2tdTrhF5nRrIGBRF4V/6RnE1pLdVO6yfGulzxkxuVQt57CJYDBUX6MuxWrXJ8UmHoN
Kx9DD/NOFMvxuTgThehIgzh70HODI0B4avk5YJLMQj4rZB10tfkGjSZ24nUAKxPOGvdMs9ldTZwL
6FJe00EYCDFTTDSp89NuxVrJ5hMNUATt/c4bCMFPLAvTP5RJEh+b4bww7qqZD/sGu+oJWoxu/Z/C
u1phN05rdKZoWg482kfpEXI3nGOerV0cdZmp+rVjEO/vu4WM4Jr4sm8J9/YOrfSGx/23tOOXRwNk
SAXuVle5+KIxut259gF3C06gAURpSy9rmlYwB1+zkeRsxqVLSLCROJPOSZYhFSLokL/c33bsGIqi
BHg3ikyRoT2gYEypzUTMj30d29BUZQktcnHzMtZGe6Eu2oCs49kUrDnrCyVhgmyrQreHVjaxmpLk
eU1lYG0U8yuKnzROQZnJ/FVE60DVkOnIBWQMbylNaPextYXe65YiUAQXVfvTdn6lKESbctT2qGYg
Py9yPdduwdvqA0JIoDQmvJ8+K4Q3LNfPTqdI8b+1i2vUGz8TlfzMJRhdb2jlTZOWnkkOmR8bZftw
BGGR/0riZubgHc7YscV63QEYAicbdjhFypejfbUrTziOhxlNfO4y1r+DZA0YvOmlNmbHJm/HO3z2
6Zg1tRrfzjP2yE0togs6g9AYYLLRK1RwRLzs+l7skqEOeEh6loxdWVCWDdaot7Sm/p4W/icSs7Fv
Fih7O8lTPzEV81bC4tytFbUUsOCWJHoMZPkPsMkdwmaCSbRzYhGHLFwzF5Bl5UOFqvsjcI9hvJlc
NsanWu0L11Dl8jXqK/ZP6D5R3Chuler8n64RIz15JDnqpZ7ZoeitdJmJMN+T+Ko+NX8NTsjqLdKc
6iPAt/QYflHxrX14BL+PQaS5ZqG7fLOTd4FsJmaF5eTjDvKhQPVjKhYBn0tVbO1kO9NqlL8i+oAh
6E1DqnepHoFS5FK8O6Ai1NrvZK4PmAxSdq5XNi0xEXB2Xayml/0bx2roWo2I0G0VmFQ+q+nJGtAK
CCCgPiHfXxqeCSMVYnS/X2qBfMvNhjoBhG72lzRtGa2iB48H4uyPHE+Gy7Vd8EIUHigDJKn4JRVU
bh+/xRvZS8sEklplxH6Ec4PNdVsPUWjxw3igqsB4e6J5o9GuTnKOi+7dkzvmsEhtRSFMZI0/2yE0
3B5mjb3lUw9klhMez6rurivF7TZYfCcY1HT365GFeoVswqXYrWGsinmW6hbYCpz7cYpnxvThWage
57vf7+e33DlZ7EHyH9E8/hKASqWcuAl1OwnA3IxrfyoLA7DdohoGKs6Rhm924ydP8yHliTe/0Ci2
dcyXfvA3k/3KW0SE3zz0gQLz9Kb/5nLVJLRTH1X56THMmPRPbokF01SoRjm9+aRjdIBtLG5fQVPI
JTv3XYy7Plf0UqKk4I4SLZFTGitnpdSg0iviWcJPvS5kIHlEasQSKGUn1Tj+QvXzgXSiMHoIDAhC
Whm5qPXNy/S0YtQpHuWUnFLqc6CauLieVJFSBu+WHoDSwEgEKrEavjdwsRyPpbxNvbS1qzeiyZDx
pAY0K/397EQ79sdbfanzaqqZKt/QzcQpdmWbMwQa7ZPLLR+r+S2PQ2Ha5zH+vnGOJBwL057qKwYU
XwdrFoYLl+j6cDV22SX1P2saE2CrlUQF0b2u3fl8e26bULgBoonIh7znVCyyBcrvDPRFOCYfI9fY
/ME41rDb1MXh7+4jTP8V2LIbvV5J7SMdYMoE+1kuzNRRMHRNwKizPdf7lWUpdGbCJjGBsXTb3vLn
Z/GyIj7+Ox+NeYK6GXbIfMlEU/tiF1DBly/fEWFxfeXFvEh+JYqeyQUy8eOFIFwd/nWdkZC+iGJF
1xeoYIa64kbaxsoiK8nkA4NGrTi5cf2zMOerBgW1Q6XNrfe9XT54WtwCnMJ2FVJ8ksBg/jZjElHY
nA/9eR3qMSpe6y9/HCRSbm2D/cMcSzM/FdaPxmlD0Kg5sVXElkHOs4ZceCe1aBcbRFbQKrfxT4ye
9DYT5tTznVRuyq8QD3P/sHwvuYikeUzWHazFT772f7Fxk2HOY/y2pHhmWuQyASZJ0NxIeNKTV/PU
Tg/dRPTV4ahvLua/NuTjNzjwKZYjo7zEUUjzo03S6CCdr7xip5BAmVZs/2LTNAQ2HnEnmLJtgZzY
VjXH+UGsNsBrVyDO1fRgmgRYmWSppfNL159CCpb6k88/AR5XAfteFfnBNbspbNnB8sIfBCIdSGwp
9k++gznOiKq6iNNUUPcMif5+CWre3c5LRqbQXKWkqpWt5o9X28Do2cIjENndSYZiLEVdqc2z2Quw
eGOyGfCylsFx5/ZmHOE8njAX0eb8Ht0m+wjt8N1KsA/cofniQ2Mr8tBxkGbdjFZJ8KWK313zRv7q
EgQnXsmeCG+yp2qyAY2gFhq9wvoydG4QZAboLYKNzYUQOqdwgJ2zRs73aLWpVvLtgl5vkVx0x2JI
jj70A5NB54t2Hq9PE9YM6vy+yAyvb/NBuegKhNe8Zk5ce0AAWmRbJLil70/vACncPXnEG3tjTvrX
9+hJXljSgCFn5ilg6klD2rTlrTsNDpPSPZ951y8hy6aoNTQOzVP0akQYvdggEG9/kFT3vgt4bCot
h+kPvsYHlulBKsjIMscFzCoJ9j9/kcTBDmIDhmUpkDZClo75BbsFX84/5h9F3ou44Trj/iV+zCc0
Bkz947AvZW429kY5yUcHfr6tBBQjf7Zs2p+LCjI1Nuca+3lbSDhm546Aokmbbs04QP9zWxjVLfR/
gDbkwrz2GsD2+tKOy1TtbTydP/GpYrHSI9jo3YQuijfYhJLWveRhuth8ohrn7suvRty0/9rs3v2K
aKshXmycL/gEjLcrpgCWrFFseUrSDgyZD9Kv1MvWbcBP0aW+DqN0PKfT3nFsdQtZvCkQR0f5FFn0
fHkm4Qsa90BIMXQ6JZswA12HBEG68ZGehe60rdLVaBq7G7DlhktmHbk5YP03089uCFHgN8hh9hY/
45T/1FiyzHJAvsDG32Q77eU4HLzTGVYT3rRdnxe3qQMcaLRkwlmLDIM0zLNsQgiwoC7qAyfh2IQ8
ALV9PJEz+55fLyoZoAbehLO77Bq7kYJa/d+CGCHBHmUYsiLDnoxmUtH57OouuabeMYah7xUTjfF2
letVFFLMaV2HmmPbHFjG4L9u+cpS7G/V1lppn6dv01oxwUYtNJzy4m2z3mdLNz2CbgiKIHfEMb4n
Wq/tF0yD5gdMGmYPMs5c2vuJ/2jyaB0TxVI4Ogqcy8lUGlL6RLy4iwEKeQoHeAqYugAdQaykK9ic
bM9SPuHmDWlr41joPA4TBO3WzL7w5FavV+7xfU0fCWLbgcnUIROk4C7nJ0Gb3cRzsvrESQiwJXcM
KapTf65clPFA2zweEcegkVMG8tP0n1kW9EVuRCBWnF2Eaew8QxNNKRS2iGHmevRV9PxpH6SCPhNT
n8UO8f9XA0GUPFkDr6WRCWcJonhQ+GYWyXlSmHVihE+grj0VaRLmWhvaUGqK8dQoHldOUQhB1xQS
xm53petu1aTZje6CWJUqWcYlMpHJkg1hrq7QCMmVxRFqdoCCrWhPhSE0dYrKu48LNLh6SgvTFkyX
3iIpme+ft2jX0RhbRTsKi+gEmNtLlk98yPo7UjAu48hke/+TmLTTCBf93PEABeGZ+RMd99ch6lfu
JsazjH/WvCrjLEhR6zda9jmzLWXvzA2dBWH1Php7OFaFdFshZzEhl134MQP3mCTqXQ8pnTFFlEOg
L43qcDy8uWOAnuf6YoGdwwG2Pc8q4+HiOryAvFZfghiOXJ5P1NCI5loF4YZ/cIjkNv62MGF3ZD3b
JjwaM8fVy/d7jareNHVl9GaK28b/bi2NvjwUw1dDKJEESQQmR3atIjaAWSpXdO/Vv3HWWZxGNlg7
prJ3FlSlL5BfikwmSo89yQVFRHm2Xvuvv77uB699cpO+5x30J8LJftLP+Op+RwfhgJVPSmOWnqvI
kh3VTuAWmnWx2e4x7QzLaHMn3wgj47JBWdh7Twnx8Pe7viZuU0GxuM6qHRRwc64lbJsK6FIWHgXb
4kX1rur4g265uZTaqLrecw6+w//w3F3+zS20RtndQBBsT2ndDZP6n4Vr5PQv85BBlc4X79+APhkJ
01j4rOR2wPobC+RgKBMzbJnoNmzStN3g1NBSidX51ADsiKCO/GUeWE7spiSGSBknl3+a6sLLH9HX
K3e/lGpshoIOF7SMnZJ0h0NbnWXglk1nrbzWLGv39clxNV4taH5xhZuaK4uDEx/k8aahdH5bs97S
bcK4p0nxmfkQG61XjK7XjnnqGspeAs70/f5V+eSngKK+D/6MORTyi9jtOPXVXPqeJuyFXcaUb4Da
qsJW+lUgT4i6pbrCic3aafxGZgox5fGFpRWi1wd8b+TCkSjrnmkjtJPXIZ6yr8stVYdUq1VA4mXt
rHbJ7KQSjexFVt6XTZ/bEyTyalXVvuFsAcDhqasQTppbqt2hNPBKyn3EEKXymS9WunRRm7mqRxYH
VwTUz2LCOtqZN4G1iTUGzJWpazbAKT1TM/cmvOolRc1USdHNd1l0zkxqeXTvBw3BysP1+cGlAECy
YTg02tSH7yoyDiWxWn5nvhqFMnwj+b1AUgD1qcX6SEbSinf/rLEaBBtpLCwMxms+eg08gow9J39j
xBcfBIIbvMXrlhDVDPDLpMCST7ZGHh5SwVhmraf5hN6/cTzWButYVkssvKu2/8HAVHMBHO67Nka8
kaOsA1ePzxtpD4smJXP4CVEEDaXXn8GM1AVx3fxHc8KyQsefi0UGciyBrZtYGbV5LRaECBNfsyii
n0GfAAVFwgd8UGzRAXKVXuyQiZTkYV8YJ7smz8n+IWW8H9wONPhv5Lci7BQaFcYBu15AEFcBZa6w
5TAqhxmhe4KF2syyHlL1x94KumHUEwOOl0A1UoUStFfa9pi2nNk8ywPUjHgKku7vOKhoQHwClnZS
LSyd1Hpi8auE9wzzrijGMYAhtCk3QbPAck+93ywJrjcOD8D8OIbyrU8ywUdxYfPpW1788XBQW7tL
64r6HcsVVeKG2TEuaPytZlDsZjqAmZXyA0EV1c5QiNBl/eV+H/vmDhbLW+c1W2zNFwRU6IfCo/r/
DZ+a/L63YyjLYj7qxrp0nmM9NxmnxYrx1Sl6n5OVtRGxA/g5IfX9AVNEfKDrb6ppl5YnTfS4arjm
QvCDFg2oBnjHaI/ICCMTRLFhjTpQY88D1T6MCYtnnlhCo85ZkJ6l6grMWVHSyhMRcK6WGH091Din
I0xkx1ak1a4KcTCDvJ0Emwdy/ehbf1NhB1LOy+LX51YlnrkwgN8gv8dBOZPwZAjtV7BUhzi3DZRR
z6v6+vnlRTfI1qAYcR9Br0+0xJdXbqX39goaZbfRzG8IwT+4ZK/RvUgLG5LfCdQHfAhcplwjMTRl
I71XTRagHOKCpbZYBLM2SJG8t9NW3dR5uQnuqM6QCpnDju568JpK1KEZky7oA7UzkdqJj7s/Aed6
Nzu7wK4PrtCXSz7uIk/OC7V/1VNIeJ1Dt+AT3Ro0JowMq2umAiADmlHtkT/nKPMibF+E1VFCzzxY
yh1NbbtH1Mzak7YwtzZpiBew9tlXkPpim/BcFXkORfqBFFm46MUSc9rDCLxcWXhqe50mluIHkTXK
o2q0MEIx2pJIKzlduI4PHbaXRaWJtVwAwVCAUnIVCzgQh5yx2NP29CpdSyjEiv/VsBEQvlG0cA4f
pftgRTrGuOP2z/oumAVcSKLvGakesGvFqatXdmjqJ3TpZ8eR7Cu17HpZX4+IxN3Gt2T5pD0a32Om
XGpcMFWYrmCeAulkoIYJdx0xP8m98mYPjosZCu5X5ItFws9+2BdWNbX4HNK4nVboqw0Z3FwIlAdg
Lun6xcEh01rF0uCHG8xhRRghkXFa05F653pOG7U4Q3W2Q9hb7Uml0iZxsm4jZ1sqNR4BDYX358OE
RR+JX429hG4TNxopOVsHoEIN234KF5mcbGqgiI9HCfgD2lVumu3h/35H90OwtARPyRwtrHEpcNBy
AV+Brzv0WNz7L0wRMgtiX8AlaOXFZ0VloV75oX4TXt8o0VChnv/LScm7D5ttY0G8If8b+3yuISX7
KZf7awuZassEiLfYkSOxqy+XpjA9l9uQJCcTDd/vPTJ7ltk6xLquV/EIAIUkesjtINKn9O9A/3GP
giVtoo6cGH+tb5JV8iuMQB7ZuNjgS7ZLMTMKGJysnPDtimIgP9WBgjB8IgUjrKxjdPIfv0qwIWyu
6K02BDVVPWlFC1iPFIsoQg45BnLxyTmj22Cp71SbNWVEPfUs9pd8hpXUGPwBpeoW8sDa48h3b6Bk
4jmEIy/+XE9yCN5rOTqc0VGC/D6LuYk+Wt/18IyieTNmWNpRlR2EM5LxxE9O1krzH2H/hseWF3OE
T9OKFbNGoZh4KPXGuKiOd/NBq0DoddkQMf+BvAkSI5EEG6bKFkgoKF2bRKekAIw8wPMLbHFGrvBG
KoRag51nuejM/HXMW2ZoFje/E/aWw/sm3bYr54t6xrkatFW8TwwfRCW702ajyxgYdgbVJoFpujTm
lfXnF6zf/UD9wKrFiddsgeLASzlswywymaopQv/2lSpXW7bgq2OHigf1t9RSeF90jYB7YQ/0eGVv
ps5RG6IY76vFW29IUBbnnQITtf2e1nqxFwVc3FL3NXijBy9Krh+09bvRNtZ3b11g2Ce5ouVnMs1V
XclamGIS+wTN4vxYJNcCVR5QpqpFGM1SV4AbjkOkVfDB9VAVy4yK6y6cPXlNGaq6B2Mbg+7J1xFN
fDGX9LnJT3lWvyh47tzeQ8PjgkagHrnH94Jq78A3jB3FVylQo5eb/cC1vP3yYVibUwaW+5XtxyaQ
hFwzy56YktqIefvsPxxSo/9cKIKCN9gNSPoK1FIDvrTD/DrEwfga11y7SHUj5mxr6L956m5Qnros
UyKDZILBQsLNwdHsfdAAcqydbW0QZgXD7sTGRGjGX2T0DCRm+HfNxccR0FYmAKbe2KX++k8hhdqb
+xq9hlBABMB6V4Ieiaf17fJZ3LEqrr9D84/34xk+7oQB5YSliPj19kQS5wzA2/y3B9kWP5b47I1q
VVnc02lVG7/W2dq9DradgrM6X48gQ2fyuYWBg8rJvyDNkUof02bVVs159G92Hrb7sphEXabAI6dH
vvd5Gc9orfvUx0nCplbpmaSZIZaoospdZpPkVuNFb812nE+pTg4TlnK0zXoXtFmVG1gaz5H1qMfT
Cd4F7OAkxgLhfeS0T6c3zZZy5p2ILErlHwaPoHNiJJDeaLxQS9enamq0Ezu0oaSdD/71WTgVK4hI
tweeSQdPODXlbuOlntv9WFFvz+GPDySfyKgD2tyfsRfP+htkfzj3WzRnalXb4+4EzXVw2ditc0E9
OS+7CGJTritWpK6KrL2Fb3l3HP40E/OyI9QDT+Cy8XEvpArqbycKk1k6evYrrUduLrVPYTFZ2BGS
cxkBQENfH8PvRRXNDXJO+N1EfoHCCdjAJ9xIT/uDymLZlkVBxHkE9ziyBhw75Ej4kIs1+hrII5aX
73nKYpHip2uic/KcwNF5aSLakCzzvdgaMnai9v4b9YX+eAk3klfVcYRMGdbs3MguCGikYNEr+V9E
nD7JXvFlnmdG21U/qBmuI82EQMMbCgpmxGsJU9XGxkZsnXO/b09RAoNzz7oGFH8ixH3Kp8hF+l3S
Ur+LYpVQXizsyppSXOKovUZ1HJ2hUg8wkNa+X4pPqjUbgQQlEniCrRu+7wlJnOrxfv30CR0oHfhl
3fOlzwLaSslsE68XByJxGsuH2kWjkSEHd1eRcIUpFASdw9S/OgaIdMzwSbDrrdJI+93ns/AQmo9k
MxzKtaJ9ovziirljpG7DqBg97WeDfUNsJ4Rse6ZXWAjzFytEyBMJFqkPEXGSipm9jb/vi2T6svFZ
1hgOYGkEhulvf4iO3btOmz09FR/G4CqNxvxoTNW1IN6KnfZ24DlSJvJgsCi0rAMXlZNugPFvE1lw
/hW6HmluMZRoifuPR0VuyX0iJO/9dVBhEJQMJYLOcvze0EyulSoxCqdv2ID91J6rb/wm7ZnNVwRm
YbbAmdFcAwXGnz4HnRBsg97GlSdPIfZjpVSlova5Vmiy/oLtKgQ2Y0tJFjI+C7yp/IulMQxul4+W
x3iL9alaH2On+S0VHsCuPde7AkDugJU4PcxCx2qB3X/L2Iy+owMn47H2SiRWwoJMNc1us3zQeP4N
YLc7K7gEc+zC3sDUrC9gIPT7k2DyoAfiQtkhzZxoP/GL2rFg4qx64wg1AgRGRQLrW6QUXeCXfwZ8
hvX3/vPRinY2oDpaFmrIMdlFaJxcWbU3mbKY4ltR1jBqpdM+pU1yTT3bZwQBn6hnfTBiDL0+YbuX
wB7rQtyOihValIzCRaKEXg1ZWvj+Z317WANFwg7fZZE58WmkPxSqu6165UqEkSs43D+W38n1UVah
QrIGwxJplJBcHQpzJK7a3fNj8rNSdDgehc5Puj5UtlR4rjH93PhVUs42w7XwDB/zu7KxofcHGJYV
ydGnRhEdoG0oWYMu6EyGppvn1gL4CTBU/Jffu8SVr5c8eK9tEiZ5b4fj+YNYX+uqIWiXt0KKRECa
MwckTyg35qscbbpaFKtobWdFMcZLZUsQmeXsi/ZsMH05Lej3Zano1VPMaQ770csEohVphVdGOCGj
ud8KvzNyEDY5Vgrb6rfd4mQY0uXCYg4betSJUIeA6KV/q1j+yArG+b9GIYShgzHrmbQIp621rTQ1
UmBoLRrf+CLWye1DdYr7Vc/UYWHl+Y5Eff/zAA3q7s/62DfOrV1C6EPYX2CMYiMhmeXt/XyboLI1
F/+pK3xmYmQNLPjkrtAmCLLeO+Suf9ot5SViBP5Hpm5UydjW0OEwMM2xRk7iPbX08KOcBkW6PR8E
hXKaDNgIS/UdjqPzN0dBNatveCSDLpD1ZU4v+nb0DBr7IbUf6Nr3CwDCr24rCc7XRAQdsfaemTnk
dEUqfyt/PskN3M8+SGQkN/uvlBQZEERw8Bx+WB7ltRAlOYMP//vdJV3OWHMjf3iYcaLCvPQuwiKH
JdBuZjgp+A6+RY8eKhRxTOgzFaolcmLyxQ2YmXWChKnZWWY26GInm+ZIWaxlICZ9ea4kntyjZw8o
8vy/TBhHaYLEFzDHCQj4zPlRhWMeaCQSyhw0ACFBIiaFcpoZl3mbLUIE3FFcZnb06+huJdoeHGrC
aLDPnRHcy934yy4I5C+0uQMV9In0zkUODEFg98UVkq4ffep566fZXhNw8gYSRGQ+flxz9MqkP16Y
VE/WlsLIhR47tPdWa49UqmJG1bqUQnIzLe4r/zNeSYL5CzL1TWNcoWcoPNHBT3QMCtAx2VEL8vmZ
+Ll5AhBaRgrYilj0ywL9CaFcux5hAg4rO0wRty298BsT03WyFw6xl7p9AxsN5pI447DYBqoxBbqV
0S/Gx5YabtbjzM6b9//EMvh6Uza448sLhLSEBOQ49caMl74sQGl2+PsRlWy8M/MqRXCsb5kVwKl4
ACRDiHm0g+u+kEL2kmbO8BXss9NXjjPQQ2qYgn5Y9Uf0KULOwFrSG/Gm7YNzg1x+0Qbsd9OnHcqN
0gozO38YliRmgaGIElk6ClrKUyAC4kI8vDzsot7t+7+o1nFee17m1OSp3PoDVmRhEl/i1RzmmshD
59ZWIBX4ddQvZqjZm5/x/IMfdu0Kdhie2exuHA2aSVte0ZDY8mjUEj3XnRXQt73jAfdySTdmzRyE
xZfZ5cw0xkVRsqcpyhkYwcWKsZtodCU8DqamUiRrP8hi5m16sofHqlIPZzFKRNors7cjgvvf0ej4
4O1hEcm17DioegzUVeR1nY2EIPOPV4iwrVN1KVyyrkoVRM4P0wCjlZ7kfEoCNkR4f6OgdFGoPFCV
cnUEk7NOHyyi8P+Fc6ahc1MVE3pepA23uPlNQGYFTONKns+m6OSZ5HWp051Cu/hki34TPzchfsB/
aKg+C5umUiZ0Qi+NoF2vX+DodtuwSzyvIZlxTWQdiIBljuTDJJC0i15/WHss9928wMS5cM9DM2LU
leuJyJXFe4cKM4KRF06lrOQOpHqYhiFk0a6QCYNiGlIkv3FD6roU6CNoSoDcdcXavFFolVk9sYeb
gcWD0wdtCCmyZ3tl2jBG+pTin31g7odRaiDOuw909SSv8zNV11uDaaItTkf3R37AYALSJbjSXTmv
3ARgWl1WRcRUDB8t/si0oqwadaUfRwopOh7ZgKgvzU/BG0MRtGLsV7/phRHcAXOi3hP+ClV1R7uu
6SesEs+BulmIcSTpfXWZvkigHoGSZ73VGH4RxQ5UFxHDEV84VXSxR1zKE6gSQxMqkviqcmLf0EEX
KYUv2UH6aZzi63XLUxTNy6W0v15+2/U/mQ1g+1hEiI4YB6lZrSYtjNkh/adhW6XrQ/J41jHJ8ImQ
bd0FsB9u5bLrrT+Q8ryzwpGoTfHcNRAVRUls6nuN7SyIWTT/m3Jxlvg3z1bPnfJ5v11ThWUSAqMy
uee98zUwZIvYYqXvyF1oUXWNcJobKa77rjEiiz3PxlcyQrO3u8fWnyF23uMFJV9dT1KQqmaWYA56
oL+WFPOXC9wdVl1nWueYKuXsv35K3/WhynB/1RO2opEgW7bQKQ4Ch8OPKRSzcpJ1nIO2mbWNnt6O
Bb3quB5P/T5FRS44Z4KQ453DewBhKsQbYJ8Mor6R1fal7OGp45pVntNjXh08DbNThVaxlmqB0yqL
7u5MkVXEEApq1Ycf25YrMKK0Zfmrs82CMlgA3fODMKN3cq8wsnw7m2sa7vIcjFhju9Sm2YEJo+uT
/JAgMEWMJ8BwgCytkVMhZcV2G4dbnlUZ13wyb5se63HwXQW8TDo7Gyd3uElYEP7AcnxEIsd9Q5pZ
3le0R9mENArQgexmt+Jz/1FE20RGIzz/arIqmDcXa8Qd1b7Zb5Ro5+0OmCsoP6Bi3e3yIuLzS3Fh
BGod6u3jnGGpSXgf+OaCq6v/M45e2H7Tlv6aJ5hmE7D4l1ZKFILXKg0gR/EkkcAjDL9JDHWtdBKF
LBNWzJdgUtL8Af/hHCCSlNq42wYxB8F6YtdTH1zUEcTZNeEo5QnQwYI8AJB0ZibcoAEuqEALBt5f
6Jf+GIw5q+jKvPAmfbGBQkDvgm3V3tN68FSi2VgnpqsB19HGmR4fOdUvp8x8pRoH36q7ZnGt5BZM
ApVzNrynVXaEyZ/SwjRz6NDGh/Kv0uJaSqjYUv2E1Wgg5YyUprT6eM8ur3zLPGuYXWao7nPlqXDE
RbZUJOWNXRBBIs+cglA+p/kr0BeYUOYmr8fv3jSt9bZGvRo6ZWDihA1rlEIKV3BYf7AQgbSjn/w9
jVc6a+/kGAc3KHwRttj434zY6SPmie9eYirVte8O0/BXOy35esURbvWeSozmhplvhoRwLnU/IZy7
5hLPbkgclyU4akGCwqOn+ZXdvHwI/cBURo3kMpY8oBWfyjLQ5Heo54y5zjIekyfSEE13vEKZei5g
vWdYZ7dPh47gpwUdV/HfkxzeuyIhjRn05q8L5F7g4XwkNgcO75CL2h8GIQvvfcxPOTumWkwQmGdb
BFeRa+KRLGxgTN7FkpM8DvIL8lGYtS8SSv4rlbGJJhsmcgONxHErS++0dMROBgJskMFVhBLD9C+T
5pr4juzZ/ZTngOo3PiW/XxORTkKyc2SfUZMajv2QIwRjWA5+RAe8vxZ7ydb+p0+aWcKOWQmITRY1
9PaxImG4+hf1bgXOAxBjJID843jCiU4SUpy5laha+FAEsu5OCWucyLLrgj+AXMtFX0ryqpOoS4p5
/Gw8X3kaHNe7iIczCylZ2QjrdJnHS27X2bYzY7lb1v0FD6zmEAcbSfqctb5vTsL2917TrAA/SRKn
vUK0dCUH8XewGbenYqRCnJggh+AwxVCOKGG6U4ibFfGLf5dzN1qR0ah3R5+4bdXbs9C35/Ska/pi
ujtWl1aJ3Lx31ZlUHT4XdxQwyOdYICd02NUDyjYjFy0l7yYBQ5YD1P0jQIau6o+GageEkuzzSt87
gbNj63HsHzvkGe4TtUr1hEaR9SZcN6IGuFBlTMcLTdScSxxOh2JfZHk5r6ftsLvAg0jRpRwKchUo
++ECU1EcKDaYIcADwrZGU4chFIWvMK+wMP0Kxs5tdXBorEe9RlsIbfSO99VYaq00KbJiPvKtMlKb
QikhxPCgqytysA7vv0Q863q8bJGtuRIRnBEgwf6Ap2UPIEQxrKFJj0q5dcdExDVPYDvq+KNFPlqk
DtGJcYD8hpfwJ0YHo02ztF0He885OhRHW+m+AWaWzmdB5+5ycGCGU1GQHHqLg5BDvA5VggLUPXXW
COlF1U37jXp+luajAnuioFsB+awQX39Hd/6GhHLpGnZFR/U+xjxRuT0RDCibTk2ZHLEpbKAhQpaV
YAuHAIMreSBgZBhRKpFM6RfvnAcmNTtSpzNyl4Iu+7AiilZMhRRERPfScrMxbbOMWgPUdhS9Qsct
WVsu1sjNKHCkTSky1V2Pzaq2jemEfH99q4aw9gG++Wf6Swjs2goo7sD+QQyKAYGWm7cRqruUY4zF
7CB2mCYwkqdyedNrSBrW/uGSRqsFbD2HYKGF3vVx45OsiTg+jkEdPWfZ9VbvVpoifNPgh7gLa+Ou
rp+/VBbBV5kx118emphUOogtiMJp/fZW9xW486WiIlCzOBFMAj2A9cExvNSIz3UGxolq+yk2fq4L
huwwnWy60BbPkN8Nw5xwUzfSug1NC9gmeUtlPvSOduQVcHhW6T+JQvkevTXqv3I48qWq7gMyXZo4
BBVGsSUgMWMOCe9g48zOvxwZdXVzlhI3P+4GFyYN/M8ZD8tJxiTal0H4kepDSqquCaaT8XDe7PgW
eCFjNK1BS7GVqWBxXaroQypReyxGq+CIonOcKID3U38ivdEk6ZjK6FLCfGC6U65rEjjFcvHYMyC+
GFB6dOqsw0O/7v2vVtGfI4DJflomi/qiAa3jaITj5UxYMERVW94Uma+3sfbJKVxtjh4XiRvUR59p
N0nVdZukO4M6MQRrDrIt4haJ0uq3qdrG5aMZ7R/mcTuvwny1iRF1U7gP6P3EjgkQyMpyf1fchiAg
XyLXmOIc/ZrTizIDb1iKrdveiF1Xv0b9BHIYtwCoH/bP6et99RQyd0jAzdZnN1Gd71mY3SMz2xmZ
+Vu1D2O2Xk2Cm9Im8QjBviGMkpfS59K4GOzSMN2qcb/BvyPEb3etvmDpuXzUVBt6kpVV9imAoV1Y
I5LIxvH5TQQfd7a+FtffO2tVF7WeGhHwZtI94yXZ+c9D1UulAzWNeH3SyBqCJfTcn9CTC8LFyE1B
PY0Xq6bwqs6iNVJa3pO2NnDxcgY+fkvd/nMcOHwzAek1EBqmDgOe3MI2ZB5oVZggdCWQ3RHu1mZ9
GynVShRMA9X0VF9QkWHo2mHq0FrFqU9Ox3atOk3NPID55Pal1pSMhDreQzjopUOl6LGm42eDhkhx
h+ONVd8XaS6RId2ezi4ssBVEH8Q8oI+hEjXix1+FVhKwXzdfFRK/tFDNc6a4csRuh4bqQdukaEa9
YJ/hCBXVBJCrwUbb+AwysG6l8OE17ddX/7JcQxUjkiuZyd980f80YWMKRSiTUnIkEu0gC4ognQHX
kpxWhZa3rfR/dyxa52pTTnv2rxd3i6XnyYhTfcoPIpAagPgUl+UeXJH0+7pAVoL70XPEUhalrKm+
jZHSSDziuV2H0cXgXhD3QWdsFL4kz6/oweJ8PAPjyk3iFrkYEHZdF1LAKHh1trMHCrSP5n04PqlL
XmJ+XYmPdJ+m5sWzl/iJ9fy4L6MXZhDjB7gy1zYwZ0l7U7zGPWRc3R3EHqEDM7cKePkCf04zUb01
4w+boBcsHKX30WNVPHK78FJgfY2ipt+sq56O2OXGhLMkY+/lTX16agrc0odHWL8jUjNrQrN2D4bN
V/wYuRMc8NZWKTW16SflLtCfPUfFKi6b7SENbca7nDbHZMAwdCDjkUpbzQ4RjnrYE0faEzwnOKQN
cv+z5YdbktrlSsqbB2tbgXayMoS4mXH2bod89PQye8rOukDdNGTNPa9HTzQFPknXjQcM2G2Cw/10
RoiZXGxnH6f26d00IZvJJttQu52INRWrgTePQo8jIszLFkPTnMu0GXw2U6aSa8qW9sF6Vv625vZ3
HfMcrv+JV4xsiTjmnYKyUrQGMuaI6p1YtAgn2bjFf50df8a1580REE6LyGmfoCcNEbgH/QjbtpQI
DV0W4+dwng8hhxewxPzR0PTkUMoazEhZSOhARFsTprsqf+nO5RZc1kBYa4L08qm0hiyfluBHmBOk
xtI/L+GMCnPenfnYRK9/vtEVgZxaRWK8BFZu2V9a/18A6JTvvP05TiPv9ZzzfFxSFvWYV1yO5Q9S
Qs3SnrvfDfmHPYv9EgvkuzkzuoZ7V0EGNVnX44UXYHRcIOoZ9J9FPhkkt5reOt0EcDkBwkPa6WjN
/Olv+7iH46E151AX6sh5EHcV2hEY8uUy/7ErbxT0cyd8hgkzY5yo9opkghm5x9qxSMq6r8oWIT5X
Hp+QGoGQYf+eIbeywLlEX+i7xIQUsYjKrAMkWOAxfqBzijiy2E/HURjEbcG7OGXdvw8Wp8ykZSdG
FyrdcvJ9b+/qzjYCdBDFjcz7dySCaAGigoo7h7yE6DT5wxThhCE3hV3Hmi6WHC+QMgYNC46cYene
iY9VbF0/J3LNXeV7Sekdh8y1Z72hiZszavIAo+xtECsu+xxQoQBvqVRjRRirrH5fuqLXcwRL/q1d
TJwZ0s2nCFJ4NWa3cy6dpGviJSMMHY8JQvlIRhpWNcxF2mlICaQtjh46JnNIKTN6mmsuV3qFUSyO
6vNf3U48X0oS3oPQ24sQYm9L+m3cIo/ljcHZy15iQviOuJVoFORmumpM7ECJ8nZaybv47WNO2B51
RXYAqNS3WWExcMtUfeixVdxoL7rS5c6UfBTpTVpTVRua90SwPHQ5cSfNxhDnnPZFp6MKI7+JpR59
Z47gEoNkHaBurze34CD+6wx0B0/4EX5SmqzxYO6atR3i7Sz/TyW583NI8rm5J5TFqgWV0yILa/jO
XHOUGBaZuDHTQGsix2wcxgspoWS1w8sbLVij6hodrRoDQHif1LzD2TF55+UJ/XJTfWRiul9AHGuj
LsT/9yqbrj94NogvgnVQGAAl2enAZnvHSx7aXtCcWQK0olaRXyeDrnO0SqyWYlwav2KqOnicvPOs
jf/y+ewDKAYtJ50U0zBPaJBEmOwwa4rP4e0oddzGkP9kdWaP14o4odvSNiy8N05qNSrN8E/eWboT
8UX+zlAMnOHu1bkIUc8UF4zUn7dl2Mdjaq88s8LT4Wgb8p5c8H6QaYFjqwvI7Knwjm/NoZ37jzyI
7vF73dX3L8p2m680pwBFRaCOZbAth/5CTu3EDhX6Bynvr1wgWCYic55my542/jitTHRqJ09sdK+c
VkmtAC9994c34pERJEfLTQSvmiUc1iy2Vfoqp1mF0Zv9UCkZTpL0Otho/KL+vz9S2WsniKbc1rzV
rJi5cOJQD+iSuxBqF9zUL/zeMbBkbX3vPNWOwM+8W1S0x7G4+Iy/+w1Kv++VhIcgCuqjE+Qe0KhC
lHFyO7iMVdRBDGqQa574YWgG08AConi3jsFC5hwNMbeULZPdJClr2v6j0F+W8IQnBRfgcc717cW8
+DQi/1eH7DWhOaF6cqx3PG9AZBpXTMlYE0EKu/8EHThTaiaSzlX3cW1IgUKXZpyTy+vZ22Zm3co3
9s+1TDOtXmllx74HrmnpSOQcXojlJGUsGYRWcFfM0Ba08ERvd5uLdNPci7jIRzmujgCMGRpIjx2W
L9XiXlUL+/lwHGmUlnW4Rln7FBjcvZBLn735k5eC5jvBkU39yR7PAxgm/5WHRrxAZs497bWTO/uG
7iGwb3HEYycG0Fk96uc5JL6uaoO366E7C6X/A7iJXnBQRUb2lcKMK74xZUEKzZE+0bcTO4jx+XbO
/ZbxYP2XeOcCFdVmO2jXkQwSO4jNrS3d7Y37apdMXuVKeljN1qY2esob7MP8qzgFsPgPvMcXVhMt
7NAQyoRAe3Y+tILDeIVfFdO5rXAK6nQswafBBKNfwXlRuipd5JTBxvvfuunJ+pGEMtO97VZ1a4fB
Y6ImJlXYz1vgwGMOEnCnGAuJ8pe5TCLUTA+kruiHQguKTj4RWerow8M6QALsz3CJGxqOkLLVk4Ij
u+AkAOqcTvap/NqZlJLzjUBSvYo7rVnGtLyXjTBtE9KEZI8ITSPQSdSQUO3dDJz+LlRfi2hDBVYG
xoHhxvjvo0A1JT/tWv78YCsOZw7L3N+WZ4mNo/30cRWkhy3X+expxVRIDlyyz7dfxZT/avrv8UBv
mrTJEp9o+n9TGX/A5JAKLBoGScl6915DMQ7RGl2M6IJiPZ5Hdh2OWsnGGFeLOndbgUkQJGQ2Zg3r
zlRG8EIA5zEVjBYrOyzJx1xHS+LcGRyvK+p7ufJXzhVtk/rECSSG/HaGGwwVtKk1ppaV1cDYgwgX
xrecUsSGo64+K6Dg3Zn4AfSkFwFO5uopOrI/JE/e6TGpRrpD4Vi8ByevaphsXpIMXz/HrK0r4qpm
IQCqfxjJjhor+qKUjAdtO03l2HKaL3fCddhX4r58fOQMw9n0D2vSHsILWbt4LODenfU+jhSOYoTZ
FAtwH/Eh94c8jiw6RuuaSy0PtHFpEDdqRfRFU4ojyLtA+S2LDvET/ZKacG1jWlHTk4BfezwkEQyw
AMPAF/pnm9C+S0iOSbBaXbbclRpBtTOAAR9+4OVa19ddwSJCot8yfJqNf8gHW6BKrga5jm36BlbV
dQvGCr2safI15ZY3K2WXIhpTa9Os5v3Ci/VQ2nRj05YEo8kxNldME3XUd9lWVzrAR3TWyaZ8SWRS
91yeeZoeEKuyW9sRcu+HjGwCx78UlIfH3eMfIBxjfn27OZW3UfLBl3aT/iJ0dKvmz0jUH2FKz82n
Im/9HNxdu2h2U3RulmPKKWu1l2KrjL7fwEMXKjSvAoi5U8k6Jjksl4AkTxDJr95ckHTw0QlXR6ub
WOutJYFiX+5dJoNw/0L4eiKPQ8kurh6eoxamSGwv9XL7ZQ4SRiTos9+Iug6JwvPt04fSNM9qlmAY
ACTunyLQ6gY+0vGRFRQl7OqSH9G31yaCGKBsV4mHoCQAT1nrOWRlWU9MEaYjO6SH6q6VMR7+Or/4
YyHtfURtv/UPfPL83PId9/a9SOguJwy+KoqFOB/1CuH+23Jnv/rEaFwNXGuwqeXhE8G5KEJsISxG
ppLioJMIhW3E923y5e+M0v6TF191NQhAWHOPA8yu5yMIBHB9OE8d2sSbPZjujMiKQG9sE/ALVx4w
e71ZRI0kV8iJFsbmnCvrBMFuvlDiNs0pduZipQ6MRrbw/Sg7bFGkfHOTPCN+xVNLzVmzSc7B0HWt
mybC295XAIvDNOiZWfafVZeCoQU3pByTylI9ySpoc6cjeAhwAU1tn6xTc3Y7QNYBPFNZE7UTU2t4
53uoQ/eLejozqfZDCgpTGjSjcMfIbPZMAllzdrcIVed2HpUFuld9PovuWMadPIIctnJkN9Txso6k
52NQVMuso2iU0WPNIo50N9HYyQO0CcWr5S4OmyG9xanVmkxfzHd1Y1nm06MTJTz7ngkn9KC28EsV
vjiyPo9Zv85hp4CZ2GXnxQG+HP8yWPQxDp2jHPW1QjVlXc7RNocrMmIoh8Wm/6O8KvLd6ELiv+G+
R+KENfgI0WROWpEWukXQiGCAg5l/OEEjeFzvTqa1eoquwI/YiUOu5eW7fE0U3CyrLV1qQcNIng75
+xg9A6dgeEFJ2zUHIV7DIRygWIOEEJP44fi1sJO9OPXsII2yNocaoSSGl0m8SuMKodmzr+Y4Gf8s
gljWMJdDxLLHPNKiDvaFsJt/HEFCIyPSRyyOgXS3UqEo6sxQGVq8uIFLaytdApEfOcIBTdPb2ssW
2JnPLDPQydyMM/irVUuVYjR8LBDQ9rpr97wWRYWf521frDxtrMgeZfza7/UJI6/CPcmxmSpFj8EC
QbtxnJqb5IibZ+hvzAp04b/0b3geisx2T7HfRIaN1b45mu1uCbMAvwvLRnQfOj8JHv2/UFMSpXQB
bQMBy462Qm26kfKhNR+rJcSxM/XoIUETVmlK6KsWeTE5UKOMFxyB3of1BOK/btyqIacDO2EJiQ7+
h2s5uOWuUL3ArNZ+5X3DP6c7vbhVUaqWBEEQv6FMnceN1/LF2wvME1jTde7fP1YVzHHmA/IeZBV9
060HhcAhDFfDsk4edeLqdvaYMmr/pqr/328uP5hd1IkCWRC9/zBd6n/1a6kpW47N4VX5jkgAw0pe
kiaxe1LHtGy7iayiTcwMXjTnUw8bZ7gxLNMx58xcshaQd7ArIZtbxIMZb2A84IeaaDk84/sS070g
aAt4lbI7YZSz4mh7DgVtcpAgHCRQhL6yeA/13SQZrSe4+ifjxiWex6CALXjP7sRA8yXUbNdSeY55
/tcbRjqpH/vZJnuOJjsEZ5ML1Bj/ULiY52HJWsficITh2L51ZheobLC6l6esUkivQfPSMgxke55X
KwMh1raYlXufZRCBqJfZRdUy+luCOt2oth10YapKN78n7x5L7tcFuOE9s2pQ/XJD2opPSzWrSZw2
CAh3AMi9c6PBnYgpR0LYNVO2xWn9+9wGgeKYuo5wBaRf6XAdIDSWQFTQgOqotWy8GR0/mDRQY9gr
nVDFQ67wHUh8t8L3e402a9pgaHaoy8cif3peu1iJw77sXquJuuG1wvx8zRJqt4K15FHNTibABMk6
T+mB+pqChT7JxwCytqC7kjMcTDNcCUOMxUNlaK8/1SEgTHW6d37v3UwUBNnmMfpZX+2eSDAwF7ii
UNqLhqnzGaBjLXvQts2vDMfoPIOb/neZkLgmx1hU9yR8VVMiK2B+3+N6CZP+zVj4Hv2DKPlVSj5B
WC7LSvlrxsWq6gDUQBTP4KJe6QMDSxXwwW5V2Kgb7pmqSSgNbHxaN9k4pDKRbxgmoo/Xt9pQcAH8
Rr7rUYqYgTx3EbU2z65PhyK7Lrs2EKJmtzvsJHdcziYFhaINhZg9acm8cIk5Lpafv2tj/VQrsc/c
R4wIrrP09TOnj5EnJdfE05+jE22A0r2pO/BlVI61vNTUbAA8nS09MG7KdbK+KWGCtwWv3tw+L0QY
uZh7U4PTMfUXsK8Dyi1jtEbavy2oFXRSQnL0r1xNSnu3iwf9RUIqOuTlQ3dkK1WuGLCBCIV7etWf
t769rorbzxYwJ9Oye4f4f5AlE4xEfw0Nm0IihprL5YX5EojohxusFZYXQYZmW5jL9b6kCnJhi5EW
EZ4K8uTaaet6oDNQOz97C0noDLSQPB9+rMkObgayhnPLRtdfovx6mE8fLWLeMlue+41/6F2mIta6
Qus+xTCL6X69sBw2E0squYxgM+mEn8fwBWW+YLZ+aeyPT7XyUtHNF/f5+Z4z3wVwYcRNF9KUoxhJ
qwkWGq9VvpAksv+4qYaet8Uufgr6Se0+MqG16Hpvd88AuNvl0NKUdbG1stl71jsWfZpT9QlMcbLZ
/sBKPF+fT5JZjjEMLrvgzyJ8sR+8qnP7RQ1kxi4mNlCYRombKy1TwBqSMmBlj8ivCvoxYDpmzjIt
pOW87+4fBNthHQgwF8GwipBJFvbmSOGMHlSwHBUuIoMWSgDa7R2sswA49h3Yl7YeqBLRlqBeM+Ut
Ov0262RyU6KIESyVkqr21McDxL9HiZSM6vX19nDrqKI3SHG6d0SDl1vSOb/djVrlYjlepqElErmm
tsdhyZ/7Ki5gn8HGteSNwSDJazwoHug9QDBcmu1uQxd7VnaxwfalS+VFPShdnQeHvLiiVLB7okx9
2hf9Ox2V+WN45xSLi5qnffGxKWiUoVXxjNmUq5g+bLdKoV6h6m7azCqKmHTOxpiA4JfVnnlTIR+f
wghVfDQ1AAFGWEs/aHiyWb2VlHCeQMEGyH7DIyPkvj2sgUk9fR9RN/ErZphDGn9UObCCaQOpjV7P
PwEL0iW27r/3+gAxq0Ga1rrTfS/6GZhgoZYhXwGcZip2ec+2IqDwxe57n4atlnSNX05KU6MvSsUc
t+a1p4p7+nGB20JKNHIt5CZd3y6J6hGePSB6WC78GBmeQ3uA0+EIwdsj+7l09cSOZ3+GTYUvc6fw
PRZf8ugond5N3F0nQPB6x4eLzrIMHecWQkMLm59XbaSpqH5xKx9DsjGbolDRz2ZVSjUJHBboGfir
fpWFrxdcHOClgOKKZ/KPBZpVY3N5vj1QeyY/xQfygjY7WbDjTJssylPC1HxsVyvpj9MZ5muxnK7D
CuqYA1HotoAxWCCRpbNP1QG3D8o02/VRGdvL4CA1Ujz8LwtgFZk8dUIsPFiLk9OqP7TJNac8GO7U
k5uck9cYXsSdDjsgK6gXMC2sTF1JHU2mBTsIvTG7ML6qhfz3vv5Sgw8ilIRbiPPVd44bMHsc7Etm
dswJjFLACBPk2Uxyou+3jMG3Yh/moMuWDOjI2aHX7u4uphi4NXsmJwhJB1Y/1ouheB0ZCgy8BdO/
3V2PhVuHaXAoGOpsdfsxOXq3oJv0eK/px7829gddWcuoli1k7+6m0BfdZti6RNcLDhIy3K52TjJ5
DQnVVtfxggcfKjRrCUR7KFq6hOyilkYQeyR6Kh8mNXocF6AYtN4REbgatvWtjU/BemX72OInqlwo
8moMDeRwUx5aWkIORaOpymutnl0XTvNEM8YucaVCoAYMrLESxsmYJel9JGuYoGhbz+49eGNgLCGI
eR7Hgi06tksyLZJA4nDoTYfyYa36b+JqA4sesGIIcqO/xtN6h+QFPsQgSOIHQKiFU7TZ4T7RVA0k
BKPaTB3JxMs09c9CRP0yu7+OliU/pYFn61XBHYR9mAsSr7BgwHVFKPUz6m+tkMyDxzhip+QyKsO4
LFAyfWKJEH9VuioUbqlXSk3ZHIN5GFiK7/QBR3vFlew7guAcRzh5rrJ0cZ7NUwXjw9MNEKeiAmS2
Vc/c/WhvWvYsktn3lXxycAuiYga/M4pGJpjTUIEpHlV3RjG/AdDb9ipzgcDxk6gvMH20OrKvxbFe
iVSWA50cGYmlsSnfUmxV5slFCeWeX990dGzDEoMujJ84Tjs/q30sVmEcSY9arpOAna0BJM5nFDYN
NyZRK2Rrzs3fXTYkyi13MMDaLFw0LHPbSTDqUutL0rOa7FI3KYegIruKKRwTogJJTZmPUVI5wQ6u
oGbuVYWCLlZyAIS1pWpmiDjSF9clhPYV6jYuwvOrvk/vYdFAmzloN4lYCDbnD1htlMZ8qxJJhdgz
IPwzgzophI6KeLaeJTPqFOxtTUijsBiwcrAYlxVZgvGPerWa+ujxlCAhsJoilaSn1Q7/+YxxY2Z6
Xt0cSZdDGY12s71m7YZvukYFxHZO3Cq+e/dd088uC36C6CnUeSKeUgtMN60wytuYH6thGaGEqKLL
TBAw6EmbxLg75AOFYRHlJD79RBUcIxpol/Q6op8daPJx8EoNyQkDGffZrH2M9OUJMinHNpTHYNg/
ir+rXtKreQ4jJJsTWL6ctlYSMp7KvkFy9c65d8aFCHE91Ry2N8BeAL888YD8ypne3x9fY271+pv5
9J0aOxBxJR/4pMjKTvF8phi1TU+glHYiutlzVlqIfjN20bZ10trdqzNpb+EQWhdpu1WH5AHS5zUw
/Pn7zyGgdq+nodYP7W3aJz4YOIE3U8ETctyZoYFeMKYXecBxVuJf0cixoizkDbXuxmV+K8Ti5wLd
usngqCcNAbJyd4+rI9mcC2c1ftCZKOsnqReu++WZKTj179L8Yx3z3u7u7y+GFy+ekDaRlZeLsv1m
GKHTSCdqNMiBlmINuheSCTfQWNCfOR4GsIDSv51G/sTH5ORRzeNqpjj6lz/ConVWs2a1c0pBBInu
186V5Sj10pFHDnuYxKvr+Xct17tKSx0TckI7VGwOigCXDi3RA7LsnWKbl34c8NNnymarY/awsIRh
wbuEjqBeBlJUXkvfZGktv4vG8xVz27KsZs5Nbqv/exlcS/pt6nyI09E5j6sxchpvaQFYp0ajBB3d
A2uF6Pui3C/PPRSfOLrtzS+/Ew7w5H6kbOZ8pswxRaGQyehk1EB6wH7OdubL4NiT4ZRv9r7ZYrxK
z53CAw5NnxUhxsEzi+RzZEa4TV+23hGuPFwhTz1yo40EQk0036BQ/qhXm0iVoiO/xZWroOycafKL
hpdD9lRxX7iLW56bbvoXUQlCekK0rs70e2Hot2vsx5gAnm5a25aG9EzKc5B4nuwGy2motGpSdkpL
IpWDxu9cDPKjrZ7LkmbMclxSJZU9qFDe3b7xu1oSJZ4+FgjvwQkFE/2SsP3cosN7F0gD+qv6H8HS
PKfIAazViJQRPgq48Nr9/ttLtCCBMBfJAoTp87BmhBLPuLj0xUzE6RAV0vmYaM8FZkE+73Qn7uIY
2bSNByW4gycVhIMPoJ/JvHRp8lhao65Bxwd6yHCvgiVEKc0gxQYzT8nw5ucMqYOGUcXfB8eHw/ls
gc51nfDT/yBwQAnLDWEbscGbggJU6NrGwqcPlKUpoxUJejaLgbpUOufleHgyOhM+upU8CdXIsfdN
r+W4qU4jGjWAaObe43VNrJe73DU6HHVh5ujrOVLXAoeP3YBmqEWFcP3y15HyyZJKD/dQR/Tko0ew
0ZPA7Jn8UNCR/HvLaJ86Vh0EC4mGK8yvv7yFWdtuQAfYqlsQlokA6BfYLr5mWD/zeZOcOCMwc7h4
cmjyq1jSdguyNPEbVfCs+Id1SExyRWCE8lx5/8BQWXYYP5V+U9xdMFDquaPbu6TviX0YfUzSLE3K
Lff07mhSQ3NelhCWEZTg36770RBQoePo9SPzRmXi702Elv4DGr8ImQ+eG8W3FwRJ8mbedD0PB2sg
oQ2PjfUAD3ZcnpgRmZdcKxQ1rPUs/TnjVbLbh4mAQCL/q1NandD0HKtYItXALs24nCnajDZsxNU1
1jrR8PiUNTyoFzwC9sMWW/dH1UE4zSsNmeIbfqY21p+I9zhKw5A5cXJTtzxxynJP3VmQ0k6essUv
aaeKPM2R2Gdx/1LSL/H8xz0bFhB2CzKWfB1HukFA3/VWxA/KZuWqyUzBQqPIsVjmJpJmNegZEsSH
qa/W8yaKY6E1X1f1pzhFlo3DzPhqb1J8eYnf0Kia29Kbfx7ZwQ4K1SnZXBWGUZF2ACNT40KEThTC
/BipAVp0630yJa6mINkWJDj5cdGVjPJvmJjch4uStYPJQH2MPRTzgNWIYMI0t+JnlrFRrWvQYc1b
064eVxxO7J/4JQH3orYbLY21CUQfsLPJxEHRRBDWG9c6++vjU2+lT+t3aiUuaIbZ4iPOJISJTbZQ
H/g9/FOpzQEuayNeyAJ/FnMCucasSqlHmmWbvltiD8qzJ2mnaIEBtdbef9Xp9doBfIgXilLFRG0a
xi9Yrrn+Y65QgTbqY7IExRY0I9JwkLqtI+BQQ3SFRzU2hI5TW1DmfMFJwNqa9R6tyKUj8ipu3i0I
StDo85DIF+yfkFaToQXI0KXQa5AyGZuyLnkwc20cD84Y72SWC6ZTQgJ/TG45ROmZlOTeQ8HvRrhH
s1L7NF4NG5CUtqQTskaO/J+WKDp6TEbHgkdm1IOBW38m4DHgCoQ6o6DJW/Wn4HEAqSPl7ZcpquDM
r+cY1oLepGaQ5ZzSc/SJ2xdhq0djkkPALaSGqqHXVBS6KfCKx8LJ+d/xrypYDOPVJfKdtnSmMyK/
0qr+mAW2pbYPnJULm3Q5BnfZuUUtZyvN2qwRjaTM7d5TY/zLcEmZ5FjgpkVULIqs7SxoGk9EUuUX
qUDcAKnujvrEK64rj4zrBH8y2k7GjuXUmugN6l5vIltYaMAmc2wmpp6dw4L33JrOHLR6Y6PK0ltW
6O/JCdDBrEa1sJ89ssbhEj2g3a3AGhoRnMT2bhGeEf39bdkvlUqxwLoes8Y1tulv51XwKjoHENpL
ORaGZwgMgKH52gDBOINXOgdAlLu/WckoXC76dKh2ez25fF3fBVHAPMVEwRFlutdWV+PQTux6Mzqt
DedyOIvSXW75VLqoUvJBAwMiw034+kR1cBT5OCAQM3KenRjXjjVzu0B84fxSPjdoWINmthRMo6bP
ovUSo2Kl+D960cJEVjdYbp6PUG88b7c4Cpcgprksgz8EOR6BCDVwbPVd7aUcZtbAHHMxrX1qNPpX
gEIHM8gNGWAtyWV9Fhtg1RT8m+eLb8r4uo6LSfJpAMFkwBtuWYBAjtQQ8jY844rlmNVOHBZm0bNZ
vJtqwAN3Sx4QsrH/ZD+tUu7tgvO9A1NnRu8Ubmlaz3rmsH2BOz/fSl0Lqdv45uMPGuA6Ra2vr/Zo
+gU5zYVcUb589mT/uB8g+wo93heQgpOP0wj/YgD1Sn+HrsZ2EznghI6hqWAnjjmF0FJwnBCKm+mj
NX3bNE2j7vnwrbTbjN0zyRADzF0afR13qbt1Tqyq3RZom/AKzpt1r3Em1WXQF9BWtQiLlSlYxYB9
X24EuVcP8BfEWj75IVYQzxcMkA8XwafeQXZzqyRUg3XwP5DbOjWcmM5WtyjMbVrK7z+yqdpqlNbB
AapHQ/O6HsZZGURPdpoFrDoBKmazBItK+DhwKkGgEwJnR3tGIIxq8JfdgxRwJ1uaI0nvT3VlbbYR
0OdDGxwGoCl2tXDAM6SpeJrX80iTYeK4R7B0yIxIeGT5JnR31BF5G0KCczKZkpiN5xMJ287mq7CS
GPd9v1kYISdY6jD7XkJuiKkUtaf8KFfNODgZdStCakTeQYZc8rgxNExayopCJVeZiTB+l5cA9el2
gvfRH0rgqr7xmlNGSo3s1tABpXTpw/oF4Ky3itp3Rz3/8IZkJa47/MXKS+7gYjli3yx0TogQqnNM
FA73g7N7evnE+CUpNfTSKCURVNwC8rSMBmLzIFBsuJ6p7Wwe1Kf4W3EY9EFp8HakFIyXbL3/myKf
aYVRvd5GRC34RBRNSPmwZzhAarxLg1j9+K0CluPzOv0XgAOzOxbCcpDZ+38xH1lHE4dryjBpu3q0
BCDorQSFarNbE/rKEuY5LqWDW82HzvYgia/sGlIG/Xs/wWOTP/O/6fhcNUxoJvI4NvZNc714Mi0e
oJhS12USJ5aGWAvxfTD2Ap/8u7ze5/9U/ttgwfjde2w/KHZJWMdl64nHt3t34MIYsmk4d0h/uGX0
QnIGL6uxI23L0XKx5p96cG6cj+WXvjX2TCpA8I0I81erI7Qg4bPANc3EhDKyy8nGcylfycK0fGNc
k3tSvg82fWO0l2azP4rcXMM+FOHTgaXl5AoGimiRcjVRd/Rwe537N9ku+zcxT0Lsa/m1yx5uTwYC
SVGT/5JvV2KoqRedwtL5xMXo7ri67KEyfCkFJ7EcR4sLjwFD6cW7Hk7ghxWKnkxyhfmb3L2tzbLf
M9CdbFILj2LRHzrSM7XgIY76lKmV7tsPsS31sYdfYGG9Aa6CpRtFVVKsOh24Dzc/eNAQacqsvrK3
fNEOISs7A4LyeHlyMaVP/5y+ySZzIruE5SWbFd/DK9kXDawnzon0GUKf54wnawFdIMELXKa0a9Cb
yP8JQ+75jgWPDjmqMlHGWLD+oGw7uLM7nZkloOdA4tuadC2rEEdhKg9xUu9cxDoZYklQqzMqM7Gy
fC8I0G9rOIg419mvV84GKVwMiLX6P0U5PfRWteyfPVyZfxDcfMUDK3RvCwEisnAwotCLwIpgZ8Mo
5utqc0wj2lTerlnGt+ZYAcXqlyuOy/3CFjSuaeV+6/1lrtpvig67FbgxyIg+VNMtesdXdjd0W+Go
RVAyuldfTNLOTQ5uMkeUyTEkStxAvtfSwa+elo2Uo8nK5Fen4Kiu0tidx1GPXV2xH2KbJIbhR95B
/LZyr9z3ntrR1wxGotJjGEMqpWNz5n0OsYbpvN8kMDx8rHtqm3njWkt6VBZlCq2cezeZ64H7ldPC
+SfifS6aJpz1AdzFontxaWlDqcWnI1V//jvIDGoCwtLTo2vbBmTt6R1YA+n+KbV3kuiD8FQaQ7dW
hYEBj0lvfMZlIx3r7KV7dd9YXITcKX6UMRcj1fbD9QFlHUQ++9qNpBSHSCengITNWde8u3qWfQlP
uNFhvalrZyMFQocsiFY0IQvFRJ6ju9/tWnfRe02WnRVrQRi9MC8K8q//6ExZh1iZI2lgjIviVDP7
6bpuNebHWHj+oaIF/TuXZMh4HSgbMBG0FxH/NIsBypDSv6AS6n/BP7cb+xrL5RThz+pC+1oT3cGI
R+Ul0yF96G4Ep9gl3rvLdUDjPsI03ov+rXI1EpL6c4g2eX+CJQWz0mQB14+o3ukzlf10tjVk5WAp
9WCkD1xY/13nX4sGUL0j9IimVJw5CSbCDrDKLNd3IHadzfi0l2e04Myd3Jkx+jhHTHV01WizuJZd
7xSGpKDnn3sCeFx78+q4S5lLEW8XPYfd/HqX3NRJ3rLy9Pv8lYhsylYcW01gVXayJD1x72i8AgxU
NFELltmoCHIeWJhQ2NdZaBw/uRq7p20+ZWHwJZ2puR7eB0W0NDklHuOnRZNhuYu4HCa95w67U+Tj
UO5DuM3N5zW+g8p182l+TkKcZuqRsGA5qVnSIaYlIwwJRK0WJV2Wy3KgUCSx3a9yOzWkSXqlXQax
7G4ED+aLPeT9NzJJdc5tj7okRFFcgSvKSRi8D8yIkdFImLbxzh5+gEUAabDzt2mZFwKAUj3afRbF
5c86cEoo1/I8W5scT3Ubr3MdUoIgBfNyY4dt5814Lwp3RIunSUjTAtCtbIrfsmLeNLNDzQfxsDhe
XWVuTL2IecQycY1+JHO2/IDo3X5Qkon4jFKFDIHyd5Lwlv6fJ7lX/WAs7sZsnJfEQbMvrrVc3l+8
Z906BNPXYbWSCzstGktk9keJpPmLeN+IKwBYcyg5Kg6h3U48W4Qcc34+D6FjpdgJMBFu0nqeQZ01
DMgv4m2dAiSsMEWaVuw+6bh2DO8/2EmA7PY6xSwsQBk90xEj42fIsnVu5clQzfs0nGezMljYaBzb
3uKVqordYU54dK/QNcaULwoe9YKDG+CzE+qGYGlScoeRscKkhHwdhhEuK1zACQ7/sW4oZwBwQZki
/tT8I4IjZRpVHAhdOX8eepa/EFIQiSHI/2F6Qpb56snfsk6naZwqNknPzplqw0gqbOab42ttj6cc
YUl1hF1c/hKyrNToiPjP7NbD1NXX8IMYI2uCSlsCn4BCuWPgcjL/BOf1iz5k8JfMtCG3D6WhH8Mk
lRDMB+wOOfz+j3ArBONI4uFoQsddlHNWa8xUQ37aLLwUpn52Ewo0U1wZAjUAWNAUNffou0SZ9XBt
jrzwXN7iqlK60RGCslh8Kwj2NxgxBZn/0XCRnykzgCffs/CdtYAcTBPqrWkvKacG5gg124Pe0aHG
8S7FBGXWGJw63lllYLgczJ2VD1ltFR3vBfRESfNRSwFP+T3HgTlDRZSoX1isGojGse/xxDMDOHwG
GdLkXw8dEgWW+gZvoo8QaADsYSlzhRdHJ4VDbsA/f6QNhi9bYMgZFVTwoCA+gN5nliUfEMC5EzkB
lHDlXB4sr1hwkr/L3QZ/7jZxokVi1Fu+XoOnksJ0Eqq1Ee8SXHakulNsOEpQ3v9vapLV4pPQeeKe
yEGEMh+eYo9InsBBZAeKg+VIF3oW9cPPSNczrxKgiepFjc7A8v6ePKWf/nRwx2991/wQPzRRmh80
uFEfnHY2YE8uDjLKtU9TgG8TIryzeKZpQr0t71ZUL0+/RTk2dGSD/qb3LA1cppu5NDVI5+a4SAL7
/wAzGHJLa6VH4ZuuNXbO4gCMJP/CkqeIztO+V/513daUz0PuxoKbZgwzHaQ0wqMWgyaSJ8kMFzDu
/pTEbVYKXcD4CMpmcEe7q9GqiuaiqhIWzyDMXuhG6atqMReMoAIgarGrmju7suV5R00q2azCzvLw
oagPh01x6g8BXltN2Br3QzJtigAJHcPUENJ9bBHnSr+R8WAXcvWsq/GfMX4idw7zS/0NOZ30Q2Gc
MlMZBARqd1ISQnzMuGltQNsnkx0QI07By2Df85Kl4ndhSOcbHxsohYuby0qKj8E/QDtx9nQFZY1p
/xK38P3cF32t75+Fv103PRUyT6VqtY/ses9NI/UC95LkwI3nsNhhLp7gr+Jx+MPasMAHng1cltYI
6Jn3Uwopj13DFqn8bqZvuieWqxDU681BeQWSOni7Innzki/csVSvbzFR9ct5RC6IVtCOiZJaOsLl
a8iPC+4bUsdbrNqbt1vKm3iX+WsDGIj/RJWGf6ntdkmggphVp3EKP+0Kyq7QwsVjprnqGOWEPKZu
CZr3fnrX6a6KRVZQbBXOdW+jqeg1m/lcQb3UonAmImf68YFVkKkyAq8dZEV49zNCYoYpxoh9hfL6
gZWc15r4FR/WLeQaPl0SPrd2nqGRhSrNxSrmkKYBkawwHVKlVU8FlV6hKuUBlaeqn7fXbz/c6Cn6
eHkaArmBw9vcwZ0GU9ptitrjWS+UPmQ/RcHyGY6eGJH2u+GUi39LzocFWJToSgjPMpueI70vRLiX
xI1xzjRkG7rrEu3yBsJc+2i6D84tmZ2Y3Y7ksCmBFzxwnh2/VxDk/nXg7RpTn4PMu0SQTSOXxbDx
6/pfqTE8P87lW4q6qIfgXcH39W1t32uIGrzfbg3+Bibu+M3FIrWY+nH32V1s6Cb1E72kQ81t7ram
nplxmM7PBkTaoWWMjSHaGbJ7+BSx0two7c47XjfWzRMjKbRug0PyRvBCgsilQof5I2JlXVj0P8qE
3AeTkDcLJmtscTz7H8+QlCJBFek6BsEzrsrA8NCHaBnjEyiRY1dtaDh1iyD1ww1ysAl6tLiDGZSr
q14mrS7pHmcqn2gX0IezajgS6uCExncoq9edex0f4jbMZm3VMOfl3Yqi6TXqIqdpMFeyliVzZt6A
r7lJFDkuM7+QlNjjlQ1cGk7Av8mb3I67FnHnKPAGZKSQc88pqaOytSwG6OKqhaeIDnyUTBCKig1N
yAUMkKgancQcDr9QbrZdIiGjP2mEU14qfReEr1K7rE1iPkmFGytZQpkeMc7Orv8cV3veVIzDAOJ2
23Lkmi3W+KhDkXhxRxE7gSV2RzeAMwRvkLLiLN2WvQi1VWT+4PuHg58O/QULIxiQELe9zJ7+vdbW
DPrqWW3tkck8/zMiUzQuegHN9IqzcJ05J93ZXFRKVxMcsdXTrxYmmPlv4GPsDPMt+OpUPKDwamog
W6/ar50lE4Z88Jl+T8i7ZimPT8FC4Ir3mKSgz1NopINNZurDRMcw06wT1a+CpbrTSvmdulf7b02R
zs2sdVRgaaE1MDaQGH5wY/1UhBYCPhXHM56lDb+/f/ATYamwAFYPazV404h3in9QNyisVPKvJ3ab
aXOafF7opLhJBrUePMEqoSumisAqzHASn3Gt2Ef6wofM2ASXYQKW+M4Wm35fu+hvi70D1rFe3cL+
UhcQBuHh7C8/FA/x0eEwCDqkzTY/22zUVBnYBaeomc4czIL7dguxSJgY/lDIdUDmCwWZkgpOf9RH
pM9mFwdOYREh4d3qTm06zfsECbdDG9AtkBWBmgqmXelZgX5rbyeAVD6tkO74lHFXNq/MwXNUL4tS
P9dVKn/Bh94LVhwiTOLRLZ2MsPUpTMyKzVEqImC/2NU4P+XLGyQ10cFr/MJg5NyDTLZD8qn9ZQmI
MIp4E0c4A02QvchJ9KwwdJ/V+Bpn4yQc6yYfJUVa/0lIUUoOc5EcvueSlJir+6v+eIPyyegT+ZcD
TjtneQWFk1HWEb7/CW7aCNpkXRp0bu2HKSmRBbrQisNMRsdwQWixbME+kY8ep/hhLiy22DnHpafL
CIEs8lohIOaPKRGeUvQlrCoZLGOR70xImD7ZF8aABlKzuF/rg5DNrlcUJgeT0rB0UDBxWYitWdWN
kWx+omo/PZvS8h8C+Ab4t2zNXyiUlkKrzek6U15wt+iUOkPgRNUBE1M/6wWp3Vm21CvrMOXrWS+w
BkI66MdQ73ftKWpj9vZpLgTDMTV+3lUHCG2YABaurhb0AIfU3w8BmBcV1MwRaXva7KTgYDLuKTL2
gYTHMp8mcRR5/iPmzNUcHlkU4c9xn7apx12QMxNA6DJOdxW+wIMhC1XzZiIzVwjK/aPx9fA4sq8E
8OfygeP7hI0SyK6CcRJU0fIXqMvnyIZUG2s97jtbKqWpJv/9Wpy+n+rLOh0KIyFKTiyD+oU9l8Et
mLeqqvkVu4cFB8CfZgN6l3QxfgWP+LyMyS1PV5kMCOOVbNdQE1eNsPDRFJVfGYcPrecTJXcJRQzb
wmf3AZLeWm9PN9BHb453Mxr2/tf32/YbZNmavopDA/d8EkJpFnqno4vrr1jF9C9liZCmv5mZ5lRc
zv/P0npM9LtLD42DiUm2kJlE2W31Mp8nEmspL5AxCtQIbbVp8D081j5q//TzP0to+PDymjFmjRzQ
kfffL+vyZU7bbNYtSLLC3pt3nbo4FipDG2JhU+X4smsU/qw6C5NGzvyIbPGaAa/2TRht4xz7wy8M
W7JdJDG4jkwhhXpDi1M4sVwdiuJzv8URaS8m367126xjb1sj6sxqwFVjgOByAyLxy/+J8Syg4dz0
LjilF9+meR//kkpLY3h02yqkBQvMzGLamjvbVOXpJPAMOrWZU1JdNo1geDmqsV04/y/FbGAHBy+T
DQb+YDS33EjKJa7X6lNUJLZSbb2+jYu+vLbCYGZ49VmpzE483G5tsOjXd6OgjCD9LmA4hqvrreiP
VGKVSdHp47zSs96k4rvwxL0rpVglQxjO6pZYQArfIoW6GBKMj6Y3ZcdDpxGU8q5qKwC9zgur4p/P
g5spG6ZwEsqI54uRgIpvCi6gEJfPWRKy8CxSEvvQJ9EpMbS+yWk0Gk+EYb0PbCpTTFi+I+gxG29U
fQc2F+0qDa3nsMT7fgdjRDrkTPi9zBOOlUvKVIe9LEzdlXCeTG8lggetz0bH3S3ZXV0KE6Xx3CL7
1+CJaMAkno6uyBE6OkzhNz0wPbZannb2JXasECOODq2mZWG6Higs8DUIyqx1x1gQDBIwM3lBUpZB
e69zKkbJUC6YJ2s/z+Dc4ENMnbNMRSgPIZvO3O9ZeveNicAHYoQNUiU5YL0guA00kAu/yAPi8Q7Z
4AH1/WClIJg6hUe0yG0iYyAIWX0f1PTAbW24/GIkXY2Knnmef1akxOpGi8xtlb4Gaer+five1p7t
iOWOpMTkzNY0UmC3thSjpOB0GyHc2iF53RWFIvo5KcCofY5Ir61pXajS6eZyX15roJ+7P9XivZ4j
rfn0ClB4Yyvi/DanNWHleKQ8ehuspy5k0Ri/aUiE5BL9TGuRJHCnY6s2TODTTiXUf5lTWsBig8Xh
keJi/XNCPXEZpTjnbDmTALuXOKjpmeK21RZhP8mHTdmfCEC6Z6BDWg9YACiaSkNfKoZSEDT8CQEo
h1DQ9DssldXT64TyyZu+gZy+0P6dARIfQByFI7QD606gK/LBKOxJ1SEQ9N5wjQhilXmy4WOwjBTq
DM3u1/skqdyFfMkSbiRyZBpBy/SKr/8COGAVBGCxIl8Lfev8S3tdd72+90br94YdsyRGwwtzkz8q
o3rb4ztz7K+EM/mPF5bO14RGmgM2hOwedhS0qHTSVpGDYVkYxsS6qqHpjEYkNV9R5hsPQzk62hmd
4Zer2KvH3tvHRZfgoAjgsD19PKKfPsGCsE/4cBT4QPhWT740ceAVsQ7RqH1ds8AgCLPFWFtM+hmB
WRkncGfaxlCHCifCAgUjinvtZ3McUekCYTd/YL9DI9SwPWxN2Vs1oQW4szYGbu2bBtkKg/pVQIwo
Rfrd6H3VPU1YcEFX5Z7sHr1C0qdOq366mtHrXdSryZ7OazfJ72oKGjbHdMPl5/og34bovYKHkq/C
GFhdXccuG4IxP+0WkhxLxA89szZGD40dgzhyxihWNv+4Cl1JK1jZ+Z5KI5+fD8/1Ix8s7BSb/yw8
f5oZ7sR+f/SrlWJmef2ySUc+c51Bx1Fjv6gFiyup5XRsdYH+k8XhLfoVTK3l5sOzoj4KwYbDPl0H
3edumzjO7vuRqONO19ZiYO8FonQ1tkbSIccjAGTYUyfnRyneN/4VkCiSBValtg7Y9KkYPRlLECYl
fMi6K/bQqEemnVMM2GeRJEKMLNQDDggqe886PNzwzBrU1gtei9+xyOOxwhFiC2Lzq1/ezDqP+NNr
OIrg/KcQeslgaEOL0VH7vKrLSnSg9T0WyxWiC9T8X9HaIOOgnQlZK+u7oWStZz9ynq39NyKAQSa4
BEJwEVBqoq89SxI25zMbr+AUq1LsB+bxfoXCjX5ApU6cOF8+5C+7i7mXeiuDkcKL5D5Xg3OcGfDB
Rz0cMeD9JufcsT9KWwVPUCfwlRE9mwVc9LHckvHNqFyh8ELtkZ6XXimIHu4Y1jNLgtrIxg61L6lD
y3dRwL0lr7yPc6ulJtJSFWd937xmW9+Qaw+z6pwLYWZ2avnci6WsxF53PkLPz3vQ/5aHOB5sALVk
JXKhHPM6FeOkBpSppqUvTUjPkmMeQOv5yJo7fy5rD/Ai33jzxE7WJiBXeWcWYxWTWylkTToWRD7s
r/oqzKaNXMnUHwyrD9ASA99j8qQ0k/04fcvoX8YH+8VqAblChhfH7xITcYdlfLwAXQwLDaAp8FUc
L+5Dd2GOmNtH0n1vCce+Tgrt3qEI/3/bSUXY4PRT0IiTcJHDBnrpgMbd19L1XK5EXampPJi2eiED
CHlGiUohViBXpuuismjDv5UJm3+In/Qare9uoRBbnAqLuRRmI+EGDhm3y5f1NHyOpsm+64Tdo6iD
9FieJMbsCONQLkHg0F/WJW32fIAK88gdfX5AGJVPnyEw9wRfAyBCZqDYUlVUzRjxdjhbgPjQHCWD
GkPfqF7HbJKIVVnjhbPRMAfFni2JiNuTmbC3nWzoEADlQMYqqGXV8x/epdj5X/CPAzqGMwpJNyn8
MoB3j6cAj7N9cMOwE7vLE4c/CSW7JPtZXtPvyRwAHHcvoYec2HdXk6yHyZiqzXsQForBa3sBFEXc
tggBC0j8TTT4qHIIGtu9uB+3yXJXHNCkuaCOdxR1W4oSa/IMgyqV/wHEB7iZ7uw83aJc82wiXjtH
KgWLH2rYqYCM1dy5CEYtB508cIcF7vK2K3+KRGxBFY+gYJ/2WLbd/qCMyV7ksBXBcXudG0PGpGiB
6wc4KezxMzAZmYYIhvvvsrxvTIZQcIqsr6teWjbfEtEiXedpGxve2ZO+7srOfwNP/RnSzdXLRiAK
8DDYUIkUTdFrZb7ibGuFsXwjctyiM33ElBZNB8PtIXstkt0b/6gHUwPWduexK9SvlLmQ+5zWjj7S
YFg7RkDSPoDGLAiWylGl/SQgNxRAiZT3DaDWfA8rUryp2JKLrv0BzDV1V5ia2agTQ+jmjRwQ+tR+
Dr0DqQ5OlCi8yKWDvIw7T8GtrZeSaxpho52+Aon9WcTDP4L5qYTLJWJAq+DIHvbvC/E1ryyUPqCW
CGEwUDkCEaN51HCSQ3ggkyJYBPh+9lLtXPaDU7IA+Ht3cGCd9ogZP7z5wbfKxJkS1fCPExjjfeyI
zeyMS1Ywj4i11kxjZxNtxpzAHyafD5ksbUR8ogMLtYHGQwxADXYxMEl9iV0tYuvxeL9vVJPT+VDX
bLuuMDglO+5XtflG8iv+/hs148Nk3yvbLVBTJok6HV7F50zQyV6PMkMaQ87s2JEyRh8KzFvuDmZm
u3l4+gpOWMCynMwU4xiEVBNMOlvcwewjKD9CWtxrys7SExmiarTeHjFDPHW2aJ8hEoQE853b2yLE
Hh0ojkqEwV49zsFiFe5BX5p9B9+6mwat/x5LCCD0gNAZP3XmChDNwns+pAilcFazjlHAPmXynybc
+jw8f6kDngRilc+1swYiaosZDMB873s8fNtEluBCsZ+HR8ZUh00WbcJOLSrcLc54JXGWe2N2nqQT
PFRqv+j8KvSh65ILceG9tITurViSyNN1oypBakyYJmLuH4EqwC8ovvyNn4k9r4DRw0/9U/2D9x8t
Li3uA6jV9+ENxrzMAi0j0sIhNJn9SdS0mm1UZdNSxSJNjUpQXw8IMtnIfKf9fJe4pDR5iIaw4Sey
uNU5Y54tXocbaBsojhqx3Pny+Fj91Ra6rfOrFLY9LTFg1vbTznMOATkJ7niKHhE52JgIeRsZ6dN0
o5nIqOaSK+yRs+3L1sfcMyJKV1gVlrlru2f3yh3Ey2ONK0quBgR0hZ8t4Ony9i/BdHIuLJ7sYVxA
8S14Ep2hw3J55bWEEL9YQ8Sq4+UW+O+1l6d5k70mFoFFtkWV0SKOWNNVoISb9FaQTscVpNTuAum5
eprVOltIr9MAXoTcfkMmjlEmy5UmGlTxWHRS4uUSNz8oKIjic8IXd4qjNWNzINf32tWvfIhVLYSi
wg1rZgzYd5//owLWvST6JzFjpZadYuDifSRL1Sb/uBP8jMfAWtsceFBCDHl8JO7PtKcesxITj4qg
tB5pzNaTsyJSDOqJxU5C9qx8dqDI0kAeF66am2szar5vRGSIS4q729am3/fdrxeZSL4KDWnoO+nq
6O+oBJ3Td4OWumAZNiMFhfcChO7GaqtVR51a6B9RptygnLyEBLXqKhSDEc+uXWeOt4EfCEvkotOf
VdsLDIE49xUXqxKgdD//M2qNwA7cfJT012rMfIm4DsyAnAx/bjnuc+q3jD/nqcTb0gGR/vkONZtH
bltoBd2+6/YFoTpiqVpSmNes0Bof/c2ovnwGi2IYabT4cGithufPIsuGpubjIBP3wOmyHXNQFJOV
Swbo1oNi+kelmhzM/tJFQ4EU7IDBm0QgOqw7JKlgeu3A7CaTZYdqa0bmXcc2ilu4ozt2Khu0A95I
zx3bGfe60GWlW9Y1pcCP3EK01dVxthPnxyAQJzPgvISo/CSB3YZV5MgqJ4J3mJ1A2hTXJ8zdcKLo
Mdput3V7uAJwjoqinLJIGDpks6nyhmEKYAASpoI4gtpyKN+DJa7yJPSUAznIhlEryFlSAGn4Uuj5
eDbFvFLNQCj5bcxaJs3my0nnH4sLPgwgWQRL3QQtTvMp397Xw/sSpue9hv1jRWye/JTZOZiXI41X
rwf6oq60USjGY9Rb5JZRiQvnePR/mK//aMpulp8GRSODJldpn1lBLqO1VWXthrzNiKV09/agxTf5
rhZtJ/KML+snM4MTnCkL94GR4QvluWFWrrzsl/wR/IcMlAuyR1yFNJE5z4XCugWV87PyAMGGP7fv
9w8OLXvz33aCV/YEmbsRKD57GI1I8F3f1+t+E8JhzFl8FOdT+6C0YKwGEyahAtiMFUePZb11Dwzn
lLzSqgjF0ESf5EY/0UyJotlcIszvufSSr3CIexfPi66zPKOs/GCoTHpaEJn100Ms/j4d6lNZFccc
hERHWBViYVS7K9phu+v4dIVbLfgr8QEarK7QWmMpasCPumEipdbOssAUrB7iruc+pc7DW85wOm4E
bKs0RF1t/2QvDzL/+K/zh7vYcI9YUgxQUxFennZStQQCw++UcK3ihbvCfSOYxf58wsj9SRjqUx1s
T8WCDtIXtdBu9QIOh8BKUTJPLpHqI7MO5wlgJXtVO0V9ZaEAs64HwQLDM2stLsW2wb2SAShleU6l
RBuJIeURq2uKOZFmu/1dQOI8WoV9WvgAqnhtAFde8U21qXhd2ReO3Udt2OjwHNfTPJzvsY7wA5Iy
BXeX3We8nrpVwuEn5gUsk/yyitV5G7ts5t9RlYzyfCBF2ybm1/p9/WH/I9HrxjljmczMxr2SIP4b
iBYwniDiiPw+6cRzITc5xBoua/AGuEDiXYKRLrkbrjaCLw0X9RF69vSCUeQ+IcmUHgvj2FqIFROP
r92DwIKA76h+yNFAraPHzREQ/S0iHvu7KmMQPXtEzBfv/m8uRTyfj+qcIdZ96VXmQlQj/6WLPOPg
9FtoVm0xMreJoRxnDsHqJs0OvjlbWhyUGJQjvCTLNjzYFJp3St19KvBCcTgQtLidOpW3Xobevill
Yx+SL8ZD/I8xV0dPaSdP3hnbNpqDIzUxiQtF/AhHchpCaxVcTz9oFMofjwE+9prJeUhnRQ2z7VR+
r4pmJv2vStuwc49O3z5mi82Isz8fFM3nIyqOICJInlgejDJHN6NfGdSiz5KdY3C8RW0vrLYox59z
Ki6QZ2GaCLzRKWAsfqOnqwKtQMnKIFF3P86hN388NsOmNnH2wKZ6wnhUQ0lwLgLPyfnAU0PiG5JH
OSrKlHPvQMFJ68bZKovuG+B1c8S9esLcpN8dNjXIgtsSyp3MBzN+okq2slCEUeHeAxk3lrFRHUto
/7PmdJ6gk/ihn8hmH+sXH4cE3zRNcY479WuuLEFTTiiy92/GQd5khReQF/J5yg5jQQ4S3hpVPgUI
LpNukUvB9a7Xd+1CMCrzjo2KjHa7M8uyyJ+at9tiLuOiNvjBjlBJ2hX177w2IT4lIzk22I/RLBiz
S66VIlm1oPghigWO7qj0UzDxrwsFTKDYVP3JN3rBa1COUgEHyyspEMlKiakibcx8JHkC5JKKDaBe
Qkn+KZ8liemg6uhuocO3UY1JTibfWmxOoxiSOrvvsNE/6c/BqKqfGKTMXPqKTGV2dGijcsWJG+tN
PXlYTk47J9HOYPFTx2Yx+kJKlA+vrts4chYk6EUn0b7J2cs1qrcu/k7PvveJHquB1TttG1wA9/WF
2AwmQnVpvXKcXYy3v1SWfxpY6ZuYJN7SALaea3UomSwIuEUACU/d5gG8ZFVPKJWthqI9DFPOQF5c
jwFWOw3NLh7TahtxNCJwWce3ciXR+YnHhc7JAbocQATA5dG/s1ll9JevEfdeN4dTnlXpH+Go3T1R
METKzVexjIdX/ndaeb5JkgqmXLna0t2ea7zxnR7gq1PgRQdP46joEmO3PHkkesMNfPA0/CAMFnbb
WvQQHsbbnhu9jPyMEwvdXR8P1q08svab7X5F53RYGHggmHTX7SXgZuzJFr7mA+cdpt+oGeH6quAK
26W8AsZqPf5Nsk4QvsxQzSbAiBqMaeVW0lqicFkwmA+bjwMfEMo+ljie/ws2N1+P9KIQA3C3GXdJ
wBqv74WqO2/eDbiEZMa4bSJthv1aLJ9fcMxTlLY7hRH4lk2i7HFguWjWoBGABZEUimVmXSEeczaF
9ihbY2/sZL9zmGUMDgxkQ+8FQOXuBErOM+rrLdzB+oECLWuVeVrTHmBU96NlrFDojLasCJmgN4hb
nMGTyXgiUuhQrA1OhfR5em7V8IuGm+iWuS7ait5NY06xl8wYSUf0CxNuaAPWWuR6SNPeV3vLC0F1
NJbM+YKJ/duLYHPG07mSgOJK/8KxXJ8kyyCABQgh4P8KyG6Q0LHK6N+3Of4ABnVwzRyYOGmwDHUZ
hUI9/O2S1aSF5jy/i0dJzbvTS8Hv78YLSsgrpKrFsoRfRaW4a7A+hdAvVat7E/2krvdd/CRn2xE5
WIK/mPRX9v+Lsj3KFWLHj+9VTNW3kGZ59TMdh7fpXnZcCbTkuB/m3Fryy6RJgywXBWg5dvOSKuvh
YBrE3LDRkaHCkkJM+EI59UdH4R3Oj2VdbBldEFe4wa3vH8d9Os2IjiSoVcGYb5jcNPwRNBBUDsSl
N8xHPMttZVIvn432J0BrDSk6k3W4Nvby/DDoKlsx2hkkew+xh32CmZ5/8sB1Mmmp3w2ZP94PEMR4
zN+kNWfLO2eh4zJ0UkLUvcR5tAAY2KcKf96k1HBEEcphg21m8vZyUP2QxJ+sQH2Dgu8AaD3U3PbN
DH+74m3hYK/aiLPrSlyMdSK0lo8Ty29qsCFy8cPYjk/OrbHgXTV+36n/9uBMwakchor1+m+4mWDt
c9Qamx2cAu3KZdMjtKU2aqxCD+SectTQB/91q2c+GoJxN46bOziCU6yuJlueszfq92kLwCcvqwTC
Ufoxks+3u41j2FWf2l8j1c4FjuB6U2OaS4crT/o80fGW2kJZULhdl2X8Ek20UbnRejLld2Z7C4vO
oMDDmyv0NAXJKbyPYtD8Ckjjtgw8FgAAA5UrDou1Q9XjLS1voYZKL7BWSB5eZhz/DekZdlAdDdIv
zBICY3H9KHb8PUJJviNRU8Kpec1VMn/RtZkIOIxzxNnrlPF8T1wKrTYv2j/xCspb1u+SnoxjdcQG
iM9q0EDfcotXBOI+Ah21gW5QemNiOVIJZ6iWPODBllwS/3FE4K8n/4RMQNez3kfdHFf/HV79+Pak
L7UUewk6sa9JcoNAlKmdOw83prMylPREYxsQkG+iVyRVTMPODIzB6SPHh5GuVQGl98wIWs65U9LK
th3Da0xaDLo84t70wuRWMY1zV9zlkNxXttSCvu9GkWKGhn+zRbT01O60B+CoChRG0ZQZAtQVDTHI
7eD59ZCsUdLOZ/Ir2oW+3Czum6LTgkvO6PUVLKnnIBqXAZYd5yp1bt4RJiaC4CiEPg1b7KFZ90Bz
zgGsIjKFBf1L1vufxwBN8SeSwl25n9QifeSxIIBi1qCkkYReiSgkrx7BDxCqMj9MmA80SoBAIP2Q
55r88aK6adP0Tz2GEatpp3q6eyeB0czmlJ5VyL+CIc2+x+jsJLscGzF6oeYa4RqpuChM2ETR6cKP
rQAilsp8mpcPqETBg5nxgpwV1F6zSrJPX7+WHGYxzPqVFSBAX0HwjmXh95lnqE+cQwLfzLL8KPVX
CYq8dSbNard7wkRme11SppmDvP4r8ubDolSRSQpPxgdZHLXPZmDCrWsF5YLlCPJYlnGginp9muhw
wrhjQLE6oM5df1U38gm37lEacNLhCz2PS3UsOoKO3sj+/IO8VG/d2Xypnv1V0CyqhBv822Z4wlgR
vxVThgn8v595LviTpkdm9IF+Th8FsI4Hlep4s6kk9h4bS8TXJzyi+9m7F4Wzk+NN1ohdHk3kFqS3
vaxlIDKVcl4uHNIPS+ViD7szE+oVjfEO8NCbEzWI21V+yN8LvF20JmcvKLXI/XKPL0O3mDiny4ut
99pMj9fkLfpy/l2SPIRS3Vl7SNQdp6C62KE3WFIjJcvQj2VaryMHMuIHQd5QfXWAp6CDy3tyj8rP
yr0hr/2RqGm6sneZnhRyLAaQaB3EmeOkJvgymoBgNiuLlFa7ZvOmup/IEQesyuxPT1DN5ugMtZAJ
pRIY/T0+89sQx9jYfPhIVG3BV/YRmCWKmnk4YztdeBmXeD2hBPf5qkP/4sAwlKS7hejkOust/ttt
NAA6YILUrxinVKBkrQKwdS3IlrmcGJA0y58HWfr8KPUyuseXS1ltyuTjuBRCgHDI5WV2VxQDgbKo
G3vC8VVH+xw0yo46+0MPkZKGwBg48gGqjUAod/BLNsAVx9YXuiXNVrdXoJyN+B5BLcgy80pZ/+dt
+MsLtPuvYfZmhHXs1hwIcrzS6YZZD04LPmyx/yzb3SYPBEjlhqdIVT91e3TpAcit6xd/2G+YBnV/
Y9At3HB+KWAk0IHt3f/yz2pcLQogojocHNswbGd7HXfRJ5/V3CqE7NORC8U2ADZx8W10S1teN/LW
vwvHLKSu27zvw5Mk/y9R8PXRx0aM1Qo2NKgdCOdjSW4p9gpLIhheZ8RLa8iwt4nhzhkLK8EAqJLa
HWaDLqTjeBMgEYNYAGqofvvojw/TQ4JC6jXcdPrOvuEMpMY5XswkxUu9tE6icRAbsUFnkzFAGV/D
bm5f/e+U5v+OLg3fBHekqLTUkly/be7JqMDm8G5bRePDAkC9+ynmA9s7nr9JDzoDOFs39IB9spUn
/mDEtABrD937P0VUK532pmMfuty37w2zjVCF3mbsf2JDCvTiiB89PmVHX7cbPtINIIUKnka281VC
q9CpU9zfLCWCxQ6JEwHcppwjvKceJ114+vCW9X4OaiuyepoPqldaBWpFh94dTH05s9bVBJi893Tq
PVH/8zY3RLYgylR7tWhBe/laJrJPBI7OeAyzppe80ecSK6XHe5OB5mKzSmhJiuDbyoi9vadB1b5p
1JUXrTG2iCoaZk8b2Q3bhq+xHYoSvU4X5UtSYc9k5O0JHJeE45+1XWfm3wGOV/HclOMf35Ed5DDZ
xOGYZMaZpslfkBug1dhaNhlzlj1DZrDtf4efu8WlmIElVztcJQG6PGjohubGPUvcYzwLmzuPLlEy
MRcni493eT0fpsJLOil/bhP951LvWhrU/8f4rjw8hxi8tnK8THayTlWTZg/+QoNfUugiNQrmQbXN
m9TmVP5rK52jx+IJUJ+2M8Cr3ZSQ8WRcVHiKtoFKaUSKdwTa6CwgK0IvtkaGDIP8w34RSqlPek37
BFGKrAsgrRt6Y08KOSGC3gT9BvV2ipmdX24BRwzhdehiSZ9zqkbRU8uR5VJBjStGdkDe2gZan5K9
yLjwC2z2OiqAQzXZ0QhAfOCk3Iy25JfToZGvVDr8wO0KWH3ziikBq9vWwpve8h8zS0sEH+NJvJDo
zGyKsllSqL7NlGOJ3CJIAibJoR/ib2vDvzYYfevPzeodHegGVNXtPdnPY9H8GDOk7bttxPwEC0vr
VNg2L14k69odRrNCcdwa1DB+RurSFE8kKv3TUEgMaeigvTzeHQbqRNIUiPS8O7VWHTBOoWsrPR4o
+7hcdbx4YdQ8cyMI5BsEIHy6/CzAu2wTpMNpboOZPNU1uHQrmMWMCENZjuinnDcnuGWEaNoOi/8M
v2dWKmLeqQaDV5Gtg2XeB7dZwuZph9hsgCesO8bzp/2xbvoSI4IQnUBi7LOGJQCl/P5ezBG2fAy+
MsSZ9qwkN8QSWMnN38hu9gzJqsXPt/2wCQuyIgVil2SEbZOUqcDmF12P6cAoDOwLSSgpzSGiHGlr
aneLVP/7QECbuhBiJmOjwO0+kblj2DLzdDOMdtn3OkAqUSeKypJ3xicyF3pZyrQmeYaSNTRhiaZ8
a7Vht+fwfJEA1AV7mQUi+xvckbGYFeFkwN2lfJPiW716Bm7xWwYUnQz3FJUonudO3oEXD2cfhdCm
swA1zh2R/eDdO5iKxewTgqCzZBeTIMhQvm5dMoOqGfrzdSpGMJZyS7FYDT/d0HX4k/CpMmPg/uNv
RXY9UH4jmSRhCmvHaTnxYuCwN9JAmUnX9/zr5EkGe0Fkc0QiKQZxkbYEWdKtOsISlXbcvf+DM3ky
Ux2T+4duBbI+7Tkl/4CkwEhMlg4ljtJiAAZZTHIvisia7/ywA+Vc4FUm4hQ097g75uBh/oS5XqK6
ACKZMGwZJY+XoDI6x1aLBEaGlGJu058nK6QtFdtyrt3v7/aJVeYILWp504qV3s1tskjfHH9b8r7A
2+rHyz3nNW1IT9QDyv42rlkZWHuXFJL/V8Y6Dpn7puqsC1jxQciKvML46pk9a13crXNbE+8SY6wz
qORMvsD4JNhRcOB5OzfnLuDtwLSyWFd43tAsjAflieEl7IRd99uCSEBG5EAklYZ8JBP3bjMGqS66
UONSgOQxEv4NF4R3nhGdLoEEXQmKvEi9mJZHTbt0j8fezEd1yE2md6DmaAcbgVqDOkebXjY9o7Aj
VIDrGl+nytyP0cJY44hyRPhdJ/JBPNIbNTg2Iqqsm3tcDf7F/IUPGz1tEjtYZbtJhG0rDt8xZlCT
gezZ+Al8oL6pCCzo5D+1HECL75aKU/AQDR0e+e/8bC36M2d4hN9gf2myG07riSfGfTq7E4DyK/C7
znQP8CjBoIMHpwb2Rwlnq0RlJtsIFqcFCIoKKfxsK72KoW10KlmigHDBO5rL01Z4dZlZ4lqfUyfl
BLgKR6WPm5urh9NaNlHgwISMQOSOW3jSok396JCRRjPK1sMA+Y9f6YjLRyxflRnHlQB+Dn3dKzxd
s8Hj9xbN5TgKnJwJfeKf3YRf3CO4lDJU4pV7yUCOoHiLm5OWaMYlIblmYYiy8LuKh3N8Lwr9mLHW
/wEPoOf4m3NFHl5TJ6aj+7xUVRFiAJiMbdXbX4smsw4qRoFFvgWFRKxSeV2WtVEL36D6UaeHhULM
3f8s8f0QU81mqFloEk9BQtOlBinxu4ymR69q+XcDRF047rsoaJut4I8wWrWHDOWS4nG9LfxIfOkd
IFlPnJnhl4iOcdCPbiLnGPvKWPhtBEo+Th2q0rKSxTNWF6W+BHHheueVYalixQjsWOI8Jrh01YTZ
DiVXu5Ej2eK+5pTvsm49iQhKRVj87RF/EMSJsd6a/aoIcHB/Vr2nxLHTphw3zrEOkiUrk9gafGZa
39shqvpZr+nrnhWgYQafdtwHGM5zpVFmLGAPjQUP3swhwrwi5CkAHikFM0vn7FoFDLTylZigoNd9
dkWN1aHPw/bdB1onuQdFj/msomGbYW90TPmyXhHgIDOl20ahTvSBPAIvXVbRoba/UbJV8MBKcn9/
v0TwR2O6QUwNqIsLZHVrXaVUa5FpuVWQnQHvyOM1woAbUIT1qrZwXaPtn0lnsoJ8VGEvwy5aWTHq
ut0ywvGjdKDJbWp5m7y4gFQeMicGWuv3DnvpYGGiYPRo+wx+rtEtNuLe9sUnrt2JAtNAKLQC+a3T
aDBWF+7JL+aLE2kQqmrgv0HAxDLTBCcmUdIqS5C/iuqFUdvwK5quUE8j9qiLjE7Umd8Obb2MbjzE
XSvwvkk/iTemiAzl9HMiEtDtqhWUcYxxhBK3yDdvooXmasyGmtS0YLHtIQo8nfGXzFY72QMHOwHv
gK6ZfP5eL4OUGyrR7UAmUo0otuVC/TXn6F1SHTu1jC8AdNszdRm51vlwVpwgqReNzvJVgSF/aZAo
uE6dYRWm+EiyJFdV03EXU70XAabND4GUjqXO4Ga42pI3M2HoEa3qUfb3PHMg5ZAByqhNJ4o35QBZ
mIoox/Z0yVwOsR1UGy6qWc5aMNgWcAQxqn2bbB67ZOMP3M5LfnkJtRBLyyNE/TZWUh6wOYTmLlDg
NKE0KnOYbXYgDwYjSay3hZiZ5g4bYGBfVoJO0V2IuuhZNSr61mENyjU6xd5+H/hlPuUhKGd+w0dR
Oya1RDc+51MA6Eu4ByWFXq8d+ntSbu+5nZG3QrzFtSaxeLUvJAaeVPJoVNMork1r0vJeXaVtwkE8
MIlb87/D+7jLBCZG5ELf7EgfPTCKbY12MRxIgG4/8EQ8rat56CL9MsJQHrmaaeLtIauKQXRnbmXY
VPn4WmLOzxTavw375gZImlnBbTyKOxSqNoXyfkAa8fMuraJ9pKMgQLNlx0/WNcMvjVXPxu78o/Dc
sPTMC60EmhBZiob270RQdfnd9qjTrYH5OAD87JNNoeKiAmE/lQ6OMh8BfXcSDpy9Psv9ztgzIIse
r0vtAI/kiGTOLGuqShWpYJIllJcku+m3+I5D8Eg4+QsyRJ3f6Nmvxr9Ohl+9bGfbaUwtWGKmbvPJ
dPpSpFS0QzUcqfydIuxiVY/MLa1Nm25oR/8UhLYW0CIvPIKqtpOULzBFXKmkK3goyOArHtMeU25T
tOW0GIfPwNpVA7Ph0d7/SHZcTzUZtX2P+5naogPCqfjXngpwVeEa7sa6/L0c+P1IB4x5k/X4xprT
ZXviNKD+4+KvjS8O5hxub3XNuyoOSdHmuEU1Z/62Be7o8eqyJgdSVHRi5+CiggO30cWndDOSCdD0
d+f6GA0MwBKngTpYF7iMFbYo1DlQDCxOVRC/S9h4ET+OWI4LNzySBKPAx+6i3p7PZuTz7cMv6X+G
ry4ITO+aTWF+fkphRFAmxSHC9Lz1aCLribxFzLkdfk6p2kLQz1GjEs5pX6sZs6Wm00ppodIysjth
l7+DmWkuj8dDCGWDcaIBunEexzf6MnQUHdbRgPSPc+jgSNVbv3TdVF/mBX5Y0CYNZJi5IOGnUub0
JdKMtzCFGKjlNWTf9A6YEHPWLYEHAX2DdxU2u9lu3Fa4pgPM1iwairaGujfhOROg3wnlcsg3gvR/
8mOMI3YgqmhrcgJMPCAiwj/jZ0CABcx6uB3pZcoiT55qjRZGmP73T1+iGBBfmbJAxiYICxmtfqNi
Zcl5v6onusLeq5AqN65IpJIGKRlqEhffXELgTa9WsoAgCki0X8G5TyakWh8S6T/8AeoON5Mjs2tO
91dUdBuqsTLkhAuU8jr/lN/YknsTs/gk32qj3gCBcaW/45Aiof5FtSQGf//wqh/7f7BLJEyeonuA
Ea4xJCkPG9aZVWrmVxM7axwy4u3bFiNGZmIH8NhNYYxLsorqigkE8riZgpG9LIVxmaZ/fQS6ESuP
iskXtF10uptXTiujWiS2cjfyJqn1LM7NP5IpQRo6RHfcY2TR5Lqts6a8mW4LhUwW54Af04JA/Qg0
cwEVDhB0tCzJ/emFliIbwLk6PMIhoNO465qGVbTRo2dwGCLhTkW6Lqw4BTBupebxyTaI8F+T25Eb
y2PPMbamiDP9cejq+k8GN79m1dvUkYk0Ct08TstnzIa4xXMcX6UCBmI3TJYOEljGZMQOEo/b+z52
df7SmZyyikjkUEcfSQ7H8gzggnfImWsZNuDFImuFPDfrJKEzD0VF+DSccE5K0/XAd3YCPn6Gz3Ft
cN2+Hh6Y7IMebT+noHXpkq6iVwuLY6k4CYmrhjimFAMcAzf6iNxJ+uKCmSJy59rg4eB6At7Q27Ec
E2yZq0CT2/KKq6qn/6xaF85RTPU/lKk8neG7rbqlueuV5KwJ8gG6J5ILvgwTVIiQ0I2pnR9zCz6O
NnsYgeAM7Jk66bxXDtw0bw7r3Biup3vi2/APV3ewVspvzT7lfKcLUq8taPbYi319fKl2QDlnH1iR
DGFqq50Erhfa75gUY1RFW45gD8U8vE7o14NKXJZnAidfd+ltoyaZgvba1BoumpEn5FSJEKpIafGU
zSyC4HYO2weHMi1ayV+IRXVEVTqrqyVR2wmHSBC6DsIVtq7gNwgvOQR3s25ogy3VR146r7SBNqJp
roV0Hg0PUl+gaA+f6Xd8sKx7gWo+sB5ZpvDHU2yGRysTPpIlOydx/2XtOv9IvkntHTLvz7bGEVv1
Uvl6i2ZL6pdgt1Dy6hGCROFXd+RB0NRd//mvyfcZqscR0sBDkveoCXgUdpdSf0NCgK4AbsWcC/Q2
i3BwB5qnDhMg1ymRjzCo9hup7zTJK9sFfUlLcT2A8yVXyDEqEps2RuHH2sLUtlnO3nt+qPIYcFAF
ko1zKjsXq0s0U04KBSkQWaZ4m2sP4rk15Eb2482xWKoAh27q3z4BKemnSgUKEtbVS9CpyjQrS1LZ
0Ib/+1q7kRmycjrA3uCj6fhYCEF8uxJ3tVdxoCxS0RadJDkLcAsMVpVeZ1pRHK9srVNYjgT8+uIb
0QNzvRhCPD14tMmRNq7BWUl8e0X/3UCL64xR9oIpjSuaY87HQv2d6fB3pckPdEsqEKomXN+9nK88
ZuYpudcoeozvcmvczrjJ7JOHz1IoxyiSsJGz4B03clqDLZ7Tx/ZS/kArq6Irm3Aqxw7ATPkP3U/w
CO6LCNCFHysUPd3YIcNn7RwlMj9rVNn8/U5uIegtV4XQgvwVnkHxZA2FYDdjDe8yFVsK4ysoWojw
geO69YR1p2fOdKy8vSoernHh5PEZX9z+YRaFSCU9a+llcq7LhNR0OnnrfELtNUJv5xHKJHotdk3j
jIc7CSnsvteL8IgiP5TF6dXFe5XnWDY4sfyh/2aMF7tKQ0oQsnt2NIf310LKNXWeu1+cGz0cCmFo
ME6amFJvNUPSofQXBvWxQBpVFxSCvHCiJsfj9dXAWaRt4o4+zrtrxj1IJKdDGt2ssN+LBBmZJeVT
xDYeq97c2qnsEP4Z0wVplUbMfeTaPjMeEskCIin2YPaVj5U6JEg87yN4H6fOOIh6dlG/A4kE28Eh
Gg6hq+cWk/8Hig4IS50QQaTURwXKRmDHYoYfko+V0Fiag+wI+gnq3n+QL+rh6hUVukPpcSVLMdgj
iz+/ngMJ85+EzipsVyEJxLr/9oPksYDdsT9WrMMWBEyyD3ST2790RdUOMUaZ9uxzaYg2g9W9GUjy
tE9SS6/X2nuHpM/JF3QYRj+oyFP6AMCUdKCTSjO1EOzdjJEhBEt2SzY6fTkaXEMeSLbVix0Yac6A
ZxOAHq+0jo9XPflHWVWgaWvSHj/noIxHak2DKhuueIZqPJnKC6Q9Sds2dfijOHWEtbgGS3plPlkq
RNJmf2uaAio+jrowUKCvDcZUamhy59egIWTDKh8D5siDT2InmZQjDG1K/B+9rSkQOzoURamzABGH
SZU96lLSLv92mfjdblYBLyliMLrV8QzoZgw+43mZkT3CmU+PqmAUm8NUjF1SSpe796oCph2zHeBb
pvMm4ZglN5HhUdBA9UnxVpDaXp0jjnPk1Hi54sVxKhrsnYY3EU+ycq7EK/T5EKvVSn4qTtTZNa0R
UqcD+rot93tgBKO0Tjb96nV1p9+RurIrayTxR8gtFZ/gJ/rIlh4MWvI+2eQTx3lhCltLvq8GlTC2
7AToM8D42UUmoY8Lf9pcv0AsGynAVV//9KKIn3pqpyYFQLp/e2KpGXu4P9QYNfN9Cq7gZBTnSdt2
ZDY1tXPBovUe4t3K2Os7YlY9tebj2upl20jIzf9iqh57+QbvrFgUI5HHd9AnZbxxKz4CWV28jQYw
vBPieP+dYeCwjBp9elAhsGl+v4eyTOx5wXWJwJgq7bcWIau79nTyreM34qY/2SXKzhkn7a5dq++1
Vssq3Fko72WB/HrB6ReI8A9gJoW84dzIlvdF6EUtIRPpNXbi0xzSyMlAqUrkNEdIQkgMYEx+ctO3
G0LK4jeaDlnTPVxfgKkKTnlHBYkb7ezaEB1lNGjl7RvPGCEmVe5cMyFH3QgSffmbF9+br0qFxpgF
a86RAEPGsRz+kRnQvTV1qttGw0eso0BxuK8F7DJ++21qeNKHzAL9evDjDFi2GLlg6qL38uHlO6iK
mGkmJKK8/xQAlUqK7pqJ5A031rCHktQujL4n1R5gYXRtom4ZB4XHCnl0k2bJGngQkNO8tt8Ow8f3
ECioyH00k3JxOFpASK21g2ds09gX75Iq1HF8sXidASwYWEo5Xfm4Pma7OViaW1ukB5MXH0K1suKu
zjpzkmOAOQwcDLNGt4h95BFGxj56shAmMb3cI6DUr1X3DI9pR0I9nPwXJxy5srdGiKX55Cg0yVYQ
xMssxcbqBCsjn38iI2f/O8gqMKNfOkDkYVJ/ZSV0WKl6ocvyx848ZPrUaTCygWHC82obF0jfgudG
fQsu4L2fsasZRu0qy5BjiYxS+NRFE2/1Svp2Ep7TLWncIvr7NyPyDXtdFhUEiMYdu7arYJnlnelX
HoKGfCL9V1CIzX9oLc85+Lsvoa61KVLJBysPNqX2+RO2iHackc+pBug/v0qnDWQ40YRqTvriv2hy
7G53o9acRB8kgPMz6V0xVvYg1Ej9t8Dw5PhAnEZqlnbSNg4wL199mV961FAXpnoC6mbXFL3uEkU6
87fMxORZ9yPeE+fGokcyvZECBOmXKv67fP2gGbnGFiemlFONYtpB06XnoGlFBBpajxOEHNgT7lXb
C4fDMvzyAmEpMsfGHx/Y1BTrV2Hc+pHTExPyDa1JftlKtM22aXuI8Fap5uvapE1jtU0vBCrfMWHt
wTnwjyxmg8f9k8TrI1sIAqz/1CFWNOi3adeynRNBtFC0i9qjv4y1TMYDidGo6l2hoFslq+16LrIx
WGDJGsGItYUe+uN863yOS1mcPDCD3d5/PkAGbBflnb2LUuEgayGv0cY2wLqEJMjhp5m0uwUPPlAM
5X1CAbUVgTAVAew4Nmdtuv0FAkfTHuZ2OTTSTDSIMLBzvEL+AYhD61Pi+g8herPSQM6nKr8psFkI
9DT4+mYQV6bssA85VtrNWt0nehLRz3mhnMZVff2E8bnM324uI0rLOYYPILW0p518gSnVriXw5yC5
YgE567sEZDl9QRRrrrG5BVyRupvNYqBCr2D4r8BGtgxwIXSSOOWRRvLgscJpFHFbEm2AC4XXZAT0
FFrmzFZSVYkExtbFhVnymo5vsDGDJ7Bgd6w1Dh9Wq1PGYvLA5VHDtNDkKAWJSjVtQUFoSazSBUA3
VME+lCGvO1iKKK9JdgaGgbNUc8PgmYF/6jkgIUVvxmUQkkTWipbANGr0PY8u4SBMtHtFfj4NdlHO
ns7ugeviyGEfuvt/PIHNmRXEry1g5qkhmbDnnWvldVK+CuAT+G/7nhzu/D/DPXZtjcL4qfc8060b
zBg2cj0K4RS7PVzIAYKpBgBovZHhgO4mxAG1QqbphE6F74bilurPIUGRQMAd/hyliSHde4UDBcTS
iRdbVvLKGHU94aJiEHMu55c/l0auILiZug2VGCOSG6mxNjD9lrT3Tya8loq+pBPissOTjv6va+kP
u5hZAR8IjFVQNPS3pJIbgEtg+7ru0wKu21q0aqroo1MZWPE+fEqJ29505+u4DiYkDx1LpYT16ud7
bBxsLmasp9dy/jKKxmdrmENciCTNcFEHvWUlQnsqc7z4R42xCX7rkFPefORHBU3pjYgniLF9MMW0
ygC8p3IIjhF4BQ+TIv8sr4LXQ7gwebcGfQi2iNLzSN0SR2z4X7Jlj9nDWjxH8lG24jtK3dhVCEQW
VKkKYUND07GEvImsEAOH5/tjiYox3zWcU2IFv5zRRmE8ATANkpCC5Vn1Aarfgit//NPiop6QPiCe
4ivWPDbARQwWP/V9Y1TJnMBB/gDT7hXXbkwEyk12cn8aoYJlQIg7I1Fq7LRkeWsA+Z3DhUoQdC4h
fAkEZYsbl0Aet5DXHDetrivY/620uJPq/orEC5z1oeQjqHG/BmVF9XgOzD2q8Xmn/P3I06yRIhxt
IeBrULhOyFHQ0kUmkgeAkSiKDVQH88/VICx3GWyy4Y3hHXntPNQ7IdIclZlHftxZut0NuQoK+DbF
lCwspkV8CxbhSlj1lY4f4SqV8qC39NXHGyRj6KXURX1XxcjOBshJRj454a/GiEGB/2T24RbrInWj
sDnmFLiJIjoix/JRDSjb5P56u7f1Qi0fJzI85f/e7zPD2eUb0Xv0OIjF2Cf+G2ToBX6Im0Ql3l/J
Gg/fHc4bOaysYvWfDEw67HAAUiHkoob/T+VyRF/NHySRW8qte39aHTGXLtva+syZD7yiW3PcrfZq
3vKOk4Hhd2y9F5j6U1IaLosAwtLZy7JtBureRh4jbkHeoFse+DJpVbGkSc98NmCJ104/0WybJXKG
QJ76vxfmfb6V5L5vd3b6eXOeS7PIyUxf/dW5QTiS+2vYk1orEC7b/XK3oOJkxnMTA549yAhF1G/0
DieZss86cpf1nWXydOynmjVOsRq0x83TTLYQkaUwy7AqQ8sWl9mOxxtVKLkQeiZcnsqWDWvm8FRk
FMFg9JfuRvHRyk0HwgRJPQGt96kuuAPaKN2FiEMS5yxDn92APKtxEoFjk6HRAg0W2WMfgIEUvpDu
Rppcv+D3f4DB6CCELtwckwE5BBqr9p/meEeGt0b9W1mYnlcnM4OLGL8vEbvxzluzGPmSQSySodiB
XRWeUrYgrMJ0IUnSqnDMaIT77/OaQBBNJvKBVvxviokraasNR9ph0pGOvVnWoPz6MKl/l4pNlHY5
ZlgvDXVwbFkt53xfkWnLtPM1XGsBjp3Tm6QifCKpCy5Txdfom99UtYNgX1T1TUe2SERr3XDnEryV
40oYMvoZq8IsDkMVLU2/ivrcdjyDD6Xpxh4GSSrvV418cOg5p0y/5zgBa0f8Kb+K+neVONPh7hNk
wZOTJNOf4nieKmn2gwu9BGj0bZj6WL860OyRxo/3qB4Yo2qWt3KNA5WkZiWuyWIOZ2u3Th1VT6SS
l95wJ5CEs5zQXIx3bHuHHGIFhc5VORfL5kXKhvnIKUNSkYa/Wdi9w2IEHnqtPHzBFQMXZzFUWRVY
W7QHC/5zaZ6cvvF9uqaRR/UvzZTtQFF2saSzMW4ae3pyoIgYp1CvcAmQBBDstV90velniYpDyQSP
IAA9LOjs8wkhIUX2xtqDe41z5NVfSwFIJ8xHpbipx46INv7aKogag7MX52cI5XJQ+cIfyfvtxWT1
3a1gTXLmmOW9rdI+T9OX+XHBtyzU/wYi7zz4MfrKuuXyACCSqCFrAmeJ/2GbKU9HG3Hl5OaoRP38
n4yuS3W1vvKrxZTF3Wecc6TLq9k1Z1n/7RlUxWokw7S+DsJbFT0YdqEPXB3p3uxwiWqI7BzNOEG+
KgCNj6i01ro9C5vIWwLeDhZXxWDXrSZjvCFV7WKQFfySh0eP8i483fXbyHrqnr6FyouTKwGOJagw
qrzLxseYPYMBPExwKRbB3ujVHa5D+RvriGtHTjOMSb+QNWQqMwPdCcq7iy/Bkd8BFmYLrnLLlU5y
dvf6ZGyfasWLnc4+FLMOTQfEnccGAj9uS4dxO4rgaaQdzjnHSu49JAO92yhah2h8yQ2NRDmNYKCB
qDlWZ5bklVDy69Mvfp0HKbLQLFKJkTLv96g1cRIQ/+wYvypKqbOIhq7KNVst1ztgQfKCJzsLWz7w
NwtpLpxX554WERTRQMr0BE9Mk4JmsC7Ca26Swh7YY8s89yePEnmUmjXdpPwhEDHHt4GZGBfeCp+k
c5jg7G/nFJXd8LvYBzSuAS0ZVCythG0VZY3h/eJgZmYDjHShHVNrS7XMjZ1GCnpHpRpgrpwdD/kA
yZw8wH0MbCb/J6olgRUZjZ0iogZ9VIIQ2g1Id945nIzVK9yAvVWdGLPumO/tvC+4gHp5ZFne+ekb
DdmGgkuNstAncgE9mHiYfHe7pgF8F+/MRjIpUIK5VUr1uvMFDxSpBu5rmZ4F0P+mWxOcqK3E9egU
4zD32GFOjpYe0JJ7ygkHVbQSwimTgl2LEkMAXdpu/xhwk2H+K4CYwfEg+yGgrE8MGLTwkKGSisoL
7NcVKcKZ2t7Ty72Gv+iwh0HR47Iys9YyC86tYzWmMpYgs+7N7xC7/or2yK0DNsSLhUf9KuQ7S1RT
skilcgc9Vyx6i9x3RycuyNqJbyoabM25N9GuGdSw4fJd2EuYYzAhc5fmoSw/3YW5c21sS5lMNAVu
GGJa1Iwul/bH+Y+QDVzSfbEvuzaoxqEiVxNf7M0+I+entXkl3wKSAeN5L7GER2eo8JkbksxeJK8d
KFV7/DQm9bC5cpD9aMY5zWf6i25258Muw1jWDyRuE7W7Vq3BMYPUEL0mGdQhzMewEUVO1Ic7AcDU
GwWRRllmGLf94Bn4IDAHOtHEUUuUMoPK5tuGZIiUkAM4BqLA0rl75pXvRrjAyQQRAVISnzzPoxaY
N25wcxxLcr6pdODomSxHyohpvna+pMezqN1ZcKHV7/UwJQMh9VveMtQQXhpzbEIDM318P1bXLslC
ktajpC++JN8ruXl38wvUj7XRT1vq5aY3BZJReCH5vS/HqDCSoxcWQinXLtFb6PlLExr8LMEM9HQW
41gntolfyhBdy0Etw4dJJut2UaFGqlpVDK4Uw9moK7tlSX3YSb0l4ueQYqIGyZJPKFq5wA7FPRrN
D0OhwNeIgs2XD1/U0NVip9vucFGkvpvN9a1na7AGM9/M3KhRNlu24QeSGOlC1FeXdMnRW4CxxKXR
m/IVaoEpCcT1BenohkxmYUlhfRzQCkNMuZGf24IbhoTRPJ32e1pkBC1OdVIqYpZtzgWcrcv0ZOgg
TRKEUnd2v/OuqHBm+wd/0cAAk9DEWBdjKraBt5BaSGy+Vim/zT1mW59KA0VZs8mvTleiSNv4pIl1
AErTgUIoYw06dM+cWaS9T77CsjzooQJ8zEAG97F6wDlYuYGIlknQg3t5lTZugzIrzTx2znnhdgd4
LvzmNAfBmCaoUPKIdHy+PaxqQux3lQlPuzjp+VEJ4OevD2tl3LuT0WapNiXU17Xw5gRGMoyOn7pA
NgRMX52mSceM2OenMLAFLi3/upgKhYz9AX3f+E0GOdZ7KoEHZPm9dL3CE7BU5flDx4U8W5YyvUpy
mN8P8pMsZnVwtGejEV+6cK9tierE1D9Qthc54VvahqonYVal3Ctbv1Acc4yNk6uZtzJC+sgpM+qt
sEtJqaDW+S8vnD/2FSS679lrujw0VTRXkpp83zLmL2K3TR2UyFatfZh2EmzKgCchXH2ctu0EEwpg
zDmfzdh7jLKKIeLfwN8BuzT5iGF9z8SCuTCPxHf9bQdyuaYHqxtmbT6j23VYCf8otW7RDDsKcIKp
UUcH+OAImSzuFDKJVMCW3gKWhv8+eDl8PVn1JctplCv7TuuRrbuuUsAnh0k50j1vhv3A0cNRV4w9
FgtIH1Gzf4cp+tBmEIb1PFf2ptma3Nm7yJ3qMNa+jOOsflKxJHYz/DASkpyyGnaDeedDT/yaISIj
eTTMm+dF1EY3iBjbuokcjOIxzNt+IA7T5VB/hzOS7nW+oZuRvzWTl31fknpno+DjCLbfRta2THMq
7io0JzUR+dl8HbSVgNOSjZclAISIhxWQqQp5VmJejKPW5Efn8ehDF+VfTRvWjZ1l9nDWnPlIjNDt
pDT0FFExC0t6Bet5h1udp4QSN15wGG7RIIDnD0UT/4gZvSdQbN5BajFyZ/aZiMH2Z19i3oNNW5Dq
iEa4Ebc8umIiGn1rMpEanNF6kmunSkoX2F0lXaSzyoYm14QURPn42PgFcoTVcZGX+ONXwO0pWwbx
8w7pTOui0LccKlQohLjUWeovzUYZkTpJruZRXe/G5r6eO7ZE2jyOwhEcHhgIAUPsP8+LEx5+ThmH
PBO9BBMBtLTexUVfnNsiH2GfwXcNTwt2o3onIICoadPYHSPVdyihPA5S/YfCO+zRHtCbX7GqVfFL
H+i7yM5/yViqEjP3cn8RKTr0qFYLFHeCDr18WOldVAmg2qNQtNlBnLja+TtS1zTuPX0wSnv0tWL3
zmZGi+fnj6Ovb0ERVWQuIzTXkl2UcIE0CtiZKF5LBHlf4UeaZARfw8FcD06Gsr/raCxi/VPc7euf
ZdFnppZkMRy0Ji+13BiSAkdjv7OjhRAlYjA48/i8Li58A87Nnpqa/UCzPclNc686LW+a2DMUjcRn
G+GObimIen1HYl5OxGZ8gSIjqwuzif8uRsDiDhGSm6LbgEOtqBGZqczXK+/Aqd/7tUShHdUYd4yc
3ForUDPZM0QLVcbzZHqStUlZ5ViGyMA/HgNvbnlSGCZcGhxFiPMzpKg7ExtUoaxHRsQ7+hhT9+r0
Wlm465RpQBXvdG1qlgvtAojE3xndFGw9GDmisP3rjVk0+0NoG8bfC9lmohn9zR0C1Qz43AP3eBOl
fL1onFell7z4gUmzUTOt+gQ2u6k9qSPbC25ztoIoQyvpcrwVDs1qBT5tSeyD5ja1UVwDSYrLUmcN
Bb/CTBd1dqDusK2O1YnVN6+cyfHNO0WYkRJS3ihkKHTJeohqlXpi5CmAHWXxyqUVVnnrHKynUPUH
+n4xFGz/CQ45Gq66nBVEe4MtU3QT++46/aJ5Ayr+xiL8rhui1H6dnWXrXK08QGkQCz13gZy5l6Yp
efuYVLUU/NczZ1NrWpJTvaCTmV1+gGzpkDF03/Dzec8Cwfbs0C4p7dSxlHJx/ujHRSmUYfdavQX+
zJOE9J8TxYevpEfQaGAmGvbJ/Hy1qE1GGPvnGCRV5Rz0HXkMjt1DLG/EPCySktHvIWO+FRJjf0q5
ZKl3b6swRZKrWJYyhezYnwcgpVSMpT0lhR6gT6bmhJ0mE8AM5iqXGBZvCeJhR/IjWLwbzvs0rou7
BTir7c0o+pPJi/5N5ODuphFPoDDOG5MLFsgZjLxzskhih8z/C9P7LV/HsSHqQFUABat15//tgUzu
QfUAy7owuWzLwG4wG7JeTAfgPwCXuJKpuPwBSpQg4Goh/Hwq/0KCwP3EGYgvd9NCjOUVU+DUHzju
v4eKpYV1Y0zkF48Gd6onauNhxn8usSUV0MkDJFw2YvGGCu2MV1Ngl2vwSC8/4ERQC3bTf20SvOV0
bYlQXeh/yoAjSObvqNjwZ3DG7ZkBzQZcdL0YV3L1B4bbDrIf3hhAOjZOdggPO+lqn/46+VWIAv2v
8MTN9g5ocERD/smRjA8/UF3ixLhCFw+wC7qoxyp+nBBK13Sa343pXwuqy58xdXW0oCXnOF0JhQFj
I/BXtGwsVpSn0dM7RqtfctYE07C7VAxzH1m5GcCT5N1fuM+NTa30L00OWgtm+y8yPLQ7jTn8aMo2
CNnXZf6I+fS8WAIIX4R5vx5bWdpXjD+qgLMp9+UXxEwj/k4RUetGHRp7n9tloZMuqUgjtV2XowPB
Txnd4OTN0nLtlOlkCA9F0nyu3r2ryBsua4n0e4zDAK5zUhzCSUd2CqjftJITb0TZgol1Gn7fWZc3
gNa1Jx6hew4FI0u9KPTbB9gudqvK3KL+6YqTuWyj6cLhsZcVGHHFT4YtPywHtz5MceAdVCh1QTrU
3aOvNUChQVbVHZAzfOgrNpwFcCOO1GMl2FneUv3Py67NUMxNpNNrfXrG3AEdRcm0YLWt/2V5w3Su
MqwFpM2N984NeKZezC9z48s787/D8oA50u8dF77Wo1NMFeTc7urwFlQMaHXP953jVKu7Sqkcp2FA
m1uFBJrG3OPJehjWon5bKb4ai/iL0nhOwXFDUH3tMWJWbe7ZfiqwD+5Y9yfwy/8L9fX9ODxrFmDp
gWDRRhLJX/+ffXQD6n4eA8P5Yxl2/jyPm3I4ISHFXnaOrog9MWndgoomr+4vy4IB4480JiioIZgc
e6ZBw2L3GUPQ/A2wHm4+kyxB2ZlUJy8i1zMLtA9fPAzxgSh2X32Fc4NntbjfAMgKvKGWtj+vGvFQ
CkQ1NVpoDZ2UuZF4dflVyFpgKwzHfKdsoeFz8ElfjK3ntnwQ/siwyqrWPfjRP7Bfg2XctRVIz5cu
I+/Cty+YyQdLCARur+bF3r3Mh3SDlryYPdaeYt5Pmo1qvbqbz+jt5MmWSx2thckS5kjQHmYt4XAI
+YjWf2lG+Myh/ka0xpMuwuxPmeFQhRcgzixryFI8yCLIsW+7pjP64Brwb+EP3oEEkmFcxo3yGy7W
sKlSxYEjTDq6lhYagjO2deBle3dAclvX6x8cJFU8XAHleSo/kwNpkecs/1BVjwcAgL2B1Ah6S4Xw
Gdivw9eiiz01H/XT6Rz6/ttqHIi4IixgryVi6keCwOCzzQkN9RBOLRPdtkIHLYnBPcH6NEnWXYW6
1uzUoaO2KRA+IlWsVMwn6rA4znWh+u6Ftx1pQQ9kAb5kNpvV0FSYUSEoSmcKcK2+eEXATpLwSUJ/
dCOzosn+0BlqNoLTKyq+w2BF2JOxJdzBPb6T5nGQ3Nic4uNEq9e4F0qcNBHNi7jUlMNPs3SFqvKL
4wNVKKn2mXGFaV84OmFwKrpa6MJE6P/kopDNYShiRuBodBXjU2lIYrWnCOdF7Vg1J4i/xnucW+mL
Z2SlPcDXIKEuOorcngugrayucenDl4ircNdOYE957AHrZ/atigrvViU7oNbRBkxnHIfwxni1AQPz
9TblW3Rkkv6Za0WS+JiBpYjqQI2fg1PHkFue97I/FSy2+3oJAR1cKYoEmHaeL6WI/yqcruUrmnYN
WNpzUV52ppmneZAxoq6KIsnR0F/eAEAjQGr+mhabAL5lMnIs6bIWx+H9dtxH2kQR/rawfBZsz8qv
/bVx55GGevQwsumNp1uI3MIAVZH3gfczchhxM1XeLUG7BjCwPUkPrLj6zF7sFN4AQ78dBZmqf6ax
pQwLGIaQw8LbxAWg09SNFbhYSSQtuTKwwYgrIAFwVVel1pLGx0haiKLQrTsSoU0k0jOf2oXYBon8
cowrB4KhsNWYkGB5Kqb0sni9EDFUMvRoSjAYB47NLPDTos1UrXrh1sON70QJ5nUJ2oQxyc7D64oH
vBMW2cw5utiRqtLS23lwcIUIUCAAh8PYf9UB7ApwK0MXCnhgC3sQ41bGXyg1mMsUv/23AfBTTl1O
EYjxD3Ck+IVGHE3T6wDRCixYIF0JLGw8dbZv5m9Ez/JULUn2wOysxfTG8SNgq6m5rWWWpzm0bmQP
3LJED5F5znL4gLngV/iwRJmBj/j/WaaYidhNWdffay0tbDaHvSq0FMMxKf4yhl7Ux38hhTV+QPlw
T8Ec4vqqcMRPv1wPnFrLKymud0cldJdXoQlAo7u++DUK+guTK2Cp40AfC5+aJnJtqqOumvBfJm07
NJ7zz3TAksCoh4kuRWSmXfXSslWKyw06iT2cW7PhK/FMAoti0j2DV46emZrL+flxjAv5bQU7/mNA
sz5HuK9oC2GzaVRzA7cgVDmXBvcMTwoQS1kfPN9u2mGJqyn+1rnTQ+zUhCFm9KuPeeZCOt58Aw/r
QcmI5BjBHoH3DAMmL9JHYtA7G7sOJ5khTQp5/31qGnyGEUaLIbZgCU/o7olVHWlECd5/Mp/hTR1A
sM1QqUJBb739K7h0rsK0dmQKT6NIHB/MXXldYncSRhptoejyTzVDrgGXsh1Hl875JlD2aGwII4yz
GFArJ+U6modCq8Kh8SCMa0X+VmJ2oFHx7k7N6DwJVjgU8FGXDBF/pz28rowjYGQr2wDYhZUSub7j
AWffQYJGzWv9KK1Hs4vg75ij4n1rQIsyXvJJpmaLE3WFSWeB5UlVFxKgX2xEzOdCtRk3ssKufWCL
MPNlmXcZny5UrXAzkGG3skFD2NE8zoH5wNbdzGINF+53xiYenqFpZtrWGUqDLZLUO1PfzM6Y/v8V
WldxqB7wTGvHY4Aw3SDbEnwIpbg+ps26c+7S+m55KAhcUqaEKlmj4AVSdvEBJXm05Mtix0HUboGZ
7coqvnEBsdOAS7hbvQyh2//cfuKAV+MlOvlswEv1Z69zm2AbvixMy8AT8yYAno3YVt8VrDoeWQTt
hB20WzZR97D8brVZ8pC83tT/Arnx9qjX9UBJEOUeXuzmwqn+awzqz3Kwtgw5Wgwf5TXVpmEe0RCC
rscEtAOJ99Zlj4A2mqhgYNVY1vZkQU7DfL2NEfToQfG5xihR9HmQDpCXav2lEFvyQZAKIoLtSc4w
dJ3N+U3lyHBA2l0VqoceMqodqCBPNqUxfG3Fh8fbEfuNHT8dBdEBzTPnfoQitGZDRNVXCPdVLLsC
oB9kmTgdP9/BezX6uUmeaydG4Rvs4UYXjelaaCQC14DpmqxvhhLilFdkeU4AB8OzNhwSl3gumy+R
EdlC8QLmn3UTbHRyp/NGrVDgSCZVvXxIhPbD3A2Ju6ybizbMxBHrI4Kf6qS1XDi53elHojYWKIaz
zkIwagvFV08Vj11HCS96KMyjby3M9+Tz2HvKytONbd3rAD+TYy10+ETndnRpAfMlXoO5JCawhMEg
iX3m+BVuoJfynst/BiBw5nfNrdtXm78YmXbbAHr683VdMVbqK3uVqBd/m4JLzML6taV6eKy60q0l
McFExW0Bm74q2bTm3vQg1OGk501e4Sz01fRdnSHMHOacHeADWq630AWMVUXwYHv2zaocqlg5+ZZ8
y6zgBPGrGgZM7C3SZubP4PEDvvZ8APm3B55CdIqo6uvylHOQIcoZo60xvkts+xOqNe+W9uo+WTG8
wifG594TO8XfjXs9vCPKhSFcy7U61VdNA5eN++h/1fY7vaUN6HaeZYvgUzVB6+0cvle5hBlYwpQa
bFDYhtgm84Ek4zpkUL78niKUT8P3Zbfdcu0Xtbbk9u6bW1PZFIuWyDn2rEcu1uaLVGsVgqU0IAHT
kaiCwvsJvLm1x2RExlE8E2VWxt0e8aVme+EFoL7TfNKcNyI+g9Ly6/A2i0akhr6HH1aGo0UhwiX2
O1JbTgcphSQm7dST1TNoPTa+Ch2GcKvvX8nieDlUodzTnG8Zj84MQxQI8/eP3rzeUKLq1MVKt3oN
mS3MmyaXr9cU4O2AoCjehT1/oItvGuRUqE4vgf7DcHntNAaetWy36Eo1Nwi4EzJUFecmno5225Qe
YcCIs+3PlKL0dwcctJ8MWBRciHK88YUIsmEjmj2WU8hK2t/EW9VPTROo7umA3kEG4NLPg8/l7O9E
sXB/6KC6zDgNDxEHe+ITzLlsL/1aFBXKSE26gojOosxWgHVwQot7e1Nv5IowlTwpI9TWPb4Y4itI
n3k40f3keP9VDx+8GQ+0IGprGbo6QY4s3jxrifs3BrffldVH+GHC3f7JU52tCvftQIKg78Ec8H0C
1gm1XGwD/bMzsgghC3Zu2gvbSVts4ss1bYVh2ZLq7Y3zdJOyWMj3yneh4g+Q1IUioCsU20rY1nX4
ASB1Zp/EIZYr6XnjQC/7T8T9rk2IX+W0hzFrlZJakbs0DGKtJdIbqKyO5ghh0lXzScQlWN453z2S
pDK7SXErXqGYqdZDtNMQH2PvWm9w07U7Pwjiq92irjbfRPjidKwAlfbSSEWqVMGnyKaecmiPIDA2
OtklhLD8BnoBmUw5dJ7aJNNCFJxSBI3AkGeRBlIMKCFEO07jQWq/tZ5SMi9EHj/0NXTQxxdZXPEd
K8J/zovPodIaGLogr5YlxOTDNf1p66wunlNrVDOzN+qfurGcjTGfazISvI4RKEK7a+egAMMX6d28
ZTai66/4zfFSkHf2c9QNJojnjy1+45PQmm80ESxjYVjScJDYASwxcrBp4yOvtb7GGHdynG7zbjQ8
38/cxMN4yOy27tBq9zkogNW4fzZEkgV8I4BN7mRzLk4Sv/BA7BgI1Y0+6ZeGbkulypt5h8p5KBLy
ivU6nmRp3FfkC5skC6nA7Viaf1236cE8Lsa7Qk1xjyj+WeQoY+1VdPg1zK0llXK7ZvV2XPnEvBGQ
hq/RPmLBX3Wcj+LI9WUaBanmuSXoaEj8WBacBbXQpdD3MvlSZgBzfAaqRk6MFGCO8xHAaCxhv6kM
CKKgl5WyHiIHZTYhMKxeADcBgkAdmfzfPbE34d9jURCqC2rZZDRwoedK0oXCt5DdXOwV9knbqcmo
F1OXHs9SmPA34BJb2Zix1yts9ZzkNtV95Nn2DuSJ3/yppCiiTtU0uYVpBaAFXE+bbI8tL0NCSB+z
c8iU7umiK8yLI3IYRCVmvXOqVBTMAh+NVXzLh/aioiNXSW3kh6+T8idIrVI1JX3TVv1LMqV2l2xh
orw5EXRoXiULjVzaOyZbt2/buAbp2/I0T02dZrNMVC14C/PjFQS4b2g5AgM41HFUFuMpXH+KK4LB
kbZgzXrpLFjOgEJqLXKee/8TSjxudFD7HEtjqrfUPb3jmKfxkLv2ZI2mBjQSm1YeSVq+38lSxJnD
oMhMLZT/AfMFEPnu3T5Pf0pjL4uFQKe8vI3cZ9RtR2/cnERlgW2JpBhd/SGBzEqCVKMWpSu4sLYc
RiudcXywpS21NB8HBwACmKb72+D0/jPJid2IeEMCAQLA0U9H3KQ6Km/aZ7rNx9FgeSSFbJGYpo1M
XTzyoVChaLN04vPpaTF1cqF0anq2G66KYa//RwjT+F19jYhDq1wV4GEAZ46UhN1ubImNQMQD5h1s
Nm8FZKwXXHhd1hGLt0mEm/cbOe9tDRM52yDMaOACEzaxFebWLMaBbIJ0dC8kMjZ3cJ2YnETVteLD
NCkh6jSlXBIC7RG7NrPbf1XUDRXphLv1xd4dorwgn9Ay0HcrMS2yQoEJVZDCxQ4Pkd6ENHcy2gi+
03vBPn74j2oWBdkFwIIb3uMcTN7lXl2uCuX+t6P/mQ0d1gE87QbxJACzFYni7Tn728llS2TagjnI
iKfQgyayDAG3Zn9vAUbTGEQhRRn6f3lvCQjZ3Rd255nMorxWwfqPnXWrtgbS2QDdjxb7pPDztQl/
iM/eOiytNzEbb24ybXRB3PnlyC5cFcvjUZ2arwi0/fPPPTVJZcR1M5uezImS+h53hjmx7bkBiCvM
XO6sPHV6ZDhPbJ85DI21a2bwNjLBb6H2m9rnD3nmAGWcPF+9ex8BVfVLL+cy3Y1ROH5ZAV2HmxNf
JOCknMaXUfVF6X2TNuU8kRmmb32xTonN1er6WcZwHOlJphGUqB18N5cDufD7DMpf0bjqJdgsvuaJ
pkRwp30ZF54KJKGt4cfF2YfXlN65OMRF06fCz/+90DyJQYHEDPAihyQFK9zJGVQU5hndpvTqVOG3
Czq4NL69OfFYCBnEXdOAzfPRdZ/qrAwLFROAPzovbHupQa9Bea3YljuKxoBm4m0eSuVW5X6B9TkI
sZroMBf4LFHkZqcC+udYsBjcerApS9DUfP41CdR0Ar4xSjVoJQugxc1fdPqJezkzUE6nad6UGaMt
U2/+X4lMpm2pR8bxfJUGLx52GE177ryhVt+kz1XoQ0my2b3P1YXk1H8hZRpSbqLh0QunN5GoQOh3
3b/bkEkKtjpgU6jTrpnpS8mV4DBPpGaJnhZwLdu6Gi7vHG9DwlxylR8Thn58kNQT/hkUtTl3/SWw
j7UyRzdjkfRp1o8xYn+cH1wrq+s7QRFjmwdznJzgViBnyCRIdwD60LzWlu2ndp8+EprUfgTIH4p1
fMobeBhE7d11hE8HcFVf1iMVOEFIiG4nQnmk9ok/XB967dnPAVXmKvTcUGaZTCFSNFQ/7AMaYvnH
R/KHU+A/NOCK4w93kF5vRgUrqnFvi1uJFjFJqzUkoapF3VdCDOXUV0ZbD41nFzAU8n8KacwqIxSs
gCEYEzS7sWFPUAwT92nLs/8Tm/CyejugQla2j7yWqTAnp202l/0Zz1q28T9iqPdn9zmOANp2DtQF
s7PP9ICFFQqX1rYcWDA0DJkLuJh2S8twPmaoiSAvp84sItwYDZ7d2KT1mU47RROTEa8MUR5hC8IW
yOj9HvbWqD0iPhUIOoSMa+Ah1q70hcS2R+If8dA+7JE1Y57BCnkxAzC06WsyBh9I9kEZXuBySNGE
qWlBdSF296qX7Ke5QVlM9AFtM8l3B6ldXuINwfCiEegry0Pcx0+yr9EgrJmONj4/jtNOnBXT5WjG
ECgq7xy/xlbDyOtam6NHZSiCnevjADzt96lmlSVDS0nm2grSMsBuceSP2R0Q0bWALbv6OBHbE3vA
J/bOVuQFSc6kndGxhZGZysSmi1daXdzOA/Pgce5MEcKQYMnfA2D2FfXdYYlSFdf6YsPL5azKvkMi
g3JWsyXTzG2XXNsldeGk6d6r8ADy+ZNTVYDtMi5blJ5JwNITp1xmsCqX+CZ5U9cLhe8xUHzbS2ok
efCh267bUKaNuYu4kNiEHSq9eZVyhylhLCUeZp9MFjQSJa+vQpX2MKlYywFTFokjNu1xnpGFkB2k
9Yo2ocnSDNosMAmJ5/m2uzG3Y8eCFVIGQf2iKaoiQZbPAys96JQPwDswrJx1dGpuMJBY5fJWfcux
ngDJbAkMY1bUg0f25QszoVC8lEjhXNIHeguF+mCemRRjZMz7X5+K6khww6ck4Al2pBquuj3ANg7L
pQV1GN+KnDMNpossNJ8UdymY3J9SosVLao+zv8MKhxryxkmAa8/jFDqlI2r4XJ7NH8pg7eE7eI+T
AFwwcR/Ov+g6a4QVs7GRdOhae6GZ17Gj9ULEkYksUCUn3JfBYZaSFuAWDsybkZHdcKnuX58SYDgU
lHwPiheOpJZqPLuJZOeJaj3jJDarFTZGb6kFQnEL0hEE7DScJjtlEt/M7J/khg2/76i4SHtFcVxt
mE+u7+h+FnLskjmiYwB4PvoSRyX3qzWMqn4gYOiFLw27Nzld7k9+Q4/ux5eb3GjgiziOKaOXQmp+
MVw0JKevWoZgzxeyTGSgeOS8AQ3wuXSwkPHbPNUbxZ2pboTbhH2tpipmlQEzVJTO51etjDqiHUTO
RgqgzI191rHsBflHZjqC49uOYuyHkAgEFnRKo2yKLIOT7gKXmb/LQDaBMQbPkby04OylHtNOiEze
kkv1nyTLjI9U1Efp8f3Mo552Y2svoSL+/RpofA7/ISVhmqJRVKuBL62qrTwHHioWd6fyNoMsh6bR
2Twzt/ESW1anmFhjI/1wBE1mkykE9twqhIch5XLSTCqP4YgkbaYczOkED9CF8ItlqNlnX8cVNPMv
xTcdJx8u6kcvVY9UxSzsg/Ga041Xwpzpe9uIbrALF1HuEhL0bFKfS94ieuA9Nm804H87H6OPuubQ
Rf8WzqTErfHZX4HeRa4pJ6CCA5nkuhkNQtIzmoxLBJo0D14Bou06isHRKSLZNbByvlSLS0SCQLuu
hpeW0PzbeYF/amUxRPTZdO9TOLKe4NFsRAGPS+6I9a2LZ0hprM7qANIPdhFzk3YbCnn9TXQHFUME
w4jzX/EmmqOuLhO0zKMosBZkq8jm3tIsvJOuA25fL2PhMLsE/Mp5FX+WpGKiA8eEQkISRwXhYl61
mV9L0mFhaELK5kqcFj4V//xRXccaLvDBOxjEF4kJNF5AJbQtEkbbx5pOKdJek80ydt9SWkaYBuM1
px0IX4TkDplfH2bVG7vdTov8ef5E3rWCzeTM+TciYG6uCX+/+gxLXgQ6WdYEh+mJqszMzsIa5fjf
ev3jjFGlDpDUqRYQ+EKMtraRMSk59HeQhNIe0hTu7Ihi/g4y8uJTjvgzkGQ1dilfqDW83CgST+2C
qYGCOEYYSL1K2WpW0KH2IKNXdXUHnKeML3NxfNGkhulDGk898o9OM3z9EMevWhC+gDzR80UWe3S2
KuwtVMD5IaE2pk2H+Gm9G+9NJE3viHjSlDmpQzrFeKYo51fsZLQ327Av4fRs/kQvdKsuroLLYPV9
ul/8BqgPYPJ3hZ4/IAbu9tuV+PqzdbeGdcDZelqldQ7cZzNccXPv8zPpLaklECnxYZfOC7ZqAKoN
1J9/trnlwN9Yoz8xEldpbRGz8JOtTMJFYw4xkfsjhws11zrVSQJaujuuhFFAOGaON+QxOXc7XojL
f/7HYeNjHukH/KpBv6UVgs9QjT0w1unBd+qViukAn1OOMes3ZVmYNBWGI27o1siKFpg9M9kwoEy1
63wNhnMY/+QGD1WZv2kVbAG3lOLltxbFFYuBH7EvbijNaVQ4tPCtRhEmhRqz7yPHcr3m57uXxn8y
NDiR+b7EbWMfT9xuUu8ziP1rw/NOY/pKtBGClxgRowHEs1ucdbEbzy0uCtkTSGS1kj/jh9MwHvtJ
Fa7e9r7LwKQINF5p6hzo3rtf23Tb5LcZI1xDenz5IT9XgJz7AJQu4iRFszS7AFwC04ZEjGZn3/kJ
MbvlsTZGT19ubGijzBg2MvjcHFMEVlG/nd7kebpYy9bTV80ONNzmg7puXZoVbO9gspKZhoxEBlsy
qvZ122mWn3sdYeG5wDG7d8sHpBABJezHsA1Hz2l4A7pSWlsSzcUwjfcmA2uCgZ5y4MAhz/HhvENH
/W2nQtwiNBre0Ewgj0aNfi00s7NNfUz2xsyEC7FMPPsDZyoSpuQDME8e/r5hrMrvlzrxX98+9wln
vFiVe7NtYfhnOD7yfXMvVM4ykKg9qIOdZ1XyuHDDWJxU+NrZefwj/TigQ6JDi0se4XGtvqg6MykW
FkCbMcPvkbKZCeSnbS2Ksk6KvRkofll8MVeedGTQSht9DAdWT+IUwgMLjNCDdR7TC/8wIE4fytsw
RRmtlkFXGhp7+cmF8dsOFkv+I1OxPvI3WuZl/VgkinU/c0pl5rozIxXz0m17HOZZmIdpA+SIDX3D
J2TpDeXl5C4z3ZdncEMa2jqlh9pm0ypdqqos+DhqJiHUUQB16woYtxWQaeuI14g1ZUAISZ0/dTYY
q9fz31MZThUvTrgrB6PcHguqi1iRDGWYcdNmqTbAhtI+FbBUzvy3RhTVTpk/M3YCVwCOGyC68oGg
25vFtiLfky2fp7l5ih3/fygfc+9oYtFP1jLwlBGw53pPVIXW/1SCW/OfLdSpkur6iLYBWRMX2X+5
A9ji/E9Ga4XO6mUqxHr0HArSrQ0G3uIRhp8tPZ/TaPqzonaOty5rBSYPP9MbIEoAiVi10ghy0iWG
aeQ7BjIeULlz+fxjjtXTQKfA71wqapVK5QWXfQ0Maktc2Yh9W1kVmsUoRUsWs1ND76xOgcbGf/Jt
cBiesYaxT5IIfXQQSlsAfOMNvjAQ4aGMrr1y/zU1vho56pgJkgZqsqBPKO3c9qdNaltQkX5/xsHb
zH7BVsW87IChZyxaLLH9ifqyppB7iVlPJI9OWUOItNTEm36Mj6s2wtKtqum5dUOyWCPOui0xm1Gs
SG2px+saDXdLLfUvysaHkFHoDH9aa6y4lXe6+kObeUNjgjW5/YSADOj91CLHnjw7mh9oEeAZU98d
udE82KALCAVaOK8W5hGxSisIbE+zTTG6IBY9TShGJ0isVL3Ixh7sB9k58odHknTmUdFaJTQIkR1U
VIK9tuCX1dQMAAx+K9M0hhOXtZWNJuAT3cW9xFtSlkAEi6EhcUNAlKzMsbsiVq6aF+bzy1mmKqc/
gqnvPpb4XZ0U72bdNzIdc7YRH3u4PyVHA0KeD5Xbir/bDnDEQv3diDKIs474Ye+JdShiUS1j7s36
PfwNDml6sdGsi42huR4l7kF52TJXHdH3qokYZFzuu8omlLEoHnAKC0Gu0L5RGU/sR2EhnxFv8omw
dLG1AVBvvli8kMUS9yBYbxjoXVMsuEq4Tk4pqmaG/A/q0uwWAH8qHTbwhy4pizMJVCuBO6b4FUtS
tFFY864AZNBnE0Kg26ir3vq39fNC7Np4mcyvJiCei/L79jeF5Q/pd5eA+IoEATxfQkmTR/OoMp0D
0yVM4TOkuzctbE2fPEX0NPfXaZNSGtJixuJtDrQ8EB89CbGIEX6GsS/Px6UW5gVtYShqt5RrshxF
7M0p+7rxkiO2Yr8Jto711UNn2Dh4L5Me/6z0JAu0s5IFXYhzXu3TiENArAYIS+GxyPY10xNXdFGG
+or2akT7UHDWE3FwHUnWxpLcyVKME0X8agG9jnEhmJyLrbrYGpe8wqWkCw2OzkhS52yssimZ8Lnz
G7HsV4xCzibnFnpQ9PaeKBJd8E+etzFELOQwi4tCLvFBdZ+lNQ7P/OfF8ckFX7dqpImZGxnmhw17
CMV35tIhSEy1HwyBTZwpYqUIBQ2xUj8JSP2E+k+xq11w2SMDPtwFc+ihzb5kRdZL+ltW6yU/OzVH
TOCxR+gPsO4ABWC3GK5DitMLj+M7Ks6dSiGES2fHLZ4iL/sHx+aqoiaPguIO4GnBcnUG86wcbosN
2zGPPyQxEyCEFbY3N7HvRSjK19dyB1BfyNe8gPS3ENo1LNKf6HBNSWe5wLr6GOGEuBQZkOcWV32y
5lfufF8vVwFuo9j0HXXZAyuu4Qsg/MRhNFJzy52hvdq6BgEsG+SUR6IbwPbaEwjyUk/8ySK5FANM
5JcOQk0lwwnXi7JtpQXea2GNNgHjv6ZScku41A8gPFYRkgRHTFiV5dJ3WpOjEgd8zOl2B88NXqQR
5pt3Beo/FPRy4klNj3fPhQolxMKbxhvqu4ruG9VC9Na9ZTHrGpvH++wPEGDMwsuDBzWtdEcQy6lL
bGY7h9xTIOSZSGy3kweyafYeZK057px1AN2eoLI3f0e8i7Zwg+gvAImTMTy1nXoziQ8qJgIJpmw8
pIbVixaAEXrIRqAttKhcGd94FGHUpEc/VoLiSUFWyrMIF6JeGYabXILnsA1Xm4++7EPP/auJo03p
jtcL5UKaxLYIIgjujrwcQiFqkVdkt+6qpLWxNRfHegRuD9V8fQ9EYknIt+KpeNg5a6uEVA35u6hC
Es1JWBxJQgXRxGuzWCq6WYe5rzSX1G8vsSW2XY67h6HNUxvfcrMPNIin5PrCsq5IkJz9ODvSmacR
VmoKM2ngv5ZRJMzQRWPYaM6KZL+7GkMJCQKNQHSm+D0fiF75MQ9c/addlLU8+0Ipj0kAGvAiRfmS
nmxH+RMu9DQ/09I9hnkGyR7LiGmNdDskC5AYBnMfDZhUuzqVXOIb89+rxH4vz4bpeP3vI0qCgTFF
REN1cU3KOm8dDkfzCzguW/2C+yZrUNNByOOwyunqXi7dOQrGePZT1nv/+hO+I0CWOVODBKdhDrOc
T7EybKiIsYGByu/Br6rPxIs6kllQOMDmgaIkAI36oruH4yzH2fCoh00eL7ExoVyIAd5n/qwDljZI
B65XzLKZ1HXaV4zJv3z/k52sQxBz5jDoE90F9KgOjIR6iZfD/NHj1tH0tOwvbDmXiOHLQzAb6PzY
ot/eJTR6VlvZXBKdBE+zR70BQiFwwMbTPCDr7gt308gVEagODambjwGvwvtW2ID5yGkxR3Hl9iBY
C64lB98+r6bfItTa0dKHcSZUbwgDC7hZ5R0buc6+K2fKQa47VMVLM7CuqW60Q98/UPel8JmCpk1K
9d8VwwowCt/ck7wvr4qKP+BcUkTjDrl+pDCblnkbAGyBrBrgoZ5QAWj9yNd5PW+rnFBrFfcP54Ke
/WfWj7fTnzOQXOfbnuIsKQ/yn3ym5c1zAYCq/Wx8oc6Upbk3EiR+ccShHSFFVe6LYE3gmwpOlN/j
qpQG0gcUh3QBNpzC9Qp+5ilWJYnLTHOyI/QjxKbbSvnE05um3wsz5TLtf4EXUTTzgVe3PXOMj0v1
ssHFOhU2GVG2nhO1jZUxWl3K/33FB41S5V9zpbl05Yij+UITqIGGcTrvfqzWzzvbiEN4JUNyRvp2
S1RfiATQnqe9HnrPtFCidzFYZ7xQ/9Y1ybzk7LNuw0pTtHT8s3uI5Fv8rPJIMerSzK3HkitNf9Cm
bTU9S9n6NfBf6FhfyHibIZ77UNZh5hhdPJnAxytoSVY8ODe/ryD6W6LjVswcrSlzLSkXIgXx9ZLm
22woGq5RZBX0DZL8hqz2/F87a0msgAqQ2Mt7C0R9kkUh31KNPEP0p0eilhywht+knMG5fuVyCBBP
CNPs4PLbrE5b89xFPGRpjsOSN2nNKUKK/wb3E3YUFqnyAYqCXTbmL9MdmA3Ay6cVI1ivcJ5hv/nJ
GR15S/XGFIFuWYDRWvcu2J6xYO+f4azilIrCu1+Ap7E4+y8jwLkCFgx2F67rTGqfKz5HkeFvWwMu
7wmbZSO5SiokgYiLfVbNRV6bfHGdHsY012bb7QZlYGUxReSdMDPXrkX8GHqW6/cQbdba4rx6NEzv
Z1lhvYp+ejbZUluPC1ny596RlEwEva2DhvKuH3FgEHqm5adVVzjHFqqCpWniUxwaDA8pUeNhoOBp
CbuXmMqOfyZvZFoOePmGsmQGNclpHRIxt8p2nDWAtB+437FaWtRnm3HX56U9PrZ1eZ7FCNHnR0jB
mLc/5cUD3DuuMvuD0v79STtJ0OyoZ4Wc3rDPoir/PP9Emh9A6tn8f8b2BejrY1WhXi8iT7V6XV4u
peNa9Gq0dFOvM24fjCSi77yPA/05D06jpkMB9ntyr14f5xuOjNz+siZvwlxaJGt7SLc63f1VBK+y
CFNAmEKPhtB+EuHp384DYyzvGDg3WNTFjKbAUUw2+GPIEU6z7h4vuQ797VOmzCtqvvz3RsolWQ0J
jtC+KHOytBFwTdSb527dewckeOqrNOsqzfVhf2mjgatEgA5+PiZQUffyWDWCgFd2hpBRHAkQYa27
0e+2C3cJgD2HohIYl8MbliLJaB3aYIUQWu5HLwS28kGdpF7/xQQ1/03zO5F+ZskLE/XEOmpenhK4
hnY7kOVAbB6HJtdd5v4SDTayf0oXmJPpOqJJxGC97mkhn1WHQGL/2V0Vl2mxByMsY8WPsSV/TDgu
WHP4k87XEm7KJeKL+q8Kjtwr43Ns/DjDIMDI1/GhF4OkpZMV63Rbo3HcNqENwQElqidSxdy2ybp+
tV0oFxy4e8px9LksOcuO03fPqkJU4Sbs51qcbQ3L/A0L5vp9el8dGH4btQd5yAsc/aG59IVoay/f
nsSrbuuNdtgpNQdRjFj5F4OS8ZClcohzWgBMVKY6IvfiXUQeuhNr8Guk45phv9tP9QnXnzlPvAum
5K3UKjuZd3TF2B1+D9HkF9CmSr5hswtCTncD739eaGh4ebktgeOx8uKszXRkSw+vZfsUsvNB4MZ7
lEGGfZCIFkQQg1ckuic+uCLWvAGQLP16ofCYl5mGs5dcAf1Pl7o82Chhz+5zH02qn45P44ufd1lA
4ctUwRIUUI104CMOHiVxQ38GKfUXUQpzIikzj/5obMpyxk+Sa7bQ8rHn6qT5WAO1BNjma4LrGLjR
41H6Bw/f12a7c2mVpwp8PM4Jf8noC4gABHCW4FpTeYMNAu/ffe5G4vpZ7X3ytxlRy5As6dr8W5u5
k5lADSpqbSUt83Q8k1X60nmsg5CU+8gp78yy/5YVEPK/v/+8lmzk/i4tvBooX3uSkX+otS+AP78x
Qj1gf43thk7gDGW+LXFhBkheSZr9n6843IOtwyPeloqNDqYOtv6UEBGukUbpgCzNE2QT0cODGgxi
yRonRvSSGDjiVa5O3HMOBRjAN7/gbk08e70w/NpwwuGlI5MUYsWrS+Sv+EizWcwIPSAMAeW8M6Wp
ZFCfinYkEDzPonZ56ipQr2aex9JifKXyMGxoY3G/oVPoTN8SxUxe3z4kcmZraSSQfoIVhXatihRH
/PaCtDGzRpoGmprOUAbyPuHEpLz63m7LrCrcDw4wIWgG9oaVoCbZEb1WsbYgyvPJGOdNdEUd/YJa
KyzTmFHozQlYB/xNdtEylWWjXTZPr7eOwaOInUFqtQG1Tu9qRr8nSVJfjq5WS9NTzWeGzvAjNhaa
RkxLLOWqZSFqBxCdCrgu65KkQikSJxmgCYORno4HgU5D1KKTWdO5dgmi3DNf5qBCvhtGkKReq974
dxvcwegCVpG/9tcSQJYn+ZeiApo5JhheOtyEnZXAiQlt4ZniuDZ48AN3hlfOlaYVsvEQZAHxI2Bj
qtqC4fyueUrN19fzro0CsRWrS/laEWgBJ34XU2kMiW+eWTLS2QZACGvXYZqM3h89XR3eyBX17oAM
eOhZO8R4oKxV1GE0JPWxsopeAZXyawiHBt6fuP/xev9PYpAn3n1p9bG9LAJ3afWPtJi3hQSHlTaM
kGpZldC3KyjM5O8qN69e9zp/0A0dtFN6Ew+O6Zm2uU2kND2zb+1P9LfQu7jBmhV6x6Ck3N9a0Fh5
Vz61ZPIs+F/S8qt8nRnaWC2XW/mAvenSBpTHVWYypor990uKtcnTOAuC2u0tLJZK9Fg41SpjpkAy
j7GD5amwh9t3thzd9PETf5qrffmb8UxBcXd4APsqHKMz8Hu4d0RpJdBigXj+7WCAI+JLYqLMIzN4
QoNg0EDavu9HNcdmSxQLsm8+qjI8YmD2l5MQNNSHPSm63iQ4xd9rKpsRN7HflVZuCDWmj09J14+W
AGR4WyBiLwO7vPzhb/HHMXxl/BaeyL+oIztG6zKK9/XboT/48CNNdlhoC4OtWESIupdvhcG7tzLk
o9P9ZOk43MrFfdqFrf3QPHOJzf6KbrlbGHQVP1Q/Kj1+EfAoYXwdrGNm42yGvKLrplegWk3YUrQv
0Weo5lAjnVFMNGc8zyNoEDyxB4DVBOvciaSF0ziTO6wGG2xJNRjRS3ABlBwI6W9ZW1+LZquvIrMV
T747AiMjvkWKalzRxhATojsY2H8vWG/eylQ3o+JK169w1H9VyvQDBBFkf0yF7ITYH6iVlXBqcFj9
FbURvQGL9AlX4UPDXyUal7IbaL7HnO0VfudmBNBKrj8eULCmkQJpcdVmQznTcGWHFgFT/f8w5TRy
Pu4jhHHOrTxxa24aZ3HSP+UWDMbgaVvNR4kiG5PnRnGkI9pToXvdDCuCz90Hh2NW+/bObPTPuE/G
kqxu7nWQmMh47jncKUie6R0ykJnsnm6bJ9YJc9Zvg7yH40IBwAqVyzRRYuF4HJsLyLsHZQbczYYs
C35acvF75+8HyGzIS3Y/stqioRzNc3K2i/LbLs2md9WoTh1IwzRGwQvQcIsPSWTGLVTSwub0C2Cw
xgkAlMTe5kEuXEVNLtqkgKSHp2eWO/Sqz+KhwaBAXKl2y+Jf4AAJ29d34HUDZiIPg6tWLenHF/0v
BZSaNu0lwgCyehv1cONa9H3drR+uHt8D01ZDE6THkFuDbRSLjo1CZiDL9WQZyFiJETUZgYPvRRSA
KoDo0SohXeN+Qmhww85dTWBicttCuRFuaWTlzZx09r5jzCCNDIrZZt/6w6FcSkGGN5rAddSepyfR
3xrdUe+6pEKjyaIGX2JJBF1AsSANE7nuPOtJ7x4TB+MpDWquOBaQVhmjANZ4Lcb+etcQOlrGzQjm
HqiW5CbeHLK4wk/dFmN2RQ3nY64MDBjq2JGbrVYHYcUTibxs9p16nhCbaKhxu38vyiYhFbNSTVDT
5jKTQeUi376ll9HnnjorLzUDhy8NkrwaBVdKw29DxM2HlSmcaUVlRwGJGl2Dy7khGq7Nukc/gsM/
r+pZgkNpom7FKfwH/915bWwPePflZ9RfgsTg+tN6ziEk3t2QQJDfy+/vmL1UZ4tGmZnMfXvebA24
708FuHxFf7WMrODlqd4AdOYXk8JgQSEzGpJaJi5o9UrTFfVpGleVLkNwTr+Il6ZxFlGYyZA1HLJL
XyciErcztiknapOAbTBypCIt3ssYUtIEVn9NC6co+MBb5vxHvs+y3cuwVS6j+Z6xrrTtPTsB1Y6i
BciRrNUHeQSgqsLsZuK5aGxo7TF0g8FO65u6odtObx1oYFmJcZH08DtFtRomNv8Z9igZ/uGapbNl
QCEJX3VluVQI7wBGbx5VinEohr9usTfDwbZrsIrZET9c+uU5lLxl9OoGfbF3tPRC6NHnT5toS+Jx
Yq9psO7UzcrTlPYyMUzaIrGhGXCTlayVeSaM/Mlsy9pkm3CxEnZxo0tGWUoXBJioQ1cxsITds+xQ
VHFw5QcqY33NRxRlAXu4bbpttop8ZZcAvE84l0KyvWVKI6JQT4F5bMuT+NMiU3HH4xtyN7rw9Prl
dHAizF8LLDZXFAL0Ctg0aEDDeLjCL9wzb5Fv9WL9AM8FmEWCciFMqtzRO+fjIAoas2ZC4MpZ70n0
A0+xG5xuCT/jinydk8Hp3tPn/WgCExlV+rryzxt2jF/kaMypA9s/C8wZlsiRSE0bqFzcdXqwdVSn
eRh7pRA+8z45Ew/xS/9KDVv1M/4gxoE5BaptqiQ83jMoGllBtJ+E/ipZ0TtZJ1CiRREjGtXuBYh7
vMVDrMT8yvKetY+gi0CA4vF7l+7MaKKTJ4Zg871HjKaVPfphJ+q7vR2GGXuxnFR+ZCaAYfxbg/ak
6miHvx3qJBGuzhgew4ynSJpoQiuTLuk0ZjhhFOkrr9quK+1gOsK7P/oEv5ot0kJzNTHh6aqp/hMD
BcXvvLN9xh28pA0AXlPpQu1JxD+dX9EHFIGXJZN2sWZi/O04ITOQL1BarympS67IbsAw3vh4qKG9
ncLzlMhfwCNE5UO0BtU7CCU17D4dDbw94coyGlADbqSsuGtB7RQTUTR0QaXd+wyf9CI/LhpXCmGT
0nyki9vRUM1Bq49cG1+mPCE4eVXJj6HvcKiAjqGEqz0n9PIPart/bogqOTyDvwDiPhuqJPSOFICt
sYeL6XdqIHGQ7g7cDQW6UblRlOSmIeyfECD5sqp/Dv/D1KRIUdpbOkWbkU9OaTaUwYQS/o8opuWv
aSDAOcQkmvfxIjg8PFp3tOWRMzYIdzVcJGkAJRgnNtdXdQjO1tr8XXCmtjC5ONG9Naxq4YeDYj3d
1yxsT5IFoShmmSA15sNI7+xMf/9LqVEVRi18xT7qlB6p3953LHMzJfpr0Bp3q53p/3GtcgfhRRC5
114reTEs0jC/5nsQe1R0/i60+cRszKfjsExRk2t01kahipqEyRM0Cc5a30ZFEPeZIqEE9LHP7/Ls
rz+VI4HmIUYIxky3Iv4zdu9klzulpmPgZteq3LRdCJnE4eZ/gJkqGXYA6DfkNfEA2MtKMUtwKfup
N/ofkUWN79K0vzmVNSjm4kqGAaar9pFn/oq3GQlWwBwpmclUgujyArEzgrQL8lVeUvEM2nqmuINk
fxe7JNuMfuSv/7hw8RucMeCdAWKcG7sYzL1pKokoHWHSYsgRgkeMi3YPbEVzWdW///Q3zzrL5/iE
Fbs/ePA5vCMdSJ7FFlg9ho5f8zSdjH4KYuqsc1N8/dvEmkQ6h6vENPPH9/1KUxZToI4BRH9js9BM
9Dqlvqr5JHUlu8GbOgU9SNGXEDpe9JavldmQ5PH2Lx7ZBHoKn3XD3swqGUOCNDhEepcJukEnU94a
m2/eiXRQG0dlPuTkLCquFUT6WbZWamh0YklEr3y2cd51z2viMI9wnf+fgBQTbbITxh3DcoAJ9lgy
YMSzjZX1+lO0l8qJc4Bw92u988Lo6w+/oD7rHtzYBGxqsMTQwFpLL2/UA01b8Uy9nolCyJzqVrDr
OBg0JM6e6jdhnSeKMtjceXbpYORhZcDtpLma44JKIMRaml5PqntSK8wdQp8D31cj1YkEoruIYJL0
CSG2u4zV87R1eFQiknZsr4ejJLNdC7xgu9N5mdZvvHifTD0nohXag91ktZ9rBwyinySvH/IVNw08
OQP+rSXNcti46Zq9ILvyLplUJGLx0Ayb1mmLqFxARv2j4jjh14oP5eTMMix432aHY4fHDWKiIV/9
O3wHOR8mYVNZ0h0pbAzS8PYgcb71xxcA8OtDo+F5FEdWZUdHfcN97k/dZ6fyptkkzfEgdXDzN8uV
eYScPUw8Eq8r8PsJDynrg3NG/kgfsQhBSdnhX6XmwLZWl4Eh6DnObdec15CUrGge5WM0tK0SuoHr
Jca8Zy6VNkk/dfUDZrK60qix/EiK5cT3uu+sklZ/Nnzdi6co/rdYIvVZjc31YE8D3WQwTLwCDEnj
3qFL0EkvDYvVyY2prBFL3brJNPL80xri10LdxbK8immSh17a5NC894qCSsks3I/PcuaUwc7IZP8v
CwfzcnZY+bZ3KHKs/sKRSXG1q03yNyVUnpQpVM+UZik2ynGqaHA7F6g7bJgB8pGOHJUqX79sBx6r
NY5rTXU1QekyGEohgxJ8+3KOXYuBOzqYDD7UmpOHtMZ+wcs8czRQEc94pxXOvGjT+RC8xLA0j6tN
aWmI/8nU1Taax/hR3ylMvMq3O1EUcH6bvh1VQt8aQNh1rTjaUWFJ57ckqFVg8hnxh0BjyGo5D277
qZTRdGAVlH3F57PmEe8i0Ge2F6s/SEr8OYfrSWagrPUgaaPa7K0hqFBDh3pXHJSgcqcNkp8Rlv/g
5tNyt7aaEIqkiRZT6W3ha6wOKGhkJDjR5hIl+z1QK0p+2dnoXQtonraoyuGUQbQ5BE7RJvv/MerL
Uu7FzHQsGecARHFJyPVKpWrq/KDsgegyGkENUep6GSA53+PydLM6vOyiE4xEOrpLtn8CSRSIuHHy
0JJ4GEp7sluCo06edXwx8iw7yBZpPlghbMme5vtUeLc+R52Ou8h6vEXZnLgGga7+AN+Gu88NC9EZ
2orIZirazlRMXSvaWa1X0m0Fy6C6CsKPZum3kSJx9Yd/YpyjCnpITZA/OO4rEEkSTcg+nskOLakC
KCSxaU0I2rztAdl1CFsyoOCex9WWP0j1sJdD2ec+o65odCpgPbbfIBZA4yUgY7sFXbklQpG0orLm
t3nSVDbYOoFj9irL77T9nnFC+vpT84C5jlZvX5r7SEdmQKWCIVvRAX/8Bf9nQyx9UKxXQmBVon7V
C8av9oL48xHOPGnMpLUPINTQtE/dXOnDamzKCNLWqihIlcBvYjW6vPfstIBkY+M8Ijlk+WRR0145
UJvsLYl5HRgHUx5ZjAzZeZcpt+Wh6tsg8308Di2XrtD/fEzqyiDIoPwx1eVo+4gQXsHkF6NkwIIB
6zTAt4HdWz7e82t0elxS1McQJXD0tThQXzwu31RS1GpbJuGGZsTC04LlK21ITDJfRqhQb4/ruriA
QPsKfT2WKjUpKA0QfXUiJuvwt7JVfJGj0jZxKkMWUYawTWrs7w2mXleq9JtGLangX9dhyA/QEi1p
P5OIInaFQ8mraktuVCCHom5Vd9NdvEEzQp77UFRptwTBbwl92u9qcnZYVxxm48uF3lIDoiMbayjY
/S3Xw0oIyE3StHo7bJI4AmlbiTw/ntToukkxxKvK699iORA+LwtmXn7Hr1nBtux9rFxJHLa1i1wV
dJcJ6EZHTUT2dZl+FnV7NErjcArGNBAtDJPmp1AwEcwz9IJUjv0CKILmseAQsYCHZ7QpI3tBJC7D
F3tRHobWkx5l0uumpIKdDh/RGypca69yFz/S9IQR1cEo4jf80uJUAXdwrPYBrZVElst9yKgooBha
WkENyMtDPcYMJae/cfRdgkvcEd/QIPc/uHJu7I8dFA/rBaTd4TN8tAFA6gW77PQP7wCfic+khwd5
8/jofUVcetkUeQu6vafkjDauoIo5ug8zwxkQEmvbWYznwu4ctt733dlcv0V3can26+lzn6VVlWRV
p0o0x1OcwSA5onIamaydhc9RHTWNixvaHYfxwHCRAvi3nqMnwqw/7RPM1e2fapEXn/BtxCJsNYw+
HE2Pj1M+huNa7khVR98QDZCGNJojHI3ql9+uEkwzd7madkmtvKMqNNBeL2w1TnvJjAcC0sDXjeXq
z4GnQq6BDeI18yTnkbxR1qT8Ibt0UWWyM2D5GmlUCB2jmZ7viwQIRUozA/bgNc+BAGrSUX822dab
aMSE/a3jcB78IofQbPIoVbqlnU/mZyWgKuYsz6fYZ8OJSFH1W5/KmkTZwOrYow/Vnr34JE0UGWQV
/1dKrA9so39GLjS0eZqgqukAga+HdRG6CypLvuTwMFipdkWUMaRC3YaLPy2U6awnE+fUx+46Sjo3
eSeuteLSJDq0fCjaNcduNbNeO5/TwscHhRBLR0xf85z11Yxv3o52wZZcjI05OZKH2KcZhw0ZWr85
2XGaQpLSnY21U7DDarwT198/6g/a9GqKPxlfyshyH4M5aPvb6S04dPFDbuIeNjbADAJ5g473O3aX
ngvfftfNuN6QRoPVMmS7sFytOAIUPsZYbZVTtqMOlVY8N3R8oAAULD0XU7hktH438ulg42LtZAeG
j1SsN42peFpdkAbhquca0678+Y7VqWZwcL5RQLfUduQYHuwIPmXfg8KhOr1mSdXX6Pz/SjOmSx6Q
ea89fILP5h7bBMaPmMr8XjlKw+E8ALETVcZyY13P8fm+pXf2xpNjRvuTXPLdc6epN1WxkAIYNOlT
RMmAqxhQNqahD9BKNUDXvBRP0/9QXTclWHqPE4Ha/B4qHTL2oy8q4WDEeQsDA6YtLoG6smERyUvJ
CDOUVp/UvX+6KJVQLNLwJP4DH5MtlkMfw1SN4y5uyWvvoqzM9Ge4ZDo0jcg7uA4DRu3n+nt66gKg
DtZHDcPQZQPtEFME/ZmB1F4J+PvtADc5DeAZj1p+ivq/TmBRrdcKXErAu5r/ZWpW/bA0b+51KB+4
0tQ77YVLoV+fX1X/SDI78uSM8BSYmex/d26L755534F+rRqGfrMaHHsJSPWGmGTTg1TK1GhTovWt
biQsR++8WwLMDGBDhX/3lTk2P5/od/i9dpCTLSe29PLIE2XhD0xxqlrDRA15voPZZefUhkwSxRSA
6tz+Jtd1pOqTxTdU1zYJ1TQ0vfw5xVVZWRKycCtf/eURK7UUj4Jgr3NwcITPXRDMV7qpfZdSNz7B
MqIpCWcBuHmjvvoaZFx3tiTJwTt0aeXnpdU6kPLkQAM2KAf4q1gfzUUtVeGXPZ0Kam6pod1n4aoF
LezwgzNrLjEVCQ9oKzytWnYyYmpcjEAn2CD3INws/FRPiTvl7JhN893Of2IOZFNEr3lnuq0u/FEL
pLr/eweyLEPwhnsIXW6zSvCceL/oG9+cnU4vFqHw8IJmUaHOAj9ZLYJ0/bRYyt6Ak1zw52s7dY8U
EWoDpq8wLYombn9KghgqciuoWLcKq8tIhfSoweGQQjHeKPfl0zoW0pQdRT1lOhitqynGxRDdd1D5
dJ1iwf84/729EQ5frzDNyj+wFWvQrFVaYm1bGukZaILah+Mw2rJaH1+orW+kCVPeOUmC46bFfmRv
un9Iyk41dY4oy8rJwHaZI/wyqdC4ph2vMo/jA7hL6ft/7qfmDVNQJ/LzFV5OmvCpz/EhutM6VJ1W
NTOktQX/xulJLEIpUqU7/aJwrlygE5XAGHTKkHQe6LlrtIbRUr6nrwfVnu+MxnJRUg9DJUi9m0dZ
rNZqfDspOQnzaNUuKbd922D6RxeeAnm7NSpkp5sAs6XbrAHpZ2+gm2SwwrKofkL9L9Gj727Q5wAQ
Yn2USvP/TJtr/tflvH0SvCg/vgqIbN1o/PLE4JrPu5PEC8mTeF2Hq/nTN5sppwmIRD0P65lIeAwp
hl2+9SXeB9RZJrP+KLOIYJebwZUQMKpdK/FDy1huKlqilqv9sI92m3Mh16qfxgEumwlRwPQsgyQF
t6xl13pQZarneCH3n3KVuNQDe1Y1vx3N/3FO2KqEUZCqDywiyxrmYn25Rzqovi59oxqHKrQkVUDQ
ETRQdQ4ihQ4Ii2s74bY4FrmdnZhhtj0gmAP6UDqQeNLg2jgzM4jWGk2uYF3KCZDOKtdI23nnAGvm
IaOfPzpxL4czjCN42pI5v8b78C3h0cGX+kEPEA7HPqnVJKIaTlFactEZ832QTzWXnbO6Y4ObAxsT
/VIOPzxHAloZvSp35kVYEgsg+djQ07WiCX6PGye0drhWW9omQAGNxpkQE5YJwVW9GlZZ/JlKoVkJ
vE44ElW+NxlfoYRELepHDAIFeiqIrJ1bVuqjYr4EO931OFa3E2I0rWdnA3y/lD0Xk4aBd7wVFcQr
nAtlbaGPdh45oiAvE9KVpidyjC6OWI3AlMhTiBZjMdWKY9QzHg+DN90OMW9BSexy+hH4oMLLxhjG
VUFvi+KQiTuHU3wDxV0lSOB6cBdJbtvclcJi8e+xab7MWjHhx3FW9gdqDoahqs32o8pts/msD/e3
Dc75D9/Hgx5DZRX1A+WOKxFqzObQRg4xYzP86+/11mh4CEuVGyKa0pCu9+VGmlY14Dy9+z+2IRzu
2CTJCiolRCqb9ywRTVeCp0aEA4DzNSTHqDnpK+muFrqpRfLl2xnGhwe5BuH8mFiNlQqJhhb/A/ry
ht3pog+FwTbCp6+8llEcSSGteyUlK3tFty4MHHmnDcyPIX+NMO/m1jR6tLz0QF39EoJT5N9KhoqR
YMO1lAhxDwoK3XvFym6L496tjBLxp3pbIHZK9CSIE57y+ZlY2ERhSvA/17MLJNnTtyzqOqG4O8I4
QDtPKEkUmFDs9OrwHQ1t0/dU1JJLcWbjBGvJQBT8uP07vzzOFXfhGINlI1/q8BxhZCaLAp0UrWh9
SvxgMukTI1lPQ4rWay4LQb6pdFF7dAZaDRNbaYh4KX58DgpHsCUi760U8kTknWg2fXwDuVR2sazk
9st4vgD5b1c0jPXM3W1KTA9qk7MfaiQelja1aeYc5ceyfyf9xh57wsX0gvyqrvZrTpWdvgRs8Q5R
fmUkDKeE6hnUkeJW8bLvv9KL6FODUp9Tklw9th71Sqt+H9AKVUmIWHDoWqIP427q1xTzgQcfwcmO
jvb1XjJEwshTeZ3JzQVe4JLvfzfYAJcC5JDf2bOJ31hv3cLKtFqd97FyLXf3Hv/LFNXtk89xBTqm
tBKlXOXbCUybMtmifP0Qs+4Duxo1lGoD2CuaiTcEC17QSU8gptdkYJ9XQNV6fQm34uSBCT1TnCL/
EPELueOWVxuo9oAD3u2rxQyo9RNR2OPeMZCIYZtV2c78i+xKFmhWhH0+j+WFGhirFXBHBytR3NvZ
3frr1km95uV4XErH7iL0Q8dCRH48elTE+k5CAGKR6hwQvFv2m8YJ8y0Y67RfoAGMlHAFrTCHbgB8
bSCuAkkbfEe6Bo/zxBwOFuQrP/Lrq4ceTurjaWtXsBI15YGuKcSKsO5LSGV/SOQ8/ilueG/2rKoX
NvqAqMRTAxvm8D79BsJMkkTNc9BPlAhmEl/SQmN8HfOy5AXh8IlSshqHWy2IHoqN59al86aKWOex
F6g8KMXXrFyYYOOT9yc1DSd4wRN9A2H4i6EoWiX/JpcWe2lxtERp2gXVZ/hCXQHxGMg50NNRoKbp
Z3uw7ptTUZXEqn/agH/ZZCgLsTalGRd1fS3UUVS6LlGYT633dJeua67mSOz4MPaR8JXCcwhyvr3S
SAtQf76SygVcdLB3lPu+KFmlO16hXAmbpnKCANzWNlY+S5gWoljin+vHk5KG38I2odD+ZSQQixJS
zYh7kXsfqTKoWGkpUno4WR/ROlfIdbVetQPeAQI3AtLDi8StgU+1vxx5MhBh+jMa6EfaIhujJTfX
U+WFjPYovnRZKvigj9iCg2pKMJEmGufMEZ3T+iQbrzHB9ISLWqnd30HHLQlKU2Gx5Fk2aqJAkGF1
ATLFoC+YPw7XBzDyDhWuo0mQl88m3PSVgeTvNUYynAAKRNoL/vLtQX0bLX+GNV7Sw39fWZopxaHY
TGYfRoD2vVJ7OTMKE9sXWxrfr5pvG2cVg+6WKZoKDn2s2lWf5vDFeW7adQ7wwRgC5wCbarHYE7/J
Ycx4CEDWzLKszmSdm4mSTPYKV7/lt8iC++sDdaU0HDhM+37JSbanSmjnKctYJrZEjJZokEHzxSBZ
TVQctprGDf3l01Ac+m19sQQuB6g7zAqnca/TuZooefLRLQVsXfVnyqEpFxO9jrKW7wwubqvjbXhz
LwLRpobHa7C+OERFznZ8Lr8zzKWkE8mmjufm1OphIeDD+5xxx+ADv8dnD7EtRnEjAWWJRflIJwT2
+hnIdavREbCUFUCKKOcB+HoaV6lGalaHR//yBIvbGjrmbe/RnmIJPBJXtc+ltP4i3BgqyjfQGgOd
8cFWqEWxrLD0i2ro7N8ceO4gjLs9UPzPg5HLTaC0xDOcQIDtHbFWLw3HUW/K36tREplFxYOEFgEO
XM/+q3Y1fT8pszsO+i16DhTwDGI0sA7P2sNqLRDRRdR+ot/LJa4TGew8rvfWZN7beVyUf05XAksz
JS1Gf4BCSrNWQNhAQHo/qdLPngxcNByIjfa3sMsl8rqqnU0/EckQJsYAR+DsGxYDXVhPrDxg6j8E
YWkn6fOrJ5fxMq98YJMkKGONqytqEY//W7QkW1AahiNJBcYePSVOwW/9Uz1zFm1nga7N4260ioYT
P/+TFFUKkSSWQyc0Sz/xlrIyz1dtPneN3/0US0VQbeSHyNV6YnVjUbORXyYJddFOVBFo9Hy1aNkE
q+lECparvnCL07jW3d2kWSi/BF9ntMhmZI6nyTQFRiEq4PJIRYNtZ3Wp+mNjL7pmIIlfbhYl+4b7
wUaPfx1A9jBWnLlp9Ieiwe2qc89QIu2N62Am0g38vfBhbXDU12ULfhb9f/MO68STs2Rmx/H34YGc
sgGHAVOrh35F0MiMCPRzB1dBt7iQ4k0mKAkgsKdy+FOZq0zQR9V0J0bIrK+imgm+WXAgFVqm/vOq
IEsKTfc/3L2LZOZZl3i1yPx56gOXda4igIbQsVWvb+dkYWrbam/YHSCPeMuNNilozz2yTx74A4X4
V/UrO/gb0zqEhnZOAURbwtZBQoIqF880vy0VRaAObD4TuhugL3jAhEhYaW/GcRisk0DeuGJKnB0Y
c6KLaCKFXU4/+NpUJ+Y7wCWILVYuVAu4+youWqnq7qHAactUO117Y6SU8zBTXx+rB+FIZPvUxAoq
/DqhtEg3c6wm+4TojuGH6WaD7GkMzCnCF9mUwhC3hxOTwoexPtksBxWg24P1qwdabwU+zc8Z9/dr
8D484llyw2FtgGRANP8AbFPixQNivw9MkGxFLSQoD17SwDAql8pqAkjgYSQpaFhZzetTNRO3W9U6
azLHODbb3eiwK1cUMPlm6jZlurZb7HIdsYdnHyjT+DqEH/1RfGoUSQrNB2A8kok03bxnQ6dfH7aJ
R0bjyIJvTz61DC9K7juiMhwFPYXKE1xYgXgJbEnnoHdqWnTPLJTpgzCJrt8trC4UveshgAI/Nb62
zSo4w95Ah0PWvQhYRD1HReWuvap+nkmwkukcelDWHutsUaTw0Kz6dJA2Rk+srZ2X3xLhjVuCsST4
coVNcyM5lAeF89WKY5HhaGmKK32dAH0Rq4uzJ7T2Zhe8Rqwi+9mch0KsXNMB3Jefzu9Flwb/QP9s
l4qcXlrqli5LgRqDsU+QfZd5nUgl1cL/+CnzB7sdOddyPpZPHUVrOONeJJ+8NmavRTZroLW2yYgL
ZHfPFm6+eAd0a3GSuPZTqI4xb2LDS1H0tvkI4gWTCAMAqZaB4H0VaTx8VsoeyiamdlZF+XmP2y+d
jgK2IQwvA4ANPhlrpCxvBnLa85w4+9WCiBwo/6Kl/Wus8Lz5GqNlhlrVmxaDBLP5ssh/dc75M5K6
oddzUZsmnbJnMqC6mxFy+qAiDZz0CSIOTLrYuZ5nklViI4h39Gg7soH73MZSYrU5BNjWscF4510c
btceSHBlKH2/awOnJA+mYClrrB/OGwtYmeL90IGjyGHQBgh+WyQzTryJhOcJNoQzzg0+g+VzWug1
Eug6sFBOihy3Y88SMC8oDBCjicy0RyGLhgmIw3WAtWgun705dt4DZSNVr0ywvGjE2J04y0GOWUIS
ZZMgu5cUHpvuDgNbdNFMtJFgI0+/pi1791dW2LzV0gxD4XEokD0MPkODrI1zqbz3PIEiONBvxCi4
BxFSq3xAl7ZtMROu6CAyJNQD4c3ahgBK/XB3+Cb/HHZLzMFtiLN6K6zY7OfY0Ac7jnu+M9yQWxJt
5/iie8gk2pFdr3u8tbWpumJMg0wRfnfSKgDnwXk+Toh+tCDb5pvZjWmmO2LKT9G/JdsRlrzSCaoQ
+IWwav0zLi++KEuE+sTL+1BT4DjFup+psd9Uioy9qW5iPLnaloI3okxWmUCgn4LWxh2zXT00Fp5G
+CnnwR0diBhLYc9yMi4fidb3G81HaivUL0tu6IWZMSxfBYDUHSnkRHcKeHBURmPd6wTr0zYKc7ze
RCKhyJeon9maXk6m2OzVvWUKaRIhI0tsbxVPLxa/3FkDVqnxGwnsEfyezob2dCm65AFeUY+Dp6lq
yv4m0dNLksd3vFaBTJoPe/cAnw4AkSQ1SkFgLWwgNO5SYAGF59hGjLZgpKFGMB8H2lxSsdUxP7DY
aX/bdQUnK9erEPP85DiEqZRldOF7avvah/Xw8Dj8Cwi7RZOgt5jRrWuvzZvFBr8BwuCGUIeLRJaR
aXF2mWvEY7HlbiFUz+eWfFYg0wFR+DNNPweqfJsYD9L6E3uPqaqoZTHyG38Sd60+xjTcgZjXgyk8
S6WvHQeJ8ktLwfImugxaQmUwoL6cfAY4S7jdUDplFIYfS0k4t6cLa5OvCULXhwDwIeW0xbcrFPXS
J7F0i4e2PNf4OXUD01nXIZ6DICTKm2fUJaW/9Jnk1rNezW16HENmhn35hOjJG3w65EoABcthpuZr
GP1/Rl/6dJJhZAYJyjOf2lqNuKznlJAv1PtmqPY7fVCiuLk0d0OFG510zL8O82kmz580ixsAvVqK
nbJPwTgbO+5lQ0v9uE8FFU/Wo5FnipnaHvboVMMMRkthmtx7xG48SrSZ/nYMyrK3KH8PhSLFncin
jurXrgRqEaNvCBtqCGWR9F4Fw1H7h4UkgsmsvF3YT797BKT6HDiW05K1gXLqX/YRxKWBHUHD8LsT
e5EH0W43iy/rWbaImaQ3bBWvrw4FKi+xX6b3/x8qtHBrY6aMnRnhqoyuVtMr8Ul72EduemHjMvqM
EOa8X9NRFbNgiQlGkA+MVKBfgiC9Rf7PHPGEHMB3hN7Oa3nUzWLHbsafwz9gOjaunrp8Z2LNd9EX
8hqgkOs3xT/TSnsXIZjTAIETJgUFXvik5Or08yCsRc86/odZFVBpqIE6hwzjke1kyE8faJX7sFPE
fxyRgcbYR2xV4XVAhGFs9++R7YYvgwz0hEUXmeH5YeFeUQB0ehGQQ9HIbATz1Lsml0y71M9dP9iz
4dvwmXTzAFUQZtIvhGrKhYxe8h97ZXb08mBa+hmAp+5V8ssAZbRWv2zwrlXfmn6ZvgoInQV0Mtix
rjl31uDVrAmm/PnaViZtaLI/DNiQFxBTW7YSzGaBxHuOnQ9OV+nELztqpQZV5juDMBR8b8ALU41l
vFPbRqliXhGvd46u0Fn2ZVG+uvZokNPcGCV/VlTo7VFPxA09AXJhZ9qQ9lhwmHfEqD2UTbCLAM/E
/bMF+C858Ji/e64SXBkRaW/b81wrt0Ti/XlBPayBpv6pSH7LnpeBzi+6qeGJtv+JH9M9LpSMXhyH
4rH2XNExPITDuWrYLkkQyGNuN64OspbudoNk6AgjsdGJpg7T7Rz3OxbS5ruRBfRRu3rE290IBvXH
9NiQmhjumppIvRMjECgzpJe9EKtOPWnP3SUzYDJkWIcpysbOp4XY5CK5C4qsSzxrMbbTXO38Ox3T
Id2i10XEWWi9kT6/DeB6YJY592RiGROvXuqkVsFBe1zgqZB8szt17OEeIne4zam/LUm63Cmkzn+B
xwBgi2eYc+rm+xu1AZ2fnHZT2izwPui1aruy0LOuRP2djOrxJESQL94svg037w0Ak2qWDme53GwA
1z29WtgJR0hG1hhMND/Rwl89KHesSPKWfTDH85msjvN+q1Y8rxyo4FVhVtyWQvvWkCqkmkCswHlk
55xAzovZ86WnQpa17cELNCy9kjgh8D99EZmlsgMEknfV7gyNqkNEzwk4oCQ/6d/SXhs/cB+loSVl
aWiSJSGBWKlJLMRC3C7pTAD3xN2Okg8G2S0JRD7gYZGdLnynZfOUOrNvN1zs+Ui2ETGsG/wfLPcn
OkGefGtwWhMWnujMBFtFtHP4mHybwzzTa/y+t5xe7/M6GXfyqcYsdzu+yMG9lUlVzJ8MdySpOHTE
Qty40UFWZHkKgeS4AZVl0zlOgyVooFatx/zksT8lHP/hdENj6+fvQgKlGRsDPLY1UqTs9leysHth
930nfiGBidfffwornM+5dviCSVhUWWNHuiKI5T7d6YaoLlu/ndgE40fDzfdW5ydKTIAfzUzrpJk4
Icom89STmWkT1lYOZ8qkE/3dTyOdfQxAvlFJXkdzpG9SVTMXBd2uYNgSDsj4G36Gbq56SNBPU0x9
OtLhYohrjT1rhiIKWf0/PWuYdHKyJcIMw0kOIgmS8mgbWFAH3C033aJXSMdk51f1i/C0iPtdaVJf
sBJfiiTflkZY36Y+qSRWfd/IJxt8ppPaibVIaN0uKHRQqQ8wXCz+vKKdmAVavYKQ7c6N+KTAjdnK
VYe6jB/IzgvGDdbgCSjggsAo2tFTP5bnOFlcNJnz7loH2LvLKXgj0OXBNgvIkmHQK0LV7lZVzeCX
kksYCJ0J1BnVvnQySCgRlJu/80xQFjzIpT++71uqJz0tyefqDf42AHTRx6crrdlJfGKPKzzcevNS
Bj16bEKv5t0122/WxI36SNqmiFCXOeLpDugsQrsquL03XOfo5MdG+tr33sLVpJqoDy1VQ1sJNjy7
vp4wZxel/chmMI61mKZ4EXEcmBSfpxKeBT3EDH9q+dtFRxNHF9DzUu+OL8oXkmhmYjoZHDB5JxsV
XZlCnoef+C1K+5cbg/SWwgoVGP5qmN2EM6NR0tc9r6I5gfSj10t1cqg3dgESKerRj0NjeVv6NLMZ
wD6EbXoGOwSb1oS2lidNRebPzNXnI607116Y1gfn602G/2+GbWnq9GvTI/14xulmc4vk21VLKTZx
bj3rOpQjzmubsK6jkfPY6ZEFsLRJKpa7VsF7EWqoyZB/IFxJeKII9HBYO4CwQAwHdQk3IX8lm2NX
WJSQOOP2HUv2afAJCTzG+WUU81CTMOuIQP6U3Xry4PpjvskyO9OZrtNgr0dkwwFImvUVaCxs/VgD
5D6hMY90aWnFYoz+/sTHBjcor8orKWgOJUfIpokDApw0b8hFqX6vpM/aDbAaTt9NmeoLSAQlmT2u
rHTWRIYvBdPIczYTrO/GP/J5VEkdVvBotuWpCzPdRYz/1Ez4UFnnYIUdHPJSJzjgYetGgk/WVAIf
q/ak/yjaDaL9v0jw4pXt6g0cxXNH08NhlcF5wJyAjy0JqoN4UlHTi0GBUY+MZsYMqlhnvKr+I0WA
2OjrZ7899G8YeV+STmka1l+jIIBzocMCv3twwSNGbysokEruYq2CGHNnCyXxilfdXGWyo8iBHg/7
Xb0HeN/x3b1tfJFAgGRuRPsrHlgqeCRroytPmu/PDVyg4Y8opYFCQ3kPQ9geVh3g6Q5JC4HIsK0h
FST1AL4J8/NxY/ThLOGudVT+EIvpu9m8TwIKO7CeuYx48SeU7I0d++35NCqKfUeVBZIYjjUTxOh1
J4bLDR+zo5ir6oml5Qn76SEjf4anZ97Hn/Km+RfVEamcEmxDJ1K+Dh9jI/k9ia76zaqpILGA29+A
9J7xeSdEf6Pc5PmpIHZbCQxsisF2RFuytqfjDs3soPF3DruU+ES01Vt9uAiqHDYdj4zCCCBozH+h
CrroIRUL3Tzpk2HBC5ZN4BhdNlSvxY6kZPGaarLHzjQi/Imwt9BUGT4zk3+xkSWpev6eteg3tSo9
8fsNc71TkdxkYEJ6XXtAu2k8Z4+eLG7m6qJGOppf2QwEQJnegpvZd+rIlAuorva+hKwgOETKboMg
INZr+6mUEekgk1fJr2bD8c6TpJ2g3xHB1SQOX2CpFVY8K4eW56yshDHqhPQ6irW/quFMHJ+dcMi1
0juxHb4FCkhIkswm7V6v5mrRP5IBoSoN1w1oQN6KQoZ+O3jcRSrSMOum8XTIXbN/WxgXrgvWJpqy
VfUk/qgquRmpiLFGX3CeMdUVmcsmw9Rb/4/gtcH/UqPbiXpOh1S2FmaKgx0VXrJOK+OEmYCnOkK1
rOP9QpyXLP7vRo3eFW0SD6wGQOz8szDsKgVfD0TqcMNRApc3TtezVZ0MZz68fj4MV+MNTQXT1AHL
XMKzaDtrrqIAe4PTYvXiov5yb0QiyDu7lsVmOcx2qWCFKGkVhiHHA6ofpLPmLiwXFt36eqI+3lCe
bpBgp+KZXMLnLqIlHhX4+oixnfws4oB3OkD7ew6ZPk5UyUFYPFy2lksuWuA5Xf4m6AfZoVhimstz
aV7MwGxHqL6x+xlpzu/qSJTAxvXfpl1h8KWTo0JRmDgdsxYYEGLzBzLX4cqJqPCTyFoGKwOGvwz1
RHKyGgnHsfDW0wpwkblGCEWLtZsYtRVQQTnO085Juh2uN35/MupnZAAZYcUGQ0Mj7kU8w+s+J86U
yznkm/DOZD2MdB6fR04CBAwzcc17XtD3eGcdhXx/UDH+B+Go+9wq5OmO7VKr0MtcvvjRGE7p7XEe
6h0weYZJz9fOpbfZgkNzZlr6dLZ4ZvWNKD4ce2TT+MI5Ww6MXrk+KHzUPjv9I9ormaf9R4iiyG8D
IrlfycqewjX/l7MoGCdP1foKenmwgri7e7gCQhm4U+Dj1WvyfsIhxgxrZrLFi8gzQdaBW5BG42CB
hJSGreoylb3RLC7HXwhVInvuP7RiQEDvN9VGW0A21sLTvAgDxNkqWll7O3HT8mrM8Lh0AtWpUqfe
28Zi5iN9hQUl7HaW/XikHDKa18SAJWhncpO0+9QofqqZ6lCjXRM6pCL/O7x88VmZ3vn3c3tHZjE+
TqOzegyjYh7KF0pLRQN7FRdVZy4UbfTw6ne8Sj1/AzrJeZ2CFLj/UgtDhVDgCEyNNze/lIucTW3F
DMuTiTkUe/2MZMnvVIxwR6urPbLQnaJuU+kdX/IGkwcvWOOYYhFo89HIgVfOA0vRAnuCZVwYgJbB
0F1WEV96ig0I7q4qrLTSfPcgj1UuiBStIOzxVeU+jnu01fX0qVlhD7kMM1XVaweJ2uGt/a65OH4R
hhXSRHCYrI1EuYcXVnuobzrxekeLtKmi+U+YNHMX56R2m0FQ4B8Z9USlIiyZCq32+LRSnrPcG6gD
W8FYMKv6nU8QhZR7gjWPDd6YmQ6CiuyRr52XHJ665HeEaU6JKWXCJXaVxoxwfHb0VZkublYb1b0B
NHjo/L0F1qc5xcjMl9JzAzL0gtzoJ/EZ6XSo1y7VbI81sfTgkuOHuSe5c7jSUn6XijkhxuATPlN2
SwhWPHSyCJrnx0xmFPpMplQP0lvbgyEV7iJKt272WFYGYqz5NDVkopy5HnE++Gxc170M7lEWnt+O
CpSpwiWnLQnyXRAwvt8vxvWmxipspg1dIXZTYVPtubxJmWirSOG2FtqeZ5orfX6DHnBZ8AjyBl2e
ZDB4Pwr5Sdyu2soXz7q2Ei1Y2onZsq25FgMeqq8+IjDZdllnms/fKyRIJ0iuwjCIA0/4EO8ek2iD
TUEgis/2ZLzG/7HxewLGqGY3TrtJMOP/5CzBpx1hJ/RF5xWghgh517s/qxV/7pp2ugmfL83kCKOY
Kg7CmDem0FcWSbH4+ow/b6b3Oetf8jHfICsA8AI3uU03Qqo6BcniNEPZ2sELHhxV6zqhwtvYPJXa
lr0yERTnCzdznV80xbl0Lixq5kaTtCrpDVN/sN2XUUPni0AeKZSiQEsUiDjFx8aBQl7CetpgdOL4
kDv3GBJLliFJ4pVV7wnY8u83KxR7g5Xrmj0j+9jHIeyaYGbbKTrET2iSLhQWdScajMVq0Hy26VIO
XjaB6QIYpJIBW3ye6D9D/SfGaNJb6+OpA6L2UTeffokjWv2fYHDTFjOT47uzMY0JFmNUHnDep5gz
/b4eJYDDjbKQQ14fUwV78+aOnpGpC8j/d26WfytlMlab2cOQmthz2wt0qzWOwh25IjwIhd5sqmt2
1pivRRXn3jvU5KwcpW3orwXHz+gH6XdeWaHPF4BLBdaXGchbWEYXFGUOVNu0wdDYXmFV1QN19qhv
t1sIRUMLY29GYJjfITBuwpsaSt1hKnMJWYvCBB15//1D1DKYnT9jSGAKgsghgeo1PY3AKir5Egdj
lXh9zW8ioxXy3Nz+bzY6eQXGA6ZFa846tBUHxAGIlkNuL+TYxsxWGIPoNCeAIp4qv1AIIoWsrDEc
PxFMuIj/NTsAF28jsmiRyzwfNWT6BJ8JFeKw4azbYulyYrbdTF6Y8cBMxTE0/BecDihDmKJNyxZn
QBdvvFYZlmY/v35duA+TitrGsjJH3CKSgq5cpNI+FZBRL1tgsd+uQxHCs9g9seYjyCtaq2GcfwNZ
eYa0XzI60fR0EqmtyUzl/dANlMpvuXVwLnL1WkC+4D7+CW0vRUo0DBR9TM+/MdaUd90VRN5w2Qta
Y45n7aPbRBJR26piPrvMvPAc8OxlqEoGhC2IkGVglAS2zlIKkWjDdIfu879SCdi48SS64Jo7NZeK
BYiuRjkOhPlGjqtdAH4VKdxeCdypx1KuRc/1ORaK3tXtbq9nWFlegUoptjRYwzBRl0hzInzjlZmh
9D5bn/g2HX4JOWf1wYel+ws5BWTfYS0EJx7aXj6A5pqssUlregWcY1m37vZQCat5fggchXWBGMkP
nYBDTnKeR6x/u2o0Th+pSfSPEGdYXKUo1KM/Dc2OE8aSnmuJV1qTSJYY6iNHVBQ/Zg6ucWDy9Mor
Xlno4nnpUQJsRpKfsUhh38dgNGlup3uSfe5C4HKGOpO+JX0GnjNZFSxIpSWFBApTg4nUcqHcQXPk
6w50XII1Q23aesviKeMpcMwjP5zouQAJIM4t2zavh+UBdBkO2EGJ0Lt/jbxEPPHvPI53Zj1v2xNU
oULqiDcygYurt9ccKdqcfwn0QnpqV/Ru1BzQ00b1IAx0vpJPjEa4EBv5u9n/sG4ZlIZO61ejXooU
qB36f9yGWJsTgROHaT2a6brECZIPjFO0OkszUa4bbXWBPYPih9O2AGkIS1pqM8BopYuBgOyHBK1J
AtXPzWOECzr1wWGL+BrqHJ749VsddVYFTXW+r1eBoyBqa6tZyPHJ65VxfoCqv84xuYZPtWuGw6rG
Yj4KzGnozk3NL3GIB2jDs2wfAEFr2FQb/ZYBZTrniEmcRqDy02OV4ZAKoxGPyMjuf7+kg4gZ5zYQ
KOX5aFgRzYNVSLuT+vy8r4QbgPaFjuScsdSmYCOyYb4a4LQderDo3khtTi8HDodd4gjsic4EOawQ
2j+rNer9N8oiAHAtVjo3/3wafZkhECVdHPTN3irRcWHZH29Jn55/R4wbyRu9MvZnX49ruW6QloYx
qSx7wNdKTjVUyaOAjHwrjs/NeGOZl+Gh4/Cd8mUu85Qeh7YzOZ4hQDTYFqyWq8i6wAo50hjZGS80
drMaLhGrmNG1w7pEefhHFiaPfnFkpOKTczMp+ERF0VmPp/9tEFKPn1yaAnGqN74stZ/GTZtmNQK2
MEVER0PF8HUBwyhgL1h4FP2Ytn0/3+0L3DMswNslg3IUqLMYIfv4OWMk3iT1e1nrbqUedalDPklk
UhMTAmt7Wj/4QVCLcWTbizYPt3GHnvm36fZvFmdnnJ47CFaa/BLWFFrIyI4r0gmEFsG9ErU2lsyG
srwCczJeA6q0p9BFlXqw/5HxsKkUa6eRN9yf3gABgQC4fo07OyVuaLNig2QCSswZZ8nb0xqkEQUJ
QX+agyF5cNse61kztN/Nn5Thot1GetlUp9wLbIiiVhn2lCBaNrRohoea9n7JpbXIL31LDTc4vUbU
8vFgpqUxBKRIqZbtdpncKON8gk+J0SfJ26xMSJ4K920EJxK5rm0o7LL5iQwrc2tmHkvWrGWVAKBe
UelaF7Wdp2MQ8EKtoj6FrooUTXkp/f8u6L6NMtTjch+IGGHA10+vvOeAlcIwbRBJEBYfGl2pnuux
2qmuUfWs6ai/i5lp6y3mTLYNjJRGhbcyfX+QHGqNP9ouhRkf7zjo+7iCXCTYbcDYmwOYz1RDN01n
QInF4UoFklxuENTnsbZiTXOsAIFR+Up8IphmI26xRi536ywXJYNdRri216kjApfv93dLq/oAUlAH
bdHdtl4AaVulkPSTWPl/dM1xcadg6tSlged0tBKGTmYJlKWw54njBVDBfj6ziLrxnjI1IXBFgUYj
gFrsOa8SeKgPHoAb876vVFaWocKBQcPhiI5MiCDamb1k+GkGnh6AeX8m9C+QtHJ8Hc+pqCuzPjTn
7cwhTbsy3b5zFd0lkqCohdmU4lrlab0xfl4Gf/WRfpZUVPfUrH93fHpuGTCMKSWIRILQF05o1u7u
X7bWCLte9rqDaedKqsvwyN19EvIAhOYtM8vtNLgph2pqL+OHVJnKdnyWkwkAh4eAQlQq/s7d6sUa
Do83KF7NfkWPVMd0ZW1xOMR4P/NnNvO46HsD5BhFo7UBy6R2NuNd2VQTgJpLJxjBMGGH5kv8YJF+
wHCK8pCMs6Gd8HJxhjsKXNtKAblJ6iZZ13saerWfgAgDS1m/Xa6g62j+VgCfip1irAZqeqgCMAOT
aoiF9NsWf4uYGs4waaI6LRxTKodeeIdA8uIuCAWmnMeCnGdv8wqu3hP+OWmJxaqkPejHWhe5WSuP
HAGtyWdF+Jao4KQE6xHModHO7UFx1jAn+Qz7vdl+8Yf6/aFtsCQrmYim+Xbmg2amU8c4sVR5CYbM
Z/60fIoN4850QiNVSf6RnEmo9HSxQXEN+29pgG0Sr3GK/0+BVA88oFx7LgnyJoLy5gALJfsD5q3q
AE8TuGHzOpkbT/X409CfW4AnIxaNeBn+iPdXhK5sPMOHtTY6SRF7pOZ1CAqp1xHMbqHFCqOn1gcA
9EPyJfuHkIWAC0rzcUkksZnwHtvRXlt/ZuI43x+ZVNavhK9szG5BWMw9yNoIiEuyOZSBzACAMfDt
BFcbZclHIh8eytRVk/yymfI5nJmwSpLGanmlWCZRixMDj80Ky1u8hcaPqKJCT7VhdTcL/yKHV9Jl
+nu/T34fu2ONNZT2XKK6wD1UM8XRZUQZlkg6BUe+oLAUzuMGi3e4yyCQo8HrQCCJLkPEuTR4vw4T
5bhZZZtWvVBf/8uupzHbNbU4xLj58VfmavJE9dVsiallwEAx2ix/bWIK40rdlX/lY/O/qrSI1usA
6Sf7nPkGVma0UWEgqDxbLp/D8vmvxzWgSeuaqL1/wJ+Af+G9fo1j/tnL9VvJ4mMEtuDuOVbXv5hU
zU0nP5+NoO8Mu5FllQT28iVtMfWt3JoAtlO02PD8jUIIrO7j391DTSZNia13qyhHPJkaeTH3hmJ6
iiQLtXosuaf3/yfReud7Sw4DbHu8ylqa396XryD1sNaNSbNK/c3/Y4HJUf3+wJEW6TONW92oyMjA
L2jQN4W15w6Jl0tPaetcMzpFxoaMZWTF0wVqRZlDXlmwiNVPWTgVmSSvnz3PI3oV0kFmVN/KCBRj
qO1Q7IxpPxgmlbnkdyuisCZH5eYzOaqtf16Y6Rx21nY6dnxBZoMkwsXxYpc00wPLTYJPuh1vklAp
FtnlW8gW5GaKW0KT2ebpP8D+KePDJvdOfp/3DLtw8QP981ja9fgJDXnMBngSR/Zs8aM65sAAt1L6
HrpbsXVfqd3tzaMD4+JtL/YrsA3IgtcyLksQaAJjUwUPBuHGrE7uwaNK+TLu60P193oXqfd8GjZU
BNMXGpk9OwUkMttlHHC296xLz9w9LXmnNPVisUPsYXdzn0fQBFwOkxxN3dxkG8eeMb6N9hDVg+kP
B3BMlNjT32T1VcCExF5svWqIaxcjN6dXtdDfB4VF5gQvEKcN/IDloTnmO/2QIr354d6fuk7qIqCZ
q0MbLCPg8jPPDY4k4+hkiRHZ+y+9JOEUi4Js27tsVdYEzrZo1v39YSxyatuZwM6Le88hBbWKftnV
EMw+yLF8i9RJI9oZw8E9L+MFAk+0kNl3MvA0RAlBV2zWPudsd9V8XqKZI2AJAmEBRkBzUjLeF0XR
OCqnII83d7edpxVbgvrmStxaTw8sOsdLXNvEHbxDUlfkUP92b047Cl3skxzr2MFVW4Xse6EZWAlG
GZrhY6zAjaui+hgwqyfXz4zumZ+fQWngF19UoddIXiBviSMlfjzh10JT2evD+m8YzODeSbzUmaAd
AAJ17/MYa7lGP9Gh335yZ7Z1u+dSwJAi4WAJBDGuYQMRdBOiFUNTLZXkNmXde2Tp6P56DeAok7sm
32aFq0SGZ79oREcToFXqfhu7mUgEPKjGU2q8i19MiCN5UkskYkOi2oPQ5I8KkogWrrHSk9pKhoYp
DYkHze5S0ed9TNOPovEefopbUQ1dsrLw+okK2nDaQoqVqJepBjnQ3nBsq6raXnsd4bq67J9k/T9q
jDRM0V45ipGw2APQR+D/dqnJZDc18bNGMXRvFdhNM+iROFIuk+DmakcRjWeRNzBM733RZN5hqn3C
pDCSaF0i5h/vkJO1OfZ/IF/WLjlWLZZ/TIRCWcbS/yewsI3YVXA77W/IXd3f4jUCCai4Xh+WynfO
07kEDjqcbf01ZaN4R0Ml4JvEE9b1YAiGY+m3n/bky4eObQSFj4amqNycO3swZJh+e7KozXKhrtPK
iapexq+fqB6sardFsrSgy9ry3rspsXnqaVre9RjdTT2614OizyystzmJgGl59YKUQTe4Vh63/V3R
40wcVn1Di7KbBA2Us+VV0Gd7sR6SgXIZ2oUK7XeaiFMcvsIBzdZskGSCRiTY8JqJ+pLYZr5R3UNA
oMftn3rOMnMq5yhT1RfJoIT5gDFFsBGf2XQzz5UGaogmBdRi/693I/PsMt4s/VGztUnI8828FluK
UMJOme8nqdK09fyxQgUYtSfRZo10EKb00ihU5y3DzWxFOBTNnpNDaJBF2NgHDsdB0hau7NfyBvyR
U/bYxtMiBznHoKf30l7TBC5EeItdzAscfk1B1BcdCnr76OkjlJaj5OPDWenAE1ab0Ai87ETV7twb
4Ntg3hqZyL1A8UgypZGm/ZUu8j245ewFeQa54GXXE5zVJJSBtPTqncvBYSqFQw/BvYG2Y2UL5BfS
QYh8JgweXOrTF8oS6JUooiJJxS97fGlSkAXHPnv8zLoeDSAisLgbwx2cIiZD5lB0rtz3/dA002if
p+sjB7uMK0UxoNyy7P65C4/nXooHiiGR30TlHNkcZ+FC4c0zHZEvfbckfGqvPO/QvysoCMvA8kTr
OUto57wurSzFzCJLz6/mO3uVUSNslh1CSHvMRTz2P8RKcGtwSFgHVV8NVWH137mCVSDpQJkK+SLg
hnJLWpkZdiPM5VeSiZOW2dzn16bfnIEncskQkhLwtIx7/LsxhTEu8cGIWoobeCo2htjup658bfBQ
exVTHyMAmVwhDxalwOjxTFGsXC0P00P7PLwmh5yyK9Oa+FjFaurw76mb7edodicFEUROXrfeAtef
M7q8709asGw3s5fqauYtW3FZ4hsIv2wap8MUrYQzD4tj40PSxwk6jcdtOrQSmBcWb3wB9EKZlxH3
RYFwRPbvwCzY17oTVnon01yhOjcEMz/uGq/4kEHdVUD03WdiN7AiO+wpLKZJPljH5EqUA8+C/PiZ
6NVvdOWtuO9kdAhjh/ewJYH3t/cIgP5Im5Ae+Ca3/mchAEWgRgqriI7Ia1dbZmZkwVJ/skgSJHqX
X8Zi2kT69Haok672EL0nwxm8QUreaY+fcz1I0q9RiAwP6VPdj5kZKOagPvKmvA6ECNFfejgw3NHJ
30QUatiQAlU6ADSmsoecsZMSBFqxIVSIq25AB6HS3vwQRepFYvTQHvstt33TRZyXgJ2mxGwoj2vM
xGHf3LVaTdg6msgPuxH43JbmwK74iG5DB78QAspNEwFQqHUlLXrMnh4UCu8MWi92LYrgomtv8ByF
eGzZ6qdl00buAB5wfyk2jwIJ0QeteQN5dxKH6aHoqDCC5I1Fxwve2RIv2I4PwQwFVlr/MgpZ6gQH
XFgXVAUu+DWVxyc40AA7EdB1W2qkfiQEkdSKt0g2kN5bjYf9nb5fDsUGh7zRRAjAcX6vgbFXDjbG
syNHWlAQkIxSawvZ2Jk9TcaZgobMIRc4yaSwtpYygo0QdZQ3CHYI623+DGoiE6kPACnESK6zlycj
93SoBM2fhknaj4+5nWuwsSZu/24BoMS3cxHyt9q6ANp/76FZin2j/iZS/RaWHxVAjVBhfuGmikU+
MITaMO1E4iCCwh2Am4egxXE1mGV4lwHQY/DesHAPDLrTkBRBNdeUlEXX5IpdnB2M7M6t7uJ0tME4
0JDEPFjDAWa//lqE3zDkm9XUmQtUJ1hSida+clJWcBANG/dkSD7dtYaEYofqvAlj0eKvVWLP890S
s109T6iMi7/Gc2kE7QF6/3PJORRNBCtbz5rRLkB2dAqoZoWlJbQ9XThecDXJ0SghMz+jdkYWGCHq
2oBCiteFncUDc0ilOg7gb4uslWKKsVTATAj/H755pAvCRRP60AVhT4NyTqNV+QAN3vnAp2zZEkQq
D1Un/3CREa4DM48pnNM60UHE95r+xejvYnvNZpd9C5b8li7LulWho8CzoYYQO0aRiZnLd5tFbkQn
wOKUG1SPa42/1bud+8xSUtJmb4iiNj/znR/9ewFZp5Kob1+jx4PqS0mWRNHYKCItbv7NfcKRrPTK
GtRTEvxeYZNSOyk7Esgk+ODdForfynWXLlrA5PkxFPXuNtKAeAprNGcI5842ieFrthYFx3SW9xDS
1J3VuzpFGACAw+01TjykFADhkuu+tZoOhg/zPBGmtEIish+XOkQtuObUIGfQ5SqmAk373QlIe9tf
7pYaggziNADUa1+G0mWUhOUKnnugf6A6qMKB+c0m+TIy1+WHEerPT97z8J3V5lhMxzRbNK7YYU+C
/5u4Drta7gE9JbVuI2euS1HdsGf7+rCGewK8Nuw9iVU+lATeERCTSfAZhh5was1W+Z9SoFzoAN0C
IyZkeboz4g8/L75VKXAf894s6og2gzco5Qw2KgXC5Obzn3BPa0GecGk7lIkcsXc6dvtYtjv5UHvI
3MOs5YFJUa2IZkDI4cHDQVbVlNeY0HHpt2dcaoFiwKChqe8uMXOrilJpVNGvFPzdpHAG/JsyBGFw
Js2qhsJpe1QsNNVSRIo0DbF1Xx54ZtMmWj5GeEUjOkzg47Nucf7cDxQw4z+bmU30y1TxRgn2aiBK
c4v0IXxl+n1P3Hr2oUXWqy4SSyoeWGW9dYCNhOuwagOcvbGjEJq2kwIa0spzpNh1qVOLw3P9o2vN
38VGNWN1PACVx0ro6PxrdgG1JIBj4o68S07GAdTxdMW5tl5kRspsoWMpdArFEiT/RUoj348AzmWJ
Q+LAgGX2dV7cX8onAas59Yu+8jgmm9xchVmk2BVmVK2h54c37l/xuGbLlBtAaZvRNUHd+9KMYPV2
DUGisQdXC2xKRZ0bcseeQU9r0j7j00vSXwCOahiv92Izs5SJ5JJB7CKY+lvybpWSS3Mwt61s+Rw8
ElX+JCJ1MwUaRjXmxIy5i8o6wMOooz4MunsH+H5EdmXCIaQXRoevVyQI/WKcWNBvZmwmq1s96LC9
z0NLlB6yoqXY4RtdnMdtHR/5jxKZd4b8OcXTK9D9UAWzRFOsIM/vQ1kDdU55zBDNuBItk11nx17P
vqjyuS8BIG+l/ZKR7X5waOTAnaargVvlJo8neTOaxQodgf8800QJEae002v9vjl7wwUaQz75+d05
lLb1th708d2d/LoY96vg1NKZuv90KykcPtZB79ucj+ptYldUgvd/bKW8NVGSbSosG5wYJAidYzPE
RUIrPJnOS3KeezqGvLSGWFY3PDpxyf5RDYM2wgLlm907L3u8TDwFFQHUzT/hi00t9JlHBzyXWuJ5
f0fLM0ZFJWf/2YBYZ3YoTu0J4ogS/L0HNp4jA9aBwLu7aDeFYbIE3Srrv9DT4Y5/+e92EPnKl2gR
X+g+epVpItglxlzXSUwYqR25t4OTtWYAEkliGdFotKjF79w9xcKbEo/kaKr5Rx+5P06FXf5qSVw7
hVF0bE17iY2ZBF+EkQ6uiJ/yB2x9+Hw+l/6yVIDACN4wciFHRE2ALGmNAnd38gUQHPYze0P5t+YT
KBhMZEJbakid+FkiEZFoBcnDuszYD9CDlDyFFWej82aPOoGI5AdiM3X/SEen9zJr5PfhSwMxcNAN
Wc3JBIE0DX0lsGTeU00QQrU9R3MuRJt4/g4TSH4kudC9w3T2UQMhERYvWUoeG3Gic/RNYzaU7sGq
ixBOYoxhFcjCGqfINziCxRsesgucQvR6DxyRpbP6w4ht4sETVs+GjK1fFKZtv8bzt+YiqSWGNET/
S47zNmi9JckXqYLJK2S288rGjbwoeCo0NY7UYIKP9hs4HMZU+boaC977FkukvJQZqNg2+hiJdpQo
XlHkzeOJPoU4lJj5CQJz1GW/6h/Zsk9Ms9F5uOXV8/aeOZwJIWdyhrOuhtgdZY7MQvJ0x8xLL6fT
VIoPIUxMUEBvtDWDvX1Kjx1NgYefeHboAWJiOX7lqVAHO+SDIedqYWBy2BTD6sQesNhzmLPxueb8
S+f7Z1YhN99ApLtykpcO+MH3bqQSmxhN+UREFtnVQm1tQkpSvQxDryn8FWkZlcIapS3ptVa2uZv7
sl/tUxKSpe1XF9EZ++GxgNO5fTSwy2ZSVrBqY5GqT9etg1drk+qcFWm6nxlvHDUYucW+q09B8mFU
U29sGuMwgDswRZx/31BD9uVCoYdYv2Gafnmpi03Kn0XFSleZN0cnAX3U0uYZIB2QRawB85K2/xzN
z1xRTlXS339F2giDzVBXLO4TXs4Ux3QLj+tqks23cRIhNXSswoJERBgfOlfsRcgv29nUj53lzK1Y
Ld36gODYXO0ePuhPB7LLbusd7PRbO61bj2ql2x4bYU+vWL1h6fs5sEUXD6rZUCR5AfiuyfmQtknm
Qbo0o1iJptbpqO65Drr6i9kTaeYVXqCtHJQ/rb8Dq7jH9PHn/CUEqBKIHcRrgKYuQRd6UrRrI8Fb
c4hYWYdwfcQhCLpwv4pdomfqtjtxGPJtAuaQd0SoOOe+ctvfUeLGb8iyKpEeSlS8Q5Myg8x3pJAz
4yTmmmVxPGvuWMVh2Mmrqo4QE+LJSKT9HSk0e4dMit8jrv8AhKhmVO7D9EBLwPCF9c/FT9uME1Qr
kYBAZnLrQjUnjX2l1empRyyUUXxfhZBhpBPvh+cW/cLvOURiHl7onawKJmG3IZFVhzsG7zLBWHKO
+sNqUWqIJPkqp/oYjUd4klvnvqmRiS2qZbGCjicXTsvAJJlqORXOlQ3ssco+IrjXdhC0TDMFUfkv
iq4Z93NhCTMYtg0RJenaX+9V2W2hqaAECL2GHpOeuL4ENxJS5CuMqSg1zM4EDiCoZjAYzKATOWeH
kqxFU6B2Ilgo+eti2Rx+jV+mDHgMctxbHwyImvi/2Wri+pgEQePuTzyioOvrx/THqempZgTQG4r9
8GjVrAcb1akUofiNdmeJFuODxExO+uhRLHQZzMCPgh8Uwony03NAuK9cYeKXc2lEY7kDzwn78+hm
OIlfTZA8ryYYolIzIN/G5kp7oQJpmDc4TNLsMiIAYM5I7WUTGovpUqrObrAlevQMGaDSjHUECSZh
uB0AiO1P48tB0OyUj0Al69+1M3zGvm/774G+Uv7lpeGMnxnU3vQoqMwPbpkZwFrYOXIcr9VixgLr
58H9xqpCvq0PqxKP5gv89N4OLbrP/zYiEv2qfqhIGZKOAfT4nqKfV6HZBiwK9fGylrter9IRS3lk
LH2hG3hNM2/QbY97ImgAj0rIbD8DcgeLSGLhhD0S8c7aXUfqa9kbQ8gd9AEXJvT9tkabg98DIhsk
/ozqldFW7k3NQl87bISBredfd+PkAOawr5IBDOzyogfnTvKS5JayN5Uoa14qPNmIYqkvsmIc/PSp
+zJP1s6cWUBUesXGPISVbRjQu/Yi8NoHGxmHV1Pb4cBui1waHYgdt1rQguKyGdsybiprxtZyHi8N
oSBchHcLx7GEIWwdQtcIHN3rJe9ajMyh1BfVTrDXSezjQaoKUzB/N24Ggk+CnVJo3UqqOUuvThKQ
0KfLDOgpd7TNuian3C477CSQgNm34hRSN7cVKUfM9BG8xXokXMw/Za5jRdE+iJxgPwCE5DvjPc/D
TyOgak23veMExtG5CnrXgo3VCDrSehv2rwUkcKkylcpBU8oFi2iNcVbP+oDn7V+3bjfgHyICpi4Q
1jebxV5MKLr0RCLG/k3RXlBTOdlNRC6H+uCmFU0JNvsbIyXjtfuu+vnSwyszmmW59fnN8Fu7ybpB
dmDl7Zuuicsmra4uI3By1EOPuN2tmsffw2/DNO/DLhi/2PMuhuMBCHMAJGsCoVn5QxULZSz4ptmJ
8zE8tcFKJxCM0bWuc6wQy3+UdL/iHrlCQERQ3UxTEbzSYvVX/rgLEzHU8rnsur+4S7cHkiHcTMRq
5GZ9ov39jq+ezycs7H0XZ+QSi+eOnazfrdha5gve+K7we3sDTj8eMlV3M1gR8E3ROl8uvP411Nop
6W92Mv9XvRkHMoyz/lVuc5bSLsc2c2WB8AN1XJ3NBqpMcQKqOgVjToNd95q79jRSvugXeGW3zO+G
AHJmhmeB0UtnEHeEQrPIXn08jYlzM3rcQFuoCS1z+OAU99gqRLqRIfcmUt/LZdQss+PDAojebEdr
0UbUUuRbdFzOMrxEYaXAe85doRzHuAWQnrZ0WvmM6ySlrlPK0ZzK/psTK/vDLBYq/D+cRcY0wHa7
ervuKECQ7kgmBqOSpTz9kyjcgShVLsDeoEPI15hF8ZlBc32uzBrtP6sQUhkmES3Vwxv/BSNyf0P3
/jCzuHci8YVTNyAo/bCntDcBcbPsTTTFRXW+3/O4P9p1mm92QKThRLwKnF4m5AgCAR6ATIvtfxmh
QZtgYqTcxxEUhrDoO3o4sATDFduisYXbuo6YFHlHYeQaUPBi3g0yFu2t6TYN122NDBk2mJ70G8d/
hGNX2AKpMbrlBekZdSeQEmdOAU+fQLKB5+zr2Wl6KVIKsFbCgK8f5BLfk3WN/MnA5jSg63MIhDQa
XUHxkTw3KfDeFU6BSMw94n4kupchJ/gMDVphsrqcUBggNOisky6AQbgXG1dmbIN9MYQc6S3Q0s/Q
CGzwQ4+PuTHbuqKAR4O7nrL442zjFo4jGgWw2UunDQidTEA3m0GMhClwSdnVUGgUNr5RUlpzx/Ry
x7nhUQgBOGw6rZglIxatKoS82PC2i5Ch/FGlPHLCRVCHvPKMJ8uYcbBcJezC77xFtfldTp3xneU3
TLiSk5aIv8PKff8+uRLnVA2P2uBz/dd3K9Niak/RniABxxBTo67ZjWusL39SG4ZngWRKZE1OUSa6
Oz2D7XF2BnYvWBgb0jceVqsDHaczJ1TLTqomi6XjPtIUZosJr/OTXH750YuDbhE84cI21kjOVMbB
4JTOgYZhvA06k73p3SaSAyn6GQT3Pmakj2diSr+I5Is2kOa40H3Q6bJaf9IBNIrQzZIOllESqrSd
c4rsJ048AEWThL0oCd9zWv4INQrgySNLcDfxmLk11wHDnCLWN+6dtfdJ6oh6itO4j8AFdZEkMhG7
Cf9yx9FAhuFNCmRKKj2Ry1r44N2ryfkczNAZjfuZ3bbvoghfM3ueM7iR+92KgK6fBfKxbg+A9aup
FdEbjm/iXfyHYxwvCzs21cUOxz2eYyEhpIdKwOAjClNQAl8Ws6Wtmv0RqMA47/IxhBSexHUQe8o8
/DXCnBLmuB3JZWPJlWZuz58XVSJB+5zcgnEmNwuER4fFoAjMcs2VO2RUaOsFr84/PgMSIVTM4Mri
by2A68uHgoIPX8FVfJi+VsaaM/k5PvdEzWo3DggvxjA2+hdHzxQr27rY8UZr1sdfVwTnnq7OV7BZ
cC7F163o6yn6SQii/vOBHk2E/kyxe+s2EW51HVvHsT01BwFpyEf7OJzZVy9v9TKdqkoXlT/tFL/g
pFOT/jcqFtm/CoWaUbrxH/sajaOOoYCr/A4hgB0JXGLrQ6SsvoSQXLY5oFgt9nkHVQO5Af/ZQzzW
8sDeIv33DM7Fq7OzPJHTNJmGHhGvNDBaCVPZscp9Cp84Lf2ruwr51IqspQ8WuGEsj3viW4lVgnAb
gmoCCvwkdOwE7+6v8ku3ZPaecgmtMXMiV+axTdagPa5fzy+tATPH7STjZ/IUZPsreN5S07kSpc0z
QDEzxye48yictcgldIgqLDuJnMXmP80P0P2j41bUqbWr5qUv5XW5f8pGc8oJESYNU/ddH9sMzfNo
6dD9US3lR520YkGXKIQHtwRaVz5ABJGEc8p91pLhOX3B8xDf1840O16js9j0wmYZERP6kZlzDdQn
tA6iHnjdstG6SbTqoienNHaX/i1dKeUDiUwoKHR64Guc5QB+hOiJBv3HZASW6MYcZxOLpSQwztzD
0IW/vLP35MyDlnyQ2vdQkeGe6suhJqKvabYTnmfaXnIl7Ygdc+g0jKnqvdC/wJ+YquwCAzZHTX9Z
nBbZVFeEfjXCn3EjTKbY0OyHMNa3QLrwhZdGFpZUH70Z1uErSCr+0Q5SJYlX3rO7uG4MpbSCCkbi
v4Q2LlTi0uc3eDEh+D0MkPQVU5wcnesX5MggbFiO0NPLQfltxCOVm9Gqcu2LU0bNFIBQLtgp+xSU
exI/7J1AjsaTrIRkH7R+84W3FTWxlNC9y/40n5fUwZSO67xtwNRJe7+tpJNJQ1CI4vIQrmhsiNqj
cH2eelrYVW4xggl+QMvMHS3uYKHXZ8+IUdmFO/ixOtAQ8/fi/GaT99VzTb38OJr8Jecf8M2oZXUO
wbQSqmFKRfJ2DNyMsJR+J6p1EXSfe2GxyVOUsIpek2/Iaet6C9Vd+xtwX+8B+C2yPuDop8loCTBg
Za2WfsYpR9ma5AICtrG67wd1hNXmHxeS8eG57NloxLXUlh09vnYRbTc/zss+tIJTxAxF8GBfZAeW
3xQdBoV5wd+wtOQCLn/Ls8FsSjchY3SOukb+2p06Aw8RyTy1/PFKGAcbohOd6s8tSLoRIgrfzXBy
73p8u9HM0Jfbus9ya1cDgdXjF/9o5PdkU+QVXuvmwCAHNReMCwlzhkAlNodR51KX/aKXISVcgNg9
3XwlhEwy6mkUI5g4tWJZkz6TW1IzG+4pYbh3eC8pLMPRLFDe3jI8bP0bX7DoI8jESQqzWz9MmXEp
c+DHQ/tRYJfKp0AmNRtCySfYgOarWORGszR5EgOvGSet6wp7h6eOCChuqMTiHOzVCDV5i0Nd+U6c
xBtS7WXSd3hrnxhxxpwp/LQwE8Cx5TD1giBGR6OwXGS/o5tUMRQe78jQoHGVCTHsXSzvjwiUorSf
1+tZtDcy/xoGQ9c2rT1RsV2wEy/yOhXnPXs5x/wFZtrsI/GnBiYTXDRmzE1uUju5uFLw2HgCp5au
fxwc55ww0Hpghx+gct+a/b2Rl9cwgASuB+UShlvOhwFm6ISYAMxiaIJBw+LHYlQsg+QgYsuwZIlG
/RdGVbS8A6CbCkLFhyO73mYz5cFzDUK/AcLhj81rnRlWHoB7CTsni7AHgK2KVlbjijY4TAnfnu+5
vrttSkq1juEZ9R0x9goD7v7GoLAzFKuOXVyS5sq9QZ+fu26StPPajIZ3u/oNTy4U2rw68HJHA/zl
WuThOQWJVIcyaGDURJbWEkbxRwwPOIRAkldJZWwRQqMU47gmK/gVM93vRTOkZdzOQgf23gYIcdXT
AU6wFUshHFZTQtya8qqd5FGdSvqjLsaAoZLnhKwX2xQRGiIHpORhbuQZ00XgLAQk/iooH4Gt7Lzb
1PTSiewaOvu9I9lldAQn8YRVb6SXidaoaE9ZEOJTJ78FLHCT+U46aMsJtBSadzkTohfeporsZN3a
WcPcpobUhAU7+b70mhN1xAz8tvAm2dl+VplUly47EAcJpJGl3rHYtbOY5aJOuinG74FO1vIF1trb
KYDhKIjf+DcAV/M3CoC/s0C29+mW/W7LVNCxtuPvMN1wg0gcf3rM5ONODuACue4IXoWpkrohuB0P
fgI5pVUqP8IyRb22DBs/ijMInKl8ckMExZ0Fwt45KmlrU4h3SV2Ks1MsKr9H4Ea7UtmGfQtPP+aJ
Bmn1s3zAOXiZ99ByHpSE/WJi2/8M4zEreBx3NLRhbDg8mj3t6UiyrSskgj6NENJFQundkwDh3GRw
uL85em788m5RDPto+0QXNVsM4+7EkpyNg8vQFH8oyl5WpK/RBIaVLyJhu2puYJ/fdisR9g4TJBox
8FngyRd61UMct77Oi+n5Yre5qqTEiAHROe4bzEyH3M+lVS74TyRKvLjdPOlmqEElN9akauDXU99P
5VqPdHQ2x+QZ2qkGfuql/YW2gsio6LOeTQ3Q+id85KHGpMLDcxGjFpU8GFtQdzjuh0qsMHrZvo3e
pynVzjLP0+NCnlmYO6R/W0vkXveuaJDmW4rKaATY9p4dbIozKrmp8naZ71yCxN0geEhBT0/sRQ0b
eld2FjcW31jgLk4njs2kb0u/vVoQrDzDl1GllRh38dyLYQICzix6D2/0mcAVAHb5GpUDGvi44gDC
mQ77zv6G/VcbOVROpZZppuHIMhCDPdeUInocbX8i4K4VgwkVTS4XQDTy9ndvtLhXh4JSuugmGkVb
MqlIiW0w1F6gYpJG3HAeHPpJztnGqq5Gi2o5jy6jYrhlOsNM72rxibgELvwzTyWV/Wzw8jkwWhfn
TmtHR6yQNNNoftniMzG7ovw7eXC+mzCqcnZmEDka44CoOLoypq894TUieozuUNHDbKKMtAuDr/47
FaX9tAUhJy+fn5iyrTrDyqUyYyFq1dylQKToUbPK43J8TOXqhIKvEU4KJF65BelQEMdZVTzhp/HF
+3KSHfokwc449tbIK9wAQWj8G1ivBPSiSFUCJz0JDEeHMG4IpJ0qBtmkTsIcL6aN6wayqKKcqHum
mqy/sWFdMx4RyNtqrpYhExPk2R3BuV01+OUk4McYnnUSQ7sk1WWncCVJJUCAUoDz+JLgwXNiOyO/
A2MOWZw9x9oA3qbRzGZqfFUoKytNPOc7FaAJ3aW+fvQle03CQ3e1LrwRdcSzp9eu62Zvd+G4ndyX
mkp6QiS8V0t13DLBBV2em/9N2miA+W9NBXpGQIs+bc3WHIqgegw2e2dQuhGGoAaleGrJsSYSBFLa
mJuKRlwWHtyoD1tK+XWYvc/oBHRONhKHBeZFZiJ4udL2DS9wUa59d7Gb0EV2YRd19JYk7cdYN/EK
lF/1LKe7RXGb9Nu2DI2a/dRg1vR5KKbe3Rk1yVqAMv1h7Ik24d8IV6+oZvBjy4OzDVgOtO4gXk1a
WcATNrIcW09pp4KWWsdAH7pslVXnQqKF1T8BNsZRKy6jkoB91C+DBoMcerQ/wckyCeY+AMwSWDdH
zK9HFBUJIXUggYQeY8S9qJx8fLPk3h662BUubNBd3R4Y4H8iqvHVM8CxvLYVZD/imZLsgMiA0DsD
YbYUNaVvmegxisyfCd8KJxo+Yy3gNXyfWxkP175BqIzAMJGOHBU7vW9Xxpe/k2KP5yrLV64W99ID
NBNfJSKgBlpXNnBioZlVNNe/8ancz1G1wfDeTuVmyxuY0tVHm6ZQCCticPDWTfd2/ShVOPaJcSgE
jFxpmU57CV3h/yjdizxPzyTFPUJMC0it9g/5U+sSKfnTR4a79r1sRQL8GMN7pigXQcMwo5BBE2W+
i0pLncnnTVD/B0uayV9C8Y+jMZMsGU4SaKSK6geivKmZboM5rMJX8VJQePfzNHVHnByHfFQOAAzk
GVEdeWzOTFopzZXvh3TCz9GCcedIDaeyRhFAwA3/g/WwU9CuaCKUKQXHwS7amyJJi6YRjJuSyn3j
S2mAC5568NwqyUU1ieyL8NmfHYpyUfvzmycjQq5mMr5Lo00fNFVTK1MnKNQ1l5Bqw53139BHDN/L
OpY4Y2YQylYBvWF7NnEgkJJ2rs3j259TBX1M4nFGLQo/Y9earDvp1wx5CtuqwJatAzWJsPnG4/3t
4fojaShm/YtJyegaImNA3bTtY3Jqbb6/sJANG8teY8zlBTNP2NZgOOanatsiSNPAcDECiK37Lsh9
4IJ4FGhHGkyUdBdn9vZo5tkEeL9bTZRmKU/npfpAAPXQotteOI/yHbupTPGpllO5TOmdbTGw2pCn
U7WdoYGs2kAliR+EQf/9Q2lDJkn2u8UVDz1xEOno5MIRKozUEWNyQ6TVglk/oClXzHFDOP/WQSpx
s5SSV/zdAzXHnPT3KCNhEXmHGAYnpbqbs9osqw/WIz5wbbnj7O+7WyCiePCC9qhlZdVpyrdkqx5s
y4XRYhupzrv3vIwtD5oGkFcE1eETYKuGFnt4Wzx+ILLnEN0fY2Xzck0ziIuUd+VQ97V+E9Z1B40l
gwb7jrozfiqnOlO4rl69d4T4dRyTOOOZ+U0GMznoHanZePx2OJfi7fsqjby0xDeRIU+bU1MNiZam
/We9SNfT3HT2m1cwT4Hv4+7BQwJCrY18LLa3e5SXgmXl+MsIRIjkft3OwIWwuI4Q9am9qxXkxI2H
Vgk6kcKQzsvl4hHfsNKlDMsI9roTujdF71qSuyurA1utEpn1q+lPLSntPeMPEZNlSKelk2dPvYkJ
sgAlAsVtevY0/+aonLYYYTt8Catvsq/ptw1QsEKa7ul7PXPgoZtjvfOSttlpJWF1RFCLwnN9oO3C
nJv+6+jh0btEPxb3apEpLhXzRRBJfoAHxfKm2A+IIC0JG7KoWmvMKgx71hHemjlqu6HiwtIylTOD
nXuGEY0wYEvBWa0CtGr7hSxD+eCAGJjxjZhtajdSEaGdbvZJODAB/nmwxnKMvaOLQWDCtyVhIlih
NLsohjQ5SQRSl4VFGAkIvXSwQgCVB+rlIneIy34lGuefy7yfYC7dV+nXGVzj5APqWY5mdVWYPgCl
Bms44D6ubV0OX8we2IKTQY5cdLpgI65KiTCXb2Gi/CA0BV/urFSTpjB+Qkg+fQEOiKuMJ7Cr7T/x
HfbYsMM8GIfNqFtWZlgGM1+ZbhRLvQKQ/i/vWqpxl5i3nlaVCItXPXA05siSIhyZRJ/ghPldXxFB
E6pj1poAmVm/YT4D/5LroKzeNW9HNG8e1w//jIoWKHnRSOILGP0MtxS4z3qQlANXpihbqMd6rxAf
Efy0gkBkqe0BCzr5fzIAn5OY6KANEcCH7H+UYZOAXM9yZURsiBtfbgdVoJcAGuJq2WzYnQnTjMau
+MF3yzABMv5wERDqsEie6iDrY/h7sKUN+JnHBRL4p8pnA16Qu3Fx8M6P7HPT+tFKtgfHD80iXdRa
TzQn+pNII48XAUHb1X8RPSqOwcjlHPik9c7NyUud5TD77EUxSPRDeVwiXXSmU5ClQj/d994lEs88
bg2EX4HRVnIT/VROU+2fTOqlWzfPfY5CYf15w1JNKe19Sx6N8uqUHEMH7twywtF0e1YD4SGGBEdo
xUCZuJpVGEy/FpmiBE0SDueynw+SLRxnrWAKwlvQlCHdXNlAFX/gnslVEN1nbRDdgp4llMTmK2r6
8hgVYuZwZ49VZ1qwCjHASPCXL/BAf6ZY2TLHhB2IaRAwFNic4xv+QDkOK7SKmnc9uuAQZorkk+c9
dyL1qEdWqquMiynr5BpxnQaLYrN4/IRo8up7xptLZKdjnnziQrEkWHxDSp/X7maTA3DOVcP6PEvC
2q+p/MrR8zRY48KxwPvN7T9AROTTfhxdmG8Lv4c6EQIuW1lL6EPkavTcQwPQDVOOYb6lQvNzPw3y
tRJ9FZWdkEh8UdwssPuJc5Qb7jq7rBAKHDrL591NRWDFYBsw0bBcENANsiax6dKvhva7+euMfoE3
4qw0CoOVXqqTcUHPkYruUgZ966l7feqOLTOXp+WaIqlt5bNvJCdv1BbANEPpSh7W3cVhwvrwI4C/
/uVwNZcO2u9PgKdm1kUZfHF52AkvBWTdVr28JMziLRoAU0FO1aQfGYwrsCBonP3Bdb4Av4+SsDp2
KuiT1vwqQSx/aIL0as9KmAkwDSBQKnqW+59Y+fSQ57MX+Qjl+X2Xgnh8TiC3mh5hyKq5zQV/50yx
0/a0OEJyoAnU4YaSTfkr74s5KzGWkqzo64o3Gpb+RzUVq7s6+uthlGCB1qVvde1cKyIjgSIwnain
vr4gcMP+O/G+1EFfvHOY7rDLiVwgDJZrC2oS/GrFHHQ4oVAkUDkyMG/Vl4pK0t7a46UVAMVSiDs3
Wpxavajkns2erZd3VH9HDNIj4xGgpb/6w6HqZm0KozI8mvMXav8oi1NfhK10Cbo9YEokJY9oLUzv
wTlw1GnMTlF1Djf0flNhTgVddaupPqs3p9g5a7qs2TSCXmhJtkbM7Ufv/uvcpIf1BgUgRVtGGOp+
AkQWMpTJUJRExaUVMBZbemozpt8jp6gFzrfcqpDU7OnIhpiGi/sHl7hjm5MldW6LswyREWh2DFpP
VYWC+ha3ZfVgUkLVWhospjBnPPPr+WbNwcXhTHMMh+L3/g3LaxsYgbLzxh+VR055NezjcGuoAULE
JpoXuhtkK0rtBPDwNFPttQSXPIzcn7F87dzyxUjGaQEO+wII5Xb6oz5Ty7MLfG45FQwhFYOsCAH6
ZnhdT8HiHocNJYR09p1ETimGlvVf3sTglBVTZICm1LAhfUJZqSNquysudf0s7/EIMDLFhgddvRit
NbfuSj4MPIyr3XZLINvtJWIw7GJUooHH7+m4z35DhyXBE2YMhMuevtqE/EGT27ExvoYDnDcFoY5K
Nzujee7lB7pv9UXS+6MHphBxjKlKYkNYe0kMgxRoRFQ72fB/eOkvbi+g4giri+jBAdeo1SauuczM
i0inyH0N4JTb+ddKd06X4zdLXRrpQmAPacPjKpopk4lBZU+hcEJDrOLPTikjkQew1pWAl1/gzjbA
6JHGI+RRyHlm5/zh71Kc+FpEcz0/nvqw6n9mj9d8jV1G+/eTDTtFwdp6G+xMsflODKxid9IeS4AE
VIiLE/vfKJBz6GglbiFK6RryTtf382+8YHAszSsnIv4f8KLxsLYVZcEHoZ3E6C9/yK/VlxId3eQS
DSxqyxRC6i0C6UEK2Fy9TvoG4sHw4GlwTqOJher4owbQH3Bw72ZPCC/2LzCIpE8Ii/BdCGbYeCH2
63U6XiGKQ3roN5VvJZPUIZDXaDpVyF7HppBWzTvSvH1F8y6k11WFksK+rdC6wMryLppBgsD8moVC
NyXMeSEb6yajcmIiTaflyLoREjgbFvoVPCZ5Q6GUlvEPh7oIWGkTZ+986iQM6IPrHIVupgr8e992
2MbjuF1hfhC4/a0pcUfuBIBFCl6UE8HAPF6LubiembwqPcSYpDPu2YGApr7LN3DemN7z06w0gY4Y
iHeAicoldvDKzVSrlp5mScjrO9DR3aSeeNXU9p/sgJThnNC2p6TCXWOOxrRTWTT+zu2WuUzIFFE+
QYdZTrFwE8KEHZC1GTwtlhThyxAfYo/udR0+Ryn2PmNBGGB2gDen5hollR5IDJEllqrarqa+21Bu
VXNY9M6+gN0DzhYkemo0W/hpVTDVrxrLTmK5LmJYfcQjHnCxcIAxcWcV3YP1l4q/WLMgyrE2C4M+
3oxBq6hlCUcHFcxTgZt4PU6P57SAeInuzgv2kgZreUkJlRmXs6Y1Ur7jAo4KOP/6u/O6ykHSE4nf
kXDUa+xAXHE5B5gfqJ4z2g9Uct+RjgIOjAGhJQetE2lsB2IGB+uqYHFLwcPPde/Hx0yzQBnSBjnF
HtIf4IAwrsJd5N0K7ytFVNrWnIB4QF6L6lUGa6V0YDJKGqKPrxqbiN9JfTZSToIDGMvUr3TBN8ys
cdKW5PKYos0cCktEkEzn71b9FCN8USOzlSnfcZNMCrQQxzVO+pQoNqqxCnu+R/16961+rkL+ra65
eQdMaeYavAwYqGJAWWoop9JDn8QJZ2KBjNRyfkQxjTEblZyyofgb3PJCQ63BCJUwobTLYaFzWQpS
e8QXKtCozK1ef5FCOYC4fE5Lr1X8U6kaonUPE6ESMzd5XlUtMOsToZPw1YE9+r9T9MLq9joruxRE
J+u+ST0vEpTRsZB+ZZaQxH1VqZA5+5qF12SqLsBT/0dKsgE0ipJfi/P6s5SQLQrqWcY/nsPQkxjQ
so2wJvfSDqAPpbrB1d9XT3WkzsXdi/QoLp0MLFzZchBsRNn6ECqQjaBa87MVqvGPme9sZhNYuVxl
qQexaY7kNE2TKSFOggRoArQpNJ6rXJGX5rlPwxWGZjmdCnUIPGef5garUFbizTDV1Hg80Np8g4Pz
s82/W20OnnMGMIrobAbCsHKSTeiIf9asGT8eq0i4aMpJMzIPR7TnrjtsnVXEN9UfDRqMdNBT/Cke
gEdxV0MVb6j6JEdss88l2tVqf+dogj/HmkJiDVq9xUAw3N6X8S7Ixwagh1C24jesgVsp+pEpFkwd
2dDLKENFQICWvSJrQgstqNAy5zQxfuGSafEQzN5SHxvjdf4G2YFS5/4ixi3oiaRiwZh+7c17IGHc
zXYufvu4VpGZayWk31cznQCzK127x1pPcWbILnRWMOLPhh/heBpgr3SUNrASt8VjVULp+UEBMFe5
BjgOonAG7T/VqEeUYnsW/io2e4HxA00tD5Jk5MiLUF2zJ/XzffyVpqkGY5GqoJCNJoWAIs4MflO+
pQ+toO9mBiQmTcKAhIicQ64gxkDJlH6HGy0BoZnel+VZpQNi7GHz/KstF60t9y2jZS65wgPe5FE2
QzeBsjCZoqqhzF6al2cYJ3i4fNGi5s+lGzKXlNIyxy+VnkILl6ONG0h9SmdsX9zbVIzfhMgASAw5
qiRvipDW7L6pus9/ktyFB8J5djG2p+FZ4r5Yt033+SgXqhZJwL23I5wa7EG5PV8RsucZoXcBx7Fc
6RBni6+bB48LlRwWNe4XYI9dJD9mdTz8Jq+3NBwOroLUezaEmcsywyvaj+yOg088OcSeLIHAwwci
h9svQehreQn108IgdNRAjjd1V2D2t3qcEbDRG+iXes+pe8E/LHx1peffUHtJToARLhU5TD+ghpya
7htaVsQu2mZZh/V+P9ZO2GGiro2gpZ5dyJyixG0RGKOmOfhOUUa7IwYI7XTO8LAFhvfp9eeedzUN
jOCKbAZ2mpmkDjOrxxqHsnxVg1mNSY5Tpfl3D4C+S+eLDjPJseG+qTOt/w4zW2Xe+AlQG1WdwUCA
0svO+l5NY9zvhYW0F254z+tBBFnpXBgEEAaLaQqlbbTHGm7VdlXFqZY2qRHQYoVBqUG0nqcSunv+
Hx8hdpCM+NvIrYM2rAXWy7zMwqzpcJxlsORhU1Pw6O7lC763+qtOAyCSi2EsPjaVVrfMzuX5Neov
SYZ+kouLvyiPujnFsDguLfdsuuVqxhP1WMeHCzTev2T1X0Z78ggTPX/BPhsSmUM1zOIczFquEkM0
lL9HA3jUMLKZvugbUUBBD45NzLPlkoaBe0CAqlNklb41uH861YikrzMfe6gyHYXYl7I7r2JJwonf
zWeYvsEyLA2eaIRPN82BUz44CWs1d/DAgyGFsFyPr6U17TP7USNrjUkZxVhCqjws/jyAGovnyLRw
mHDEOPvtUXxzQdTUT3CUKKtJjUgaH0jk+RxR5UrevqsUoAThJ/3NgwBNmZJKNkggabdKwBBbHFnk
D8ZnPdtxhUzbQVhn1s+R5YAfTif+FUR38KubKu2zBf6N91N60VvvCDXKXdktBvIqoZFjGr/AeXmA
UqfJ2o6HUaelktw5Qi9/rGFUKX4sPttA/pJgHqCg4dY4CwVQ8Zlrigi5fByy+bZOxhw9tYj7Kk/u
i4CAyYJ4PzOKt7G2kJdtqt3qSVedXpNp2IDFNUDTStTy34R91qdFhsKhTRo4llHod+gmKUuH04Az
5wB3QdMa0aycMCnXkXsrsDGgnrg8CsLlT/UHbV3nhF1KeYBunjvmcAqBE5pBZM50nt6PiBwIrmbT
aIB59441ZIAUnTETUpDF1gk/nB8MUXLXlnr4XKWBZj4w3bdkFpmFBpkZq/m+GQMxOrzQjB2qrBdc
J1RXfa+d40Tj1QrS9BzgiN82DHrRGXxxXs9ZHS+p1w81Tays+eoZeZJ803nczjBriJSGb0x6mzQS
2JX0q1MknwX2p7AwRnUrLeIYk8iYdEpSLpivMQjKAwFrEUbxITQ23h6vEM1Nd8xaTT6K6BiKOHlm
ikXkIp66PwWbP8zBjFYRfhzCa7BNdEQvf7iEKrgRrPPtEoMUMCRcr8OcMTSvQF1xcVqDxGqS1Ncr
s6460N29a6MP9nDNRZaquZ3JjaPUP6zeldgwS40YfozYgO/2umE7/5Kbk1eYSUP2bE5NtowJyQS5
+XZ2TpVYQvxBW2nMD2atDPjfW1Lac0IOOoky9C5QJf8Pf57rTDBfm1y7zIhrIVC5nynvZzHmseyX
S/h37zhrClA9jXuHfFqeC1YT39fYrFBVF7LpqfdTIlquKwAvItrG2MzQCFBG/fRO4M5Yy631Wjem
4mqlkyEbbko3xLXK8y5iNdrUqTwnw7aoBhYAnkjYjNuvmbU5JusRxfZKnQk0YSrFUK71Ma2mgTSi
ZL4AY9ptI8eSR07UfDf7FdmFKuz7TZgKe7YV514Bt3x7+WCDjb8zHmDd3dTkTq0CItTizz3Bxihs
NC//+IwqnxgTqnlcce7FLbQ6OW+5wLn0cfcnnXbtkQzUm0wJdB1V5YfVr/QXUKDT75esTPgkUL4J
aIitZGuH52moG0t7HHji3BOkxFj4WWBI4PlNVTOzcFNZy0KccPfDwrxtUXJsTleuYvlNBYwedcDI
caX2FuM8quMur4W7rfsPGhnticH8qUNz82+Q04YhKSRUJLzZU9WPJIcGG4EvbxrEsv/MCf42oWx/
XED5FwDysEVEll0M3NZXVyh0EsveAVkSRgCYdyu75FFOOPn59NygyHolxz0Lr/UsiYiRcRKs/68m
oP7CGyWPXtMOHctBKcs5I6hbk0T/zGuAbBPMNXUgTsqhMJL9QeY7pkJkA/yDHE1E7mOlWSd2I9HR
ep+9g946dJqWT+/6jzS5HyS4qM7r2qDGDbLoyVDvnvoA/CZN1PhJ4M0039D5TaVcQUviPLRQzeUj
5coTpfCUgiNYMMU+cWb0nhw9OQdVSxkC9B/zs82s5kvGttsFDOIYvpn/i4wHkG/V4jOObeIRYyke
TPiJURMaccbAFvgLuz4x64TB24IjJ51B96qKSMo+nJwIJkdzEtbaeQFlXW4io90wgsCX+2ayiG4e
7w9odqsBF/IXmmM3EjpmgYqEq7pM74hMJ/6xtP3MZkisBHpJgX6SCZFCLPKnupElQivt6Iiz/b2g
mGcgRNu/cTfgMAnK3xmlA+9jxMmYpY7LI5yqtsWUMPXvZWk+L2rgL7OaAzasgpDKhKUWR9ivdTXg
Ia0GHjplT7JBmYy6KOdYaQRgR/OdTmLcyLNYU5d12sAlPb1yiE7Ra0ofMVAlieiK3Y5KMNH0FUfm
tJeTfugAuTP5tJenXw2fF5nFfsxu1BHv0IFdzUZB17K4DgIfQ0uTyipgi16CkHsqvyBRaZNu+ZDD
/TV1icvl50tdu2vAEZOmIuSLRvB/0bWwkmEBuztCMStOGhe8bItpveFPhhNBKc1+qYS5eFu5+RZS
wJDTut+mqiZ0f+iRFG0Mc0IiQalWzFeGK3+TFEG0UvstjOlR1BqbD+nfxMd9c8uXQvliugspsu7Y
RYYkp3/TOfKwW1OSUz0xJyrHtEwoMfjs/O4kV4Jhr4N0TrJe78ZVBkbWq7NWGeG1jBU5jbBRThu8
phJHH9MclZeKeWokhXdrVXy+Qwwzx3lB1tc/QnB0/b9FcWmy6vboiyEj34TuaaoSL6cUXaUgwOct
vuZFI1OEwJUVOWU4rd9J7hsv1XfkkT4mRnRzsRYS5Gg6wHo/XUhBOPoTMuAHzeaxbXzhhFF5yqcX
ydG44f3dz+uoVFc1nnMdjpKA4BJSo/icMEJoQ598F9pMmId8XajEs1fMNGvTc0TBKD0PNdQ1GIhS
Nl85Wz/mFV+I74fq4d1n0eJVMzMoNENnwovAuQrOvAOE70QqWzq5stifCr0TLJMF/zta34SdxnOx
ZZUM+DdhIcuH/pJ4h4dot8IYNCu2aNA16ri/QY1OpXsdVO10ok7TH1U7N7ZBjKJXN+9AJYRKy+Oo
oWTuqXnxT5yr8oI1ihswMkqmOlqItWBbhRG5XqD/M+5lbIzIkAQnYlHgTYA4hpIXr5pP4RLwG8xs
lEitBP52AB7w220htUm0ijcMf6qbKOhRC8zXWDHk7LEc1ouloqY+jUV/w5Tj8ZOnuZaBQTCZDfZY
o79Y1FoJ8/3hawm2bew2d2AhfkIF8LVfi0J5LSaRign4FWoZZ9eEz1DXhF65/LuV7RvXgjF8Wwp6
Eak0paKqwsFLZcIViLpmtpc6st3pSgClt7wn0wedrYLE+xaUkVlnpXibIleIN1DJ+NEKjKv+Uz12
8BfNWceWjRiLBc52wUltkGNthxPAeJby5iIHRdz4a9vH1e+JWBeBnmphlWDUBUdz2OAlp0fr2EkP
YNjCbp57BinzObfpJIHt+lyvyho1cqDxO5Pb2rqgyY0lezxhvefa1AuAxzXike8du7DyPmlkkHN2
B6BTJLQo+7qrkGR255JFImn1rjBXNYnH3JQdlcYrJBHx8VX3gOw7+n2B8tl3bO8CQ1WVUKZvcfrL
fPq8g0vRR2UCfGi1UZGhMt2uS1Ru8+u0bGhGdpuAs3jXpx8Tj9W51V7cyx/kaaCTGLpFGb/nHiC/
EeoxtL5hG+LaZiVR2zps630wvS2o9UojFjoG+sEDLiU6S+UFWEdxRaBkRotIZnEGtWaTz26xDKnx
GrxT9EeLTu3w8o6IHe9s5CXTB/4+/an0JaObQmeFo8bScamlLqKAKMyBZbbuRfu6wDzmaKwsDL0k
s7bvoYAmPW0O160kNN0UMtejIhxGfy6oH25y98Wzu7DcpoWy1+tuUVY55cRLPlUTGZfVWacN+cqa
Wi8SVrXDoVwVnYY+xc1dZ7XvXx15bqvXASHowvxmRAUBCtxzoKunN71a7Q0TkPBO71DOnJ/o7R7f
d8YUA2J0Ak/zGEOHgymszWGOx/FgCL403JwWMjpizoWjlRZcFgkCL58PohvlGR4cx9CQxDquJ9AW
76l+8RKRSvb5iDIdfofmbQ9ZcK2EVDZnRUXz2vtxPkUSLIqeIK41HEKqn5i76QREdVAzX5Bg/eqd
9PAdFoCeZ00E9TX62BEHOs5l20CUrMffsZb1O+68XKwO1DHZDRyhhynI+BrqSXPr/aGKzwOpQfTI
agEZ298zMChK8Ae6waBeaUqkr0GnJmUlndAmoD4E532MpnncFtKRT6ygLLjhWnvOQ81MAtIaQUqu
pnDSP2ne6ofPxoat5pbJ7KevLfPPgBQNQgJesPATVy1DMMTrFqNlDYpw+7eKcdMVzQcSh7oJFbLJ
ErLv8wH0ktp1p7Elr/zy6rmka5fqDnT4wEvsNk/33JBQ+RfQpekBr72efMF2HDhxcScnGEy+BYAU
IZ0x3Ol1sDy95fMLZkfgvVNCbP2erJ9lqthOSdcYJcfTfKcF2rrhoyGqsI5DprsNyv9x4fnpu3l4
RQvi2OyYd/k/x1rycJq4uAcwqv4xWHux/+YZF2AKnyFkbNqJ3eht9v9jYjr5Rg4ctfYeozPIk9R+
z9CJ8W6AQ8OxZEj6/tAA7fG2xlbe9Ae/d5qcQGjAI5Xh08aELrH1e4FFOSsKqAzWamtdm6tmz6PR
/pWgfLljNbVXO+S0Xie3Q0mY/HXazOuWuTTZxCDCvbfZRCLqmE251/bVNZLmTFqlVQqkTjjGg4/4
106uHtJqf4P2ag4JkdhXsBPyDsaSsBt2HKKFhIfLbXRGZARoZuF/MAsY4Ryrez/rqMmvfnT2T1Zg
kUbcsUg0k7mDInzPR+MgMspV15gOs0ZcM/3Xixsrk4GfaeB1iEJgFo/OJJOYSeAej3Q/5OCE7uoH
gOcKyedQ9okMZC32JouwYkF6ljlh3/o1Ml8bkWmpwrg+gpasKLxDz/y3CZ/K/DviTU2KwX63u49G
107b0f5nBLeecisqQsstOZOUXiYoKN+LFJcODdKsx+4UqKsYbv0GUOBeQKFyIqK+DbC+H0Gb0fCM
8EXPglslojpthwe3PRbDfoiFkT2zZ7Mi73BKlEHt2lQdMy/SgbN0l5olAuNlpGrkIYyieaBZN8FC
qSwECBO4ZR22CRAQAzU625k8oU6YhCtNTwnSGjXvH56cl/SURf7+rwEPS1om5uzMo1GIr+lRxGAv
hGdrzxG8rDjo7K4WvmLnN9yhVqmI7PUtzjcmAUsJpSSmj92MZ5y3frKrUASzqIX6dVWxCJ9KqD0A
X41BHEsNv0TxeMWooPWgQTSkSbIVWnix8/6gjX0pTXDOnDQZktaSKUoEnD7vcICoWLdpBbLHZsgF
47ntnguviq1CYurYJ7C83PzsG3FRQEkpLPDmFRziBIDJgT6Xgp9mQb/rZK0iVOwLz5iZgG0o8O2C
26ELV3+sMWZbHy6h07byjV5FGxr2Oy19d2SN8nNCcVeLfOl9AE0sxHcek3VI36K3Mxn4gM0feRzv
TjXDd5og58i2w68GrVd3lh9+QwGMkYMvRfKcRrMnhpg6Xhas/Eq3jgt1PBpXgM48+imZDP2QLCin
FM933WfP9bpNKfbSDwfZd7wiDqa1JOxnwR337MYi5t87KXHzTxHmDNhFPhXPaXSP1KzEuiB2Tb1a
xFjS6isLlQPZoJ7qbfY/WXhsyfhP0JDZvlgNSM+18eX+j0gcL8IFS1HD1HU8vwRiodmFFT2bOx/G
jw5B7ts8f/2/Dt52FZAbvwb+i9HB8XV89nIKCUc0cqM5Hn3Lub9mziscwqoRQl5jUJxAS6csB2hk
Af9Hsngr3DFLp3mbzVidWA86GSVDl4BMqf0Ns0rfJbbQpm63AC/qy/mEfYVO1aeVS3uUHHJ1P5jV
mMsPyJILE72miDnW0TY0RWtRWTLD7RzihsuEECnDSI+7DRzGKEG7vSsHX3lX8x4lv9ytKmXSdRaa
bUvsld+P+zkQ7KTN7xy3mxvEb4s9Yp/+0I472w6J2kmESMtvvMG725JlKGu1vFPBcNJd5mFm7fCY
Ysns28DdxeiX83E+mEVL6PDEXgfo1B0xlaJJcR8t8Ge91Xx3x3LhUsyArmxUAhiJaP+V241tW82U
zn6TPBB0W+IESI4DeyFHqDPcvql8ppSF5E68guFb+eVlp5wNhrrQi4Es4VUGw3hQsrcPg+smPK83
lvGmx1zNz5GMcqRHTCIaO7x1bbLx3v1D5Gw11DI/AuDyodLpMk1rOl5YhRnXPh+pWcLFVgs0iTPP
T7MNNwmdBSPb3TGedCJ0mAsfQWFVGkn1zl05R+0Co+u/STEahb2qDEw2kgBLGGnC8iyr4rQWLogO
zyixOTWXIDxUvo9oWAySRb7KgTbamqU11DoA0vOtcyIXk8HiOv6EjrwhhIlS9IYHK6SOJh2TEjIR
aEV5xH3v/WKbNad1Vnz1HiD6za21zyqYLSDq733RCyC3tqvUuhNEpgnj67xtuUL8a8CjZvobVPGq
3IGxK4IdswPmnlUeugwbhfvfMtuJKb3iES/PMLrZ+jN+rzslZ/MZPsfkDlEO4GiydZXR2KPBzg5a
DuE/8qUkmbKdurQAhRTkOIxPy+EJOq4Kt1whpbvVnmBkUnjd0OKr1XDVuewdjsPXyp/wu8F/Deb0
ONkLDUbmhfLnGbABZYefpjv3b6c2IFprQ8DxGNchQuFoclvKDaXs1G6bkRTKpVOl/zziHemBIzTV
O/1yYodJnP6ET3O5JUzLWEMRYlbcaHv9AINnMz2UXRbq/NsGY/c1rJ5+httbxpwHGOd2/pBaAYfj
y2arK2uhC1bFx4DdD4mGtNiFFR+nXHvISI/ZmQP+hzbkdzb5hIKqXTx95tpzbAMKozWJbohwiCED
I7EFasFKToF6q6kN+xZ4CqsPRxK7e2wk23YSSxQ2BS70Y7oJEjM+SXW8Sa5C4w3QxYYhr4a9Yowx
mZz1D6aAl5Fx8xwCMLfarmaPqFrxIMjVhptwiLHDJgL0jtn7hO7PU42pIZ0J5hHFmNxaGSfnWw3g
+QaFjbWwPSRa9pxU6G1C8F4zIXzYYU54S3ZGMpBrXI+UDZUPFRAWMbQv2FvnaFlp3AL9fiQk5MJ2
qRgPmPtxShG+WiwUliN+t5fmqy6ne5GNu9v66EsF/LD0BTZJkhi0pqiFeUE3ofcPtKAAc/cfOf36
RwJ+L+VEHSa+EwPOs/nE+BDohKbJrQ+7pbS/P7y2V6Rt+FGzGuRieTmR91l9Rk5nXBiXfKQNQBxg
ebqnZcjMSZdhxbo4vcm/aEC126X5kKg224AErGtvjhG2xi9IAWyOhc6mUhHiGCap3vSCX3Pau45G
JJdoHGjiXo96fbkxPRrEO490wx0U6wAvGErbxw4vMnIRPX57vK4idiulu2PpNhMrN45npr+SBWtl
upc/gIZ7ZDCjC1j/7mh3tt7FOjwJkumX+qiN5GLn24kvAI+sR6GwdvjL90VBQ/sDPo0fmmmwbbiC
ofJrwMHA1CYm1xYxOCqiuNPZFgrz6etlifHTDn9zwgpsRkVmAgHoX7ySpj10aKDHo/cmQxEx1JN7
K/16gjDup1FoL6d5wmV+HfwZv/gCmKmJD9QIrzR9GkYN7yN9CqFk6dXIgswdF3oNyHhl3IevF98b
Y3yjTgZAGxbEqd8MgFtWl1/OL9kAMtDooTwCT1lEcUdv2un3Z3tpnuCKXgU7xehoNcmhLoVaxbwy
jPlQABEKac4NSI1gDmTCChlrcNFRsV2zaXnlBd2CZE4AZpKpVtoDYl2YTLNwhF0CTNs9jOHftYaN
ABnXFLmwRvqkt0IphDVGjPEmKHmBFlgL9dNzqfGt9md4Uz0Hm5M74TVBA8Xl0+0YXwanLLYqV8+b
50m2ZQywmQFGulacbfm9BNoknl1c7wun+Bjq5T5epGvtaNsHETVyoxo1BRGDyFkeiF+CgJ4GGXjR
xb51KQ73+0+cksUavLsU5YHU7sudvKCQ6B72H3fNHAGDc/e1DNhouqGhACtXClSLnjIJXpaZhFI7
Mw2IM1dLqZ++ma9MdgyiCWH1CHb84WERP33iCd52n8SEW+FBELoUhPy6AIFWXyZ0YemJTC+IBrj3
mMLaIouZrzrFQZtgydnvtQyJmKkhCnHLCVTdMW2ufNwMv2gyJdX6Tbjt9/BzZD6P9qYS57uznKzn
JL/QISI2XG1Sj4QJCuk3TmFeb8TSsWQ/6/NxZNxyH+dXp25MmF/gAhLktt3Die4OCNn0rSnO2hRW
X9dcszlcYWjLoQncAouFQ9eZpUQ5lzBccDYVNBmPFk7edA6ipgBiU3Km6D44HmOLksS2tc76Pon2
/HA+UU701xmntG71FhdG+hDk/VnYD+3XB3Q/XKjgb2kekg/XNjFkvT8oh1MpK5wZIBVBL/GUOHsF
VDGKsw4RsU4wgACTDLhTpazaaYTvNZqP+Ije5sfA02vpPIHneVC3dZArF/ZA98f1tsosIGOXLmXq
DKlbkB6zaaWcfX81F5J9eHXJRPr2adlK3vIPxwvTLVP/RKcCSmJo1C59UduIIopgal8DMYSffXr4
WJ6ox1Ai0nSY3fylNrj/YbEBxSDI+uAir8gSiI9h/3b62wPz995t1vq6Jjs9/UzTxXS60eAGL7oa
nLxzZOuxDdJt+4WdultlzpBibAMye7EhOLnIcuu5Udjazf6gQM/fPK+iojf4hv1+TQJ4LCeXrqS7
z4VfCw04VwNt9TktXDHuI7M+zG+DGfGEj/5Y8YP3tV08AytwKLV6YFWtQD1nS8P0bYUkLO5tVlKe
YXhtgIu2R0sThKRSwCv18SN335dozfommtDDyqY+HvGDxk6O25kZM+Vp55fYEtMJwzsiqYODUVaY
qfpFNu+lzgGYzCeT9mH1BAm7PAdIFoJJt5Up9hqRFnycV9h7a9l6eQ3oqUEUJ7TIn9k4V2qoCrJK
Poau+jaf9/+ha/wGS2R/ALm9bWEA2eS+fMZokJlAykX7aS6RR/Riq7MVsQQN1FPhdcCZsgFS/HkN
fVMY9iCz4pvQS1E4YeXXZTcaocw/LEFNPlZaVXPQuu/Xp13lrOStyW4BRwuLIU8oz/XoMwjv+dgO
g4LcfZCaqg1/u+MhajnvV9YR260rw+TDWI3ipWgqV9lLk6Y8DcXsDjGXzHEewoqBzJECkG1bam2h
cql599sQPHnKt2BQbEhkppL1EqzOjNsctvpjmH1Q8AsvSt+wqyxn691JRiGcQw/JmSRgZtDTxUk2
93VCYv2caRqGYNAhiKp5km3GLWVKnFktHkLTTmvpQSTBh0LGyYwCL1Pz+5wBKQnIdYo4ZUSIEa6k
vlSw58uCv0pBKeio3zGCd9ovIUe0TACFoo15rN1fuLnKOmm1VxUDgMgfvfrg4Lt/a+wb25wyA+Q1
p31xAOxWcj5MRe8MXXeERyXzlFd3rv3qA2OzBeZrYNaem/687JyWhRCDQvH5euxkgP95T392ZGPY
ycs9MeFY8jtw0dIgyFL8JlDa9bc2poaM3vYy8SiJywIbP9rLnEUFyLx63bbDJUr0maVFZ0grBzEm
9xY4EKcbcgEPPY8qKxUAc2ctvj9JhHC9Sj/DHFWCVn1n/bG0jx32LRmEpNqdN+ycYmEQ1Rl0plpA
PW1+5C4cICTDcL9DTlUDmjdY1P3vsNaEPo9h/mfoHUuYBt/xHF/5kil4pAto4fC98f6/SAW+jgv1
+Ye1hI8feIO9wgPBXHVLGype8GbN1yVWM+yS0TMO+NlIyahMhoOWodqE95fTsyeql/S2nKnItlgt
/1u0BbxQFFA5qO58nsnW/pT9GrQD9xf4Kh3PmEe7OrueZkDClaRWmOUiGBbRfzSU6WWT8Zo076Db
oR4Z8gjAetBP5GPbtoOCHPG9kc++DJA2/g5tu0Gv2vUw03DG9pnfUSR9Igki/ww0oSyy4Hl1D8dd
IGsvJ4GPSsCdIKrAVw9RIiPa60A6Bo+N2pv8os+mJVMa/MQPPS2HsdboCaSGxhy3ahpiDWJfN2yA
3oxRgPOTpPv1yd7j6+P6QAahFpR4W7yTOjMdazIO/VFclb5Gtg/dV1mtSh4vvvZzTGkF4Z+XDiJx
llEhT3TX/M+k4s3RsaUgOwBJ/s6PspO3IEoYpvJl+O6SnQoI8XB2GKcJAovc73umk6BZWw9xqxWI
Bp3AOOZa5XsG2ESr6+iD1oARUDSGF/PV9Xg/6qPbJi9dvyz/UrMjdAAO1FAGoELQdrEJ9CvvubEd
Ex7Srvu9VKhG2LhWzC6t9ywEEyaMstLeh32+aR3l6aRuZFxUuUDDf98FYMMNJ4Yd2NWUkwKhr/rU
HT7ZQFjzTA8qKe0r2ip1nw5bmEa+frbMA1CD4/L3RHKY8THsf/+houEvSP9WElJp23HARGzhhYWh
Ii9VK1OM7HoBqG2xRpnK9GsshkUdhgxZYZ/algkXY68AUMxxYA1uFfk2G5BMf796Oz1DPZORs0SU
neBls9wdy3EOyBxhHfbbdKJf4hXCjnmgBetxj2F88gs7DNtecRn44gXadTi8g9DPra7x4kz8BLRl
WTAWxH5zhJKGFmLUV7HhLO6+6KwseP5MpNYNyYoDYmmAjoonvvk51nDCLh/+UzxK7JVa1g9BDLOb
dCeRgHxDCm2IoJ6JuaTUgCSfPFMqtRMk+5t9Q1piLj9CcIm6I+djazvbvsERPeTvn29CHVg3A2Tm
HOKU7XvUgd4nofEgzeuID8rFUwUFUWicPHHQZ22EOVIOyn1cVFwgy063ReVjFYw5sXjEBBgCVvn5
q99+PGmRRYJmmb1+fd9hfmjT0THFPux2h/JCAgXa1wFbrnJnJdFev9x0P8D6X2P1p6HcT9meWHyp
303sPnRFG7f4miIWAhMZdNjikOjMEkWJxQCh2utfcRQf9Maydz6nTh6Jb949iP2StC0QSs3AUMd8
n7UIACqm7fu1rt6k1AiMWSafYX4Uij5+E1+cydEIIXbP/oHWm1j5yvAyXn1rKgdzz82qV++Oc7b+
jNLn/RxDB6eHyNsOG4wpi2FMefDSK5FEVLubuna9W96F+JwweRzMlpyk2g4oPkG28OvlcHSaIiXq
8USnfrrWAJ2LMtfI+mVB4sVkLDRdatAreJVaaIeRfpa+NmICJfcrhv47a7tHnztFYeR5hkgcvjAa
PdjFtuXTI3GrJkkd3+P2sVcvgfQDusS7NKxrhXjh9zYoArUuv5+xd7Vtc2zF0l/Fb5q0Hob1D3do
hsaC8YLsWlxS2QJ0lt62Ca+N1nUyiZBv/vsCly10N4lBn4AWnkJiBaBATAJNGZhySpD8rowEZNro
b9ImWMsGyb/oHO8ErhLxVwB/Oy0wFCBgYddU+m1lDtFKb5stwG+QPhUosC5tbD+416xgSrdQWfmj
uElnGziIL7m6QFbg4CarUS9+efoTK/lkSaj+HnMBx/wFk+De4dUd1ec+k7LRU4FXfFP9gNs8ma/Y
YGt4Vzo/GRosGjSgqUk3LRE2EnVDgIXA1wjdPSaq85bkbCanRZu3jK6uc7dNab8bJOTwPtdcOUmr
uXyd0SjaPGgjNMG2KuI8MI+3hESa7mys9CEwUH8PdOYVZyCQ4S+MgzHWB2fTkgPKc9KHcQrlUVYa
K+xFhcvHoh/U+OUh/3U6UB+3LjvdmIfe3/EHF8VHxASZqzM5OjeKo5JB3Xf2voKMbRX1cpRNmH0p
9urqW/KExjjipqG0P/LANFtJ5BJFFFuPMHqQDo6xAUK+KKpBUh7loem0zCql+Za22iJayNO9wY8U
thi5aLYl5qJTHBJpwJtGUIcKlYdR8C5UXSzxQc68nDbWhLgicL34vas2fYukR1pGBH8souToDqBU
84rihYI6CsON5OW7yJkPudg7F9DAixx14u1HuGEDc5nhAA+volgXIq89qVXB49Bk4yr2sWzP1V5Q
kQNpbgiGhTVOmDMceKb9vkhhhJVYwh6bbWgMJD2SDPUwYh437Q/xrH016VMIXSXyS+YNBE3zpiiU
/cglQ7ez/6t6scittWx2slHHPFj/QHfarqZSrrcsUDtS4hcXNr5r73ZIi85w9wXRHYH1qB4QkClH
9rsW/K904Urh/wGCtc2I4sD5tkNuQJA8kprBl6T0g/jElgvzLjOj+gl4tR3qoDcBypiO/kh7/d5V
z25lc/Eze6gu/3NwKRur63pRQspiRr2Pr7uaFBwF6ICskbvnbf7eW9xeIURiu/XAe3LcPhQgU+LA
QDHgmnUOLEctMgcWj53CIHa6BN1mDTJHoF/YxEUBb9uur9Fvqau+ZKG9idM1lJJMwj2ZD62jUrAL
up4nyekiZVpG9Z1/ZoGhvGaRwAAuMNfSDlmuCIDPahHNz8NuBK60BGUiT+Pc84GGEjMiPxWoZVkt
leRTHgt08L6jyuynOmENOHF8b9BdgehX3gRuAMPttBJTVQO53n1Hv2yN+wo8/3GnXSsHDaphTKTh
VXBji+ftAcZs0WOpymkB8IofT1VrQlVZBkDHaK20UGDhZWEijrYqjc3nQLWunJBVqYo+xiuMm9iq
0+OzT2DGWPIg0YZrQ5jLH9Fjpo5px4jopD/ldj/9pksoiKaxa+Hga01XHTP4u6FGDEwLOYlfIglh
mRcj4aROzGjTUHDLAMkHVcv6O1SWOCvKWmCzjyk1ejjE6GXLNkB8GfP4nyfF59spzp/EPENu6G5i
2OXcDG18iznheLrNp7mmsruFByK5m5wDeFblH4QNfHflMi2n4QOh5UjTxPiBkHRf2yiDC2QT2+Kj
gFTFb8Eufp0hiFMQTGOf13i6azJT0+OCtFL04uGsYt47rlmR8IRpE2aXCOD7eJE2tzRuLgMTmuKf
raj1CLJ/UTXv9eJ41HMRsa+l1JdrcCuE8KcVlSyNqls/TOH/CrKiKu8Cta0vr3C2zOQmdAfq+JzN
REWdd/kX3sRF6YDZa+vuJE0c8fq5nzGTakv2xdDcPX5+xeRdmXrgRdwB4L6EhIdqotZjdOyOsDh3
u/pSvVaLggwHua+1gi4Mq5xz/gUn/AwKyji9R5Dwy02MBZyUTas8uaN7rVZS1Fq1jqhLFt7z5r4a
zR7ojUWwc5CokoX6QvKDvtedvjBEQbC/gnh/onqO0NZZY0yPPXFIeGLMQHxbPs9n7B4GjoBbTr6q
qe6XPcBZNFrrMMDuxIQ2mqmtRXduxxJqQlv89j2s7asHzYihwUMR/WrfSfTQmQQpcrS6u1r5tYzE
zQ12euaPGBGpndY1/Ml6fvjKPxyGd9C/CNf9eDBInGco7VopnTYf8+E7Izy05/zDndVFaj34xmpm
5C74a+bfEFbSNvE7gqjsOZ0X02cB+6bdprjeKSoT/GIQkbprAk5i26fw9bxSVvU+TL/Xw77WW6/1
7nHm8gJ/6Jk+ZfwpScTJJX/8omjkkVushBBGfrIZoaQP83zQbFHXjoXbyZEsnTqZrxT+hJZxLRNI
g6W1yab4uZ3mOrRf4fNRmPso6QBGsOip9ufg//9C3URVrWw7gBx8r5Q6Mb8JgBuJQOO+wNAW1kM3
dObTge+Z6ieZAUQWwSoT6ATSS5vVVsr2NHBYyCDpPosIF3ogBXuB5INkBnXv7oL3KnS/i77tan+j
DTflv5/CUlwU1spPi+oW/gY+XdW1W7Jk8n3I4UquuymRphBC+UCPA3rd53jbvGQETO5zQ4aw4vMT
V9YbwyAOMsuSoW+in9J3mSwM5m2QXb+wOy3ImToaYbnFSVNfU1cT0DTHAM1gSKEhZ9YZ9VlTjcBM
G+s8pw+5zJt5j4w9/ncEBnWCH8yf2Vs9HIoJ1lmECkarWCGzRfDiLd1qjwI1K4ubGzC5tLRl3HUy
UjLi/PjKjCeqfcGbk2tBershg2avbYJj6YrNrVXgGM2wSlTALqoYqFUu5r5bIS2FHG0uJA2N5jXK
lBRpl6xtcZWJSRXvdmMybNGqrOrEjRoF8dagCJaOLSAtV94O2cBFoFgqteHT2KYVfcivY2oXUuL1
i80IqaL4SFFivXiUPMoqI+yVPc4OQpAOzwZ/3E63SL/PJFAywTL2d6QlmD1l/MRSUYr5vmbOpKHj
NMU+E1y4ghkp0Pcf+Q3yWYCIqcYQh1kOhkTtGgYeL2IE8ePCN4wYNgM/Iyhy3EouC+NgrLRXPbC3
kev3xPKXSsDEq+Ye025nvjYqtwpd3LCLVaUXjqEw2vMBD/OJltMKwT2xnKNMyzrHeNhH1UHv0Qsj
HHYgOhiTqUvxAcPZ+MEDl+1frfjDu91t+32RrEQtA/X3pflg5yi4bGZc+GwMJUzyPrGL41oDkXhX
rhojqdywrEBWlGor6ti11FC6WVyd8bKbmAAooXlL0ORLI68LrU82qlIRdd/Z10vAN7PXq0Ta6sGM
wTgvN2TMankt2Q6dYoUE+BuCLo34KYfByPrJm+sS02b5ayygnO9hYnnBERayBM+KzX9P6Sj3A55D
gi9Wf1yDrvFtmuuHHrxsS2OIzwWUDaYzgIPybhXHJeSXXHaa9hwsuEmFYdJFmVUssvOzbSUKnIuR
RdokcyFkLBrp0lVQGW6VoGMWPCKj4oRZ4M28w+XfppXfcPAAWz6ife/29VPHxvppcVMocBZNR7WB
SVhkz6J4E4Y+7ui+Djdppujv9oBgG8xkZpQVM1EmeclaM/OUIHfYBq1UcuyieXKhlNUHYpFa1XAv
EG7Vsp8AwLQowBWb9TZNanHYVMwPlyXlwGnPstECAmaWrYzdtUrxkW9XN4kXLes8gUpXhxqt4nIH
jM0+KJNTj8NFSQpFKlQ3SIzdhK+CAYV4mUM7V8AmHUbAQMF9FVAHUldXU3umVumzxqt1zwzUExCV
S/uCpNWDezNHX3Ykh2dpz8ujS6mhbYai4JMSELNfqCdCfUkl5e0J3QoTroImQQM4CNm/Duv76RSW
w5YaZ7K45OXaYr0n7NTcjTvS405wMa4HqG/voD5XlaQNaCFgsYbrjoZBbYXgv995oAeax5TYFLVy
wqaro2Ioqt/CpHaQdozF1B0wXDZpe+LYjjUtesiSF2W7on31+NH1V5zUDoqOgxDVRxqxUSKNFBKh
wh2pU+RKF89ufgMh/c87a1kKlnrKuT0DFJFXFp076KLOfkaYTZtZFFKrjYv8L30xd2FzZScgSNXZ
3E3pMVgBoFW+EAJ9Fc488ZTBs0T7Dh0KjpEG1aIrU/raFXEQVKjOwInH2/qp13vktiy7OKp9yYCQ
DNJohuRmsjBL+wfbs8p+ifx3p/lWRDv8V5uzH5AZ74JKGzdv9gUtoXjK5JS4qN4CUVLZ8P1+fmDU
1Xs+A6cPnVbzPWpHvenSAAAASXNCgcwAGekz4jCv+AxL3XRFsKVQ03v4uHf+Yy3wLwzXWDlaI+ye
bIg+eWtJpudSZCKa7jIBVmeTzWdStz2ZjptwxZCT2+ahU716DnPAQOWVEEdF3ZNs4k/pg9o/v991
oyogUXEe89sVBvfJ3KErkKG3MtEAwx+ZWCj5RY6C3fnfD7Ize3jSw0LN6lEJ62Ac7v96hp3aPDUd
PHq3d/uBD7wxd8Ted6pYfN56KCukndOnlxiXnnjqLD5zYpOsQzgAhIkpBPdx0kYBCMGQAYgeZjGW
tSdoQ/hWDJQ/gZeQjAh7pZQER829KRD1lbT0Dep2HkpmJlUGAzCouAudAg8Majbx+znOWug+217H
eHWq8B5rPmTgaLkF3BN6IFef9s+cDe1guEa82tVmkLCZsX83/Jf2b7hMdOzyRIXayKm9hWMWGucF
/ucUNpOKVfZUVX0hSDcDPYA5rSWzuhl6Bfyp2QQYXP0nhzIL9MKa+017zD3wGCzPfKSPaJ1ZdZ/U
GsQM8uoNHpv2IUUld7s0bWd7+zeXaO2F0toWD8tnv+wHzBA/L7a9gaOKu7I/tLEN7VXEIXwJUePP
S5EETZdaOn67tWsngZbdfmK/kqQ0iNTzK+072GGDxAOvZWdX/6kE4vrep7cX8rGLOZp3obZiLE4V
PflmE8owmKLfWhmRpQVY3rAayYenknV+iOXadl+MDdPpYURCc0I5nrxdSCUO0Z+6SbExB1eu/GJs
+eHujw2LynfJuz/MDXr14594ARqEGAXQ2+oEXxUKCcA1dFsEWoHd4bJHGtdAKkDFRb7KlIBSYBth
Ym36aDH4GiAzjTuh2HbAaQ7O10VBXNTy2mSZaUj/XW3fzyanIlMxEe8TBYuQ3KN6vgxD7+2s6qUk
Cc7wvrZ2KMfK+dPF7J1Q5b/T3qgrMgOutyUiMGfi2rq5p1K8QsMhTHYAYoHm+lYN2oyuayQw5ko6
CWbxMHV9H4GpbOa1nU9Gne4Hbb8YSb6gpcHVgXX0ZVNroPWDhtGcMdiQAng+tTvgN0SJ7QcNEom3
Ze4nIozuSV+0/Jz6NuMYfQifXOsDfqdkgtph3C5snHIzMkde2/InutP61c3mcn4qqvgfzH1Zjk5J
/Pe9PUJA4ixLJmDQtxTKsFKERHK0oPk3j1a1QGCdXYIXrRdLhpZcnKNhr5zh3qGcCeMf9mK9eUm7
UbRqJB8oAXTC0QS3+7oqbXXXSlPOsNjAmPo86hVlmFXfaF/4k2eUPgwMXrxN8gJh2u9gpwHyaz8f
eR2mbeoHPqH+uQwfEAcHL0DDZeyHXVXBRNs3V9Z9ThONJhkbORC5qeRf2hs2k9FmlwrV+qLNCbRf
v9RKarqB39e5FNxUKsJm8ZV0NFcxWDH2Z+c+eC2+VoXcn6KK8WkeaPF4WoRZW8Gj1TbmFRgCfgck
OlKEHvnjLb5lxC7w38EcW85/DQe8qzXTb9wi5MKXvyRoyYcgafe8Dfbgw3rM24sjGZZ2yjKaXXDL
o+KjYIppnAc/7dP+nJ5P/e0dAi2JCuVkdr1M7TxXJzLC575qOX7ZL5fA1rMOi9/0aPpzqcCuc90A
jLA8NiMPBOnOSp6VenIoUm4mtHNHNKkJIlwdCZDdQVhHwqs2CScPF25Ds+hfTZII22kEVpr/xA8A
l6FmZ5zGCunuQp0QNmS4L22Ujg/5wl58AFrDFOSJfQEvfVGOEOhKPtL0xEUBc5ngMslBsVY2caGQ
fxhOeACzzNxwUCrvnGSRzUtfKJ4X6QMmS5bPJPksbYBXAQPrfx/J8wzMMiXVJ+DnBSiTBsMInn84
SQllJ/coUTmwaPE3dDFH46iU+RSaubgZFnpK/DIi28//qRpy1J2JJDFtHkma4yijKpwtzu3dtsQr
kK/fDAUyW/xkVRdqw2eLGjw4TDkrv1kVBoxXn43lLMyqxMRqMmEq/BEdMp43HnxQGzkAkpWXKmhc
lormX/yKkliS4DhizKR95rxUpugV81K8k4PTARGiozd1Csj+GBxb5X5G8LpvV5T9mDO9CnoFZUWP
fH8qgTV8LOv/3+LEAVXEdoe45QE49FaE1cxkG4YKdh8Rx2O/4BqXpUnE3S+ZDZNiDaXQ5n7SPKrK
yNXrXUVNV+zGZb04K5qO0V08si+CAwU+9bpxLnxMOCbsaxwE5kDDsIJfD1ay3T+61Ty6+P2rB0dn
RXEgqKGuUijrUz0r/ZiXuUuFMuAoxVZy3jeDljS1wELQ6kybf133LHhcYQnRW+Epgrodr6sIjLpV
Zh4LEqPH1EMlohS8EEvdOps6UaQ+ovPejWrVZGQSy4+QlCvXYMaMA3kTrIhbkddCUBDaH+vPbrY2
FBYYzswcd6RiVSTxT9+6MqorZS32ey6WekP2IgGvHBax1OAkHFtGcIPD/3gajz9tq/OF7JHoJm1h
KuaVxEKEox6a3EAecn4CK7C58thUNCY6n1oA6mLwBpiO8TA/ahFkJHzeS/uPvdRMcVR61BmpcVTV
rwTF4rRAh6BTQgG6JQnASNK7WZ5Ym3c18WqmnkLh6z2nE/JMm8pFDPqdF5nPIBDohWlw7M0Ov4KL
G+v4uh3w+4T+rcVHo08tSZ3/dS78csxsSbp4u+vsY6RqOvSuiSGknmdZVr+q/7E121tzNP0dnwwg
65Ech0P38ZZT9A/DYQYy3HXCKjLVctEBc8lsBvBCeW2Qw8190AtWppKOLVbOkUtgNP1VmWdl5qVn
DcyM8DwU4OabkSuOgEN3tLjivW4SKzAgFxgezyi+LqxMXFw6utm0ciB6vM1IH5AIHFkLNebjfoV2
9MBnPBUy93Wpax0i1L/to0cr5Mv0RIwSxpKGNfNEaCl7q7P7kOT761KUq/1J83Nlhb7+1dys7oo3
LKCa2GCj2ktF4Ihr9rilz5b0XftvkVg/H1uoCFpRkN00Ef9xKQy5kAOBzLfvMTJDaNS6r+33PQbY
wb3fxiIEFiYtTm3g8deSja5tVrAxu5sDAowMXnP9F0koqHQ2D5IlMDoHzClXnBYByrwADfAl3Uc0
ZtO7yb4XqUaFg8G8kOV1TeOedaQ1J7fIQXWnzhBZ6LThoUfw8RluQ4CJ6taktJvlcihJbseWlr4W
7t4qOqXI2XMSlnGx6rUlzO5hw8Bi7LAWCdvpIsKCccmd2HNQiP7Zy+xsgeZfut2WHB+lsdystzsX
q1ai/v9Y3I6LRQNnd/Jrv7/Sh5dmn8jydioD3VVtGZTbZfUlx0rEkah7ti6CjE6mjRptt+Oa+aiz
p9FOX2izTtt65G0tfflHdF9SV31z/lUrGlSC4jCv+9889BQ45oOnkUPeiDmdSUXHxkVQv2zeX8BF
yA2EFSKleiVfPwRci524WMxFlpq5obsflxXEd+Cu4glfOCovD6OdyHy9jy0w6aLRtskRFVh7ooiA
YrN6WRxwARROY8nX76LpI6MlpYMfDElDNcNvthuGucdlMNcvHfWjH60+RGiA+ulX01wyOGWrt6BQ
z0/D2uxfRastfApi/pcVxa0ECbUJ/W1FAAfZrt3em12qkIUGwjgsaFky3miqEWp9iLb4RvMCqzf5
d5Aj5NMd8jfiQ4ioFxJY3zgKkWfOUncLbdflq0C/Wu0XiToHfhmTURwa3276H39EpBG3SsrAb/Aw
qDS5nNWBuG4aA7hYpSjnQV3vN/OmzAP27ux9abcmNnSyvMPXp9ZZVKMGG7q/+AyOUfJZ73QzGh0m
fFo8qrxZWxYIglvhts7e90KHWKMX6wqqP2g8Rfiw2AVfM7AiL2+osZmlmP8Zh1+MNjONamwyfO50
jtpgKh+7gNGon0/CBCda6igPkjp33Q7zkff3r1wgWHDXT+tyKEIQZ9y1lJMZL8NryhsxoEVlIdqo
qC78DtKKRyrrde8NsLu9Gd+iOIYM1QaNCUrqH/K62ZZufSa2bA05RpzZX84smAeboE5y7hRqs2Oe
dtLcZ8qcELm8fyB9gQ09FFZ0seG8pb8byxaAOynbUML4J1MUl6DihpDVilGsVL7QP0CkeZ2QNVKE
dFKpJtT33HsVb8HUUKBBzMzvwZUFiArVvgKRHZNdG3dL8BpD2/PYqj78zJ9lKo7xB4a/9JmNvBYQ
UVuUGEyza3R0/ImOK4Apy3K7Ipn4HDouW9gUTT1AWsdElyMxZLAK0bHls4US/qLQUBULzBa8j3q6
BPoWIVZvtfni7kAmPSU5uwGaeO0vfImY8hikFfUoqvhcz5IJOK/nGTwJtXjHQrukIiDHKZ3yYraW
9qSPmg5QMSfxiAfZH22Bab5oITh1WP1MaW+NS5kRfnT3n2N3CS/y88oPmUsdaGxImgsCVs/UL5R0
YK/wFFrTTFBGS57jDI9mXLCph8JXA06abstosNBaiUkN3qePwlRPNN7PDRs7veH71JjhJF0Yhd4w
RC3yepSP4MOrcc18cugohC+lCAG7v2+ROonvoDFQ7mbABhEcBWow+tT2lM5rii9Zao9XdsgiRBiT
x/oYnl6d8CtOet+5SNKU9AzEqmoSpwXPJhIHU73AqbjMl0uZojkEyE7zJRxUpHzNbyglUNrUPo4f
O6RfgBesAPOpuO5sYDf1DWb/5r0WcAEQhMdqWSwChuRdroxYUty4NoGvJcIdUelX52dP5++jlxis
glMcIbL3cehFbklAayBB3upC91TvmwqsOns4JUiOp8ddZCK/MUzhrlsjUH0k/VtXI9/2rTZLIoYV
rZSsQfROU0S4fMJAjrGXj7vTP5YHKvkS+4Qpt/7iFFCdKkY1lXIqgxnNY5XKd9RXfdnlKimby+5F
lHr950oArzIhBeaXmOeegeWDDC29xwOymmIyhW5zdofU3fTpMY2Wf5LZ4e5tdouwDBEqJmxXUml+
CIwO/OmW3Xz6zW1NVnfECVzDI2snLTJw539xNhmSzy0aotVk4kiHl3lLgT142PpBfz7/L0Zc4Ioy
Ll11gA/WdP1qqJkghcpLvc1AD3v4futdZcNsM6xDf/PmIYVm8UQdMiakZboDLzudGArzPvmo4w7y
Q8hInVd8BcoopUmRcIjtTvQ1JeGz393w2N1e6UJUlFVvWIl53slZH7Sj9g3MlL71Lf4ylZ6t6ZYD
v63eg64DUNI+pdM/2h4yvdzjs2mY6TNQyOco6TN9xE7+TpjF1JbXTRFVMA+lfALan9Gi6dcJqA4D
U02K966a2k50MD+wOLUwLo9pIQzS97nR2siu6uZHi4ZfRiLKNQ1kilvtwREN0yQgGchJQJ6riMhz
4f3gYeqB25PWwehRB4qfY0K1GntDZ+RD51e3LxMw9TpaxZ0deGi3ffwCjgLHGE2gn1UkD/G1phkL
PjTEkQH9OFkOcnO0MgbMg9j0aoXtTFwohhrM/G2jhCK5Y3W+1Kd7LaUtni7cqRZ94MDMOX2yizCa
UMyBCnFX5MB/7K4RzI9NPicT2t45uGWRWMYV6eVbOLQTzdbKxaqn0H+Z9mdoGv2/IyLreww73My4
bN7QhzWyCsvkBt0Mqjc23a3D1Px9ORiY2feKqsSXZNplYXxKtdJjvxjeN3p2YFq8orKk7rGWkxQF
anb2p4Hbyvx7Ao3IoD0W+Gjby/uVw9RjmETs7jeVchJECjDE+SG/NOYvnnW7A6UrweR1QKjuwUJJ
5M2QwwyPxgxx6Vd6v7/qDJLFl5KYjfJeH72dU+tgoFWY8z+v8k8incgtZW79EQHAEiMQY4y9fO1F
ijO7hSdRU20IKZvcaYQqJsMz2c811Fn/eiIC4cKx+3HmqfbFZ+FcpgOjXGoeSJY28nbOJJRVECOm
y5qgN5YQHDlo9TukXANrto12oW2xAIHhXpTGSW06uxiYYdDDK73G9Q2ofoEqN7SrULA3PxZ9lxVm
F8jmHoZqOeHwFVIFaqE+AcbGo+uX06xlSFC22jRAYDRHj3SuRTbgxjye1H7iU7MLKiPpB2XDEQLk
NS6AiHM8RmsZrwLGTk7HLGVrqLtRNZF8KRy5RolCbyTMej78JUigppg61Lnq6MxK3EPqDdoBykB+
y9gOOzoQ1/JEHqtHez6huZduwDlrNyCwFVEX0Ksk6Zwke0RPWxx6e6TQcJhBnChJakEq+32Qd/ap
mPgPNDOizGAqiMea4kWPZ3W3wX6PgfTfKATBYjN2MaDKfu1MloCbD2IkFbWpiMRcJmoOPQJBdrpS
6f410bHJ6ruPLgrJdlC6mBwyb73nAIRGXjpmWlybZkTIuNyt1Ka2Ot0qkRopmpfkKSqJp2EuFQnU
JsZvIZiqBB99hWE9nNZQVBJvDHqFMT1K0lPjIfIJnfhaq4yYNLYNRAi182CBfjyJ/uour+cJaDgN
Pu0t5vLA109+V94WqQM8ggu4Y3uDVbIARhrtDBspKqGjd6PCSRa05FpsbCga/cUvWz5PEXroasMy
lLI61PXdtI6lRFlMNgWSjWlRJSQKnTm1hE3XpQraXwTqw/o26h6lfqnjNxldqlQ396LdvsShWumD
mLMW0DSNa53qZ6423N1hBuZYYSkkxCp8zHfmchXbmVKgAmqwCKv5O6Wk5gnWsF9dAx0tEdYc9/bW
EHLsikTUukOwoRUdlTcm+NJRvdshdcVNxZ6wbU49EyqnUWMwnkqdw4IzxeCe7d3NVRFexe0QfsR9
IUj0jyLZwvv5m6+REcuYktwI8y70+Fps50RtUp6uo+WKSUc6jhpvETovaV14C64yuA/+u8cBOJEC
jia0yqHkcqFH/94rm0I+cryAzID7AHgrccxUd/dQ+WePrjrT+qtvtM11j5KeTRbErgWvFmHFjk1T
0yOfTZa52Iq3TsyACZ4C14/70i9fFYkr8KyLGMeXieI/PFZpptnLqIDz5haV/Pli44Iu5jmB/7Bz
eA0GW9/HwWKa2qo77fSpKw4IFeykvxeWgz3cV6M9XXVFsqcGkL9CbwsIGjgAciXoVVL1snBJuoYm
YAFw9TReFCuZg+SCzMxEype7N7zV3ea6M5mBwLErjmvBDNk9IReVkIjdnX7SpzijYDxs9IEcCrPP
mWLZDzHpLURr92+b9MvIufPlpis86VnYSgnyPhfijOv1RSJ/Fj8WVMsK7CXT28QIO43hCkLezmcx
4t++kwZMztyepxFIy2PRoTQuoU1M6Oito8OEkEkGDAN1TYcvVsjLpGFZVgYiPmc6Jwq5XrAyO9Ja
OOQyQVc3+TQGSILBrJaMjOMCKiPY3QLKV/Qh8fpdZB8VhfTgq0CsrmTVikz0baXCIfyON0FTThUr
UGqmeTEVMou2dAL7dfMVj7O/1R+jTBJ12wH6Vbkp5AMIcWFYlk5lmD4D9DBtm6upw16zSzHfBwrw
266y1AHYDDn+PaWGPBOl5/EYqpXjfAc/vX8ULG8piVYeBElcla8u4N20I02qQSeA6zCiNRXL2bX2
Z3YypXkCHwI1656u+Tah7eXXF76lXcBeGnYQak93UVKrsVhsWBYhNbHUpXF8v2cUCese6dInkM6t
nNJu9XDMRq8APg3ytuOgbHrvoctM2GITFKnaiGvoFFXC+CrhPPqfEC3W6v6pFvujxXhxYknZCctX
ioXiw1xsmSAZZivD6JqdxQiBZRmWxRWXAfAMIxD3GFE1cCBX3HfApMHbZ3PKWtHsddI9lAW/SdD3
Rqk8wEZZGdGW0wE7lxLDNg3WthCVNtKuoGe09xU82OQxDc3b4PkXN8KuQKGyfpkzbzawc/ETdV/9
Tm2nwBtwy08knhq1bhajMsfz+85gfSXrr+abkjTUk8dH+2CWqsj6R7cJet8VLidGfj8bBlcPq23t
v+iYcdpNSh65UDTip1MWNd9zo1dP7JxFBMh4Gnybv7VxVUeU89m0bqjc6PMp9LCYjoDPhScaLSdU
5PeZFOFcaYR+5ymK0AHuV6uZTgkqyJ2O0HcK+rtgxp4dDGfzgchCng1gExEknqPm9sgicUumWblk
OsDL8YHMbcvRQcFGgGNWweoPpmCj1Qh4rLhRV0ibXRM5fLTnUN56af5lGRe+3MQMf4wrCpVqcyKT
NaU0G2n2mrlM6C7IbFEhfiF0591z2e3vw/iJGutj0zBJrl8xDxNfto1YtqwVu5ZnmaiXeIyzsk4M
XIjEcdKHPyYOKpYmXYXT4oeFPeXhlirz8557EAB8QU5Y9OoMfjxnkBGDynd3MXmOr2mGI0Y4x20E
7axm6RjFHO7fN/l4xWTGf/QohEZgaVdaIid/C92vCm5UcAh+J0DEPsMh7tEtnkGkfg3sLXNmqFIy
K6uHOBo1hl9eUR/ByrTOHsfZMOsDqUiCIQN21ei3qBEht0527bjttrzYvhX3djmXMl/W8KkGBpvh
ds0C4lO/N6f0m2nGQkUlcNvhuN/UghrYlsv7qw9EOJvsfRZfISfuU9nODayR5GugP/1mZdkj8dSM
6NYBmPhEZr9oW6VKqZrypjHGkfyn03rRhMpKW1Wamz9v8FkHpF8XEg18Zgu2Zle9TV4tqx34D05i
2LY3MFOGNxMdMaYstrqnXJ5dhgCigcjIqBluzs2lJ6zXPR78Lyawcc2zvYTGsfyqvdbGZO2pY1v1
gboEu6snrFZThiGieAi+rcHgLIyabOBKEGcci56DSv9bepOcEK8twfRmr8ajbcTs4GLkPv8FlLE5
4xJ6GbHyLdhFncJHatyfRPjw88Pq7e95qvNOxWAvadkQd4g20CqSYLa0JEttC47cqjcWw7MLHCuY
F8aFcGZu7pMWXIsrg3uV7cL8JabkDboObGBfVjPMgCqs4ONLk/gfcJo5MStLJoaQFiO6gUBH/Gy5
9WOemDnkqg129kv8DAOX1DFy5KTKcht0cA1QK6hYDXfknfNW2lIVlsT3C8Z90UWvfgcC3OilyF+m
1vekvsFzL/Oj0nP9hHXAj76EJaZyXXmyFT5r/fOmdeXKEXbHa+e1f6lXXCgfwQfuHk1WIL0TygPQ
k+RTRDKxK60x/4QhZhzduGwwlMg6UTet/5vbgski6SJDK1On6kK0Hrmra6qcUqeDBTVOJ23t9eCF
sGt9kOOJXvTrxwPkmF7PrtjVF2hHSZOuOL0WBmqHLpo0cj7cG9jQksySddg2o327qPYRKPCyBlha
2miq95ZaQbhx8dT11po5WJ8xU8VKxaUzClsE3qvOo91kglFom67ifZ+f9ZiMfWn9q6L3i1moog08
jeeAJ6VbQMNWEcr67jWZj6cuI2mW91HWhRPKJ5mz2hVuyefHUYE5WVq3E0z91SY6hVgt0Wd3Kwe8
e5N6WS3yE/zsECSUFL03C4t7I8xIr+5udwea2nPwdGUKRhmqxWYP427aHW8tvgRWNOxvkXXf452W
BEjkLjC3lhHXxjymmKRFlLe2EqxmvgFfUFYVdJporEHV3PYvOGBHhA3tKdkCDNldtVIzF7R7TwbB
Hqa7YCu5Lgfs3TYz+LgGL0qtj9EUzWHdnUSNKBdZRCszUUU3+zw5xn9AfxuNxppjOtq6xufgKoJU
L+HRYMJRxh7D+RAiMnjbWKgt/jUBWaerjpPLKWtWH0orN0Ux33FV1bklTFWHUtT2ja39Whoubye7
A8zV4fC3wiaJ9+kcE0onP7HdtuxFwzIrTfF3mP7NTgsWXbg3hULGRoDvB+Yo2nRIHCN0ll0H/+Ks
y5B7EbLIxsrfZPB38Kgj+gQ1mtMO525nbfR6gnA2p5k0g7zgW82hy8P+LkeO07+dASl9l0XWZw9Y
eL7S8jouMMVwp8SjHVIOARJqQGEmzH8SsgpsGH9uD2tNsiA3MheYsm7bZQR+NleN9svB4YK4GMyd
YbSv+Uux4kAkC2SqXUVQc5n+ZoYIqQdnGvNrFC0iTEzayxiSxDTv4jhQ47b9Lfcc2SqoKfInVQsr
Brc2bmm4zBxqez49W+KAwiJsJgSsrUZMy8QQ1v5nkPlUN34WeCfvILGchSDk+J2XADl8G3aRztJT
/KasZsjF73b1wIfh1dBKJBHW8qogIk/QWEVNqHJwEr5RACJZic9QHubZHWRfDRHI0gemYtwHfQ3Q
3TYa78FhthoMFX+Pf6oGJkopAInPO9v5niHBZY5Bsy+gcomlkeW77ox5hrvLZ5Y/Jn2IS6aNZgUF
oFQsG42GVenDVUY2MAU2u4PaWkEmvP+s7+7onu6L+mrBCHGMSaHzqe96o2zjgqGpyVdKpm1dvPG0
mNMPU5YkOK9ZJ+bcDofNPdjcwQ08+u0Z5a9X5rTSr0ZJ4p3Emxtgpj2pVd+QAmd8Ew5C3UWX9Vmr
N2Op29BGzZnw+FkAGvb7nhATuc0kM6AXeNJOKUgL7WB+0pQXecMn0k9n3E/8Q7sa8zE366APp3ME
/Vts4NJC0yPTRyTHvoOFqLM/qeu31sbT0wxsFVyTWdTB147lg8I3h4SrcZU0c0Cmis58rxPiyjg/
meuFD+ngFCEhAhtJHogpf8VdkOq2OteOrGd31y3eHR0JF2gr+Lfnz95RXZkKRa2i9iU6wR//ye7X
1KsjRxI/ZEFq/5DMeqGQ62Xr+aI4VBIwCLtZk01e12CjVbZO5PuqcYpT/TwHkIWKbnwd4dvUWWy3
uSgHmtcxuWPNQqb8jozuDo/a0cOZ6bgoGqgEDhFw9e4rNKlaoLl0PnFTPlwsa6x3YBgY16hR8Lk2
QW0zyDVenR2CpPgTZNz9fQaA6DEh9cL9hcDsOEe8Q6ZJCodP45Fb7vYnSYobxF1fMEWBIvzov3gc
l/Q37sCTCuUBJDPrWSQrIhgWtkwTKVgvr6MGZLBKb+g4cCfLk+OT93Xxivlm9x+VAIXI8TrQaoYq
A8BZM10tSB/d/Pcs6sL1bhj9nRpMlJEoKEv8mzht9E1a/NrMbbWjTkBdQZ+x2g+30AIe2MQPjIsn
L1AD3ZhuiQVao4IhSDKZV1txNStHr1FPNsbMaGagKAq7ZhQAe5PiJPWW2ANIaog1l9UT8MpKGi6M
Fu18EMUzqNN12X0vk6q7YPHKmS76eBnVCIt4zM8gPt6zTITUzRlSFRCmZjAn4L9JzEIhzOALzO5Z
3MUE6rll9rHXNu2rU92271nJZJkHXNeJzTPsT8+aTPyhxDkoCdkwHZ0xvyr8VPGnnZbHxeOa1PCA
G0Ps289lWUn+CpfqefqsfIRDacDCrNeoZquU3xEqVqvCn6pfRSpBEaoDxYCgwL65I14rHrLGxLA5
80BSVAmJHm1j1HBystn9VRga65kx26Ri9cJgJwLHKNi1umZrtF4bakp9kvAiHne4phoYHla9IrvR
wRvUazezfRBSCaZH0tcn9Ld0u92Wka8Ov28yJc6ChsQ1zda4dNOCzXh8PTXxKaWix4bG6ICZm9Zj
hYIHB4ZI8CdtcWtxfMC/6OjmrStd2shmW4WofQ6PsXfrSN+H0kC0oFHIYy06r4dy7FVsQdtO6hFn
pay6DDRyZiNWTjuZi5U9Ii2tlgXhIxGBc1C4yDGf7HGB01w9M6mburXGtMvBEhXRMgwuWidfUrE5
zchIuJwPbd4IcLEOjve9AIErNTcirLdOnOnmG8OfVQMNmc6S+7buoyMG8EdHnVOXqyQsMsVX29IE
UgbzkIegyQhNKMcpWxCB+ew/qzCy9c+8As8wrzh0L6Rd1mrjk3EBJw1/xdlB9cH3+r9U3x9q1AAW
MbKTjkOjcJX+ls0N5RmBs70C2US6srZ8ksW6Low0nh2yJqWUTRGB7DP2JDJxqu1GpBWDcz7VlgZ/
v5kW0Wgz5ncp+NdoX3enp3ubKQIFRE67UkRqk+A79uTIZAuGVB7G6fzO3mfQgkrOr5Lx5G+Y1/yH
31q4MvDdDw1odezhL7azHGh9Wzjs8pY9VtHmXWQ6zjAj+x/dpvON/C+97RL7OMhJxjAUbGLK4Bkg
wlnCtt7f510Ce1dldPYBuA7xnkV65/sO0355nyrC7cs6+bN3eceJArxrotKgybLwOSSVjeNXBPUD
1kKL+G4U75fhqXt0uFVYCjSdQSPQdBc4xQfrU5TA0hRktIOiHq1yu5dm6rmCQvxzmISLaE69UzHh
I3laiCKyQowDz7djP1fYFDWogtki9xqCGTpbLZ3tUmXJkcgOweS01LMJoCp3DxVSbuDibbgBEXTs
t25bX/aSIYyPFxZXtExc04OHNy6vWZcc0C+ZiZNLql8H8Cq9OobcYgHRCewZ9m0Ia/VMrkPM0ZlA
iRDJSc2ZSkGWEbaKfveZBnMobGJddSrftigHuh56YmVW+SNpQiM+bBYOFJfWSNrITYOYiqRRF+fh
Q2cXl4iD+YuIaYmsUZtflhzQVtHketzdMATOSOnYsg4FKndxDu9EKlJkIFUrTsTRXZLP92qQMR2u
POwd5BE9W1VVfxFcy/Lg3VyGgcipDzAsrRdsqZh55s8WqAMh+cu72EI2Z+fKhKC/KIrxRyNUMdgz
Eo2oMlEBwj8OWvGhx/dCFpFjNg1c+rgRPsd8yZfo3gPlYos+iQo26xojspihvxHCngrBiSUzHz6a
7f3dA4w0KpHakYFcUG23dWGrzZ8ygWJ2qvVUHizww65UkcOL1gmgtPmOV8AsnNGBJ1/njOMFgsN2
b8K12ruqLtHpLCDxpgKcHimSv9aOo1SwTfGk0ubbcCaoAmgnAMUN+p357eS4CzqcQQ7whMIIW04+
xZpwLLXe/HuSxCWkH4OOIiokPohMtdSpIhByjY8h/isDeJLBmSdfGFdY58byo/1uXVXLggii6/mY
YjnRoCd3Ux+YUYioSCmu1k2sY/H78m/WcDASSEQ9wVmuUi3BH6GFg+S5puD4wdIrHzaweJOwisRt
UpopQiL6zxhKLPVxmU5tLasT+HQPIhZCfzE3LPq6IwQIx1OzQAcK36RFGtAnpccWB+ayULhR7JPR
GopTc/V45egLWcZo7rRLIJ5TzdZfEaAAbxvY9hdYO4hUKJsqPYwzEyODXHoUMZZZpwDB0sAbrxSj
Mct7hueItq4+ya0+KK1urzlPcJvbDbEEfoSZ0O0dyxPvHYhaZC9Pz6BbQ+UKOLZz+o1Nf2Yekxsc
ZIKaGacQUeAAs1NBoz6WUBXKekQiuCc5zbP/y+CaXb0hvLXDLSJlXbA/RwH5Emjy+0B37EwT1xUC
3e8epRH/4rs9GA3L33x7XV5X4tflqo8p50As3cHgBHr/HoaUiLWSJ7km2VIbY5n17QBBuW4ry4oF
YjZniH7VCN0V+aA8tz50nFTp+i5n/RaqU3bKHcFQ0+ECO5K4t5MDFw7SYzUMQsph0Y/UibxQFPhg
DPVVZrwUFox4Oxrpw9vvLXgL+bqMWQfBcod80tLtqfw/x93tYrJH3Ad92FJinqUA0LBgl96DL+2R
ABd1iElvtTIcs1xLJ1XSuEeQyun9a380ZLiGQfDK9Q5btBBe8Q4PwYXc3czIVZ8vbfXTZVMJlO2k
iR4Gb9SpOuMqwDxMI5JSrrFBYIZW3HwuR3nuddYIVYtCIjGABN4oDj/SXXvxMpfFrGj20Zd8SGSN
BHe3mNJ3TcYN6nnBblyBok4MCGH/+Oisx9jG1mzgo47iUP4xCLNA1G1Gj0Iz7jvXIkueCsT9O/4I
1g0GYKpJiOZmOoHrLlrPRBs1iXBVoMqtuAcPN3jw692vayiGwKKMAfvMEq+WhwBVZMfYzfv44WQw
AnAuoHRt3bJnc/+X9K2cyRJEYWX4mwU/Th9SlCqyJ6DXrQY2lVyu00rh2cFJJkslYFlyYrYGh4ON
1qNeyonE2sXYjvUxT0wYEF63X8W7BLSTfhmT2l2bBwDBS7h989xLUPkUQuUk/n7YHbl2/K1Kt8JX
p7LoCvbHMc1zQ/Opryd3c/fdWsmmolXCc2/VrzrNPiw38BwClPLAwROyzMKcvRW7+LeXUPi8V4mo
+RLotmPABsma72319bg3SES4s+lxKuddrJJtnLl6Pq3WoCWp2qGS6X2b3CNnKRwZXathdDMir1kc
t/NnI43UlIgkZ6RxdCrvcYXNJhChbbOWgMnSEsCrMTqaZUjlEu+QVeGiDYwWi87JXc111KelFkL0
VCpCPsD3Hrr5RBVMwFE1IyXkue89pU5FLuaPsX0Vzf66OU6tRTBvsRQU7XL3soGuBDYyNmEbu2Xh
rjCCFijkpb7rwGUs1rjVMNM4QVxrO4siJ7YgaRYs3+AQ9zK5enDY0GkpFT3NQRny0cYscXEIwRj7
pdtD2+3wLSjXV5tdB+yiG9uES2/pW7mYMxn5ALXUHAq2NWE/ngHdF6OM2MI9p/NS/R541EZZ3FMr
cEEUqMFQGqCtE5pfuVbperCB9pqF2REx7Kv3eBbEgGUTer06TCtWTBBUZ//KdmVVDFc+mz/PQWvT
OhJ+a0jFPfwvnPVTHNLzgBUM5G5MyTwhCFYg7MZZUyMJk8UxAxRopDqJy51sGJwPXloojQft5wjT
ucUKnD8h/0HSK8lV5UCjD58QrBQVbINxBoC6ANyKUGHQNHnv+cVrG4gKFOqBUcvDH33/E4pGgZdl
cZLIc4rJlUHXK2hjeDVLuV/c5urpUwDtqSaT4K7F6NAo1eLKgjIr292qGYx6rJSOktjnJXTDphKr
/M39kF/I/+BIncvEDTB45DEZC/JGb1i0rUqpJ/dKPWhJMG8KDnM1K4uiufCH8wes7pfoe/xjxWUc
rtY2nwB6HHazgWw21hv1B0L/m7my2d0rbKIR0/aNU7wQxWSmdqLrjPr8XI9+JrAADtZwok+7sj7N
U4JKLhtKisGurmZUNz4U5MzEBIpIEqqVRYmai7HRBa8+DmAo80gpGaFK1RfeT+/PPhn/u7aa/xyk
2K6ux3vgpHusHcEHB4d3xFq9bk+C2w/1UHp8zNSTkTOCniM5+9VBZp1r53VZiO/Z/76eVK2Ctu7e
G+LAnSUUBYvHHn2NkSdJmrRoyPR4Nk5pYZW/n4KQNCU+5cPMwP1MC6qDxv/L7bCn15qZfsoNT/r9
sKca944BazVZFzis/2SKzMZTh3J1cZqh1vVYLGE+Xhbpcu9ptge1fZjQ8lc/dxOr7WEnobjtgqyX
f1kCPEunn/i1YSpkNK08c7H2N7ef8wpsIc3/t4ZGmMIa2F6o5vjIOrkLUl7+f7m88iIWY4sF9ief
PFR+HffGCsFeHKthbOu54Sr0X/xikg6zx+54D2e5untYwDlonAZFw048BFQAEjEmb67eu3bJpYsS
tpapFmk16ey0/kKa2abieIaQU8qzQ7dXhP4glQJV1wApKCMLooXbmvQMU5FamTmQN1d000tcgwcI
81Tv6wh015PhYuNt2hNq6u0BoYPAMrLfbD1tSGLZFm/88ZlorrhhJyI3icpgNq7NDpH+3418e9SM
6FHSD52OrtUS4iIFMv2y0yNPsclF4LA/KCKTYWDcn8uj/2yc3mDspSRfLM3bwqhtVmobG9M26S6a
54DvGrMZeeHouFBOlnGm9x6AfCtvzInHl+ulfe1TKeXSAbfCQhQBjrRH8dnk5CZ/mI+IkLwJL4BM
UTLvQZYsNdg8ne3duQOFmzFuv/fS6+4TI1uLB1SWDiEzmAr/5SGQH917HHJ0OudRK0RLs/fmL2Cb
gaURx+bHFbW4OJNyvs3XbSoOIa482QWplUxcUm7VxsuMdr92DyR+HAFBxlzHKh/cFhGexj6r9Bg7
xCHNAe2s/xw0Bag789Kf6z/Yj0f2gWZOH2wJda8WWPEC3qn6ZQ3jox1xJYuewUKRnFJ7ZpyIRnIa
6v/L7AOiIkv5WqkuryjDKy9uBuPSBSvTYBmnSHpJy9nR47tBEzWiDS1s2KJhjiq34kdMFq5VqnFG
xMzFjz+ZJAc7e8kIXV6U0pyC/m82LZebSJcvUTmK3ztggIw+A8SQzXqGbmixgeR0CqLyOFQOwONY
BQVVgl3z0R8gtVwnZWr/+q9RDR5cWezw9of7Cz32yqL8Uc0IkGs9+OuZ0iyW0oKpXaaI+TZqqz/0
qeaHo0AvEAyMwdtzpCUVDicor2IWyjIBcENB+X75UAAqzFQyopYmxDhM5CpFL5fFpRMk2SMYrC66
kRMJrA259ZmHG+fhmYqW8FPf68L+g+6Yv3EgAg94BQKXGiYjpAiFoQ6oZb6J12o7J3JUBp/o5D1A
JdXlYywxtClF2gIbJdwNDsHgzgBfYR4Vm/SJCClpqkuLUSWoJ2q2D6PccWQx8JgRArYVAD6a6QzW
StXSEH3pY9qKrgKBxNNR29VdWYtGOOa/sgmhTecf16v0Sx9tbTlz46sSYJ6Dv1WcWlHaNy4ALfOb
G31hd0gacQ8AmUzPAQSVQXSXl3cLf9j+XcsqBK29+hrc3Blp3j6fIVaqE7GFqm7l4V8buiZd5KmF
3pghPMt7DfMBHlByIQj9Jvh1VDNxVSubGh/fcz2ezVcpbRW+e+satn8ZxJQ18IoFpjbndvToDY6C
7n1ITMvYpf7cb2lf/DFIGMo/kUVItBwbScREiNAtyx+Kc2CkLNQZAprxqavQrPoaj+24BqxCbHSN
htiZs4/FrIWs2PPfaJQRpR6UQkHzOErP4xTObIsUM6ORa9wp/Fu6mHXxelJhP914HkT9Tq29yeST
QJKpk0nfcVLhQIEhNWCDTfe7Z/V2ryIm96lB0PX0HRWzNbgbWqkcWN1xvIz8Sqq3xDYmWIlq6NC5
5i5GWw86MnXfw5mOGWNHXU1neo7/+GFftZnP4Y/jhSk6ZiE9WX/ydTvjXvphgMGdvz45x/miXJ+X
Eq63GSEnIZLStGtyrTrJqpzrR+g/y3gakTRhoWfKmqrbah3Qq4pHGjwi1mPxjz0uzQYLXTIJBt+c
BrNepx1fzQNAi6qQZKSYdwhMLkxrFxlRgt+GyM5vdEU+VGUPLmZ/R1P8lh8xccCnkcG1c0cuqup8
mstjQtiraDf/rM+je0ylscLAuSd8vtSVfbuy5h8TO1gdN1iWHIoNW/e96VKGYu1vHDHX/AYkjinN
WmVX+MtdD4HWSlTRtYNRhBkjBCEuC8SV44Tfty7e5U6S0WQoTzqlYap/4jDwQtqzKzzPr0opMhEa
FvzKNcJA4/o6yBB1DZ0I1UiotQiiiXlKLABjxvBqMMlQeTvC/hBNuYxA/v9vRnaWJcIgQilClj+u
2FLOnD3y42fMr7XXpmbHVXZIwzdtc8tihP6fAFV4Ooo8M65y3RcOxFHkfs5lgVZCFnbW6bMYC9xS
Ke7j14O5QQx5Ga0xmwTFXGtSBFug7wFNpHCw94+atAWl2N34GlB+jFt9n4ALhzYRV0Zp15Y3T8hn
sjCdOpxJABzzWeCx5ydsbxXSwY4CWFNqOCY65aUYBd+Qrw6JTHEz9vMmLc2kLGIw2PtTxCIROs1T
FlfjEASz9lw+lUw8pQEPo5F/q1gWFp7mTNYnotw2cS4bfZjo7uSDeJpubqeQEiOaTxr3PGPu4yY0
EpKCSLGlGpGHNFnqfpXQtntQwFzop9oKd2eyyr2g69hnIHCzWDiuOzjZl0qTshOKPJ+C1ca4BOBn
PZGEthwwWRyiRQI2Lg6p3IHDvL6g3nyMmrVO6WP7fzO2MBCxAWLDkOOYOWS0vgYD1P2CPrOErdpe
7uSDXtqex7dwwu9oRq/Nm8qptK+VVbcSeyhwsgZQsTWQBqKboIYVMyji6gwPfAy0f5eOshSLV6No
VBFHQE3j9h19CZKgrSdyMWWYJ6vihzf/CsmLCApGdHnF7kNOKpZ/SEUHlw6BfAOkMbuk9FRv6laN
RtjSy944dyLnzraCPwzH0Th27uuxG4WupcNh8u/Q8Xwh/H+YncG3dZg90ROpZsNjBG22WFa5s378
ofYrZq64mfQ41pAR+W7hM9gLWzJBMOyGVALuBWkalxvqOAEGLxuQD/xU1DiJo47IccDAqLes8ulP
o98nY0VvyncIrWYaIyppEbDaQKx8Rn5x41+tQMhNHAnQRox1u3ytf2xzaHGh2/yU7l4NlRyCWJrE
JbnWaIFRuRR5Jl2VnxJoGbyOEbJd398IxicMJgDHrybgzFSw+xXMf7yxmsMfIPFkFr/xUX58YV6n
v27y6DU2O5U+I9hFKD6iuXqkCm4TL+qVNkeuSx0ZN4wb4+ZY9fpLXLMM61XiIz4+AnsS2LcJnGmt
RLamdxZXx/+mIfmcLmP7Ufl9QrO8Vrrm2E2xf2BfwjGm3bVj6SZpXaZXH6S+DbgkrPeT3bFbwNC+
O8Juh6LRMSjmb7ZDnCaNNHI+lXEZUsHU2/9BmKUwR0lYmnERolE2N+PoJe32moRUm5n15IOL/vlu
nPhouauam7PZNOyVmvggoNsJZU9MkFezCsDGOek2SPZJAZLgGM3uv81IXQjGW2SY52vwMUr0hMee
IxuLt5JEKRwRhP5bCWM6YPeqF7vYznO27LQrHal6lW4oDu9+3p+PYIylCuwJ3TnVPEKT6jX8PmEr
mf2Znr3UPzYNv1y4ZlLIEc1fqoCrIxYFyojLyfTt94cPpIoCfx9oFPWqT9ES+EVRS6jzMOqBSyeY
v0LRfSzZcEh88MwAz+5TZKWbIGjhZ/FOULDG4kjClQ6q5ezuovaDn9pLw8/v0eVRBGV3AIAC0aou
xfMinuBSF9rwHpqDVkASsJdBz3lC2e5vAd5AcXIPtTmUnJjbR6C+Deq1cttZCTBUF20YCZHHOZ3t
r+8t4Yc5nYPiIn9OiHzuS0HYkcGjM5MFUgegHsCilNvOPsK8YkoQ+kaozHBxHsRV2n76FWWgYR/f
MXCV+yoaUHPKFGCF7JYWhax0gssyAuaEGxjdKsycclBhf2+STzUheXXo7Q/CqCVQLYIt8qzQRPBW
yBMPsr/Xr3Bp4qRZa/LMO9L51RVVB3+99XzoItv8ci9K4ZYxrC1lkGvke/Ck9CVtYHvvLRSzSrcl
NBpVOg5Mgyu7poL8QQJrEsPq+D889zPQ0z81IhZ+B4ajqtxUv2Veb54RRg3HAKAxYI2LP0fPpcXI
sfHXuLiVHT1tWManddZFqIggpZiOwanBjLQhKbk/bGaq8PVFb29klc9TX7B7IIgIudruEzTLfkdk
IWxwVO3BDcqUlR+VL/r5TYMbfl/Z87MYKP+rQ293Bmwa9iOGJHLIh84A0yvRnBL1XEUXVC7dSnra
pa0sBBjJh9B2/sSlach1IfaQdRMmUeXQu6f7TN7C6w8ssD5s/q3XlyMWXFUwQh2edOUrHbku6JL9
pttg0DHyNe3qLIwPSjh7d2m8FId2c/D7tiHuU1Dm8KKjeOkNJmSBeokmlus3YBEiTVhv1P9LKgMk
77lsca6yQZMD1qxkj1DNkM81Aruj8zvDc16EcS33Ap1jAX7nOHfJK5/7nzTk2OSko04vkZC3bqok
LYIRx2Ubti2yFLJ5dLemHRqvMbTuyFRfg6vyZDP3ywhgR6RmDfNOC+aQEl370v6zRsVzZyG5Fo92
kHhiqZ09KbfBkVh2T3VNc5X8RtBxi+P+D5HJYUXSe1QjSC/jJKD7TR+x47PJyMeuyaTdXo+jTkC0
FE18WuxmGUwEPwtHOreWsxygBC2mRJ0rPFjUNRo78fWHK++zJ/uL+YENwzGLvWzSOPZq6JQ2fprA
waHuSvAmYTRBoUeYQuKz58jlEFdMQjyLEj0dRUnGJNakbzJkQMW26RWVXTrcv9pkznVJgW5UhOlb
LBwMA3VsiXyeIi1XyGRGbE/PEk5UQK8W2Yg5EdG2Ib36SuYuHj+ZG1ZLEldAk5iEKGhCaU1a6xeg
EgFNoqa2bNg/rQelLDf9AMklb9xmbJ3vDn5TzN9tI8RcBxLL+/Jq5Qs4GobUHgCqC4/hIDcoipA4
RuS0PDPu0jAGEdu/mIO2xoeYBvxySpY/mE6b7KoLLyslygUIHKfWWsaCU2Qj2ZEDrqT9jLnf9M40
QpE5g5Oa7j+Oe66iDTyiLBY3RVLpsCz7eBCH+xa2IQiygtQlNVv+MfQdm28JwQn8IipnHByC75xK
SsRMvOzJr4KcA9BF265gu+OcmX/MkHdbAuqYDI46d4SlD7J2SDjKF8GY5mGF3boFafkPm0ZadNOm
sYu9QD3A8LOapcdBH88w9hXQGpbDNRNOR3U2Tx5u/iBnjI4dwYDaXbnabgCYulQGoSMEyE3Ncj5T
WlAb7jRSWc4Lt9CjzdpGrC4VePXpfmljk/pJoCkewkKQ1k57sgl30apQjzNvhRuRZhPJjqr57pTz
mWRAP11tVoDIblVqY/HK7H9gqMax4/iAIrU/nRzouGgtCRacFbsr6/t8FVGcxdybJaktxWd+sPXz
cP5b3CWV1me6qE0Qwmty/N9SAApeaNvpCP5J18CQxF0hZyeFUzuqp9G5Crq6DLoNKGuRbpnXiBIm
K2lD3aH2USDyG9gXFpiT0ruGaOdGqQED+zA6b7uXZJLtL4uH6lXZ3ypYwI47BBjjW6m+4QHTeyWQ
ej7YeFjgSl9VHhmyWwJPsLE2WvYlTqrUUa9yf/i/TOeeRLHfEvaWgMVXpYhrrE2clnvTTKj03qe2
rhxMVA1G3Mc261wMsxChgjflfNC8Ds6y4rqomlhx4UPCDXWSuqD1n6cQuJSI0qP+fkyIegayW4/8
IdlSHPTg6zxYEuEo8W40nTgGc5rey62TcylDxc+yd4cQQ0sOLi1r1G5h2remeIAJorNSFd7cxFMo
CrVJ7r/9I+ejku3SED/NPTQPvMrDn8561LpD1EPhrdbLWj0JG+3nhCRjN2WI4C9v904Qj9oP2gz5
6rMENcqpgymJ7E5cPqhtsLRnDX21K4TL2ODuqO7B5Ft5DDJQe9bSofuqiUXkrQW6nekhgDI3nHkk
Kt8rDjeLfct4AQ403JNGSaXPy3ZuPwFWY+KTK4N8+8Qmf2yvlEhL//4no398VHY01DlVIno5CaSU
37UcpQ1nFkApTj/fLvwMdX6oKcAmbQV2TDQuI61TAC1QbcZoBcmLz6sonY7P04pYgqVj4CwjR5Hb
hfejqIL+ih0S1Z8RDlHvcslFJEd7IeZ451QANAxtpkEijBlVhvG1QXgmtGebNo8f1c2A3WkdKI6w
g0bnzemsqXBAU6kP9Rvsu+AFDGB1UAitAIiSIBrUBS9tfJE0J50/sPk8eDs9tyDdG5buHSsisMd+
JevzicjVNiWiPYpIMvaSDUfj+bdlVZYczU8Y1OQt5oK/H0qe4jLDf5rWlh4362ta4GaaTVVCF0zL
snSZqnHxeMZYwQaFe9Si5UMdaUJWbF1C4dOLf2XsLu5T/jHJIRy8HJKr60Yr3LPdTyYxDzuqyh6/
pIV90cR4gqrvmcKvdsvQTtfJXQ0nLwI6fsKTcl1hl+DUXpEHcqIbbwsh0alH244xcb7Ki/vup7U2
cgF9hPS0BbtiRFwWP4ZEtD7fu1wXwHGWEvsycR6dN1EOvaeMF3sG3FL6rmfD3teeRHYqtywW1g6A
kgC1EDIeM26XKGErkVRCo7A22JFX9QfWD/B0/XCcUP8tQDU8xaw94sY1dwa6XtV0S0+LtZ5CL1T9
dwL5V5K60MmeJInSgVtV0+tHneb/p4Rq3sisF4wO8I0Ddpr6PnWedD7SN/bXpmg1OaXfr3Tsm5TT
AYvGMS+iJbPUu1KQ8+cQIMOcWTV/l3tSMTFxtbghZmy8J9QlRxLqTpoLrVvcV6tyFz5uZL4fYbT2
LduJEJw6fDLNr/TyBqBLijatyt0Y6yRgTRP3hmbEq0mmf/UUF7oCmwA8j8v0EjbDHUA939+yCt57
j12p5mO5p5ePHA0UzinzS6qrW9C4L3Wim6pUcJPaMy3Fq7MIRB4q1ssuCPoBj9bX13CKshChHWWH
DdB723BdwKgM4zzqHYGHqu4F3ef/PZ0Z9OPR4l8se6M/AlJDwzI1a1LsDDxbntpQofLz4UJ1c7YN
yd8kedIogR2yhdV2lkOozuIRSsglD734prT2rYqBI6CyVNDkhajK9uRs+sq85SPmh2v06G56yM7y
TmrPRi34+zi+9928aym2yzyiQbNPL0E20W29Mc3JfgNtvHrTDkPy5+ep49d8FSlymWvb/DsEZAV6
E1WlS6f6oZsktjHajVf0XilvDMuRaR2y5JbFaRSlxz9GZC8cDXA+UOU97slxN+/VB4fDIer0rUpG
OqKRr9VrMvMCpR1Y1GE0jo/3qD0jRUJodtNOgPxWlX2ASymhHDJHmsWHC/2UA7Mgc0ty139qiFrU
uqRC5DTniqfWFalSkxKov14laGSFTPcB0voRWyjnRXdLnZkDBi3nysiSxA5vxhN8vybC3hit98NM
5KbhHoXyHP9tcU3bwR2Bzq2C6uveTd91OsChOkr0mbKlHQS45vizto5WW8pGOAW9EqjSWYvLDbbb
BGaftyVLaY2A4e057jwkk49NE+W511QN5KOujrEpr+Y3Wb43zqGNq8sDA6sn2a2oMqMNQx9OM+WV
5ZUnPw54DpA2hPQFqywa8u6dRXmiojD18/+KdM8gSsbcWKG+y6jcfcw3SPzMtcNNXzCQcF1BiiHC
Us2oRARloAxGwP7q6mb3WCuJpyeFFYK7aRX9/bC8R+bNvnbiHNsiAqoSAWqgWjCPqpFkeTQa99Nh
EeyHnmykARfYAJRgbq6e0bsGYE7m3ToSI2Z9ZrwCVuy3vqzdKeAUCTE1nOaEYS6IY/cfnJRtTtKD
xgHPpzY9KAo/k4RNk8xu2idoRK1uURDj3NrtqOsyecFQ5HR/fTtysxsVeoMKZ4MRwpTuzO32/ZiP
Z4tIie8aKmHs5dAb9AZgppMfa/GSdY6IMtyX9K4X99P0cQFmthvr/IiVLArkbS6gHFfAagTMtvvY
CVF8cvvt4Ge6WiQDrV4PBufgM273B7H+K9N4AgRtijetj3aG2FJl27atog/Am4LNQglv8OJVMoHH
TTO1MWSogcRUMQNO2UcR8gmYrXWmPsoqoAmZsxAJzkA0xE8tclhdTPlaFTPV8Ct2lDCZJJ8E373b
90GUHYq8v5o01szwsWKZaznR0cqLMIqGo1ALkoV8CNWXkVYOQqfbWvQEIz9DOhBa5B2phZRSRyPM
KgAyOePre9m38ex+9KEfp/MiZ0xrv6rQWTVK9+o5OxEKHqYkK8MOOPcJOm5IXybsTkSqohOPvUIq
7wuKQKCzmhiyi5HyPfgrLg146UrRGsNvZS/XzqtQ0e09Z4qiRUUprIu4fyy7jgtTXKCBDGYV3sFB
F5QC8S9INo2Y2hbOyKqqT3eGX4whcrU45F5zvaCuAdxyC++rIpSILkFS8GkP07RgNwxzTnbLE/6s
0AisxUxhC33GnwgECFbggcGoOyVpVRDl8KTrruzLUiAim2FWjIPpHBZ7cYZTazCdnIPX9iRyPyfI
v91KInWCGyoNsA1nX7RGkgequFFlKIm/yiXsjCPpNYcnd1XpMDuCDxLayzmSUO1MM627H88XAn4T
5Bvj5CRZ0dJ9kOVvon76e8STtEugc7WwxDHdGs8Z9qNmclE+Vm8ZJM9Z15pWF6AG1mXuWSHToK8T
uyCaCIOP/jPCSEsGZW7cneV6/tkFTTlm87NNdKXeS1TnHGLyhDxA1yFuntKfEjonrP6No6u95KXJ
hqyvWaPCAo6bUozm/taYf53WUxlTIF3YDMZ05HQW1zhSQ2ZuOcocrtgquREoF+r40ObkXAnm2TSm
nqS5LliEGnRFVQ4phQ6MlyBZC569KQqiK3n/SNDai2RtjwcuPzdgtkODDXrc5/cTdx5op8fEEbzI
lYONfp8W8+rKsLk/UUA4sLEIryVEar1eqxPsUNIcfs2hx786SgsL0c8BEZXNVodSAX54o7rYVqCN
YTvAK7GRSZmEaJq45zTieu6LC8cacv2J6QTh98GltHYqJNSH9hWMYPK0cmpmNltjnB4nG2dfcpcX
IvhX1geaeyXMo/8jJAGf5GNt6hO2vt7uXyqTM1711x2LvM1Tm/j/h8L01qyQdK26Rzh+sMVGvskO
MHoKvsm5Cljmahy7ZNBJo1COd74QLHKKEGWKMjpk7lDU0EWkT98v0S0WAAx9v5Xh0FYk397XYpxQ
pCmylFPKkr1BiJNOTvBEp13GJ2jHHZ2yGiLskdHFi+pxag1HBAnXits0v8IhSho+2aD3XoL3RSQO
sAWq5c+JQbUH/c8FhKruZdRlGeGaLvt3j4/hxJwRBVIsjneIMywsicwY4Sl1g26QYZ7yf+Q5Hr9Q
C5Jz4oY+BQzAIfszjWDHaGVY9K7bZYKcJsfLc/i2twtYxXzqcRofGrvIOf9FMhTYGMofPmDcwtLd
bwiT7Pmsz0bRUFWSmdy/PosHS75qMrxBFTm78h+jdkBslcrGZpsju2UFFIX0O3RY1vewcIypZPCh
9QZqj3ziOHZ+qkD4wpwjnHRx73FgMbo8kF2BwXyFjXL/hLs+0CE1dzA4VYKp0mXamV/Zemo2Bj9x
40HpWf5FctpDKeC+LakIsmbcTzErJM1Xcqpihp31xcL/rbtMUffZK2Z/QPoVAxr3Xsqyiaj65BK/
X0ioc+NXr/mY2lvCb7UFOgVSJIb2NrCDA++P+ZPJcb/35hbqNHEm9LXUJ6bMqNWIomFlMzhy4ZbX
gJb8hfDPkUHHUAPAeETxIrUh7Bent06yiJrDPcUjeORZmIh6sNTJGFKWN0GgeV1oWPUPU5bmGLoD
PGLIXkGvYFzAb4VxYwLS4I6H2Oi5+CKVO2jOs8RBzWJXOlNIRrCliU0CTtAVFYu0zcKoHN0k0LYo
FjxEuCdngojMnI28XtSb9xMUMMWDf/vVPXevJwxqO+9FRQQextBhfRjH3+rzYqZTcnI0AFX1Tu6V
K4j23hINDdoUx3wLVdIlj42jfeUkWid9FGMzPJ+j5vzoSFYrf86ZjAcp45gWeb3K9ap95MUuuzGt
aicLs2PmYanS5EI3YYABOfXd/Z1L7zB+ONpXi8/mmGASla0KrqDGkSMAUFMdpcH74H2GcKMnO3Pv
qvAGbEWDRdS4B4xj1VeF7cHTf29MXTWO903PHDyul8drbBkil7vexjRMFlMHtqmXtKRYCijhq3Rm
ZZOQjbTumk0wYdft9ckW6RR3T9uy4tEciXa9R/vxIJrjXQhviQI5InS7BJEaUh6IUxAtB93T2N43
7qLuUJCI7n7SlKRdnlgDJTP6OEgTk7/6gjYunhaEdlbXJ79+AGl5iXX1mqfXG/JenTedPVBnznzF
xfrq7Lk6gw7uJcVgPMG8FKZ0Fuk8G3JYjDF6R7x8rLibq2gTvifyxRw+EVCEmu9/cVKItI6GUvQl
WhIwiz8iY8iriWHmuPJHtWzyPk3uFz6XN2JUVMKW6gTunhrC5jjvu4u/VGHsZB7qtF5z87GKYfnu
G44A6Ef/jBw4mms07UaO1ccPcdRvEP/JS+j/1xE/m9SCPVmCFAfMaIX9HbdF0gnjs2luBhUch88H
XuFPggg+Wpiy5F3krC+R3CFFyTCwOmEvUGFhkuo8C/a2/8EUV4s93Kb9OCZAg5zvX0R3uXsMdnNU
qps10S3v++ZKcugKYBb3+vHea6TZ+ATwjgi07V+7vCcJ+XYiPLJRmaj442hDDBsLFGvYnsISTFvM
aqXq3bBN37vDWaJ5ew8vEjeyk+tAjl5ExsaxQ3dN36o8msQpVXwdWagFuzXzC8RvIcetLP//XQlU
M26BlKZQyjE90rHmLNBvFGhL6CZwfWe2pPrQzIvEZYPw+AuwUlgfVwKL+dq8eGeRmWrfwQtYOlR/
vWjkcb4KJaOTjACiL+3eF3efdJlVTaHJl8qXMQHG4Bvj7mEhWuSRa9ItiOKADQQW7dAig0vTGE4k
5GlEYjjcL9HgqvW2laY4B0+IiPzC9P2IwNe9HsRzJmC94ULOg7661nx6DYOK6hbAlHW9CooarDSD
Uxl2wurbMUv1uzIsuzLfhSOda4XdmyAp/9NgQpFdCcaLThczV6RQBCNnCRYwoS/JAEfVRKqoRvHX
ToM79phDiyEjP3S0hL24Bj5EDCq8rC6IQL6RjyHkDuwTPuzAs+8g4+MvGR8b/Gzh7aueLJaVnMfk
aWqOjnsMyitDI6Ct1YHO3IjW2Ac28KnoaN4FzkWKRUdL3X1o5qufNwzoV87TZp9LGbftZruPwcpB
/OcCF0T2wt5/ScnX7DN69VB1FbO0IyRIuouq0ogncUNX0wPyaumrOXL62kLZ6Xt+qtCY/OzkqS+n
XlWsPDFn13xPErPlPp5+jO93GmENdevJf111kuCi22uA47ulmgaxWXS3uaanhjS9NJdV1RjDzWUC
k+/3o3jawBafUIS6vkugGaCOB4GxdLvDL/JX8jR4SW9MrFe6ywDrv/zj6tdb8VGxiiAwTpUuKH6D
ioQHAMXi7xVwJqas5afUdDgWkjJ4adq42lopA/85lY27l2Ty+B95sskBGrrl2n/sLlBLgS+cGtDf
61k9WjZXq6vY7IDmVWa7MrQJfSlGqCdrN6uW/02+cRgSujIv4OfGdTW4c2ulJZ9DejlatkWQ3lfX
FuUCr6H358BGYm68ItC6Nc7C3RQabi0vtz6JeA0gcOlAMwFfrw3Lzwv8plYY6NBcLMOIPIIUpZ95
wMrFRtkSi3X+//UpmLDvtxo9NKfDuVZwdLxGGIbza5bANqPq5tKwcMKsfzBOdm8QC89bLsMLbMwp
sC1+E01nz0WdomZMzbLycUew528Qv4kjMhY/Qy34TM/oOKXKE5z2DIyk9r0rwsoMtvxllJsv2BP1
6v3BanDd7BxMABAuu6YVMjDHKIMc5D+IkHvXD/jFEyqqZKzFZQG0iS7Vf6KOmIADisTyvAV5GscQ
9fSz+jYVkTGhEZTrXYwfgwywcNqxMhpdnEV2bKKWstbwmbL9om9uPCb4quT7fJroDw1Epk9dVwkV
HVT/9kAsvLkEi4wKj8btZ4XlTpK/Tc4ZrdaZq3zDDLn3FHLao/lXKDXJR+7D3pQpCKeTWUz8o8Kq
hjcksRQbRMVxGYNDQoRc0WHlSKZS0J81DZVzxfUenQN1HnWEOduQ+YAiNpY9sG13BS7rptAdDgNR
FPTmdrRN2G/S3qo2IDH3jjyW75H9Oz7F23jN2VXNn1iHHw5mnEBrsIvaJ99gBaO1fKdVuTgirW/m
6xG+SqoBixDFQIshuprXJa0lIbf15vyIVTe300IZxyogKiQhZlFR+X7e7g/uz5XMrvE64ObPZdgJ
zxsxCAuuc4h+YwPrd6eb+q7ailQ8S4DOny+1nmhoG/KX3QO+1455Pa7R6Ku5Qob5wXh9PUm67q3S
2FxBtkgKd4raqeK881PtuuGk7S96yqAMSb3YLiY1WYQjU/2aTr8+rnV5zVUyqI6ovCKXnRHgkrGZ
CNfWokinyj3gTTZ3Fx90w55DUNBi/xFb3pKww4wjEcOg8SKKKP/8ZUJzeWr+l7FuInyHdiyTJ+jC
YAvQNgezg8C8hPBBu9e4u8HkVDEFBMoJtPXeDbFPh4yNdYe9cLQ1XGzophf5aBCoa0c70my6CqvQ
3hn+X9tsUh9MVepLsIYrfTMyPyWV0EHkIs3eFZiZpE5z6qs83BLI/vt9PsBaZ6I5gZPsxENqF+jq
8SDfePnqA18Ei9Nvm3vm3D7giT5mKWaVYv14apu7HhQYUvOZ4mShn4c7gpkX77AwU2/RuP63CLfE
E6mbg5UtXwumP6Zmb+4C4XWv93V5ioZ1S47R3Cta2KtPzxpvFtJ8DiD4FHqp7/UlQ1iww6+oC+cE
jkXuDR6l0A807EayeVP/uL8PFLNiqLiZ/EX8sEvH3xKU9k2WI4yqybbQVEtDlE9C1IqLPg51MwnL
dvXSuL6tC0Kdd7Vf5xlizv64gAM1QvBToX5fI1TIB2jDqO0mxS65bcPfgyLFupXMKoC9AZRVeL+3
+w60XJvqDrxaLmzsVdgVwK7RNYf3o2ZENz4zvXmapMIYPCzudd21sjnvYRZRA/WX7lYfRdqhtnqi
a02cccpHQsFjebpqeXvk3qih9NfL6jcYWB5STWINeAcZ3nPJlho9UQcxa42T5/PwLN2g1RZDrCLZ
Nx5Ws6SOH9/Riu3oNWOXrsHNpBdNteikpKgjM09xbLv8qDmRNLpvqcpCWr+MyXlI0bBDpf6LKLNe
sPNp5BoVpREAU5RCAmoKL9RXqQrvh4LR8VpKVY3Vo7AtpOuwlCfJfRglxRRXm5RIRkylO0t4r/Lo
CbbJo8RsEqHyTpwA4UBk7yEyBI23tT1XxKzLToGfOzK5jMSkoxNZDz9c6HyW9bzJyeSuHL/bDtCv
s8b57DGrKG2/LlEtckxW/TfqUP+l4cqipQIZf7PXHTMX8T9f6UHLfPCvaLH85bKLgn1/mjYaG3A3
c6WPIRbvKK/8cQ7mpWwoojj2UNTF/wK9/HrgHXssMThOSjN1dSqluklmtbkOrbGskHSR/tEZH7FX
MG9IZAVq3ks+zftuY3dPYnjYwqrO4iguxoy/prE/oQtf2aCPRXg9zzR2XbraBcUZ2nXvgiOWn1Da
EA7ePIWZZBOq7vzWxWO7dRV8/4YCuugntXe9fMNeMX/5HZ0eWS7pW5iowvxhxx0H/D9GjNnzF/nO
Bb3PEkCZt0GfAoB3le4rMd64G+9EdTOYj0SjCTqgwk7PFr1FxOfE1FrWgg5IBDkCHbYdIj2DgQLL
0O1bjdgcs2q+B0RzAdH8iPrYK/mRywMtBZNYGa/TGoA4S6g3blvbGkJ3htXro4zAz7ImcKODiz3X
NPLQjztMjP3UYJFovtWib1conS3wp2kmy/xPQgiXkeRmOna32YRTfS62UiklseNwteu+mGd2FqLS
dWKs5d0EOda0XaRBEEXLcIm4jSiCPEgCaGDjDYi+oO76DNbRCazAX91+3uopx/ym39z18jN92cGO
cihX/eLdAOlbN0zfCpBT9tFmRC3WWH/tKjB4pyLkFUCoSQpgi6p+6Ecq37nrZbsCkTvOq7SVB35B
Sd4SYoO36qllAmn3kwrF3IUcUDnLg1P67KO89K0ZpsUsc0P1BYVQE9ru4/kciUXf5XuWwEzgfHQ2
74xJt+j0v2z5oIGQqg2daeruXkScDDl2LRD3fZIAukYw6gauS7K15tepvUAXjKxQTbmknKpikkHo
6eacMwjDLcqvdjFooI0bdd++JdAIh5cIGTIKtKe4gkdMjjul6OSU1eU+gOfnjkgwqW2L94pXYy8/
cQfMCZut7YW5M9gDh2KBDiRkqTU2WRGF1OpCw+fDBXnK+x43ob271kgCYuBZm8Bo7p63lIwpzwLL
Gt/u8VCJzmzWr3GTfPvrouLVNKZk2YIyAB3c35erGNQ1zjdX1TUF+iD/0GIeFtIRe5B64Mprxzhw
mw3/3bAJDqAG/74KFxhjBqbxn2M9Ey4+bScwrAE9UQoLKmb53RACIDjFnA5cC4jkMepZIKsdRkmC
21vsVUSY9TGY0cpuCx+/BSyjF+GaLmn2ajjY9POjL+xN40CIhzR5THTGtHcwTBbc98YNRbILMmkJ
VVsK1y5UYQxLSCtkRzmGF5pC1a2dyNCluDapKgclKkVGAryiSvnCVHuiTVBdpZIFMtSpr35+z7IE
HYf0v5Nsy2ynaLlKUNbDU3RG0FlqUBMGx9w8Pw3FLv5cpsVUzOerFd9EwYZRkv+9TGW/c4TcDfOc
chLUyqYIm3qh63oW3CfSH/7SkwB9uVUgov2eXPiAZbCSrq9YWhkHdIu8fWU+DKcfImPZKksGXR43
yH8ZlFNXFPlKtNPmsIi7R+3lTpLBN1jggOjeEXWn7uoiWHlP4UxM9X/X+HyfN8DSqqC30KSh1ZX+
bPJi0deFFqsnX5RBr8k3L9BS1w/4yh88CVeKINc5Udor70D6byXKnYrybN1b+ugLTudp5S66W0wV
wGOnQiLHngm6sqWJ5Xhgd9RNumUcFG4c1rUfqpmtwUCbZV4KzQLTY/559gy7y1/MGDdT7HF5pQuF
0MXPJy8oHyeZ8ueAEs8OjpoxC/vdPvRJL0DsJgpCvfq+Eri4jnQngnq4Sx+yRl1rY5wOkrRCUO9t
Ih/vppwswU0qCQye6NpvAxP2+osaxwyltUbFBmLvKnpibizekksrUtoKCMfn0cJArrDHy7BodFo7
SPce+P3BP/dFITzUHVYADANzhFVWifWUl79Hgirvtu6F18a3z9OhkE3lwA/kFpeoWHI+BM157PsF
rk0/dKsdaU20yycWmNr8njiH/+iCOF1fx98YX//JpP05nF5vyy6UwKwAeSAs6n6wFnEvLk5XvpcQ
wKy9Sg2zRn/LplmSPKee2suOQPldYpgZ1u9o69WnTnTTEpT6XxMDzxNx/nO6xUz+YG5zoANMibgm
DnHXKXUD0OAi8l9lgHQiI2+a6QVGB2nroHr1mWpZNI0+WWoECRNda0wSKdc2r1zqEEaJY1lNuiC1
OrGaAVLilwKfqwcA7HraXSJP3GbWpYqJK693vLogKWL2pYdBm1LJ537f8dFFsNhxniVmS06G/9XC
t9SJDO++/uSttOPBOrwA1LZQiR3M0LvktUXBiVAnnEORdqZChzkbS0KPW3k82GJAcZqs//uhbIst
w30gsFgirMTPGuZIB7Y/Ys2tnwauK8nC7nmAaTP5MMPxX11GX9sc9lhr+1ZikTgeHfgr7KR4iONc
eFmWw+nezgj43nQEfhtmnUmrEzr5HM/9WVawGLxaAiR7DPDlh7eh9DXH3SuxfsxF50rrsCZqQN9l
ns+DYceZ9tfb8KprfhI8Olf+btvBem5nJAVVYZCN1Exxidcn7QP0CAdC4if+y8RD8NeOcYGVL0l8
RiMz9Kz4F946X+GcNH5/pRWSZ2E6bc6PzJX34SMceVxQdvUCBl3+8wIQkAGY1gHzp+M1pcZ7sOMP
QlUrv3trUcxkdQJ2z7iva4j6EWcbhUDavqFQ7xZsbYvqGnz3VLWz7/WQ2qj78Dl6y7L1aVDsS5jj
ZtIYpWjIcTc901NOFb9NYfJrEUgU2UfxfdoylNHKLB7X3x4kirEe9eAp4277HYD1xov+We4+kAaQ
jj46iDV/tEL4eS8GQID0NmrzbsL7ACPzXH+r0mg72xbZShIfmLuLFwZoyvXOs3dCy2TWffbXu97S
PPVdhwnzkhTZl/hMiQ2Ks6safa2ah+MPh1BRe08uijvhAiVLLG3mrWb+lQqrAAGBkSkui94TGS6R
fHimKjsnPt4e9fwLeSD698J85oOnCOP6QSDdJ9Gan+7zCPq4TNLiNGnUb6Uq/cCwsOzjzkPt/UUm
sBfJ7SItKiZz+gVbyATv0f+pytHFRW7XAGrBO0j1pcHB4sJmjCCUxhygEUKECuLxDh70xvzMIR0R
XIkA0SmJFxTBDPCNxKEJYo6dzb7Fktpg5pFAnPFebugmso/a2je8gbxOJo++g7GavCUV5BCL9qn4
xx1d1dOkmvytMvd2ij8eM3KgO07wXxgbxyoYnVSCXGx9i+fWHkZ5Wu44MbcYnyBipKkoGgKqlbzB
fMwwiC5P5JJGx/m6G3mik7uzA2QFQQxRWQ0lgrOVOhhTiiW989gdbVeGSMmkvFaX2fKD6CyXFwIY
3ANpuww3RpxZ6xKLJi/PoIlwiQ3Nd3bCE79kW51tcqa0jvFy5izjwBELcYYme11Yv774Qes8TBtk
y9WNaLuoO+QAip3vCGdJI9VWh5PPAfKC62ngSKDfylPdXPgkAkDTlF9SAbJou2VgKcsRoNSx3SwD
GjuxlsgZDS13hIy33MYRyHnpStewB7RWXxvEY9fFFvpaSKbn/vjVRAnHJzQHe2BuqGzHzp0H3FU5
1gHCay5UShTAiMr1LrBxMOmJ7CuVvrKbUmnwqYVROnRI/x8svnHVzv+VTZzy72E+BI2yWWk71FI0
4Lt3wlxUOQ9CcqhLWvDXmFuTN65hVl65j6zl5ATuok8DfuX3IKFpwNQ89vdLzVuKkBdEuNQT1YlD
nRIs39PALz6vO0gp+U8nlXwhuAUpG7RcZ5EwoNpKF3ufQV5Dg92CsYZxQkGMlyxbgR9H78rJ18KH
yZjAX189TZfDucNnDZbR24GMfzgLjK0z1g4Q/uQofkTboEIzXe+POpgI6DJz7mPWrJIQfzdpZYxU
+xh/7rAtbzXd6J+PgM3tVPISy2hkjB7710dSwFmxUGEM42a+vsHUb1OCedGZPwN6SpXfOHslKyT/
3+VPkOB5c/3R7cZ0PvBnBjNqGd8NkHhCCTew/38cdumssUfCuEHOyJF961s+NExy9jlJbb4iVLFN
BnJlY4AYntimAGut92HSIaeUY9efKez1OF0DM/WCvshSFCtAhCaQ4N9TB99GC4rv/vBymdrAcXVr
uT8DRorLW3q8sQduvuGGb0DZvCb12zHecDrWcXkd+lfc/YBvbyLKWglc6uA9Y0KWfkEF4u8gSn5p
8dB7UZqRBTq/Gfkiq/31vhUHooywRqOjaRT1W5FTyhDgo9GVeT84rn4S2hr5EQ51ph9cnsB/+nsm
8IwTm/kHzANhDykMsK+QI93Y/WfPi/WRXxKZPKfSNJcKjj+vV13RlBVXEjxbOk+WTkYHlMW8LgEF
tQUg0WRKB8oGV0LmzP+AhjTrPPhaXCNcXNZf59NdXuYLhk3oNeS3zwTfygEHDtpnxdHcry3NA2j0
gsTg9uSpWFThkxrAyAmoz/tCaLDP1pedaiI/Z9aF6Uov12SznCb76jK0IiC4cJBTFmsWexl8Nyqe
yixhe6D9EATdrlpzrg0Iu3STR+/zJTGN0VoJmHt1Sxv/Uzqympv22xAOCMqePnSVKTudKVI95PCr
dLyiNbaNDcF3eg8jZEIkdO3vrI5Yik3+c8IWyLiygcNvVL27IAZ6RBerZO92EIeW/XRHg+WF9c3T
qAqi7Og8M7RkMC+OHBY0dM3EqOMK/NoXqUJCTGeI3o9Fm50JVM6qsi4GAd1dY4FO5wAoLNxN9ed0
e7tPuDKkBGqzkSEmwOBjxRsCafu+At0HBeBVU8ly7R5zSXkX1p0aKMu8dRUG5f0y+u9TQLJ1Mh4I
25A+4tllbtrc+TP5v4JIu7C0mylfONPVov9CvYqrtb9k4r1JDHE2oIl8BwiG/sHdAiWCJXtlw7wQ
OP02M+FH0Zgvv9cIbyuAXDhfkLa3YdHS3JU2/T/7g9nIWj/aS3gg3Jiayb3nS+tKPzIepXdFnNhO
Z8eSzqv6JNs2EB2Y2uuRNTLmyO/Kz5KFbRTK3NAhloff/KWdYrf8jWgQ2HRLIdOFpCpLiQGcSaRI
i2ElDRl8GqJIne6R35kUaRF34QWXilJE+rvhyyH46RNUFHsQ4qWgswTSpOiVkl56sAhVs8Hh+4uC
W4p04CDKwrDaWctyxZtLQj4sw4LPv1LMFbYyubblKLGeQKe8I7QXIXDZnWjBaJ59lmxVspSLvD4R
AvvZpsWNRruAmgIFnoXGz2xyrpXd+dTCFMWZMf8xRb8BKSOnjjvzbBxhmh5gj6g5M4of20gBRTqm
KpZoWDLuodQ1g58HlyogKgeyv7ucpObX3E3c4W8rwPCaUFjA8HGAY8gPWHc6cGDotLYQGzhtRF2Z
YSUkHk9UKKarv0ER/nCF9fJmvmjp4zOOUTnHtktg8CTmOVd134mABLYfCKeGooKAwItREEwdVGok
Lv3EvkOdRLgBiATAfsoa6VO7bGYNUwUwAtpjtcbwrIvN364ivIj8713t0ZfbXQJlF++zAkJmHVCz
sF31DZ9Y7e9NcRdrS9Y/hafoPuW/mhF0BnCEgmOmsYpIkePXRpFvWRxycoa35JKLHLtrU39BnsGj
1hFyuuubiCbk9AjQ9TDSurbJwKtux/OVYr5QdEvG4imXm4x2DgAQM5YndtZVeJFWLK0fV0JYz/LQ
oDk9E0bN81GtJqTTxb8X+DGeocoyQkzxJHMn7gU2PkX8aeQnXFHitojmbCvXG33hTd8F7pZqplZJ
7N/hVk0+Kl71hLaPetI2D1qTOobU7u9Okol8CgbLPg4TXnCV4TPpnFDAt7KNswBdq79ug0tXPoNe
FAm+qDYS3bBLIHAZl7HGJcQv8qZ77f1e8wPzrE1jnRwVk6zsWzOLwpSmQSh5FTJU9Z4sBdOdnzNH
YB5XFVgxmMtLii8IfcfEDrKZNG4XlE8gpBg2uIsCMcJ/jyAAe5LzxENbGYTtnyT/l+BaMNZVe7MB
9BGccJ92NnvRXsU+vDUxsjhDfMbNPasz2fXqIRZ/+O5EqsFtqYs1yaIiCQJ0IA0op9iFwtJ1iKQk
oFyaevrSYDFJGbP53iLwqFTVSAq/AvWkFS+ez7JPUnzjuuHkBxGXRj8GVHhmmt7Ez+BunPstiQuH
40vuRHDrYTQM9WLvZeeMYza0BZlE6/6Vpt6K5ePkJRkxgeWOzjIcW7Yeewcy3Ml8jbCCdg855J7P
wW3LiFsOgcUlVzTOQoG0/KhxY5kBcNiZVKMxqkyId/Bjxxpd/ZO2HFyv+G2Cxi0X2fereBN4g+1g
trz5b6Z8kHqckxRbFQ/1hxTiWmnPeWwq7zb/Bs1vg34SgqoceDjzqihHBBysRxH/2Ol8hgpzAgSz
cIJqA2Bq3tBw1cd21waHHyaVoYQ/7moyPgyAvRyBaZQoH64K10mWzxizTq2xrRo3caOr5le6P2rx
ePS6DdZfiG8ZJ+Km5bgcuJe16J85HhkhO0rrVGH+BZXpKn4leA6IxiSvKmIVGuzQ9ro/kzxkbthT
RqMlxNSKtwaorisWgUoQl7UfEs07vDAaApRAaTQD0IHqEzWpOWRxNlaM+vDlS/qp7dNpsax0pz4e
9i8JhNvRj37xZn5ymt+2ZDBCTaaTW4icAJE1+jNxaXTPIT5g7wYWmVb4ivtV2WZ9KCRaXoOt9VA1
hfrYG79coD5OmcCCyupBEUG2OL5+P+YlmyaXwC0pV7Kv/i2jVyDHjQwga9XC8NzGTAURBdzJr3/6
ktj9oUawE6l2Ue43M5KAIiufbJfSui4RBtYVF8qE3NJSmsZY0algPWcqm/kJA5lgKPZRHzIX2/f0
BSpHqOHQgWbi8ub28vpL1gMqxbcx3SuWMm9c2Mth34RsJHKAy4IOnVFUnr9G67uG+2lJnFVEpzax
P3W8a+bOCRZaY7WQiDnL02w+OaSLaml6/0q4icGGUSs1YRZxvewVpPnakSBp/WwI09SDr3o1N1p+
j/BFFbsaNpJhTJzJHoKk475l+8Ktk3o4HPkcW/G5698SsyiHqgZpExlnLxh/72NcPXXNdSXjLtZW
iMICcx3UTzCFk+rRQXcrYuAjU9S0K92wSI+GXgPEdXWk3qSXdrt0tLYp4LV3GxL7lvA6wHcLG6Ob
qQP7rEtN01NMZiAX98qDPBiO0ebkHz4kIrasmo4t2gPTVhzN0hvWZNxK3FoAFd3DSZn5fOUhXE11
zIu/BM5lAT3ig6+zxPi7UU1mY6sS9OsvI3lbPbxFY1PEjzjBYMySUy8+8ZqJ0wCUQi7fSOGnfpH8
Y57tNQVW674OOMNyZwiyYcKgRYut4sM7nNZZyvWV1YdjffV9fK5UmfuLQyiAWkPverIiNrC1xRyK
ABFpaGE019wuc+1Rfs09M3qO/XBS+TkAA2q/gz4G4GgNJsv9KuSx6a3kwzxVzPlOj9I1rGU3XyEz
uE+jEg3HJ2oQUxyxRYfIlP6lE1RSa8Zt4WRxxVnhbfnh95AMWvUwqyZQlltvqExFJIYki8rYnJ2A
5TM0XBVUsq/ZwbpZ8pOVUzgOCsjBT+MDgXeFFgVvEX5Uh0xUXiU8I5TNcmWjto5vY2A3OIg211e+
TKsn8pnfUSwYtH8PM+uCCu1xr7IHM4Vcf+uRF1n/zmlO/y2BjfcA1T6WTlyGSxpiytkwfvBABdMl
lAQgUHWliyYhwr9oFAgtTLCy3gohmP6UVWbOqJgP9AMyrYTDJYQT4p2TjCpyyrlCs/tifAeLce+U
HPJifpZKSxpvQqnx1SzGoMJ6WrLpenovVJvqSFp/qa+3GevIXURNO40uNyJXLtvmZvQ2WcskMT/G
Hy9jhqTFy0jppfrUMdxJf37V7jlgWH89845fTNgogkV79aWfwoJyzb2Mup5TuVFp3EpXj/weVW2Z
p7mH8Dk2DzFghgO7/4PxeDrYzazTTf+mGLqEshgKH51ZG835t55wR9Ligq16yk67mouFJh3GmDSa
/gCX/8QIILr2YwXsNR1Jmi2KIRjzuU1nHZYbLXKD4hnyHFtOwLFytG3xq9b30ps8ldVZRoVtXibP
fZ9p8+nrZbvk7T4rtsYOj7/T4f4eI5f4P+9ekZU+zXgm2Osm/LoaP41OqsKFwi5+cfIp7p6WolbC
EfZdXST2ejqDprTWg+9dy0bLPt0hMuD+MiWRquIJRwlsz6NsxiHD/JXXJppKyz1hWhEcN0581uBt
bBM0rgKTo0I+4aERcF/aiuIojcQXQZnyT9RAfIy06Mj0J2BgNyjy1ZxO9zkZeCiF2SXwpNfzFgtb
O9Wf5sj4jzTwFVYXSZleR5d+YdaceL8atXFkP8K/UPv2j67YO+ip0SYLgK+1QnUAhr3/TcCCZM1p
Iy6hQ1N6w+rhCW+TdG94z0Z5m/Irh279dA7Agn1UJBqBBAWpCfwTRcKSHhUyTbZbdkjwY04yaKPv
0oub2TnF196W70AWqteiVd0MnpAnIY1vdmJg8VUY32Rqxnxtoo+RGf5thQ073Db/xs9SSQx7lM5N
2CMwmr4vLIgzANJ0tNmCKUo3KJKiwmaRWCA4Z3IBR3pUBIrGVFIbSo0jCAmYpYiVyLTzvZ/0R4lO
xOGgGJWHTbvXMMy/xeKrzlgH65jOTnCBQplXqqAqT88ezFSuRb4HIYdr1rVUC6KYQxPAVXd1BxiE
rHENod6j7q+5UaIxw/KVlvw+Gun9nzTACacmRURHxSB6t9H/hX6muzqt8r3ndPnXi7OhE/7muXA2
tG6M4j2oRcZTf3Paa74D7c2uDl4Lirv9rTyj9PloTAh9IoroZj+WnFihDTKiMACchewIcwp04qja
acGq1KhJ32Nicygh8SfjrQVSEZ5O6ZnuY3BZft5ed0FZntiubV2qUfS6glr8CXt3VihSTyFbxBtG
h14h1YW240J17tbwGtUwckmNEc+f1z0YGGB1sSCWZLD3Hm4Y83J+jBupEXVDM2d0LiN8qIzUzaL6
L/sLTWRRe6y/suVrBy/KxleNjedBd4z3K8rt995hUzL7PKPsFagHedosmYWOIds74P5/KQCnhPL/
D9A7oQdHPgnHnjesvW40GEbNDxKp3gHmcu3y5gxul0IkO7FapRn1Rk9jatcik+KAItUWB+5xrpBm
0bLCRTbKtEGuDhEmjdScgrTwVIDQrzCEy3Q1yUtnN97jU/3kO/dkB87dJvdHLJl+XcTB/a0Nrhid
FirIhQvemBJA7AlZFMOeyTHRlK7QW+Knh1ylFqeImWVQTogJPkhzQH8VUjQ+tnyPaHqq8hlGXxTx
f411GOLntC3DPR10E1SxW1DyrFwrpydWQWrxHrsMHraepSKmfZ4UuKDwec/4EzCLEExKhyT1m51I
S1Wjxcu2EH7VBXCVKQ7GswR7zlBcIGUemKc6HRGUDOgh7RHJCTmuCGlyTVOWoxX2Wzt/NDdVXRsp
6LRl0Yd9e08NQDNvPZBevLWQpruXVIWF/xdwTXIJBjpSYA3EIefu+H6g+bs7B3SuUCf+4olZZmjh
cmgwQ3WOuDZYMUBeMxFhTx6l9naR/KSrP2m3wR54UyXa0/7XCO87DlIEeGR4b87TRUQDpIElCUyQ
Kd9QlMZemkmkxQ0bHf0R+NsiPqC6dsbLwX3iw44S8+fkc9Orwn954IWannsv9w5/QE/5CAf0KNUe
AI6eGTy8BLxwTSW2xxVzGsyyPTKsCWlwTVfVHXheSkdoT/q2Vhtpd6CH3vYR/EjK425Ajo/lx9sr
kCghTrfO0Dv1hrPNMNYLZA9ZaRL513qiT0ijL4sAMI8E2+KCx7VDoDXUxEPe2+fMNddfkN2BOo59
tacPBaw8YdXiJTsiTVqjl5JeUFG0Cf5o1FarQwuddguBHRSQCRmI6/BnS4PnOpcAEKewYasZmg93
37sN4s4VxHGE3ayN13z4jIbrPhwA6S9pigDQYC1MOINtLQMfR78kw11kD5UTOxcSccQ+HPeaGeIt
yzwk0Y3oc/+LdCKp84s8i/bo/UG1QaJcxgGzlDpTbbPDyoACzxC5iLyJSEGm0lo+4oDO6Zfj5lHu
CzKm9CyrkYzMxJA9K+XIog1QDEbZThgUQt7Kps4jYOPzEcLuT9GcFnMVNyYcS7QSyp12bY0+iior
XABbmraNZvn4omTRSMruq4rYE6trPxU1q/K0gFNB6wDVJC/reBlh/3H/r2hVoyx0+Gh5/SaGQGS2
O2nPX0hrPMCr4YdywdzcrKevxtGCNXrRujYqbJfYudRoJj18ogRcABIAB1q1dql737+CTsh9HjOc
0LBYfJ+X5UCfZKubxspIc/fE3yVXqY+b5PZAbPyX4s01GQZo/KBXWpWDDN84J/SuB0lIndX2N/Vs
r5yCRd8jIju0hiwDZlxvyJzaR1f185Niq4t9Uk2QnfKmAzX7ruKerjd573qRPHR0eS0SMaT/PhFJ
2sKEZ1rGf+S1HJeP0gxWeIuJQGyfRB/E6H/2aLikHcujrQauoQNb6tPOEeo89bFQqgOqH+/4mnWq
tmm6kD6EuKaEoK3x+5D1UtciIExVwzT7J3T1A0lBSXqJO/2t4M6ktNSnHvE2N0ZZPfNyi1jN4cMe
Ap2s8syp8jRe/jplo4Kvc1T621FRTYfrJIkoag39uvD6bJKJ4KYCrUdIhgnlzWVJcszxLfueA2oC
Zt8NvN98OXUISPvaX2HyK/vOgQYz5vokvG3/eUBNe2FfJpl+KO9GrzKB5IfZsJfJ084yFMCLsSbH
4ii9b/3LYR1R6XdimDvmzEL0qj617A8+l+6Z1QiOU2tgYach1OH5MLPL6garmNg7gQJQbXY2hucG
s9G3gIqp76mMrMVnT6k1W3sBIJVDShTYh72QNe0JspTx9jrbU9XHKWlTClfWSd+W7ivHDIjMWX8y
VQnecqJBtawNFgQCpcR0QI/vAT5hsEF3wHIZeAwACod9EzVV1C0Wat5yXEdtZWht9XCCSeT1EnrW
j1rMawLcY5cwWV0kKRyHqXTAogLllDjl6fHuEtVt7wcpyX9MOnqPX0L87spUbVJnfDkW3SUSsTha
mp5kLHuUKKf5aQVfOs53RkHR2sMDQ2zGaXbm9ArLZIR/r7FtrqbZXyZbplQeTNjY50ueIa75imIs
VwrovvRk/6mrEgCfgCJZZQb2vLNC6mC37ApIIM01WraUYorNWPYUJ6aY+4q203YduVdyNXtgYygi
IT2VCUB7XZKnsaKVKug9VMz6YWpEWQxbE3kN1Y9qDMSpGK+ZT4FQDSudDqtwFZhUXF1LH83AutIG
4amkC1ifMWarbSHhQiEXQZyj42ERFs7xboS2I1IaoKwAzyB5QkEiq6GxkC38SHyH0/AQH6sbACvz
tvek3+XB9Iq6k28vTUdKvIzwO9dVyqniFX5l4rHQIlR5qqi1tJq5BHbBkZ31Yg/VF+TCS7lBGGDK
Nf0QRQPk1MPaq2xxnlS36JsOdVaqodF9xc9tlRUOj458CV8pOIz7KpIGkMEspTk7V9WImf7VTunv
jx3kZcpyu/m+Ft+RmthNdALP2Eso1i14fctN5OWza+a09DMcNGr/zSNs/LEwVx5rxSY9AJO1zvtV
M2lSD0yGKQZlLtpWbIZlN000OzvUJAzSVxW+KyrJuAcvMLd0dWzmJF3uSjCOhps+hlUcJPXuMqVJ
QYw81QCMhCNhlU4Xos06kLioNiE/tHRPw+4R2BC4q9BfIlWqX/GjaC6JYp2fGIhJI/s5lbL6Gft0
Go0I7jXSU1rI34vY99inXrUoOkzYgQlOwL94QY13yCqtvEa60Tadj7eqLE5PyvnnmUdm8iZhT9WN
LidsrrZgTHYrly/2ogzTi2L7cS0iKatd/9QT7jWr36pwHP8HBLm5waQpl/DbaoM6FTAWF4WgznY7
9/16V/89+SEuSz3or76Qv+uohXK9WRUfX0kxI85syvvkEdSD1VLaEZuPPeuCHfkFE9qUgg/lc3ll
BC/ChaIA5IZ9Sp7qWQNEAruO54Cp/vzZ4+rclR8+mSISlq2IhEHwUvLpOSfQdUPclKPkbF7sfddE
Q3BXovEo8g/+QXl8/v6Iq0t8IS6ExdNwCBbJUNg87XuGzu1skwGKrlOiwjlNMVmgZZl3q92PPeEy
INgsmLX0fbfiv2gunH5fIUGy+Ie15bN9GPjznpgKL5LmRVnR2tpCxpJr0kNf+i8btq/T/vmZgvin
bdzI3o1IKXNLFxU1pEELcxOyg7kzPs8y8pX18z8hGFXxlE0t7zlOMwExVECYFp40ZPaJk2eDpGEm
mBSuNbvcWoh1Lyb5fWyddQJH7AdcqKJYB9OPT6uPgvLQuB5J6VGKeLty3EHC/2gt0rMkKeLrPqXV
eihEzWkEcn6hU98NzEP4PPIIsgUyt8VKKl2dBlNZtU3ibvaOQ/Q4fWriTQYXboXdiTH4+tpT0B7M
y53oszFczOk/gxfWHqzpRlLtDSni/6dEkiBABtDrqz4bAZRc4m+24Nv+dv+bnKIwt0v9vjF3C+gF
tQYdELqEXUFHava1dqO1cugGywWr5hVpc9KYRg1eU+YV3PrT28hAdac0yc630NEBYhlo5/KLt4uv
amRn6bOX+oo41RrfGlLRlKH9VmUSVmRsB3q1291zSANn8oDptUgNwksJfC8oEqdEBk3F39eOu17z
Bn88m6rhGQq6gnkoZVTuOcHHlKNE9Tpa44ye+xy5yYmc2l8gicdfecozzux0aFr+WxhkR3OBNYqQ
Cecg+qvZZTFyFuy3uQyr/iQAgNf2tHf9a7C2hrmyu5+IQo7MlojWKLsfYepGLZZcjJR5CHLEd3Lt
vvZGEo97XkQbMF7e4tGnHvw0U/3yxcI83v1GtOWoKSVt+nr9fplj2vlZ4fv7D64aHoG4q4sEEfPK
7bnlHT/+2sQOZ2umP3bAG++Px5zJAca8QKYwYSi5HMeym+TcpAGj1qb+ixTuIh0jcw3xzn7Q7zHk
tq8lS+gYt2lZUJpDczHqzdS4SS4ev8VaBKp4l4F1k574ULn1AjL55y7RxulVgQTz7iPVYYDvtW9t
yOcZCAw5GYNsktkuZ2lxRMhvHXpSDf6qjXak17gvjSKbEGFXOJymxEv++u4+A8AYN+GlHmRlOITW
31sIsbS+Jvkqrehc9OMfvu5IFxcUDxDmp/hCr/GBoz9qQ4kv3xzQebG/EEY+uUV1eKWraPnMSjGG
p6UwIcavLgNNXx5qaeCtfKvhSB3B1extyNAUEOMfJUEphFbaouDMF++fpANgFsogZDz7BRciXRBd
GmMCmN8JcaE3krG6eBFv6wINiNftSnVvzCJO71vigYezXnj3KjOrPWDzCLEGhcwWUNmqsNnBq83x
aoOc1JIJ0sAGvnc/oz838euGRDodofDyZZunVYyilYZGxzQaZaPTkHlZkzSgnJApBwQ2MKJeA5Sj
AufkEe4WFZVosQnmtBm957RRbt6qwcB9NYE8lArld7sSFZXu13fg210LseXfhA/3X3NaZNcT7h/k
JDAIKQxy1TqCvRuhIDxGwAWCh5e8nb1tPN00Bz5RBrb7/zSlcbcWhpei2CecKB2qtJv8blk6YyGi
hF6mY4J4Ef+Suh3MCs9x/nR+I0mEiGOi+DOfSXluZ5CZQaip2GCezf3KtioA30b97nPD14Jfm4+a
CWxFvawgyqoutW5SfCQwTA+DY/z9WPEi1TNFvdZwYiGy32X7e5xNsCOGKjAvtVBKUCaJzlxarpOy
jIDMBWL5czuQm/LVjibcTsJeGEK/0352N3Ljk1niIbdxREcMb9wCNCpMmAAuwpFk54OYiWSEeZAh
q50gmNSxmgalZbrY6D+IXK6dw6N0BIlAnqMv7UAY/glaQBzyqCupgplxwchPEsl29CJ7MFVQfudR
wGeh5ncOhq4KMSwMhZVh8FGTadLP6MqzSqvWHlErXJ6D9x2TggGwCT4FrpbsyOJvYm/Ca5Df8X9J
JznDANzsnRniEQF8StOPUMTTkPDLutNLJiKDWcqmeDb2W0VJyOhkG5a6aByK3Weda0C6hvI1/leS
qDuQ4b3f/3nXHr8rsaCqPAfJUeZI4EcodqNsTIZNCINIwmBcf9ePqFZIbWIkTE9sWVN0bzmf8Dzf
G4zkyD0BCUx0Qff7LeuGOY4aphzYmr3pXpal3vU/75avQpp7gKmy0BmnoQLEQui2D9HkKkeDcnWu
XSv2OXsE8rVW29xipsmfPaznbFLV14WDJ8UalEO7qVJ3Ymk3rwIAoqV2QZ/sD+NgyUrXLV+70Zmt
+KUYeGZuZ9dCqQC4ROFMdugr6Ux26FArAlrpuiaHojT0FCx2uw4skZNuCx8KvUMW2rX1gStTn3Rm
ajJPqHbXWqQZ8zzuP44EhQBBPDIdvKa7b6wr1kjmQh/xWEqWzCYLb9inRbXZP/8v9WdZPYYh8gwn
4x7e3JGh90ETtQL/ndPWzzw0OJv0CvhYvh/sgRczGPSqBYKMgNwCvTLzAX4LOAwACV6W71st8aE3
4GCU/4u76QAhRlEhkw0KfC2U47caLPF/gSGiJ2RF19XFAAxhLtcWmuUKe+EkoOXP6Pt24Lo3zZBs
AdqBHjQa41CMCU1joVI9M3k4KRcwxwZHCawgQP/BityBxuSLV6WgkddYCOzJcWNZZ5xOgo9BLnkJ
sMxflajzGvm1l8FXOOM6ty8VZvB4p2ChizsQiu8xIZPOuwESPQhvBdtFoPshuh8PTvfZmILY2FTX
gj70QtHFsYHdUkABFlGsvVYQl+ax+hE0xvjH0OY3nkrt47x5lkCUusp89vGJiX74zxzXwWj/M1Rl
cDenBzmJZ9g2YgnnCICY4+yOPOXRjRPajRN9iVzlZshA8DXrDvbTt7CDNWCBHaiRaDx204O+kK52
1+1O7Il3EpFHh/uI2GEoypmMeD/lc6oXtCIg5ISrxQtjMPXjCMersP++QO9SSy/kufSaQbBthLV4
4nz4q08HKfSdiBzbELj/FTdqRPgTSiDK9V5jaOQiscKYNrU+nn16jyKHcaQ2enmxe0I6Zzxvav/H
BRZXEvEI+h1JgDks5Bkwfy9hAan4yI/dUqKhxEWc2YQBufrtNC4FMCV6HE/iIVHbUjDYhZxJ5ZNP
9QVECfrBZmTM8CPOTTq4Owjsr12Ohds81NJwMTVfhbUz6QgTOeBfpyF5zP3rBLmPQ9zjOro+Hcaz
fZGKakZ4tGWX/wLeDPkbS8wzaZZbKsW+vbEygzRymskhAqJZ1p/RLVHK4WdsYbnb2VBJQ7AxuNi5
CnQxJqn5S9yj1CyeVMaM69DuX8gBbXKkN1Y75RfPV/xbUio9GFQAgxtvnfPOoMpj3X4mu/O2u/ch
Bt6Px8xCgQywB06owoqKq4TquMmosw24oPWhRIfbwr6/w6QLKOlY7K+717kku9jmmCud2vjzU0zG
gsmHUuU2DVy2FLTkdx80c74jN62jhBVJ570RfuWCFV0mcTQHRfpvd8gJgoyB0au10c3rHVOEpeBM
0A8MOZ2VM2+gBn/hExFME2Zd8rfxlUCC9Mrg24QfTfwetlxMbDomElacQWuM594EulDVzb42py4E
ZBx+utjtrlVcbjQ/1DkKhlmePLj5FMFouJfMcKqxPcQMDvQEa2Ff5W0qgbgvj0TVKgdX8kLIXay9
UiW0s2R4ZDXnomTqPGheemfdMnQgtVCG9BrnIRr+i1KgDxWqNOyHibenRCvBZjs82MZE92i0NomY
tUaj2g2es7s5I+pnlwR3mVgjg4CcQ7tT9m0YxhE2DeTADCzcvQaAyaemVhg3mDxmXVS5MwLgLlal
oTPAr+LvNvBugIlH2hPA3dJETJvpdRoRqTjJI0mMXz1VXzfKZXuquY8Vh7rD4v0ZnvWGCf4Cwwy6
JrMXtrcaXCL2/R6OO4jhIKXpUF8SupPSkwCZMEuYq0EHUqrFfTu4yPGDpOThJyzzJy6+6N4LPbqB
meTNAtuAQk87ix8alIacW4MFVKKux8CRAUDH0pWd92YlXSeH4Jd/VciHe26aXbFcMrR1GdUvE5ox
oI86Gty8amVzxts5yv+adG6kPMjK8jDru2EZqmx+DTGZS8GG67OlMGhmMdm48TXsgRbRwQ2EGtkm
piBvzGq7Tb5X/Pc+qv+NboH15tBxgvRxHPRFrIqELgMtVkpsdbTkgod2LRNAfcjvzsPwD8EO4+n8
Bza76TEVtSoxz+d/YhpPRgwtY+bTosoXfCKg6beiZDZaa6QmmAXkVY/h2tpseD6eXgw8pZdiFIbp
HYpoBZS7UI3o2Efu+bZBfJkON+Y9SEi7MIY300qxknrEj6se3JD1GkV/NbwGUZUkOhH63GN478zo
p2ugriAXrewYx8N4QXiUhrQTqzVMapjkCU7DdLvC6PxvqFI8yhMG/DwZzhd9zLVPfIRpBk6wcxju
UrLgXROCVgQ/dPKUdAzZO4bQMcySA83cgZUymxbfYEfrC9vg1YsrfnNyj6Aas6M01btAMbF5iliz
UGSg9JZVurmrQ2sLYi4Ob/xFf622lWCxh7Epab9DZYdhuJqFbsEO14ao+U1GCaBbIMij2WoEQDni
RqYDmhfby8+iUhVuHRHzoHkKzD0AU5c+UofrFIDAyGQyryeQI6AjQMP/zsu/W24hrNiTbF7qX6jo
Mok6gMhELc+2OVJz9ETWuhZ3y/q7qmVoolrmFbF28qvdoiV5BSgm6nLxynSy2IX1592nxJerPUFv
M8VhYbCVhh2DPTMYEvD8OhGUAe2as07/36nm+OUyOeXEKYR/j/ehN2Rmt4XncItea9KueY8cc7lH
IkXT1Qk3pi2QgO3VjGLrxa6j/gvif5CLycsFKg7Vmvq4SBp5VJPdN8zLKVpXKyM1tvYlxAcmW/ru
bwGZE9GkhKmd8yEnUqE00ulO1nJuDrYYckyhw9Gus8zBY8Zf9UsGY2lJ1N4akDM7KnYQE8HA6koB
KoLSf8TGCLlr6ALpOQsGz/kgOPNkv2QK738iVzD78ZHMDbTTzBqxE+fPk4cXn1utvM202ZMUwE/0
I2BYXGcz+lMbNWKtUVWL2sbHc8v3BHswQNeErIGdog7CXLmxhisVD+fEe0/VajI1d0lp0wlqL5mG
Ss7yv0qWXGy6M3aMtazYUQczbNg05hrs6/p7U9J3NBxogBRhytvZmN9iL2WhTL3ULg4yHfu01pri
MH4zfdLNAnwLS9XjS9b+DGRB06WkNy6FRZ+VUF6vRGU+q0RHrz2hBKFcpb5uRMdfeccZTtQYJuCy
rN7sVqvKW8MxlK4NhG8V1sj5h9e2egxNiyJXYlYmbOpONtsvc2V5JIDcPBMVj9/rNAKeeEqzbjrg
PMKkKLLA/luUS9uxFzYCvSA92fylG6NsUD+WdD/Xv5z5L59MyMg+RIzSMIO+xWb3THpm+ihrV0aC
y7G6hd0LK8O410OJVYY62OyAKGyfiwzw0w3VTxq8ESLizDCmAr7/ldXer0DKJtSlRDSPXrjaWqTD
DVJHz2P6Jo685ccQSae91Ed/sfP3YxjJIefYZ+ZAvhQLXl7+/Wzi2IMnGA12+EZs4l558samZM5w
GJeF0//0i4RagZve9DogWh8UkXt4pF1pF9r/cYaMY2fwZB9ln7wwMWDtta4O+y+4qYu9GNHLL77M
8p3e/59pY9HdBc3NuG2bEYuqtVFop+U83h3aRfTfMVb8QEveRoVmGluDSNRRRPRQOf/witryITwA
yCqEdW1oHnckus6uHOtx6+fJcAZCklBx8Di9l7IeQJjeowcvV1je/paboB/2LzFgfe3TXTD/DFq7
6RbIHSZsPtqDBor5Q++vVN8jCklN9k2nvNjl7WW1f/6DToQEkDYDBiz82lRjKNJhsUlFGkdCSf9A
mS5/2W29CzP1BATg7FzGbEwlsx8+eUD4D1g+cNwZ9VThnAKpvXklHJTeDc6pQCqT5HP1VjxcS8Io
vjrOdGMFB7Q+k5U1S2/WqKnezlXMkNG12T1Ri3r9wPNv8CmGSBcX1lSOqYw85qnPkD2Z/W24scEY
UceoZCRTFsXqUc7ApMqyNzDwaBnoGAgmrgcVCyBWw8oe0/Y6kuYqBdBcbuSTL5pJfBHkuUyTn0Gj
EUd1UQz8UGMu+C/bt76ad7c0SfJQYoI09HdQCnkuNGzktjhijdfr+aL11WCog92DKa5P8cbG7gpg
Aha9Ik+b8uhDlxQr+8KOFCIo4pqWWnMjH2196Ypx7g5bB83ZEeXfxvxi0skh9CfRr8g4OOEpk6s3
ePxzWofBFwXtM8yzpn4hMV2w1pTiopGbEQqfdsZBRatjV040wBGP0gY68XCP20UHPqDkBFdDeo/4
2Ur3i92hJ4YVdjn7WBB1Yn1FAYOgEMMXAlnIqAy8FbyHAg60u+a7qJTVYFv6YNlcZsbUoD1MOHKS
fl0i18t36evA3eBkh1+1Iis8K+frVlh41UjzDeqbPIplLjmLpJPYMhrdOtsFFZUTZfOEin58o7Yt
CfC5/wir14LAWdKZID+wEwpGyEG59Z8wpUry1KTxEj+ecIO76h4iuuvRcbYLH5V09gn/DgtlosLU
te3sZ4gptOAP0l4IT+FtopaCTtkRQZDkY7K8Ws4A0XRiy37OD3BvzAPi9dIEoZNoFz38Vtk8SULa
mZk6g2YWB7G9mtHsHN/rLTwJXnmH+/Bl2+cH26t45zMGpXvHVHbWkwU9G0wo0N2ZRtbi33mUZa87
cGYNCUK9StEvecweNUtrr67/cl5OL7JBLwONBNMV1OGs8tLqavwspsI2bBgBD4pXT9aGPVAQbTWi
ierk4xNyO5o3oMRFsCAbozSEQU8hukpcrIKP0DSQ35Ij2ELRCdry2lZT6FVkfZG9ShlRydyWI5mC
soqzb0uqildQDhgHDD8AftOrM5Z0tTEQn22GKtkYXHFuOv42GCogHwwqfR1nTRpwf7crYV1OY/ea
kuCjrAGXir0laGWGaC+lSNJTfXuAwAfWTAu0NgFNMjbyKue8QyOLtzCOyz2fbVUHrjGUVGw6ltv7
MxYAbU5HgFwHO9LhvtkztDYod4K53UrbLVM6Xq+yp8MkGkRzKVBI7x/KoHHsSV7rNdmwbJeDNO+C
U5RuubxYmM0zyHGQEPzePBXw2eg1nXI2RKieZ4u96NnIo4LGYrwshiigIUYq86plfCMlu+ATKaNL
tH0r2PHH10lbf7mATB8oWqcyiXUA+M+6/wKah+u+G88rtBY272xineRCS0zQueT204IteS8Wi3yF
5CHYekBHilOvzH5PuzSQJ74DT6UDGWhxx1w+UM5JNNJWosTEOzU3QddfLneUSgrI2TlTGPG+N4fu
DVrnFV0QyvG6oYa/ZAVao3TWXN5SXN9csoOwMdLjX1VXVsiUBuCPj+wpljbz6h5ORAeusQsp06/r
WznjPSru1hvSEJAp0I2+F5JNzdOtYtfa/c5OuM5UR71e7OO8PEnmTEyB4Rm1S4YPDqULGSHr1vBZ
6+KPTAOoWSVwLwPPy3hSSqMtkDElpMsg0Epxo5i/wZ+N/CGxXmAbB7XEcqONyI8ioT8LFBo+IUFb
ClbUAlQ8NAhu/qTISLwT6uFgwdab1TrLCflzpOk8zMtIYWHcEzI9mf6LTOvCpIdpI9wS68Htq3Vh
6MPPmV3B71Qv+oWgLUdur1ekatrK4uZNQf6cuHvd3DwJ2AnSO/XcWwNHSA0/Id6tdrCzeRQF1FRb
n94C4H4NGRG6fMSGzvX8YTNKuw+9IBqHMQ6lcj9q2pjjfkbbYtxhuJeWi2b2IfyAuNjYFpt+/tYS
DMN+eJVsXZxwdOSBw/OOLN+8kn+5Xdd+L010sNTvcmc+SZrlGKPuCcmeloKWiLp6KN4ZxxO6JJ83
Ei03k48YBbEpEdtm5sG4FsseEi8bwMxDfOr1rZ79zlNDCr1SzeiwWlx0eWf70/9UGgw6tqwRwb06
g0NhIbDJyD1MWs8MMLOowzgeXPAltKSy6+5cjU/GgLaaSyWoLPBPQgZ0Pdx46Cp9Zzbgv9733lYi
I3clEaG0a16yy9/mAwX0UTXwBZaKj5AB5wWU6jKK5HoPO2jgk/TCWgOteSLQeI9Z8B2uSn8zhKFr
r0M3+Om+vryHcBCL/143twy7oBKfJuuIZDTlsAqaKRWrhw9zsEgeLDZVJ67SLryE3IgncP7adNMp
GNztLd9hEl9ZTsU5pTDgrhtnmvcp2ia2DDlw9E/0OSpHp8JnXMyPLX5lw8EwlncmkQTBGREMeOtP
VdW8p5S2ARMx2RKExMP5scVxbL6ybX1GnXTVBzuS96jcH6KBx5AdR+B+fY29lekIhS6NTdxFCCig
bgs7fTa9Dl0wqW+B3mXsrZqQJGzCxGi1EkSet+v1HGXg1muDpelJqibGeWYNvZ8iyk7dGSsXq9Av
0cf0MykewfpDQ5Tmxy2oo20l8NZ08AvcTmmGxcVdwda4nXG4G64eUAfzP9YXT9X/s4CPFIX42Z0c
EpQdvzvaxe8GGZYXq98bQ+xvn3UCmLFhJcQQQHTiTz8mJV+WaO8D3Px3WWYfydyNR/HUeULTUJSZ
hJw3MpX5FC8kWOR9yah90iTtMBOnTJ36Rc+BSZlBluGayx7LtEb5tQPcGMyvMa1HLG1Fxsy9ExL4
HlctEhFn1n4bzk6ouDVrhZllVq6MtCj6D8SNk9pDe4rJbbipUXNbeGmP38If1yhyJNCcx2VeKPGw
GHdoZ9L589AQqZAsFxehk7imcdBJlTEt+fQ9gSfvEgvgtoLLQ4yfRPWUZjVONjEVwrOwnZaMsFLo
ILEmng8zxvHE6bMEcoxotgvHLyR+aUl5Rd5e8SzYfZmv6ugRrZdlZLqWesf66JsrOQ750pa2Nyrg
Lfcjzsk2TrRTyg4IspjuIvh+nu3xZ08Cm6G5ntZA4z459B3T15+7RU+5CwYAwPyMpx8Yn4TEo0yu
inWTElplSnt678GeP274+NybYcVgrFfijq3gwtWsgb2Ji7UyfrKbp6mH11IKQJYOhZXotGANqlNz
EcOYdpS5s89uhhVrJo0Co3maaYSE36nSYZ/C750rH1KFqvQlHUzkJNvBFaFFV/OaisMFGSSJAc4a
oregtppmB/BpF9n+o4BINolXPAkG+bG6B51yiK/+VYC/+k+U2jGn9FlfBWZWEouS2dg7fWmhIbf3
ri/Uhoju+MEf4jJWpJ8821IL0vc8V1+RQfHmp96jXBqagjd6aHbwB2rIbW45fk7qy3wZCEwwYyMt
TgR+5T/qpW3a9g0lTDzd2hFSSIbjS/EEP6BaHyJkbY/Cwn9JuWN4jgEx+bylWvHODpTULwW8yMpG
L6TBnbWucN0/6iTeQBbv+3KdJtJoKPrZTa7mFrGwfzOuzwzJIPpNguplORYa9JqQKVdrZSEkaIYc
wskUhRDcx87NIs/JzA0eeRCxl9xoMFB7i5xrDr2yk1xRKEfyOiaGmdKnxhlJ0wdEohHaYZ0Q7OaG
Z1XpuHlOP9JFbPc7RnqIDjM4DDapo0DCP2OqnvVzOpt2cUoZbzoCdfOE1LDktvRfKa3GANHJhu0U
hLAZK9e24LZEmuJJmwPIUEeG9tI9Kgfg6LfdbaXEqlSuS5uKVshDRRWbh46fo/+1LRAHXw2EaURI
ZoFOGBzDK6nw4TXNnvgHfjaWYqsnA77m6ol/hdAZt3wMrySphr5aXmSX17b9b2l/HiItW4N9GgIs
T1IycEkLlpGndJBmW5eOFPjgrVxe0ca2md6Uq3++LTCSR/BTzZLL8bU903vcs2eEdwVRHs8C6ieO
QTIh8NB1JYocycnLlLKNmxsz3Jy2ljJR0Zbn6xRsPzoW0nIuwrJZwiAVAI091tNyxzFek2oTI0hr
GOlIF0OZD8ibuA2/b4nT4B/geOeOIXtnEg7zxKEQhFunXrX6/C/n4hR2ORSUBOLj3CfRS64bA3tt
JLiQUVmgM7AvgwrWBjaG6PfXdvxZHNkdSaZRqTbKEEnKZvgSkSTXJrxokZul7FBC5rQ4OeP4OTlM
6P6dC5fTJ+11WKgPnk1VIO21HSXHD/XGqXZFdk+WD1Z3PJg7sEz9y75ehJib7O+LlHQSa94PUVDv
ZnMFtVy1sU+puUgwSqnf6+OLy401PZX1D9nLJbDAgX71dmynCcWeioVpVKIL30iGzd2/6rxu3TxA
FlnnXc5jsheyLTb+Jqf1XeQditKDZ4Jutyd9qSK5/xcid3Jt+xqEJJKMuKTr9U5O0Tp8sY6PS11T
KqW54ysygSf9lX46mvBSRCxuyseEOsZc3dL17sMzyJRo51EpIHUewZ05ZFgBOhnKulNMt9rTShyT
TYIXbx6PRTZbWs1Yg+bsxCaVHmlT2UAFaR20FKrvQubJPILLRZSsDVUIGOiIgxopXUlGHxrZmmpz
VgGmyGrcZsutvSXZXSEOOcA3QqMnNKDj0QQQQ77M8WUtASVli82hp4qEJJP5yYL01WFOFnSOZtmk
8heWHBMAac19EeGmpv/7umWa195t9/4vgsmcFwWek2t34JiAYGIPMjCMy6yxpTICCIQF3wXduHAA
v9aezptWIs8LZ2naBn/oAq2X16q4TyCqbWHi9io/dwI5T6BKPqqVhc76crMZxgCiIXCViSvsJt0B
6FMtW3cZFxNUbGr4fSQlQ5ozH/68ykuoeoOeqvyYm6uQMt2jHKpjZrb15htl7IBH2FbKNIFPLPgi
3uj7LbirWdy5gBtP8/qV4KK7+TydyIRwNTWGSWIqRoXp306aghnDxh+UipelFy7vTyGLq3ijXD5P
p/tpt0lxW43sUljZKEY7UHTkYGUkTMTtDpcesExpWRgsu255hrNooDwMcK8AAxbhvFjHaqT04EAD
IIkdAXPOzFy7A/benNbIZBk2+p3Lwa+uo/YnaQI0q2nuRTw7nnyljXzD47ruataSES+226qTRU3f
S1MILKBoXJPNflvsCXc3TUK4ty1QlGbr4UHd1QcchVDo9UQmhA0syyCuK7l5gEi8kGf8AJer/f15
96D76869EW+7NRKFSQHN3BkUFaA/ejmeVMCN0ST0LoDasOluqhHEsITZ/SDeVaq/6y3dQfrq21o/
E6yqcJmztX8qrW1LpySQxhUvlZNVoOXZQbB7wLU2p9r1R/sxChT3EtQN0cpU8xFyoa0Z3+KVotr/
3uYGWvuvZMkIhDkaBCrB86RlekxJN7iUV/FKD28zx43TYpA8Ca/QEvy4FCJeZAqcsxy5s5IYnOQo
LgNZsgDw0X8akUWlgWEMYtIGriulxUnZ1hfox/Ip1E+WRkgr3xZzuCskzNJPKkdxSacRkxK4kGUo
etk00cvVwwsjZI/wwLWlwThKghKcW2GQgxdNFSB6cAq2+sL5D78/hhXUBAQMwjksRzRwFkV33EgF
ZnaMNj0LxC3s135RHJrYiK4WHSOlvG+BTXOUMqGv3u8o9A45EWhw0eqnfGXQAJFIVXrmUiDpq2Zv
2XknMHL4/KmccVfdD0vo4rgFGH1ipWMSO15I1UgC27NQXTnmlt6Hso9XnixehcXq/WP6SgDOrDtj
+MEhLOsp1lBpESffEkQC2kl3lfHhgzMhhab2Fr3bFPQ4B8n27I3OuVrCKACd3o0JHDIkw5GJYDRu
ZpxJoiDblL30/zNgos0sPWGbTrh+Y84f4HX4sPtJIkapPqcJisw3EK2mBaKk4nULIYFXV+8UaNEK
ra3nciJXokrs/g8FQkl8sqqj3mKE1RhhabSceZl4X6PAxCwKx23tkOrWLgW1RwIr6mmD/ZXntrMz
En/9SuL9FYThXpq3RjtD7afOXbKHKvIgTwcA0Rb8fzJ/tfSayYMzfibZACYCAZRchWyimTlJu9ux
IdIpaXTmaZQcohpAj1CbvUM94goJV72ma6SYkT7VEGMnmBGWU3htlvw/xVJOqkgiK4X1XRhQWQ4l
pW/eHh4WJHn848IEizZiuw4nXeIBL5CGBtVzqghY6W+JuszoBYrpvL+PEEKn3nUj902Cggmv0D7x
eShi6S+RXkDR6NonLyXSpJVlOUJ00hO2T2iJn8vAdOpLXHkWb6JqdRVJXNVP0fDE6uX6fVCJsjO6
gbyXakXyBp+qOSLomFTpXx4bZsl1aXjRyDggCbQ4VA5Jw+imkCeLpUr2uSpxj22NK1nawi1Yyeto
my6uaNGCo4a0WNzdjsKV4WwTs08Cn+mdsVychJUYFSZtHOaCdUrmqXXJrrYT86KJqIAXvR8Pb8IE
+kMMb9vRsWJo5YR6EJDDQQxwclelwFLOgCssTgV5mVaaigZGJNcHlykHC5xaZtNhwy/Ivy5V3nc0
IqfQoXrrsGsXVBUIdj/5v6eVvAM8stjNx35HSdc9Hf+JmNby5GvUnbDNEw9DdO64jOvj0kW5l17s
1vHteYH+0fHLlxWQNVP8M6/Y1P5X+X2gyc6mX9IC3a8CYBjHhescfKPmaIHl0u++m4yuQEPCsYfs
YLwK34m6W8syORqcJRHeuT/WSO7GmKCoFAnRCADxgo/QIAT/GzUS5T0jeJ8ODEf5bSDdKxPCc/wf
H09EkbqqJPtxtz0Kcmn808rTWvb7JMyOpxc2oYiRJH52EpxqUQViyc8toCglTk5cy5/MbgDkwlYR
sJ8MEBuX+VGg8V/BBKnc6TNLEqbToLwfQk4EIYnIXXzxoj2f58DP5IPI8kDmZWkhduW+Jr40TxGn
L3XQ9nLr9suFJ5d0NYvFBV/qwgPjeh4M2m9bW0OMFXLIEkZQdE6cucEAJ9OVijBmQ9cgejQ+KWwu
bYKBbw0K9/K5ZaNwTqpP+OlJxNM7tl0cu3hdBQBXFDdjygRocU88aXOrJHu0KUqkKIKTEE9ebtDE
mDNgmKxJ50MIfvVMOuqcIBvciU1I7/yca6AUrSzPXduyD6JhcnRVBMwW0v6hDtf0QxKxqaCFl+9c
PKRfr4GEJ5DaBQswA7oAsxoztF1WTlKh6BPPRz+viI7vQYk1UQrnLIn6H+6KFc97VQSTG01ZMaHs
rXhSz9oANi5Xn3MuvsFgqd6yg7zIjkJ7Jw1uwJZ3KPrY28wcvPSOHTyY/KBYq7uhT7fNmrK+og3g
9pb84A3sQwA8SxfE2dlwoAn9bnmzAD1SXOHIiYApgFseOkNOU1Sy8OeJGzWcp+ytvaN7xVxhoy8x
8qmKBthIFMs7A5a0qLNax0OJFsr8Ryw3py3ZWGDdTBCmaF5nH/WYlIZs55iM16Y+i0oaOXrbI49B
EYl250ayNy8b6j/Z0NKd/QDvIDSQB9cpor0A8KBg8KRt5z3caTKSThoJcryc3RJ7e7nVbwjUW/v8
J3tqYeuPJKIlMzREcw6sDPd8FDdhbKRW62hgau88fWPkUV2YvdXRrZMX+pHjskFT7y65dlQoJjA2
WVMgpSZsefUfYmjl8ghTTIaQfBU78CpOElEcH9cxKdN/XOTUlkU1xQpvAeaR/ZOEsAjgUZUeuDAm
2aBfwQvCBQJmHwIcd03FDgaPah9mbjaFE1PRlI6LPjemFANueUdc1i6V1q95pR8vWXEov3ieteta
1dJB0vCYMvyqtavO8Vg9jWGbz9u0uPMXhNxJLjJ8h5ZAjtrZcWTIIjk8v7hbZau+psU0B/oqt1P6
T+DUBATxOSCJcNvOZaH1nBxQtP5z5a+UhfkWcXdaNJHRxUyfIJcL1Hkfq9tQ/PAJwzxIJR5lhJ17
O+v3ASi07E9/crYllRurSu6onFyMdjaX223DE+1xzahQEf5QrGCZ4XU6KerHKfFpFs/9wfBaq6eC
iWzAeQXD/k3WD6HghLXuKDjjSpfnK5Zios1r7hbOgdHsUdseamAPXLby9FY1F8lkHEU9KrdgEOYd
/oXBu2DtSQWxudX1TMWxAPsc92vQJugUWTreHspXElNUtVPNGSj+QY6o58HKa78nYoHWnx7a06IR
JszM8kR/QDHL3xpvPLMzqdSruSsyk1ReFKTjhOLwgC0vHvhLKSRrzjlwrAD+T50fCGTbgY7C/SNg
oY+xiEvjcP54DBPu423iHtsgjUnP70YtW/+/QPjw7SauY+oy9lxKDs/UHkoI9lJQLnfQd9EMWNKV
h18aocCDMFMIOHDskl28ABxrO4NHHmq8Cxf6kjR3tIynYxpppdYQ63XqqRID4NSZ9GC+kk6TccFX
/PUbqYonYSYwHx0CwVw2CUXoFszR8+TTSeBxz2kDy3xrFs3x+9Bdrv/tAYvVeWo1H2CKVsfHMwQA
P4sCsrEtsqrILvGiCHObZOqvMnZzTVs0ioTFUUxOVgoW70dvJMvgWwkvjE5guYYnby0YFWB4OI5H
Cuvuck/0kKk+IYqC9awXDbZDHqlEom00+7C80/GedOWENeb5VTIcioUI3zSle14hV+RtBXyY2rc5
yBdSNSp27OxqJ282DWtDI577kr6k7W6XiA5Cs4sgGbSbLqIhumLhAdu3zncUXCZMhgR66ZPq6B1A
yCniR2ZUxmErylxzm+Z3akcgKMBwCJxrNSJq3G7I+RXV5fhMsE1Unbww7Jm7RhgAb4Xu8f2Gs7tH
QuOmfT7jFCnSZI8cQrBieu0y5e91mlzrrbCw+P4trOGgm3htHKxSWZ1aJjN0Z+kwDchzGDoH5pai
ukeysNPxeLq8gatq+UatjagJ5x5avX4HJwfwGGCyppROiND+Jd3CeYo7HcwRGrg14mSK42VADS4k
4yeOCW9CNZEcFcPlY17MxHmB0jqmT91JN3oswjnpuXcBZLJX/nBjgtuDBR88YFzj98aXyD66extc
96pSSNPIrZncLZzPYXH39XpeH0r3AgJp0YxhKgQ7HLzjeaThZvy1m6C1jVSGQ/NnZjkH8OWKpI5L
VahOxBMWMP2+HN2W4iS0WUNAFBH7H4Vb0ByW7OUdoZ1HZGaKB/rKI9uc0RIF0mlg9lul/gS7Oz2V
aZGhP5QcGI74Wo5dPBViHfc3IphZKRqFtF3LKYjMekg6AUCFfTNKSKGI1nmrg2zLN5ZjmOuyTppA
+FcCjla+fyhjOjjB3B+/0yy3hnzX+8vwa7I3KoySE9CEok7EH7oISBpsFfsfmRCSbfOOGLzYYQg7
IelTW3iRDJa+7kwSCSsXu6CzaOqk3q5pUlay3YddtuvebNJITY2MUOBLqN7qXpeXOb3B0wl8kuBx
mUtyycVJL3ve8jJ9c2Ns6l+3SFJTJSxDf1uj+Fqd6NFBs8z5ZTLSTmkNro3TIkZ/kMnTr7W0D856
ZjtRExw0SEAAIj3TDehh/S65U0JRDylWWrL4IW2zXa1LQA/U82RrpELI7QKuU/1DQHoopgYBmo5W
kjV2aLTM1ZqelMUywszEBo8UsM/r8EjbJQSv1BT+qKEOzOjHFJotfcyP7lfsTnK3QIopVGZrHB3+
VIMHpN0gFfxDFkVwBBtTtsSaIxFny091Hcsb6X1mIqAqiDTxdVcSTidPL+Q9YK30ci3FzgEcKebg
GKC1gzgwYt1wS9PDDBDAhkYOF+RLMdR38r5o4qT2ECvhrfsSWBiqYuSnbNKwWQMRiQIDYWHkxcte
8VUooHLc8TcamrFVLr3ocl6kEq8J8uLWmBFvqolKY4tv4EvqPiP8pt8/UHI6lnp+n6NK1BsyUu3c
gElck11zE/1o1EkG3hGcPtiYIjWgnk9BTGypzi4yjjB3dEy6VrtG6lYJeQ2DXCatWfOhuH0oU+tp
1kgcuLcai1aF+OpmbyRdScuB+209wjBGhxNGf4UYg3bCC5R39s5W7UW5WpMkq8Zva12pr8JCi2nY
oVAMjiPv+iMraXhXTZ3EPHpem8Y2OHdn/2lgeqtuMv7zB1V63t0YWwhEE0xeNfo6++1u6pLCpidX
O8U0HkrIx6lE+wPFae3mYUZQqwAHQ17o9DTqMi6WA/LoFyScFipIj1bpr381v5cWxqXwIwcAWuV8
8IpJIeXzCDRjeYrkxvC8qPhgSRABnPM8+lpgF2iyoZ5RMx5mtIOHiTpfxSDkg2SR9CJ9bE0QJOH+
EMuL3EqDvtqFeOosul2s05gjoeClHszXIR+3MuS5NkyPxybQscNKUpf6bJ6OnmVw3gdYDXWx9o6/
QVyJZUPSVQlFmuEgqOnGuowtGwOm/WeYYTf4JnsALIQExBgIy91zJHc2VmkpgBLxZ/WLnSLZBjzC
dSOAyzVZ0+PYTKTuFDsgr5+vCIQY9RipSt52ttnqxPzbd1PFZSNuQVPO4jYIR4p3iY6deICmcZrd
vCzA8EIGTUN6SF5Hw5KFXzQLp+fRzVw2DhBa8H53Aq5xEn0Ekb+ekpPofVvtBM0dCjd4EelgGblI
p4H/cPUgwkxEgjTjVcSYoblN3fYfJcUj001K67xX22iZJdywYYfU2ryWyg5ZHpX9dnLSHgrlgxdN
Z/eiFzPm9SUTVvJDzz9Mc7vPjOivqdvJmS9MywK+uModE3gkNFZXMauGzgMaJXJtiyGxbHXiKn5C
b46TNeew2meCMpCQxkSemSn1f3yp5qRZORV6QV9VaVQW6+UzqVPp+slikpyJAq86SM7y9G5T769B
dscjwJEan+Ipk9KNQiBZKeHLbs/btvcs312x0r9z6vrOserOPmv/ekGctsWvfXbWnFQfQmLnQ5ps
itjC0zfe/j3cYsyiHZZj88Gp4Q1HhAKBquA94m+XFJuxVWcmMfzrP76naEtZ+wgiD56JLPEkkbD4
yK/P64Lghcaz506Ir6zr4WtXP5nkVSJtrYMacRmi362OBkPPs7GvsxkBfCF9E8PNQwM7xfzBf9fD
PQ7Bv0MwSxTCyIx28gEULahlwPhelZmHsVNU9khvwmzVKxjYxZSTgIIfU8pQ0HIhquTYWu0G6u16
EsNsI3wprVG+tp+lBqltQgIwDl/Lwj6rp5DdlXIixTDhCKYh+DgwtFMZbJ/MbmNOe8dktj7B1iIv
UcLerOSRAq+6Fcp6yHBshO28tw08uY1l1ZNBKVQl/kLDc0r42vhYL1EtzgSyk+V8+oIJkHB00lzY
42D54DXAsYovsZGGS6USY8cgYES/HPTJnOkj+saXFyBPbstJ/2bu2/7boOroK4A5SBAIjEbZbbiN
nprA+rw8h0AxHx7M3Mmc06QShgz2JlNNmelgMldLfkBDKvJIM82YmUNtRxfHsWVnCrN9v+HYHAk3
pUlrDfb7MdP9xatNSfhAHAqwSitrxLcA4SKRJ64tGEUsAK12U2FFRDCWnMaun67iJl9GcLJSLupN
q+mQ1g8LOKGPjHBuYr0/ET8gB/+vfX5LhgJiO4M+ho8R4d4XetQqUPkk/V+t/D87SEqYSyCW/i5Y
IQo595IlKdz8VtXkf0cJe48b7Ep10swiulq1IBCsqNsxNZAwxwnSiJb9yn3NjED94BPW6TNQhbv6
ABX1XLvwDIo5Be3glelKXXs2OozxGh/iFR+oK4BzWo7dx1SGfjqFmuhagTmgQi339wCWQ6avMYM4
D992XpJoeUthrx2bNgs0jGczg+a0A6syaMMn9W8bPLxG/zvkjJsNTlQzPsdPMjg5dm5IKExjH2U+
0jfzLhhiMKqO5sJzU0/e/5CmE5Dlc8u3eZYInYQmci+dPAlOlxZTMFzYj/qo5LXd3ehwzWZgNocS
9k+sGOIw+pEQ9lfDKvmshRAACkzPpyn7qbEKqUpMNNIYuU/8XJ4056q9Eg0r43VZr61/JMneBARU
XA9gkU7EOZUvcKdZb6/p/E7rtpLNg/x6DXiHrtTT9gUOB/wYjZNYasDSWwX3UT7+YZgZQ8lpeGM7
v9kXxRO26/NQ83BQej+ITepSQh/yzcqrMQTLFXDIEvYzDrO0ZZ1y2bzQXfts7dTIIvZr0gfCzVsa
8CjnaiH0mtTYEqwZDoYEX3yEsYiTH4D6ESle3VdqOBdxaHWWuyxmcRihj5e6zLps+4/PrX71ntIn
Ar4U3P5H3aO4nCzzWwNEfQueUzzuKsAdjz6xkat/XzJSGo1tZFhfJPjtKcBU63Lz1d14W4ZAD1HO
rlnXongqUSY38Fu8VSVzrowBCQ6Cv5+fXeWOrBwUf/SYBD+IO/sBYZuT1CZ9m7Ouaw39EDnjYgGM
Niu2vI4qzqMyWyOdCbYx0IW4G2TpYhKNq69VIS8ypLa1TOsx20hiUxnfOfCyOC6gt93vo6bqWrjY
rMn1XQXcVYGTSVNCwE+Qc4fcN0kAdgF6XNVvXD33Gu/L9aMO7D+k1+aHfIb/09Wpb2w5uV2/1VTL
bD6TR4JavILQz8X6Aa8ie5pRugoaq85YSwYHs5Uk1c5sampMBG3NQngMAtbe9E/Ozj5awTFxMPW8
4V784xgN7BZyLNqeRaz0QDwVNxTPnWRIsjKBCXpJqIZlp9k5k8eAeqduq83baRNfemhup4ph0FVf
CVVE7T1FcSqiDOPraDOLqbSnunAxx+0bz30o77JfOzVcOqTHz/kiIlKjPTz1GdXW376y2+dGBgUJ
GC8+bE8PGyUV4VdxdjwMkhwVprJmW487HYBm2nDjxvObABWR6VbhPNopnSdCIqGOGraYb8xZgyP/
3uHJ0N1M2zwv4/6lwXlRJDNwVwM/QMRh3SFQtsMUJVXh9c95dju4vgnI+FzX/kpFYMARuVfMUQJp
4DMVdn7H6EWR9JzhpGOzxB+XOOpiuHlzRv/mSrIGhrUxOgCey3tgDGRkCNc2Wxkr/h/Ivlj5UfSf
w4QNgXqUJ/qVhjgzIclu8QaevXAZ2ZxQ+GGhi+QVSNtZLAgsxn6gYsuh167MNIUJLhnFW9xFEg41
bja3m2KJnkWtTXM7vUldHfCaVm3/ULXvt1L3Ky85mfXIOlVIJYY85Y1h17Nu6ceMaoiYLOMDkMJu
C6nd/URa+o4HDdaqn/sMdqXNf8mDBBkJwG3Y6Dbd4WETWtBqt/fd6xVLqVU6CZfClGBn3gZom5Gr
L0cH8xOgPNV7PzJ2+G98GOR507ROtcMtLMlNpCm3thAQAjcXpUQ8s4H8jqM/9Cva+EGaPmZ8Cnbi
hfu+RQ6SolpGb6DGmOUEK+ZStpKol7HW4ZWRbRvbjMSbEKhWezBsV8iYCv5ryhwLdcIir25b7Wzf
ha1U8/1oLW0mkkp+gv8G+1BONKhL33bdh63KTf9LwaxXQUEaiu9OC8pw4U2tIxHvHuiv6JdN96qy
WO6H6nIpM7CCKtiTjBH/wgGAg+ch3r70IWXiZK7vp06ikrU6P2gtif6d/Tm+88LBpKWCOGiQb4ig
WjLcKjoYPylXUpNNgjuC+/8ac8QwPffvrxNxdVnUoMhNC33GvWf3Oiz1X9TpeqKiVwXnfRhL8F2T
2tHsC3PUDGdUIGqf+/P2mLiE7FdZkLxR6WfSHAmY07T5mNPNu2okDKszB6SHdcedgqps1HqNBcqj
DGeFHhsqGd2ve0vpb0JcKDWzq9nRyTuiv8RgP4MRj3Y3HK4Bf7YuiPSG4JeKk4Pvdx3p0nQMQq/O
da45bYHFmM758RsgMqlzdBPDL+S3h4kC2rclYm8pmI8g4+CtUk/4eYTC/S3d7Xis/ErJyLE/vG7y
wi8Rl2pFXnB4E7i0fjqLaKesnmSbvJHSqmWTF5AQbiQajwTjEXryEQ9JSzOJATV4YBqVaprZexof
ttfwnC9CQHuqmmLwCXu4PmZq49kasLJjOdD8lSz6EQ8OEuD69U4oDy6otq3Amh5kb9t1dsgc70CK
R3zLSrDe7dqqgO1fRz/vdy/TDBSMPHoDYjxMF/JFGNUfH2jx/ONGC/JYzfwXP2YS7JEXFLFCkoEq
3Bulm3oOqxZCSt+ILVgArPQCyUCQfSOT357+vqfJJLOAZAevUJonV7RUEGf7Dh9CUDWlrSnghg/j
dImq4q5z4cyTIzH1xiw/nkqr05BzzJDMl2G91VquplXSaGOFbRVBxxyKnB+urBp0pao1pqJSW0vM
Ee1A0OhZNdPVpbcZkaNGHTspm+8o7kZBWg/KzIZwZ6j8E/On2YtYOyuMpDPDj4znt2Jq4Vzhmclw
1nmcdY8c9lpu3BuL6wj+OZf+eAYkLeEGmfyopnosHrL2bo2VLDKGxcmRZvdSsa9z2gUvqwrCI4Px
423/OWCqrGTEQMGXVExFhOK/aKOEHmxJ+pt9csn9pnDnE2NPH+2jtx4X2HAjSXZqgms+mOtOCg+o
TCks0FgtnRsCpEeIizz99DFS9yyMS/qC3ZOivQHgQlZsR2WC2oTAUcl6FooyF8u8C/Jmz1IMhQiZ
usXRyja7nNWRoy67B+tIm57ax5ncaptCbjXGGD/XAMmgKwKnuMVYBNJjbkDTOmYXJ454QvvXGs6H
X9l+7uDwV/NgjTZtZ0LStPrY5fx9Fe5ZjWJ6PFmdhiPJjJAO0uMI0ionQniCVALzGv4lR8+ycIkd
9Ka/ZwjULIiqj5OswjFw1EEuXz5Dy+wV+aKd+LbhLmSLM6nnb5gnoGyYpUuzuGBNcQNQKAwclUVG
0Yu9JzejDPBgq5Pss6w1/DY5g4foFeaW7YXpubO38V8YqgR38xrNvMrRMJkf/Kwgb1O0d39exZ2Z
Dri6oFpMkGB4juvuiv7owkqzS4AGZFAi6xoKCBWUeqJzDBpnZxcoFISUx7Czcv6IlT0fHzXgvd9e
opAETweJRNWLqFzNZ8M4OOSsTDqSfDxmT7dCz5gmex69DVPhQ0cTzZdTq2itn3GEqtb+WyAp8x3o
x0C+88FP4TNPmpeE31dWkaJjgI4h+DGUcYtra161Kh0fDlnrKH3DeL/BiY8/OYE1rfQp7c+5cYSF
6FD3ImpjMghuppwX/D7K1syalr2F26Lqv6TLBO7+Q0wo1r0v+AHG2ieljDoGDKVaRtcj34SiR7KO
Oms2lu1QUzJkkfeK8966fqsyrknmJypjyO7GMkRpJTQKHzFlel3zt8yACR0dYg7lwxOV7N64rquo
zvR/kDFFQDsU24nxhpeaBZjZlUCBMuyTLCjutnFWPIOKhm4Ds0U6Byx5rqycFDwzrBBWyMGqW+sO
bJb9XumZwOd/FEreSMr4bc2d+UItye0u7qjUDFevt5i97lmoJVUXcdtmfe+2ocaJQK4rVhPgHU9x
WOb2ue4qOyuDc+rEcNZLTynSRgebTHcxU/In8AagMo4NSjQ5z5Rf8v/1hKDe4pOKQquBBxA1SCsw
ZM5pNhbY0wUGzmQsg3uuVVoL8/hYZOENLNLPBq21bJCo2Mxf86TM4lO4DN1h27qzyhylEN0mgWip
xpNwV+QdfHKQJxet4yS5Gm+SNpT4/HL5EEuHSFGomGnxa90Kagsh6R1hvCMb7iVMMoBIuPPQDOS2
oWkG+tooHQtEAiiQENrosl5lxfR/NJWxCZAbDQf/fhCMnxJihf3+/hGGfMMHKJYG6l85859U9mVq
LmnXQJg+lJoTKRtMZEYjA+1EsEOR48GgjXC5sQIw6kq+Jz9orXvnp5gh/8oh7xy7O7Cmls9n6nCe
xGGDu782yJoV89ORR1LRwjgOhozMRu9AR5hY0lsTMTmJ6gAMCHEKffWVe8jyZsE+6G5jdEJaOhIN
S/layhg5INvQ5+WQjPSuGcvMJ/xEm4OR8jDjK5llq8er9BIsz1uKyEHhRwgk6cKGEGdU0GpdV9Sj
riHDAvlw+h+g2uwp9Ni/drztOyHyw938DhmJK6LShLmfxFNOgjKMwjkeBK3K9StchsDTD/7dz3L2
xyu5TTh7TdbokEtiR9lNCGKDHj3yASYvH1i4JGZ0s2GQvhxkYuKPmlax2e92yPxYMPteq+EkYr8s
PTvi3Mf4Bry+khG9/VKpg112d/1KOde7oNAAsjS/jc9oLpJAFpg2+eZqR8Qx8L0PiAxx528Qsk+N
rCJNLKE1MncSnF8IoC8YV/UroKSWGm9pSKe0Az6OvKft7MgmEf3nPUtB3YoGXwWiyfgUzpOMUY1L
fnkmLysKf8qpFxW4FQgVPpVdw5eE99bvkhPNslpDgY6nOrXZcma8EqkUnCSq7BabX4QBwLK59luA
qPtDaio4Rudrv2mzHc/p01hQ7Vde86iylpId6l9HMUyt5LGFJGXVYlvqJFYWWXZmZF/DEIcQ4n6c
SCCCZ9XWuFoNBEU8ODYrAHBZxB3gu9hQ3+1B1gLM60o6Z3tfOpEp2m4iIYaxAWj8M/CIM6c9sBLV
AoZUEZPAu9bvzJ1iOA5dswFbjrAyFrrAnd0kBmJN/Ph5QOGG3RCste+3KdXH0YxyvtwNTMsWwlZR
kcO0gf7SI8tK8FBwJztt+mfhsiULKxQb+W5qwJLMqBjsrwu5ax0+k5D5RNiAn+wm6ohKnmucXTL/
iXvuwRbC27tyAuhK7ROHarcDSq5Sn+ETum9tviNxD8hQ/HVqy9O7WyabCg1WXYyJZX4fGfLVviB8
WM84EOcok/kNSmWtniClBTF3SxzYePeFX7tZdmFv3JccUVXAAh5PdwzeKgcKe2oBHIMB41Gctv+6
fcU5x7bCQroAgPiZ3ocPcL38LR8cbNJxoWx9obRsApUF8d56xKQcAyaZQhzsD9I/bDhp9dnO2vrn
KS03Z7FpfO9U+htp0xwY+ufHDqexqovQLdcqH2AdC53xi5Ze8O3PHtfE/4x0szPTHL+6oc7tP4zf
VDbG5tPSfc4PIVXk7JChMfnvaFvGML1+MXqYE7BBmz1ZEQjH/nr7QmrvLdf4dBqGJ+0ZT491NqjK
HYP7qq79fvDIaPdwnLtsBRtL/gJlD32lFM6j2H5fh83Ofwace/4ZuVoChb77amFxa8biqQmzb+ec
MRdI4dT/SKv4LAcCVKDQnWYJQyaqHIzPzx7qTB+xsyIMQAq+7YIFePNnzZ1kTZnq/pcJ27M4qL9v
2enWC0HhYJ7JZHHiL6EQQ3TwE/HeGLvqpS05XxzILOJXX7cypt3IR9ibDneKQxemwWihRaQXSD6G
mSii/Ea8ivntGcZQVmu2pjEeMr0HeMjIF1eyBs5TgERYcsCquFCelH9igS+Qbnpd+gPU3zf9sNc4
OnvooWNE1t30Xu9Yx5ZC0YHkEIW7kmiBn8sfZm+U+k/8oEhUeziLi7ceSHQrtmSkNSCdX7p6r+72
NQToD9cnHnR4+7Q3XhQ21xc31Xun3q6GIBpPZISJ+7T+kvBFdDZwucdz//uqbuH/AlrVNmin7fjn
nlyQDtegzdxhmCql74lZqgsPvKHfhVU2bnXL+nmV/sTjLOKANcTiEggH95QcxnrtikAem6yHDpsq
y9E724XCjghyPk3qukpNQ4jXkqsDE5IvSiZhdhNyFepTOq0Py5uOdRxe398p44qzyEXVTHJNQGzW
YGUfaQIBSrYeWY6Tv9FPfH+ef7j4zyRMv81O7YS9D+sODyLGrXYqbo9EWPmd7Bb+bvu3N3AYWXD6
y2qqOo35fN4PWZGxREJjOlns15bkg+eq7DSNE1D87bmkMZzvjP4gh8itxjPq6hqqJGsL2a9KwcCS
gBHvq4AOd37Evs9Iqr3RZs2SNhT2WBcPQFE03lVhe6LfPcMj6azH7unPJZLJWNkSF8sgTHHrI6j6
pFGlcE0BPdrKQh/F6lVbNRdcxKhUvY7fV3kcliRRqy0U4/n7+X6xyj4MDe3dNwf1UQ6DROo4JKFW
lvb9Qtwu5XeSHh4XGET1KE1GtXPW/PY+m8DvrbfcVxZ+3TqW3kPoyICt2ojtvVV3geSwtmYyLLn0
hMsj6fJDfKnZ9RvIqBAXbCR4qcgzGl3xpbvgbIGGedge7DEpb61RD3Zbanoy8iN4z4n4mE9KtLr5
tecFRPdzhok24NjamEJDNjnKD08SC42L8Fb81EJTf6E/QRrkHCyY/JB2sjlrF2PS5LykuwW+dCdM
EX+0tOb0mnWN4agedEizmiooZw5yGnSWDt/9cqHJ9P8ZE82UUMTymBL80yKjr3a8l0kNWOiPyS75
MzENs4iNx5e8KykpNt58AsxP005TpESBQdrbc24bNlrg9bHiqD8ZPMzPTZ/Dc2SII3jzndOp8d/i
D9/IBBbyXf973AFej5EddD9AWunqgKAnC8HMoiLXWC07g5saRxf0PiVJ51T4Zu71DJaM9wYqsmSF
guLJzSswQ5gphx5KOz8/iAWW5d+OF+VLVaIihyfktCQTsA4pFJ0mWkSn3DAM514pQgYZDbr8OvWK
9/DdsXPMBzLoRssKNcIPVjOom0aOEDNQodiuQz4EWAFzVnjek0sYfhGUvP8wMWmpARO1mNuH8JCH
qVs76GcfbEKV39p9R9xdXsxXuJYrMa15wFVu+Yv17OSlXvOEj+X2j35L1Y4Ztb85IyLwKZiccAS8
A74icZVwJs7jBtjP+az9gI6V4yNKh2vsI6V9YOjdauJ4iwZRPOWQx9zlmQz7CWdKzJ3qLhkp/WTI
fXfa30nS/3ESSWXLCbcoNKjfkUqc1ntX5qE8E7b7O5luQEDz+qLrBf4pM9RJetpY/1vr3+NqPRpf
AehAkfOaeQQYMHUe/IruuAxKRFzDfi+qBGjuW3DgHe0PnhtoOZFpF/TUAMto3vYZNfOlAKXal+UZ
HGxjP6//CubYyCUxOpy34h1Y8wKPuaa14n21ZWC2cxoIDuPQptabW2BgNaLgIfF4OUY3AYHgqIqp
qhhP4V8sGMwoibOfSJDegnWY1o/LpcDBrw0UbJfD/Y4DlYqrvpKHK7MoI0q8QGjM01Se9hbcHPCo
n77yujKZVbYZDT8Q4P17F9GG5HcAlD5y5ZVa+7fFGOo/5/6OWq7ML8R1dx1RK5GUn5R7nkfL1wcM
I576tKKiXscfWVGjjSN+feU5UxzthZSje07MlRpbcFTT/rs+n23HA5ioKbIJaeDwzOzxssBn6im7
eWu1GkIz3v/06OLvDr1J75iHkRnT5U8MdJVYlISYrDGOermSkh1VSG0EqzwCtswTGSLgh5Pkb3CH
AB/n/tZy7XevMZ+V7WEWXdCu2utO3MX6MTUoyFbNysi8SfH7+us9f7SaLa9IR8jb5IKbhQjKaxwU
f65T4k+7qlsF0ntO+Q37Tkop71y0p0/IcQP7NSDlbJ86xNms+YzQEQd7+9H2cxj0i7MKDV3/wqx/
21Kh1y0JzYt6zQMrGuh9ZxYzcn0ym50flNUNiZxBMni2J2Hg1GRZRf2ns2VayGBYvfseln5OT72L
rRaOna+FYK31HkNV9nTENL4Ws+HJy6PCC9ICdtMjDnp0dOB264wk6s54ZDOWRMcPEUysjf09pXKF
C9gjLbbreURzUKqeQLyzjrOTcoN00LRRwyibkegc/+rnr01sPQVDXZmlIENg2mGcKAUbHgIQW+xf
+WHf0rNA3nxv+4WzCJkXeKkS/1Uu5gy//YddsZdXSGSj7sVdGfrn0Oo8NlcpIgazCvPypCaOM328
WtLQJr9j6jA7z9UheRFym1kr7spSWh8cJXjlM1cRJhIWNDuBJ7aTHtSPQV5Pa/5TDbp5IANAdx1O
fn1BTYfgThYojaMCH0LZzcwnCQDJhf32tYZjDKR1eZZhtwWFCCDjZrxGXEuzp3qX/8dz+lB8NYfs
RK97tqTzQ6WAc2NP4n3gOnuvqYzg/cp7bHjF2tFx+KLkcneS44jEHbZ9JlBXQ7W2QDdWA+aUtGh8
sEYNGSmqoiynNglCjCLu09127C4jm8P7hyw2hYzKKk1sZ+H6+ZvMJsZCL8Zdli8GDqvbFQ9roBVT
RdQTB5BjBjyloYIx/Hh8IwKRoiOyAMOAGANyLCmFolJtjJA78wqXeGvDzP9g7BmnBhOTlwUEmnUm
dsD2SrFuFIksC1xqwYDKCPzU5+KdN68yfOISyuPVYwLMyBVeXU6pnmcTaVYvN3zAVp+QyRjHcmYP
PsLpYCbltHrqr4L4Pl64XoWMWjsM+QQbiuofM7DZgFEjz4MVdU7WZUNNC93iUb1LtFyA5WeUyUi9
O9zYFmBNkTS16VjidU1uD3Jg+ZdpXn4T59SWQzDgPh36wOvEfMLrQ4y/qKsrGK5+l3flK4GG1kRs
1Nhvn2/9XNhko5R9oFNatii1gIbwD9VPnnKgfroeZ5htVUG80h7sXLyUMvQgbe3vn5kR1jfzpdxS
UPfR1GemlqNnRYvLyk64plV5z3omvjrPPll7SsWf9krjRXyrPCyexTwPLlWj8jgrvoI5+3M3d2EG
dNypIwRb3JbdvnIkPbLiV3bovIKesfFPpB2TqJwnxdLBioE5XsqbTWuEGpaezuE+0Rli1hJsXRUU
s8YCl6+xFX2zAZsWohPdU5S4mWWZd/L3ZSo0r4nGzgFQBikQiojomQa26bRdS3Y+vH+qFiNkgAbg
CBTdImELrggnIdBONXEz0iSX3HW76O3kzksu3/oZqdENtUL6j+dn3cShyY283w/28D5tsbfI2csb
lYw7XP/vpRPh95ebBdX/JdzD0P+QNtHJoXGC3lFpIdfP/sqLHxUAY311U/Rgl6xQdVqBEX9hpKTT
uC0kreGTKNO0+SS+DUGPRbldqtw5YVVrq2NH0Xg6A7ixxkvhZe/+Y/T36nUtTVS88sSm4NWJ08o1
d2+lEaui6t351hl6nIneX2Fke5Qg9D+f6cS7cgXEp+dGUcrtgbFAL30TklCA+IpkkmZKnKDMdQV8
xg24HjFwpcmfE27L4zxdF/yNNXIIj12Ovw2MFioVMjZlNO7/Oav/9U3Zro4FDx2Txf/mLPLFEcdS
qVcVIKoNLk9ZdSTozsNUfRE2vUXZms0FkebR9paRAiCWQUTXW8EWRx2k63kKM8zxpk0PwA0ymqQs
jKz1H9vyh3A59kBcDQFWrBftVR1DSyByFQ2p+0ymIXcST+a4Za9pAKuNA4qZvGrxpKYcXNmAzH/Z
3CuHdprUL3Sq6qMIS4SGDDFEPYuynzBNGJ7pxQpLv3Ukge2sJ2oXYAvTgSRQm3Jk3nrzjVSgDoY2
z+iyx8ljwAq3h70+zgBXs6zTJ+HfWG4FF8PM8IsFb0nrTfz3Y8iJuI/GZyagn/gAzRK7szC8OXC3
Rkat5epf12xPsen3OF+/D4fvQg9PAheq7xXsQp1j3p/OLL9jh4fNk2VKX8kT8klpmtZBHYgsyfGj
YWXX/NbBCPryAuHzs6x+4FNowzMNKEKpW3zPMFaepHASV6s4PJ0wgDL6CaId4/tWmKPEq8iphEFG
75QQO0Ohc5IoO0kvyIbcHqIt+vpDfJ7OHwWe2xKTjCzmfMJ/T1O41Ym1X/SlgOryZzNMX02Ey+dL
Zk2eSwukBl0TkzqXi5J1n7vS7v/uZN5C8fjtOwdicVG3aoK9/ycZkBAvR4HvZFYVZRYNGpeNGuso
t13wWZcufl7XCpdFfpMeTJWUmIXkQt2ny8FKg/u7qrXMwqHPB/OwjqsLJZWyCnjb7aqDMo6ByRMW
p4aLgebzf0YcGZVmAIbZNvkiS7ZMRutZ4KfbXeQ6jzR1kFLwxiU5SjOJNeYRzWOrxC+QJq474D7l
Fb1OxC3IjbeI14W6z4LMbRwoXjdtAKxTchg+LaVdz2PM5UKw4+dHezv1k1YskRTkW70KAk+MkZyZ
1KWWsSw/8ksZ4Q5V73ytlHq9RSs324hUtWCPzq12pzXYxAVH+BAcSaWIQv8H3U6s+PDs6vR4bili
y3KTEVozJs4qoeRWZxi3gu8Ts1mYe7wXGWj5lSqgNRcK7Mn3rasSIff27gIVrKq6HVQS6TOqhwD0
y5TnTEjK82SCqZOosLZo70aQDnyPxeRD9R4giWJkjNCutSRnsSgoXk45+TbVNCpkMmDYqnfrJuAd
87BLRUuwAEA42T+cT/vQxSrn3n2jG76Z8M2/Pe5QmQ/zsrF/h0W+KhDCNyk+2nHL+oTSpg1QLM0u
qp9htd9xlXQaJ6f3MxZxvecp2LuidA4iFbzP6SL9JoBLJh9aRp1hlxLm0jAfIE1G9+E4PB737PAj
sT/KsopatonDBJv3ti7u3YTtXR3jZ9tCfYSrwGZHGtgYi32lj84V9K5QqDy47Q27Z8VO+xkQwH1K
++13lClGYq6g2i39ZZHoUNPJ570XZ1fh7ZuJ80DSF3QZ1BzDXeA8gbTWueI1fX19HV9xyLmYvfgV
gJfbFi4YEqZsBfCoqioqi0OGaPJ7HErtmnPmiSqNFNXD+XFmJFGRKn9EyM52rIktBf7INYMNHSd+
QbOBL4i9r6g3Vmi195JAfKLDfIA3UpAjW02+OqKGjYz1PkPIJRn7ni+3nNtBgI+eM1pyTtJJUAMU
4rHNPcq97ssob/bkw7os41oyA6kfbyFuVqkDf91qM9k82hrSZF82HtDTBlz3BBz0MWBap0eK/fk6
0Iz0ZlGfavh3tK9OnVGT/xHs/Bk5dGhlsTky16ZUm4SFdKyfJoGU2wpt1SnqoW+DvwrGcA/tBWLC
BKIQT1aMpahyR5k3BIl4g2aPcw9qSyN4cMnz1/q59hf3tOW7klvqNZQhfPZx/d/bHgWY1tzZMzWu
d1LHRBYaUy37jWNI6+jbhcCL30XxMExzwkA1iCTg34OFi96qt0KimIEyDcwM2ErlE6GHTAc78dix
3DkECIOzWty47KgtA9rXKr7yDvJ1RhWztlBHMt19swIDQR4oAfKizI39L70EPz/GHXm5MGf4Pqqx
83tNUY4wY57kZYwbyiPE42Dle0kAx/SWQBKon7IJ9O6NckTbpa7wfmAua99irTREwnccv3rjmuvk
3Zab+grYQ6480JOo/IgOhQ1zBEuecjafwdsX3NHjObAP8ijTNdOOqT1VIRl1WUtfAIXvVEpJRcuX
mVOXmkcG8ceSmLepqx4upKV50RyY2+kNmqKonwecIoqH1G4vIQeRD2JRpEYj+8czoxVHJCA5xWTg
1oQGhgvxrco9a4FtLMz555RMOf5RdWQ1KhP5Y2Yf2FWYQ78Mo1T+kQGbf2MLizfx4Rg6fqjUdqqf
oXzgY7HPZUWr9R3v9EFFrHNolZFz0F9rEPMb7ygQTqH/2ItsC6HrX7UxzmhahadOiiLBw4xGrbxD
xSA8MczowgslJ0FD7c+O3UFag4hlwsEt4zxSsthBzQVW3yKwSunx09xSed3T5YEdGVRt+PXbw/dq
wuTEpNww9ftR60eax50RLZKk/Dh4eld76hbO9GIgzel44Mcwf1sSl4+hM5Jc2+6GDq3jINt/ERCY
SXeZTdkKdYQThoD3neMbUTBf9RSBVtMUHoH+nK6uqDMGVrNTBcs5ZnU/gVnFi3w9IlEMPiPlnfbI
hQDDSAoPwug22b4si9R//663FKdW9jxcZ7E3Omju6isFaGZ2E0ZDU4XE/jUZJifrQVh9vMLXh56R
DEPL34rp97CAh/dBTK8x58ALRdKK7fD4wwxPtNmfLli8pIHLsDzHKZyBaIa1dYGxDt5jg4BKQyPo
rpAdFtYFgeEKJFvIlhHH7F8Xcve9XClua0JJgPP/nDAI7zDYuwP3tbxi/ANjxsMRcybznkADEgSd
aTLTFQqq4pNfZjR0QZxfWbIuYXSnFQLKT/VMVITV2Zz/sKWIoOGa+SBWi2QU0N3jup3La73yUVTh
oDRUWp/JOnu1DTnFu7vXe2Di6cdDzod6BhoUEe3lAnR7yNMYZlbRP0rE4IrRyUp+jiYryqR6FkOH
GXsTDoJLtAZDBkppDj6+Fo+vmpZiPZK+1lcGxLnGLjmhTHGBnwCCnLUYa/b1E0F0ZOz1GyRBPdrk
S/PusRlCFda5nGI36c/90dnZUH4tPCk0YzEX00O4mKv3yMl0+zTUoeXnMZl5Nm1Ld6+aE6s732yC
OLYc4KVtc6ZJ0Ls4ilNywHvNv//0rYRzQVmbphDlKbU6p4OjJpDDOgHM4BUl2czpM1Ohp2fbIffy
OLA+9gUttRpkDbZWexSYsp7d7D9IB0iYJMU4+4dZtgNhkl9eOl+Dw9Lrh7e68+0JvCNMafvi0vzW
11ZbSExPbI0RBxAc7fSKM64LyvFuqvA644JI0me5pjaWPlKbxtht5t8Hoqxj7/QuhBbMfd3gzY8E
6WeX0NLEq7+8koiNcny94DbZzSELH8z8wvUVN4XGWWW/hNQwsrZq8uDY6ajsZgrETLSKjLFb+SCz
SOk/jST2OTTdr9/QaPZoYHzj84MGm2KEILpobjDa/jHstx4JD67pC/1Z0XmBtcJy38t3MXmaJGtG
kLwpAvtdOjdRwGpkh5C/EqsBAGSXWT04gWh7+AGA16uF18GGfG8AzTfNHuXCB5A8nIECpdPmqqLq
fPTKxTgPQUqLOuy4rQ5guMtp+6wTGIUzuYEXPqD7uBhaQUxFCackUILWeiTdsIjT/aGgPe7/OQt8
6E6CcMg5byJ3W+jIEKwhin39XyIKf8xGrW20A2jVOB6vus+3GPpANNXYUhn+mEc+Ln0kWQFw1UfC
TMKXVk/LX5tGZT/5efb0jAYrut91l2xoZF/LwTuE7EmZ/vh0rbQOPUB0SbTdS/JQBC+x2M25I78j
FQ+0HUnoCWjlnnellKa4ElAhfPltrHxorK24JhMkTFGz98ynEDjgxMsL8fCsil0b7Y00cSi24+zm
5xmxUmR3GnsVGpUJkqd7U3jmPB9mX7lzz8lEdiez9ZkKNGl1BWUMPuHXPehZNRWpDk/3iQ3nGPLr
s0a2WS7pdP67m++/enyFFzYaqRIuDBiE8pBlHnk/ZmAucPoHM5PbhHjRX0gLVS62kjxPA1SV74Ko
gPxzip0tADoviuKNjDb+TyRub7ocGHMEublVsE/QDfvKBfiwwqahvfA17zNPT9m1GXUA8M/xWkNC
B+yfBbJVYG+mKXc8/fkuuL21Q3htKNp5uVrubZ7XergRujXGniZgPXqoKVvIM5Z8vGK3LmAz7hJm
8nLaqRugycDJyLjZFDQN5eesdKbrnL2J/v5T24RrfEhVl3A5hQsMikHaxHzjD5+mP7oKsZ0C3XAT
wjsnn9Fp4H8Zny/QgULypZjmoYS9vKzDgCupBzcI3K6HvnhnKJ1WHYAhIonfYGcbOHKXM6Tr5vdF
mnjGIv3g5XatcZbexMGLcqfldxEDyccUr+kqpQly3h1urk/NqAQb+1zH5NsLl55/xY7Tc9lgWOYC
tRA5zPEdjsD8fOafPj3XjzUjZZxnc4WPfV1ZDxha3ZurFbZwBA/8CpiZX21S0xZSHtOIA0Hioj7z
yeIC/6kHo6cTIYIXyZNzm1o7IQm8X12cTJO8Ql4xxX1Fv2SN2vsBl9/KMCE5aUAUMsXD5m0JNPs7
5KA1MwigmAHy/o3RBs3UxN2RMjb0uv1/X0xp5SrZeeJI6dDoiEKdxluWDCtvJmpHDAwI/6Ldbswp
dQA6uNGBx3plB74M0pY4dfs3J/Io8lnkgjdPfY72SUJ7GwmiGmzwOB+Imc7yxCVAwMvoQgcvU0kG
2aUI/MYTcwEbpT62/VNwsOkRaDZmR1zHaD0A1N4lKxcamjlLnKYW+wK1zU93nHC9JYf9NCcEvfSX
5XDwooW/08DWtWYhTkMvj3Hfqa5QOonTO5duikBLHaFOf8SZzvslpSAeBZoS7CLzclaDS8ob4PwF
BdycscETfHDQWbPicoQgFn/9j+YB0DZbA71/vezgZQhgNtKxzrH4LQNPM29nh4IlL7rZS1u5DJqA
DSn0AheyeVj8r0HSfEGGweC4hd68mJI052Rxx1pYsePWIKIV57i3zoV99++ymWrKlV+zYxB3ze4l
bXFEzwURPefQgtQ2GEES4ttEwlQlteeZoAZLXCufNqWUJpHmtzTJJNtx49Pp3WJS7UNz8cd8aKl9
1ZaNtCSjbmJ8dzECEZPB69BgFwLpq3FFI9QlLOS9uaUV5C+vOgLDjUuK59cKxuxIfUszZrx4D+H2
+YLa6RF4+HxcreK0hsB0Lyhx+lMZJHK82zg5WSMZ3rc/kPKZatxK4JDLLKiSLK9gRC0JIgNSn4fs
GILcjdujq+WQyCqJ+i9+lcdZUW2HlDt0Mp3sathbM0VUjBvYPstIIZY6xdZo6/s8sypGdoVv+svQ
QMgl5vGcDxIZIzJIdiBMzEktO8cEJD1ZhwksoWyVY6CgCsuISPjFah945cYfuDazWRZ8NTsFSD22
IpEW5SaR/hX3CB6vZz3hpquRL4YuZz8pt87KizhenUubRIzVNdc4lffx2bzu4HQLt5WDwRcOP8zv
LILcr4rkPwrKTyefJEbgvPPCW56Bb8z1DpeQat+rvkye0L8aUUx4qrHk8XZTlYevFsa897c8rqe5
w04+3vFfvsZhdU0g6S91QjXqHKZ5ZVyU2/u/lP6hfGaRQDvaP5HSgCrXVHCLAzDCa0Ytp58d/dYZ
Rp3jAvSoyGEM3zptAOAo2Dd6FsTcjWUYRZ5aKiPQnUyCnHWlTt8G+j9w7LoQyzDNMp4BeKnrsRlz
RNp5yVMvrOW7T9dhOCgVD/nbOZRsr8XdE07xj/FKHfZhwJFeR0TtjpanjbUPP+jHxTrqLxmb7HGu
j9uCS29Jgdbs1gRwDTSFEETJWZR1w7C2JknX1J3ZlSimyw/j6bnxt2X8vTMU7kv+ge6eVCCZcOSU
BQDO0IhivNfH2QfAR5BgEA21szKpKmhBpyZtlrP2oE6tr9z3BwlKd2cbgv3Fku0yl8Fd5jkBakSx
enH53HXT0dI16WZnHSEfwh8pzHBiSgdncH503IKK9EAi4r7CWrvdN/jF8mlhFB9zNUaCwMAfyDuK
ddEql9385jw5V2gM43SbGTf+ahtTPec34SU+3ZXX2Eg5K6jm00jd05FaVuZKTFr8iAzLdAqEdzmu
gO12BZ2IKIjKU4cMHTs/2Q+7/rED2ZHLjioQ4RL8fCLYqTyvuffHr0N///h7gHkMfq0Z+z1f1QzH
q4fCbmdolQSf8fyjeTDwLaGQJL+mjo3bhZ7eZC5YTtE1sbEqKlF95hqNreyDiOP3Qkah4bcaNEHk
1+/lvxJArqxLuV9GOV/ZaBDu8Um4U3HrcclAWIHKeEGsPLoV7sxEbgFn1Kd2k62+ypOuq/Z3tOZV
FDDW6FXdA8DZ4q8QmfRfa4qjbnjeK7ybuJVBwMpnPHQSdfGNTsGhK9fIwmMdmLHmke1dIRpP7IOF
1T0dLRSa9vUEw9612Njya0xI6C9v1wFL7py9rLkHT32ISzJVQvz8muNZsQ3jxSyaTcDgnot3c8W3
wyeJXlMe2vVdI0KhSFKV6vQ3Ob+pNq1dUoIPgERaTjJUMK5jliRZkRE0yITifAyxZvYxOXqKeaDE
cchRthdB0oPcEktONa59DwGlLCnYAJvhv33NAUKSQA+iigW+kiNm2bt1oCkMhJqQSmWiJr1Hedwo
11D9ciAB/Y4bmT8w4Q1g3QoAkjNoyCvthuOgCUIrW6BCp4p8UU5RpW3Hu/996B5fHXdRXNTM88jE
o5JyyOkndSAOjsXOxYIDMs2mHXeQOnPH/fPCsUbynub2qatUbzDloIVmpp+5tR5GBOH6Lv+8f0DY
N5yfSpa8//QUNnPOdMyoegJdzqfKy2VpZ3u9MbRM743xy7zPFvKFlJb8inBnDJx5B7U2Su8b5R8u
Hww1B33vSTfA1DbjjyUk3lOUEVJQBKDvKYZne7bHrV+PalO17AHgxzOsp//3dCnkth0+0cgHm40s
8U4jfaegwX1BzUK+2tvaR8T13xQMCPK3PaVjZoSBfq9uqwPEQaeSSkolJMG/c1++XLbUeelQGFeF
J30mGCZ3yHzVCYSNx0E9OCITFoqlRrf0cCc2uI3BcvFBFy61/awLEsxAiO524543yyEG6l5SFmjk
Vrte08gnwm0AsmW7Y6htwiIvI8so9t/0PwY6e899HTumn8WhGkd1CS5+m67oDQbqAO+ey/ChhxFR
Wc4+McNjdumy6diect8fHggcokq8lVzapG+akArUGaVTXNGZACjPSABGejfBctpWarQ9OkbgXZ7e
Fhziu8vqL+tv+2Oe9Gn5FiunnApaUHkFfWBCXa/9R61DLRMj24BsmdiX0aFCyK8UyelnAlzT6Dty
2B9CTPfn4Jacp1eD50OiAuy25hFGKgmHBX0meu+Skr6o4NFRJ6azwTy9e5+YOlBu8QSizV0bm4Pf
UCkRqI9M8XbWb97zRQq/JiS0xLzkp5GhiLldGZpZoZimZmc9ZgiaQJGurqLbPcbFy+KeQp46MVV3
q65JZO0LKGWZ2EvMJwAq8E7v25hbrC5Ek1nuukSQ0C2Rcm/qykLCaIH5fA9xWqHy481KYq7bcG+l
JBnpYbLUyqqZaQBizu/2kAm+5p7W/jgD3mcX3SzL+EAJaEHDkDnLTf8/mGC94yVW3DIECM3VB5XV
xg3GK5fAODsJZDeigdeKzApp6Y/m55dZu9O4swo8PmHwD6RWRvWhRDrhB2Dih9GpsTfm/7ObBsdx
+9rmfixUSAV7Gi44VwHJz7OLJXfUix2ywoM9LDcBf5aFojR7iaxWr6kucSyhZDYJl+cpdSlcA3pi
ze5ql2ll34FJ2Dch5Lm51kOfjw9FE+xLjeAuEWw/JSpPmPiItFEDQvgoTZFhP4EMRvOfINXtJ1cy
Vj5lLqxNSRii3YbsOQQbJbQIilozVcWgy9s6Xuxuzc8Jfc6NjbRStMPaEDNrvKKIbRwUc+oEUm5S
YXmRPEDJg5kQCNgx26GC0F3ILC4CXjRW9fUrb8Xr2yj17mkJe8OOnZgjLIqRV8pfSGfeb0++M2vw
FBE++KzXZ7Ooi4z/JBr61rBots4p8AifjaGcgYEL6bhcei6snby36NFxbGQxKbjbL/Em6rpPbtfv
lQvGyR0U00ljR54/FeqH0fNHL4iwpdsxqR7rwV056Kf2c/6+ex6APUlPoqEBgirW+GcA6oBzL0e4
HQyH5BJz4Qk763v109HgGsDUtHL/mgx1S+eyBAPg7CaHOO634e7Tn6Jd1H+LLZ3iIshtAc/xKoZ5
15OC1HKM2rip/6AGzOMb3iZEpUX0ppqXe+6XLHIwA4qgBvFdlcPkhTn8wU5JkDi5N0DZOPwHIJ3z
mW9tYA1Dpuw00KgCOgMPPvF/WAJjUKfOPVg/ycs9uZxiFwzFc7/aFl9vPf3naXfl+5r3Hpt5MAed
GfiE+XxiOq/UUPYH5BDe0Pz8IKBaizEazGiFrz3cP1rX7ip3d8qdV7LB70Y1QForawiVOEhJS7+B
KzzsTH+RNHLL1Pm6+6VAD0YdTiNOb88dmD7H6zlLI4OGDXVObR7n4PNmRstd5JsbQBQRbROBvSeD
J9m4ObtDEq2l0sT1CSRG8TIyUHqjmSEXOaCuP4AxVnfZmhT6V9uJaEwMRS6i3IusNLmWdMWjYgdD
GRYEFcAduNI7HPaOQcSi4Voy+IyKpKgSCcIRMdw1ZJz3S2HG6WrlfyVHurX9htDHs3vhvCLoCzXW
AMoY/9GbSZjUd0SOfukHpkzyG2ga8zvrwqrna9NXLWd5cQ2hPztJxDI1V4IGGWd2va3+Dh7Ys32w
/tZTopRc5iAYqc/wnrz+2mXRhbiohMX6UFOdt7NLErKQ02HNL8m/+STH2pU1Q+rKrDYD6s0gWrEf
JOiAcubekRBET5A+2wALTCmiZdfACVk7p5JsFMQSEAW/FTQLDJvj01awo+XuSPjA6WohM46BBrYV
RbjnDfAKkzhce8zXC+sjF0CVcVOBgYiNlqluvU1E14Vj5RUo6xSqJr9TlhHiPF4IFZGcowcLhBCz
zZnZOjW941FrBNOS5Lt1DoN6lV0K+6tPLlihIODBDSaa7DECMxKtgMnkoUSX/k8rG8bEYq0C2Hyi
sQKFP/GYrRvi0HtV7V09GcXsgfKdFzovi/en8k25Nuf7MZyXb/auDWcym/4iI39B6zSmpiHMGp3k
L2o+g7ibYLW1GZQNR4dj/OHJPvVnVvgwizaRdFmYTDcz9Gnn4Kh3IWz6+Gv6CX7sndWKesrCvl1Y
aT6U3Q9ERVC4z5YZ4uoM4FMXxU7m6ECK+aa1WApo5aZy/KgFF2Yr0ONHgx+EkYo6GwQBhcfGlOGI
yhqUL73KkNzpOrY/TYd/6vJfW4JUNNlWkdwvVss73a+lo5NG+cvB1Esmjq4FBExWRKlXh/zbaVVS
KVFe0RO1AMX2NcR3LNSuyEFT69msyVkPoNyUe5cohOfYjuiYwlkS5hAbjKd3lNLeUv1C+0D5ient
tbg6FdXUoL+QECgqedLjDAStY2r6wTSQs4vE3pNUlL70ut1BZ56Ned9XUK8HRsn2Vx5RYTYwJWur
ExSBuJmonqbSZZelFe5rGRv2bKvLulcE55S9f24uPdGKj/HSWJBN/Fwl+HWkLqnGgsiQFroXt06w
j/hTueEtDzXriZ0T0+iWt4/7yNQz1LPKCHiu3BpScHai63h05K334+wMc7BtSDK7fpv8C2TmhbjY
s8r7UvxcNO/I7DAloRyJZ9W9fX2aD2mkn2eS2tyuVv0xwpfcu4KvbW6Rf7+9eWn72Zqm71ZNY0MR
S8FnhG9KKdMqlttZyzF25DPJ/rdqL5QTQkHQNKRHOYDdB2MDu+TAmlW5FGeWvLriRNUN/6zWoebA
hPI/TsGQN1Ixa2wDE5UtDVGzwiADQ/i0YaXjq94t1zqdwBtNNqBM0PPFI4zVH/elhzQvVLNqnLiB
XP/+aRLdmwjAbl3nb8uxcBDj7EMFq+4ionOTgAlGHRLLEttBqk0AInb6RJbSP3x0wTP/AgNwKICi
u1lybrdogYQT8xRfA3sA2+dj3EZMKnHtnebLf1kRtN4trKWq5M4FGyWPT5BExGJKiJp1bklgMAYB
/HXHzNz0yoJm8TbVN0IsIL/nkGDmI7pcPY/YuCf3GhcP/9r6+ccYtNOC5p9F13umJXK9tJQcUaoy
Jcdx7QtfNOKy1P3PFgQwSialbbjKJDZ+bQvR/CF3xCYlYuBIZRRvKlWNoExaA+2rurjYq3tibXPU
EaY8I1Z7x/u0FwV/5Ig5IFO5Z4FymrLkYJFN3PFeUxGJv7/WsO7WrD9Wv0kO8jLCNtf/O8I71VjY
CuGb4b4CgLIwn3zXjW1B0cTOB79cIB1nkgeeuqrMw++t/euUZHG7Ealeny4oLmWEASR3kT5jeaMt
QZnuGLjjxK8gGANbPzxwYyM7/v5IYNG9twOMsX34FWduxAggZATleBmYtD028NTXXHcQ80b6I2ga
gGtqzMIdhebu2Tzg1n+bClJzkmJdWhoZu8BYV1b/NiefulAXZQLqP3S8x+eNE9vMz7jqKuL0p5R9
UGghUvcIw5BYe6f+YXnrBe0EAqYHN7ukzQbUTUS3fGYeX19pnlKDAGS9oFhysOIaFnm4L/5NRSbQ
zRizSJLasDgFvfyYevxOHHZzND1BfceyBpHuA3llVqg+y8RZicuElHkZtbwz2R2sLOxauZUeZfry
5ToC7F7M8mxs8Y/Q0eN+Or1yFkSSrfl55Kl1ZDFr690B7tYJDuHV344m03DMhAXXXhCA7BiG772N
3/+K2LkoqzRyHNQcAntpn0v+LbGPH5X95tTq9GMNWNrRdBd3vyY8s7y189IYIxgjwbl3bl9iOcwA
5HTiuZ0HCXDMc750jdRaWc2Rm8AqcyJLm2UZe/hd2V6Lp2Ja4LLOmnJk3819QoTjBTtXZ6rgn9Cf
EeEtePt/mvQpvI5A1mHJn6MnpF/MNe3o6y3OuX37tNciEMIoi55peWlkzrlDBFhRrIutNfXO8hD+
IojO6AJRf2OrNh0/knfFm0FNeaSwIyoI+d4TqAshUK2weDu2oWJ6mlw4sNQ1VENbjBvT1snSFw0G
QHanYUTFj7kzegsSD2aCz0YDiO6MqvHoU9aJpO2GWaq5yLLW9gVUJ+tcJVtomLL9SupSf9Kq2k6R
dK26iOhcZKJGnXIAy/xTgNmgia41h0ne6BjpC0M4jl7Xw7l77wpAe7AaGNEdp0FFEFQMJTTkkCP0
rwk3GscOcNEBRLTtAtY+NW4nf/G7JlA//+xJWCG2auugI+pFlyRciPWXuBvO50zdastjnZd71nlQ
AD3y5wyFwNIUUgP7EKt+9Vp5R4gsSwCL9Yehwa1nCrrDs7y5/BV7ayrVmB1KkUqsey0AnMwtfRbQ
t8pRpxu86/rUZaAGmkPZdJjR1e+2yHLgMwK1guapwOOk9WidhlcnbZPmDjGwUawtWBQ2Gquhqolz
RXXZqSBw7jPQaItZCfsfaGiExEx7/TFVL1Lx0YIg3hh7wcPElPPH/YW6k1EOTQPkKbFN7NAyw4wi
RmgVLInu8n4yR0ksyOOWiIHjHSGbKl85swnWeXEt2x/E1EzjfOEI6CMV2Yo/mF4LqbGZO9d7txI6
6f434bN9rJesSB7tfX43jHDCJLSUKt8+3UxJuD/zNHhougErY5JA4cKAl6LfO4fCXU8AKGGHT4uL
4gp8t0Txs0Ckk7U++7mIkfzU2QberwIpqbJSW7CjE5GpghuG9Iy9Dcd0sqnZSelwIIpmuS1GQbxe
3YKIebLTGif0/Pb4SHVX4wVOJervDlsZGp8gcnTq2SK/vR2C2wBrKDzNKWPGTG4FjvRy1DqKGzvW
J+8Tw/vfJ3eiN7fNeX8OShWaTdypSNVdLgs+dcRmmEFLqhJUpnFkGATbb0KQtL4Apq+S+yILBG1C
NoCiLPfZSXRYCU2bJd5BOGOQqYi6F2XkKvstX/I3J/aofI4eLITAJkGLfPP5dOfot5xhXUoa1S25
SZwF8S0etivf7f4kucTLPiDElYKp//5RNi6E9K3T6dZhFVFtFclBXIT8TWfJjjg1vLKY+se9x4pj
TWNIXQF/YsS+J5TOXmquPomsEiTBDSHUpM/c6u09Fsa7crggaMtERb4sEjcPtxfy2lnPaH26i/kT
W5EoSIrbUJS3kCPyz6Jv1bzUG3A2L0MkoGED9lv5ZApDyaBSi0AbJj9atLWqAi7Sgfok6djJsXhw
iAFKsfD6T/wO8ejPyVjbXTnwGykke26UBP97yFIqss849R86zTXIYFfPmRZnleZBmUmPUi/ceLoA
FpqhjPpddACLgbSgcg7T9zeCB803cnJJtngxfN/fW5uuelGH1RKF8k6ORiJ6OBFKxHHC5tLkYx+k
/0iiBkQRHMmBU4tzuHl7oDHTcglbn54gjcGiUOTH/Z0POAmL+YaeaVGRrNEVFckC9AJ+glGkBsmx
z51WlLeub0U9w6MjTbrK4XO0KxMe2GJllS7TzWQPJhxyFdepckmwJijiFwGX5gyTJcEUM55fVC5q
Re309tYqL8rfY36Wq7o1Re0T1GzpObjLbgbOovJPITsgAhph43L4+XzkBkpOTAPCnPUnFXHLZ7Ej
rIir/AVMJAv8ppwcv43m/YBfu6vw0WnpuMrthTTDWUZlgY3Q1TeV79qs6cLh/dLPdi7w8Hcg16hL
duy9nckZBvCVvLlVdUBG3MHE9NswyhmUA5HszMCzD7SHJnsTchAx7z+jLW+YBAdbr3VTGot2eix3
/bUHcGzc/u+vH/1FgjlGsWZoWtm7P1BcRFbGC9D/aSMJmktXpvQYBFltY3cm2Vk6Iwbo+35ZaW78
+9DuuJJxFxbe4wA6vlQsJb38hQoovmQCMJFQgq50r6349Cx9kU0POBKR8nWtiE6gIANJeQSGKPJa
G5Omr0FFMF990+79dB3bYCj0nmEMGqoe3VIkks8ohtH1TSeGfl3uy5FuPbvjZW27Tdqp6enaFfWP
YOgjYyix/vmRF9vU7fRwmh1JHugqZ5o5i8n8GcCVElxSf9/rM+8uo/OvkPHkm7WtnjxIHYZG4w7M
w3K+K4eGpkOKE2jB+bqY3oUicGAHav4wkZQcbWR7Kwz2vLD48ASi92a7U5Mm/YoSx1N0sBCOFkvG
XaN4Q9YB1NuU5wEcjwr5+h5ZKgm6eI1aycpYHxgxfMfmRt80+dGqinOrsMVOUvH85Ay6ce6Pciiz
0CF4KM5boWBT5u/JK9MHHMGRAwbpHbY7WJ1kZ4wlRVpnrjJBwj28NgxSHjHJ+ztCvebb0Pn+HpCQ
kzO4AXlkL6ds1FmtDVrbU7K33dgkT8ofbwQUWWFVx0p9Ub6Tz6lsqhgvH/WBuOAJNlrDr3hroyBd
2aTQfM7vHndeSKO+Af7wBLubiBqlWVGhEciBlZ+OfeTcmL2SjkIN9ukXtxgXpYbdTxJRb7HdULaP
VgF/SlcdRCHGal5gO0mi2ciNaqrLClpB8wtgbABg0SI4DpM4UABNcR9OQvIpx5ElipNKdlz8px3K
TvHiUnuNtuBGXXWeBKxhQI0/1QDwM0iL7w5MImHTYYePwqRRdwdRcu50PvtUTgz760Z0fARQPowG
Zn77e3Y31sURHgjRa9hrt/dFe36OYhrx1/21uaGZtuRCiF2YvWDhZuZ9L/4cQp38M1Y/XemhdE9v
xHb7pBdCf41uhJMKn40FUF9U0yrTLKAmbRcUbmfSoGUCcMMiV9fb8LBeYGXFSDTFh0rmjNWXjTny
enlpVauPwYqAOe18iQJRjecoWYZZox6Fk7EFuCvWpZDVnCNckuyiGBpqhyXRGbJ41LNy9Wt7zfJ/
Cf5KC9B2jmDsaxCmIOFjZn+klT2hThZ7KwmfMPpfP1eY0IoXSUCizwDGuguSsma5/ys5O2gamRfC
DtmL/kVccEi2afYVPUwm1xuSaedCLSnh3F8sG0i/V+vLojDjDljumMbozWduT1om00IrxhxKj1c7
latfqqVax+8lFXeFD6vYsdnOg1QepCMZVPUCi60FHmHqjF9qz2Vul8qvNHBpI9aMw/uUgyk29Hrj
nPmMvKtvf1ajO+s+r2aRIC9qyhNwPbqh0KaRKaJnEHdcEoGlX99dZKGsiwfsY86k1FQP3hSYnPwo
1PNQbZ/N9SmsDmvI4vDxnNwXWbGFCwjiDM3ne1KoG3m+7g6pMGDYbgXzC6RQAAk+b9Pq+CPGvHS2
/+kBoe3JcRQ9k4Eq8FOOfo4JwsQBPWC7zgpzWC9dlwTz8D8mXby8uA5iNW8cz0h5uOdpF58YtL3r
Bvklr/XJ3s+fxjUgShEdDDRiKhOdsGCHx1aMJ6Dql31Ymn4zVmhZtVe1njXN0R+blypuRQ5p/zlO
Xr+lVpP09afSpuhPilWGO8iOhPVIKD4iElKRp8RPMBD6022jwa8ANhxekz6ft1hIBzO/V/gQPTWC
2qh0qhJ1WVtSmxfKFY8JipEVRYkwERsW4QncVHV6wHaPiSpk21Q8hpdpApMbqbhioSRxOWuZkBRn
qJ2c+Vb9YcHnIENL8rbB9pvX5BgyQQmXnh7vX7acO/JvTqrO9M5pMAqZC6UmAHBgu39TQewnmXDJ
NGDpAjpCo8ZrR9toFYBFxt1Im5pbAUz46GM37dUiAoHHWIs2RLAYLHuvODVSSo+ynTc4DDr+nPrt
jbUFMscTMGHVWND/FpodfnU5G7Rc+PN2dbfEzqUtrNf8oU2nGW1WBUUALX5UYBMNg7aMhGLyVZaY
uTcKUiifbqT48Aq4iqJVN93O6JuzxTT+qqLPvszg5hkYA6mtHN5E2eTlxppBgsDffecqnVy+zOKu
/U6KbersDJ3mRhzI8vpVQBhJ6uy5EMRI/eBdm48306u3DCtZJrlKXj+OU/bdjeUmZrgL2Scq36u9
iQUtdW5y6j302Tu2w3CywUGxEcVSf/7XICI3dF1Xwdn55s4ApTRGKn6XQrlr8xN/GrSyl3yPfzHt
OaCRKVZYspSs9Vbfnr/WlCpjRsk/dWHlK1XA4scTDmZFsg8hZ2ZcOkGbh/JVXO/UCfPteeVdtkIO
5eXJ2IbPbSmjd477snWcgzDNMhzhd74gEf11itKkNFAIeZfSBdIH9FcceKJ2MaskLtBpNKWnlmqf
SH9DOn3d6jSd0KIXfxRbZqnizTkE9UnWEsM5qv0PbZAB/JZ0Ig00oJc1hp4dAoYawRNPdSr+6nPD
/IgwKYxsDLtGRRdmsA2JQwPz8sRjBOTXeIWeCqkskY7odmdCF22LE6IKcpynSNMAAbq1EGVyhPy6
cRv5nKuzB4gmRRFACHtY2uvaURhoyPNp9poxBL89cPW6+zv4b73Pv2UDSHqF2BL50SMipDJYwkwT
X+08wreKfhzgvPQcCIpQBtxC0c2uT4dfaBhaaqYVpTxK475vZtxPecxWRvTS5TL/w72rysFI5CBW
dJeZAYn5qtokOLymA3qPVQSm0sTXS+CF9hpgC4Nv4ZNP+xGM0HTRHNEBKXBEQpaOWY/L8k+SRxqk
qdF+97lZfzPhbl2qZMZmKbuGCUyl2GVOr47dwunaTopCZ01gvwEivY28FtAqVbgPw7bbJLjaLS33
cnW7a5C2IZ+5v4Z+T1ms6f+h98Uvl/sIAyfIEKEa5PEHJzDfpAvd1OvBswaByijRGH56r9RPkEwn
QBHd78A0NmEhVyVmdppNiqyyR5vnrKA3D7aV+D7lYDMBlIS5CSZZamhbn8rlejv+fH/hbqZ3xMQ5
P67MG+ojrpUUDQgI53169z/FGi8UvxwK2KbPRMzRgCLid+XyI62LQTyDA6lpzIDfhousenOIJKqL
xSoC/vCnmipMyAHjA85dZSSraAClH1XPLK5Djn0pOEeZKaaRQw+FDBA8T/Ej72tibMCftd3x7fot
jsfXtlbIVNDAJgIf6TLvgE+wdQqrB52QVi4Nh/v8TYGHRvq20Hze6TKoa3+jFCHycQNTXzEXM/bI
ZlUmTL0vC1LXXmmw731jSazJFMMErB6GwrFfrSaDMZxcxRdfMinvojNZSSEFJ1boalL/4UPRq1KI
RvFazHKgHK5Klf38JFWdKalUQPoIDYCXr+YhTRwJm0sPGJTCJJhHdsYB6RdGNoF9RLf7O7Xomy20
ivBpv/+Ojn+LYIpYEKFL3+1DHJL7Fi1+IYfgl0YcrpWpXjTsjsydB1q3MuOIKYmu5blzzPzlmcFv
emIGJsFSWWmM14Z+vvUhD33xtSKz/jmANyeViCh0IWRMKutBeYUTZt+aTWVs2L58CetjL0JntDZJ
F304IWxak+48Q+b0xlAhgVrl1MDxDezen3J2LI2RUD7uhS6AIMCtOFJOCtxUkY75cDT4mitPm1xi
QS7EOP9lXo1EUCN/mzqvbCXS9BSAFtZ+3t2TvuOoun2U+ovNm8hGQqoHGp7vf1MqfIEL1NCGqAEu
AQryNPNBetFZrO2EzP/SomerPYHJdWWQXW3j2pd+1aE3ES2mXVcLHFGnbt8PhY6+UtAR8yOdrx6/
qAqTTrx2m53/fLJrK1At7grNk2/Gc7hAHBorhSva8H9y+qVAJnHV2e+M009lk3v1FDkzavs8sqZo
12ZTSVaqXalCUzBPf5EAvVLt6laagDM3F4a1TJKxV5pZZErMeqf+Wid1c3bzDFUxSqMjeNhciWrw
JTfWkueVQ+Ije3eTHaXXNeBGG5N3V1Na0SThKgOivr5tYqEKIQgev642Vi08k4qfGp2/FKhPtLxI
LueLjwiuyFlFLMsCjO0of6ZQ9V3+7FA6GioWDRM4Pb4zqx9yrLB/rDeqcH1TtDhaRuGBspNW75JW
XSVtx/XcTs5h16akxQcK6i+BR0JcAaqw8wcv7UJVya9xj3WfHzC8oUk/WDARnpSGcm144uimGsf8
co2zVGJ2jVv2xqxb3WDtPzrnj51ecv9yjTTGF736kSDSgACpBU6z9acjBCrflooy+pJuyUMxeVwa
zpE87eHM//1vM3+tCeML1AaHVQ7ycNXZDbUkkxBiUzV1EOCbFuNuy/85Bi/Sch4CyExOmo2JqHf+
XuFi4kau5Cy1oPJYj+qIYneznnMhWpDcgtLjgTDE5OccgyUVSkd4XPYsWiYLdLq2j02x0tMRjFaO
WrwKqfJgJC0B1F4YuD3iIo9YUffuiODL3JiJ+4gu9bOMok2+qtePlj6C/XbWp/Qp9oee2Y2s86TX
PaS7zCsThrlT7c1R48GeG02YD+JFuZzTMADUjf3QTSX8w4uqKc6Qx7mOp1wKSmevz8HKpbCuJpc5
eXtuT75OUbxKDySGne+dO1bQBendm+eKvkAJ6zpMByIfnTvQtkzjr8NnWHWwX+DlgezVEfdxWAqh
huWrCe64GkRy20u+HH6kZVu5E7UCHduNZxSkJgBdAUyMTus/DRgtdEzmPv7cyFCafoUr1HBYYnss
Cnz+klTavEkzj3V14vg9+RGbz+cVQYeMrYQkITbL5nta2jcEj2tuUA24GBgwzuKiWvr8/s+3hec8
MPFiSRKjdWYpb3gZA3yCVCxMo4cqABrz7Cdv7YgV2xCCadFVN627jKd7/LQqOmJzfmZIloDkl9oq
hazBliQxo0fsLHvggdYR6Lvjg04WG6vZ1qMKqdMqD3UsQFSybAMTrn3d7zy4zayqvb6GlPo9DF0Y
jRsqFNM33QVR+bRbbrM3y46UOZwCu6R8Cke1M0MQOPtEoY/h0MPwygeGYsVhJ57penBl1A15ZilK
3V5WohYLRGavpIWFUCxSEikXLPSk8DFcDlvTnJGR9NetgQJdxP9EpMYLr8RiCwJ4FBd0kC6vmgFI
3P9sDO1TAvZ0w0b+94hSUG69IyqOPOIUtu9hFa+Auf0k2yOOMJqbKpIE7xkrI6tqtkFf5aaQrX2L
QrXFv9Yclli5v//PL/t+dlBCux9ztcCaNEbnZyg/RUYjMrYKfMFPLd9NV4PWVqKFjKkwOl0sQfdb
bT1vAlMa9QwEsPkQPUXwNODZd7h0KhGJQeb/h0GtAlyG6ciMl0N7JqO2qMvT/BRWBqWrEmBMwqcE
7Cw5t58YUXIZjovOZTGMOrABMzY3RPXjDvA85FG2TO29AEEsvnTfM6aJzcF9S7Qm7+auii+h4vS5
wsafGrd07xb52YI9/zTRwZWpsFc8EmYwjEENGam9/1JtN6iPsdi/3mhDhh8VQBBUGbWYfny5QBT8
bWtUiC0j4mbTp+cujaOf7U19l+7OHH9vBh1vkXOlv7ATLWntPi1qiWVYarVUdpeKb18198fI5PR8
h5pHLm01f2cxzapKjHdsZehfhmOG7u0/xKaouF0kqkG/1/kPjnj7BlOK0eEjQgzuH3/WaoQia62l
Ty2nkHFPd7V4hJW8n6sKALSbdhQophvxmoS9/6d397X3i3fWY+kLK29E+dvLzUkS4Xg5+dgwSA8U
T6KoPswKvwepQ4w0/hwaobCnxYuj60vOhfcX3deIPJvAQVTgjKYJd7Zav5os0VpC7CxhcL5y2EQi
ji3DKPmgnMjeH9GhcURm1jLZfOVY0mss8+K0EPcQ1qTdM2FnrOKAci1Bi2CQfoHw1s0E52tXIsTq
niZzbKg7vY8/dI81TrrpTAL/EqcbGuOiVWEYt6TkuLi9YDXIcV3tVgyneraX9G1AXJyK0fR3BCI9
0ZlTJdK+XBGaVqFKZ81Xnw8jJlbMxMTOTYxqEHZRKXGLqf0te97rfAFi4p8ZUzhFyiPASb9wmC6C
jWhPLEgDSzcfZVp5qmTXeMe2HjfUW+UbUwSaYEKH9fWL69u0zXNdBPiUnbiJGc7P7KVke5vC2QRr
rqAWLyEFDs9AjOVNDrTVRfRKshHAYyK53ubwnHuC4ytieckAKqSUZ8wZTvbGrgrJvmaa64ewR3uH
B5kKbYC0LecdMfZ30iGjU/fnn2oyXTDKppPcy+3SAyyc14aqYy9hr+jvhFalEssOyV3dmtfQYWFA
Ap1+yg6zHJK1A7EwOJPobr/GMFw4htslKBJEhpjnI3cdh7e5pwN5QUa8wHHxy24eMs49VwC+ggts
6/WYLTnIDuV24EPBVpIxk+TCekPW6JYpQfw+aTpIOFPf62cKWvkwqn5lWFra5eNQXE+ateVFZQfj
MRSBowaYVnEJpyCTmCJAiPv6FY1YaOiK7PTdfyiU/eYBFmCX2A3+eyBbLcN60+3nEy9UG+T7NXYe
Ir1uXg1KE74SRSsrWqkXCbOI1MXw+Bo2DsFZ0XEkBgLINwIygVZzIDcRy/irlwnPsz4sRKDeuDy5
q9flXY1lZ3L8gIKad4PB5+EEFVk0kA9TOCgUIjr1Wz2IWswXUknHpoOSSdn6rZNIJJeSwnAdj5am
3LgWbjPsVU48WVvsUYb2VA3sT9EYMr+zIeAb3Jg1PDOAW94QXkx6vjK+B1mhJxSW8KpVWEqCNJVG
22QPLzJfp/jzQUJuOngXv6AZe03N5w5osz72kpGgrpjiyH3miO3WUV32UWSGio01WAvRL7gl1o0j
QJ64t98bX8FDXx7Un2KIQfZF94Q3m7Dsxo5NK21i1NlG06Hf3X8pjTnZoNbAtqPlEQ1FJXdeJrSv
Q3b6fnaHtVEff84B9vmIWTjeXYJtZhZwJnU41W2arwHS36jMKH9j23qOu5LYGSLoGaMpjx+/AqBs
SCztv1of8JNwpnW2XyVN9RUg9hAqeBAPNBJoeG2MTVfga4QoBJncGuwjBYVOO27h6gBxlTMH3y9h
1U0wBmY7EwtvMEKy9pgZjfzoMaJvQAYiTQwtZItWGjtlT/xBauM6jN9CT28x94VH/BvPuNOxl6tS
ZgkZr9kru4/TGBUKcGRBoKLpo7uR9e2hRF9K3OOm6vbtmAZV3nx7725HBAjDlig7wsoZp7F5RAW9
xYZR04crNp6XkiS7UTzEoWl051c1I4a96OX3SDPqRl1u/3Was7OBCo+wqHjmBp+7z28989wfDp/Z
TbnBkeTh/q6JtEq8v8HkDErX09Zsr65utEXneER6q/YuJ1BWgjnIrHisXPJu3TQMs1/xwnxRGDA6
whXvZTtaHERXbz3cBp3VfwnG1avysGaCyjOmGVsyPUtacK/3RFU8WFujfI6vWXuiyZwQ40UhiiL0
oWyzNmgl3DF7CWsFOq54HgoshT0ZPpDuIsdGWiD3Tf2sv+p7Lw04/gOUNEzog5n+v1/+L00iOsBx
qgZkFyjBuHrVhvt29+S7bjwzbDvENhCh2sCW053E6BwFEf/WRSbnywzo2Z37NB862W6C+CGhG65r
GQDm/F8YYk3ibwXgHLJRUQ3+vTVmsG3x0jUZYElU2X78pl0WPbly9PShzIAax5tpw1zIay9gznYU
252X/ejdo1hjDKws1Sedy2zF1uCJX+fT0OLE26CWaiZmsnYmcnNWlGKkFEe0/xqhiZ0JazlaFTIc
Wg5eEdywFOXetOjVbD2IZnYYbekN+Sf+vOZxDuHE2hDPSfy9/R6TMFJB4jcRlA8iwAxrn2zE1nN0
7yhaXXS83q+3FbAkFVhC9Ep78Iahpirlvy3q/rIxTjlQoowTPdB8gVYRSLyWnePl4YlyEIigKZ78
2/ViXJHX5TDKs9EZ0JpTmjMWBZ/FP6K73bdK0QAavtOnhp7QLCiFtyzInDXDNuxsk4DiCnfE9fpT
IYMyxGDhWpfzmJ9cHD13FwOXshB60oJebYSzwPzAICipj4NkMEKPr7pVYItPduNobg8Dgi7ZxqUi
bonYCZF8c8I9AcDiPyk2grR0ttSrtTZpcn3TcDgY48Cb9XcWItHAQqLhGL/0hrpov1p2sJnyZhFy
K4f8soxK5IZJZNttRylYT4eOiIzpqqG/yUAUCs7+1NNYN+i6qLR4VicSnwMqXY8IYyJ2R9JckPJ3
sRy2Iv2BjeANz8hKUoEVZtEp8YrG6UKCUw6w3/XMpS85Ww3TqUlKLNWP3q6rhEGHdbOIDAEZ6AcQ
akh/cw5EiDGHauHE4pfor9yHtD6yR55i2bk19qxlGH52as++ohAJ6qJjiuPwlC923rubUCeYDxH4
foXjMBZnGj/s9jODAtJd+N6KDL++avzpX/9CeLYpTqEZkrr03KV0XGKfJ2GcqfPOOWxfuYB62HNe
a4PSNEsYHZl+i9Q+Rb9YNkzFROyy5XXBXfFRoCTRyCwMeHdDFSNMwn3fsnRO1dZPemoVp4V+MDa7
HkH7DTUHtawBH6txrXOGxjkbfP1bCLFs9sdhsggqMrYllz4AbhXQmiYGmL/Aj5ru1uE3T8eRhnIl
NU5ym94tcK2EEIPhqHE2pfIyd/4o9Wo8h7nT0BvE6/ZdnzbrxFyiMsPuEYRL5BOVF1a+ENNUNAyZ
lbw68jxe4YbUFZL8L5MuVeGCsHVbJ1UaNgG0/uFPJNDGOmu51zEK3A74RsgySyiCc1q8hMoh7I24
LxZ1vVadqVcgT4mgddinVYEV+54yqkzLzHfqafE0Ri39W61CnnEsr20Efnj3pap6xRSktLQ9OOFZ
+NYa/ECburhBg5cqB0oZQWmDiqSqSmGuZ2ABXPmSMZ9T4cUvwxqqI/CT2gyk5KHwkxvCLH4irkra
g8mXdNq+xMnXB80JbN6v9nQEwxTwvv1pL+kRPy/gq3bidny/TWRkmqL/g+u/VmzfJ+oK6WA3FSvd
DO8E/oLqnDoMuXjLC0LRhGy0i8/XIGrB4kSHMh5IWkOwmILm84DmAqrIVvUK/hKm59BHqmRYWg3p
QRzRm/LC3HvDdrziQnw02+zvGshLVUmc2TvyAlvwLXbxuxneT709VmcgfDmshcuZMgzh3XbPB7rJ
YWWRCsvEsSAaf6dX3eAXzKHyTe5hrrylJNQXVPyfB8pjLfebH//xHxtD46bmUvipJ4mmSimGpVxm
TeV2ErojhHlFXNLHYHx5KtABl4aS62VeNIcyiwp4gVxMFbfXY1iLWhwXmYiWXi/RAKIsoqsygPJT
zxBV5GiTTlXqNUCIJj3VQ0Pwidzp7b94zi05kL0m1YLGkWAO+HPobzFazjyao4BKHifw2b072gXk
MyR3ync8wttCN1yUs3t2A4N4xfcDyw7pF4UNC1bt4h0cepSoONT7+9UIWLwoRwD1npCMr9DuGs2P
c+pfwtYrn2PP4fQTddtUkC5Z0bFUnoOPEkJKVTKE3bT6jUmSEAgBmC90n5M87GK+O7KyCc+r3Ul/
Qh93XBSZZMd+Y20lZKw1I8JiCEP3+SeeORRGapmaPV9Iznu7Oa3E2Lx5Bf2iqM8EPtCnzaflEvwt
B+JPn2ASFrMIv1m3hE7eJnES+0cRa/0fEqzY7rius08BwfVwtNb3xpFxH7Ojajrx5rEAmNVEp9uf
e/5u0E1ht7La7LeTVtxk9Gl1V8ZQ1/CmKWfhyf9qtMeHHR9UBtnCstBuA9nmqnacRxF9pC7MS9j+
go0nkK8hHBYxtOh7XuyW2jRXUnsHhpUpzznJiZtDW0/4jt2GsJx72A9fV1TUCt1YAahPagrxNFBS
93j2Ub/c9C4Xt1mOuE4oSZj3ZTKZ1XjOrdk0rhzYpsxn7j6Cd+WqKRvd+oCNWzUq765yY5UrotTq
DaMHkrK8jvYOxuOf9X2fGSRDN0QKit4+bXzMy+ysaKxYKNsTtQNo1eYr2E+AUVdo+2Ier49M95Mc
T9KUBrugVW2z9LTszOzGDsXGH38supBNaUo8YMdGymGgDx7a4PpB8X2SJi9CicElEKeJDQFjJKy7
Klt2nDAvlU0LaEat3i5Q0xWQfc8oHCqmigwOCbzmLCzdk08Y3IEWGwNBosnwo7OZboC5SmvcH1N0
b49Ew4TO6N+2TAQsmebg/Bji2IxP+w869UOil1/x6Szi9EWv3yy7lpfVbMI+CsJLqFOgiQgZ45ow
ubz+/Qsl5Rx+wq5hNciap3MtXTWnAHBlX7MDD96W3dvjo9qDYPrAqhZ/7lnYmgwSsTJjpqARyOfZ
78o9JGrPe1ffb3frZtZ5LyZkBxMkyRYiT5dmKu/hviBGuizzRUOs6y0CAgfwcc+WWLi2ZhAgxvvX
c/dj+1jRCte+WqebWXN3FqL9qty8j6LeWWI/ZK3UQqMQmLWoV52sD6IDBCGaBpSzhlpAigIjWljL
WaPc4gmKfhwizcZvHw1AgkoZvKG39ywnk0AFtZxELISrVwqlnN/nvOjeDTvTseuyGfgfVkLRkq0u
kWLHBCYZMI0X0lx5jr/09fz4pY3vieQcT4zURizQiuuS1eJUV1aWVYgq6i+/4TUFQmYeAlivT9K5
vds3vv3H1/CPwoc2xSF7UtSV/vJ9uLwBDLhH+oMvIm3iC34HSF7JJkvSm89UHYRsnvjnCzOjY5n8
neNvTdTr11CXnTub8PYCKktZu3ZSa/lGKWgbfJzBBIJBSeYWcgnG+iPqyNfmznYHv1OHwcdpPHXl
vQB0Afn+GhtZV6jd42fWO+Qtc/hdoYKw9Pj4Ls+RVJtEPoaqnHajA2FgCtO+fYjYBIGbf30EMpdK
NqhaShpJvKYDH/ywE7Wd/vtzzmwcly4lN7EizTgpHP0F9gBAIox2e8v0WcPlYPk7X2VLoNT2v1uj
Jc4Jdpl9pjpkxVZOaUcDdldwVqGD0dMFS0frMfxqzZlCYV4E4e9Lw1mRL4BFm11GLbYblw27o6UE
qD5dzOgPcgC36xbJXA30CVy/2jU0Dv6hSYDS2ciKNxxIpN88HoVV4FS1kerC4kdMrw7hRH5A9PB8
p/r+5tyj0PNLqagtEWBY5Y0wySR+Oo5p6iB2B8gSABOpAL6iE7r4Db3oyf9A2j0NAW1G04/gabqm
K8lP5JaQBibd+8Kk+QKCveixr9E4wzZQhukMcFsHykED9Qy7NwfF86bTgpzPSdvt3BV4wYjTWe9W
OW5SjmXxidUVRMUmRvea0uejVUEKpFJQuzP3wBmIMj7lPvPNFathRCUpyDFTI9y4+Ns8HLdJcAsa
w1mRFjD3t8Xpwr5jFTWnsU+Iln+19ADQ17O2VynP3kzoqNfSWX26GxhAqa0BjlfQY26lgXAfB59J
vl6TprQWi9khIJuLaRP5p0T/5Zb6HifK+CbVNs0CL6fdyCiJdZejqAXKdn+19GgEwwMG8riDXPMx
7jJIFaDJdtAhlzGgy3ppxP5//N14+3HpQRdCwNpOQRajGlBIwSMHXJZS2pGSBrAhMFyPqgzxBxa7
VcLIxGvjImC6ZQotCMiUW3vn26vyQk8Rm278yMWC4NBGQEtcSZBzvhSu0jEBDxD+obRubOLTPBCM
v3X7eeaDsAU2LzqY34WAc2J9cvqooYt3wXHrHxJ/E6C85Vs9X56unmz9Md/JDTwt8hB2mfn4Opfh
EX6MqDiscnE5jo+v3kI74di9Ec0PSBGO7ug+vNeSeSVTJMmTBIE3Wn2i9XBJxbSPH2oHc/zcIDRl
SbxFSj6KuGlRMMwhkbiEUhmI87nasISpdtivJbekDDMF9O/Rh8ITWaB8RSSI+LZ1M5qfgRQNbnAF
H+2ol07gGTzVZXpN0ZxhY02H3RAfLdkjYlwSOunIVw3STr5h0BkG1YvkyYHzWoTX3/QoC2GdcFnn
YF4YpMJxiChjbxSU+exaT9B4bLspBQdri3UoN5jGpYej3sHmm+sZRK9ZPd+T1danMBzL6lWc2IeF
rwnw0pOqAaNf1oLki6cVwWaqmyxIfXSz77WLy18Kv7ZJZE8JGYRXhpgvbBlCkImQQt3oHH7GmmgQ
kNsqTFjuqNTZNDe7wDIs4cNSmQn0KO1qABkde5iU+SDt5YOUUR0wwbkYqfSwtY/xxCUXHQFO+XF/
TVWrHGNm1pGbVtMpQ5ndWL5RnKu/U6Pt4NC93/+8g9owji6wBFyr15ACeBYMDqojidq2TDPBv2YM
939Me98OnTdP7nMcwv2Xy4PWsC8Qm39zzq1RyUcxUP53PHvZ6zk2lxAxVfGwihVXshUaQG0PJR88
1ShgoFLMxcg6a+0YWVj/ggcMC14z0MEP5a1jbBE69s2uQJUM+1HOMAckvYLGNlq789noa/0k/5IT
ttIYS0uHHyHSq9mlflmtqBcTRF/cLC4RVWzoGrhQ3uZec4Xy9MsFunFmHEvXDxWZYN3cOMgBjJab
YpV/fD4XZNsaaRoGfF270hN/ljVFRMkfiqNvFhWzBKdyPpvUCipm9mwa95tR7ZroSRgqOH8ouAFz
OaM4j3r6zQquk/DTToDupOqN2JsrieEAQ3cKRud5VOpurAVd6mTV1/mFJj7Dx3f3S6RKTE80jzEW
CWIUrTjwjlnoC/RXykm4djag2NT/jF4y9hF+bzqok9fTS+2mk07K65HJjqkFi/CF5SRSCNf+SI9J
GXv1O8E/YtpZZk3YAvRA+iG4U8X0fhlmVICeBP2DqCDJq2/8QJJ2NZtOWG0UWTMbNuMBngMaFSWm
pxRiGn/4nRy4iAT5GOQj94sz5EMXr44mROx8hlwVE9pUdT7PU/lcjQ9Fi3idR0ffftkIxQYJENh4
+ODZhcbqkSXpu3yZIG+FUUDzZZaLtQDJZAEXTfW9Gewshk0kQH7V84yWyZXUwhDT/96sY8UTrCXL
uUAVZ/AexUMp5DhL6MwXWKT/Ny4UZrAw99qkkGrbJwYLb4yPAu6OSKlch+dGSjtM5Qs7VN2JXWot
WefpF5o46MJafFNnV84PEnKRETM8nhmM+4Z86Ro9+741eTeYgOzH9p74Yw2LJCxYy7YpbEc5K+nj
WOsxvwImMAaaIYDNOpiSz6wdHE+SH7IJ+62uAqnRgSGbBnSp8J6ZAvVbfplBT14KqIxZD5i8T1Zl
b7uOCkMbG442+GKFXdvdaeujJIFU8wPathP2li89OW+uIyEIjClnFIOJP5FqsvETOn7JGpUeaRtY
758cykciiD+7Y/gWjzykIofHu2vamAj0iw4EYIEkjwqIDGyziu35GxeFittSFKNHTzXKsy8Ra9fy
5RVfJHEySk/R325zz6h36CSnhS0jNDSBclFON+FSMtIvxIF559iLSuce8ilBP8TsM6kez/+wQPYw
Um87Ons+ZKuXGMLcOM9ltc8gLfa4k5ogx/kIAIiNp3SJJgaPq+zz3cv2YHIlV5gH/Z0YpfxyUhCn
lY+AvznpptN/wbsvdgr7vXQLulrmIoouAIuqVZmGssdQikvUF5pnHiOgCh7sZjYDu0vPzs4/RXsk
TgEIbYL6+CABnqeQy9UVZnJVIgSWzptlIrjnzavmdeogXuxyYH/cCTMg+3js5QVvMlsEUSogjNj5
n7ikEM8VJARVEDvUtLJ7t/Oro/OTOb5ovMUtxkRkpH/Aa0xwRjjLYI1V5M4Bw8VfS15CgMBMHP06
kgoFGleiic4DDgg9/gYZC5tYB9+eRmdQrUJd6MeHAT4OC8PEPU1e01bxuJe8ajm82iorXdX3tOQf
2vJordMRjf5QFCDOTMvRyOe6bHtBKY9taMkrUM3wX0DEcz14jT8CwAzgN3AG2O/L1yqXQ+bjUFLq
DZtcOlg74MI9XZzY2xo5k0zeBCds3sL6m1RFM/jgThLv/VAJKg0DxzAc6vRa+DA6e8BK2arCcqze
L+Jh8R5pXSsahoiZTkYNGQLTIEr9CspTFcwY6bInfSv7cz3F8FYPsnslgvHss8Ff1N0lVApBtYHF
fka3CtBwoUI38NUg6/L6yMqn5AC+y/K8Q2wcfuerhG2ZKafAhuUf+0DZ/cW+mazfnWyL5quxJpRB
eFxljxvBxbmsZlTJ6pR6SotruVaHC3iGsLctbizOfz74OXwnoV1I2ns2eUZaRi91d06YL35D+GXS
3Z5z1dl9iIa62+KsgZHiARqRqwHJpUMsKpXUdLTGJj98y/u1m4JwyGQraL575sXIkq6UvXLE3sPi
W+X0WnczjPqOAcygXG49GUJehM1xCYhgbMuxPlZUBuknz90H/euxAsP0BU/uxePzU1q1udqeQR4e
251/U73ejK76mwsXwmliYh1rR8T+aAo/2/O2GjAa9OCL27IOxA1DmfJiIGe+KUKD8Og+onMsCVjI
rkN7R8JwBpRIV5SApHLfuYagw6bql5sqW6K4Mylw3B2eoR5Ega3SAHalBrJnsFE20Wvpnt3Q+mzy
gsHlIWZIAU4KyVXjBLEll3Ul1WoY7fMq48wf/8tSqMcg6S//TukybfxX5jM0x/ZRBxP2S6HkNmK9
T+p7lyg2AbcJZRisVv1uZcuvdD9mESPD5FcY5SKY7eS+IJA3poxZ2uGUWLeRTss3AKL2fAlNsiCn
iQ6MVXchTsNemQqYldVkVXvQb6aztqrMRW/VNy2jCRYndTb0CdL+O6dxZngNzsxHYBhlQALmCXle
+U69y2d0egJCeczSWFhQk9ChVP7C9zkuLXez8brkTSu9rzHpx4x/MACxJTpIzrNYvtVjFSAYEfVT
T9jpv0Y/Iz7FYvUBEF/Z2GvmqhkcgiiH1fvziDCaL41N/oessSm5ClCGlSiVipMtqL6U4Pw03Jvk
KsCqyN7ECEa8dbk/sKuFi49viMkKeSeN+12yGwtO46pZgPVDAU2/JcwOHLkrOzH45hlVPCkEyyne
G49XuIJr7Ts1eoVal/kxwrQsYxFrgRiWhdCKAL2WYkY3mUeu81kuZNaSDeXepnue393p3RuDyzbu
m2u23K4P3L5pOqW1j97V/ICiEPbp3Xtu82kIaWfXOkpsAQTIbB4oRkdiqC1tmVEnwyW9QR1VqAhY
OIeMLC6v7s+D9Aj7Ceuk8RkEu87k/x+sFNya9H+oiHTyh0O/+IeMsOvh4PKQJZjgR14nAPTJ6C2Z
zZbS+LuxzsV3BSzvNcW7RqNu7+O2QlClkIO7WlagLqO+Tlt3L/PXmFmbqwixlCpwvtSNl/HDx9Cg
572NdUTIaKbEsMOcVU2Sv/CJ49DedjVi4zOeoY2sNdHqDGyHYjCEIurQy7LkDbRqvF4cvm8yKgf2
O/7am8f+ZYUYXiBIkmBq4/73cDowKR5Z6mLGs6/Iaurf/kr6ddV+3Ve/Il4cMsSGwb7dOMGqMhFH
1VFPEJXj9q+dVRkBSSm9NmyWwtjpgM0olRvUhxGttUsybuBTL+su+5ZmMfioRb2wW+MTyXdY3k54
aasXh9/3V7C77bWAyfIhc99c1PMrVQ6aavP3DWb9B0inkATQ73kb7aVsr0KU7ItfbNOykoxe+0l+
0Ti8z9WyO+GKjQViajmikEtlT99+Mksc90G+CjYCU8u1f70actWvubFeNikXUMvsYoEH69Chi2Hx
/BO3NEbejqgvHNIPpnBDzndsyCt4fxz5lkzzDCygkhnS83yD+bpfO/FsJg64ug+XAhq4rkM7SNxi
UHnTqa9nS+p9mB0GgRtME7dtYvdVJSxtMUISWCTzI+lSj8h+HonFx3eHrzvEyU3Hjf8nDaPDy/td
/KxAo9UfdpSzz7jW8irOCQ6LtUzNyK6G+4SlBye6cx8OGWDsKsxQ1kRcW8OLm6RijcfyrE23mNJg
VYloCMuVUo1Z3P/4xEwIIMASLFyQ5pVxAFF5GyuDgNpLoBuZ+TQ0z6Yvbb59A84XrThOMeYLkKu/
mxvzo19ed08SdU38+BWdthFxhiiomDnmBBq9mCZRApv5hGF0UJCmzzDQXuxf1ZnktQwOYg7e4CB2
QKbfg6B6QRHpwjzG7yP+1QBjspT4IlMHI08ZiFOXbo7CUBcQcoAcOJQcvSA8nLzcJNUEptFO216i
bUbco9B1HN4wWMA35HbuU+yg4tHkDAh6oF/xAzvOtUCUo0NTTU7B8WdHfsP11pf4s6zY5KaTcyfX
S8+BOyEJWId+zTp26aYdevAHTtwdaQiOLIEF7WkNZD2FZtZOMk07CsfHP0SXCB28VgT+X8TEf/p3
HXVdH4iNBgNQ1vdIppDKI2N0JZ/fzIoEacFTzlAz6yPgVZ7Pqdn1OOfl7SFugqf1knN55HJtIiYB
KttE5OB69gAp0oJQsyq3VhjDIrO6wYkBvYjuCFqj2g3/nbHPQL85d1pDA/b5cewGF/GLQhyFRGuy
lMEiIeYpxL8IOhEbDTHWOi0i5CD/+Nipt/5rnnoYnSbjLm3MptW7sryQecNYZ5fFmyKsWunM0DVC
z+OD+ZQnG+lkaSU3MePAA6hEKGHSLAo2bSciCPScyhHOIRRLQETQVbFIq3lJAVdMnD51JoQfqRPT
nkICCdrYMDKa+nFP1ocuUCS8JF1dyDkXLG+I81HlXazbwt342D+SbeunP5nTdaxUBf/N5z1iMrYl
z/giQwcUPWM97H6YK56/8tOzl7EEsOCiQ0xML6j6H64/hQ9pcbrPMKgE4NNcm6MHco62dZhZy6a5
OOfUxxEgDq7svp5pFFt6++782c3Id9OzjoPJbR2r271AJw/FmpW8u04cHijqayvBvsxS8YegGm5q
w4ZgXJw7AJTohV8tKC5S5jDAZC1i3mKr35ajmuNcw8YxoGJB8PK+L/TO4bT0oJCw83Mqao/10gMk
iH3T8U9DHHSCitreLAoerjKEFRgBnJdh3T7MMKzUmWAqiwBUUdWSqnTBTiptALTX670dJjA0II6R
Xsmco3OTTvZKO/+cyFqX/5puHVynn7m7K7ogz45A/fJf2MtHhFSiqQET99+CtdCko9ITsYMY4LHV
C9FnEHDGJqpDWB6RZ3yBs/HSG/MUhgmEIZULoBrvErEmkwq2llIELsu037UIlytOgAKf+qZv/KJs
W0l/wRsNUTOHlYUGmL3usgkXxAshKpO1S4Ow36yT36oGKRG3cRUvsjyz0mQxawuImgokXc8bsHuo
GGip3MDDoY2QBdeyEcUPFekL3O4JPnD0idygjAT6POtwFoRy+nkNUDcixPecaKH3+HgQM30sRPER
k4fhGAQJX5t4XuZwNAFkQ+88nA3AiqGlY7uGuEvqxpeYw8iVHfHLHePE6yAuwe8QFYDORMSLZiA6
TXsQb0QUm7Ddrl8Pa7aMKjZok9YD0+ztL8c1v++TVZuC20ILOrmPPbemz5f0AoiI0vpxkAgIwxHC
rtHYwE/rut136TFcKOca9R2aS//v5o25bF+fL04Ysg2hSO+CXf6nBrkxwmn4aQZfPn938UCnt8W3
dKkoQV+L7xZrygigMdqDRN/UuPf5IXqyCue+CQD/wvupZgRDfVOsEIbeJc7GzasvGu/Em4hRk2eo
LK56voSljXb/BRlNTP0xC2AixaXDg41Hnp97kcHauHp4ysRobCaukcpx6FMGehMlUOmxam7wXERe
6lQzSfEez6Pv0jNVQThDrl508T5FfkPbz9fQcL866tCylGS3+pg24MY0wsgoEx5oLetQ0ltWHnss
Z+foMOkyAiZMwhbxeN0gCdMUE0TZyL252+75FNxrZI84d89wTI5B52+i37iw6m9lyZKCPliMDjeS
ZzsV+lcV0CEu+03MpIWaoGgCPrVx8jeUgefJpoQ2tAfUgMD7wOnnt6Kbu1mhEvYhQsEsxfNI9/Er
dTygdvAaAyccJpZq19klQ+PGxpBRK3TBFdnYFIeaxOwEyBMNHEpTQ0OjPwd8vKU8TY0BA5AoT8rN
eAFtaKqOVOBumvLe+NKIBBaRfIvkfYQdE/7n0BtJhhWc+fenW3VJfuR9YavIva9RnlsHSii1ThAl
Ina9Kab9Gf+5W+BZvFIv47EiER4d81eUMXpQrU2wAt9HJfDPf6CzKHF7SaKFHQPfWuJ41O/zYCOv
erXc3nbCxunZzf/4UUT6PWz7WxWt/asrcfDBNbTzwfE2yHMLyJkswOEdB0kD8DSwxd/tX5l1sRxv
pDlvYuqa5z8ICwMO38O6sLUDZfEy3RuxBCoMmnfcvNZebG9Lvzds03hmEYHtcbI6PV5i4fYu/ub7
5Tu2mM9266R7sntJ0Fz4NkB9y0QG+37VUi+M1rgHdztNn8P8TJBVS7OvYAVNkk+YlVpBCF4flaWi
PcbfLEszaVjR/XBXtav3vkKVWes+cmZ/ml+7z32h83Vr955nf598WAVVbjFSweAK/V0DpY4jz3sV
yo0qQ63FuZGHB5BzfOA9H/oSUfEc0Nigzn+CykHkVG60/6v8GLtG8kl+fR85AJyqZ+hOgGktSrsw
HDwrHHjnZ/jesc9t5lCL308Waie5OP7q8KEZIEpGzQYBvKJjKqnkzl8a4csYvpKGa8x1KLR81YL2
yWpxuDABgGHGn826aiNwZKVQDFxM4ViFltDqe9LvkVwg2ep9L52FrXSDIlXsJTJnWuE+djcJUdNb
tYzinfupsnRe1ArR2wnexuKM9650NTIzWxAj7mBe5kfMzyojLep0vPa/U2f+k/aO9IsFAhuuL4Mq
oWgESe7FIIOvD7EZZW9OQjw6/kivc76hQfkkPSB40vt6TTSqRVocDphQmZgRjCnv0HBaw/KovrC4
K/Y/o6JkWYUbn2scVoGlBauVBzfKxK5QaoQUtMZ9ZbRv5kqcSutqtqg5icY/M5AU748Dn/7t19in
/qdNe7vI4w9xWAgCKv11EzmPfY645oft3vsD+Vf5Llcfu9cxuxyooY24QPFH6uygEUXGKI5jZqu0
3X/S1eFPrKVhFOdrqNHw7NKatc7ZHOsvSfOQOREraR4zk8dpz2tf9xewsZnuwr2DK6pwC3SxDM3o
ae/AuLsbfoffgi49Zjm//bCdwwt1w7DmA70i4Kc6xQkx6b5D7BsPL/m0zI7SJJzRSC48rzDRU8Vi
ZEcS7HjJ6ndkXx/SMz4vK98lDHmiZ3L0oI60XSt9ESrxt3sYkcVIagGz9g6GPxnpJNvPb2qSAiUl
Sox/ttPNgdPIoIB9Ne2dyCi/RKAr0uxzBJCrNIEbqaVzm8+GE1JImEgWuef3RZlyvcBpUJjUtPq2
XNmeG2dxRCp4nMflQ7Q8RdOE216r4kSdtzoPZjyjT729GmVxKI91MuWzRoSlTyRQ9ZesxWYbIty3
G2aB1vj9O07ggMSQFlhy+0bXsgvXWvK7EdixAQvZdP0xhRu6cVWCpckyLIy6UuaSK6UoT7H1jqS2
amD3uJeS2oCdHNpk5DJlaDV/BG04kSIQ16ChPxO180yzKkE3a/cOnkqjeUHk0XvIEsCE61GKNKJ2
Hpsk5ClwHfpAbbPMhIw1Wd0312mCojleTDrZ7dwGK2oQ+U3VjitW12D9pAqq/RQUoO2yLfB6hJLL
j69bvXhHtX2st/0CwVAyYF1zZpG+g4amIkr8Fm7Q3muu6+093FJoLU7U+iTIvqN2A+KnuR4kLVmF
zHZNH1hTqyt28IapX0SEt3B/EHQDNgC6b22nls276GmNI6CWzMumVOV9BBNlHikJPSnIJCB4nG0F
hW8Z17vxWepdWlzEa0sNwbd+OWYsAgdvIAMzm2XMUinFldYCG2qwES/6AYjW16f1onHbYYGE/J0V
/CQ6Y7A99sV5VYx8cWx+h1DYKSyyROJZKzXF7pszzi12FTPEi1OKKwbMoh1KMNBj2Cho9cWxaNdd
1LC51ghJ+tbx8jmuHIgpEXlL9mjruYiDt7r9WCmfX0PkAhTwD/negW8655d8nvvaAADEBAW0L6tV
VuhoHbRFF0z1D0jnngQ6vDku9Kq2aJ8A9NOmYe6wwBEHX4H2oVaXZZ6BfcGmwEMN4NNdvgFcFe2z
MGVPLJgyGksRn2Ymj/8Ax7RMIgF8w06z3oYTPaqfx+ncKmyGczTbR6px7mr+0Yio4tt7b1AttK0Y
dBNHLeP0BnYttZjDb1mB+dvBUPPHJSJs4zVq2FzMUJct7HH4otNANINbHVq3VJT5CxWSySJjA8S2
KADRHkEygI2oZEo3KeSbDJ50uukpYOWCI+lfdllI6YZx7CC57cremG4FbyF40MxmgaQox/57tcOF
1CEhvyEGCitYmFINdKAsOW0gznEQe0RYnqfLMzITO8mRFjMR0CW9l56BBxJaX1m0ftwzeJ96J+HR
gRTJFgXQhm1SQU8E+umyqU/RQqsZdpo94Z/GuGwFcnsbrxrsYES/jOhkJ/QtruiaCC+VITOJN798
7uc76SJrlYI8orJPP5oc75lZlzxI6YS5nZxCApNfFlg8tlXMx4nJYT5zBHR/Ywb1+PUjMCAUUVyr
BwyHiELYmnO/Jlgu+nvfBVvrEeruvO+1w/iYZnDbJ3y0mHE/2al5hU6/IzXEwi52VsMxum6C6UE7
ANmuM5ZwyIcU5oyv90D0ySQxQ0LOdVRErwIJwDup0BFEVcqlaAteohl9++xzjWnPSE1CXqzfVC4K
lJ1XJ+Lddh5Uvz0crpehkZa254VkYXBvoAcs+yzfqIQVxLo7BChVKWHk3IN0MBxFbrjM05TJtSaW
fYnIlp/RTzKeiOWLhfTNT+hyZzlRn1arN6yZUoTkWy9kB/fSyKEYKuMI8Kb1wGTX/Ty6QL7Et77g
I1o5kcvoif+k1C0++1FcvfYnYF1VbyMxwwsussFgxNHSKvC97wynik2ruwWc26r0HZ1a+Y7sXF1t
CO2bgDSxODhpMHNaOcQ4+e3oiVU1nJ99Z+DxBrO2+WOUyK76qq9dFqJZx1MHNjQae4dMhHB/IGfL
FgDY1knong+3Eg7m/Q03b0iVpBntF4V225x04pX1uIn25K9SIu9Lsjb4MdY/ZLAFtN6Nkdy32acH
J3nOZr0Us1hQQHTcGhEUvnPXtFbCOrwvNQOBimp2iJFZaTvyFQfL8848rfm48b41CXne/6Bxoh8D
yWf3QTJBcyebniBARsVd8NGPhpcZbGxBgrEu20MlZ0yTHqaX4MFetsCpfYAILPCq1sga/gDQbwWK
WazD2lFXVpW4EuZhP5YgC8kOFNIaSkKqlBIqVVLE44XINDSbFbB57eKLPgVzKIO/ytu2k57yq9Fi
R8qo7w8wMx+BygBx6an+uXp4oRX29aHFHR40UbGDsCscKrMbcqYx8z8vL8ArVrrVAf4f+9Mf4BQD
EgE/Kw1brFC/GvZZWf0PBQzmyX0XCA676S5xgW1eiYnQcja5OfqKziG5fSrBxtBQGCljsHuI6/Vm
Xl/MsYANogG8D15jOVw7Uq9VU1EvCOlylEd8TR+ISIQVtNP3fZWWgA93nDQVvujAdVmvqkDVJlqX
UfsZlqHRii9LFEhdLIiawOzNZrb7MU6p0AKD6lNlwk24E8XiQjjaJ19ttZPpDGhZRTNNER8AP1Hs
g8Lk7OJxORFzQKmuymSsH3krUNo1scgK7INMVT0FC3A+FagsKWU6DMxL6gK+sVvCVpuDyzVP60PF
IJhuHyajEGz7btPHDvrjWbTM6Aq7ofmbkZZz/PPk3qHvd23QvIM14rHsNE/4KqJLa3Ci0wUMKId8
sFt+frCtjWa8tMF5M8zdfG7SZyX2EJ2zdETPrK2pWasKpvnKKEbJBqUKKqYVr9uuBBZ7B2i0vNJA
VcZndbAgE26e2Pc6jiABe0IuONzvmitFnlLdcn/jiFMKahhW2xnauruDyujR0fA3/U+Bri8WRQhi
elxlbz51GDqgkY+67O61KtgKqkguoJPGS02xNG8jPjIzgObqlU2SOlUMFXFI8EgoBSFfQYqWa3M4
3JnGfG6hi9NKqzmmIWRyd5j0ofFtbp8bt+MhO2kar3yBHWlcQLXwLcmQ5RwG/7tFnC2lzVnnQ5LH
MmKojEqpuAqIUZFMlAoMNWuE6PQ6PwuJtRvvzVFwOV5Oey1MrDZJPsth1NB6trMNd9Tm7PC3VpTA
4QwB3bXY0pZuvnYyCEtEcdf3vFW2gSrkEqILAWLzWFTDfIPtGIAr1fZdL0AFnmxVCHemPgzX85yY
Lx+uxgvJw1583iqO3c/8lIoGQep+MhKL9zF95gcgHjc5JJKI05M6+5R5OlmpSVJF5ID6vvDpxm1w
taAqQy7o0fUAdiCFx7x4twVD9gWLEEkn0k3BHTAmpRJbZOgtr5EzQUFUoEoztlLhcKlbTfw65+z5
qtNVzh2a7IQ/xFSPp19GXjLh4x9H54gSgjXnnvFpHRsh3CyKB/6KsZx+TbKpMrR/pwMD0O6lRTTD
WN1HwrsXcBJuFOnkKgx/miCyt3+B6E+PwdEcB9+eUeXUZk2uPimdl5zLoFk6DtTgR9qM68j2aiwn
7XB7ZeLV/1oCInaA1wDS759jLRa5Ue2NHNB8ZgFgVlJfQiGMQhIih/Er9chNuWFlI15rYTg+esCr
TR0EKrSkijqZ25XLj+FXfgT/YFdByf9XtKPoz22VT55wgP4OnnGrnzub3NgGtRzc1NfpCKSy+vCN
PDoAcYeHPiGv9oBVaj6nYtFVXng0PRps1PjUl1unmMCasxljASvU67AfqueMvY+r3U11nRM9RR+G
h7IWye8dEWNuQsZA7soxt0movyhPhEUYFhJms5cLBx2q1XeobcxX5U81efPk2migK4WYCvoxZA2C
FXZiIokh9gU6fNVLi7TX+sfA/KFQstKCFQEyyHLE1y3aokQP8N30WbMBTxprx1DkjVTzIDmzYEeF
wZHZADXO8macbZxkTHu9sPKpc9zNAo2PQdATGjdpJPhEIipMLFcTCfIelJu7zlYALRYi2hg+orr2
BkQmabsUy8mTw0S1L63gfB1TMJNAb0+43SsZscYEyzOJburEiWTEKu651OnfL1Al94EvAK7IGd3K
ILcmPNgwevpA7N1tVQds8BLZmgi3WfhK9RvRc200cOvGDu2mRWW1gEmFXtMjN5a94207wQSOaId9
2rN75t8Jr6Shb4GY9UtPinNVkrVJfSrvFkFdCRhOrJDrvUSWMH+x1cUqDY/d9tibN8OLjpSznY7Z
l2Vet1Cmn2FRXHHEkGYPgg0bL/qwYA3trhQLIG49AX+3A30pRQeClTfkfXav2dkSTzk71TIsYOAl
38jTbZZcxK1j3T2qQeZHpeZbqVk+jFTK5F6cwzGEPXpFuWcTwvDKgwrAcT/hWCCxLVuqtlXP8/c1
72TKaZYjaA5ozMqJkKUwvcU/Bix+5G77QY0K6BVbbxAC1Pp8cYZ6BTYsEcWUzFyPw3fNsfLYApNR
07NEg31hLBs7FlJO2EnPzgnu084a/sMMu+NSoyr4qbwtoWjzkDOTIYMDvDICup+hDSKkds8Q+st6
MApqiN29FIsv6vhYEKs/znk12GLTCVnvHOoC2HqyQTm1xoeI2+M19QNN7SlcjJdUY8KuDEaE7mLo
N+t74uk2dc72hOO/aXNPZA9WBLBSR5oyv7D6GZElst60eOxG8UGhN9tQ2+lsbFDiHWdMAGrm8wGq
vzNRlJDd/vQ9egX+tUzDWuCiuDZq1lVj6UKj34LNkFxDng6tAzYeYk15yyAbWVTZM+PN9JX2dQDf
z10ZAXxxDDXo7Qz/DRJVvfnKNZK9SkvATYC6TinT0YLnB6EwIlAa5VZBcUAT0DZ+zxJgZKbD20dc
zeMccmwbjt4rjKXbb0AMXvJOysy2HMr2JzMLT0O9B9iPJL2zHeWmlwdJwuhjrvJ0nmo1uaJHT13f
59ljd8d07Gw1zUGoucXNb0MsPudqsp7UfKFN6OFBRv8mTq0iZlbkR0r7o3xmeOXu+Orw56A7gwLl
KsHTNT7NwE5hFES5g5qublIbZlKv8CzfvT4UOYvHXN7XuaUdQM/rknSObPvQ+nB1TqWLNCggJtqd
h8XtFnysSr/ydSrOIxRD+9xvVN6fs8Ev/15gWosSO7wCqDs38I6Dqq9A9126EToNRoLJXvN0VaZX
BqixqjwxzG3cWdGa3jfGx8VejiEyaxY9Mq68nZT4+gIKPOVArhgRfL64rHD1INGBGE8/9NoDSt4q
knlhflW3+xIMXmKF+wlAFZImKcFV8osfrDtzayPTfIJkyUnta/9lMlE5++kONJ0BG+hHngHsAxtJ
BulnCJSADXcD0Hu8SjWla/0JMrreE5xqI2PgYkqIIttu+JFAi8d45tQ7wZFat/xlOkjRI825hjrn
YSQadfbhZAppbk+qMcWSyHE33gTUbphxa0xeuv8JGia8djXy6nfxa/5BqbW+f19lNPiVL0wOnNin
WmtoaAhJ2bX37BeC2q+y2mXb1P3dUgnAqqPYfzwvmAlXhSQp3WMdRVDTIwv1MyDWjjWW37usc9KZ
86CcOJMsbTU0Ftr6fJVd38IetA1X82ir8NPaLOQ23TdrLqNYkepCJiFrlIZojBS43WN+wELlEIAa
ZgwxFbP8bd0YyrVd3PxqFASo7ZQ29uwJqoi2SjZM+cQYqT3nf2bwDIHpIrz0wAM+fQFH4f2Ab28L
Dh1cO0qYOCLVeaEs2pEiPJvmX4YDwMfHFHpEX7t7WGlkQOqTHk0z/81c9NA3Nh6J5qpmXGyvqf0t
bGdSkrYJT/oUgCt/QKzOJcDkDLm7Z6pWcUNCc/P5fluRaXVI9cmxsrgYE4mKXenOxQf5/JZKpJHm
0BOY53Rx9BzC2kqMLpRDBFdzwaFiyWtHCoWj6EMHxeDh/73QKImZhON/s6GG3DmyZ6kll64E90jJ
NG8MVNxMG+iisXeneOD1HgOPJ5pGun08npZEJ69Bf+x/FIor7+SKFgRIbPMIcXmiHChMllT6rN36
lSNQdE+e/0gYl8U10vDBddvkEKpeEbEHNz4OcmUMaBqce0uSVdibWI7B2gZJKkaCbq+Vud6iHjpt
UOZJYL1IK6HNOgjh6xvriRTELgK9fb9uDazsOHaD8tJzB9jV9t1URWhQwXvjfNtT9UFoZf5NN9bK
psWLoSnqG72ocOyW4SnVLd3a08IU0FHXsEGvy2uMZXzElwPboRsXFGFcMF7xmD8/67saOeqc0zOF
zLjnKOpkBVtxcvaUakI/wgaGP+c0TalE08GgTzq/DhgzZF3yu+hhD90y1cZ3suTSpkFfOOVslP7o
l6KSu9rqPPuD1gV+f1pMDfJOBD/ZnCPcoQNFjgkOp7LeuoABdhhYevdP3p4aOal4XI48ICI8BSxZ
p3Axluh/7lE4nsgVB1OKZ8ARm6LK367l6pcUQMbhnxV4mPKB09MnGiXX4I0hlIuOsZb9MZzZk5tU
/KqZzQxySTqb8rsQWgSq/8HsUYEmm8+RE7Fr5cCO2GpBxhxp8x1S0O6s9WAgIbo98Rl/eOytS0cz
exePH2XK3x6Uwhj32ebV9iCgYO4oCfXqVCNDFnU+KssU3vWDPjehvdxMSEa5jtzynYUBKueqQobl
leCOa1a03tFGa9ZRX7zCYkcPOWLaPu3WMTBaHG6xopvYDXCSqS/arAm1v5urAI0YdRen3u9yKXcb
gtjaJTysbgO44ERx48LBcz4247AuGc7q8RudqawzOQdLufK+yvVIpjfna37pcM8OipzJ1mtK43z+
EW9PMPXz4tGR2khfI5CCDtZWAdQT4Vg14wPD+UtGQHaMJf8lzxy3LbFwAPbU3hjgAxSH6VWa8rpe
pWL/YOdBSdZfOg9yhDcYPpXNROTxpPLglLxJi0hROaFmeXL+N6EhzFqb1X3dRXm54QQ/le1LZRCO
jVzwiVv7PXR7pBt3nyOHbWd2rNsZhrHDyjRUN/WtEpnCo887YRB0+sZylSCTqoj4kSVf/I5VLUaQ
ytIaPAITEMDIwATojk0l+vMnyxzjAzeQGcKDaBYdeLQi0zBaHFKiaXCZg7li3xCdkLba++vd9iM2
ox/lvX8O6F7mAtRUn7ECPb2daTr40xzJPqqXuYxsrheEkVC2wIvtd2CYshp3As38wBRrZYBGDBmw
+6pI4QLiCLtR6TMagb/+WFLENFSpAnWGDO37Dfo5cmDBrTa8vEdP81TrcB6hUNfAhcgK/fESRgdH
kre2XPXzZvK9EWYCpAJA25JTwuk2+p/VbGUJslnwc5m1rnACHqThJV08m9FxW1e0vV4KHq2Bbihx
Oky80c1JYLx1EKJ1s9d2z6X8AGhq5zJG/O7onaIhVrMlCHRSVQApCjPuarcmtiR07hoPPBkH25fs
TBqwubrdxJdjJjRNctGiHqnDU5LhnfTXruXZAw80dZLrzJYaWJRPRVf7MH3MIhX0JhSKdybAbxjY
whlJgJ/zZdKhhECosjFfXY5wZtbFJLyvGeyLMSkinMozTcUvQrjuFuTWXcY8z++BrE0J58MbXrQ3
fEHa6kk0J2k7YuUkHdgk9qEoBSxNwAvoRGaKsJA6xMql+FggZ+P5bR0G22x+9z6W+dlePNcCWYEI
OdaTusJRmFfx6gxfCYtnK3uch2fPk1WUkExpYZCYzQchi58sHsjjxQwTYeyL1uwHekG1S7NA3bB6
FuTzwxKvOAUjIXy+u5MuwqAaO3oR5SsmkAKH48BpJFb8ClxJ3mCXNj5nSSFIDxApnqMdfmSy3HTj
C7AzNgvwYQYQWZfwgyJzi5dsWHwEypjcFHT7m2aJ8ni0berSRBIg0FN2g+LKoBP7qApPXbPCdKne
fjQrBSu7DUEZFeTV+cjKic4lYBpWa9BU3tkS31niZpe5eTE3M0Ugpp3ZWbpstRb1Qi/+rJKSpryz
67/j54LQyuk4rbp5wrCqWBLHQbhI5USdMThLco5cyPZ5MYWoemwrqc4ryW+wlrbc37+44aymAmGi
lBmybC2PhHjf3OOfLboQZoVKo2ht/Ot4S32VuMPiYwWHC61XLObasWm3xvDr2kDntww/blnunnXk
i1QaZzok48z+QC5zciuM5mMglgPuYVN1HN/ISJoyh0iQGIUnju29aguhsZTgdbBBHS4LysaOhZ55
M4DyiASTa+oZBXWeilTIuaRMr+3gwh1IsKlXZBlVqAGQhCzz5XGF3z9AR+5dlQGCJDcPY7lJBJ32
CnIuBQQdTSx0atFOyALzr5ELNgEgCLv4CAcHiJ9/sAOuqf9h4K8qysbndFj0bV2RYXhcWVLt5tc4
eXFr8/AWmayItoAzrjvxdEsLlDO7Nnbpz9yxQ4OAiuNK87UBern986iXGp11TUIJGh0Q3Un7zogo
9anr83CCaRFo13415v0qnsd2bV1ylviVue1QmXqgWoNSAhflX3YXdxXFwl3TfabWAMkcrEzp0gDk
fVdQZUF8PYfCIJyyF47RglgqxBVMY6rzb6AbqJ+JV76tl4Xpy9VcluCUROWrc5P9FpdqsjUlDycT
OH6y/KJwB/h8nMqhqOk1wfP/P8KWEO94MKLJJIz78uSzrM6eywuZCe7cdkUZaYSCoaoVA2DJuQGb
QorEaIY/6Q7N43d8/tgidko7bED0wYESUNZy+T7w5dRRJZFK0Q5L+x8susmR/7nj7BC8s2SzXdF5
hJIV0iZYV/th1Y9xl++ginuvxE/TChOxSjmWfKgT+mvOPDc4R1NEwI7IcIBYstRoNZGG08poF/Cz
8NS442PEssX/ZxpvJPaVkAresZn8ji64WKybITL2UXbqcbNLEuKs3yTfSNmION4MyRzvcL0xlhRA
FM5xziKgo3QFsN9V7dkF7rBt54a+I6cm4TicyCGFnZpMp+at5dRz7G9C1Grx+8hOseB//c+3qRyw
Vd2kYCftT14WSvbPmpHyWaHG3y4j+mEJcH7ROnme6/H2qfXHraSul75T2lUROVhayIscpi/eBQIk
ewz7+HWjZ/KZpqUbQkHbZX2iWl21kvNMvHVDs6b5ouPVD622rJmNGdZQwBfavfT551+82S8AyH+7
/mf0OwL0s6sGaphCXDraPXj5WYLH3oCSyEsu4PWiLvNeJpiDJW4w+BF7R/2p1ag5RJH7t2n8/Lqf
kDGeg0X+bJKl/wcJxqSOgmt92/jLQpE6cdl9q5hO8jgMMHlYeuEcjyDMFPUU4i5hHSVVpMqBBupI
xK0wlp/2P2yP6bZXgD3LKWM/zK8Of9gGLMk9Dn1fn7S7+jjmBTiYyoPhshZtn4S9YN60RIYz6ia8
A4Ye68wqLdnxpsW0WFXZUdF0kDXEBPvIog1q8HF3xTmE+B0C3CV4okuL9mAqV9zd8ZwjMnVtCORz
URxVccvEsQOOKQI53W/i4QQESDpYXeuEoLiI2ZaKssQ3wwFGIFcBe9Pbq178jCqK1V7c5sVUMdKg
1zKud3t7zDS9GveUgmGXFQEIJZixaEAjUs3QlX5HTtI581l4C11ZPaHgT0XB/Bp4q6V5XH/nWIdq
9CxJ29I+kYn1UcBE+W5RhTbbAZJZRo7dtGAzf4MBavXTUm18a4OqLnn2kk5D5+yQ6vNfXqqcDQbN
J+wJMqwPRfs19J9mX6+UTfBO4PpecNtvUQfNDTRDBJCsvknT37EoOWWBn8/vW43s0AMCAyCWPOm7
LRV0UG//EM53TwjB8tQR8AQoZlWqb9euhOabvMd661ZunZNZ3sYWyuiniBhtOM/KsgF9jKhLz7yP
WoofBDx9Qc/uWWRA/J7agE78rP0GDxq99sgofNMM94krFqy4KrfGTkViwdGzO9p9jJD7ciwh8FkB
TzqSVxZW1g/ZSaSycribZlalmS0TBh829ktw0PGGyL/pTleujl+pkKfMIOjv/Q/Y90fPBGffnnok
M/e5PxUj02/7dKntJg5I4UYrJzvjVxMNOjFX65Lcdtxg9LFJt00uaBeMe3Yt5bowXQwfGtOghCoU
A/nzI6HtmAtQ0GAYcLpE211duL+b789uwZBoChbUYEQM4GmGGHkM32k3vtxagA+P05pfZVPYpwmK
8j+xsjRbXM1VEismI3+VKUhfVgA6vkdtFHmdLCH1yhsEFZHQkGlWQTIaFq2kD772+pnlcFLBNKgR
A5CHEkazcDWBZNYbce/6YrASAtK+1aQyTctYYrE3Jn3596D8AX18nYyMDoVpidne95+kNIQcxwCp
J/70Gz0hKW8BK36fEqA8fIgcUuykoPpi6C44D8Af1zUYAK2Wt4YYRaOetqgblwDRwh/USqRL5Cmh
PKrB7NhezUlYaf2sHmYrFLNfz+5TdS45sQsXetnuj7Th8REewBetYcB1EjiMyzazgDOiMgLoMD4e
xOZv8NsYf9hu5bQTj9EteS7J4NLNe9NWUJnbYH77zPtAtNjax060BPCF1gOrN9hY2QbpSKEIyuhK
3C8kAhRw1hoMr3iFuLqs6UmSgzXEJvO0dbWZVmjOeKYOnZw1MIFDvwlnz65gSWRkWtvUmicYEGru
v4Xl/mBfzOAETa9N1WZNGHUCznjcPsQLrGPyfSLc8pb1zfZ/oogAAKgnzvB7ACEHuM9GwDMEJIWV
RW2h077WReBJJMOa5ldUadnTFbwbkkyFkl96C1O45tF/GdL0QpRuvzGmEu7Tygeo1Fi7LfCiXVv/
nlU+rP11jajsICxtTuZPWo0jrZ7eWdjOMviB3phUI1voprj9hKBUYDGWqKNKNfnMIyqYrC9gCkCl
6IBC2ui5/jlU7hu/XT+3o1ALIMRyBfCTpGLOUkrVRnFIhk9sSS7Jr/l2AkKlQDKhf+Q135jcTJjO
b1rmOm3xAYU813uK9K5JXNDiV+OarFKvb6tAg/aAuA44uxccSuV2moJxBVIHVoFxw6aReQNrVzqT
b9noOXWg/4KNf8sgL9qX5dtFpMM28Gm1TVdBGc9X6sq3HfDV0tHaiw27KwGDZ976tiO5oFcEa416
NujAFXUNkzwAIiD+vX5yQVWjZlyGaBmTjYwM6HIbS6es9/N5ORQZQjxR5GXihOg8gL78KsJF0Fob
mtP+NRCyoi/F5FaqLYMP4P5qtdA4LRbIYoloqs6OnJn48J3D0DK/Vr5FtDd+bkdP6peGlUiQHnX/
I7eoqTVezMLEWPdBDCDvq1O1hWa+CtOBiXORduLSyubth1DqHlbKaWXhZfj5XmyDnJ6Nd3ZX436g
I14X4mcTLKTaSjj5fm01f/TKZFoK4lTwPSOzsNnJWAxY6EIATcl6eovxjjI8abTavNf/qb2WrtjR
CAJULSDXlYv63q3/h5Q70y5rNX+hFpvH3i6f+ZzgY15I7z8jkwOhIJxyVZQc4REofJpdzCOlbri3
rNZtCGw1WjpUcPQdKQgqaBtoAk5s5sUKO822oP+sF2/YESqVSoLKa3SjKz7Kmn3w71S1j2W/ZR3P
r0xAhACE6BCEmSkAOXIzy6JBxCXLCibKtbppJId/dGh8Q+cuUc7olRX8L/Kc/RETjgRBjPAJIenj
onAUu++L3ILbkQRPeE0ye5BmILFAVPBh3qfZrG/eTmWE36+FUCw8IZTopjNEzChxfdR5ObNc/tte
0iX7fsMlXmFCREwmBa4ABpsUTmFcqRegKUlSrm1t80E/lIZcMCmN8O19A5t4tjGXsI2C9UGO/IB3
g5ZYvpzyRY4mrzTW15mCQ63T3pCmyCb5fHjhKFpqn0lcwnL9oq+L7keg0ydEbR7ICvfYY5hGn1Xf
YC3SPWQQi+Tf5qjo6oQvLzeKvyNjItpFCmI+e19KkQi77dgH/6JKq52+JFeFeBW+NDd16DLKb0xV
M+2lr1QYrlty1UwGGcSmhuKHs3oYkWAklt+7/zP1gUlMDxvHKa2I/FccxGkHdoF+NlfPMR7GxHGp
0rjNbiOFMsojcYp9m7Tc6GFLYF2peVHzrW1ZUDTSZaBoc3gin2A9qDvUJ3w17HEgf4TkSiH/VCQt
Sqe7KFaYGk1daV02s6wFto5rnSGL1g/0lTfPXL5t4E3oMGPdUc7Pf3rc4qr+kiTugWpNlFC2H+jA
i9yUuOkEu+g9rVKYmjwXnqeSaWgKHUwIjWLjsChApH5fQr5mxqwb5VhY6gpTD6J1bRpBS8yogkUu
UZeqAk0i+c28YmfIMyRc8MzB7eTeo73TKJ6TFwwuK2OIwIOu3tokiNPNJf72n0zXuOt882IqyIz/
dkYnVqQ35J+/CM21NJMl8PEOR3HUTVs6t+c2rWOiZfGyof6NzTNqYymGTQglkRbMZEvVbWhZfw70
8ZXmuahorvKIYOiRfJzSvOpZ0OzdPewUO7e8m2fFdOpkPHke8q1jMUzE4+poV4/lpx5BsHS7jRNY
G+0MNQvDS282/uhd4PRJAppLmksUfeylM9khSt341QcF9hgyZ+GuKl8dIIsNhYo8Whw7uIu/h52W
GRD7ys+t/NxxZZQ/jeY4Rz7cBZT8wsdEvrWfU78kGnAJQn9GdB0vHPZXGGobyH3H+WEfo4BmxsX/
A3kqkFNC7SrK20ziBxSzpj4QJs3cgykYOkthi2Xivst18UMz+SAP9cqwCajaAwVfupU/ymNz1quK
5SFQtOaSzgMb4kt0Aiq4rrmX0z+8aF/PMfgZUbsxaXfh9wjZNEXcFE0YFBdWIAEV1YJBg0bV7o8X
l9qXfr7ZvowsEDRkbXhh8EZcK9FETI3EnyTnyBYMIJr/F7xXh/L3NK/LK7xZsbODIgNaJOeBWQBn
g3G5x3P8iDy1ojVk+w2QP7MEQNY9/0l7Bv1nELtu84bhouCJBiED0MhI6CWWABkSmuZLvf/7Afya
m+hFqXjbaNwQNGusFzOVPMRtBOS9wnb6EcXXicUIxR4EP2v4c//Rij0Je73suVhrszUSBidBGPsF
xxcEKwNGNK/XxtR9q2brdDH5bj+Ef2iXu5BwY687+uZfbdV58fYlvDu2o/IuBKsbfPEYMlgMk5WF
MP+kkn1yulM4OtRicCPt/M+AYalSublkSeiKmanlnaXEjgRkSqphICftSk/veUp/m9++qrD+2DaO
kKe6euZnov6eowGVroabazVXiq+2sHh53px8bV3yaDfObzXegMOrI7dA0loF2y559Ei5IPuhzGE3
RwqYu4ccKZJtQWLGSDcJoFfwG6m2gO74MVPsGvKqFOcTOXuKjk/XPCtQQDvJOT/fjaP7VeUF37RK
4HLdVS6j0kUof4CRuQOk+WH8QJ9HsRNSx1HmqW5s1dlVb4Say3NQ0u/wpNSCD1Y5zNX70eZsQ4Ok
WkTrFPBuJ4cRHK4wqeZAEE5wM9TKiluww8kbFVn7l6LjUXYyrMNRWyrxf50OY5ejs8upXOKg0Zsc
CZptnnfIdV47ynW8Vf/r2ddZqay7JG+KLVuesY9fdYLOPRpiCe6TKc7GiRAjgvSG3S3iRMSbn1a1
chKXw4dj85zRscOGmTEBXTx1M9siv9niAxC/N7aoGfqdqbrcffYHfnJIJvABAzPcSOqtVGXPaUMN
5P4dw7Dd/aKE3zcyUTIKRWsJh/Acg3YO4oSoX5vur5/ArfUyS+mwfgCZbWTjX17K3DwmhAf+tYvw
YK/PxPIqVZd8+X9lrDRWfjiaGpZXRbpAHS/llpYN/5H1abdS6R9hzo/o36eLtgL2S5lOULFEbOCZ
vD57RhL/a6P4ZrApgGFdVDmwukj+bw/qqBddgInxKPaL+KOUYyQBLdD/otrQqrUeSbHuzXGuIUcK
p4nJcoStAomRPvIlbHwlnb9e0GM6+V7k9jvZd1arQ7vfwqhd13qU/X+DAe+xlUukreTHYltArHBa
289k2a19mp6jVpcTZHP6K4jS+3vyQSGP/A+8NRfSg1KFCjnG8yeclprBwMCrp1PA9N/AIcgcbJ9C
ZsnKBkwvFjOcHJbQM6rzsm6bW+4LH3jj3piecMBrtlQK9+0r4mo0qWrOXUWiciUYe+owEkgJF/u9
m3u4MeDcURTjJ+wS0lt7GtDTOc915IMfZtTqA0aWsfGkG2gGB1RgoRBw2B1g+QcurBk1jAoaLYsn
Y1e5hkCWogjsaKDiCTrUBI9B6p5T5duq+lanUL8z1JJx9Ez3rSGn8rLCufn+ee91jG78hI7gUe5L
68leYwokeBLR8a/l64gA2m3/08j2Tmr+cwxuzlObrRRT8Jf9sJpkOGJCJRgoTajXs08CC/AIbKeO
Uv43YpbsIM9Dh11cgWIse7tUOkxv6wzPeNnJUtCg/Nf8qVbQ6hzfmzBj6MzXhEZQROPD4DZ8J2N+
gB3leX48lz64X5utegT3OdbPtlBGlp1E1wkb0Ae7TI2kVUvTPq7p3xrR+d0XJHuW586TsWe0+FGR
gys23ephx5LkoChcs4uyP7FVawYdlRTBiPLQXA/nUWQWJ9y7huW4AtEGLEbarEScX4burPqzawju
DHo/ECgKXfW2m8Mt8BYPnT9WcIhSBM2dwAH9wpIDbGzO9v/MI0/0l7O4HoX9Qu/O9FkVOF3xH10q
sCEWQtffypcD2zId2JLvVgpPSjXxFGxk8K+XilexVVwT7dA4nIMd2kEESAayIvrCf1VSWaIvzybe
2fjNETGOUIec81OcHmIzio5O+5lm4jTyFgnf3urWuAg5PCh3nIU1Kb+fFCmkp+KpYsERxeM++JBu
9eunFQR17sxQ5m+vrnMSPU1ve41whnmvzX5BWDngFb9ErnysRgPOoMnVeTIvRW/U+VBuuDlE5jHd
tOSWroqrPr+HIijyFzPKaCKaeyGbvoYWV9eOxa35jyyhT2xW1iVsQkAUY5CLJnocVqpCGEedPQ6H
qf+3lhOOoPPTVpyMYXWVjTk0OuWMVhBAdbniTS8nPyzM/zJJ2W49mGgzseThmeJa9VVEgvfs1QZH
910shYJYBXZvhEi7jpIESAhj1NP3cfMTsKac+HC9tpeiyusr6isqISAOL/FTS0Nmevem5Slsc0rh
7ySnMTqCdyH3233EDBbzH1TZ1lBN4EFGLDzZlmcqb0gJdaM+S6QDF2xammwjNwRd3IxqWjUwtjoa
qQYHoqQWGxZO7hy+6QwZnQD6u2px2QlGlCjg7Cp8SclpAo8IopBNeStrZzmFh6KD9pwPCelboj2I
DCxEzYw9rL3hfjJ+6rBYsJul7ONISHVwsBa9P3QWeE40Jw9Rlx4Wccm2dQAg5y4rIj2TNbZwOqCt
LlayFxqLP69kpeGpesCaEkcpgd87M2m9lYjVznzJOANYH8DzybqfBMtYOuoVkUfPnlGPmESB/HIe
mQ27UkIq77f9T1jmS9vuX+Dw5+DAFgpQyBFuXnr9/gP5M/TOyieKsIXdnNnh9Ay/cPJ4DchX46kx
afyfh4Rk35l1xgFrzAvniDwInfyI01+eDDnxvc3V6Ddp6IrVrVAYfQZXg3RnD+c7qWD30aWXrYni
omg6wm6WK8v7PL1iZ/AtZ1lg3olM0xpm/MXfJAIkNKt/9MwQOucdw4nyw/vCdeKBfjkt0oalymkC
4cwYYwx/QSnXHQPq052TJRz8AVrHV/bKhqiLDLtWZ9XS936FPQ7RSFA9EjGada6Us3P21es+Bf0i
FfrwlkN6ihH4D/ghSOyoZUI7e/2gleLheBnjAY708JPavvylXjTjhUFcs7QHcaXaNw5a0PeKDDLL
Gc94sso/krjpOtRCbPz10B5WCqxECqf4WiLlC3R7zV72Gr41Sq0YVdi4kuTgy1uTocGiZlZkxDq5
l4SZKa3ttztJ0LbWG3QpFr5cPwS2LsODCLlJsqmY+2Zb4VwbPkmXSm0O6fWD/BdFGtWrMYifuekG
f8UOm/4JeLs6NtFhQ92QYvnTFPwWw0Hb8C0f/G731cIwk6Agdv0i0pxqtUvse2+Mjk//NFVxskO8
WjL/y3II1PBuz+u3Y/L0b4GzJJG9/OAd6Ipk4UA+UJPjqfciHdWlP88bEnbphmiownJz3aY9irrA
bx1Zc1m90fU+wKrLTKqd6Rla2fwmbvjTBhJvB+2cPQ1UUYcgcLDv0W6tJg72xgiKEJrrs4y1d56V
UbPCOj3MrLxQb0C7N3/7JdoTBvvq/ui5lZNQs6tYNAu11L7lID/0ncP6zxdi+nkyrCFnpmnHTga3
6z/ajYnPw4W1pnnjH9zmIoSybSD4eCcIhkYj5kLUHsCkgeERs6bQePn2/OJpURpxJNWLxcgGnCQ+
k1C7a38j9WWiEYoGBr1tc2qKczx+qzVn9l2lNoPs+/g54pGHL9qQsLPyN5AMnD54RA+Vg8wsdHqR
TpFt14/r8t8AenSi7Y+GgZ/GJIFOMOBK/Y2wMrrDCypIouz2TTwC8/Z9sMsouxslUzZ1DLrMQIV2
myim4pqAfEAQGQ2GLMg+HiX2N2SpwzUZtKzH3wpmxGVlCO7jQQXRI+5heY8JavSZYqJ5WmkE9aa9
5CoovIpFRfUSrFelf32SCN7YHG0lOJTC0LhzKs6W8qdVyaNWxlvqo2jqOObKAjjj9D7FWdHfSVfB
OV6qG+KaFxz0ieqozEaLzmZCRjiQdBzXApDT5rHypXh8jgMrts9BzUnkOgc6PiSshLvsUfwDthF/
JTpjqLxUrN1xm7XuOgoZKzMCbzvu39DLQDdzi6LqqPrQWtA4cmaTsVFNTwxwgUFrkoFx8iLRJPtB
32U9T2kbeVy0OoZWoEesOL1sBXMw2Xsp8AEwpdbbIy8oO3DgjEN3trKIQt+lKF6jSFnsNaDUFSJe
P32Kmjop9TvTGkg8FRTIdFHWPLk5qQyNAXa3TrdCeoF42YRZXChPXuXeDbKwMImva/gicJ546wjR
klybAGkbeRPZMUtXt27COfY0yz1tDs1AWjY+CIUk+6j3AS3A0pXFhwXjRAfC22Oupd044BSm/Mqw
dwaefQWtOsgkq9/gVQDo+1TySdM/wNI+RHsq+YSue3e3b2YiTapNAdq+G2z2X9CcU7HY7booS2v8
deaBKmc/tN8A8V1yuE1THzXZ2QH8HeDVY6VjnxMTdD8wICj8qyN+BldBSf97ImgNWq76xKmWlUNC
l0FQcbUJTppKkzq6CmdgGngtwDQxC3o/5nyj5nFkX12aWR2KybPUIQ8ng6fIIbrWvWRG7+GwnizS
hdsnyjUTfPtrEyc3Gl1f7aPFxGMYdMliRpYvqcccmHTn6kpjy8tx9dAG+540rAIbsNo/NzldAeM0
+9gwwIjewI3KnZVUYG40I9SeW8JTCOGKJahMT+q9KTUE3w9gs/gBuQsZ/pW0X9+4opUD842rnDGY
8oXe325nphPJ4q58CqbDGOMFQQoFNdL62ywZR+Mm5qmqDH2aDakIbSffwvGS58jraDN2Hiee+768
4G9ChyQodHHU3KkiJiQVOd/2NBgsk8pzCaRzN4ZZGy4I8EmSfVebQP4aUuqZf08R7kxL3u/+3boS
UstsCeLKPMA+WMJv+ZoX6kzuA/m29wHcg8TiM8A4WdK2JlI1iG9w+QA/G7KyirWpCHhoYGTF4Vwl
vetak6mqXUuksVpl0Y6dTSMTd0Xz0+XluoV8TXwonQznrxnBbPE5zPPAkdVrt4MH0nTR7QGqaT8Y
JL5wvb8WSqeVs0NZsrkCNnGYQ5dLiHxgqUkF5WIF8yN5YDlaTyaF8RIlUxxVU8xbe3HiWGBvjNAn
3d5fWeK9OxShFIhafZoLayWD6JF5BKio5vCiYCUbZBIIOfaJ8Iy4SCNYrfZLYQXxA3tSczQ8CfXF
ISnclOKFTNnoSmMnCWTbKGGosIbwYIhcSw7lCL45W5zk14u1hr4+7f7VBcTlwSreSJSoWL5Od4Pe
Sh2hRR+HaZfOa4Vx/cyarzjOEykbC/JM42Vdp5LNPYPcNlErfaapV6vCARqSPBCAjsDt4Y/kMBj3
XOknHEoMS+aW8qNRqY1DVY4dbxLZYYiKts+1Y6xnoJcUpF0zKXWu8umIsHlIp2CqSuKBsmBpj0Dp
jquaaYbKHZSHp/dCiUIQGyD9WFNngSZbaZRzJqh25W3TzrN9CQ+blwUYBrXvklkrd3WsR4ZucXUd
HioBOfC3hxL76NmBcZzxIL3o961OX3R7dfve8XENtY9UEoQoGtx0sOcjDTbb2uVqEdH8dGgMk+h6
razuGezdtq91n6vwHoKsabo8HFVJ1kI0xOVRJoVobrgiamjWiAxE4rpHcMfoLWtOS3tW+61zuRPP
c2VMcylZMa9r4zAs0gsP18dInVoIA8qenGAOVKB+Ep7crUOE4tHqdZnSSK4BJsHNc/uFWFFKlWkQ
rMXr1TbZjMpXvl3pYY8xEPpI/CFwKzMGAzivoKVMTHVDSGzHr/QG1CGEefQUUpr9Oz5PPqg3WQ23
kyaDLzCTlD3aM2gXXZX6+R8Q9vXAXt56FpnkrtjPjZxpMlvByIYRzLwFq7CjHhM3l5lRcOZ/dcn/
ouI54fSos8EWk8ohzTi6njCkRd1OPCUGubmK66c1cDS3zt7E0W1Pyp7ID4B+Gfp/kqn4D8crQDUr
VaP0Jjk8D+zAQ/zgfqJLiZLpCPXaDqiM2K73469nFDU1yud7aoBBOcj3iZS2QRup2wEbFmAEuqT8
exqc8jrPlJOyVFRJD27sO3gqukQY5FJ5upJjrPGPxDyvS3d8xqFaO8ij7CilH+kynaKpvkG0ypmO
C3bZaKl+3kji8tvrLMn5TmXY62Zq0SV37mm9zJB8FGaO1wHsgcXaLD0rf9wNdFNdoCy6zE6rL16d
ku+6oGAYed058CdN05allgj0q3VEGoye1OTLCv0gQK+YbJmYfv+DStjgX/+7zU55C1jwzpu6vK/t
IUBMiEz5to03TllZQ2ugkIKwm0apNX7BJYvPclKoPPztwSYpBHmIpubj3xGJVzc2CuvmlVwsaanz
0IOv0yl2SYIQ24B9mWyq28gYRcH5LmIZauRbfufgM/a+90L0Wuv5yG51Gu2Ay8uiNl+d3r+MronD
OBg+8TDdygWTzCmPZJsPs3Cyj49jXfXkaK842EswMLAgWWkXQPvrs3yxdI+Putte50dIfKW0ufmb
bI+T8WyLwgrSHOWkqk+PT7xA50JlQT0OTyTMtD68mtyD5rsP6A1xXUa5vcQKpVdzxXw2U0O28gQ2
wasd6kt+Ad9N8WrYecFSyHl8aYNh3ZQ/4+mn/1vxjelM5erwdE71zujgKTY32bPQcWJRZJAez14s
0bRq+ZoWwhgGKEGCtBHnER3ZoI2ALRQXpbb8kYrt0Lw1lU2HkD8xliBsvBj2Tu2EA4KN2yUf9qn0
npSIM4vUNR7EI7yEVEloN2y8zyKxNy+zi5p2NjYtoZA6h8buTCiksglUOlrK9cDsOOvsZ7swz9Qh
p8XmADlJ33siH4iKxjzVSGE0Rt5wjsu2alF615bYEet1IL2hU+E1MNyMM1D7wzdmw9h2DY2INO0x
oZHtWhRU7A32Mk/0cDRK+y07EXLh4/sUz8QNc3gw3lBsc4+xtORCBHyKYJjzTazR61pZZ28efXO+
tVxjP6KyRnqxt73Ua5lPcdE9Z4+34T5PHqjfa6zkWKIxTNIU0I4RpBzwAV8QEGXeAuYRjceA6S6V
4S7k76AvaXdDo5uWDeo7IR0dcYhEf5R6qgPBWCq6Jkr9EDxef7/W/fbdHTxDkSzIOIMt/uVpZifY
f7QnQB25Ls4ZqcTVnnzbDM4ZwiZ65m/2tExerBXBERz7FmUoM3+OzJVdvxHnQKMO4w/3YuOzoHqJ
QZioOhc3eSapwiJYAOn1SQ/y/g9RcJdvl0nW60rRBcxj2qhBo6J+C5DgYScsCwOIAOFHCH38Umhy
TXlH+fVWQOahCyXZTPTh2r0hib2FyN0amZ31Sv8Lm4wQ9QTp0xkDNSyo+e5XjKV9vshx2FKFNrpA
uKJ97UgqyLyNnp7eHSes5Y8BJRD/99FftuKKC1rBxpVXLdF3t4pa+IBN6ScMP+OiB5MNZk3BZ3py
moihb1dgwK8Iy1HEc0EVmSFjtSUulBXq09RIBDLb67Cn+ywa3x/0OmyfBzMerWxbmSpALvSrMcvs
aijccI/u9B4Bi/65VMexKgp9YSHAP6whGDNKiofNRDddY7KChSYbR8f0cIfQ7msNiM8wMEvgvCHA
NP8bvnN9031r36biuZEKDtd2/+HAP4PySLW3CODWl7kxt90Uls/cXHe6/cVpCd4L5HQZXeh4QglT
jHGzol1HJ9Il7fXZHE7YKGS77fflcOHcNEwV16Pf+y3ir0D41zO5cuxo4tQzV32QFUmPLn1tUUIf
U6+BfMsvidLSFGAjx7WF0E0tfqs1WV8nmdxcZqWPDVXbGRwzjW0wuIRi0Ki5cQ6ejdzWJDNrGp5v
KG9cfjcmhiqx+q6JTnm1/do5QThuW34TeiJhYmdipxKJMCtsDWXjFzxHjLQrdx8YUUGPOpF9U0rq
uRVaqz1slFSdIl/b6y/IGtG37IDCboyi1y0HbfI8rAz7He046HnVWME7be2H6fK2bhYEwYv2qYPW
j9/it4kES5OSY7CxsChZZ0RJ3H3gjrWDan9IoIIUfm+/Berwycc3rx9aEwlZzCpZIqWjdToQwKmI
j7fam/dNfZ1BVKDl7Zu85VTljfFJtDUPmk3XjBDE3pfo4GXF8o+IWSnm7NNVkkdxfqE4hV/Nwe66
2hkQQZH/1Q7e2qVwf1pg035UGckXcVw30SniyRLmBji4yudvpfZlik/jBIcsrnDxqXCvE1jbR72+
LvyDYpeGX+EqU8V4yJE0Gdb7Cs8P7oKRv4XRlOqJW3aVAJ4r5N6L4zw38021jyKXZAp0y/vSa/nY
u/2V2oXAP+My68OIEJ/UdPdZ582z+qMybzqd5CQpKt9ttH+y6C/N72RBKSwJdE45wZbSOXHcVCI8
xsWEcVmOssmuBxqbU9HzQ8CFHDs5X+UpD19OKBTSuuvmmv0G3B4PHHI4F5bvkNvoEx0L4vxXEII8
KRdCx3fB+mThedeSynMW3fmXg9pAOpWsqM8gznBG3otceFZhDrULgwqrpkiyPxdZ/2PsovWUA+Rp
BwvtNEshz3y60lasKd2d5vRqri85ZSuGL+qF9TBBQzjTxAwzfyeW2cPdIMcpLBDYFXfORzTtjgPZ
P84qQny/whIKCaZIN0Tzof/CdY3ORdwkPJity/IQS10U8+DV/N/9Vhn0VMrr0aghzNZUelFi1rKF
IUelHN7ZFU2bkdOFltPJrLkpKIkj7X4zqTxXzlE7UCWQH1VbrIv5vkyYzbXB8AhC52cgxbSgmsgT
yM71Fa3YVusvuUgFUki5CPN5+8BAOsRxjjYX2SeX9CDgmorlPPGKUJIqnBvM5OjtUMdlpENkFAzO
PeiSVfLNT0uNtu21wXBofcyooUpjIK/pU9V+5Kilb/3Pei10inEZNQHH4WruCtqj5lS8C2xp9zds
/84veaJ3x06jsIhlM8ZkKf1lDRY0XSedXlEJmZ7hJVosxrnhAntz5NB+jgGPI3+eeeB3rVGncgV5
6qK2xymbf/9foWebhc5/qQjZtSyU90AdgXeTJZ1JbZqOWGs/rPjJxoFjH05d9YHH5bxvw6CBlGr1
oa47qNVAF0ty3WKl77+LQ14U57HtvucaB2C8IzaQGcfkBBb3O2CZzo7iG20ybYMppZWJGQss43fN
vLYZdn9j7oysE2w0J6TFRiSVXQALrBHfE/kQLcwiXNEgPrad/IujXCt7652ndVcOYUdh5MdieUQh
2zLmz4EIVU1OAvOUqWtl0W8/Pgib+qVluhv8Ly71MwBHJL038LddYI33OVpQ0BlNhi6/0c/BTP7v
8vvqH9IaKXQOqxLgbwyvI8C8MvJ+P1yD737KoH4lGpKwTtJLPOYd76vjyBXS+9qGhMTuS+5vQkeA
kSLwYcx7LMJQ5jW4seoCQ9/0Ta8JqB6xEM/Ht5sbamPm//9tBlvjw0P8JfjYP0AwE2zDm+nZAvD2
ETZcgeCeILMX669749qETBTb0YTcAcK/WqIvLcBwVBJSHI+RZjgQf303YpZD9lwzbGAlfq1JKUVR
IhwieHgbvSQAr8HS3RpRCnZCbYAwTb6LUiufJiM+cHR+IyJpTZMglWmwTHCYxR0RYAW5ar10GBcA
ICGt448HTSv5vG403i9YhcEFDWpHhiplt0cy54W8JIhPRKgvPPTCmtNys6/JsFRFYmpHPU0gfGk5
tNMc8ijrBfbZXRWVMmdkJ6FnpHc1IvUDkB3cCcFYCNHDg9kSjeKVP7Q17O0wdo0m5qswStYd6sBd
CsCQ+Sg7S6g/KjjZticd44kNY6nKkQ/XHKmb5dOn1bhDMV/oQKjq1Utk7+dmngkn7NyvH9to97jB
E2GYbmmgsJ8aPIH9htDdh/i/8wQztPazQlICPdPEopLG7KxbvN+gKJjHiBp13HO+36tH/wnID1Pj
PyF58UNE4EZDfB7HnNBfkOT3TQlhCNlBLscbCavJx9nlXSJP5EHaHS15pPezPCAlmG1VwcaDxdAi
UGfKV8fzakmy9zaNT7aTOZxiOuiz4WfT0WsbNDS3/F3FXCNl0YBXY/SNUyeANTSqHtd9Kkil3WiU
NHh9p9fMTBDylKvGetqlDEtux9GROD/cLWgQ1x9L6VCJ0Wd2Ojhe+FraM+g6hHrSr0npE8DZ5fLH
LVoJbKM8fStzOoMSmjGyMiaRCkt5eOH6Nm9N6IBPCZ0LjTTn1FHj+pYDrLEeQbua/z6ks4o+gnHD
soDIpSIkv5sljAdMhqPjNEt5anYlC2daBBl67CuSCSnRN1e6Zsr/c3fQnSxgkgAka0GSTuC/Y8Cz
NbWAfs0QDBf+acIBgrFkbnJObn+eqExy1ZJmxLLbUwIwRKPHR69RpLcoQw8z4nS11GsbbiPcnKXp
crQYIdaXcmYF3HQknSrT9rnML+AO5OuelFLJvccsR6tnywU3hymu7JqzZpp7H7WQFa4E1zzwqoM2
2W0HZEVBynnT7Dhtjhk13MCQJclf4CH0A0ohTHXy0qja9TijWVyZfoEpbyVFH3o2DqgGA1f8GLv6
KBBImF6/KAzrkq5pU6UsuQSQ4j2IQdT7S9Mv6eeAP5dQ6ZVdcZEv2GIqjYyxLVA1tAtSH0yc5FBh
ASBy5h5H3mMWsjasPtRV5C15oREwF6tAgPZvQ2OIywE/UOkbKrp6agEAeOmC7IGwAd8hshs7pPpc
GajP6Gx4/ZLHS8fOh+ZVFLPFpjkqZ+kIyIgTujGgMAgroCEkweyF7qnZ3FPIiGM/6QTSLPFB4aQV
OHXlcJh83PLjPb4DYXibBWwdmvy3cvH0IMPqPDRGcDOYXgkTgrdpvWzZ+f9CeAkj5yE+6tIFJ9L5
ZjVfQTsKJjlSihvtdZbN5oVtoL0RuFHLEyhGKrMUlBaGaddvckY1CTyMvl2uCzczmUQysnyawyWt
P4SVaMaNttC9BJLOfs0HYohh8HHICxqQIXCLOFYlajBisW79qlbbstr93Rr03uUGfAIyW9exLdMH
GXuHfL+dq4IAKs2Qhn/DjOtkIXX4IPpOPQxrGVFVdOecld94+c1wOIRuRcs1Wm3+UY4uYDOWRLms
sa+YycYLjSKVfcXpDXB13LZllVDOPkfdAVTeChNwU1/Zry5lYxOfnYtug9vo7ZCPacqELshmddxX
VpUDbpTkzXM+5ngws74XK0jTAkIWPAUgNJDaKD3DV3rqCZAy6rFTho8Ny7uaFyseYL2LY1IwtxD7
Ob6s96RM6KWCoK27D0m802u08Rp0ZfnwGzhIq7vE3eR29aTTJlLG6EN54ZTWxB4kjIWOK4dQPdwj
JZxiy8jzr+1NX7EPOZIWVxO5e4kIjdrZ/goYAL7dyV3gft+EIkkPiobhGLim5bUSNV/4qFJGqk14
QmLkl/avQkaAzVl67L+a5RqyFLHEMEm9cH6cFCxJl9Er1fqsWeUAwvxqoi4Xu5OpKMS0Cxhm9fhG
iIoz9S3Uid8Q5G1+zX1jMQgZkw94Ad1kT2V0Pk93rlq3Le9VSjeWn3cxIh9Zsf+VavEK9Oflk0tZ
oNvzqAjSs3tylQRIP/9HYHO8e+Gd2/8ZT90eXaPRcKr4gqfPDo1hlNVNx+hVHX2uj5DwcjjY8EYY
Lh1Zm2uf7ilLgf5PcOXiCsr8UDzWT/DU/SXcQaprGJENxjO9ZZq8zq75HJnsVyWu63Sas2FrviVT
4Yg8OB+H1G7vmidFyWeqMFfULscNZlnIGTaDyBWqVo3PJJ1Si35GqyXklQ8ptDJEihtYAnJ45LPq
NVZKdi3GpwqK1kcoRZbUv6ufXhR3j0/RbvWBsbSJtSBH/gltwY0QiU/inQwCelYGdiY7SEak3gSO
PyZ2slBiZs7/MjGaRjA6B7HsYcJt2YcUVFcWrlqk60Wl/3baVHHsOpqcJtv4XPyTV2QLAM2egiuF
rPru+AcNIRINdzFXSttOhDOnqJZURZFn4poyF4Hn91edXD723XObnM77ZMKHOTBirj0y5UQM5V4M
5GoHfPv1F8QK1wqnTUPDAh3xPzba+N12v2bmoTGBqAqvk6ZNfhD6gckuQ56/qQgiziHB63D+6YZE
2AJ+QGPOoEnVqt1rx0EMKNkZmfhABAkB5WO88FWRe060wysLEXxQAF8iQv8HeQAGD8UDiybEEVlk
tWnRQL2G1pvbNDrYcJd/78ye3MRhBAMAx0emSRDtEmsQSgFNaankQ1zJTmjRtQ73NN7oAmSe8vwu
0LfGcz38B3WXtEkN99zrwmPMGtDVGN5y/M5vVZlTbraFZOMYmvrsibt3aHTO1HGtU3cXKIJ+vOrQ
T+xKmh8Qd5+LwiHeDBxNieSchV1IQPZsDFWCd3ryswYY0p839ORHkowaM98HgkNtpCy5yNBFuAsE
Ipc1KZoyTlZZZQLFL4vIGrObC6aAil6nBduRHYF9uo2wLEMqZ1BrYuCd3OwD1gE4XJhPcHU1nPc0
kBIpF1mHlmDbeqYDAZPQH4aIK9T9ZpelAGkyd+325ShA9xDHjt+33YmviGbsnd7xT+MoazuAtXTk
ItGY1eGXp0mbj+E/hvA0zu1evEYEATkIszwh4ZEpuIBhAUIXPP4tfrB0qaDUVklwFvuiB0dV1Amr
51pO9QgWxNa00gDrndeB0c2QNrdnjbraZIz7xtIC44UqHFcotvzqg778UTIcZlWT7ofZPdLKVy8e
ZXKD8+EP4VoCD87xFOt9tPO2GLyP2MYEbYT1e9ax/UyUGuYo/fIpeUd5FGaGWofiog8mVzjQNtSj
mIrdSX4TLT23BjqcAC/BTP23m41kfH/bbybq1x/Tzssqw49JPDOR0QCfH7dNqyyIQxWqvksCTF2m
tp7NokJpdqTuIME1LJ74QC0eh+fcUCNXN0yfZACt4gcKKcAwnxQ+gQ76EUnd2PMq4YSn7BWLMhsZ
+YDVo24dZ+j3NIXoMbkrh5NWobTe2+rQEnh82VpZPL8Is0NlY1vW9eO7UiHVMQnRn837l0zU2wgM
76oF5VvefUcGZp2Z9I5H1E/elWuy0WjMbralum9VZpu1Hj8R+iY9rNSBQijCYDMN/hqXSist1GKV
VIq60kku1/wfeWEyCmj179CYuD2qKhl9Au0Ma5+y/VoXOuUo+gAfrjbU615ygXpMJNT+MtOi55od
yfbAwG0gDIEPPEUvVlyfm2YzsLHRtU90X5HjiyBhr0iaN73UtC9AjuwFdJRsGgbeeorHqvWH7HX3
gtm0JPaDLCIzkmGqqHekZzhm74ggeclPAeFqtZpQQ23dPTFU3R851O5aW/EqXaj3mp6WLmcDQ3Ch
Z4svcNqcIf5M6GOqQFHWMnAKoKXhw4GEbCjX1Hax0m3IVjKVK25oosuew3RS5vhLHm42Fu7/FYFx
OPyCrQOooIavuos2DdAJf31wDSKEarkunqcd3IsAb6UwW2lXVqOF8tWVCd06MAFrRjTM/oe91GVL
8UGDaW9d4IAZL4IvDj6oq5/44GzJveslFEs29iarw/uhgY5YkMW2FVqnaddKRpoMZMXkauIBJK4j
NRY9nliT4zYHcestRMI3G3/o8nhjwDSlW9P0SFw+3e3+Cd/84rsOPYYxR6WU1dU9mw6QSmGiDrXh
y+exxRgj1NGR3PrO9kX+B8wdgHbHaDb2MW8aq886nlHC9fR2Iwq5fg1aPftA4GLQvfuVE60i2fEl
sJLQHLa5SAijubc3X1qjALMNaq3uirSvbb08Cl58nsqz3E9zmY80fDiJ/g/sJqdzFNqBfSDdoUu2
m9TEMBv3+MLPSTBMdN0i6E/q7uopvC7VE004oZ3QKqb9+8kLkRibLOTn3YN2MDqTZp4HniOTVqI+
nLSJW6AV1NoM4/lhr0uY506fbf3HbWiANX5nyBNfwoCg8avuclApYwlNU2xLwMcrIti8cOJwNEAl
wlAyDD0Jze8JN7r5G76NwisX79qnCIk/nHDoIA+tF5nWBGiuUwQQBBsPcWBcSOlQBgUs3eqsqzO2
zJbRZ5MkG1uQjjXf56/VAsf7fqOJiSf6fhp5Wa4aVHfkuVd9wF0p0WZmWtUcImrMil/OfAbHsapa
fGWpBnY/bhw/nZP0K1w2hCsWxniTXcTkywkJXMDou7cRBxjm7939Vm5PlMK8Zzo3f7mRWkBcC1JG
m2OxlNtkenwJD3A+fPJh/5nuZCmvI3gAro+67x+r6KXRHH5KTHhnlvDF+W9pj7N+IebJZOTWdGWs
90+WfYZygvUuUk+cPJgqZUxfm7JoCSD24Q/Cvd6URT0OrdNPkUGxF19MZWpuoGMSZekTRQI4ShdI
FC4xmXj2JLbVbrtRxv7hYkr1i7HVUHulOhG6gX6+AIGNEUr6xomDKnoHqdjgcH/VA1WDbnLsWYFM
BX/xjaxotPHfzrOgqbcI65/RLkw+OvWuG7PtYJlzksaS6fkp1bbQLE17GC2U3MInRyWi/ObA3v0s
/77IASCfaGomLmMZQSnVlalttH7gAGIBDtxvlTRge47W3lCRiXMCvMSFhCqgLVRUlhbiNl3A4W9K
IukN7q1eWHS34rZqTLWaLP9m8Dd5sNQH4yeBZElPHHMMfnbJ0CTq7XKNIGEObkq8e6LgnlDdg4kN
7cjDwfZAxY0+H+MrhxcYc7dSHB9hlX9UNGbFlwjp3dEbRJw0QGYobIedl3MVaN8N5mv4SDe9+AuL
Xv/m6ziF2HhBaTLCMrI1XaKom042QqkU4wx8w7s3XCXCGcLTsdofgVkJgcYy0RffX6ZvTSFGisb1
TqYUQbLGfWvk/JqwBJxiTO33UgYG4t+O17VA8gS0BCPT6NLnyn9sIdws4VIk95SgC4xnlkL6udwo
BYItJD3JLxOtdeqFz+SUDPtEhfTK3QdKwvh8+9WHXMfW9CLJDnHu2MdpoglpdH6NlT2ndW7yboYC
5jhMRoOxa7L64I4zTaYoZWTc7nvEVbfrMacO+Ej/Dyx2l8OqkF7vH94MAgIakLdm2RrDFiF4nFy4
6e1+rkTawHrZeVmzL3PVXa/tsb7NSlZ7lLfAuAxTuyJMAwUYKAUFIojXEG3t4kxkE7YBP7epAs6I
NPj7YOVDYFiQaU6JOHCPNq+gm4DJuZlHishMsXc2aVLeAdPCUTTWFb7Knrz3EF/Of6mtUmGt7y3Q
BWb1WDlDzapUfG10hhC7RpvZHIQc34NeOIUjPpqNW48ZwAoy+jeRw5x7ZpDUhosl4xKsR4FByXOD
cykDp9UPKNTYTSY3zs10ht9+exRRhgJ0/lIrf/8rETLesXCW+ohWGaVGpSA44nFcGJdadSi3wRZc
UZDy3mbRlZrqLUeJkpoBbBaxBWOZroIzG0UOe3Av7xuPIMTcLd/2vE4smW5H3wpIdbWsQmWRKzsD
GHanJ2U7jUMoipEL1vduDyzrwP/6oozMmF9frWPko6dQUSt1Ig7jgSP9LnDNoRhlh+X4TQHwpe78
iTvOEULruQhczrrHXsPBI4juuqlKNV7uxxUFXlIu0qPTFEwO04ZvRo2QDl7vrTScJwcCM6Sa0Yf5
Qdn6IUg62lA4lbh7AQv5EeNsr1qpLGpfrfT/oJ0YzsEPgA7JeawfqanaGBL3eBBBTgIVjGQJVjGp
BFfzAZiytAK857Lxnm3VXrNwGi9VgchvHBQV3ef00t1dohApbpU5JE/32i2RpFdwHi9qJqy2YMD5
lgl7cRy5YQAAizMvJ0QRSzomllOusD3dVJ+KQ428mr/9zadPgIyFzqPCcuiuLg8P221f/1jwSSnf
zdZ4n+eubfnC0I4iQx5L65HsKYjnQzJw9a0qRgyef01n4iNH0VKano7R3J/ls+blLoxugsSfjLYO
ynxm0FvPUf4AVAzZSvRmrhOOPUkMC/OVMYSXnAYUE/XlKEvE5vGyukAGDz6juL3ZZuyqlKRhtlYf
Q0hhZiY9DdDQADj7QU2lQs6jDXhcbLxHzPUP5USTaQHBQO6xSn/DcGjpt/O8HJOzb3NDtFMyzjCl
lJy0Rc9AEcgXoOONQ7gV6JJuZAdMScin/CNrouezY3N/ngPRhYKwOn0H3k0HrHi/uwXyiP9uQPzO
ZoM2y6bA5pCIrANSlkYXZ83A5ZLY+y27U08+2ra7D2QUjYKseICW32iJzquLKepUviwP9/8yUPSI
VnZD06kifU70Mg6Pvc3K/BkaDwv73TJEUAOgOILMMjCh/bUEx8qnbOitxpf8top+1j0DV+8MalKj
1bfQxknbsWXwvRFBzz1q/jBpZgjiORU3Zz3Tp1rFOG9JehLWAZL9gF642WfKhSynellWgmISQENY
i3ltgdxTxfdqX8OJeVDRJr4EeLRSE7ELymLZMMeYgjwi65cYI9EyDKg3PbIyCUvf5FKNvUJ3Ulhp
yD8S+/lSaAMPZzMs5U7retEE2SkSB390V5rnycrIINHCANIKvoxvFNoyTY34Q5jWSqbq6vPKACBW
68VlD9TR9itJdopy42HVxbLU2AHryzJReFgIAKdC8NbpzN6J0iIA6INqRXg+K4qVWNuikkGJwX2F
wXk4cOcFdwA+xejHbQnzX1bj4UKZBoQ8tIBKdUZYLV/P6vIWN2Wl1FUUbux21+1Cv0rVHnyX3irT
6beC8ceQwXGmsQDk9gaWMfPRWmfOAIF0O/190R2QThqxAy4GaHoyy4mgMt1D0aUUnqv8+YsEonD+
tIyvnF6rrNObQI/s+NsI5nHJKyqJx3nyQWoieDn9gdGNThfOp238ZGJF9LlUiYS84/GAc2Bu+LJO
W3br+t5eUYFxTu17fX4qxGju1w1NvQGcIWN5UBqo1ApoTPj7xMAqC/EOJVEdDGXqil1rQFIYiT0/
cTLTooTMYE1fZjcZ+3ux7VNI760/eeDtz/OuK3CpVAP8iZQQCkOukw08oOgHzJLNmJqkf6osPZ8v
CPTb1cSBOCYg6qTwsL711w0FdJIULGvoBc6UaGdPxarudxUlMOa24DF3kAjiAkiPWWD5dxZ9dbfq
MvDf+AruLvzrECPK0Z4tel5sv+Ax6v/UdwiaNmQprhYHAtbWXLLi3oaiMTTP9Pl+BgrftyxhMGVr
iBXCmr87p39jpX82F1TeJUli8PxkxDuSLF+D2i4km152bmWBEJR1pCgL8F0YWoroAwy07o16G/V9
wH+t2uLXXRlkb1Mwk+NLNYM/s5MLnVxLQYB38puS/rv6Rmx1HJVRyCiXQTgD7FF5JjTwbOtcz5yE
YebpLcIt4fwkhgZts0BHb3BfK9TXMkMPT/H0axnNbLYncCUlbnraRMAdX/ZlAUS+kQJgLUB1qdlc
DrtmJmYpdm+51L3yqbPWYD5xjjtj+A6fNSw6ujuYjB7QAuBAjuColAn0FwxdzqMzdTFdkh0AorxL
mHue7ARrXFYgj6EtREnySREYV1SgOtjFZ6pcnJfEyX6BH7JUZghTJtvrnpoNjECQHn4vuu3sxux0
VRVA7iS9DOUH30QvLzes5ofzVxbkZEVJWDXPBZRKeK+bbGhk5a/yKjwUa9cs2WgQ1DLV71nqg5jO
jAkDHFDK+j+ifEQpEh7F5I5bqE35UpPpVd1das+oSzYg0HGyZAVrT+7/VfXZLIcP+ouxFC/v0Dr2
0bOQsXMku8wQknYuuSBzXSDe7OGJbUsWUdS1DhZVjrcj1br3rAfvkmc1z1JNm1K5auyNFTYkBFKT
xIw+3jOgv/fpkwHD2SluC1FCvLjhewvy7b+3rr8fk1a25aY8jkz0slqbffK1mqsyBbl8gWwjo7Ex
Z+AGUM0lD3AYgAY/lu36d4okzynlMC7BH8yAgnXJwDNtkDem3fli9ZppxI+bQQhd39w2E0TsHxzJ
VduwYOUVaq51nCmMVEf7LqmSj7cSPDeEIHAfZn8OXRv1TqrY5mq8f/edK2BWm9E6sXiRl3HN75Hr
pbBD21xrJSDDOTL4vY4KmhuWX2VhS1AghboJr0Lt6HeALjlFTmkE9Qyp6qVacNGpDP4yhBk1uYKZ
XIzJArzcNHx9g1IJXasvy0f0D0TJhHF+acFuEPBs9HJf2XNoDEF480Uz7e40Oq+JURA+zRu5fmba
jlWmhAhPvPepQhjp5kKNq7Xj6VEaM/zqDNZntVi+Tb1A6BMpwmMWY7Z0juKrPM81zuWEQyvpyunw
45Pjre4t7/ZCKpKLfWpj9YHeWWYWG7wnp4NDWQdhCgGjfOy06Vk7Nnn1SAexm+CcptNUkQbCmlFX
CzzyOYImwAPSdH+Mh6Vwb2Wpjjxzzjy0sd26Fuw7ymrMskiyT08zzM9TYN5dKl2Ogwax2twDz8mZ
92yp3G/OkzLaGS1kptwbnhqLFAOKhiJ7wYC+zKIR7L8AOFaZ4IFBHDDoBIUEoTfF2Ik/K8su8WY8
yVsbw4YtMm1InS/tHGvWBMznTbbeXWAgX1lQ71YH9hps9VI3ihEEOhK4tGKwaAV7EL4mBtkfTaio
8HizYqrLvdw/YQuDNTOYuZKiWRWp9yBW5oU17ReuT5FolrvyHgP/JfNQHG3DMNBCKDry6QCc03YN
ypEv7Rf7xWGDmdLykYlC5Jzh4ZEeVmFud46HclCeFFFeNSZIu7LyYmGS3bENQ9AsEXXLeLCA3Rqp
zzhjSwqyAN4rqmvee8rJ6qrzKbaK20sNZwWRd6+7J/ggKO8rCH1/scrDSrtfQLjkuIgU2Hd2aON6
DtLOUzsfmHaM4cAvaSkqnzrY1/VzOZshD9aONwhRUkyBeJC9Gtlv+rJZ8zL0ycSHbX7sEwdNmCEW
qEjxmJEurF+OC2z08sYsEpXq7C8fquDtu3AXqt2JiEO5uAE1NmIprJZRtt4gZnZIH+6v5CfVnGY8
jECj7wgLDqaHA5myT2C2II7naPNtM6j1NBN+5LXaMRFyipw6fudsnCHrMxpYhL8Cv5ZUy0jopqfe
4lMZgkAyDWlAF5bhhQ9F5kXR+6XvM9GEbMtpCdpPRB5q7+ZF/vVU2xpX2lpSGeRNy7+h8oX6aAuR
deacrJxegsHHF0cH89HaknUkDzIwx65Ixcs4WsGI6s7VwPwq7NgEeiZzd0HlbhtYN3rH4cXnR+7o
KQJ/l6GSxmgQP9diOw7LpuPuodUweBG5H8iYDsVZwoWBmVRV1cBfk/1xg4XcAmlF0MC3dDJKliSj
CKOfWnpXnTMGI7uzCVtT4fto8Fl3UhiTiIkj6TwQWTBT35kTMShcIZv2N7H4cIjnVPPFiO1e0Ek1
PCcn9NhSm5GwnRyDC0TfemGENm5lagrByGXNwooZ7+kkg2AjaeOJVx9nK6pDPBHI6U3MCS4I1mjI
j88bJ5VKoc1+V+XAzh3XpmSuMISRQ4qC6a1bcLJofcvf32NAXZ07KRwURyEQcHNVl4+L3LzEGNzT
dMV+2IgxYwGHhRIrnbcbWdvlHVKQvyVgVpwmPiShb7S3p8CN5RUeEX6iYs7EXD8IK2FfZdGVmlzX
RozUm9JNBaaabpRD9hfyCWdFbw/wCKw8nCeStPwdrJvsoMawsdIII/nHvMbpG3pfKtm9LqMztgru
4mM6ePwyq2HutNFlW7ywFIyzxeS16QzLpSn7HN58jpNkfE7dDl02xWEwezT9c1ZXPWbicmVRzrua
IpyIqy0v4EpYn5YcHGaud1NhrvGVx9L36VTkTQOgVtCTSvsJvk6oobruOdUy6hvynStja2o/1lMB
c4Jyu6vxbSqa8sRje5G9u+oL3p6F+KT60P+dtn9qEsiqyoCqn/GB0+bjnJX1kY7gxDKBsBuS1gbi
72TY/rkoMvwSu1jI/SPjnoiRsqTqoiD8I7Q4620NLWdKOd8K1cFzn0/bsuN4/2lloBQm3HbtU/wT
i3ehSVSdfzs61m5mruTUwOwdJE/0XfItGzGA778/SIgyWLjd+ADDnfECwDPfnlfFV0GdIjNi4E+f
SN0gY2+CtsD057dGRp06p3M8Js2GbazXCMmQKoil29JH9DPc4pQqzl3fdEJnRbuRd7qx3fiYPryu
8ZZ9Pa+KBV9B6cUvh8QWMq/+ZdEATVjtTlin+imelUSv9CRzj02QzM5ers4ULUuAt0RqorvtJBzM
UecXZzguYC124iPftI+v6zDC38SIdlQtlAI0VcQbH6PdkoG9BHXaSoiXMT+MfyDzWq1WuH8HdJo7
Kr9xWIPS4XKRphMuQOU30HLNKyQAsDcRp5yxQVXPUFqJyTo+YwHerdlyMuxvNUGbJDl9yhsF/PRg
paTN1FNZrlDLHd8+2k5Jqh17tsByBcQywbcq6ArLwlbdAqBFhIMTlOKCQCBBESvHXhyawwkqnNxy
QqNu66fTKPTpByrZvWdX2t484NhCuMujUMsdaKAwz9CgUCnN2rqBfHk3Wk4OcgsOyMNO5+xRcvAI
zDccGUGTfSPFERnDiRKOCIwzU53BKrVnjdcg3z2RUb18/p5GvU6s+y2EsNQxNjeZXxXsVpp2fZUi
9qkUMbXIIPYx0391B6LJwyG9MNnd6pY4OEP/laImxwH2OWVvYIE1e6qeleS5FmCYY8SNjtPOUq1H
cdVHC0f3IZUYhhW3R3gj1zQWqVNaogof1sdRf7vyIA3MSi6hoaiPZ8af/F4oTqnXfM1GUMt+HMHm
hNbTZOfuj4pCuB4ud3p7+hGpU8CYUY9hCVnIvzSukg6bUu+HNrvty2XWTLF+Tg2urwgM74fq4O7N
+G7f0Oy0hwFIfilhySY56MMne6pQGz/NAOgLzOz4a+szPnwgZt0sFaRRkTc6Nt+vRX+3VqYiOrtd
EbuemRB7jv/ZgQjNTUhQ4KGAMD8yAzdUouyadc/HuwxGwksFnKVxq3EBa/2GVNtM29u1FPYWqo5x
/fvsBuq9EAGESANNmx0CbQfAi/RfE0uQ2iFkyrwohugsJWL1QC2dLvcNiA1NunhkW6BylbYDciHs
cY5DAPYYw4NwWjP3fNB59skZ14ycNWv7mbEcqlv4kyAP3rpwKsw+S9xV4oSMM5BFIj7ebZBLoqrt
vWkmv40x6sjORwZxSLpKq8qU4X3xoYkXc5k+o5G3ZCp2eWZjEYAPqpp7P9t31Z4L0ALsFIdzblGv
8MrifEmhCEM/SgO+dCmQ8eGLfntyHkIC+kTDYf+YDfEUc9Otu+zIbrzzgAnl49QSf/CKCvG1+qNp
BB/TWv5LYr1rMf1TxprnBRrovRWr4L2RevYiENnhVTFjt6Pr1reWGGToS0pQlHbBZvECWBpa4Cn+
6m1tK/c3EtZtOaxGX0ADaF3W+/8/BU3vZ6UBNLwDma3aKw+4rvqswiswHpC6BSkp+LruqrCNGlkd
FTx6ox6gGCSDqkmX+EwE3V5cqehyI2USdJU6kS/LaGLm2PSj9lAAz9+Deu7bLOkPn5UPBEtO2v5R
idAJF4kzXtdOFNszulPzN3GqxoDsaBKKmDjMnfuCPyFT9wQnh6PtDLPm6C+IQuBRbwVAVz18XqeE
TGckdaO1z0oW3MYus8TkXwi84QcRwhgRMC+115GUQRWnis8xH8cpTi79gcSe9vlzcU4o8lH53gvo
qi+c3MpX8+a/1PalhKDjM0I72wGj1eIFO6riBbqvU8T6PvUYrNJzalB+I3z54vaVLBlF75Buv+EC
85CTqXEV9B9szp0MmKDcNuSBWe1lTGbo5w+9Y80HDepy84rpJ5kzFWuX6hef3jmPQbY6jeXRwaD3
GZfmv8rx0vrfeFdUZCak3QS2gDBS+AL1ORrxzQqXNH9Xxdr1bOgH9hEhQDj/jmplh/Ck3GqM3njT
GvOI6wk823QqyT2vinUYCdFv596vs3Z07Rl6m2gxdtPoB1N6teif4hIwUHa4dqFYaCv1zfRQP5bg
9DmC2s+bHB87eXxxgOdwq6Rmz8FLpZvAZNIuSGlLo+mRSXirWtBsIaBOwK740YiyZDHCFoYeSzbX
xvhiw79bep2H3LBwxwgOgOlH82XFu2nDPB6xxed5YYzuNOxEwc1asvtxOdCOlXS34ty86y6RNILY
GA5AE9UkSxpPVtana+BR43DYlbfDe1V8yxZcj4jFy5qHDBj9iCRfm84QLACW13H6F9/bcmc8C5YH
bkCZ62VCvAuV6z4qeQUFb/XHkgvDVen66AnfgpTkewnSvS0ifnf+3LAPD5jj66B/CxrAH9QBAQHC
2tpI63fB403FegUHZEv7JYFXYkQsWtz5ySv0hTdFVCVVfuzZ7j5Yvr1CVfqYSMd1G5hAXlbquPo3
xQ3Ucrgz/CXE9UT+cnuzP36JwVi+SHVaCCdYcXdzzE5rFdSnkuqd4Tvwgym68NbcTflmSMsT6EnR
OjmtDTzqBeocQ+LHyR1/aM6ZbSBjFqdSVGr2vhaDAwzYP+tTSApOA0Sif5eszm4cqxwKzD7EwdAz
TCcfRSGGs54W7FDPyFzx3bQk8MB7cpURe70FG4rkno1DiPuZbZZudDId6pwJgkLczTw1b+HbtC0q
JaL6AryEc9KjKypl+d5LmEdMmzBNqeI6RhwDr+9yKUVKnHn4ZpCtBKgCMFr+LAZFYIpJ/UXQD75V
yONkVMxU9ZdmEQNWl8d1wTQBwEuUbNOf7ZqXoQinThqwavKzmGr2JegtLcTHsByuxjQPiIagOTCp
t619QPj1sEhYn/SlgNaluawZ4K1c49kUsSkM+l1iDeVOEKxIy92Uga0UfN2u25CpaYPucfAe9m0S
CLakDqDOqfAgt7g7F8pK2WmCu47WS0XHa58upKoyYH/V/fQ6F12e3sWb9g2cLxWe/iufvcstr7Ql
uZM46VM4XAe/cgai8CttcwASQETdpJHoe+535nWoP63WaxsI9zjg9+W/ssC/FetEu7Yv77HqnJ3Q
Zwmen9qHEipIRUhdcU9kPtOFs4VoSPTaaqv7eUWKQSz5Sl7L+Nz10PC/Yas7xYg+zHXMUQhFaEL2
9pEsmYfB/Gup04EUnlBbsiGluzhlSoMniIyRduys0beq9RTD15ZHApInsN5EevUXco39IC7NElCn
CLLOY7S+zKS+wOXYPmvwnSsaJz8ALaphAt+SVbP+VU5ZgX3k5+ZsvSrEVfLdZYbeS96aVQAXQZvC
1ku+hhzw1W8Jxb11tT0Zuq44YgrygYyiFyEkCefVnwo/of2+M5wN1wfleGsi1/eLKjbpcB9hHrCw
r9Mie9jj0jrdqTM93svpbCmJwNMlJQ0dBntvXtJqCBUK5h/vdzOmse4hrJmoz+HXU8wErgo8i69L
yDGm8xEBYU6Fo5wZ6D1BMHUWISroBTQ/ED981MylZvOyS5uuSTZpipjH/DOf8H4Kg5qYQFSIKbJh
fep4h3uvzXtHUTBI5YcGFtEP9vMghVqyew8LiCpwKwy264KMch1wgtRiLgHH872m+sM7C9iJfypA
8gMiipoz+jW1vUDAYm5xEgEO3wTqw2vZ3EznzzalGYwNkAdtl5SY1gLrtHNJRIJG7N/fi5kyLZOs
v5QFXDDCwwzYxzsP3cBZKyiKQ+7HJY1MqDoHqwJV460AVSMtP1yc83diRF3ct5sHm8oAgeJ3hP+d
lNBVZRuw6C7h1mTXYLVEwRVM8JSdI1l9lI+ZUM06+qcwLvXc9gKrd/CcFPsSQyrE4vUaBst6DAje
4y7Hnf384Dlvn8yh+P9GYI8TPvA4V0hWcdmPdyN+VetI/Q/tjsmAypzNd7coZsgDXAezbBUswGUj
HrDbyeIeW3UR7241NRyPFrzkDZXPVM/uGyDmUO4rd4KIdtqbKL1mynC4HPMVE0tY5Rgp5cCfsJlp
vRoWngm8+ba4FA8qTBIh1/KFALJcai+nmospEsD1cdat93JwYN89nixZKB/FFz80zx9ugQmgIVyv
k/w5pfPIuRnWqeTPuDLKjH2Awzq5oSYmAa8eJTqQnsQZ3jyjg2Du/twIVWGenzOJp+x60250TfeB
su2SIn1qMMVXmSvdbBaUtSCm7Pj6J6HzKVFQrf0/GK752L5j0ZZQkqjcXs0nx3v9z7ELqDNLgkzM
8UEggVCCFOTvTjRy4X33ZLSX/ZR3DxCLnx6D4QImFYgUCFpD+weLpUIx87jDF4gpxyrQfH+Pa6Co
1tuY4kJajjrfprCams/shHM//wQ1zjuUso5VNwNqH1rIhT7IqR+28otgTEwq0/WEhr+USb2WejaP
6qfBPk6a7o2/EzYxwQQuEndw+1jRfqE/dBqU8uuHHcyBhOJcLbjBD02AwjoDyF6Ei7+d+4/YB1t6
hUamFE/iF4TzNtWerTjxEDwE76RMaorPV/6qFEuCF6aaSC28eO4BHyHwuM/gOZshT4gQiDOPka6/
Jlrc0M5va/4ovJDpKuii3sQLwkLTkZhGIm4z7FLbHITYqavqYwFFYDYAqehvPZS9i70Aedx69UYU
Kk6baTHVMtt8qq+OUfDuJGgfvOKzK9EOrY8tIRgvMraULZBXnu5X/dR1sNBvSWByXIvQd1IGwR4Z
SpqTcgUvUWXfZe4ULeAB+uWCulHnW2g4ZcKGoaUld04mHWeWggStfosHfXzuzVUMaVA+5XbT9O2Q
YGYRXnOulKPbv11zHPHOSapED6PccWrf1AncaJL4dgVsGekGyjJ7rPmFVNgiX+lK8Tvnw5MQycBJ
ylNCxDKxUrdVl6Cw5i10Bvxn/lgpny/1CoTTlFMzPfP4yFm6WQ36GrS2Wp3gJartDzhUC1YXQ4CW
lg4YqGAAJ2P2MedGiF13yffq37fyT6xjdEKmg5N8nr9ZEk7FUPZiTi1ZnNXzMtVh/YGl6Ez6/6Hg
4cHBcqJwJJVdt4GHiWPejyRjiD8cVcLqLsHdcDZsxTL9+REAEEK6KzIPE/KCQyfw0bDjkdQrEcRI
0Q5rj2S8wVOG0xcSqbAhyoF6ragMIAlEdHIHEdGC5/0lIRYq0p24J1Y32nhRykO4ZZojhCSrjoIU
nUzRcEkrCLAZRt988iYTSpmCKQzRlXlloptXj57rIwo/BTcX6o8NwfCIkm1nCO0Sndu/bEbr02oy
5LryygiE61LPbHZEdUQEKHV16COixblE3QGQ2b99Ot8uNDPUlO1euGZBpHa6VH+WhH633izgmlnp
C0jPeh3tHa+Wk4zRk0+vj/DoPEoDxI3HugheVpQAOF7UJpds6T3rnvOoOA1fO8GXy7IRWnegWbWt
490zlqLOcJDvo4Ggq7tBQtM1r42idmpCeuWRHDKvEYcV6KfCBN20hnujIC243wOEIpv2m+idJE21
G0teSs8DkcuF9f1D9qUpegLV7V3aSEV8LbE+K+a58d6D+T0X6aC1ErV3qB0bydecqjD+651DfFgp
KzrX11971n2e8/ZYjsTXu4MncbLsjhCD/pECLHWLt5JEPmE7Ny3cJFued+j9P+mTGCXrIQcPUrn1
W1JE6VDiM2fW/8+s0TQ6TJCoxHgZPCalo3Yuc+PrGM4vdSdt8EcJVyVbtCt1b5Ho23Y2jz6FYwDu
qlUeq7X9AfO04KmOyQkT1cxF1GDhUpHCi7mgR6pp3mD93ouvaPFeNwbU1h0eVc5fLbJlOnUdMj6y
dKMnw4dQpNZ0h3/dvv57/cB5GzanRdmIcjGkN6woq18zlkjojvoIS+j66zcYkGHrL10hpjuDsF7f
H2xzhlnUOS0wjdrD/D7QC2SRsIl9oUy+uueQ+ZwKr6WcTA2uv20tRfcDax6uZhDUu3/cZpKlZO1C
BO1RMAcN1lt/MrNArYnT41nV5etTkOwHvGT87Gqb5N8+KPfqirT08aXuhsIK1auWlms+/28IodeV
UIOVhoKGHyIPqMXj6EdKWrMn1vTlTmmwnpkE8IWnoeIh4lLI2LNd7WQews/XpCwrXtb3b+emAZ7q
KlJVLLrK8p2VoRO5X4OWijb09qrG+mTdIODcaPvJjt9uf4CyM/+PvwelcxFwRkhwIBJTe5TmA4Zh
OivAs7iMHA4qYw4ajd0cZnyNlZHmifYTPXCDsKtRPTE7gmp+6bV4PlAc5olL52hjtuSPScTO1wMa
xxs6dlrpwnSElRCp+zGUCYbzs885EGNBedVoSS2iczz9+ZijLocA6BpIB4Sl9sH48WSH0+CqHGCh
I0mHSUamC4BhzOiCIvO3aRvVSRZpL+GBiLJmffo8MtIcSGJN+PEK9R6ZsIT/+pITXBeRiSDldr7M
w4PkrBTE0la/1TtkdturCxoWzPuqpfdnxXjO+xbUYacDnIYmLEEIUGpGXVzHlcTNJLBkig8OBQY/
Ts7q5sk1pFn6IILtYgB7/gT+XK9xAkdF3s8oDJdjsLCl5mm7I1CvXTpr+E0LF3OKoH36BEHqKU0p
+xGE3Sd9AzxIuwg7JL9JA0ucD4W+2grF3kHIjhSdCgoVxq/BJT0NI1vMWiye6+mdEGQOT4OYC4AY
cjkJjc0ru3CElYiLy+ZWykiyn7Lek1AublnJVrBiuykbzMPEA9i3oHVIocMpVtPYD4hvicjum92N
G83ooxlap2YDkEwI0igYsp6pV7bVCsHNTE9QRUktGG+2aXQqOXGEXfTe+DAEX8LyvJJTjuePE0tu
dKVOuZyq9eY3q7S6ugorxO0e8RAhUraWxrkWY3F1MdjC7CKmk2eK7/yPi1qDotZrq4+ZvIcZrLTC
WGIC8L7JJV5r3t6hkw7pU4BoDdw5Ph+FhKAptTn18xWbYolP0E1SGNja0sKqi4eSA38n806yO8I9
YFWL2/nwdwn8jln5XR/jOZirpwufbQvicoL2+B77vKeUlcrfLsRbfi1Zvhq22/DSNwJnq0v4N0oX
GdhqXbLZjaUQd8suOAl8MDjPpa8vUokjwfgsPOwY6Qngnt1LoVGB5gZ1o04oNb78zqE204N1oDBb
/bTfphSEHkocOgUMjdK7BM7SrlXqF31zAn9d5cwCibhMPcGRhIItKgOvDqJSX52cul0lIRG9F+ZY
BBRyNOsLbWzfvn471NcLqCeDztqKOXYgH4hTVKBhMDRD0e0x8Z389SpQnxJdds9oBerzC/K10KtO
QLvf8FRKF9pcOmhAwcNd21FWju7O5lE2JOaHA+L8PRBXtbjmsXsGrmH/J+zAIL8TfshIugsxTJRk
yBK6g+7jGN8c2+iEXuhbCX2PebIv//R8NZ8oYolv/NonDFOWD8xXGerx1NozZIazY3/k670d8pFH
TF8YqTEtN1Dr2XQMX13E6YVec6EI0GuN77UYXtzeIY2810kCE1pSAluPJO4mSD9LW3h9+2XzXgEk
a+h11rDbTGOR6idaV43r56EYt3UnUsfhsHwm37cY8ayyfZICazQG1A+XFeVcQFA1d2lh/thHCaq9
Z9nn5MqXXMqSdbDgTPmOsM1OJ257h/T8lPw/PAV0HZZIpNHPBjR550Rib0ZjU7HYi/jV5+9avLUu
GR7hZMQ26APg5uWmTN84Sb+8L00QAg7xt1rn4rwfMVqID/bH7P3B2qkbMnRRfUpO3lteSKi0NUlg
Ijnug0dKBPxv/jbiQ/yBYgeGtXwjMh03Ofa1ejvsMdqxO67KhR73HnpuqHzzU1JyC1YJwauidNno
oddZycLZJgvYEd4hXmM37jmkINhKhEHUItb0dOa7r/23LaucBOKxOvMi0WI0noutltY+ZrRO00lk
NG6JpDhK8diB2QzgOV3O51t5KLkdXFTo0cx/v6RZ7HRcqy8lKTYg2kSP+cdhJ/92kRww9WrWV4fF
3cMZFtNQpkLm0zr24Pxyu/9kCZRwc3r+0NhEMSiE+L34By8XX4xwBrhK+0Q23/ZvI7jNkCQZXAUn
MOE/w7xcL9dPf4GVJwFLp+ZfakgqpEGURVgEZG12IgTgE4L+2noOfab/q0CiYEUPv/vWCdmPkIY4
GAyZyDg9RYq18hIFa6AmakXYRiP1dPEUgtZOVmmaZ6Dhzh7kXYSbn4uZG30ujikEbya4JsABc+Kt
xCJuLk4nADyaIjZ/ELwwwhSIdF9PLQV0p9Vz2mMAJff1YMmL5g3jBYv6V/ZTvk4ius5w18TKnGxb
OqZEm/y16iZvxZEu7A/QVlytn4rfIjre72iBKbbN8TfENTuxd/y2zCJS5KWDR9gElaoqwO3ygWjM
CjyC4M/tAhImCDEdyI9X8szzt+j69+F+b3vydlnxF/YHNlC8cp84MwMoVzrmxIfgWe+26ciUObRR
ZGbgpJO5pCSA9L/++VEd24Z4Pws0kfsYtQ/wzcgxidP4QiDsix/oTkDW7WhImxU3vcuFA1Nh5py8
zHYMiooRsfPGwU6W8uLelS5eIyjBetkB8guT3O9e4J8CnSD+FYYvAcwCLpD2NiSX/JmSB9kRg5wG
EipGPpVr+1fJbu59fkEQ66Yuk/7Ygu9UGBIBokQ6e8C5uzspnfxUnIBlNzomdiiP8XZYHt6N1yoQ
N6wDUlceIRABPj2b737M50q9/L4wB/tDfU7/kWYgQhKqUg79dmNER/Ze91XY6Iege90OrtRu/F8F
b2p+s1rQgPNj2bAN2L7TA7JHH7HC0FOnKib/EdAvXqvaqaqTBHx/X0vGiYbsSW1bvN5Qo2yh+gxa
MoTUxA8Q/FYKrTeE+ErkzUYxKlfoOSRGMNQRYScJ7l0GG1K9HHOlJYD6wdu6W9CfFCxDhn2wnnW8
vC1iD7kB0Gne4xQcDlH3lrQVmTmedqyEu+0uwy8zNUgrkkKvmp7n2Pd2wrKnOjYveHvosSZYcf6m
q4mS/Q8BWDcr6E96huzlZam5h+WJ8RJm4SbxACsVwsyrKHKxPlQpLgAL0Iw1UOWufvlVf0qS+1Bf
u/9erar92U8VSSjgNNc1qkttmBd8q9iNWtLctjcQl9Dx890vLSjRxS1smfkmSh9VQM+B841ZSv50
+9nx2owymaurDm4yYDigGqk3qKKPczc9DMrLcLYuPFjN6TcNuRjclnAftj8Y4ABjnZ3EbKV4R4ZQ
h3slByz6nsQ+ouShv6S7xtoShWBSkqPBfiLu0/DJ5O8mS6oBXyljKKhHhpaTn0m5z07uqKseDJA3
BK+qTq7v78U7T5U0Nxe5xBrGX78JRXwqGBuRNyfI25BBtP1SrLkN6S+aqdnpPDzLLo5trWzpyLQ9
CMMCqgTF55ooiXo0o2n6oOR6gtE5TduGt+BfjhHIzWHtA4Znr2Qy+TDQ2keu9mo3o0GmP9Rbmsem
maZwNQtF86BxPNrWg8isDbwfzUM0vyPGSSMHBFJuPzoCqy8euf5NuVf7RR4KK75FxMz51yZmjPjV
t/JI4pH7j4XNOrFdD2u/OUAhBu2UFbGgLn3KKAj1Hwx0t0g9ADinoWHhb2BqHsMCso8zADZRNnci
toZoaJfXd10khrCqPItOQKQ/JlHh8RYUeDCRrD/CveO0GdTxv5AJquXxiuh+GE766wyCnEPbjPOh
XHpo/umYajo7z+Hxi2i/3qOLO3vdQNirQ1m08m1AlKRF40zt6UilDbd+m+yxl5CvFn0Ug01Dqabj
GFInQWQL3K7pnFRlioqU51pFl+GOk8WIzvL6420vhX9lSo7Xr7uFG5/iY5h7cy0C5j8TKVP0kzjo
EpzMj+J8CvrOoWw/b63E4r0s0pMPeFNGlxpbnYAbXdFs4w0T9+px4c4B0F6W7R9LVaVIpRsrrtfb
AVwDlmrwvNZIO7tRuLXpU+z1i0obZDSpJBJYgY3F1t6NMHDFJesoeFeKDsidDvJGL/Ag+fJPIzj7
WCMWzOE8QKim1dNlkh1FswHPDc5QYd74IWkFuAleBIS+yqukguj6/vMV/QT8vPVG/8SRAgOqRXV1
5xesAqGDW1IQ2PenfEBecz/WwyQmt6EFCdiSxMhr2dnPujDiNwAp2lAYE0KvEMhBeSL4xRQ1l16J
S1oSBbhhrpDj+70Lp0OTAINTr5vl819xhc5+rRRH0jrvOquoVp08ehJ4h9Jma0JqwxlMj7rC2Afs
04NBFUfolGHC/nuv4SqKG9p+1q/3C9760PkmiLLIshUbN7Bm6DQZF7uJFYQ19FOU2N6sUWr+9Rtr
BPDkU/JHsq5VT6+GT+p5cA3tyYvnfJUg42XuDHYfYq5YiWuWbZMce+tuJeEv2cs4mbSPNrtwa8n5
q/7SVDn83S97TpiklKKw+M/91wHMhKAx1HydhdW+iDuGPf15js32YaG1H7jAgwzMcKEVzxbygvkc
2OK2AZN3mLX+vEp2V7IV1+mGC+yZi1AVt8RusUBkoaggHPY7910jppdDi5EafEH4tBauTYKwslvK
I7mmprS8v8bWkBvEO9kY1eKNp2rJxitWqrncRe0MsH2TL4/rPQZoOAGobIoNQ8gKQgTn1Up7gS8p
nex+RLc0B5lXH5jnvhrDtwocMLIxJuaCw3Iu4GVy8GCVsRSEKr5fnWFMHtoTnyRfjureajUaXpmd
LeTOdK9A40tdxGpWrTtssbpEdItseGudLQckV2yXpaGcI9CHJUzSOo+uBvkeYNUzzDXWOujMzYi1
IaZmWTHsUoZNaREpLCqFo4CtdrpUKU5DW1Av1XXrWzoL8Xn+ys3l4WwT/rMOWlNZyOM8kpAY2FuB
PeoTq6uy5HtGdq99i2bzkihZIUf8NbCl+wEYUxfQotQNuHXaA/FtXZTMDMC/6oLd/MLPsR66Hh24
Rmav/1T8O3tfeWEhb4GRKY+9p/Qxg/6VgxVRTyZbgoxuLvUbORMqGE+221nWTqyW7JKQIlhDeiyV
VBhonvBZciwsI9CjmEv6Vpm7BrlOYZ1PLEg3EVIfLdjtmwqsYHEa3IijyJmYSwDlr72XhYWrCHnF
HH4n0YR1by3JMv78DmQ6YSzoy0e5DNqnJ55eMXSUv583CjOHgPWzoPo0ZTCEwi9EUsXEDJxqDO5K
G5ylMWhs39ZC5Up7MdpZQF76UJInDNJ6tjul6sFz1MXyCvmepoT/dGqs+HHcg+vYouZ9GbUQSgTt
Kq96mquGgGR6Wln15ZI1yIJG7CfFbQU6fj2YbTtG+cTCkYc3i5dddRuFUDvRlmSZ5obkk2TG0rKw
hRGxtyI/QbDRM3am7Ws4cb73z2ZAgXvd/DVhWGX5bXift8xDf8a0PSEc5cCLiU+9e/+WlsA1QMBZ
KbXpyNECEwKXas/ZioqQM7BJm6WxLSlUxLj9UHUmfEKSJuQcgpBeL+dk4k4a/1zZWxVynoZn42EF
MA4idXUT+QzuHell5vWkL6CKZQbDo49ynS4uHiK56+EJjRpyQZvYYW8LE8ZA8dUOQuZG95jqJttV
8UiwKJ5UKtWhyrfwwXVHbVI+yexJ2fNzyrJQ/aJYM5I9qUkfbYLR3XhQ1bD504RaLQwxrk40hV9a
ogzT0JIICGTKIFeCgzyky5nviWE7Ma4f4LwRpCE3DYYKOdw21yb0b0BMYkitUFSq6RF9ncTy6gxp
G/DzFxkCIPZLdFFvjG1/RUsJEetzfeksjTX433c8sxYfPJsYt2D/qILVx69Ehn6S3S+PqT71A7fM
WjlOqny1xlG8oDvJAOnRoOu89JQWDihfBzv+MAGvzxbeNmcvw+aRgPpth6rzNv6wSao+Tc4w/TGp
Kr00tP20NOhnLxu9dGeV5EExRpUO3YPsZNlOL/WyMXLm3jqqChtrhCsdoKBIby5EilRiImquGA7Q
6oPpU826CYqYE3p6dceZjy/vr/32+t3Ufh/x8Y3pKl+UeSY+r7sZxRmf5P6WCclJsFTACgFgdrHy
DucIwriKWeM/VfLK7R2s/tVJLCTnwiI5/SBC5UtCZOE3Wvsi7T78VHXHBfkZ+dpwMimXhp7uqYuk
qhJVM8OwHaZvDxup8F/hRALWCaNxrOmMfcs74FG5TzlxI+KmTCHElbduJsS+whmTYdac4EetK9gq
Ded9fkR3k4uRZjZVx5TZH67j8NLdW0FeYcK1B3assnxQYi4AN8YFaZNWedzheiIFv0hdHC0miXMC
jYoy5Nkq1kk4ps+dSNqy3rYf+E3dhJm6duPNuNzZBYuuqWbQ447b7HNLpkZ7SouEXDVXNfQAfF0x
8mQH+wSi3Mpv7ob45TUiJMteJ9UexNcDHgAyWaTMg2zbq7vXEskUGUzmynoDXs+Hli19ztRaRjKZ
hQUdOpbjPj5R3NxQzRvSmov99IEG4+qfHjgWo0WqzTlIoycQHnqLEJEGoK0jTytKPfcslZKqC1Xv
2/wg17yQg0g3Do6wbbthK6g8GPPf8ob69JKdKosl8xiHcrcFuHfCqiuCJlqhEcBWVyrxC9xW+8EW
E5PCNEv8ccO3tPOZcsPWF3MnoogdDiMP+8iRBXYVuLTl8Xctl2YECNwIlL0AR6PClMHmBISFL32t
ZEZtrXW1lFjwIMSpUsmFs4jPmXhhvJsH6wt14G9yXUkVXhzcMCJvTmvp9z/Ifo34eUMMXsP5jBpg
HnkxFkUVREg1y22yRZJpP8F2Hdn6rZ1GPMhoBAMl/chHKt5D0kOnZ1Z2EwYXcuSbSsHO88D3h5EU
gWSqmB3tYsb6H0MZZG8+M6nL+ZclLrxt7vNs4Frdzc3Qp4x3tjKxrn59A6W39w8qURSL0+famyW6
AbvgXMecnKxn9PXVNxA3m9v+JTS84wtpy++3BglVEWsjkCUIiCzIYLcZ2kLkwGSPb9W5vZ6eRASc
5ZR+xtpZ2D4WdE3AYD/bmvOwfmndsblp8+dfuNo70MmU7xLR9YYKIyg8twU4fswu1zmnV0GXzMng
m1IfwJjg+rqXywbh/ss0wB7uwQt11LFWmnIzKniE4o1//4GQi9oP+/Ak2TWHNIcdV6qKfrOGHNNu
+C75IaOmrPhCfF34xmGtR+94TJ3le3mkCND4E25eaBKLl+iFKriMJBIdbC2UpFMgbxdthZo5SDNc
dANasguxUjIUc0KFLKNoK6TlTEiQyldWCFHtQ2F9DgrZDNlTTtG5xPKZxIwa/cqrNiH8zk+1Oxus
ABBSNPLOUYgHxQErtiVYlsDRAfnqAJfmbHvhROEXezgN/3coqX/rOOeDnhkQF6AfaoLr1Oei2eMl
ACFeRWm2raId77kOSSv7Yal2kjX76IuxHj0rCum7+hqRYMb67NOkn7+2gxmACmQ5/FTzyoDEJU+u
NSTKSQ5Ix7tJTIxQZy5/zrbpbGRfyD9+lAoiEAdQH7jGLcDw3QrdqOMzpUOsFS0zZ9CmahfICPqO
yQPi+6dU7pgZOB5BIh2l8bbuWUEyguAGKonIsop105yIIwljYfU2KrSdDI3jScsn3dqj09eAahhQ
lfjYY3T97N0xOKRAX6kTaZge13l3Vb2mV1JiMXrnXqJFKsn0AT49PHgeLTIzMTCPEGOjgTq59qPa
pjW5RrmIkHYjLzynTp7GNVuO0dLXqwnO3jgQDUYUEcLuQfRDA6Kf8dn2PLjSmB4tIncGsaYJ1OMt
QeHz736HGm7sHojDdVcN/AYPu5tfgN+FGAhYRGAQFVcj4MY8c0nGHCtKK8DNKgLYW7N5M6GoWoup
aizDIIiNm8/uUMBtfwAjVWurZRnViCj/kW3CQODYhZlHz0F91oYAB4gAZbIJ0UWI671AG6gzZsBb
OazRW+5aszKz1FDSQ/bVO1ZMN04iSq/iDyYpmVf5Fldi47p4PyV6odmLC9x9GOzD3G1WJ+k/OSNh
q3nm9rsL60Vg0VFmTl3Uz30mzDImkn5PBMBCB8h1XWOGeaLrezKeKD3avckjm9ei8uMzjd+ms07T
zN663ul18dwgbrSvq5NjFShXPjWRGnEolQT+3Lwe/AR2mCg4pxPYbVNpNGInqd5VUInIcxtbkRyR
bqRSG29oclrpM8gTYIT3JvDu1f1TFR7gMnQPNRLAvRU9OsDos/85CL07+cgvSFvWIR8g5tWCsjdN
F8OMqYTygv/6q/mkyNKrLfkBtmJ2pmebICCDYNqeRIcfzS+QV5eIz37r07z6t75o2o1Rx9qZ2kxt
maR/blRgsgoegqKRBXvCdmWlD3RVXSprCShvgDRJvabyY0R+N3iXY/BU0SC+/uAlQx+/lcmZAh36
PWJ4s6SfIwmM/dYsuuUljcb9nd16jjqYiiUUUPVpDZprBYc3UTkMWVky16QNNiJxaeA9B7b0z1e3
ty4273F4SOY+ij/FKqZk0E2KFOdgf36WVenUviFkBOAkLNRd+VXDGrj+R1yVIQnD3T7DSSpEatFz
IGE1x/KYCfrxsSwc1jKwAEyeviU6W1fsr1v3vOr4y9hdIU7E9kbhuH507kF2WWQdZIuQrz8o8W59
+1RLOI1iWSyaxI21VrU+qBHHKIle73NT1k6I/lmdBBiDekSZvAOOm0QLNqvnMQ99JdM4Dyo/vI1F
hQBaP1WnH6ZS4XQ3nPb7ONtUaZTdWLAu/KiXW4m2vyRYI431Cd5jdOOymv4gqhdZPLHnuujucfvF
cFAS2pr0xdw17XWV0h/otr5P81wn+EMzuKBTFB4LlxFTqT/J5CGVyK7gWyUt37LtS1EpgIXebDQL
+K8otJAE/cKI2ks9CVJc+ZeMRS22WegF7mLfmVKuaT99FHqwq6qy7u7yTq3NHETOIa663Q3jcGuG
uzOc/bI0idrhczgS8k6mOdU6/hPHZDf1+byAHNHYcFUhA8kQjondgzj7x+TwHPes1plY6d5YxJiB
2Lllx29bs9fTRzJ0FGaYzeVmBHoDCavtJlcjg6wK4RICASUHtL38M2xQOgL4uU3gh7LgaXbDmoIr
V14uoBXd43s3qn7V8Uda3ItStaORHKGDth8nMKddLCLq+dKjdxbkugE7MGk5Ygu68qu3Bd9nlQnB
FG+mU2l5klY5A9VlCbG9g7EBu108PmAEhrLKbLiijb8LsrMgbsyxHfBPkWaLGBkp3EOFxBMY71GM
+l8qFmdUSyGazvI5dJPbMvlhSdc6SqbNB8rXbtvRFVteEcVzCUI3miT6isrlFCBBTwd5sXfDwTeH
YJl19aTeYSRFWR0ACMuGOgRq9nKPAfbzKqQS/oKz+sYfvojQ3QhHhLo2QqQ7uFdqvDDEu0yO2fEw
iOEDaj+4xDjO4T39mDOkLA+gr37LpwKX3szWfhGORiJL42gFeWo0yaOS8jidGlW+08b3Lu/Zvz3y
3tZmXMsKZPcBk3TqtuUfZX6QyRJ3oivVsDTR6VbQbTiptMPqy00W2mmxG6vutQOsRR0RLtjx+sVq
yshxjHhVASnGbWrWDb+8/GVa//HboHImFhNs+GwwAR6eDo8usEYxo+hT7B0yPLGKUYyhzXRODKsL
A9AKj0FDTCePzST01bCUFWsryKNdMC/YA3/ruN1/y2j5rVa65j6paDZcnbTFNCIBdRpqXKITTu+J
5+yn/hHUBdDeNhIxZyvdC/s2EfsRwfjR44WUEEalgE2aP4Ym2X7ol8kIl5bMRCND9DXrL++49WtD
aC+RtrJFieKBLTG/v88TL2hT8Q11y2DGsP68jyRn8rWNa1PFAegYfb+7Rr97FjuIo7vPp2inTjoE
ZvOFphqQs2KFJ2EPaIH1PQ/ylJMJAoVZ2Mdkx3d4MKublS0PJqIHteu/8cHQUvT+Ibw8cjmU5JpL
/0j9PPjIvKDKr9gkiF9qwxo1YVGMFA1f0tGtyZC4dlgyQiVIpoR+xRuenLsM1bjZ/n72+BpsWGGa
HeJFu8b0XBo3PDSXoXybVgQLR2YoeYf2uJb+fj2+Rk0Am4ubhXFk5Pz9/3p8coj/5DQCxGV4pjrt
W9xHilzsMyZtHkmfm85JXWjpyXA0RXWTHpiVB3U/6j8Yd2N8RayOKg7yff9gCj5387BJ7C+DRa6f
ADaCmMS5n9YNLiidWNyuNgorrowG6U+6ahQxUvcLDTJj30A/+UW94BPndLZ3qR28s5xGuTbQNa5Y
A53zH1LxvkN6fzNmjQZ5lsXvcQMRkpTtTwIhEtn5CjOrjueDluhWcNnKfW7M4JDA3exWl7dP886w
ew41UdyDoir+ZZDz+v3yGv5odPDaKI6/rma9X4nXaGpX8SQPRExF/CYOcQzs+sNiUUKO6zQu8XBG
P/Vc9Fp0i0hr6GES0vBtNl1GMUcHvDNQev862sGkjhNxtDzoKy1i5IacY4xHId30XWGPpziCQzks
ekMCSEpl6hPrvH1ymzR/JRyGrhJNn0SUiqSJOymrPGH8/F/A7SKSmu+EqbdpqVgH5PdWy/J+lrwM
CxSronxgqQiBLrCoOjNIttSGrWYDgR3z34ss6GTOTSx/QV03dCK5Mvz82WVnrF5tAgHYPdooZrhA
bd3eKho/LXsg6IgPmwIkvmsbt7dnudBCTqg56dFCmHYDLHkVHl4k0MgoWqC5LSdL+oqZGynFZ3Yi
cyJTJ7DNjO9E4ZxIV3SSs1l6/vx/kW3vORM96ou61bS1rAfXp9FpDTv92WIwGWv2T7PZ3u45Tp8U
tNQJy3bPWBOPVd9auX1SPcgqqDYdGlg/i5001mPajP2gs3es9bqCRflMjHlLXGVYm7Lto4vaWOt/
s51rO/Dg41s61kxLnKqYXtz5r1M7O6AgCoWuIs97vlWqvLeplsJDAE5RPYzuZQVA1KnwCsIcXDUt
sRDKuHFf+AcuYL/Jvsx6HSq+0oe8THCBQ2CQUglURbp5FuxZV0c51tCtBaD63veQQ/yBFYDDbT8W
OYHXLoqgc5/KgQBipUdyvM49BPx2DTUBhgMmIMqEu85UYwzOqPtGSrsCzh8J3IJef09HIFxn9nzT
tlm7koK847862xESYT3ZJwATZNPYGTcgBW4+F8t1Zzg/ev9rLAzouwlRVLt2OF3ngLahAjIfDxgt
g4MpdrDw+dVV0TGkB4K5qDisJSHMxRx2ra2EUGfey6NoNveAmqwY5cWxwHTk9bHh9rUV6p+im0v+
smIr/g5F/w+oeJoiTm7JNg1kn5eFRZoq97VVhGNe+FAEs7RqlllouDNxIAFABj7iYqzuWj0IeDvN
UcKStiw/ff4mrZMhC0/kgFabjjYuDxnyvCbJNsCRS9VpdsZz2olzuT8yXyrcwQt9iWQoUe8vgOby
9CLzBvmsPOCguDJE0p+07we7CAwhQizuRQxhZ0Z8BXrKqB9ulOPwkpEoj6HMCUDCc2R17IUpz1oc
ns32SQ+ztD6RH9p+V9eFOVZ6wiYW1gof60EIzLpDows+dS+cLHhvudNLYyzHshAMdEh4XQSUrv7h
VEzH/9M1ewJnr8II0LLHATDdQmqwDjHthy3G5VaZF/A31xK1xsCYK6T8Qzet/rYsm+VMTsPTiard
DIC0rzReUjbr7GR0813hbz81bAXv3/kul7lLdcpe9PCqZLv5wjIDWve90UH1d1bheOR7mC9NAPhY
f31r3YKu7ZUxrzE47isQ7ist7+c/bAB2r8QMKbGio2SY/Not/RYVLDPtNkR8AW6sXAE3ORzzI80h
W5ZE3bqb6K/cb+Ea0RtUAIJHA+7JfRToVoYD3gMLBBra4g24uiMowieY++fNsu1r0fnGdyw/dshU
kxlHf8kg94aCmRYvNvuCNWsVm/aNvUb5CT+bg1SctDq9THQcjQIP28ZpLGCsxM2ekyjx9Z1pUv1K
KF0ZyVbwvehOyyxzW+jwgobkP/tAJilFX2DLKqWVDpZo/df8AqlxhaoM4tajlFn/AHfisX9KyS/l
FPgIWDwHpXnePVpTQUyVAhuHQK6n/GkvEoD/r4tGWRY6ZxpQpZSdmcWgMsqH1gp3xHnuBhEpImYa
mff5AQRxBoSutDYeYUhdacymDTynjw/rGFH7UX9ROAb/TK5Do65fhCWfb+6whQv3ZsQ6HAfGMBCx
6UB2evPcpWB+7VksXWDBWKqetxRB5CgZXJtIoofN+PNM7ucsRANmrutVIBEq+JALhDCI86xX/xvE
58v9XUW2Uw4OH4yymhF+4JAxX8/JcW4GiF8VEQEVyizBmydYZDvGEIebFd9mV0nHGbg4OGvQbB/9
8uCkD1kTy8CVd7f36VdT9X8d+krfUlfwSeqbIEGqPNdwBOb07bmTVsDD0ze/C+ZeF4wrwQCyDIXo
LI8htiQoaGl6tzIn/9AkTEXvxbJraJJoJj8rT2m9bFnuZSVrxz29C2F0gGKquE/n0LAwCA984gUb
D+G/w1/TtO+ljr8fB1IdiBhNqLzc9auzGfdGnDiXa1UkM/TSosVFRMLobw4+/UzTxXSpG2BsRNxN
0Kp21rcLw8OD1/LyyaFfb/PkzEohTqjmFizryn6xCK5/l5r/ik/y2oiYduN1SJxlZV+lihKppHT3
9Afov/zd7slW1cH4PG9NCO6Lr2Gjne3k/psp77Wci2bn/7wEDuTlkPegf4tvIyokav4cnqpk61u4
VvholsdEQ0pPfei3MEKDyS+RaV4P1CPMu0s6RylVnMWBhdbdLPMMFCQ2b1n4afv5nozT69Dc42J5
kicc78kneRxkX2QUydOl2BH9cyPbszd+no4kYUpVDjNlayBHHDkBZ0+IbWyR6BY0s7m7kbjHfOis
qjDIiv9fsUeUKquGYJZgIWHVOSe5B8mEy8sLJb6q/rmwBKgQdkUZ7Y5BNIWiWjhEGDIQeuFPa2OK
tNPn2lzQ3LmEJDfS23LIj5Pr1/hmV2IPXk6p1Aflc/B47WYuOdbIw43M5Krjwj15sAVx2Rzh1AXL
zf6FqOful1VEC303J73TzIpIurx9Mkhx0P3UhgaB0PJKv5cjZ+zvolPCTeB0vX8UKGv6p7rAi8mu
shfQX1PF4JEt8Q5PK9ahbkD53F9/W5P591Mi7uRVN0GwLJfBDJjLT1+G9xKVGDnVimN1xzzRdGR+
+LV3qTH40xcmmL4TKD0AP9rhBU3d0LjfwFtIOASs4rffBiZ1ucIWf1aD6O9PlgCEXuDH4Xfy550K
2Vf0odOGSzUoMz7acvoL33Ow2jNKy+W3FRls2Ga+XBYKkTAYYER3KRr5vtFJdM+rNbEBcqNAGZ6s
4iBYavUmwLvJt+yNYWaAL2Z0BGSTlzEz73AmTY8OdDOMRZe0pSO425CVtN1V44ZRGtLtwneFAPUk
d+5gaQt4Ym3f8CdQ4VxhwIkGTSTJ4zFnp6f8HJfRslVg0xaMXkWIZfgvoyqkW/+vdvgY1cOdsCeR
tTlgp3mKemT9wDuhGP+4AM8iYATP1LROZOfRtAc/sL/WySy1A1R65tWPr2I/WyZaCvXGvdelm8y9
1RBGgdInWZy4mz+PLvGmZAh739cxV9tG4n0mGMKAU7blxtmAz0rLpo5NQmQwnlr+EvA6d5tH+wTB
P3oI8JP/F2GFnyzFuj6E5oSfiYOcKe0ydQcoq0zSldXhOynsv0Y2c9hD5glpnBPPUop8bERjHQWi
Qr/XYTriqbep+ubdkJbe8lWdP/BIrh2nF4ryDlVNkBSpE0uo3v1OAvryVUVsK1x2xT6Yda1Lk3X6
A7V7Dc3VD9ge79RJRY6t4JSrT3nRg6M8es48/k5UiIo1gCJAjwgr+T8fcV5O+CSGD7Cz6cQWmL7a
if5da1crbJZhFLee49EkaACiw6zb8Gl88vmGUNIQV69yYVcxuoTPoj1WOOehacWRZdh00dOydGdi
20W9bYvodJpW8K7MfUfE7mvCBNXDz8Qcyb6EIaUco0NhIy8880tvEmKzDueskAHdLi7Am0AN2uBr
szoSpeOniatvHp1agfGoW5Qdtb0pQBQUZXBgV/If21MAMM51DI0J0F/wOOlm9Bt+2AiBT0DIapvd
U8j1+VTwJayicAleFOaZQmv1akY5veprCLJEbUB8+zq4qOxmcuqK0CQaysByIhHd1WIarc+0cP7u
r7TODOuuL9KvhwZaQp6CFJnQmzH9nv8w4Y4c18VSaL4Nu6tvi3eh9WYcrS2oeZnG7Dz66r543hkG
Jjl4KTBz1PKWVlMGoXSXQ/ZQVrSBwha213PhnhsPsosbmNN72o+gA0YLVnips1Pq/fePZlWu6ubH
UGYUbeC1fQqUpEzkiRCmgkX1XeypzV5bAjAll//AhsSDcMnFTghV8GExkFYgjfweH2SYaOU1Yobc
wzix3Z7UusP9z79OehENOwAWJDGQFgKEoEBdrS3SyGN7FpfrxpO/6Ckuu4FJrax5chs3g8Q6A24P
6JpXu8lk6IJ4r9kUzRY8KlfxGxR5Ii++orIQpxKo3UGqHBfuMFA1siON39wECkLPCfc+zISdsNPu
RkrU/PRxsfldExQCoTsHVPnK0HihLPRhY2p5dZZvzK88wAsl5/S85EojpVvEof0CQnujGNd8i50b
fhr0WD1lksGItyEiW/xl3Nur1hME0FO+ziyw+Ler01LRNQOVnfZ+GX+vwNz+lj7iaMnh1vJ0+dM5
QbjCm8vp4DObFXjX1dgaidxhXF+8jnIbD8PNXt5qNsQtEQXY2UkUquQAxuPS0SkcgGK5rNw8MGOf
HfCPbUOh/170PnGmELk8nsLrkJCvNjamz+QoKNDT2jy8DgzqGpw5+LomGDcdgaWhacaUtVB3BPu4
R+VTmUp/Wfv36d46vcA7mdKk+Tc2V2nrNm1rgNHjoXVQDwKCnZA8IrFjxl8sI+TaXiES4HyQkLWs
hwO1XfF2DYXgOkm0QrBo+N3pWBKLZJBO5Ck1YXCgn01TWB8iWafx4TTwqK/HzGXDsm+VCRuTtU35
mqIcaQwxZHUqjcnakQvIAY5D/Y8TEokcwtWxxqYmc9wRc8A7rU8dwmbgnM4TYT+C99ksur+SUFjD
3cJ8lPqMTypO37Yf5Imxv65o5CzeWBwm6FSoV5O4Hjjmx6MBBkf73bf9WgIL/jzl0ke6YrUJLXFt
cb/LYqbg0a6oWSrqAmysD52gS7EyWqJpIPbfXLrX0z0E53v7srJaC78/98MAsvDouf6jkt6kKybp
0KN2fmPqS5VPb/IgCCAZhCNM9BrwyHOUwJZ0DU9kSMAsAHBqqT7srhVgO//cQA1myJhPHzRjInRX
UkCa9ih9/XHly6Jtf+S6Tn4XECu3+etMqdLjdYOMXVnNn5wpItwuLD7Yk720eW2wP6KXxjKwd3Ze
ZFbmKTe3PpmqdNrkW9gQ8cngOcRHf1bFSE0gCsylSkX/8027y50u6BUoz+cHdt3V7kJdnS2oz7q1
AvxfZk+l74qYksvrP5UZDQ/rMVCiBspCbiRivJLHs+tNU9iBGfbMYuHbaxVu5n7mayKPoFACanqM
Qf7+6LwYwNSR7G89DOmqlqLqsEfwxK2HZR/DCRhfBMJPnZIBHrtJ7s0XCkv3v/5iOr+qIGU/RshO
VqVCi5EpoFOw5pHHy9J3YfE4L6R1yAVspG+BENwlWTWkavbKa9Wej/ivQphPD/bEK4zl2IF7mgKw
JvBBcy6IXSjfem+pMgD2/Fbo5xess+RUhvklBMyOqo6oQmSW7VD/z1yJCfYOaLjtMTSHzRucHzuM
W9xMo1QVGJdB5LyOGdW4Hs32xqqSOh0Us3llnBNI5JT9HkBBm6XQ3w9V4CDwqCrGHU0jL2EVv3zg
F5D77eq1wU7CuSCTAD8ba1MAdyc/H2iHMoPg+q9AFDd7SGz3e24cOaYX/B5Gi8Z7T1nkPMcSLTEe
Ast50TSY/3P+zx56budgJlu2O5TUkZ4yiZo63bo2iuX2k6m5h3Z8UuVYsaggwFqsN/Ir35FkcH1i
dx8VZI2ko1zUxgs6WS7asdd31zIIZyS2KI3RYFCEaYZ2/DNGZ1QqreGXqRyC5gQsNySvzVit1odD
uYKZZWlouIL3ticj+0gGtGiq0F7XjAqGPv7f1W7WnUmT37cZb8y/8HNGjxStmplTj21O7Q7ti0sh
AOLR4+V3fdQB8Z6h+HFSGmp9+6rfp88oIwpHBFisTYTwvFcAL7xuSgQOngE+rkYwzCfyFf2ebWNZ
mhZmSvNK9Z1tsnIBubgtbWNQfRitqRMe7wCVZUjGEsjBmBARFcr8hSTe4x3pGnAqhRdo9IswQVqf
wFqNkizWt2RoxVbRLAYe/vLb35ib5k6mvQpAJno/iwH1VnBr6+oYI+1RI1e3TBs4mEriJepTwogC
3ZfCBkP/gxtRKigMpS8n+bfI9qMNrxGWTQ46/CLFvERMo6GSaoc/N/s121O1bWWh4X10EvkxRLeM
INIiZqrH5KiZ5Qbd3Xu/h5W3ek1JZCZOCoA+NJ3hTMxcAAvNWVmWaLns7eSr+FjvIf+goNhLMvbr
4u7ZOLcFtvT4h64wIKGFgTO5VhPbH9+m3LLnFZ7jK0QhiJHxmBFtHLd+eLbr9N4vc+XOjib0rJjs
NwUhmXE03yqCfSqXDJa9AGtbQRao48j2GU7dFyFSu1mSRo0o0Cv9YmMCljt4lCobQ6WpUbznjfbF
F4DZTKpAumEW69gaZe1kYE7ab6Ov1TEyxzRvKbX9gAMZX8S+l7aXorKgEf58HGtkF37ECHmvq/aW
4RMy0WiYbNw7BpzN68ftiiWc9kwGB4zoGXTwN6gkbSyUzkgPIJVE0SWodo2yVhhmgEAy3bXuCrdj
TnzvEXmWGwNl52d7rHFoV+EFDrelR1wDMrpl86bAeZ/p65pQGFmneurVZENGfHJTm2wbPJOBp6ft
kC/0SNASuc3hblWeEc15N/S4s+RhUPVc779cT+c0q03vOo6c5b5NA+/UkWXa1mb/3Mv7YMJEsvYr
oGJ6Uj1s60U8YYob8lZfOSy6TLEiheHpcCk8hNU3JR2dHEptvxRofPuf+SZIXcT4d3Aq7fGaR68U
kJZIYzghbYt1vdnYKyNl7+CvVjGTfmXcVWXoqlCAQHXAR8Y0GIjKFPuKvCDS9dWwHVPc6NetatKm
ei7ogpuR6Xg3avuLia04C71QpkPBWHJhO781PZEmmjIm9o/EM2cYRYl+IEejGg5/v+pWVcfay6B6
AltbXSBm2swe6YJ4Pgs354tixI3Oc7HjCxJrba4ZL6WARKoGe0lgUqDVDwyaMQLCcYW2yYgBPsjc
Gb4MZCj5gyuxjJEeaS2L6+DhIKW/9ZHgCnTOTbMymJI01XS2pg8Cv97TqjkfffgmDzo6/DXtvv+6
FWxP0RwDTwlhlBYss3DeFVm2dXauCsqpTDPn9M7aHa4K20ED1X33Wz2rQCfD9YC1tv1gxskPl8px
YDczg+GiIKUOgMp4CBHzoDYnE9et7YIkon8y6fmmKMdMcK/bemeTqmofee2/roOwLkzbWmzivrw5
WyTx1RObxHwNGkVsyu7i+6iELPDr6K5AMJgbpvuaqTlLExd1qMzNqjV0moduPvCA/Pjf+eXWm/R+
2WCEMZY0XRtb2ZtS4KSiGDOyzkHA4XH3aduT8fm9WVmQDG792ifdQUwv4Pell1JYBqBwdXjZoyBK
ontfr7CbppDx6X9R/nWZ6XoiIPqGvq6bGAELk0ZW+l67Tcwr7S7H4bAzaj50+B59yqnDPqZk03fh
mFRLc6biJnX02jhBI6Y+pOzfLFM66Iu6jFzVzK7rllkhlNkYNtwOASzXwQdFnT+IWkG0Z5PTAqqY
5+QJPGdkFZ8D0tUa7Vhkv4sQQGQtDuW0n4iF1GCVnRUWikV3kq6szHeUE63iY/o+z/voYBvqD7kA
r3rkBIoC4BwYKoW69f8vi+lMALrRsxpH6Ec6efQ58WvDwNO3wvSNrOlBfdKH9zysl5YlrLfg6eyR
WeM0nwap5LqkoajLyUOYj17U43DmOwFoHeRKTUAhHBjuBRN0KTcZjfsdLRvLayQygBkS+CGglgTs
LfHLPaJKaJE9VjeSkIowNqx9i30xDcjEiMz4KAWbjjRSn9GiGkEWBoUQxL7UyNT/Y2/aHezubQgI
D8wRQCPS/OpYsOGfTF61O3NVsqVsfPswU0oXsxI+VzDxCodLO0FT+MpsPUOHmkdtrJLSB8bfWj+K
c2NuOhIbXaFo3CwVd+vUJEEVAePX6Ve/Z30PbWhbLiWzuxkY8AcrC9i2KosGBryH8sy0Z03+ZVeN
eS2yRWw01D5jeDzwpfCvqV2mfPSV8HEpcuQEUxpRQXX7zmOXANuy/3vZu5f30vroDum95PExehoe
xt7aJk7r69B/UxDU0HF121RrlMcDP2hcdUH1uP9LQif/Y6GiRgFghoQBFvsalgkpJDQw0K39RaJi
hM7EGvYwZ+1sBL+CrEGvguFc2521dbYk6RDK/Ulmqo1EtMDs4CLdrQyhI3EJDfk7FLnOYYADbMMt
Tnit4ZnxkS3U0Kjp5DcB7YukfZ1IKWjbSstgGC22vn0I5aZozkON2SOSNNadl1dz6jbz9DckTZOn
ZuakxQPoYTICRwizGrgMGwLKNv8n63gQjQg0kWf0j/dagMJKrSnJJZEUimSRJS2TfWQLsvV/PoiQ
wclm5Y+ZIvVTBFubfeZENGwiSnwNqDhK4OmhXPvLrE6fQLYju2MABAMGCU+LT2ky9mCypnfp/2Od
PXJ8Efb1e6Nv3cejfrbpFViulYNopoR6TRQQ9j5MlHKeDeG/iFkSGr4AmyRtYbZc0GB+5foxnuUB
clgvznjay/XXCd05COsltlnjPvUi1lpqrGdH/jUn60c9Gw4db8LAr90xSRHn3sQuNobUUqQMx7RL
ko5agz5hRFdO2KpxxCbB21DeBYXdxa/ff8FE4brQOorSi4YcPGtSdJ+rJkzm8Tdek4bo8CzPQKU9
Fuy4KI160jiQ1cSHYun85RVps7ClENVvN1FiPAv1io+gROijHCRb79lJM2g6HMSCGOZiieNIePx0
3hnT6UMUg3TlA0AB3wfkn+jOjXc8rORCHJD9mHrH1zpXjLRmx1fPXoZW0LG+BQ46BcJqgTBvZmF8
qz9DT78mimXRR4yLMu3ZtPFTFW9Tx0mraZHUVArRs9AxJR8pCb8KIK/hHno5fpt/cuOcLAqNx+rF
TltL6tQq37ZbrG2O26emJ+Kk4Y9HLO3RH0tGZn3XqNA6o1u1lDeDRGTgw5lY46oypopMPkWkiaNN
diKOZEk8qz7fBLzj9m0flJ2yz4Y5qybfhbB1o6zSr9do3eAxaUTpnZUP7Y4ubSpHw8cLGa1Oq0eZ
ehJkw+Rp5qvGYZ2wgsX5oXG5bkqHdlvb8hS0U1PgACIUgZpGhF5vv4rkmmhcv2OFEaCOHQsedSr5
gwoWEz1tE9/h/o2CSoW/Kzx6Cu+pcGRgKCf4yR/Ieu/Tjpd2tNNXqBF62bdFPaebGJhN1PTItU06
AWAIkYXVMsUIxleZJhXGjJFAv/sA7o5P6VSz1pDbh4sT8czHVBMhNvEI+/BDsSp9oC2dcmrqGKcZ
p+agbWPuBGqdBeZIu0+AerkCTgS/X3Jh14AozLPctVsPHnrQrisbHWf2f5NU9BFAs7u5PHHROEp8
oCUGZLrVHXVKSTlkZYIh7fk/WH2R0wMKufyi6DPQSqBvd9WNaPmvcA3qPd3zJS3UUjxiuHe6/Hpj
QmJcfhSMIY/TvHc62v9gxkMeGzi/YlQLh+Rv0i0P2XDobvcsdkiRmfxmtzzSm1arooIYeSqOwvS1
Ks/b5GuzT4RXp7SQrnRGd/7b4fg208+OGNA3f1zWqslF4Ads5++8COVh61peW6VfV3YWa/ZM9BU5
sMaO9HkMz5Q5R4lKqB2RKvQP3EGMaGlDXMnPY6eZl8U7gBaQZ5U9HjVgFVLbo4K08sPukAbsDeV8
ITdISK2+41WgPZN+YZ0L1FXkouHI/DFFHhAGbVxB2Sj1vODrwdhxPZzGNQ8PE8OY0fRmc1gX4yfU
xOud72BFJK1hX0BlvVIWBiFyX+koPWZlW+PVb287cP6xFa0g/SPUaM9IF0ertMrTwmZeLZfc7r5h
UJp0MWCmHf6wzxDdo4T7Cy6BCizd9mbZjfs7imv/kc1HQ32OAyAxOJAgcDcRt58AMIeeCbf7RWjA
7KTpc8ZU8Ogo/Jo3qygNCHBEXhfV93lWXKcDZmtAI48na9hmD7PQ82zDNvpK+Sm5usahz/eWW8rS
NA3PebvhKAAFsOdWTzcSJDL3st7Te1f/xBgA/vXHqTC36SudKoHghxchXrP2ReUm8wBHPBtPmTV8
PGlLH0chvWXKbTXFF5c/F78mIGYypvLXZ9s1jo2++u4ikq73W6Bp4atSS9VgWhY/iO+wQAZusTo6
xrIjc+4zSJMf2DrBIHqGBWXnPTqJFmnU1gGkomkmNeKgBHwieUh/PKvmSRKyosW667y6RS3HRGKu
E7Ft5zqXsYKSbz7Ux0PH3BwiMgGVHXB5FbU/adBgY17FUyeSTB8w3GddKfXW/q94F1R8EVECjcjU
SuYCKK0YSJZ+ayHyFM83Mphws3nExHbHeIWxV4yPzr1VrdHsRyZ4dBUHPES2aPp72EZBdR0rmw/l
yyg1eGq96mW85psGRA5fLPVexWQGPpH3hR90umKxTp/TklUp4IWpabdEyZcoIpXGThr83Uujpzl2
t5QFoYOGjRmqCM3wwps2sW2F5zC/O5WGCCebrA2Z82+JkWxcJmspQ21jUIJYcsRhNCqcl71wt2ix
YHxWEK0L2ePi+hxaJGN+5HEpCOoEGGITrx0ORG+JgE3nysu4S83zS6REMuXiqrGRTMhTySvB1cOR
wHBearqMAC4FOS91EKshWiBMHsdIsC2PGRdcr4davDzbEc2n8kHZAcyvknpxWUqrXFTYuDa+/36k
HJgA7h6y9pzP60FjwOx5QSZpxqlQPmaFYWRfUeiupIIdZoZKO0A8Ma1PH0LPeKntLol8QNgyk7ff
AzQb9G+MTonY1GkMvs685Y3AoV8FRc9Pcp4qpDIWkiLgwxFduptD/QxaUBWfO3CQWPXidZ4e9whz
DGXOYWHMlZGj6EsgCsJwLJb/rO7cK8uwxkZOsKMZzJuXV+HU4Q8KdFIazAGNAcTR+h42CPHR2RrT
5uBbD/yzEDGaHLiMj2YYVg2i2IJru/uqu4elHNcowzVPlMRhMrhI+hQFhxP8msgDuxw/wRoupj0u
QEmePSlmWMZggv0mjBADaGzmpTmQuQ4xYm6lToVgEZjvEL/EvMmjiXNNmhZKW6bBJtinMRjkZJas
9R608A01g8IhHPJwyKmgstMlJBt42DpF8p67MuyYKlF/QArCgazUuMTsZdJ0odC/VY8MBqei5HIN
O1gAo3nnn5LH2LYR9xsLtuxWqyjAGyBMU7k5wHdsgvXJPDp8NIpPaxTorBaeuXa/0cjW2FZiP6in
JP+pxGaTmVgFDlMYN8oEC4ThIzxPiDNN0ubvJIzuZ1ofgQER5D8gUs0FcYMmoGYuL5mdncB03E0y
p+Yr390WBYAcJKpyqsVTOcetT7kkaHV5bwGVSpGIibX4jYV6pb04GRH1jJ/XOjtxv848KyiXtJ3R
poR5o6N6SEGc4Ltu1hFFhcpPIPp1INu9TZiIRcF4ClQfHuHN+cQCcbO/Dr3SmTd+ryslfoPxiduU
R64PMR8KXboKQHzX067qSkHujKzTzkaMMeKCd809YzhfuKBP75K4EFxUSgfHg2XS68lJAx5Q/MBY
ujbN6UnwlOKFIYSQmJ5XXb471gLp1l2owcGeUo+3b7PuDB5mIp8CUFYtVs2gRrsxcAUFqwcRSA2/
5Qokh7BlyAXmr06mkQ5LlaAWAQdgESAcgC6hoHgenLWddg8tKQDZ59DbaCBKpfEaIlSP/RHy6/Jv
AtrzhQs8kHh+JvzuA8HijXo5bNdRokBoKVO6W6oqYgPQ9ar5lkjbDDFMFQFqd1a6u9roDmA0bphI
lYs1B4+dDs7Qt+o1uyjjHWMab8Kn+mJlJr0tl7Zz+8bIq6fuTa5A746pIXIYSE6LrTCyzCK/zV17
TXRgOhl9OlFGPJq4YUnS23jx1AiDJZKPEHpOI+3/8kSALrn8/37FO7LiYKK7jBxUxkoDodcS2qCS
F5B6O9pMufHGYLFfBjgsHFg6gKHYPik4TvNTJ/3qzzm/ZSgxCSmj5kXsET+3IGXWm/wqHAzXWjjz
0mACwtkTlsZnq7c2+bZU9ejAqYsQTgEGwcoUP7B8ebaT3bmaopnHnAV9v6hAZj2yZw/QEtosOIN1
rdRwNYf1LaHjudl0b0qXlhziwps2SuZBK5tEJrf7CmpQAL1L8ZAJfa//CLAkW6wyDGYadA8+e1dL
a36UZ+7VbkfvY72jUCK6yAWHq07UiLkpfF9DG99FvKutaAIAf6diF3ZolxeXn3um0B/4A4GyYFLl
xlOpn+E18Ctu/QVkm6tWj1VNUV+fOfFMTfbufkma0Ynw17vwmZLttpbLsGx4fxTkVTSJQZUFbcr7
XEHPeZ87syEo3oqq+CtF0xLExUnAk7WZ3z0TyPxPsx4yuAxdk3h/is92oLzcQvZGce0l8sFOWCSg
Ef/ktpFxJt/vLLNZAIEhS62FiP22fSllhkrIMqPq4uB7G60p2OVbb4V2bTOrQM187AfnpYj9rZ9J
Q8SZeJHgcC1GUnxn/ZMQEL++Hs3cTzGQjlkhUzTJicLHuS3VmG06Uy43ZRVWZ7an1KZJSvToVg8M
FtVt8Ods+0rKK44J6j8p0E9Oh8/eldKOctDMqtev4Kx3cZTU9kulAbpfSxtZb+1UX0vYVV7Rx6pz
22UPy8tI6ER9XLnOAxSgSehBF3wq0SA0vn84EhwXjvzimbkd821Vl1ukjDb5apQwhqY/6Sm+DVRK
shwrjKlJhAvnIo3fAcRKwro5OERizyNcmrD/OZIcRhiT6a1ULEfcQ/BXpgcvi8v4FlhPuk2qENxu
t0cb29RflVucnirOBF4r7A6DFg4ZxlfBDqsx17mcFCLEAiQU30IMW63yAE/sU/1iln4CAfuuq87D
S77ii0eHi0K+ojI27LtzDByL843/XdlOjqsSWbCLFrcOld1VLXdzh4UErtzRCCF33V1cz/bNKTxG
6SROOw0zdjIQLfTq5DGVSHp0xxHUf2Ks2xn0whOJzgj4sFCCM356j4tTCwDHqJUw8TenFxFA+Pxq
zQ9Ffg0S1o74BNc2GwjIQRd9gGCPakDNH0lOVB5CobtROIwEvU2o/R4CDpm0/8XgY2OmloK+ZO96
Q6ubIPjjilG00OWcDa74eJ290P92b9A9dp5wEGTzXOAtnEnQr69I+xayp9AwFTyHtF8mA2BqxZG8
7aSQ9+I4pi/i1Jr8riQOubsRXyLsHga/WWsclnwGo5eIawcHzD1W1x4KfsBVcImiy2xRK7iMSwUu
B2oTuXc4d7cf0SzFQlh/2R8sMG8XR9BWSxltsHZuH2HmvS8dAVtwRV2Qj4T2ytgvKJY76E8IgoRm
YAHxdCx+AmUKnSdJDdHr60vOx+ltPIR95s+cvIwwoz+JiE9fwaSI9uz/BMctmZkVpYTeFLk3YWOA
+V3RRDqSc6tciieIMo6QFDlwSJAz9aajdI1hBeVeUfVQafzlV28p0BjS5pVteRSbgtqI5SOEMQqm
YQ1lt6tnFkAmkC4swa4hM2SL1lX4PfS/1WjRVOIUnFZboRPoCsfh82h5ZOq+afZ0NuCuF+7Vd2jz
qnUw14tyaTZ3GvHl4GCzZzwpuDdnsuuW6xgTzNckcPGHxr1dFFdkTprYyEKnHCFILwUeP47OC3ij
4it4PXHSxdZvuqYHPeYgQ9w9ALwAXl0ERAdxvUoCwIYNa8ASKL/0gmQWfDbKMGRIDccB5UNLcIEx
kh1TGaTAJ91JQOOjV8kATf/J4uRGFO0GLbs9JOvkF+xXmtGm6YhYtW51ZLALmJe5ZYv3TYfskIMf
/uMrY+CbRkr8xTfrk/bOcP57kAQnq9B7F7JlSJizsbyqa6xnVjLDgNALC3pGCsz1zcR5YAmPvFjx
kC+zrR92JmPhdq/0NP+W0gOkL6wox2NXFFGzEV8VuafQ6al8xPMT5PjuxT2EJLjzjTOkuSF2h5c8
/06MYkw5bLkgVzSk/1rM+TFj4T1UwpVVvNDDnh+Bteb6KLFwb0+jQAaiokjsZidCT0bfrl/e16Rp
n196NsEA1WINn+ogonaM5QFiP+af3dWXwbnCqu0ToiZdsYHUhiLlo8IKMweAejvIo9Vxc3HJCdzU
HaZd+6pSBauU3jKmEdEVuS5w/0fBzRvFuL1blSxjiEBSe2VK8G642iByxoKImyeeQj7vEBh00PeZ
NKXxkZWe/pfqsOe0SLZ/jOqd2a8Zivmfgcr/zmRNhACd2ykJa7EEG6tP23jPrplAPWNXDPwyAmHd
K5a1wfwBfqiEOVqPxFcEZ5va7NbeU4CNm2qkPsrtKd3WvWtT2tdHfeSHlQ7KrfweGDSYYua4Uob+
7f2EjdXAqloBqivIIXHIWgxkzT8JEUS6P/MlmpoqBmNKMRuBg/mDAUAzZ9+QuTNci+TLd/fmDxQT
5AHCZFolqSn/JmuEXvby0Zaz5oIfd+h2/dKE7GOshK4FoiLy4anSi7//LDhM+hHwsjSqDxNcAYfe
eWFqwMTE17bnuaCd4QxcJIceobb1uzYQ24zj5qTEITlH8yRI+ZJCsmgdYKxg6osNsvpQK8MTwhok
h5OoFkIb04S7sEmJGNrc1wEfAQJUxS3hY8EqBMcouE19RgNpmJ7BQcIFgrJzGuRjHuC45Mk64r0r
YJxsR4cVHgBXukXdUrZeLRm/R3RDQQLLwSDIZEEPjgS3wkFNjnsHCQrBJIwoNN3I4Em6I09W7/u/
UdigWDn3qsm6uFsJAtoFjCGfemdL5pb3/qxV8F371HVcPrGhYje9SlrXUcWs41/Shz0AeWDQzZ2t
/Flv7b6riLSDVzfyDIN4DHF5QQn+ygUaR3sPwTLVqZuuMIVr1VzUmtKx2ALxct7xXOQmpiHDdSGv
vHxTgMqmJHcfvAH01QUUObe0Ie45Q4GYuRqz45TwppNEOG2cO0K7jKy4YFWmQ2CQm5ag0x6wUNun
ocjIp4DcZOgEs60rqg8PA2md4MiYMvcVZq25+PT9UQuwg7dzWKxm1/28O3Ak1L2fNl6ljcfpEwoQ
1QGt2F6Y1SV4nYVMd6esMasEeBvHqyTKtdnrzQzcVDfbya7gBP1dTqUfnJxJC6W0PF8RKqS0S8TX
ym1+f80MYujh7NCLoK57BURYmw4IXceRqjLW4UnKrHPrYl6siqYqez5jdHS3AZShGyI1spHzSZM/
Miw0cHW7ZIFyNL+6j2IoKPgLTRuSpQi+9k9rn+2KYEzdXDJ3QWlrql/6435bLh/g3WbgVqaX7AuJ
aUfTZQCKEhjx7leRwUgDMEvw77pW6k6yELCPDTSZSTjVD7Eoj5WM/7xQ8VrJVblGc45gZlSWeNXh
Ut0j+cYPfU6IklyWrt7fyNY/T2hzD7onubXOoD1x+wZLobMjYvad8iaoOidhH5AziJb0BldoIWaH
MOFn10pVI5r2QzXuAPGz5nG7e7ui3gIjb7AaLubvTeAvek3VmUhFuJ3IpYz0w/llb3qi6htzAAbR
IyWDtb6KxPDorY+APu+7GzOg50bVPqnTOxcLnhr3iAGambzenoJkDuTSzZDH/RvSrX04/9mfGBok
7s31V5hK/z6egqOhRKH+LCrR61LFga505KJ8ZuM8FQTiwM1HrIQiak3XvMFLGRvSaiTqTk1iMnyl
yw/jwjJvymiXKc9bseiyVfKfTxiGqlIwtuX7Bu8D2gE888a3In42Oc++LoYxwnpxV8QMtYDDZzP4
TV8gEahygpRVszDxAocaOmH9kOUJh1vwRUbhTDNpdFug9ZbXNUgHZR8AoyxiiTvxmvkl5dbEporC
mAkZy+BKMkJG0PxA6epr7qK0DfKim6Vd3yCH6g/QObaYNwdjlcCNPRRu6kHKYJgce3aE1HM0Hhot
xNoJPfYrh/J7oEaJNmCxH7FYhrIAvBZqFQLyFqACXxmzq5jHgPMRCPwNf5O2cyqQOgSB9v+jOGg2
rVGBYqIjmadi64FXJ9Y+3RY7rAwGQWqmH2bsRtpdt6DGp/6B96bUCpkLkuk4hHkNdGMrOBCUJISq
fnLQ69hRXPY4gqchCyX4cwjwkDDogJVQR47H9AT0yV/L7sXy4AYcuOdWkcRZSETMObqGJG4rSrzf
6PVfzC3a/KMopApy2LwFkbf5wNuy7m082B15sBiIrG9CLAjFY5R3fc83/fT217CjQIeHL6NggrbP
gWx8bh0s71WzB29x7p0gV1kvhGgrImPVbp5KhNA1kSOboKBT/lxgr2bOOq1FNyJXBjRNf6PaZwaL
Am4uGGx11mDx3HsTxKSrxbvhilmVEhnvNqD9Q4YeiYsRBlOototnYic6IVXWvdywx62iOPj0+5KQ
T2TrMfp7B7+B4mjBxB59Ig71e24prJ2TYQmoyAoTVt5pm3l90Aa7dTEWHQAvLfkbH0E4ZV1X+i1w
96bX/ZSa+yVQS9hxO2+qP99D9JzGJOXsA9YCwzgCkVmyc8u3LiE/iW991Yh6vP1KuHMxYvzev4gq
NoMnkCvNMhlOueMotivBxT+SkBulu0dd+ZYDPCxUgv6bI83fEiGjU24rdcfU4S98x+gXF0bi6+S4
j641CO9jjDEznhJD3GfGpQbilFiPUdjFXHxsajzjIahVvT/R4DaL4w5+m9VR3iQGYEjVx1EQJPoe
Yv/9heb972/ge3p56WdJ0lBoOZr8K/2cpEm4R9kivNCYrpM+W0lo+Oo5KaL2QuJ7F2j3PRsBlNv2
TPtvk85oiO7IKIv+m4x7ybUzqYQQi5r+19F5HCIrwSemcRefpw1qhVSLbE95O9O+9xM9hNQ4ooe+
fvkLvUg2/OAe9+7WDShI+0/zQXsko1d0Jw3ZeawCqS66svAmoSQZGTdRebOrK7LkEXqms4d4VTFW
AiPXbPhtk3gWLaknXIpZOXINqTuuUxeCVEOrZsZsol4ygbUTF/73U+3hv/vWnCk1WnF7oWszRhiC
bktSbEbjFrzuJYKGSFe3+U1AvIPYXP4WoJ0x3FKiHHMRF7WmVtodehjGprf3N6LBr1Gbu/GZ0ySD
PRFZNWa6/X7hbCaFZvQOT/MderZYJCMYTU9jXZYzZj8u7crBBNt8UEX3eXRMz4Ppp4w8yfUmLe/6
aexbAhC6eS51/2X++TxEEo8IEOfgf4C4OPW/+E+h7KFxkZb0w6EET0kryj7sJKNT+65begj//I7q
HJxQUfInpbIOmy+bg1+gsQBo1AmxOY8nMNaC3tUYFDPSJfJMvNM8bmJHUNEiVdCecYymguI0zrL9
wefIN9LkkVKI3OrMVHojU16sxQkUu2fdtfJaGZY6E1neK/Di+S4vqFPw2I7VMORwc+3scmOdOIHd
nPKvclbVDMyzHSSzm8hpDOP4bPQS0DOqd/sF1fQyEPtQKn1Icbm2Drj73yWgfu+Ib0veznX9y31v
2bO6obyHlZUtpZjHlmq+1SQMsi00y7W+T1VuXeAd2jqTkYFpSkCRcFkZ2kSahft8aUKx5+Z3FVOI
zsan8uIsk1EllqIXu8q6tMaw8RixvrKy4NDv/KlOZY5fMDwpQlFND4/EHyobYIplYGsDffc/i27T
ypgdD8V+NjoslKdXt8wBGqJy89Yn/8cCQJverUjQKGiNjkNU1iuOg2WSa6u2+hFabGUqlfyjoH9n
PXNoDC04GqDtGjcr6wKWkGy06K9MZcIvl9rJjifJiihCdQFLgFteb8OJVvRXKOIFu49l7u6JcF9/
KzFLFWEXSaBfX2OXuUf9AEDgo7lgRVm0Go9XO2v3bAE2qnIMnNVzqgdSRyI81Af/8JgPTzTC3hgN
pDBmb2vQg6elg0Dgv94MjGeanx8vJgS/+P+jS53m36X4gP+Si5kA2HPGHGyR14DqFzGhBRpxMdYh
O9ANdh4L1+aS73Dd9416UM6nH0VedbUnpsMjnGM5Oe5KnVX1FPqFs7u1T/EHJr/ALstxtcnkA6Ut
+GtjvscmWX1czHsz9uMJ6h9/ST7Ek7t8lICo0j+gTd53kLypblojnLJkpfXwYZwxnWg6lLyrKOV7
vPUIEHQ84vG1jRnTPnCXiP01yhnw0qKo7acHVE4UyUdt6PWImpMma1WDFZqZXWG1//ECRqaI4BjT
Atqq3H1MdKYNS2acb3uJ6ohBWvaDD7KD4xcRIxR4bCx+wo5FIJp7T05zim019yY/GVsVI/9LvAdw
MBaoccobaRwqfUi0B7/gyK8eSuhdV/1Wpe7KMzOwsYY/jD1do4a05Ozr54i10IMwLDTscQxU8wj/
23oX9lxlAxAaDDtf1OQ6lHOSsNtYVygEtKpf/Q27/4sxBMMaOQEJ61xknFFcp9ie2BnQUU8iwFXV
ZAncLDLq1sc9A9a0tFXCZ6ZL1xs/5Gwk+VS0H29G4nPpnRLf5Z6/jN7efd91gtbU8whLWVKxUCnX
OmL85/1qwlD4AWIeQJmY0M3Ll42t8RYkwL/Q2ldQ/BiAK8E/6Lrkg7ihKtbHs62e2hUTOig9EhFU
gY8Hk00chHZTp30k1AIrJ3rpQWBjXiw8AaRuaBWnvSYrSVa4H82aofuo23yPYYGRtcguPJzCDKU2
OlMsudW7Bhv8xIzgWHnlv4AxRaX3ceBID5gvjZ3RlqpqeM7BAKgQ72h9kJQY/iHeUqYVaZ1vkp+5
GAs7KUGU9OzHQz54FjNB+2wYoxqESvOoO+/+WsWObDgHDtt1vqwxzSxXnXvaNaWBmQ/zILpbCy2v
Fi03Hgm9tJxCzV3PSWVAfHlp+SahVCOUTwE3cFW1XKCBKaoMbwCAGvv4d81yhBqzWQCN5lgjv28q
7pnYcOVWhJIW7YWDjTKnDVcoDgwMn8GhB7NpWFVxYBITsFYQnVMQqkJyDQseB4yJzp8LM3m5S4KA
Lu415cIYrcHlFB09Ev+jSLS1ydbk3tlbPo+czOF82DDhbWlEF9cxGAWnUxuFCsk57Hmis9a67cDn
bNpZNHsciBNsQPQfeaVI41wu+AeIP7qNIs+DIV1xd1Yql9SChs8V26mblsnV9W6P+6lGRY/bMl1N
NOtgIvEvmCsIccmueUga8toR9/plLc9jXoiLdR+QdnJ9PanC/ecymGK4814bbe0UozV0dPVA0S0f
GQr3ncJZfqtkbuDcrdk8wu9uKT5R8y2XfH3EVBMuxDw7E32FRlf+vgHyufAmamA+qmePWoL2msAf
+VdHtf8vxYpd8N9tSMzzf85ntegngEwGQQpceQwqmnMm6VdAh1dw5KG7HTfbw5gjv782HSkA/jrz
nbi66AV36u4brfoaqujQPsG4lf+V3pdH1zYOgf/2fG0jdv8HVu0dsXjJKWpdarZnrESFn4TcoXJZ
nDUqAf/1skDNHmTXujcsp7/eBmT8T9n0eNdSxDIEMv+NNRU6TCxd4eZS94AwhYJJ4w462mUS+xDo
2DAVekqRIiNhEw5mEAZxPuLbU1ZkGbhu//u+1HpAHc2CToxl7O+0DSoap4AD9kgh2Rlxls4n5as/
qB2gyS9f6bZSqRSLDHZRzX1j9laES1tX2mRGIK5hGDewq7e61e9w5Sk6Qexdf1aKZ2iRWQ5YNkAp
oQ5CL7bH9YQ+nBfHhKVSCa5Ha6nZ8K/j5qjHfPIOXGszxjiOtxZmgLMVr0PYxZTUenf0XVCMZyfJ
QT7ArrmrT51PVV6V7ws/b+4YBdQbt4dnJM0/394aFyHPiT7Nye1tb9cQOiyiCdR2/cNwTJ6LGMXR
jdEydhgweGllzeMiadNjVIa9YOFjCsYt+VrPu0/CMfccTi8Booli1/1Q/XMyV4ZN1pHdNb9D2vtx
O57FZIUzNQPYPOdA+WqyNY3WYcLQrN7AfC1gqoK0Dfr8xEYNIyzjmwqdu7hYirZ0ZTxFttdbgNs8
CPGcHDTIFou9ct4IToi/FIEwF7KVjI52zCW9buJ2bNmBHLK+qcHoF99UEpPUlhMfuLQPIXyXetwT
YJP9CIKaJsZMtjETshSo1bVSFLJUGp2oNK3DTkgYniHXDPTMDVaZBOYZ5X04jt4q7pixlSvp3bYb
0lVIx1PEcPah8RZszg+V323HdAhgr/coWo1gnys8f68xB0JID0m6QRtnguDZnX29SnqGWIpHXrUp
bHvKhnrGYMQoW3PVnDT8qELC6XO6de8mZQU1JcEaU9IUBrmrKVQVBZu+gUsIyJVY/oXbWPtUareO
hE1KX7ctNqJAisnHSXTkSt7ME3K/fJFYXEcI9UyPJVFFn2Dzz4CGbUxO0QJdXu+cCe6V+w49CFfk
wLYCmgjIHpPdEJjSpbX9qiYIp0mQmqjgwgPC8r2yvvyreVB3pr+0m4sW/DIyMFbfKFngEU2bGXqY
8SkMtB//RRPbd+Vv4Q9Khnsn42SQLDGWj3i9cqoyoF2AypTsXEu+wT1TBGTM7vTA/MCHaUi+9hC4
CEInQHOo+kmpDg03amYQdmL7/g9EZZ+gM1RjpDBQCUQcjws4Fu51s40j8MXuJCjiP2EJJPzuUcCj
Bf+KHsSTMCi/q2KX2o/iPAsWdOG0Lla8U6gN5Za5FKmxJal9vNzFTr78T/Cd2FQLXedKPUpl2sFw
3OvNitfUuiONKIoighO8gJgVqKoEs2Ex4ojw3QKgvTQiaHJe5Mv6TBgX+Zst9dTrZtpPtQb5saf1
8hHNRMC3G5SDArfP9CcrXtfbwdMxivUmXBm3IHtzW2OC8WZpdxt0/d3cKo8EcliEIHZt3oHAqx8r
tsz8MQT+W7nOYv3VsT5mlYHEX+1OaS4X3vl+j9rGcpDU+uaFJAghv+qMeauYFDVQYOMRNWc3k25X
EfUN3dt9iMDYEkTpUNFQO0XxefoUkQvCXofmC4HmUzn9A7qX+dc9idojPicgdqAtLEsVpWRXxu8b
SmNWZOV37sP9eGU4lWm2OU1Id6MtFTn6QMiXyn7FBbOgfC3dtU/3ysYY7NqyuC5ZVJQmQbcU+tek
8DZyA/Ofk2amfwrrHZaqK1F/Vl6Z2HDsNEyoRJJecxC4wwRkLUb9uYdRRI6QsK0Vj47MiQXFpccY
6LKIfDko3SQ1VFD0/OK/4R2h0qI48J9/QhhYw5Y0D2zb/G4Kgv7XuAH71k+/CKBM0KGTFVm8Sa/2
1GAdJFldG4G3/9TCCfdrQPh5PnjJxK/LwKP3TEAdo36jSAHq34JjVNj1dAAJJHHanH0KLZip91gv
V/rCQsQoGjS4J/7LlzBa3Y91hKfmIyIGkqalOB6rQo3fC2e8/DQHZW8GjSxyGkwgK8mvfMTP8EZT
IaqY/NnJT3awhHgFRq+X6MTVgC9rQpYW1/VHYZvg2Ntn1S35FT5jWcJ4xHYMoumFIotNZPOIc0Qg
jbecX6stYGMGyNyERmDyUEfPzBdcik5/AVUkEjn2HsB6PprmsYxJboXmE0EZvo/HhebcBQnuF0vD
iq8bDium3d2caCnqm3Km9Ij0aRC+thYaXEIlMxTSB1B1TCLMTPY0ptz57WsS9OTHukeZdUwjq0M4
J/5iNimsfOBIy/bD5rIrNuzh2Yb0DFaLwxYKFwTceBfpruQF2o/J0zh/9H2drHzqDEoduc1Psuw2
5ZwWteWHE6yxbZSszUPNkkPoVFcJ3WojcTxR96jJm035gw3R6QtzVPpJD8nIciTuBdUVWmKdLtX8
CtLCCivvGUChsbEFTusr78gIWo89FvbB9f+/6eHmMb2vlVeAOPtzdxiakyG4BnH/gUbEEs4vp/8k
puugfTVfTX9768L/64cFOR5rOObN8Kk7LQQPyZrnfarovPvotN+Tadb6OrPYmU5CdXfg1JRiU6EQ
FsWjpcmiq2sk8yVQ6uDBR07gs/KJZoCfcjjo0GzQIHc9P1sU22SNQiVeNP5PBG0JuCAsSUcSY9KG
98otAs5KCRvoxIowL0SI6ExI11tc0dlNkgLRbx35S6U2JCiXapRBFmnUJSBGmyuwtmUBYX+r9dS0
1OXvR/pD/eYwphx/AGpm2BhUU6qNa6bqD2JoMyo45y93jbQIokpSRMdlH3VAOEhCnjM4FtvlwY2p
o/mWKoq7C3myq3grwVTRIe44UBqyuqoKKKUBS4eoC2cHivoMbG1vI4Bna+ZIABRIitbaovpAsgdm
mzcUZqzYKSDxeGEd08FZY3bE9ZgOLzsCg9hzcUNp4/AtWEPD4HCHXKKTP1t6+0ltZluT9sN9apkU
OhA+kbquROTlVBeHSjbffhpvXvlqSad+QacA+HxGwXuIxV/1xsvWDaIjgRwxeua9rTDOl1TvPdk5
0rQlnypMUod33+5HoiI22H++eOLhlV2dnlKQNobvAHeKkGwVE8+/RnTBBiTaNag++B/hZGcj2UIP
4VEEUotJV+KcuybC2+vAJzMQF0m9cczVBCZVAwsDgjtwEkLU1klXd7mg9OcKtKg7twNlXnIi9God
BRrTCVedaR2KwP4UFMH/tX+LwulN10nv7jel+vdSuXXo1aHHqzYQVhLS6S6LnMbGLyETFvXjsDsx
UIb7qXCv0v6TbRp0Ptgsmudtk34vLiFRsp5kbn50HvnDpz94kdZVi7Z+wdxYkf1ewt+aIRnN+ehW
potN3bI991C+C1W2GoycHS5ayLApcjmzarOUqgN2Pg9D5vRjtGORyt9GE7y1tyX41he1ptxKcGQM
f+RjpdnVr4FUWBv+Y4ChDye4xoNGBi9E0TryLTsNstzHeYYtv1e5+7xe1rvOnANFLAVyKh8fvqwr
Z4r/k9O2uXRIoDZqSRtrZAvRa6pq/1+V3sUsjZrQodELwjL097H01kCblXS1eTIz3Nazi6g9UJRM
03xiKKK1Us6eqiDY6Zdvv8LEC3nn17CYclZVF7yJ2DYuXLtXGXgHHucSISIcd4x3hxHwlekmTOIO
NAyHkuEYSlsZHN+VFOtBPbTLacVJ5w3Znx2BDNtVbZJhSSnu1Cv9LEXmdtFcUh6ai6tu2quE6qcC
vb1qCnuDOQLvTZA0ph5WdiPdC+Fup//DcW4jg8Qm5v7Yfm4JIE4Ggm9hrXhWoaswveIbHw+q5zf5
H7eyh0aKuxy//32lXkbDQAgrk9TN+22d/c/iHBzHFzsrLTAct3URcEpLyiXQqAXl+Q8CeoVSuR84
Y0fBpNT9ZUiAhio05PDU+o2Sbbt/EVhsD6ayKRlFUe2zjubP2LUm6EBa565Ro/9KPJyawOD1uJDn
Yy9d/7i5zYPsIqy9blApnYdJexAP2EUfLGC2qI2p98yLna424PXiU1RBOqhmZGFaE84X7r81M+Vf
fRa7+facTO0RuxfyGneaEvqLJvEg9+OOD5WJeHMAEjfNTeD1CwgCDYXK6sJs4HMDZK+NXo6v+Zif
PgKJ1u9oFSp4IIkL7JQIc2VMkR8iJDu9JGN+REQU8/GXBDt/QSUAHQMCZ77l4nRALG0nXtp2cvZm
vEvmsghMv4EGVC16x4LoDjiV33rGGvVW242ES5ADFjLoYvhtcmWjsFVe6sPSad5zT29BdccgBP1x
OIm52CSnn1kDyeCCbuyVIUHh/K4M8uK4Y5wabnTvqiyC2GZ91gtFbdmVby7niaZ0jBk6L4TL/d+9
O3lO3FciSuzm8KCdgVS8LFeGHcxwlUyBdW+nl9KDXIv80i580FT0bdjx3HApJ431sdv5O62w1UXX
xwP3xe7Q3+NuVwvNQH586KHtZvOG7rsWHLnYBvcv4N4kEsWTfClQdEJ2wVJfjkFcYZvI46I2U9fR
YMUcpk5CJ5+lSCvZ9RGrSTiQ/fDdKCNB1/1MxYagAFD2nlgCKwnKm/HC9V2YisgpSUIq8mE/8Ye/
UpFZ1dRfGtQkxS/YK574Bpjoa0KjWTiUjWxgvczw2kqrzo/H0gNQh9vT4EXvdFaxOV6nu6moWwus
MvsuRcIWr4JNdv9qdhYBI1KgDxXG6g2f2qh/7FskeOlCxOck0QSccKRWNS29jzvy6JnsttBrew8O
bVSf8bKWRLw/H410xFXlMEcte5iB7Kc+ThYXaUiUR1s6iamiAR6q85av/DlCuJiHW/X0HR0OCdac
u1QZ1t0ASjuxyq+CDZES61Oe2JjfGtcxBixb9LFTLbiRR65R+iHonGJcIfZOplyBA51cd/3XiNy8
VjkOJ3jO6OMbOmXzHzNHA8aRpxiAU7PSBUxdyawuilfE8FYDaku+vCeOSH603WsatZIqiQpMqKf1
YwUezd/4DZwt6cGZ4oDzuMOVMMDsX4GN+B+AHUNixEJZi0GYEByW1HSXOD07YitPTfkfjW4zN69i
c9Sl+v11Fxce4C+fjAx7QuK2QG/xC1MZ/VSb70F7SG7XROWdgNa4qIAvxm99ORqds4XgnVedbOlL
d7s6aWKTyeojMT9D3nxsxdtecO8wIjgqMo17riasaimyUcUMaJkI7d4rBkQJt+hrYxBs8xJoIcv6
hsXFIvNwzZzYfJpoiMY/3Bj19PhgHOrJdPmHYGFVK5LxBjS68Ep7KY2Sxp7VtPxGqasFu4sWnk3k
m8JOZvTzhrgoGrtsgLA+nU9m7iAAkbE93iNYCDGK4+jUimm/WvYyqSZkwqCmBE2brc/fE9mHa4tl
l4J57wtOmId+HWy3RRAEDhX6udeiapYApZn6HDJ1HHyxSRsbSXAWDxLZ0vBXSpD2oTV0hx3ymTEB
D5J7e6CqL5WGKJ8iTLOxy4sGgrE3iZ7ziSjmlwFXd0tlrM8ycKNCM9Ams4IDwRtb5i+3KBgZ+4k6
mfwgf30VFwfgxZhNH2cwvwnGy8c2HtuOJbGGvJkSxv2GiZM1eo8o2Qd1Wp9vejL7dVnUIx/wuqDP
OQQ3Bacz9cEr3O4ABrvCfN9MJa7ogbrerRN4Wi3z4p6wcQMKNTEVfxuekcLwAX87sgnZwU+yM9N/
6btj66/UUJqDPGna9LmBh6P7TJ1WmtORo6nAv9B1tpENxK6w4zrDPtZ4LdU0ek33StjoInrOAZ3G
Ez3fzOT9sY19Ol7RGg2TurKqE3NiMRY+0sFzvAS6ahdkCpUHloVO0Ct/m8xyHQzmAhhKGx0KAII0
2aP3hcG+LioXZZvJM9/tBTWnw71vCvakZZ3UZsuyrELwgyV8aur3esQJgoCwb2q/+vcfrbF3/h14
pL3h8lBfS7D97bAhbu1SGJfhv7csOKveax4ciBkWTByykYogUatXkxVh/FLl0ShC7aI55OYeTumM
cfB5k5kplA1Do2/9A1N7VVEISrKYxhHCRxhzPmXnFJyGnLFeGBuNOIJhNS1MCcWtTvrLwsjuLULX
MXHW60bLQAar7/YYUJC4fipT0E18yJBlIiapOCj33QGcNmr4BAgNlNBGVng8wqOpY6Vd4VLREAoH
YNdlJtm613Heo413j40LNIFk4DSINtxtrxLGOMrBJFUlXtEOXtBi2kZTq7Zl3VmZyymF88qPHm58
AeaLbCinaevAgbnwR7Us68o5MKFRQuYKRzpANTl7ctEzcJqYPLp7ZPEuU3npbE3aS0vkJzGVpc4V
3H/nJ70YTTAmwXoOvdExmxhNjIQwb+nH7jYQbq/AltJDgRBuaRap3eJNLkhXVmxIp9Cu1XiBkqHb
Uw4eQYgk8Z965prk42cSlQ15Xq7z2HuOOJe31HGnxAyTvt8qxjiziXah/Xn8NICLm7puAsRKLwk8
mUxCZTk6OgHxopMfe68mFdm7Emph90l/9N/ws2g/betZUfJjarU9bJo8QZeNGmQOAU07s/KHWhy8
cs8Le0lgzg8kd2+P4WKNrPmIx/Ow1qQeSnA9QlheAP7mfYEYnck+DaGSyT0BYVb2jSbdoJo344i/
UAnszA5HppvSovEBzLnnGWeWWObYXk03BHLV2jIsblMEv9NHcrVwvaUE0K7FL5KZ6iIsQAb7+vUo
0LdUuX65qPssKnjC2hzHnbLyrn65F8FJtJCHpGXWS3e3TZVdlTFcgi4RnWqNPd6LDWZBMictQ8ZD
Bge5Tdo7B1PQM5VTFSyku2PtWc8mwdp/CBo1IwTE+T0TQJfGqnwPsOOPMVw34GW7YDXeKpSjSfXs
C+tmY/g6M5HKO8yxF48ejAWeSwb186YBr7PNDBYKY9rwJDWdYxckH/CP1/NQZH5xUMG0YdyNJHle
bN/1YXNMndII97fnQmUKS+Z/dVD3wLHKomUgKKnFT9zq/5zndwAwLXQF581J0J1S1PfxdpdWJCwg
kvxiZTly6x8KH7v7UtG0e5Ymp2YxMFoy+OlmsxuQ/Z3aWOECHcBpXKh4Ct7i4e/TJ4RwUHl7012q
a7SPrZW13ZajpvmLXz9bJcSRzaTb0yWgtPM7xT4oqimehciYPEHULcWOouuu3c4ysfqUvAoHZTug
3xeA/Az4OxmZ6p/t6bZ16bkuVcFpdE/AQ+h39PNrKgf4WechSjcEY7rAabF4uLFetc0D4DFNpgA6
p3xOPZIDwgmJjTKxMU3RHZKNFlf7Nn6ohjSQ9VKSiS/QY7MLDqg7fvCnSw0f5L5ED2wcZq0AlKwy
0VV+buvvlTXEaHs+k45PfF8w2waDyxfBlfxv/pd6+8RqiEb+B56P5T6nqpHHNRcRHFbfd1uQvNlm
yftRumgULQuriayJmpZJejs4tB1qwu878lJMHBvR5oxWJohwCil38QQREcHll9fL4GK3wR3qNCHv
hrc/y0SYtuF5bbJf8y98Cc2tDKqCtatuPEXOzASUTXCKuwcY2+S1xxqi7VSz6zRxkBZ3yA5Bz7Bg
XvKa52k9PfPwxiLXYkn4Fg1BoF8rEu9HQhfz1V/Q4UXFNmBqqczYl7ugle5PEdSBKEv38DSw8IGK
8baGKOTYVisL42MPgrLXOKtYBMguX2i+eHMkTZV8yQ1PdGzK4MSzXmJ1S/jAw4/l3oFs3E+7XeRg
2Xadg78CQNOzj6h72x/ZcbHAbEWnOs5e5DLm6LY7C3V2MzHAG+0nJTom5M93BlXWvtung4KvnjOn
LYkTFAGQepzBEdjvO4D7nHL2NT+CNry/kyLXH1ZUnHkn88/zgYCMfFjZMqEjzgcNSx4AJKxYIfIy
gnKcbyHz7a0ra0vksGd5F2RM0JJc4/P5eUfG6zA3afv3+BbMqBPFUan3Qks8caqSFTsbnGMkTRf4
DSPS3pgWy7R3agi3IxmgerAPGfN1/4npZur4NbMgfmCNZBFvTkpiQTzIP0Iidb55CpOAq5beyVJd
+DJ4FfgA0eSwoMyAjb+xDOF0R0w8mA1lY90sF0DeYYSORtI8t06R4mlm3Cg4LWa81OoeJTiDQbie
GvZf2MHVsDG3Uo4s49rCxz84W0P8suLHSuiR93cYb3a0l4nKd/OZELMiMW/jLt+7Rlg12v9+WCI1
ft4JiOYSFt4duGjlIOLb01N6TrViW5QnKKwlt/LIAjAghGSubx4FvQTDVK6SdHNcRpvFGIB6WiAl
1yUjuzlGlkHbQ2v19BnkEO0jRqmQtZsYVmLs4jdx9CZybF8pZ980hHnwbMtIe41d6DzWTNyZEfDx
d5EIhy+SGRPuit75wDiipHRXv7P7DY7bn06JPG25Yj8uJu7SEIFOTbqU+S3A58LrwtMUF334GZcc
+HO87H+vWkrvSB3I7U4w6SkYUHgzLaVWXqOPq2LniyL07o4d2JxARswzkbG460o0Ktf3mjFeaZON
FODGv2gFrwZZr0Jenm5Whv7cK0n68JQB0uoetJZKi7qNP6Af1Am/H9Q3EGJD96bL6l5qptEUfo+e
dU52dYMfdpgrR3J2Bptt7XIruS3NvnevXSy8jVe9RtDH1Olgg0ui87hO6uIxLufMduVQ4AVEddpv
tdCIugJv/OiKRJoZTbBCAUQMsos3b+IxBg6hH7hEZYPBTzDygYITW13KAbkCv/q/uBUDUndXpaWQ
gOH0aEGrwq16hA56eCUhenuDxRW1Pon1g1A8Xaoz9H38vEuZoJ4mbEwPds8n8hRC2dYlJMlqaPfX
9gf66xhMMmaS98DEjFtzHnfpj+CIwi0Stw8rW3XZM/LQ3uQH6A9bKYas4NlNEJCD0BB5lDCgl3AO
tqhvZ+9ObG+1qB5eeM1YR29QpTh8AfUa45QIBOm3WRUwCG5WQZbOZI4nMULOUaOv9o9I+knPsaVq
+0oKDbjhoR36yBe2sdpw2/qEsaEymNJwbbnAIkCJxwxMp/b1t0JoI2pePVZaYJCrWTbGxuLcBQ0S
22Yg84SOKye6OpDQQWCvy0a2Gmww+xYczqsl+YvJa2daxMZaaaWGSun/khtWYItUe3FXusTTSoQ1
CyVkUStc6iLSYddlhTR/1NKfIiEGFLNKs9ZcL7vYYXFQ0OyGVvDoDuisI6L3cmRPDX00r1QIVDVM
W3hMXukDpD1L9ZnraBTC36fjuyx/P5wNq+JoUdZ7bG4zq7Qmk/V2uyCc1oJHjdWtLfk8kAHMY0PU
HiYs+H4VT49tMZEUV/Bwb/mWIW1D+idiWEsBNtcFsET70g9L+HKpxY5WCib8jEq9yYjNA1yNfZ2A
91ZzRWuDz/wSfT9bQNXi777OrWFJ+CjVxnib5ut3tN/P8caIAQ/0IrKtwzDIvyY3mq1fosjtuIPI
bhxGUTevwDHKShVyxGyh7HGG5pK42zm/2s+WpN9uZYfgMfnHrBrywQOuJose0hIdYsTPRw5wwgNI
EGytWLYoJEQuQS8PJQNQzU+i96rwgC+WHfHDzPZeQAtA7qkg8Bb7Irsx845l5d0JyC5PS6Wu+FXo
2I1udUAlMsYMvII/kAo0NIm5U9pTSuy3Yre8O7O7FjwaeH5a9kBLYOne/YChuOaMdmYCawC18kDo
ltKVYXaHE1xpODx/vwJmxNlQSVHX8y5RhwmIl0lPn2lVeKQI1OlnEpPFbujsnXQ0f4FwdeyT0PVW
mUIwJKmthfhXZXPl83BnSUTFuDnyP5bE9szgARUIts00Ov7AKcuA42BNdO8i7HbV81SR481z1IgJ
vuOl5izY7pZuoMB1xdJXI/KhimlChHyxZ4MWSvWDxkzcW3U51ih3E2A6+5QjqAAyfBRzVv+6ebEA
fn39hmt4VRG0fNKh+vDMRa3YhOnOkrEXGZ6GDBeigtHfGlhOX6qcZUzDHqJLT0lZ0woaUzArEVR7
Wj5ZegmQ1hcIUGjpccVAIEBqk2IExog5x9k45rs9Mci6eErJ+IZes8I5mVhEepcJNT1PIo313AFD
/izB8mj6U+y4v0zU+RcmFJsAXYro7PRKLpBcaMiDrJsUuaZnpQJA61yH8R9OJCCkQauLKXE/atKv
gEwcoHaNzphW1hvJHikBpLXgD4yWzwUdQhI1lqlwTIkXq/Qx5qpeds5xlMI0wKIO0K8CzhB6dnE8
rVJ9abtHrXtj3TPxISSSHqWGlyW3dA5Dr9x/UdxlU/nc+7tUBBnOcN2amvlfytRdjfidC3G9rVZg
1lKYVZc3DHOC4L7PZzHXq6tusrPUF+1Q7ddo+nMz32RlbZedjvN9WmPHnt2FhMqCxq3zXct0uKfR
BSTUKFkfB9R7WijbgNyORsUTNfoiKfNQOCrffvR3kDsf8CqNzmEOhE43zzZhGDIBacLMVxQezYIE
5A2ThO+Frg4sSJ8L/nHsqUuppJtKnqVSHr27TUP5g4HN8eBsSwSYtPcH3OikZ4VGHzkfIkA0tfS7
pm0+Cnt6T95kFGMKeYCps7H4m9zAbHFwaQv7hBu6PrKSbA8KwgkS1CbPQa1cS+2YRrzV1NXFnh6W
PNyFeP1+jiOGC6koZ26N7HzqCqZAXNivay0IaeQ7/YUbGmy8FqtsVrCq7GUzejngLJEpoqM03P6s
GxQ+qZI6xZTHrr84vJ8KMFRBb3K/Cm5sVu7pxNirvoi3t/c6a773LO/cmjwOOTqlzzQqkB1b8JwS
H0MwIOrf9TwBzaEUB636pNd7r5+0Bf1YcCevFWTB3yXRVIyNQqKaSUNtdUgi0PKkkeXap6SeZd/P
oEH82FW7gR+CohnKwovfrQuGXe1STvRrCt1149vH4CPvPIB+7sdChxR6vK/0dJjoqNGrE7mWqErL
u00U3dQmQFLvk8E0qSk/3V1rv/3lRP1A4+sgPz0CBsb0aqoQWX8u/MDR1s+59mw5g9E1AT59uYfT
xfcw2qUp+jWcfkCrmkJCIJGngBpnLzUiCI2G7SDs8cyJuV7WIHbSsLyQexGNLax1Cn2IfkyxIS+3
3RdXG6w00xQp/nNdKMW9ry72YW5BFKynhGjkIE+bgjKjSZ/lZh+0L5zGt32WJLr6m8E98bKm5CNv
ajFNIIvOTU3oTf9nb+YUkb5zrj4tBfCwR8qYmYKiAdHg/gzXtpQ9lzLYLzuDBd2+1lUzRE2mInzg
h4SMMyzGkWKjQp98jcp/8pG2VI/TJheSPSwXb5Ws0WEhQJf3Lv1G6hAkPs+GGw+YzaIy9euGXmMo
JkSxsZgwuidsG/zQxfOeRdbRWweaUrrtu9QjkAYBvly3hutucrjjJONREn8G4Bob7iH02QFaqK+s
XthYEIubhSUAxp/Z/W7hozA8zXbnT7lWU0XYM9VDRCTrE/azZ5w3v1RDqrshbofB4oWuuMA3OIMQ
Md98LBGFy2eenMVmGDyc0jq16kejhB4ePw//Bu0tC9nXb2BS+yEBhPa9H2zKfJ2t8KnFXb5e3Q0W
qTVCEXN6WgoA/tZcjdsSyQFKR3ITbyrgc4oNtEIYpwcmiZDgNprZZoMAJ+mFtTWfOMZgjcAJeuPW
ktHfbtHImutdLFTb3MaxyBKuvFo10Q9eoZMtw1BlPMZ+NXF+CLoXtVbvQ58c4xiQc9+mczqrMNdk
1DYaEQxY/gITfMl9+SOW2tqLIENKCoHISfcvGwaOCIM8esguAwBzcZt8bjvSrG+JKjxewGZfGuVd
3psBN3hHAkaGtF+ZdFs2dZLNn4cRxOq+cG+gROWxBSaDOONqgnMCEbbCjAZuAVLRtSHRmswC6eQ1
jKZHJIP6p0n12DCRZopSWUCIRgHza6SuJHRE04I22NsMpbtjko1adrK8myINVYQCntSdy8/1L5Ov
pXQt2KGNllTPi1QDeQ+IIivy2Ig37UrTzWLCc5Wxr06BteekFmdjXZPVerPLWa3VNtu+F6WfJfh7
fEbhcbC2dSHEXgTRsxgwLMr4CSfFtMUBYBS1RgCJHjo1wuCSflj6qlBsWOeUOf1qAw5/qgfx+N8I
bdi3enC0CUJbudP5zTpLYF3PYH2qZkFspzr/iaz23xHD+NYM5qF+n++E4a1wV756wJA0szMXLtq+
RxOFSRiRMos+Ygs2qr+xh4fNI7iBNaNF/7VO61FcK+CYHAi9/RzHFft1WasxL0/6xhte6YtHQ79I
OdS4AfyeQFtPtdCfaxKpVAyFZglFulcBeLDnJu+K7LZ53RhBCxsno+8xuSNLOjycC2sFa/aMffNV
HfXxK4dDX/1xxQQEcnWQjxEsubI+hy2zyR5atgHkT8te5JJPzGtHuXHapPPiXpFsEnnb0kg75Y0P
0clQZYwUhjb/ZaEvcK1aCtQbe5r2JuubFQEwE8Wy4DQEM6VAQ77PeT1Z1rnjEFofRJHQSTV4rby7
Ki2Sg/4Ri72txPT+ht8jXT8/zysr+l6ZXOV9GSY94DXEvxT0R32ShibTBCKuKSZkT70y9mRvvrar
RAq9gITdRY8Cv4yzkthAKhDSucImFmyHiMrPYP1HItiolROUbvXpYOp7Sibbko3+TJmj3jdOSGZ3
hSYaJbUL42QTIi8qPoQkKGcu405CgMkuPpaIMc3/FgV34ZkjcNNF5tb6JVbtTQ6+BVcfCx1YzCX5
pXcAy5uy6Hgv1qixGMJCsiay4nzP32VMaLBVhjKvvXecKtf8VFjGA9KbsTPEesqt9in8qIRxU49o
P8CrQN+DyAMtuh6/8+xVfojXiOELuV6mIYxJ8oUTO/bM17bxABsiUgfXVVwXWCnUJUsLd3+SSW/d
0rI+edRgOhPHvs4FqhHzG+ltadWT90EQHUjw2y9S6lHz5wOBzDzXrvB625Zq6xPmsWOd2hRTTuh8
CBXlBJgmAuKwxxx41QrRD/ovB/dql/O5nH/Sge0Q/lz5bqeyrHVgmdvw6I1MDsL1nRU7oL/CNHne
uw4FZkNIblgI6Hq+eSJKzWUU/DzIX/FB9+leLn5z4VANtP2v8kw693aQbv66UDOlDVXkSuQZAq0O
qPpR//X1DdKt+3syUZtj+Dd3Z5/cmgKh/BSb7d4K0dWKVSF+DEkFHZRXpr3eOPtMS7d7a/fSd7Hm
+ElARaGXFck5Hy1RIWvGLpFAC0XkogLg/h+P4lJFKWHwJ8V0PKAUdmJwDDj2lQzjtpgaLp4EJjqk
chSJwF/4JAu3yL0SBpdCZdJvpaeDkM/HLuD+jI5Udc5RzG1P0wt3jgAVSsECbCqBk58wThWLz/xe
ANGkRWGShJc9mM90a8s8j6BtzxxtVwCSiN2sMW0lMtSn6Hd7z8ipn0oFnHmiuwUVdj4QbAmob/Nv
achRzUGIj85zO1GocO8JeTvJNSLQQ13Pjg3+sAEJF4tuxEV2gw2bczrWl/sKKab7qyXanSMx4Omf
Z4b+duvqD6rI82YlYf0wajnrtQ8QQAQ60f6uE2aZOnL83oOpNHzoTq1FOPcSxooXz3koLcJj9X3r
OUaAwOtMwxTZOxY+G62IBkk4VF1wrNLmrNAyhmkgu8NUOsYnfWeKpLpueFSQX99WQgF5iiPnFZmO
8pKg54qGXwFoP/zbXIhGgNhMTziVYOEuu431B8QtF0tyZy99r1XXUe7lULKhu1WJ6HldfihUnzcz
G3XsuQq+FWt5eQ3/NVSkcfcU0SJrbYKs564/UYvdgsELhJLu/gMtDL4/sckwm3W0gAkcu2ZK+dVO
h6OCcbwGnXfXyZLm1SPWG84a6JfgLY8eQig6Hjv24+U0Esq7el18PA44qeOK9dIturGMT3MAK1rS
oIRPkTXpsojXo3jXCUeNp9uogDrmpqCjvfO9sSynIEQ8y52tXHTR6gnpiZ9aj2to+ODB7VvfODsm
VcAVaXJKjBxRv2Kl7y7BuESu8TBAXQQOQNIEioIAgQiBGtj317dLKein82TRE6dxLFQ/1xVNprsD
bPHQDHhpXZsRMH+y6URsTSrhLkU3/3cYwVATZh892JBYyNkAeF55T2/o93gPeElnjSnM14qnCeLM
ClY1nZjV2oPGxVvnAMcT7OLDV1F2NIJmlbiBRVQ4+43FdXXCSRkO/Ykk/G1jrX1AAOxjSr/tEZag
ErN7SXq66x24izVCJqw6cqIt2igk4gzagiGEtagb5XcUe59O5MDiCq4z2IcsMtuwy68EFgtHx4vG
kE8C9RLawpraaix7e1nfnK+BcjqwYJNK0d78BN2SxjgEcB4bWyVE5J9drutSZzscysGZZhwIkdia
VNWV7Ra6bciLjN6bgHyFfAA/8EtfcMPdKrQHF5DgAyXOtHpZeXRN1dfR6vBsV2qbx19tyAzBFTrN
NGa3WInYFjYvRmJ1pyKd0M+V/7MQLi/xySEvw/E6XtNyqmHyuoxG2q+/XwCfTApaIcLOCKUngAXt
rEm6U0OfcBZHg64gK9lKskdKNlIZJAQYLV+muFIWS/MxyRzEa1YTIGMiHeoq3t0pdKp1Ms2nNX09
UXxoRzChy2/MzH6aNyp2OmweZUpLfIaAoqvlDOF7Xoc9qdyN2QJpLAIkAbFhV9Rg1LFdgKNB78bu
kDZysIVWHnXj4m4xbsnWVsTSWWhULNkAU2qGucVpPjPy0IHxi+9o8hAdboe5JhYwcGkGuzUgJx9D
JPWDt8cbGjBUYcSHW1j7OGnyaE9EwkgFNfE0NmYfrkM48PYghjpSVp/FcXZ6rcyFko0uP9K8rPDQ
pTp3LOIlE4DCETzUe8+i4nEuIpoPHR7RhuNGxuqitdTSG+s9pWmuJZkg27+bAaO/ewlS9Ec6yn0u
b0XpgPwl83BDQuBRItNIEC8fFPYQ9GrGIc7z9rrNTeOudCyC/ELJKDzNTqNjNi2MZDbxpGGw0QOt
JlW49ciaeW6dADkyzEn1okvRDVjCyLWAf5NLlWObm/sodvN7yXfmTIQMSKr15APKf+WPWoTJLJry
fjo8v//nEVvBC72E2lRQNkcRQJt6FnIa6AkVwnTuhjKkqPEmV7cciK2Mo9/Wy2TAwEgCIaFaYjz9
zJIkGryhszuqAtFQp7qvJg6bhCZm+am+SOQlmJ+OjrUgqpjTpkQpOUq5gxq88ip+Pe9MNmzyGdSq
4SbEaH07YCNSN6pwZ9A9V7V0cEc7K6JV8xkBnSTMUXfQZAA+JkbeXFcZ/oiUy+pd/unz1hZDJ+Ei
XJfIduv/qam0OtpfKxkhswY/dK5VLBISHjHfMOWjxHvbKqCNuZ6JD1S70nHSjX9RySCCbxx13TRx
dMpOZnRdQsIJ4QDwrogcJcV1QkL80WP9plvV26zNhdU2c3XLbMGdPR1an3iMFQmC9NZ65KPXlaWh
FOa7Gz5SgHV3/ZY7ZY92e93yWwhNxRZoa1wmR2ksZXEoBTJ3sXKlHRKRscCnJtYVIKmSv15YmLLm
hLtDarBWwba/2trmbDPmYl7DQiuzM/ORdkF+TBKWaH//jGDva6ofjzgQT5MSorX2g4qLZqaj/aQ4
/upW3VQylSbuQ1Nut39wpwbowAwFABbw4CyUpgj+gDOGxd/b2tTbb1CuUZQVom2Snp78SPerXRJF
2+JGhuhu/7sNja/2wTp5V7zmAFcRn5u1ZrqIeQqvi7cDvJ3wTW9CTbj/fpcI78aoUZaIsjJhIF4k
HJbgO8TNpOM0VMQ7CD0si//tB+gHqlo5a8wiNSrKwhYcNiK4dkLQnEWjEYJdbiTpUapN/UpLMS/p
9iPt6dXiM1rdJZgRFFXE4SC5mG60CaYqlOZeeeqSaNyocJTwx6Qk6/5ydnf4+HoRQjn7+iQGwRFR
X4k6z8LNovO8IjzMXwFXlWAVGShvJQDE/9FloSZcM/ZsjE2lWqdCvP32TVwZ9jG50kEpqJULG+Zx
lwSHqsunYQWIg+ur6cuDfwK/Wh5Kixq1Lbd5CAL2MAQR8C3UVjowvGnXSCNI8vvMHQ0dNY0RiDe8
Fv4/C40D1rsVbzU0rjtcA+OVCMCNptalGd8PEVCZDhzEnWom581F20+i/aXSWXfXNwe5DE6x4SRL
9KcGiwRflVLoGS4s4q5PUHKXJUt0BExM1O85A3057mGOcao7Zp9Uf//mOtFijnkp2/I3Iq36LtOq
m5/hOCRbjDA49i7WvStkJWpR3X4RnwuX2smq7ZaLojZtkMpNoap8Fb8i3C6PEs4evHX/rfIxcSZ9
6wWFFZhWUwDRKHm02spFf0tbCDL+0eIYoZzciewkJWs38GSwrsj+1KypLV1iWJAHWpNaulqVBZzs
7dpWMgbZFkrmZ2Ii7/hIla486DRN3AT6T/OvVs3Pd6c8V+4/BGG8vuMuOzcBznlDRR4ZNDmmCxvG
kIVPmkZ2e+JjVz0aZFtc8yE3d3XEXA+L1NYrmZ+PQJztaJFJEw6IYtlvHi30RJI1kZ5Hx+g6T+WW
f9cEMJu8KKcSVDOM1ooaNc9efHN0Tb03GYtq3bea+yCY+V2o7/gmby9UZ2e37JPvhhYYaO67zvCy
Riy+tSuJ1rrs0oDiTga2uHuTDOGJ9EGljuxQL1ocdRLR8w70SHhutBxE13zsvBU+yUAjp6pJ+suF
nrCV+alVFWiq0mvHQ+lEcTDLOKox1CpFWAqIDx958visxnhhDkeVOHtaiIoePbb8UPAYJb8FydX3
IgbCdEtPZ77VNdxLaB/UqH+6o1OJG1y3O93DeuXzIamTdJdRhUAWfqurRpfPehGRSDj0wmxvf+7i
h8PPpmwrm1uNoOIROLGbDWTRJQFQ6rmmJPw7tyG2Fkp/NuQwRNvI87njkCDhyLCp1mszLJ9waZ+J
uXkroVQph5x+k9SMgPOcbXVpUEGKtsJxQmmtV4KBTyHAVl7wARfXhUI3sWdkLQNNAzMQgnlQn7ji
elvVfzj9hKYLBW0Pwz+rvCMSvIOFUeabgAWKuVigx0rJTztixk0t5sWXbLDNUZnTFxlgudZLLlrd
5bbkfRbz423gL/eBgO4+s5gHn+F0WUxb/QMoF1XFxVO57X4d1q5RiVRNRo8hPZgrd8C5jsTfTytc
5VVOzkpwgf4Uc526tdqMdaCNHd/W1/2/8DZTrbfIp2HxexlqE6ZjFX9ur7ud5BjL/sMEEklm9Q6A
lhUKR61dJD5GN59kP2TP7sl60QpkmgjgsZinPWZ+QBvgrksUMuo+3X51218EH2KoJK5mLfIs18/c
ZlHgRUw8fJWW9Q3W2McDQVwnzPFTcHdNtUp9SfRV8wkuNEgRFWh7DHFnye28iv2phY9uXlE2sez2
PdO/+itNWZD73Fp+x9BeJH0IEiETEl8cTY8sNYlDicMB7RDun/JB/xUUEChJ+izRmvY/YshyOsX0
WNYyZpHRZiol2Ocms/Y6m4m8XRgE1yxgjx8IdJVx1m8F/KWWnQZC1t1wEh8ShznDS5ewr5dCCEX/
9HokfB/2qcdvRG8e6Dvmxl2/CVwMgTqhsDaTqCaEG08TxVYew3wRjbJS1l+8cma08NBeNeJ5WomW
TbT359Gwztlanr3biui8njsunIXuOnzGkWV1Fk/5PLT7RT7baVgb2cGYo7TrFaXkGUhSRe5NR2Un
8ND3u8qqxHuNmOhbR8j0NZRZzwyxKMqug12cK2Y0BI/u2GkmtkmDPmrNrUEV+plTKsl2Oi/uI0Li
KtB/TBXwoKoo9N9oCI40a1df7S5uxFXmdMLpnABpZx1fzE+t2or+G3rQ9YpLbbvTGAaKzQ3MH6Br
gZRjvfl87gZ0RI7IaVAilPimTXUXJhKsMJkFiPHTqdpqWe+xRdy/xe0T94ws5Xo9Wl/KkMhEhWkK
CnNRYP66tVMAe90rVgfynaVQWPmfIxTXT7xgXRv31+s/Q4MNf+uyUwQEZs1z4T8CGSFG6RP8jG2f
+CRhKH5fEa5uESDKznftSi2LN8h7MsS6W6vvP5r82dVd/4Fy/KPf5PwspbI9FJTXipmKW5tXb7h8
bJEx4raQR9mvuVybe7B8qN2NvT5gn7pXlLIGT1q5rE+4iFbGrAgnKtfzqsIiOyXMoBiG8tMAT4kx
6k4/USAN4dp9hZLCt1ZtvukaGrNkvfN06dDow2zrM0iYlgoTTwDfi3S+BpLKQ72lt0pqlkwyZmyc
Lks1okzwbEQA/CvJxKVt0IXCqDtojywG93R3EzLHzNYUKmToMHmtWNt0Mr1bDkhiHlZR5u+pZ69W
klkDRK2bWffutrL2HlvNWjzrTRZI+CW+YBn2+E29rmrvpU844sDBqdwXBwMg454gDL2dwNJBC2C5
FEiuTIjU3aCb/+LBsNbiWBxcDlJc5spvC98UJxUxP2QizeofcGEierA5CcmCPzvI1nzlbHam3l/x
cxA+bjqObfokTOXp6XuslppVhHMSKQZvnCZ7sLcJZd8FtU/XHfMg3yaSQ059QhDRCgvyOv9oTnvM
+zPtjM3OnKnmrTVuyWvC47GaKWnbkVTr+HmQSqQ67W9I06DfytEZ9JMEoURRdReI9poGCxkG/I/1
FqeKhHvKwsNo6G29TJRTo2kN0KOeQTbXjTBJIbgv68K/aFjMrDO4b0aHSnTM245KV9hoX5GGYvef
8aEH5D1LiCp//qe0fgaaQBfz5lEumVdFNLGHsnLXv6rVu//iP3UcrbYHeQZDL6cWubpOrPCMgjom
zvC63BtvTHdjlESmZ1MZwI7IK+7cUuskmO1NJHeF328aF09O6dM81bDJMiUm8pnij/LmEAU5AGLQ
i4TBbMMRqpeEQY+elf86NSdYiS+5b30fHm5gE8+PcmF7NiH6Hzw2JBOhjy+vYX2M6QMnkRIGWtKu
CcwV6w/ZXWEBA3s/ZQQ7ktJpwNnZpKREaXIY9sS0Fq58E/4z0lKtDfiESsMjd1nL4kuv8mdHY70j
Rx5dwizrSMNG4fUGA/KfRrayXbHF22spe80l8BE5j9rs6WkmgNVOrlcIUcj3LIt8K56irH0xN7h+
XuaZtX6wmthKdNJwjPkP+7l0tqsKsKcExhvY+1EBpVQtwmAsBbD8c8UdaeNUS4tIiaf3Rbu9UsAK
czFdJENx5GsIRa3vLmti54ZTACssPxrTQgVQju9xG0OsApTstEwLIGS2QKjYTmjGVWgp+uVPQmWS
yuUnNw0Y+/E54kXnOaCCk+ObxSqEXxHWGm/AFJuYTYd9V6XbjkpVOqlDhpCbLoMQOV49pOpk5Mz0
FHzbp9E4douYxCY4jIyOgImA62N4ULbIO0VfYcu8bw2tIyX2rbia/pqUNWtmJk3k+Ak0rNyclGWH
eYLal+va6IH3S2JlkX8Je5uQCYXIeiqdFY9hj4y7aoc1pzPEgwRnUifis+lt5/XwQ8he8X48HWzt
db/jTt8JdkNITeG+uzqx3eSima1zmJ7N+lVq6iGEq4fXURGpxlVrkZRRnMGQ+5h2RVs/DGkUV7VE
5LiXXtNRrTVF3kNj7wqQUF9h4YpR38gJ4A3ypgnckn7JlqGekXRieO7MSz6hjc+Ca9pvp79efKaG
J3A4wJUn8JGSciW9NK15d0PHwt7tON958Gdyq7n3yUCdItzgEGB/y/y2h0bTGEGzDR0m/dllVaWH
+0F+i4xprKV6CiCzYZX2KguqYsLJTDGa0cqa+y1Rf03EmG6qDfrWrztCv5H+bxbAAnFFyFO1EATD
D0tBdWBFjSSS5Djwr63R5CirFcp/akCYJ+0Qa6GWvmrMP8chclp0N4Qq/8XfJF93udOXQ2Ivmx5R
4T9diCPczkJ3Zm79fqIXLmH47bYAH64iJ8PrJkq6cXWetYTr0Z+3pf7nfmHnGr1b9h7ssG0zmZGd
cQIt4AIQvuDlz7P6LLib157NzX4/3LcAb7fXmIk8AzM+sB6uKshVDtTgn9sE4Oz4NxRipI9GLy93
R3S1vVTDD3T16DZTbM2kpBRi4xMhreczi0IsP1Vhz792kU1BQRA8xg0AavCnHBccqsCah1uob9uE
qpfT4HGTrtqU2F+qxE1/sDH3ark/ZAyiPfh+gZ+PBMJzkf8TyNIK0VGqnPH31qn0QA9PO3LoCBWb
Dmzy75o5Rif33DmWp64hX9ECdY1UgQX6eKeE1ocHU1fLgDAK7dFVgfhTQiUx8D41Dsd6FpctUPKW
0eUiJGsEY41wB5ZR2bUoSysAOIUSHJVUAcuJQ+MXo7xnY2pjZxhe5UkORU/unyUGR3ADC9R3ep+n
g2kZO4ANyyc3/U5xLJUYJR1wc/lbZ98v4KYT7GYlSN6L4EaEgf0/3pKxylGzwh9sT2ZwlLD5+yR0
OK8p6SbAC75TdIa+aBdxuYyViV57biUF71D7yse8bvzCV6tQEc4dZidfLbnO1ZHsu6QThUiQtRJ0
ucSfasqHGZWFgM/Vb3jT+fpLUiBGwKPBSK7n6CwHzUrGzBewEkBnTycKFJ4LPx5V0GZ+8t6HZPzr
4m+j6oFB9yra+QwwrMS3t+/kCL5DLA6odi/baZndaSAQOvUJ+fklMu6Og4hq9m6K5gpXYMmThbPS
kHcmhek/gt78vx4SfJMsUT1UjG7Oj+4lLftL/xAP7erQuMnFafaqz+bhjPNaHnxJOi5JxOHt4Qqb
/sg792pp9oPRpc1jNxSXLdLqFbNoB+JqDIuTGf2C3MvmgF/+ihAGrPwfstrmz5noq3u5vgEq3fOI
VL/McnBOiST0y1jCxK6VNk9ckhU16UUUIk15Rwjw/ueT/cm8/OVDK9TSgsiEuxIFDqmC+FxGoTjY
BivgfxxLRn657Cqqix+uCrr86PlZbNZeVKKvl7KL3SR2rPOS01fYX3eRcmP511N/XMd265D/Xhyu
bOgjouy3eV7knoj0Ga9zWNKcDceWOfMtCpEzgHwxcnLj8OEmWTFsQL603c46DNWiAF2xM8/KOi1S
mnB2UX+JRYE6zHoTBmdz9FOMD6lxn4V6D1TG4PSJvlzoMelfpqceX2TsfSM/4JTvnrow4Ow9xTLc
82pUV7xqBGlciq6Cl43QFVlcpv2lkDzZaOFm9sBMRsjQqcmE5C0QimO8wQUZEN2+1rsvCtZ2HlxS
8+tCTsLx2sXh3QUS0PT5GN6hI7FTh0L1JXAszc2coMYz8xZLyMYMsa8iNflRw6PQl6gYpZE/6QdR
om8+WXi/eUH3AU//8iPN/mHmWf8pMR2x4sNYt8THNm1anqP/QNvW9DEs7BS7cMR6McKSYPmy3+SL
+1BS9Bc8JxP68Ej8DOHdfqyd9c/leGcE2yk2a78CfiG6Udu5IvJPoPWvzXZMTsXW4q6GkcYhHdvN
3UZBPSK5nXCEG/P1S8Vky0cWPXI5PXKadXYTwEa93JlPl8xoPi+cMH8X7qbmK/UgB0zm4LTrpzq2
vVtoIJBY/MklcIJBNRk2TJJV1sPJF/F7mdCX0vmdegB+Mr/e49suP09E/zPTGCfcm6sBsieF2NOm
lOZrpc2KxT6cbFWgKwPOWJ0Bb/7xFzSuWxxflUDyuEZzIw84Jr2tFHzD7WMQ6y3A5tMup4ZeIowz
tovtuxzN7SYhBD85rlG6xi2aFN+7aT1AN3XSnP50M6hGH6u7pYa31MPBDmjfGL1X9WZlbtBg76JZ
V80Fi2S7pyAotRd5hP4/I45uKc++eaLQTnvIjj/VV5pfLrryeoDekgbXhXAyJWMVANkvVlHNu3kT
gi+vAEIO9Fnhky2jtm1P2U/Y/lJ+ZPwx97LpSctmrh4ZAVr2dIH1LXl0s9BE7njfj3xR3U2Cs/HC
O5if1oLcUHOg7ks5yWjV/vy3a830V7Y4ITetJmYE9eC/10yjM8l0cAP5PBG3OyHnQ5WEsnfpQXOo
gAFC0O5eamjWmr6tjKDb1dnfFFbbvaCzzYV3aKNfjxyYhsHI0OL5CVTAF3B+8yFnbnUG/JcULvax
aVp3BpvarlGIdtLj5Zq8fmwN7TxBtPaefbG/2/9wzBn+4H/sGVCmdSBgvkjmoPhkhC1Z7euZg9z2
f4hbn3o4tMzGswO29Hd0qWd9U05G5V34TUSI5Pr+nBBIjQPC1XhqHNzFhSgVp3s+tteVhfHZsltw
O753X43ycNHp2FmNVAuxaQLOzCpM4eDwSUDG99NbgYfafgAO+n3s1oiIzBUO2EOzk/IsN9KDmGpD
nsVJp89LpUIzN18nlPkRLlSI0qa3rsvAa2AZU7S+aMIFEZU2qmvpoPcFtRJxQKDLwhpPag0pD7UD
8CxBQHHYg95+w76S4bmzb7t2k1q7fBhms6uYM+9JRkrLAtcmPj6tybsodVQoB3WmABHkP8vc2RoV
a1zXEWc2QlxOOMrvrWuAG6YxREFrtJugkA2bkIccyjlR04SKpv5f2PVIOAFaIILcEo5Mnjo25HGA
qZiIiqnMmYQzN6fZGdG/rLizRQA4hyN6fKPMzdwGdDXtTuKd20OpPtJubY18tzLRlBjYvUUjE6tq
HHgI/p/KdycvZFVqDVTl4v35Q750DZyvbpbQ8vmEJWLXJDcT5PO3lT01so3jZqNUjSL31vde43ip
uEFV004X/9MomTWWW5F0ZX8ZBrKNo1xJJ9n1ud1rBza43s2E94Xx1rdZFh+ubI0VoqI6RdB46Fd/
id9FJ0ddQyhFEy1l7pvUc0+OPIt3zw2OWaHvgJMu03U1MI8Vv6AX7vrubvrQqAy9ys/U5Qn49rh7
lguiUS8BbHS9DHqi5VRKd2FZUPgmxR3qCKBLC6/1VyF98akOIk88MueM8CRf50ohOTvmO8fBVHqZ
f6QQt65iWM9DLL70rkiQ81hd4XTqzcKVcCKSX1GTnh27CumlyOtqRbSP7lCuSZQcqcn/cnbqLfDs
JqAO7Ig0Iluaw6LNntio2s8uNKZJH5ce9BO/UTc18G49MHb20wsPOHdGY//Rol4DUpegBX+2tkgs
SuveF+mKrHnr3myr2J0p5jMxlZM9DF2rVku8Gs8WEF3dxttVngn6dktqk1xFT9nMh/6OTpyZQzJd
DIEjbM/WdSSUEtH+NFzSa8skUP+OCrYKMbneQkFBbBCbwTdzmnL4ZN2X8i+9JLBJMv2gDGrmu4tU
qGX3jan3iQMnWGGOd0b1n3rZYswI6mFZmQ+MZxmJwb/jWmnGuButQ1deJJN+cO/gVfx6na7h8b03
dSDeCG5kSrOvkn+qvTia10PUSLQ+MSETAY6RDLWc/zHmI59XwQvP1kNy6KwdCpCSkPufPdoFgbNo
1wD32ZkK80NEgC3Z0JbtalB3pmFB+uApVpUQg7rAh+lelAYmnZa5ANOeJd3gnITF/Px+EoJJ8lNa
7GcIstnTT9i6dXSSJes2hAgnuDZVeChSCrHxWJE9DVnVwRT5Pb6WwTKXYZQDx0vnezvzy32ei19B
VEnlul+V/51gPg1MfnPX+HTxqMDE3Z/KEyP1WyveoIecH4Wn5A2oPzx4/Uaw3DtUSPWtbD+Y0QQO
+QivhGSXIm/TPEzJiby7X5nzqUbSQaHJyiy9F7rLWPmeXxbreW4c9snlvmA1T20CbaIgpszcXMcO
bM8sYNmZSf080KxqBL0UgWXxampuP2w1/BiBP/UvUwIRGXvtL3N1b/i+AjxnSP5jYN67cAYFfT98
vZQFE+8Vfm3uEuqSmYwxmIOXFumcKV4xlNg6UaB4/4ai2ZAjsbS0qfLm0VL9pV8LwdNCZc0qC2nn
LWR7Zm//TjdyIHsH/D25OK3FBW/VbCTGDkqm2eyJE2F9Zsj1mTjbucL5qomQ0h6dogfCQbuCwk0/
XUejyKFFfcFBLDeivnVoGvSZQe7CY2AB8Pil4zszLnWBbPN+qIRVjOxvtBGFwcvBEUAS8m1g4xJ0
onEg9VEa7oFbjHF3MFMhw/KDuiaxvgs2dyic9pjQ8ZoXOah6pv4ocTNAuRtLJR0HfePxG9xlL1er
vCPu5/r57bhWdGm+owzbvpLaJO4BjCXazy7LQJhAvgqtW4QpLV6+zds3RK+oDcgMa+UdNge3wD8P
R4D5h0w+2+LZazpn0XiM7vNaaP0t/Ee1RS1sq2AwLdyWCGlsRUR9ySZWmghpSG0tMY1+H07vW7EC
5Cp5TuHH4W6agVnhkOg3n63umIaN1UVOoFu8t9ZYvYfoxjEmf3Dv+CiMdG5btqLVXiuLHRMpbGxz
RndRE6cqRZYBqLjCxOH255UWtalpiImBiPwkpJ5I8xEyYwA8JmyOZ0mJREgsrfWipaOf7NSvtSFN
JR1tzgKPKGTJK9nuTHb3Nwx5LMzK3mK9DrMdtmD85/Y8K4pBWJw1tGFYZ3wRFtD0AcHp1O/37fP3
j6q/WpbL7nsgKrWTq93nIs8ihpCdoA4HyhHPnXtEtD+U5pfrbAL/aKRkQkpwq5YVBg4ms2duBqhi
/9XUbK5Sxsakxx+WHX5zTM6VlS2n36mCMUQ4mwaQULNON47jzukO7uhZT2OwZlNTKgsbE6Cc1+zT
IYnJlkcmo0K4m/3YoX6GyCW9tRkXQBlpEF/jBRnjPFD0LlylwKdueKSD2Gnpax8F15H62eNFstTh
+9MiqBffaFIFhkAZ1kY5ztsE7LNfMUFrhCyrMiEmX4Lca1v+1ticUHjY9LucdGQefMkl2KgfJd7/
pPhRUYqEnWndG0jpO5dfmKnZeqIyQLgoY1/XLmzGIdSOpeeg771Nrywn04TblCcC8t3NJZ7j/2we
S3iLodNZSsGz9fOnrYL68jYAH7yw/WYJ+J3u2sccXtU0G8CeHNsMDwVggGhhdsKsd7zLmQTi+v+3
zRWdI6w7faqQkpLNZzYBoUAG69gkM/DAP01/t4pGvL2InIkcO2YOznuVSCZnVuJrJEyqB0FjAm6b
0awYkv0HE/eC9R73gUS2THJctgAKQIwTTy1sCZzjDI8ktU8l9qyqiJEd7ySJsLBoHyuVjdoE48AE
UhGjb724dJVGgO+yxZVt4WXMHKVsz1b/D7lxfYgV8dnLgTlmiP9vziSAHrwA4YhF97w/1wQvZhXC
Qd+4VkgkUWtoY1hHZZPFlv1m/8QZ/XqEabrm/9YpUt8PqQrXkOvcMmnGi5aKMEXlsU2lMgos6pQj
/mR7khlmJqfUIR9PtzSK5HQXLEZCTwWW4dl3nImbBAQSJyH5pz6zOaMd4DN4qSWBFBS5y60+r3xw
wAJKfbv2mYrywil9n2+HxFV8qy1mAUnUgdQHYJIlcugx1XeOoQKxEVI3Qgvi827SNWapJOmDUAX6
ChhWPSWdhdTsvwFHFb5mOg9H+cZJ/JkH+YYSjs8QL/dzEH/D5wyuFxReN998wmYeKpkjfd+qN/7k
7ZUoln2YxnAVcCKCep1b025lrUFvXDObL5WdYFTZrHzI3O+aHsZxT+AdJia7H+cfZf7GueegCLgb
QXFRE8LW6da4qu0xn07F5HYHKq+i9QtsDb8mgsOfoLQpd0UhQjXb3CxbUBYeOCddSFUw8NeOcwgA
xK23p6JDCp/zgKkNbzyDNJDugpf1OeC8eiB49SfPnIDVvfVuvTOhw7/wVQ3kK5uD28KycvdekTA9
8N2+PnZBTpD/9TWeaMPfEgTK6dH0xofAOJKTB3mHSpRPfUgdkmFYVxtKws6ziLLl4O+rRqRBdoYX
vJVaDtsC918ApNloseWSZKxNrKqM870bcr6GOo/qnMXyzbSAHMwEipZoGCWRZbxrNEQogS8TMQ2h
Zl6GjNbO1aMWLskL8szItBhrsGnXf8i0nNdGMBi/jmI6vdplgesOBFOKblphVhvTj0GyMotlC2VT
eEtRXJiZAyoXq4PdkC9328XYB0XzrcMUJBY6fkK8WeRFbXa3KMIMXjE6mtv9OI7XT5BSvH6tejET
6TmHB3BIdyl8Y0MZu1EwStZwZ1TfkXQ2LP3nieUCElTuRsn/hAKI5Gjrxvhew5S8Jj7v67mrvyzY
JBm23608/T/J+pC2qW8kRcXFB/wN6eNYH6jw+HcpXv+bVST92cWtAp6/EJVmZWlKKh1W1IycxEXg
CFqwiqZ9Yte9rJUIUa51BRJS89ERNDXD+H+JuzT0QLIRk7dDGQu7QzFelP9iz1FywT6bjZpZ8EFs
bNoE+zwb/dYPFiEOfg2l8GME07HEYoERkB2UHwdMs6yMIVnO2uKJNcCckjgAmV7nWAzo9/PcTswa
L9B0XeZhrp7y7jT0myKPYtkMreRfSj6Bz8eCktHxQdQ81BEK9Gy+T87+aXY1nNY43lnuVVsPdS12
HWf0q73y4C8AySAai2gi5QRu1hOIhtFAAoQ8s6dggrZ2sMI+c4cYKbvyHA7jtEe7LRyKERIp0FcL
IDmoL8IRfDQDMfu7kX0WJhorwofgZzb7+XBUZmaQrY0UE+DBePCdgMeNc8NibQurGLtFhTGrR0rr
+FUul+fhLvKg84qWlxwwkiYC6OW80vFQd6aJvBQazwlkX/KX+oTjye1JhsVFPtIU6M6a/GPLiLz7
VB4wfRhbH+s5CisXrKAd7WDE9CKLK64rxBskkcD+U3sc6VOV+DPnR8bDi6Gw9adNad2xz+XuUrlR
UjdIOlt5nnIRiy2PpfeDM4bQqtgAy1Fp+i1+t3XHtm6LCNbUCJxNdAsJ3Ne3XbaFHfXcxVp0vBOV
iaakgXabnp8dx6/THZAvztUn1QzxOr10a9zATEEU9sVRBFBsr651vq8su0a+k4oHnd1tuNVeYYn8
5mMG+OuppqArK/C9qPfFKiaoK0AGBOzqVJPDFupMkkTfRyRoeEfPzzgjgV508ssgD72CJp/nLCxI
MTY4cPIdC8k/rG7Q/LtkjvLUvnjEeKLujkVm/b4//DRSZN+WX0mSkf8EwUkahLY2NdBH0YKo2I/r
LOlcASUyZEee6StSPSYwz72Dvr+7J90OGAe/JH6jKOdWdMIVIpZ8fmYN++O5SufOmonP6Z8+uptj
egpyDggYHTWhgPCn+CKxUT1TDtA/+7+Sc7VTBAPdQ0FAIo4A4rb7cYBN4hleQTbkt8bQkxQw1LiO
GewDWQtjAC3OTZIuCHDVhgop+GgunvbtkVtX9mawIjX8TZCHs9iFiEyeMw6iOI+7PDDkCij4GXJ0
4p9FolZGKW8o61W4E/HZDJxKpgMXw4IItd6Ur1gjatzDnm9ddYtsG8OZrAe+cq2u39vRV3HlMBa3
AzHZZ9MVpS6JtHL5eM6OAUki4aKQhAG8wR7uUmn4xo6DQAph7xEXyvDCgTpPTlg7Xe9KaFSC0K5s
BCkfb6xV31jRtixJ6CjihobK61dRN06SG6KVQhiQNJukJ9UxfDXB5kORpsH9bXo7WlbCaBYobN+P
bcblYJ0kpzf2E5Miu59XaGU4xxsgAUp6ZgV/95VKRx1pwdMDLxcEoCIk7NGYJyedAA2qC2ycDwLQ
r8dJV9vYhVfBrLJ7Z/CI4GgGDzDPagZYHtAFIa+fRWWuEfC7PAVmkeQmF7aHZB5Wuy10nzDdbqTF
23WaHw2Ss5zZDDWNRHW+Oq27qoiEtvnvGfpJwSk9vkm+5xNmuBI8x3WzGG3L+0pf9G0ViEY5JCyP
a2hWCsTf/KAmsI+EhhZWECEYxhXqUV/9Jz2qEQ2foakMRQSjb9SBqCKn3iKBk1bC1V+7jH5Qbf4N
g9i8oBiewGVoAJO9K3clTT9uH0/NQWnAyUSPRanSKH5xBUAaiyyXJRQ7Rv82/TpPDAZgj8H5La7O
wQ2EIIz5o05IO8oPK5CgsAQcsI9GOmHWNgvG1+mmTyGfA/t4XKwuE7VEhIlBex7doKruRcP1XwyD
xPqa1RiTKYCc2K7DXL9FJfkZ9PzjTq4N/nmlHBojxtIs4XRxEi7OY/etYzZ0ieVffYLoAK/hnvcK
UCDXLRorekhd+o/BlDN5z5xMd++Q+gErugJ888ngOgEBjkMjIg6/WJUgnmVRBe7Y6ZWx9qShgACP
oQeYXhwoj9vS/6Yk5jFUK7+B/SbaptXp8jPtTQ8wi1BIklG6Gr8WTSskJftUHBQ4IpqHx0cncwom
FVCMjeoC6LROfLXQ6gEHtVyuN3s3QoTg6wdi/pzh/rtCIazI/rnBRPMgANH6bOOWpQxu+E7l6mK8
nuhpwJzcXEhPTVscKz+JlU0sZKlaMfT6dU2lspy4S+GeWGBBhwb/xVXUeFsCNt41cKRa9yT4RDAv
GtuwHrlbD44g6uVjO/fk+BQOOoBDyHPpTvoeintRoAvDykiF0TqeUmHNK43RoPZMOBdfpRR5vugg
FMKuWZXUZislCfhKZIvNRR9EUyWHO2dSepWvjWJ+CW34Kuzag6eWnOIWu/R+wL2IJLXJYc9vlgTO
vmN7pSRCJO8iG3nUJOw6I5ySqpmpjOyp9QnkeD88/xnIGWNGVC4apgpLDggC0uiKqqx8ioBnbxrs
cqi9tSKaJUgfqN9rpXWXFzW+bIxmyn9AxpoyIDutZIWGtr2265ZUgxlT2p7SxrmXNSObZp8TZI4d
6JzF/ti9uubwWye+pMnwoNmqRAelzRso2eh3K3pSA5H7CQzPpKDIstwvMplycEJHMhj18PMj2n+9
0byzWMeTFPoX77HOJpHJQ1TYLK7TTjrQTfNMBnRQRULz1wI3r5TH/zUB0/ZlKMZ+jVXOx9pzrOtj
kJ49fDE/+jDfwU6TBQB22LSh0IbGRMVoDve9gvrfZODHZKYd0yzTEiR+IhD/JGVKi9YJuinONZSP
VoaDZD3SQAlmG2FXtyojBGAlknneYV5yv9s8QsBYxK2BKO5sDeRddTIWKtqdvPn4301XS1kW4RfK
/PucEIdTQ62OLudcnkjaFnDhRM6Q8mxTfa7BSMfGkx9ZuTtBiMOT7pHlabeVJ94oevRshvwpwhch
HuTCh7sI2G6/V/YN7jTB4C8vG9qpEh2C3b4m14zneOiaL1oA01sPmvaThfYT07X+4KFuuHgI+9ji
yEtsAhh1lpD1v0pisFtKvlPL7lH86nB+iLHep+AKkuLG8JbM27Ma5ovgDmfhwNPN+g8oKpMjfW7J
P86EjgBTVhKHb16J7Yk4xlW7WW30E6/M3oZ/JXJEqZQGqEoOM1fbOzJ+Yt5J4mRyC76JLRKv9T8p
6uu0ASKYG/WveQPDUT1o08ebMEpKlQ9qWvGAUXfkZoh56U15HJ45XaqbtxQyA0T3aA/L73zCAmlc
WJUjnzPduF+d08qdKL7qa0xCAiSUiSp7AYjgnFxgMOgIA64kAKJUz8qz4+ueKLxpsGtZAHhYIK5x
iQfl3Thd0NWtmqWfI/pXRNZCj+Cjt0E1bUIjvuSdZqiBjoHb3sjZXKcPyH+ltwg6loj3SJd7qy/H
AlKthHJum2HOiqIAvF60EYqaH6acuY4MzyFba6qllrS90n/WsJRDFqxv00HjcdgkPkpE3HormCJ4
dSvpCPpXgaqYrC8EuoHHcMmBlUA366hadnCoyI8g+STpYKBHyanbYnZsnnbDoWnEVJzBb8yN4ib+
aDM5rbTgHEG79f7fwSDGfJAcAvLpO88Ycy/Z4ri8opz/Gboy4uO4Xt9h4Q/8iIyMNgFKGHIiiOpN
SC8pB+/w+v+pUu3QL2mKa8RIrV5Xupg/dogP9760KZZ6Dgu8zAjC3p8kVsrMNoRVY6owhxz4kFqy
qNyUsfiu8FeLyO+Hy8Kx5/RUC2jmIAAvRNRaA4dpndq3wvypBt1P+Swui1Hyh37OWXCW23omOTpH
lQNLCJuKswtga07R04+OjuAK9/RJt7hNR2pDUSxqCQhm/NebcNqXX4tgXTha8EWSogVdaES48WIQ
40JtZ+EdX2R+bxyBcjBO8YK8JQFn+iZc2yfKSym26Lgk5GP5XaKsdgyOUGM4/mTiLgH8Frja1Ocn
DSqfNKJ9ecqCDLcP6wtdPAI210K++lA5YP/TXozA3NP/C9hw7h1ec+2zIzA116VPI+Rt1MzNLlga
VpcYRSeulePkNp2gF4SCOM+fKdJzKww5tneHL0sObCsGu4uxSKKs3Z3bfU8uVgkF86CZrrYaGAbk
y17pJAHYPdJvPzeS65iUKjBpkhZtIIKUVlqVCXzDgciFy/5K4gxovKOF4C7r6xLAzdUmhchlIerW
LxWvW7BJtBsWCHIi9xTslxvsv0Mqongope6EW/5fq0nnN9mIdZ2WvTlq3zb/0OSUHZ7h/xVwhddH
10vK65mVhWayMjA+v+Ka897il8zMAxMJU+yrbsXnEVE0aPf8aE4Gq7WeYsQGHvbEI0C4nyKq9tsa
PHJJ2zVvfgkoB/TVZs3V6EX7epZdqycae4JOJJoIjXMAyaUgGP07z7nPRusorazqIxD9mACOOb4I
iL75a0OK7VJYvWL2byTwoUHoilp3ZR4y1XmmxCY36x+eOeaZu51kxhr57hhx7/YQyaIxGoegAgtd
Op3TK++Jn0iG1Kllew8CTGnt+mBKG0dDyClmu8m5o4mPn0QJMLtw1tKRMehz9D/2M9kgScneK0yV
0reGBLRicwR1aogqSWS/XBSakAK9Z+x48i9Rf4SH30ywEnu31xQngezh69zYYto5NJCaGKYnBPgg
en5Gdtzr8ecdkxj/0ij/4Gn4CmzkOjwxNRyqblf7LbQPzj3pQS42k9kLS494q9Tk/PkX5VMcUPrp
l4DMgwuZGCmwB8xPd7c7Yxt+LXHbSFNYkt1XFzuh79kV8RHizXWToBgN/fRrqXKhYwgNqUpAPB+Y
4I2d2GLO+PxoGoP17j/3Dv2wD0olJpVgMgd4MUffE7xMPRJ+OqknYW/4DgfmnLaV38L7Cm6JzOa1
Bi2GLF1TJOI28H2wIVnoaFgLwFzVPzL/f48HTdyWO/uCAQcrrMPD7aLci0TiQtvoa4fviUiIQc8b
8FaC3Jes0yLRZpqqT4mdiXZ+CqFIiNTH5TYyGc2n+/nFIR/HIbd3giT6zJzMhKOT7At05cdVvedi
JlC4mLCgLdTrupapvyiEnPQmGSBcAecnKO3OMUjYHpC+55hPK2kR5PUncDuCIAKPsEiDocSksH6B
yVW0o4MVzX6tPYzyDRXfBxQk3NzSvB0RgOyqGuBA1EhLvTgtHNdRNgqg52EBZDpg16dEHU2Z/Ed+
ZIhO68PS3zHrbj9ReWk3Pvir8pBRpnmDKPZmCfK60stLjnHRKoLYfZDndJS0X/rRZh0x2OJiOQwm
MsLIpPSbHwzieO53SUJcXfndTwjf4ByNGtQUZaqRlWjqTmST/G4qEC9ndeboHs2pHKCGYPOmhdtf
S4ZhHexXE2hqeD+O1OFWBqWu8WYRW6vfFsJ7zedtt+DZ37auSC+InACU1AMnJpuJ3b4xq8F/Nq7G
x/l228jm8H/B2qXIauEWM2On/NujaYLbmH4EmHFXM3szQcJsiObjwOLFkZEaqVu1ji6WutrKEsQj
UIerQDQp+qxdTvl2iqY7bku4QPbQ4tyzgt5qIlrljceYirA61Bibzbv9lI/f3yBD32uxtOYKoppN
/817tO4Th9UPT2NfM/mnlnbwXUEoOVWBPSqk5o+YVZtcqHecH4hzV/EaCZoICyFlRnyU9TLtoxi+
iFr1btxIBBfTehQWlM5qPiG3HgcWjbGGC+m3gwp40Fqihs6kPx1zdclBOPfS4Eu4SRWIFi14F4Uh
8XaJhO+eRw4rrcDjORaoO7OqWxKzdAZOd1qf294CnxkeIkjjujVpep6vDxaZDoCS9rI7bfM+pN/m
iPD9z7Y2WeXt/jqdpvyHKpgglm9cRDQsiTPUDPJl3dYzDEHDVLAE1sggCBQ3LXNy/PqHZwUa4WeM
6moIud4uHlUBHYzYmhL2jlJpuXToVmmxGEDeinjYWW8UnpTbjaTFdSn2P2BVU3PTTcXK3/eQWA75
zNRYV73DTlXMNO5egwm5RLXu9huufsw6eGFyzziVfOKEhZAscpVixItobe5xPkAH9Fw7hBwnhAWf
zcaZTS/Sf8oRbEHPM97v12Oz61Ge4xy/BXyBKmJM+6MZamo51IUPQUN0JVRzwQTXi+34FjO/10JJ
iGMHz1E6hJmwy2f/EpOHn7MvxKRgolyYYtnGkC1BUOcPaPHRpWE4DILBXNl6MWXK1u/fZXv+TpXV
mKmlcELpDmduaZqnVeJxgnslPu5PrmVJnlblF6RDhmIS540/JnO9p9t7tIfuCDtO25hqeTD1+kGk
ebFblHbOwBdCjDTrPz3jKOCZJWR5zKrxCew3zaVZ6EgQXr6TYrqr1Y286WgGoqoC4UbMrplRn7hA
8B0WOUbi3Uxf1BwgxcLAL/MZFfeDhXM9u0FrBWrLEIPoXZ85xcr3ROWJFfvTipz7vu9kN1DPD0dZ
7gW+hLT2xFToO1FHww1TGbSQ+87k5En1+xLxPvpKOtjLDlWDx/1cNRVq/OJYv4/EwqEaxphJK7pR
KjTKiZraLl/N0ApHytgrYfhgAREighPvm0QqxYOZdKT1KYGEhYtcXbh8aaUWc3jerulHt90COjys
0h3Qu9sSSfPV1J+STsTybjqGn+PnYfarUgLHz+rDBxpPfRIcIDe+YS2kdlWe0cJ1a3L43UgZIaHC
ANZjfe6Aw7WD0vVvL6xm72xLNxR+0N0xyJox4YMR0e1/3SzkZcerSzFK0ZNOwEs8Ya1ZQXREi7zQ
jd9lDSbpVN2gSb0Ch5zxeSxTzmVUjuMV31AYXSfdH6x0DUIF00WNfqHLnjhS3Yg0j5eZ/1wMRyIi
iS4oDd4fEKDUlhwzDva52jg3n2GwbrpQ7JvCPh8Qh9z/xgCkla8qc2iubPuNvUOjEYwTeNRL4rV8
B+HIOU2sumlu1s1TL0JW/1bO5Dd7L+iUpRhPFx55UeQGJB5x9WWaz051WWHIoDEdhJDQ7wnJnSvZ
itf+IjRg3Za70+1yPK9D9A4R/dztTE26gd6KMJweMvEErfv86054vbN4ll3//KClGL9gGkKJbRDh
9fLDknvWPTOPoeQb6XmQoQOFE36ucRZuLg/tpz9yWaKSKCdCU3ygmQq0B54lwejt4fwYgO0vQZR4
BNPy8VpMgohpqgYHw0KA0G0gDgmeRnOGoeB6HJO4aP/RHuTwZ9vJCPAcFwERteviq9XT2heiWCVh
dMgz6hjVgmvwijexZO80qEKQYiWWKNmYkSX05C3+/mDau5/g4/TZb1b0yla3uLzZzYduh/jKFkCS
gcX2lYnWXpFMnz9xj8/VBmx6ktumdARSA209xzNVUOjP0UGqrVDY/7igBkCYcdw3euumI1v/Ej2I
6IfYOdWIDT4SIT3qEsg4I+c5TLU4T7gWYqDCx8dgxr+GUHehkPKaBit7QXuu5rs5f16OeasYY09y
ZJ7IAMAr1266lnmhkks45zLOobYIvleEL5+2O8AvvWS9e6YpqhmSawpuriqMcsbCbHL8T79VRJHW
2B280hadn9ytDG6/RooLZFwimSTZqhvnLwSe1aa++2vegN6czcBrSzZjJ0v2uPD2EiEqvQZBgtUo
W3iCqPGS6NL2YD+KINg0EN+7Cd4g1qPpmoNxrJbxFeisA5UoNJcIJwxqPRjlyH1BQy3TYO1P0tAA
eRXwjR1aQUZFbZq9LznGzSfwz4lOUgxOSLeqgDWW+adoIdscvgYk8bzQZteUYy+juk68/3JXg302
EnkTYLz7/INFTsvDX41VpmwbRhkSxqFdIkcRTRJhRhFqzsCLPWyU/1LprxIycYF2p97BqemeDyDM
kRTQABaBXUda19EkNVyelM9BDxzN82n2NEDF5HaxOw3lnAG0FurukBEclYvys+Vje4rF/G9mWZP2
bFNCrtcGXihDtw5kDJ6KOPe2ApSE/1JRFpD3v+CnBAzed2j1v0n4Ehfush9tnrNN60JLMIV/Uhtb
5vKXxDvX65YEZ1RIyRV/yrod4HMtbaLShIKTjEf3eVduAxKXH9E/jY80KMFXrUD+yveRFENDOOtg
LFVIFt262L0WPJ7sB9HrKxKY8nuebIWyC3phFKy2ixZRqPqX1eq3Iokzf0eDeVxIiU4+PUpAj/jG
9C/c0k1USPOnC63QfdzTEs+KNQTq1Hf0pO1JvcxsF1p2LCyC3IHAuzUbKf7Itnnrr7jn0Nc5Iq2T
Ha8udkAUKHLKfDd2Taz77G5D85+ivQSmolXZNL7K+RgSdKyTrR1DdPv4vzV8g1VAWfpemv4dqURj
ZTEXN1KbPhEVgZd5r8ZEExl8lKXWmvkoDSgNYPooaQawxZ0CwljCSA0kwA6SZ3SY/lBcX5HfnkDp
WkUmb6LfZxxXeNUtRj226n60voyzyxV/pPPLwqjzYtQCg6Zllx3hvXGjO8F3ViFypxLgs8soDtlk
/1p6T7RlBCem0tzTPgj4ND4N899AXzvqL7M+sPv664B2PGm1ynf7yRUu1S5pmFn+bM11bSWkFLp3
f8v3NZT0Bvm0sAjg6MCzOH38IFLwyvYfeR6iqeRpOdhTmkt1wyKMiwIRegbfmeHN3qzHjHe6QTSR
NIY0ZjMAYWY5WyY4eroiuu4jkBxScHdUsXpXIy8mwSbD9Uw79Hh5g03W/hS3HZv5A3z6/Xjrglty
Z73zj5rThCwR99bCdddU3LEh9UDdFVQ9Sszc0FQgrJOfX3w3KBITHQBbtoo8nB6yigPuSComBnzz
Td70JUZKrvUEvb1QP4As67YN8OKw7mhzLlvuQPG4ssO0UOlmg31V+86nF04F6J6jLNAkgcv6xRAp
vJXwukvqxvRxlf3C6v5g1KiPARCl29F4bGiHhN7cqFwZcfA4qGdJ2bwX4/XnfdmY7Hg7e9gw4Gnv
yxViiCrpaSstnhT2wrGBv8XpXX+K4g0kSfK48X86TKMA/uiEPopzy+utU1HY2BvQnYSDHZ/qrAeE
aVO2l7WPNBw+nNBJYn5pvzBg5zKYkiJespJZl+LT+x/95FYgH0QKZubX/5qekeArmeAaIbkDgAm7
5peLzxD0AusBezFSK2xQg9Av48OVhh/dWJ4I62STmmpYAiliPkrpoPKY+21aoDbjgy4mUdBKNktW
R0DIGYl9mtwrIEedVI1cUxL+y/l3HkSHlQ7GEARwTXtvi+MqlQF+xIXaHmXS682Qjp4LxShThFCl
ptvowV7U0KxuxZcbEtpO1kNgouNbfd8y74Ofdr20Wo1QTd6yZqpZrLTpyKgf+LKzRsCzca0FFS8L
fnuKll0KASS2Nsb6WyEtvmoQ1fwhybYvPWymzyQD0s+VFIK6nKIJMgvZ7pSzoRqstXvNU45AJGnE
KWS//DNrZlSgXqQ9E1sHyz5WVMFsQ78YfBON1c3Oqz1LzXSJPzuK8Yo5JE4LAsnwX14l3itZ6ESB
USdU4Tg3t1hx9+QcUkFPJPXSnT4itJkuLwMPS384KmDmphxi7ZjYpMTjSjmognMhjdcEZL0h7aoy
XjNrGA0hSUasWcjUVshobVpILqsbSB9rY9Je2iSXtJ26Cqb6u4YayzLqXAK8mTW+hIYj7cPeSvN8
wq089sExVyBaiRrCpSi2JHRrnGxQWTxHaSYN1aoU0qAurCabbPGiw/YVGeeLsN4AV1DYEmXGYSjd
VfQr2x2fj+K4BlWA4H9/CJMConSJe+L3D0uEm/x4BtK2JmXtwBJoA8/WF+TlpGOaVw42bOA/higH
QVVDiGKRxMhG/LMGPBNP1ocYmR2kUyyFq597wpD1L1wQaflyWcZkQf0WNOLktzMEUTo59Xh3feQA
AWGzrh2fbNjY6BY2xYfM41mPT7h2+efStBwxMOqnZEKegskaQCO4wm0uRom1iZKomIG/qzhHagZW
j9xptby0bpsccS/buFaIZkoEwu7Vm2rGXQNYZg/7Gs7wr0w4asqufZasN9YKHcah7ttVcwTtWdY+
ZsFSHogpWi559ibz27krbDZgN343SzHCrQxhLzkRvSkQfv8QyROMb9sh/RMO3OrsGLctVOBsblKQ
JSImYsPL8CHarM0Bp/FJSAA4JJ+m4aC6bHksawdN3rT+PbX3A9Z2CTXzY9CjXYebc8kE3A24uJ/Z
fTlKU4UqwnjW4J4A9xx7g3voiiRA1MtJgQv+3FyyThDgH1/qxY79NRqCJLqNj4qMElQ1xfDmEGE1
sIrSP2mRJDOT++ifwSUFRoJevEAG0qHaoxhiBwDUevIIrc/8VaQvuXL+cmQJ3K7CedyllMfSn+2K
zI3mxcHvNVhLLjPmbxQu/nRueAI9Hy5bj7Enx0Na94ftuj9431bhWT56dSXG2EJdo0d/pyyiH6Qt
LHiAMn1wfvyVRI02lPkA/Q+aRP4XxFCwDTTKchrgIy/uUfv8vG1jkSGT+0YjG/eO4sb3CZFDXNYq
cF59/eczw6vKCVGy/pTOp4KmVbq4JkBnieq6rWjkoRHm6k1EYRx/68U2ToXvkCQb2DGgRf6yiaiC
ZsbbkDod+ciGC/1sFAy4gzGIRw46u0Eemk3Wi+RHAlMAo/1cEXekKPEoc+Gw6JdvhtIInFLw9TVu
BxLCFoWS6Wm5TFhhF+6B4kX/3AAh9y5D5Rs6o/B4mBkiCP/I2fyyy3BbB6YQwk6sLBBDyEiv0Oa9
zltkYwyuT2q8XLi7kNvJdYVmZE2m8e0e0bzXci5+OnNRt3N4K285sKhTZgXWVL6+6UbFHr7ZVim7
1iRORYykBZ5dYtkkUOhebrcrR8Zdi4raVV8I8SBD6Iu4YUsHYy428enbyHVGlwBOO0Q9jAy4FKZI
zfjenFEKvCnmETy3od0m00MV3Q1Y9zqDlk6w7HGPxkLyImdzOJX1PdQ2jCrsjFrigNvyh9yQ+igQ
2a00gxp4H//7XhNj/iBv8ocPyBwb69YnQmNMozKy2ZreBTLihzFNUB401t3LILscvOPDeRHq7vON
bDQzBQsj4Slett92KYjeEh2XfClizjINTrDTnBaG1lIql6ulvAPXtMJ/ingEvLdyyzywn/nnvPPt
SDiD/3tbLCFkZvKfISii0Ousvxlz+tYtygqCnZ6MlEjZaNUESO5L5PTtlUsdpCo1qRdQHW31LtTq
dttTyXcxO+lJLWlOgKT0fOobCBrKZoIsaQLzeb6DYByyWfVbzscPZCNCKyCVGHWZsqLau8pjE3uy
RkbUlq4Ug+Vkd47B59Whr2C0YbVGSJEJFzo8rFTLEODswoO3kPWrk8r5qtjIjaxf+L1cuq8qyNcB
YmaF+VAgl/1luVhei0RwbnsOfzr00OuIRQw7No4SqYudb4zL0tIxyIG38BQ1imcU/itHhXRbLVX5
iY7AccIqaPZYMQMDNgg4KKce76Khw5HDhNTkuW3iRfgvULZvX5uqOlNgeqio0vhiKykfo9X5LZoY
hxHDaJqlDRC1vIVjajdptNBIcMNSt/AzXrycBM3uGBRkaI0i/OpmshcNK37xwwafHR5Lgw8RfY/M
xvG2Ynz/feZ6g4CYDqOK8qPehTktH9uEu1R5upA7jvOEHtn77p7BHx9xQJw7nG30ikSZo1zcoEgI
+IAfbN/tlPqc2GmprUIU5YYhaFyMvPXk86zhZf+fwlH2DRO12P2LX93PzdihHwDEV/ZjUHvwmrJE
n+qi3Umwl/n60qrMbPUBQPxABoPirFGmhWBtYLUGemUkcVXe1O1sAB8YJYK3ZVBdJ2pvRAGipT59
89SET/+pX+gsd/0scQ90tyZeuKmmw8l+FWHrI61lOFbzrA5y7ysAWL2pUVbsByyUhej2fqu3a6FX
uVAt6kzDxxUHAI3ypLTaZzriPr3RG7P90xNznGQtNTLlX1WNcxszG5ouBEMn4NyDW+pt3Ysl1NQ2
q1y86OCb16KydaWvTntcXAYTOIzy20inKprYJhfN1Ob9KsOnDJmKefyAMoD3LKTwZYbikcNV+5Ao
+c2ghNhVrvItSE3KHKqAa9UOqxQwAog65/iQqe+IrMJyzCLvHYoOZ+JdmzU0ILxwjknM7gdTPUuQ
rTv4LcmfVjeI7adwNZCkiOpY7YbGx8ORUY18p1K7WD77PbonuhabNRRpnVb2GgCBhI/MIgtfQddI
c5HZ+7kC1RpddbWXbhk6ffAxqxEhmNuepsnJfGPCYYNy1gwb+9/lD76ZM5OcXyTTxRcnNo6qmpPo
bQPrCzKI2j8xEzGo8icD6KFCZFOiwB1VOgTJGMjUqUkNQU5JC8hp4oT5xWwoxWFZw7I+VnywBhDI
0JAO72PYCjj2LL0h/CjMG/voMjZv1C4jmxCwiH4iqgmCesJwPm4aPcf2yyaxeRt+5cgRXtf6fgka
8vEErMCYHldQpQumlVnNhgzjnoOehfGPvefgYBvxH9NOgwI2+nCpmlhiDREqctTZKwW77Ee0Frid
JDuL1o2PjD6KWGID4OLpsqP6oYMID3d89s//vOgHRnRl6fTGiU9XDkTR8ss5EgwBTUeqQHpZEYdI
BBotoFJbKZvsbgJAIWFsuNLPi+46ZEPS/UH7JqXThylbrK9/KCURwAjnmuHKu5LYCA6rsBXgwC9z
IfdIpKoXUCDX2J1bD6QFgEv7flZwx0610LLGhCxf4Ihh25ecc8DzOLT0+hUczOUNV9VjQgLe2ymK
7GD2fcnK/grsRfwmlJTGVSvTvjgSgOXxISxzfPWg0V8DiAs2SSWMw9q72GVLzJWC6GEDL5Ptufbq
2Zfs6H6WsAIjj6dhe53H+aKNZoYMqgS9dfd+mOLqaHxT3pjp5JAub1BJb+6iHXD0IcKnPGIM5spY
/GCp/jcUt/paSr0vYXeTP4Iyc5/hafjsDzWCShHof6oTP2v/fQA3OeoqrkQ3BNLBTZx/w/MPNXzm
9RzmdHGBCTwk2Tpu3NKRPOJk8YfrdUN6FjwLvQgBMGjvDBQcxwWjZ4OFsn4wqiaM68i10RMsgUMj
2NNT1B1c0DF3B1oX/qCloL0qZZs7iFjlZcCKT/UDSA4Tj9m7erbkiynxka932zALkGlAsIf5aJIO
YLEB0LdDekE/k/OB8msjdyUsv8jNIazhPEkly1V8cLNLPjerazbQ5CKsJQPSEVpvcpeCVUJUG0iW
a4V4aCcnFPOQa/Fcxjabal8eE9WWRIFqWyZu07obxkcf/vvPTBruXHBzwq6n4Q7E205UPECMY/HF
NaKr2vDHe7QGSgdHuKYgj4tV18uPRF1TOXDrXa2br7a6v1OthqfgCo7cVMUUaKBs5KpbqCVoX/Jw
A5ILxtiRx03F8q6qAVvmPOGIggMulnO19RUSuv/ON1y3m6Z91TyDuHHG/lYKGz65em0R2OIXhxNM
OpyAu6V7dC23Uow9dqxS0OKtmrRkcxAJ2otkwq69ySI7P+MAGfs+2zcf267MlPLdolJCEpKrSPa5
ZyZLRkJ58ZXF/ngtaxwmjmiF+qFbU3Y0za/0u3bD8tonJfdGeF4XHpbLcFOagecfPVKbwsWJtoHE
rxdspjMMNECiQBKnskI2nFYdXtWY4f05iSCpIOoIc/rrTeOxB7plXQ2A0mdPl0d3wbckEUrngwg7
RbvjNkFL8Yj9IU++MAOvmORO20+5WNHau7OOrtUta+aNklLJd4y99vKRLr7Jz8g7oO4D90hmDlTv
I/qtDT/cp38V8YMaHOfoHE2jhub783HHATHD7BgUSWYnKhCDK5zQnvpTrYzp85rqp0ACIk/vN7WS
qphVAM850UwG+hSI4y6c55mlfJh5iFR4zc1oz8Ay5V+jOCSUVzlFrFb/dc0XVYlU+B/CEB7iwWhc
ZBNbroBeYysFCwfUjyY5s1Q6xgdUIyxwAUgoyj/DZF1TfbLF9DuT7OuF/K3JK0Fs5GFTpUCHgaxg
2xXlMh7jHS1xDNDwJ/pqECvaPq5bAFpBujoJaCL57eVwHTWn0bvAyoHavyoBa1EK8pjP4QnS+8Ig
I2d40hiPOgz/95JY2LWwPuTMcizS5xl7KeBmEUrAbhD18fquADFme5qMRHLv+a3ItfclBg6YwGg3
VFe3cjZlK5dJSrEMgTu86aNw/cD2/BkyFUDw2oJgnvT5bibiTeV3wMKQIQdvgOY+j5weqk9AOJz0
IQPS/BP2fRKXd0+9/ru01Ivmkkr3JWCsy/RW+U7DdA9GARnTd4km3i1+enxZDcC2k3WjsBfNxSOt
oLYAPHwiF6c9R0nnGfFI7QRyMhKCoH4lXnBwc3jnVnHFKdA1MVmT7bbA9MeDVeypGjrWQpV2a332
KEpHpdWKTnQ1QYQZNYpRA7ebYhzkKhqBE922lkM1VWv0KtLyBk4l674krn3GEZTSy+Swq8FlCw6+
o0tt4ZXOWpL6NOAVL/ulNRi8B0WkLwaAHuhyRbxOy637ZISsnI1n8+RE7hq222EdJO4X8Z0BV9mO
dbx/ZjxwUqJTH4KdGsYBzjyLCf/QKavUnAZzeXJWpuTk68bkGmrHKrRheS1yn0lAA07kc0G/ZVQz
WdA5VCVEX43PzPyyBDiOqgLp16aACu8seqeZNnqDgVOfwDMr9wWR3NaiJ8i39W6166kUrtEBD+Ri
LvWJia51vbU+rvJVp4diC40deB22IZrEZO0UWK15MRI04uvnqu+r58RdXPKsVlB58YqiSPYIsBcT
rezKNXZsxtFX6+nuJaTTMF59XAqiByhiqkaBxWy+24lnV05pNakRWaRxQCyf2XvgJpD/8Pv5wBr2
TP4IKsWFM0YBiTrwMyChFuBk8KHKKHBnFU/eE7cC5SX7bnL6rED3bV1TcBATzlwWlOtdxQD1XA5X
WCVSFtctpJ9514P4/gkU776fwMkcC8Tsfj8kRciLOAifI0KD8btZCw2KpDv0B8vz4jn5z8KkKATl
3VV/7NmRCWMVfrdyinZEUKa9lGJhNhWL9YS6aKdvSUlJiZqJ6rZHEMGCsveDlSFz44+1Q9IXjsTp
V4OAJaGGV3CdnCPirx5l9oV2spXEibX3psrU0xnTGTir8cGzNSFtMwn97cPQiS8l5dwcEvEm4jci
2EkN4A9OdVPr84UX/NnBorf1ySQSqQ1CgR8L4yDegbKylVV2KJ4p9x95I6vNxKEL2DfhaOYsczi3
r1Oq4rSpQnbj2bBYd2pkEPwWjTweB3Sd5sJ2HqL8gKWMIYYA4P3vPucEg6j2E5VIHjJZQ5vpnw2P
p8hQh8zOALXZ0euytw+n7n6jviPhhdp5bKRG5rsbznPCsHHxIb4cY848BLPvDPRb3b3prr2Dx361
m15WCl7mEtRzFm/RTLrNhlqCbap0dFFfIhUnYPrnUij4mFiLHNJpROEfkkgLsdTLO6lgpJh2QaTu
myN3KuZGZw6q/PpbPbK4Yzp5CNJYEMntUGVLpwv4dFcnjT+gtjmxvg6+jbQ30Gs7OzwkBk6rPrcg
nIgVBG4qd5iHyGUIEAsdtQuBrjeURF++dljCeqL4A7JHqmtU0yAlYu0aU6F9XqqYXcgAqzd73WvE
MyR+zEjwAtk2G+Pq1NnmW8PKdmaVeMxj+6ITal95O6hQq46wEu9q93OmnnQummygD3Fvg9lh/I/6
/S+RiU1zMAck6SBg1Q8v9fXWyVabYTXchMyJKLmWlpXR+LfY/nO/wA5JUbqwp3ZOl/4MX8jlbnhD
vbcUZ36YbcN04bwSChtoP+J19oZX817SshrT9+lgReeEnCv1NHklNYSHHmvJD3aQbPmJY7G3tlfG
V6dhklXizMGM4xZzHuFxo80nh8zA3+GcJj52jLfYsTuAmDSGTpLahJdyhDaAWhfc98w8jsbupy5x
IKD7DNrgyyGKshT+g/g1xZ6NsY1LiVIAUodrMH8FIaIKfWiJAFulDmwTIv15Y9IJ/lkP5dKO2uKO
/YVIfgzz3eP7UkN8qHSYJEFK8zK/M2ZJT+cWkQjM/tF5+Yc+pxABuG6Aw6o6SEstZoq7jC++dZcA
mqG2QYajViBtGZyeahsUYAmXSxvK3kk5jS4TFBovdeRcrtYUMgf2ltUo+eRmu5utfIq0wMg2s8rT
8y2Aj5cOJM4/o/iuKUMMsfATFLawr/lDyxnnpUXDn6eRsfryGxmktzo4bOSgxJojH3aMXI2XCFDl
3Lfs03zoDlRTbeCm+Im8zpLnKBdtPEViA+RkECtq1Cwr60ws8Yrz3Ey1ti3+SwSC+ACgszBR3KK0
OfjUcBrD8H91kJes+RNLPUQYnZG93vRzklVdEP6OzqYI/Z53XkzGG7hZBqB7kYq/r5SY4CK0QzOs
XkVvcMrAQgmGIKYSzbgExno25OBLBezGLIYET6cnrvLTfkClYMgiF2DoNiTyAJ+0yt7m20zJS8dr
g2TWtz6CZuoyzxKRQ74kSMhh1JoG2XOuVzGEh15JDXjohNRORHYVdYkeAbEO5Un5qA0K6/WN9iiQ
3iIGOLS5EcIMG+iN3G3aFW9DkcvlxWqA86vTW47ElCx5ecLqihuAfEPL9natRt/O9Mn0St5oB48d
t5zS08NSoxPnyPoUyzJkAT9e5Y3T9hChUuOEy8DoDUoD0OL2HNCs5jabIasZb+DsGfChm8JILaQ3
A/pVuAKZXV90ZgW99z/e8Ytjl0f9WQwDUxw3ngiKrm1Bu2aD1gKemdoX5rWvC4Qs2TuNTuiqOhJI
g0Nvvwbo/9FttGHROB3ctlXp749VBipthVqrX2a2kolSvVYYU306w35vJQqv+wQp1vkk9xUZEkYf
LshnKBgbBPsGG+u8dMtyJJzrEN6OJvQWTjy5BkyMZlLgfIWdu9Yuz85qzLFPNNlr0WWQtW2Gzglw
63YDGC/pvBO6ClPEmVhiGGxLAz6lZKUePMDY9hu6+1QFmzB+a2CTNuhCJIM8DwtJwEyuezliE3iu
JORUtNv3rKZUAmPjkuf9jv+ijBDwmRAzbwWQTVO/iJMVIsOUQZmI/f+12CYNfZmJQDWyp+OW0LI1
ySUFDoyckmn5yHRRO1xMqBCgSpyB00VRRIaSRSVrgyR3rA4rKV1meTzZ0q0VmWA1fjydjOs1DDAn
01fodbYiZLmOGxIVAOJL6EWl9AcRiz0XvANVXiv2IJKrGznpoXw3V2txlZIXKKKsPVGrB3TGGJ/P
bPdKsjpJPybF7+wjWgefQWfKTRWUi1TuSHvV6AQJq/VsGsNJ7OBKogkb4aqXbERum+h1vrBLUQ0p
CDYJizP8ZZ5ti1E8MhQnQXKe9I2K4NrFEg51hMLEWHY1AU2DR/rGEt+VTtmDX/guEboQ6XzbVZDK
bfwDrRb14BjJ1+KbCJl3EpNe7nFZ+8mBhN6E3lnQbP5gHkq0jqwD78zCmlY0bAhTe3jlHuBQrh/D
ZtcihyphJEK1ZzEBYd/LZAQamBP9bP3r9t0PZ1ckdOsKQVHi17JbX5yhny3hhTahV90EY/5CN6qP
JJOkW3J6nXHRxslWUGhf8Tk3jPXK8HblAeKkxpINZAjpIP7uL0d8eGa1rxzoTVFKc/1nUsWuTmdK
uSdnyJwRzq3eOfDZuCg7av27oI7T+9XIofTDlN2HgZohG9pDKOE+LVBa8bGlj9QXdCa0ZaUqczEh
TqXlFNjQmWH9otuVn/97bAIG3KghxcNxcM/Z8Nt8Akq20DwDVz1fsGUmemr8wnwcGsxuKrQnhgnl
htoWFNwcrrDn/RHkHX18gXu+oPQJRJBsWjZytavwxpSjuBR6bPF187zlqz96wqdgRnzFmPRrFvvb
2xQIQuZyZv9kyiUUl8QwzX7N1W4WbaTf2ObjXuGHE2yf9P4ZdGd1nyu+NVI39hbzHOKufGoyQp3K
lmUvMkyZi4ZOe5nZYjOWeUyd5my49bGtYU5NPioZjRxScYeJjol78JtWqDm6NEXwhS1X/rkJ+PAK
W7ApXIR+Zl3KkQttgpL+tIlBo+RdQK41JP2MJC7E4bAcR/2pk2IdYm6fWrmkZycexRfk4ahnciMy
YVxtwDHZOn485Al0Dj3r7sWV3dQ2daAehI5cvayYpasyYj7wq33rKUORo/+pnsYS9Js7kzcp3T1v
4fvHw7DfV8o6qw5aC4VPTJ4rD4dH40V5E4Q5bo+16LLUmcE1JbCySISmwgO8JqZiQ6AMpnPl7H3C
0spRhDqGRJLPcOr9VGZQjL8mhO3HqNUVmYs/vS+gg3XueAf0B5iigXSGfvffiKfF36RWEbtr+6x0
59T0GO2MFJYOmwYN6AH8+gVtue/WBxYNErU4HcxN7SqYEIo5mWICcgi41rQUd4t9Jt4DMvdhsSEo
gblEJj4ehSJwYswEJYxq1TBgfuL5p990OykyCtQIL5YRSIpjox6pAE99CuWwnmFbZmQOjF3fHiSp
zRaPnrdkpJBqqlFj1/ThGntcwroAsz7b3TIe5v/pD4919fCKPKwIKsNVOJHtPD5MxCmJrt+0dJ2A
XWCidjNx2Sn8TulHnhg+ayaBrBXw/pj8nGiophoE+0AjL7NA3GlZ96lEAtAsUt2ayOW07bcRBMiL
3NKFTP1GUtT3GkFR+oqjxJEf9nwqErS4ZHLCRCvzB4z0+l8V30p8Y5YNJWjFXaq8/j/C0enIgl16
X3gwqLpLNqufTXQhqlMnxJEDW3x/iL88qK3FD7b8WryrEeWghEF7t+9gsVrmA0fTj2CIcwGya4LE
SkeI1shSoEvUSzGt22XNPv0ZDClUPBcMHmfOIhGminBrULtind3sWdRyosVrTqkAvQn3AIa8UX5B
1tp/SuJw/jFxgLGixqidVigjgcyd1eJPudXyDKKbaraX9N5EVqpywtDkkxVmygh7vI/dtZ0em9Km
TkPXH1pJzR+1ic4USIwpdQwunvjbrUf9XSCxN/Rv25hlmqikAX18j+0wI5eYPm5aKQV6ryolqd2S
UOivLuqJKRnIvsnnTx/zC1zAdjiRHUMsmQI8AJl+U2Wdnsuzs834pgQnd60ZQ5ZB5wvSOs4j1qX8
qFY9J5+DBCvAsF4UgBpisLnfnS/K2SrOf8f1otjXSzJW5pCj7vgMS8ATYGQH5R/dKsULl7SUWa6m
2wpDnRYgqT0lsdkxsgly1Uz1u2+kBRnb4k65WqUUWAPRegh1E9CQZkZPqBb+7qj5I3Po3oa5mq4O
RF6t+/dybB41lj2Befh52/Y1lzGbU/4qyXIO+Spc5thEE38yj/z4KZTYnz091ZB3PDZ5juX6Hajk
IIT72wsyC9P+3lT7nu0dsdidpV43F8Xo7+bczKYpdaYz4MKcqaY83oAVwTsIh+Khd9uMkUW+p/NT
9pehZpRNdO+dFakjRHlQ2b4tzqMI8bKTYnZvvN04lD4uYZGJxVrdBLTzlrhKzS0Skvj4Oz3ZhKv1
dJSQv0GRpGtLWeqohVt61trkjDbWarxniwm6c3CpsTqOOiNgd0FdLgpZu1NGZROalYDkfmiUeae3
yuElGWQKy9/uwpIVZIYybtX4/Lg19P0mUER3L90BqCVJoHTWKjGLIhLMNpKjaVE0Zx9cxHKN4WN8
f0CZ3HAfKG5XPhDHG01QJdKeBsDN0qmmAT4RTwJQh52Yo3yX0SBMDxAX16Gh+L0x48Vmbs/nB0Dm
rccu6F9tNAA9vem+9lNsMKVDzEXgFLZFnNctKEn1AtuTtZ8UnajVrm399niYYVKQs+jGTBRcIRKY
2sDgIR8ErCHvZJW8gR89SbnUnt9cX4NCKPL+ci7d0CRord3QS2i8WzKngF0nawo4e5mvhsGPhUug
7lr74A+saxSjQg1c7XbHVxbw1/XFZe5igyiayVJplvHZxKny5gT2Vcl7c0zYB2aeTRcN45bPv/yS
Jt5Finxv2A3VXHy6jSiM7yGgqepIIuH/ql0hFC3R6PF1dX2Amk8kb4vEB5BaXLc3gxhYAiHO9o7P
r+YbPLgVNk7F9LSzlBYzErdtFBtZKLH+utMFWGNSSPa9jYYe6Woz7qs3B8OkECDgC+lvyG5d4i18
xjjdvi+ljcJCYawJZwKeDtPLMMH9bWdVrEXDvv8fWC1xSxQTDbAkW3RvjSPGdcjgwLOxNu7rhRwx
rpSD9o2EGiKetfduxKPJOlOOwt4pioQ3gtdpfRjScpuDgIyzxmS/Mhs6+AZShqswMP4o8j3GGKSL
VjUsRqYGbWtKTHtLyFWm641SgU+MumVBraYyZZC20hFcGj4y43Y+ylAhMup4EhtIqCz4nyWhtKXl
+rrDS2kBYEfcZL2n8gHNrcrTtA9SymXwUX3EVrWDy1/ksImcAuRUK8sEe4Now2HhW+cOdibQJG+Y
xQvbnW4ZyHP2qGQYDh/TCbEptXFex9Gyjkd+JeUtux6kyrnCDYSTw3aIkf9OaoUcgNNXIOmXf4aH
F6CjHLiSuRW/Q5XqBXBX9g87HPLzjksvBSGb7/XD2tjWLPucFSYqKYnVSOVyEnl6vZnguU8jShqd
GiSzs+SUjk49Cp518gnwbqRvT/bvuvneQHrGJknQkki8lO8mXJkrc5s+xcnNgwa/gjGfjbntzKMB
4LptDB9gi4Xqc857k6yNVM7tKgHh0+Nmrs8nfylt+SFIalZWHMQwTKvbw/ItBqh2HEagGXQxuDc4
QraEl1HFUmKa/0RevHeb7CxOQJpjz1/bqtOHQwaRCzteiETkGK6+Sa0QZB/E3u+mAxhPqQV8CdYM
V6YCYcLwYodxZC4BULrTl1EqiH7ra013Vov0vJ9CixFVgn3xnkzHI8tekiZzJWppioIfMllFak67
b0xQF81sk7LaJmN2HTVW8G9eZbjbZcTNeSEpRnTQxMyQPECpJe9xWIVz1yF7glco9OKvdb6fFuu/
pbr9BKZ5ZzHbfYb8i9M5ur+qe0L3PItAKnLhkrgWLLTRNUYE7avwqZb9WfRWuoY8/cq++MaeaPRJ
GhIs0XVt6oZt1mG7xNRNurljYCv2AHYJSYH0PsrtIC9TGFjlCmxQ1lbywPJiYVtzi3YDey1KFJ+O
m2/VL6bjUGcuFWFmW4F1VpAhzXWuh8JG5tHldU0KU7mABtmxtaxiiMgVpg+AIXWusHApPiEAzbUJ
qf2RZtQLqnRKopV1ahrU6zhTGoAUcRxaeyMEm97aS+JEznupB0i1SUubsuq1d6vSJ6/gbJFF9Rl0
hGl+LD1mrWZJM05KgttG75/F9G6GZFQcP6mx47JtYrcTjgf5pLpgmVE97hZFlZdCFsfy0V5JTQaB
SLiqrUQKt/m9vFVYNFl9p1Oi5sTOR12wqVi4VpKUGPxJpOtpQVND6ptDklWPExYkM9gGaYoeBfs2
xzA2EL98iO76a91g0YMYfHWZZij/8kEu8hQA1pJrzhSMDZ9hEEWuDIspZvlNmrEKiQbhDti/W377
1FiBc8mAM1GzTHYS/eL8nN67taNrGyG6KOFOSXAtp13oZxvJHTe3q7FfqtSEAiifQXbZwOlmuwE5
21Ot4kmaH/HZHdlAE0/DIAmI0X4oJ03kTebn29gnwSMmM7cgKlVILgDb5iebf5tV3xySvvWb9XQ3
lZM5fT+VmC6rfrXdv5x4y/JnMrzitPrKV3R8HujptmFnoRRLisDJDRGokk2HOPNr/hmQU7PsQKtQ
dBY6I5Rnrdxwg9mbTUX+bLRvrraR9TWkWkQ0y5aGGWO2wymPsrngylP4YOdm9HVzMguR/erTdLfd
8NXLFJaPN61c+rlSG+l6UhGi9NmobaF7Qrjq+2nCFoaap335t1eQvy+y4TEsIHwdw3bAiPbjtwb2
Bivvoqayf0ONsTRoH7H5JiSfjgiiDt1TOu/ixMyX7GLeCuGSYfCR255QRbnaZjjFkNlY6VP6F+yv
2V/12FlOTv4XwlqC5b4s8LI48mLr969/+6KXiT/VkTeJw5ARcO01K8v7grbEQzESGisIjrp3neqF
rngKmzBDhK7pptS9BXOD5XHOKc469tM7b18rsCDlaViXhYbOy2ngatCI2vHlDCsZ5bPsjZNd5U+a
pJ6yXZDbkOqIutx2SkQd1XSEi82wAjgp5klRfq7fAk1xy6K6KVXN+f0wobFRejxagF/cjptCFlWq
VXqJnycv2eciv7RD2sEQUFVolsNy+goekvMvxmmw4w3Wm44/aX7PnYCt9FrbXBguqAIoeq+wJHRM
kaSlE4SPDajbQg7iIIhI3lDtUTirfxRSNE5vBikYhrE1FS22GxTG2OuLiTpX00SMuv6r5gHucflh
z4u7mRuM5My4m/xAIi3662JHcBIj3m6KAN/oQA99tqCnC3k+ykeIgfb+MpcGthiJ82AAPFv28zRn
VeyrL2kyY+qxaOjIdEwo3/n/KsaqJd6Wih8NSfxyc572cPeQ1/GC38GbXxYS9sKw8RTruE9/c+wJ
HwfVT3TThYKmRJVNGlBiZLC3hH0jaQ9HT+oKfQN2+golAEMqcq3om7ntgYDQJwHHh7zxL7MxgXdm
guXpRUIEFffFApXO9zdTYXtOZ/w6VrHz04bKWpjbcprvzZTE1xc7Ql9UFQ6/R3SOByNj+Nisw3vT
KMM20Aj7WQI80UMlwwPMscBNBxVOBZz4GFVp9HHbsmim8msrmdyrErS6EV9jNdl/vjbkTOZ7TyY0
OcDvNDAH7hwD2OJzTWv+Tug8mvP9fLURjVvoUQVZGSCVh7Sq3NijWsuAOorUe4GpLxEiDee4JinD
MyqIGz/KYxzzC8AxLygCXTyHLcxizpaX3ux2tFGU92YEkgfm35uJsil+LCOX+Gi/cfTdY0YiQqdH
b5Oa+LGKHk9Qagl2W24Vzzd/K9+8hxo1k19Y/0T6ueeFjnWsuw8d3GB+kJ8qC8i2GpuWfAGLtMLJ
035SCNut/rdLQjxi/H2UdKGlSyTisZSLjZeblk/l0UjhAn58hgZizhlqrIw0J7hTi8EIpYlq9vtr
qRWRWjjAiSOBt/i/sz2xFsklKM4eXpRrbMqY028aM3Th5jZMwy0xfeuhIvfSPobj7SdP79gljKoS
JweEY2F3UkATZ/639JuAtS6LfBo6FEcl0FA2n9gXne9bTABUKpcLa/8uat3vH1V5aHE67TicqG0h
Kq78MY60MyWMxykqcwWMohBSWGWFcRPUDZ42u0cs0XRJ/dElXzZJCSf2Y2GsKXVNEO5M7cLed20G
h9WX8Lp9UTT/FIm7siNpeb3/HWIRLdvdDh1IBcyOQ9aRBLWfqVvt3TgpWSPTRgVp/sA2DZCSvt2k
VbHOCVieXrxB0fxbk9LB0EhLVoZlzLEXSo59M8CwsmlKLywhDnJYIuusGPGp4nK/aVxZqj1uJRTf
nQfuPoEgSGk2oGpLaiAJpiLUsOQvYeo1E5jGFcOJjvcd4WxP7ZTEIM96TFCqjTRSJBMRWd5Bmtff
umZBjExS3TwnYsS6L69+0UWbO5s9uATYM7PXveyMlOwgBQolleDkwK/QFXfiuokt23Yy4wljnpuY
2bzggl8tZr3CHDhhKQynC7c5oVUD/ZY+Xs/4XxxFjpOhbqDnSB2JLdqsbX1/8nD+RaVEim3HwnTn
rjIf/HFnkp9hAHhJmZ2QtRExssrnkevcMTz/1U1kBocgpCHKnldWhsMNjLMdzVhzCLnFrREVazJU
MA0BL0HwRDVTplMvbr3XmtANRBqWYN6woh2W51iw9bV/bF7LyvqSRE+vHL4k9QHPOL7U7rJzw07a
LebvqtW+2PTrIIV3hLEXxldGhkh9tLurb5jF0/dt27jjSCdrZFPnGv3MGn73GaXAoAxk/F5s40tD
IeSnWezOvlmA2SGqgmlwqnLvBKWeLetL4ShT0lVwP4qsO2D8d+eZUPnG/Qsx5qhfkzyax5AZ61Q3
crDdxgyxRtSoWdfKRvfMuzK6c3O/Utt048ll/+DcCG9FoKc7m+rvKsXXeF1zNmjR/0XfBUr9Myt/
FEahrNRo+qpUYfmmfhC4Ccf548Gfi3Z5zKR9FmY5wfbGq0S0x2qLjAROZRV4rTJQSpcsW+LTFzLw
eqGOX1Wm+kjCekVlszJ8iWcfMsmfNEH2Ped/JsCqdjqsGsXt+PVcFNnvzSdQ9bI9lYpFVNbeBjW4
xqHAwyiuaTyji61xV+0Lqb1g7ReD6OO+Zkpy3OgM+PrmfL4CNBmkCan7ddccii6UfnJIQK9mvGMe
uVKaUPMehEcA0YjR1M8AG4ur+EwkDNi1JIINwuq6jyMGC29dHQ1e0jQ3Yz5FGnPoj23TXabOAt1d
QbiEBqnEsp/9m06F5d0iKS6dU6druU8bjK00aA8Zl2+8jGurxIvgaIBRsJ/vCD8+Wr5UxMIBWdU9
/QG2OiFaJsKQo9GeBiHSUUhaKFONj/GS1C/zHZRwF44upM7laIYHV7HwIE5OHSr0Ar4SDMs3fLXv
KbEcblDb2SPytVRulaRrk6EXgrrqIDJo34EUE0xu5cXf3mKcFNIW2X9M/lA2XNr7ULHAe8JYsBi5
BX3rgUagF0O2XnSF8wMsq7cAfOPYYcGukRUWg6Zs1CkeCV/hL14n53C89w7cMuYMaHlFDGp19XPq
ba8yx2D6tTXB42LYYm7k5cejcF7WgHBFgxrwWRyWEqxKKDZhU9cVUCRg5auE2gMHZTbCRy8xgC1D
i1DZWH6ymNXQxpA4shk/RuxBoOH2KxFGEOTFilD7AyevhLV2GTln4wLW4sLtoXW+UOjC2Ao4d2LS
5/N92lWEXDQSi4/gLqFDGSOeXpsMk5qqdwJZAhIeQ17zhj8//uWKqyz6kCyMF+E3abjMtfRGcDif
pT6AmTkjhqfPExX9Lo/SLtzsKgDoqbJKoaGpEU1tCiT8yEgnZlPEFS7OONjPM9DAwqpX04Iz6s4Q
GHK/bDV3TLMFIhLmeXqS0/OHaf+RFb4FUJzn6MPf9f2jP3mT3hz3rAk2EipdQbrWAqc9oXQyc09q
as7asMh3PCkjFjPHooNcHkqXp18ysJWhEH+pqjbfDKS5LD8yNnYPfW32S8MmAGYmGuNG5Xq+xiY3
iPM7JGcMsFt+zECsP2BANJDgWESlaglbbf9WAdXJTAGPHAfz8lsEeMXGRsPLaKmRO37iHrNUDXDI
0LRpU5tHW6iNZjVWCCHc/+0ABE0HlS511p7Rf6UmZ1XfCQ33myS0Prp6NjYkFmIR6hprg/ZY95co
dObPvH3YFDey3GvJufeaehprY/VwPYBZtjCWvz5MksRE3c6UGv9IShMLTq5sIcNPUPVb3IrMAY2o
Fltc5SJPlF/ITVFsFSbli2uNTNtA2SiPVuMnRZQuXZiK6AdzSHVu+JNbyHFHgyp4RJJ6jkkMhAp/
+MfPq/TCXCpRYqACMBdQpXT931dKAEvLY2aDYJqGKqDBY715pvROklAdrIcFaJ4Q7f/4qkubCy/t
h0jhi/4WG398oRI4/iBaADTpkjKmhRQQsohbw6IXF8llUEwkTS7lWAeFNpxi5iGHrgW+P+oqY0zo
KRQ6t8LqSAcunXKRab8QHAkl5/A380ESaTvo8qfC2PhS5REAV+77TVxi7u8c+f1+fwkbQYrXvN0Y
oLxd2Vf1NFhwkonYSaTpLX7wtM6ecRZ8LfXpIIaafVd3a4Hhqkwj3aJC2w2EpVz14NWgEc30CbbJ
oyD2SY/Bbermo6XheUrP83IQGWa7yk7huCRoTMHry4jEtDPuWgqmSV3snqQPszCiecnGY0uBQIDQ
JfY7cKzTrbeQTDiZMJ5RA0IWaCYOu/sHgUHAJB18AZAj0ARJKoCJ1XRPZRYDdYXJN3x9LEA2ZvAt
aGiGKxmAB6k50uhprMimADzfjfpiTtthdNVWpP6zqPQ8gVsyfjEdwRrw+LtYAz2e+CPKkPMQWzZH
G9c7Efydk4mUoFBkvJ3cORGVTL17eP86a7he2N7sbaZ/j5X4D99zX9SQvkuh3wP0cW146zi7JUV6
vtwcMS35yGaETenOv4xN80+ACRwKw4uiRoiiSIRhbl6Rs+JPdka3bMUIwz7JPhpWd2D7sIVdXpeE
f/4nS5u3anrT+0iF9l0grMCfHYrEDB+0Y/yd9hD+pe+IcQerCveqLPyIZEYwSsUKQ8wZqlFa/qxx
6V/saQhZe4ZCbg0QMqe+yiaiCyQ5PuUWJ0MXcNg5XQf50sbvxregN8HNLJ76tpk1qrUtg0kvvjjq
mG2ODvuZnrbI2zgQnwZnrj4VAxwq2Ol84vp95nHrO9M+ByUxExOXXs34ToqqKIkNmkoXeaIO40f2
BbDEpwtq15nOzbX/wrdt88/uDY4RymwcYC7zaDuE1MxaZYN/I6zJe0aWsPWgzgBCS5Rf7tXuhlpo
HMhnMWKmQD9Vh6rxkw69pbVxLqR4HnE/5Cw5Zzjva00TS3r+mKPd91PUylgOjTxCgS0AeUBut6RV
a2RFvWE4hRittdiGcwkyO0kgEGQ1pZrL9vjnjcNpgRlLp66+CR8YfFU1HoeXFz8eCHFtIWL4xWOT
rQ42HeSR5HrIyZv9wDV1afOS6tvv1SgbZSoP7fySUHDVQp94xzTopqM5UtHyq7HrYsDsXXLXYBfx
y3+QNFzCUo+0SfaRlpa3+zBA/1ZycAQLPehyozu1MdpvXC/kAjBNiNuQHtaplr4B8y0EAYShdSFl
Qc5WSRkFMdxe4p2L7mADH1Z4QaHpfmBdSqqx5ErPxDjxTqchW9RW0nTNEE0kQaktzjCtd7jenZBc
QJCB0XM+OBT8lrhgb7ggrYIBWBpsEyzj3V3aclHdyL1upccTvbwAYfQYQT6Du7V2Q8YWj5dkeV8x
3+9L9aYvjDMG5ZSqSkOVzY4YvWo+ya6hL1dvgsJygzGiir6rogtT/IH/Eahri1erx1QFhG00b0WE
yKOliAiPfP9stiFfXFOijAJAoMIxOjRvys5d18hpeEgOxB6ND9f/xj2Cty/OWJSawCryzxL6UtVx
cPXEuh/kYdVfj0Z8Njw16EGMbur1B+1C6hQyRkwV8ukBwKxwb1TqPJ4rRp1rny4r9Cf+Td3j9UZJ
Q1X/VWDYnQ47o0X7LGLTpteIwPRwX5cCMDe2PI5elxTW040YALh353hvBYnwsq6NsIH4nwrz7Vdu
AlT4M27h/XKW0QhkI2FVw+GiGemjza1NANDOxWqlkxxtJWb6GPfqPZwsJCdMyh02C8yr7MBE8bu5
841uPnA9vKRPBgpgbiDrCEGlzRw/nx5s4OMaii/jomuvQxZK+X4Uckqd0xY1GEdKZLhePPEoDv35
5auhzQZ7TgxZ1w6Gp7W7Umj1aPxBE1JR9sOrnZYX/CnY7LZnxeiE9Bziutx5WCtyhFw8wHFtmz77
HMIvCfDY9/upS1oS6Lmkg2KYHT3kDsl9g65+T6jWi0TfPVC1vARo+yFIRjYshxPysaS+D3EqNpFR
sHVUAeVL6mLS90OCt0ttmDEYKwbIftHJx0WOjL9drfFOzYMzjg/EM2ej80DPt1/cowKMTJMv6Esi
ebL4TjiF0UN2JzpM6HerH2tbM459zriK12bKGL3KEKvbDoLVTDgArCFSBxA2w4FkLZ3bZBLQ33Mb
fdW5XApw2xEuDPhsV32pa3rShe09pM6m772YFi4WxkFKhb3kMvf23R87sTnfjIieFzccjF7PZJZf
1cocTS7hp8mLhX8dUDYLXD/djbsV3gUTNhX3bN1sQTuBdgnH7lAsHK5OPIpo7h+Lke/kE8wOXc7s
3upGOQjG/XvNYUzRiCJdZDoDKk54RazqLZ0Qhv8SU4kRCHiOv73WnLHWyWh8+fAatUIDGuswiCBM
9l6xsQDU+ab0rbwfwlKMIM/NSJg2EtGLU84LFWupgpaqednxFSEAUKINzlTiZZJE9gV8ZYNWzk+a
b1+OmFY021Py6+ebt0TZIBP6NbupqtHhOyJLTEbmGJt1U0er7eHOspnpPHZrJrogDzdHED0PtFoj
tqVwvHZIsKAKS/HVfEBDsOgKxlYjuoze+fMpQ4o9ZWSuaVgQV5BtOAikohitMgVGxotXmcSAXpsF
6MGX7fN6dUIyca3NkPI1qYDrsBnGsiFoxSjeVV/PetJRLhVqCXtdJfFi6Femd+JFAcOc8QladDdf
dHInm24t3mWFzgXyeDzzhFwyXKNQNq5OVi9kPIK3mefoSwKOBWyKOH10E7UI2p3HlYiEBJ5m3Hla
ZwCXeS6vyCJe/lj9SM2KNBnQu8DZ5CjVgjDaxKUJ1NsCCRqPZgtsyoouvtA+8XZxADLq/yS6zyKZ
+krfRd7Zi5Ym/hhfVWVAl0Zbr7NYKcBTgaTZmCqaeLstGxiECIoS6KPmA7OgOIje5Szw2L7Gzsm6
kh7rbdwv2oXOYBVjJaLpgQ46g1+0rsTGAKDr3gP0emLlXW2HJALq6rjZKpxACELBQG3DuGhNDZYD
8eU2FqS8L+39ocPO/QWrRNhqXbwDkfZrqNFX/AfJ/KIHsWwmSiZpZ7ndmUWCIS9dTQ25OymTshXf
GmoNq+D2e0EehRmWmIxZU+H9KUgkBO4s+NAhjhCA3ApX+fuqjfSfq3BWIt3ZdY6kgzWtZKNmpVNO
U7fzbaWr/WG1Jadlw6LtI+dmZJinXb+uS/1BtEZ15u+hWQfVhRpR1uFQwyXslMsBbLJCusU1cpZ9
KCqhyEN1DSTXbp+dYEphi7a1KuXc7FtZPHLm621yvXi6f5GDgcm5UcezOkpRhtf2XxGpZY9nLVEQ
buNm2O8XQbk9uG6Um9OA2pnTr3xHBuHsMK+ssCeEKEJfvpZB5S4xtfQJBbbMDM3+xYaJyyu65uGR
TjuJYFVClLrrQn0/KQTfqc3fTOVI1qGvCD7ZfNqT8NdNjamHGUxJq7BpUD0Ph6jLsoLKhYwryoB5
itysVVn40ubC3kg+0zjjdZLnIft1tHW6LmqKoyEric/pzbreRz1OMsZfsJ6a6pBNOsuRABObO7Xs
IlRa81aGF+nSRb5Pave+j8ZspURaFK09XaKeHF5bXOOc5U5Rs7+uk62qorNsYDYZfF5Zn/yurvZh
Kg+0zuN0t94FeekO7dABL/1n9dinKnE4+gXGVD7TRJo9XUe6cF5HWO2plESA2vGXyjkWG9xvSrjW
+lXHqDv69MMJAqiXI6T5tcWSBFhRY6fLKkoZYZghtImv/0PY6zyhqXoFts2a/kjk+kBaQuB/94kq
u4DYwbh2JKwmLnR/S+afHPFaz8SfOMc3hNEK65qsslj80DcYOpYdxpLHnlB6s3qcR08QM/A/IQja
ctizI7fgPZLUVJIrPpqdxBwfrmCpBpXDswUc1L+aoX8bitnRA3b/De33AVEty5y2ZwqdogxQrWsl
HCsge9IPXhctyILUpcWqGuzO4c7e/Ui6JWcVZVYZapQ5YL9eP5cE+4EtZo1WZqdUMC+Qie3+uN9v
nxRh3mePBLvKEwbj1ZYuBbAaLeekNQ9L/Ffj/9ak+F3QYBMoQUL6YzVuJnbf762LhbS4ZNSf44Yi
fNL6PesQjeNBxa3NodCVevj/yElTRJJUnYhUkViskiK6pEQokVUJ6ihinj9N8tYudVycaHPy1Smd
cWkfyGXtBT5mxJuyo5pqOXSLToX0/UyiUMk6c2wQ2MQ+T4bsnKP9Du0FU6t5NJ3rYAJWgiEe/rjK
UNDLZvH216IuHbF+XixkOhBMC3Y4IbSGBIqB1Dc3hhmbsL6iC2vh9kZZye2o5aF7tU3agOZuGWRS
fbfQMpNMUOJPG3xjO/AbrVWOxB66oMhUjMPGXApt7wTp+fHU8iA5r07Ebhoo/v+hdax3AKsITDYc
FG0svAdnSm7ahX0EiHlwULU3FepqD3ONqDxAkxf3VtZOW7v/YW5m71QXO22CtsnKBYsB+4412unx
jPJ47qWIxw8JBWLs6RGMZh4BuBg16/uUNILYAaGgI2DPf1c/RoRPIMu9fvtW66LG6hY2X6lerJ0j
JDb4KtwGMfxOMccWu0mQ4clGDiFcvE6V5v9IfGR3KD6S1x8Tj2sIWzIMWmJyKOyYQMYcZQKKq32t
aemkDjwgSq9R8fwmj8m/ffJpZskTvRFRkmCm49KsJQwCsbZwT5c9Hcj1fjg6KV+y2Qy3G2kePBrG
dQJyJtKSv9UVuSgOIcqrAzU5cTavnzb9eWbiib190kG1fKE/lVQIaqHwcxy3Qb1rR/WsmQ+3XsiI
/9Wnb0HPPSZZGcpvzv0V3sR+qCUShkKjoyrRzr7CmySCsOoTPL5kQij/UqbavwZslydHM5zh5AG4
qBQ665oQ+nFvo8kiaZlorpDqh5f4syCre58x6i1df3DMwJ1IsVwPdyW06G44MOYx1QCaBSgUa7pg
RmXNnWhfKimLlBvoTb3LiN1+O+vK1xSQYKspqXcn0ww6VX1zkSykrz7E5NGxtMJNcZmAT4nKUA0r
HF4V3U1UEvENwdb19AB7kRPvZ8coV1gkejr1YNjeHf5Wka5Q2iws4vf+pTeAfbO370lstH8QdICh
Yd7OgsnOkm7pfC+KdwPshqxTkIQDW2UBEe3esqf8+jOBzq6bV0WpdXskzYCZYfZmcYyix3fGz2sl
PzQdas7GA+iFdu7wZM4T7/b0VbGePxY+D7BuVCiAAm+VrhhLXTNXf1CBzWzaDbgxfirJQFk9FoSJ
3Be0pqUZCAAMkksqhGwPkTIYTbi0C39W20RW0mkPuS0UWfheP9dnlg0y1u8QjEIHOhFmJP4SQ0bi
GcSGTe9lpeIbk55VerCTtTVFYIkNZY+ZmY4ZG9M0RewkS4satZR7jUp9tjsmemqWfmZdqrH/7K6R
H9zetwpbzxvuHO8tcMEdKSqoC8b8zqErFLJHevJKgIU9XIEZNRWalMexULAh1O/CK+ArC/t1p+nu
RH2Wxl79O9aqdH3lCrd8Nke4DarojjY+UpliOAMZjdMZ9qHbLOcqSS2AJF54IQEdE4w+eN6v2RK5
Wzd+HyTjqruDQh7GPaDZTTvxmMUk0eBRZA3AoBTLE5YscTo2Ud6ksCGErpxSd8CFwT31rlBCenAz
gqDGuJ1rIuu8nwXy066XIgRbojMJjq8AB/T8gQIoFYi0VNmCyWUhbOcV9xK8QkpZMkzZL3xLk2nz
QB4FyQm4ufx3KkzsCT8LgI1yNIuA7ESSt3pO0EXMjmhHWDaaTLcHCYyS957h9qWBCfrtzmsw7uI2
cFCzxKE4MC5LfPtPEfWAC9/F+IAd0TH0MUR2yLsvBgtX71zfrVI2YhpShHMPsQuC5haQDUzn/C/k
W7wDiKyoLwaRKDMsN7mv5P7gaPF22NogRSxex2NzWr8y/eIQEuR6wsYXhcahQjtSnQPgFlWsgWKy
1gD/rSCoqkgffxHTqxoMYGkhdtpevKA3nahq/r/F715DWH2HY/6fkju8BS8U2zXTKYJCBY90C9E7
vdCIcNI/r0w9YXLxEt7FzoF61BGya+aJ15+lLgVVKZjL4T4ybC0inmwV9OuoW6NJ3refLsZNxsKv
5c7QhPEIvN9PZklI/6q4J5hdF3bEpPH3pOtDuwZyx5aFdu1Ltmh8EfvU0lJ4Uk0xzBoa4GfqAtgz
/wBFlBUmL1iJDcIPRlWoy19DfUcxWmHSZVzxyvq4RDYbNBoibd/lAEFUJyL4fs0621bWC5BVkO/B
zBqPLXo8Rxzmi7A2M2uY7ClnwjW+jzmm1T2qR98W0o+qXf8j/nOD0r/+z2FAsmyoo1v2ZXvwDIRf
5oX/uyMYvoNve+dGyHFr5KVLVjZDpghgVyIQW4hUUu57H/Pdw+TvGJbAVR9jSqfMFG1vJ9y1dwjy
todsT8w5AoOKQVgoyMfPWRXINCipVP1xo4dyhd8hPjJftSmWgjOqTRaibAJh2iOH/EJ++en/p/0z
OeV9N+aQhijlVojPTSY3uJKhTQmFg7SOdU2+RCuiwKsw0wJWdjYLWR56ArMrZUQ0NO4fx8e1M51S
pXFAFEf2UljHSb10ThjVU18Y7thEZ8ZFyu7tNFHvvv/AKcL6X0u0sXBvHxjT1Xn045mIRlHbaiM6
Nvkg4BoPbAGOtMyayp5wNPOeUP9R/s8y0WZ1lYnLdEJi/9aM19i4Mcc6RRVwGFpMXPxUA1HyByMU
/EkUGWNm8W0ssAf1bL7Q4HMQXQTNiO2iDEozsPTEGTWQ1pndSi2BWu26vGSTFWVfT7uv3G0PoD7K
kDVx8Mw2govOnfTm2FpyUJnNdJGGy7mz+jORi47yUfS7NZt9ipMG/fKZ25oPqU7fog8WABg4ntg8
j6klkAsCvGAIlECnHElJnwZwW8dWy/5ioZG2Q30MI3YHVyYvhs9YVQaYCsTUYAqxaqgu6iXw+vws
VXh2WapDRIgxnscSJ4X0yVTFZ1VWVIj3IlixdKcumcL/rLgxKLPKMKz7mGf9jeEv+wXQivN2h6HM
FjlCiinJtncQajSRsUQZUvDVbCA/jI8K7DwZ2FBjg7nXHoI3bx1rnS6qISpOP4Y4EcQyevc5ceIt
YHQ+OK3S38+/HMZWONK158i2fTsmlZZ7QxRZGh7opuCZZte1vno25TGa2fg1fqmlXnYveTLvrHYK
2WG7nowak7HWBDm88F319IqXkiQuPLeZb+BlDC8BroPF8fTK3JAoyC34gVo2+Gy1Vy5E6TDvWrGy
M1XtGM+TIXbOHSi2qcBMCSPJioB0s4WzO/i0/sosYucOEMn+I8QOF7z2cHAJmoPtoreeig1sTjNx
UMzNcmM1bYRhx1L2gEC2/vuNtp7XKbPZDy6jS0UIznNVSaUBYaFdRkTE3EpuQThDVUAadYoddZNE
OmhbyYAQLslRoUCJjIr+FA7JnkMvLuDOJMPrt5DayaPw/snIHB4X+RoQGo+uzXsnif7BP0Fmd/6Q
gsEuXpNacDU50FyPnzxlCgMSOpWq0CGldj3+FgLJ6qBCZM3LbVOh+ibKU5ThtR9l3XwJhTYz/xbP
ZIr0n+6+ynRXf3gc5ZCzRdjcK+/C3a7/8ehi8YE7rXFcCCeVBD4Eq2y88ja9q5Cs5EW4vZrLnUeN
XORVxTHWVihGQTuKiGHPQBCjuR0Ke00N2GEkKkms324EoR7ILk6C4E+DiSXh4+NIZOkdiHtmh4bo
mjvtlkJHOEjPiSML9heNmNTNhx/femyG54MMChnpWpGmGll3ZL9ojQ+q0z2//iJSYnKglKtnmyjQ
Hiu68MbBBn1XGcxN1iSlI15vhG8PgQbJ/t2a1r21/KRz1ZMqa98NphJhrY22LnS44WER+UOPOOBs
4+XmHv7HSKrT5Cg+k48XpXvP/9VWyn8FLOLslYA7bh4SF3Iq0/n6e+UlOVYU5kjEQG5BQsu1P4Tk
UV6bj3zgOdGjU7baoZmXrZW2fPwQNXm3Gc/lvdXFNgCXTNTtZBkvYYdN/rwfMoiQaUvleN4xRfVe
WPtM2uk2t9VUyA7I2hf0KXdhTGEcGRn5sfrIoHtvasHfbTtT2UFOyupv3jzbcPJU+0sCab1tHQIL
1Bv5kOefRodo6sMX6fb3bE2+VifgeotTS7CqoIGaxPdJzOqzAci01jbo2X3t0kEc/2canCYF3yK9
iUL9umpuW80nNqizSYrOlv12Yqaoe1aECqNU+g8Y9E0XSOuvhRKuiQdUMRVRL74Pkynd78S4BSzE
ohaAMGHT0ngFLJUaG5xAOWzlnJuV09VZ+Gpw2R1obi7vdRvodlg5fezPWbxnalh6ajEUVD4V/klx
RxeOWBa0zKmlOtGnv//S2hA52YFRbebxrXp7QBVdAqWJ9ghpOiMDpNSWl+D5DHGE8pgTnUjtuO3v
XCtAqAdOSvjShnnQG5vf/cT5NvhrHGpGwPk6vdXyhirNRDBkN32iQonkDIHcIjRTwL70khwPEudM
BYzS/5PwflxB2wejQTubxAUXIxcWr/g3pQczZO0oEv1hQaCqtneT7lPWKnj/WnCzZ4lPwu+s6SSS
0NqjQTHUr5Bo2gq2Sh+nZpolI8Q7AgI67efFVUog2Gg6wZc93olWMxNgmZfGK+PgfnfDHfFNlj8D
y9DcoAYk7WBVNnqoj1Zvo62aXNMcwRSrAgzW+3H/2Ip+0fbmgKa8JcxF3DEiAMpVQmh1y1fyES2G
W3jpJaEUkNHHp+fXw4lqGPr82vYaVkdl0Yq+49/dQGxHN0V2Sx5v+8b9gPFcbrKLJOmO5/D9M8yx
bFDxxeWAirgOJUdWKs1gkcKJk1P/aV3nMFvIFtoOHwdJkhiAGifpjL5t7JUUuUWWQuoBieHvuEsR
xz6I9aTkMRQ3uqe5DkO6Dce//BuKPDxGyH6N7HEExxI569IDn/TWeRZId6pxL018bec9jqMEaZAN
5Ld1h1kpJhWtNCh7n8u5mlgnh6aBRwNrrmJdMLdXOSwChluwm2PYjJm1Y27PVWVagJXKSrA/YMcy
qZh7I8tMmnQ4aJRzQHhmA0IkjIGdHMWLWWr5pHTADOQ9ltckvgkCIKrQQrX2zoXkTONunlQUr01i
/8hzRUWLC83WO6pjWUS2C15gpf48E+n5+TDwTyoXAWEifY67HW003JyAej0PmAOcB3aeaBOhnbcI
NEIEos5e/fZd67Jr07UNJaj8BmNWg49SKNVscTc9zybG+ETslMOXNxQyFqJay8TigOK5ykbyiOZv
CK65+zqnFp0KsT0Q+JIq+Q7VWwrOvkNN9YaE3VHpUgrYWEARV8Bg0/xq73Opk4XJ1YLtdsXu14A1
ET7yIsrMA1v+RcErSuqhybUmz5OyGS7i64pjtzUH/HDfRqqiY79yOs6KkQWiY8A4LqWCrpfHBlXx
wudfgTva6r+haVlqHY2thinbAp8p6UuAEW+v/UXKS6TFM9v6MvKZtRzvKkjQW+hWS0ErA+JsfBgi
QIoyMiVmnryPCv3l4w3M7WqOt9W/vtU8pd3u4rNksOwyE88ZD2yLEmL92RN8NzyKqdK6CMJxtV/8
ZaBSzr5oBEAh3F6YnCAo3mUXBSMSlsNfPduJXqpV+QnZKpgp/20qQ06+QrLXlhJml4q7fscLoEmr
h1hcmJGEGBBpLuNm75oUWnwixfjJPJKGpPz9piSTr9xP1dPwF+X2NuE6Kmib8LrkXFYvfJWEyGhk
3CAdLzOz97GI6inYdFt5I6j0246IilJWuQhpTXNv5Vzu9dfEKbbUwIl6KKe1anNxTeN5CiHNKwkS
zAFfRPWhn+IAF6N4GamBNzY0Ekzz2+T6cBVaOE+ZS+9VlUSqriDevO8eW40AfvbsYmVGBjleLKB7
s0FhTlURMcyK0H0TbNtYYqQseFVBBU/DRdc10aTTvW9/AINOEx4O/0yGYjwcgJnNKizfWitOIULA
PKr92CyZ6a8oRW3ii6k5MIbfyANAjYv17pPZlptjBfB558E1j2KUrJ3coeQsvWvTgxXbQoZjLrD1
XkfQfXY9YRQYnkwBVMCwPnkf2irVRZILonf03zfEwE5WF7ek0kSmfcgnHroeVICCRaDDC3/uwoxe
LNIw/PFdPkXuVHxc+1s+9CVOIYeiJdO7G3VAYbMN1ZV4FhQdr2tmzIkGi3mRcjD7Ii4ucsa+/8oq
JijC1JEENGJXGPWxQpZpIa62DCMl3wQPRUMOoqU+BLkUfkx4y28a+bigk4ndsZlQaHLOO1DWxnp/
ZAVDN5Pbh3NdgM6yz3xFT50uJuMoOZAz5sFi9+h/Dst45TMlCuNvIF1oPq1et48OJziJmIh4KnL0
8YFd15T4OexjNfbXGw7POUnkHoT/WgzbTsu3IDn78Tfm7kcIMSKBNFAeaaKBwJ0mJY/NLrdqGPOz
w8NyqcOvvm0YsrG8YhlEKRXF8/9P9L9sGWMyi8IPvhP5ARCJB4U+Nd/Z2KB7tNo4GIyKEjSbTjTW
Cr7HUPP8AHjv76aEqazY2rPB2EAFtdhtsiG/BqRqWHygdjqRPLnhk5ol8airKjO4HuaiEMJE2w1L
LhvizTjYwMNaEyqQ9cWDOwpz+kgVRBhdZD/UIKDjfAN9RCH14MR2wmTKqATihxOhE7wALirzF+md
I+QwCPNnnrRyyc6pe1M7k4qwDsRiVRTsq01g77FVWDEIabit7jgPMssvkIKpPxgwLTLWzCV4CMZl
fMRyM+0ECyPkWpTerVWhhUpH1qVuLK63Ts4b5UnvbsnSeR8KdPYOfqu1JrsZv8KuoWKa6AmZwrzJ
VKMizYSrHl9i6E1sMjpNYC0mo2Ec0qucjKENHqse1/F16rd8UA7EQ+vVPbJupxJytP7W44xBijq2
jDWkOeUnlobud9DLs4nDnUvhC6zd4AZP24szHuimqrk3uBClql8BJsD8IB/tkEYgmXKHxvxByafw
GKB+5b/8jLAXjh53NGfAGh40ZSDdJn0j+zM/LOHFOqC1mFHqf2kkgxwT5esWNrNCkjpXfLb4Ul89
e6wjX7sHv/j33AKX/rX1UmHQxekYgIRFji1tX0NxT34Q6B09ZHUGMKUJ7m4Jhlb2EEN0dkcHhK5I
4sHkm5YzzKNsBJbLZzaVpgVOBdLqpG10b/iBhsmQqSxQfET86D3HdbrGd4hJLmTpmxBYlXV5A+D+
70eMuB8p8RwN17zLt5Jo6knz0X82jP5k+vBoc6OWP737i1rKyCHB4vW0kxNZRtkgpFMZenucqTfm
nKifsUEunJTieGu46c6vQBjrK7BYCzOtcSfbRtwNkCtMVcbUOllbJICJDswR5Lgwy04rFHVRhRI+
UEQ5e5zlIPJ+wNJwPEOOs6Olq+krSFTwDjTzS2T29XGSZxAjIv6X+XirSh0MtPwJBT2+RRFjpDU9
CMtdtWxYI0FX20IZRYN3ubbHKU0zz8EDIFhxDOwZaL5anHXtr+pyK8GTuldpoCWDDh8RoUj46aNb
LyRO4QPqHy15V0L7hFjB0DLLm2qqFhLALmk2gXtAsY9UPkYlEgAnhHrghK/1kSaB/H92CCKIWeCQ
lCQ00sGT5BU/FeGFoTn4+jogQ3K0Or0MSmyaD64TX1Gs/5xhtA3l6hr+YEorxseboV2e5sc7NdyU
sFWO1bBmyDg9tozsEVti2l6X0xChZVgakaP3CfdBvdBcpRrcbpdx0rPzsc0TyjXmjrCMsbFOy53/
0uBoTPuP0P6mU9flZObJcTx22eMcqYyXnG3+fDqHarfgi8L8VlrehMhJCm7jQtRx5GpKvbKpn0wf
EfOe01o5Nj8nnGAvUNk8owjYJXEeBxwBwOeGOMFGZYGxtSHVbFJNEBcUdmEuq+wQGyGdQj1iJemj
4PxRM0ftu66rEPWbmj1DYsUWrW0kgIHHVR6LHh85mMFujzErtWsNt4gbTRoZ0tZXVD46DBBdjbZO
i+x+Yto8LqO2l3vap4qHoMHLnPu2OGJTbK8Lzl1hUkaKHeYMRp1Rt017GgSeSl4VWTCJNEqUgxZ/
XEWjf0zcKh+Usw4EMnMyzZbSDWvhY/Ie6TX8mUOWgKME13S3wvBol/x0ETQH9bs1OQfzk5ptvtVR
1ZB4NGELJ6mTg4OsxmCjp065WMo/kjtWEMiUg3/ND0sfrXudpQy9AiqvEBUbE43WO/RTN5jAxGDP
K9Pr15fMfVFeHj4NlhEFkz9yko75YWB6DNVm+zM+LaNZL1f2TyPwBguYqsShyWcm/1X9Er/9zvc8
PElTm8g4I5k1inSktqu6rZ53rK4RRSQmZzzUyZdWaz5Yje5khCMvSv8bbMeeHWq7qUxNFp3RNbOd
1sirGVONCKmhwjzX1Un7DkVK7bB4YybG52L5jIfOCzp/8qZyVj+Xwl7QwL6hFdju89CCVWdPcAAY
jqIz9kGSdV9AiV7HmbBcsA1Ih9SEfuokZ34gttpN2wa8Nl+09pcMBef92cRFfh9xbYiPG/Jfew8P
TvLuUUYMR1mqZ0sO+zbuNv8Zh6hjdMJfePQvb8l2jh5vTbSJKd+MQm0WWggU8X573c8xDiHArnIX
fP91risArUmg5581EyRLI9kflTi44DRlASLl2pD/pUhgBpfMy0A0gKtgGRJCEfqbYSH8+MsJQPMm
XdYtia8N3jvuhT5Ld/7cZxBzn/SuCRWuAZ0JhPi5zAM64A5jCor5dhbGQXpCk1GKbZBadrv+7IeA
1x9rogeAi2MfoBYvgvw6f5ac3FaQCxW0bokYG8CsN+388xtN+6B4beVWk2CENKyfVIk5JF5flZsN
cUWSUEL/9vupfj2VK2qY5Wv32TBcHQtQfK3J+Y3US0AtTCKYBokb6MiYr/fSmc56SPb/CvHwCJXb
8g0JG1sXnVcyx4sYFPmHF4ZG3tc0xpu0wYp0Tf+HDkwLg51yaRJq7coAJwy4RSkIjMWtj2vtYdRe
TLBWy+fBOIXtKIQsSu/nzg/Pqe3AiXAjsYFdhphGxIZieS/N3QzVRsQStVKX3kZ3KsZ3eTVlDOnc
jsUlMAcrlrTdCoFhhSsTM0gh6W901JA4x7xZWbCAPFCeT6x3RBbuYmlDi655I8lizgjpQMfJDRXH
N/pPlbqbJ/AOnaaL+26illjnbE6NAKY88+0kLuOk5zmqkVJhNlTHbfvFSFWbdqCOanxxlqOq3RFf
me3YxRIoPbPFAsVwJWocmEvCNglBg2cNDiUwg0UDKJ7FJ58eLLjiuUFDmLWmjfrqeWBM6jtN9Uzo
eMHe+6FIj5fy2Bo6eS9kLka80Ia0khdsv0/k58o6poxouuy2pHdmkdVu0ETteUD36zNbd4OR+GF0
QKC/JYx8H+mVjeqzgr0HOeZSDk+a9UyYV3mVKLMeSQjog3xJo8LqoKWPK1VyREeHuqrOP/a5VYE2
NSvdtJuHWP0EZFYoYJIdDPnNLMHK2+tiaXLJRJwL0lhv5ZqbEvuTXtBBLtq9KQDQ2oZAR/sdF8TG
Dr38foDDws9iiU7pT8+Ee84fSXDjbNFocIdv/P06zbgIKrdCuoYMATVOnvZ1JzkKiNrES+HzJKBp
d3NcB7P0NCwAAI8BROMS9dSxO20ED9zMzzUbNCWDR1PFejZnVis7NNAi9tWtASbAyC1oHEYe/smf
wWCLrAW113VhgbGz5PXZC1oA6zNrUd+7HnCpc2v32CvX5hH0nPebLgmIGfr4Ezjk/1QB/9BQTI+P
vH7z9e6wXkhQHnYZFHBSqOs9P+SnZ0TrVVTqZDxoM7ki9mYJUktdOF44zepwv8bsd2zyi0tSZ+o6
q14cd5PXY2SXN7pMRQL4RHnOpjEMmTru1+Vu81dEqJUJLjxDXJ2fY8dyNTEkkSFr3vgmSF6rfQfr
OAwGQW2XYmI3eTikPMOmyvYgV6F6sI/9zdq+wEdnNnpmVDpR9EcFAZfQykGghTmKL4ONczIAn+AN
NZg65XrvtXyDhw0qJDHXOJ8n2luUdwGGhNsc9aX3Gmxguyo2JNaDgbskeWWNk2uEqjN1At3DCyJN
qYUaNjU5xHhxW2xS5YgTa+9BxbEJnD9b7q5tc7/wcqWOSfNc2iLySsa+jAo5+8grfPj5zYbvKq8Y
JvWbe4ctiKLnPdLJvbkdMILs0K84ewkJvNjPjM7oRN8yW4yOqYkoBZKmFZpR5kxBw7DPYKfQ8T0o
+2jfNc2MuK70kFmLFGcOOXN7klyqFHht+24ZPv2j2eu6DEebUA23OuUEHn+7LX6trhdsPMM84b3e
cWyGlUlx7PnNJpo4wHjTosS4iBwpTce3IEndweQ4B5wbqeH4Wtyr54aB5ICo8ObBW9rExEYixOim
SszccxHOSkb36k+BNvu+XOQvPjEYgliWsCcmKdUjBRVzvLa9Q3j/tlV7WXKk/kGt6mvnTIHHOAZl
lR6OXPFHeZnvvmWeXYIOGp7J2b1NhXHNfT2cgqKE6oMFGI0hnS6DeTkWrqUvOVmfFZcUBZzofAum
PjFdsHlNF8AqW9Ob0yo+wW4WZ9jhFBQ9Zw+6y/r19Br8171PQRwa4D9R5yjorXGo1pKqbOKMfKz5
Q+l+2w322NhS25UGqd8S+PdxpeYRccJnA2TKwXKEHVq0Ft6GiI+X0ciyPEM/546HaEsgvHI8An2U
8CfJ1Sx7rxNg54bPnv0yHKuT4NCuaFq5wgb9R6e1EPF8TB5EJC54D3QvPAcVC8v+88uynkNpckk7
7tWWQR1ixvk4rXLXLRcKIE4ACGFpjHoEYdEivQlxY+pq/aw8bKZxUkxUbRQnCw7rq0aQ4khtMD+C
pm+1NBTQAYZ/D/I4WOPPjit5bG5PoEDBhKOCGeLvweWZRzVffYYBXFAeqQ/sp9tfODTpK1NExG+1
osLJeZU+pivNcK9jcXhx/3A2f90H2Mx/q0n7e9I1V61QBWCYW+sKMzprJoDPMlIxiP9lBvKU4tBL
QDnHKxGVJJ2PLGYZmW/TeS+Vm2XAIUBwpnhz6s9vza8Rav5yZHvSWJOLbPFygz035xmW0+qekawq
Lpy2mu2Mpx4nE5M9txsMYgOm2RQ2iwnBfLntNhG7gC5BrdWWAx0cYXeNXDBpUAfrQKNwRLIh6xbo
ngoB4CQwYAoQHOMoQuiarjON8wciKsRUu28uMZKA9C4IX8y049AUdEPAZQ1ZiAWtxcgcAQrokaN4
MM3Qp/Ij8r/r+10K6SU6qd959Ek71QqKjjwU8+v3q1ih3DzLlYwIlkAn6IWqux/p824Nq8dce/aC
OLEYB3TODckTkEAxCiUZzumirgXmCbaUXCwzy6iFkz2OL0GlcXJpgNA4xkTbN21lneT5nX4iakTw
8sEzxZWXrhqqTUfvsrwqUCxSedWmJ3jy01ixKPsbiW4OjmdVfMbbHT8B4kZiYMGsV97QCaVOt8xs
gDEwsEVx6BAXDmB95Hppb6230h6HUmXImfPj3AGRH3oVvuOYUCXXFfBFeYXVTvWrmZrgfDsA2qDh
GDBo+Lw2dYTCK6BAT/jhZe7H5tK4VsAU9RQCAAM5/8P1+C3m3K1xP+PRzBczzzW4hGMviDmynS7q
+sOzZjgjczbM60bGqmlefi+Pzt1+U0wpz3bwKUGa1t34TeLvTZbbDB39cljUE8iutBKpItPs8zoC
zCJZ+9YXMCVfid+iLz9GVRBxXm0zHrlaJB5mf3FTYD51KBCwVDnF+aTNi3rtAlFSjtJ3wEaMbHB5
wT0aaOmsDrTpP56lVnLhySJJ8cFR9MunyPXscxV+VxZ/m2UCwZ7lC0ojMNSze3mxVMdUXdzAG4Gw
KNwBe4h0pXdzr6+gmYtNQNUCg77CgkFoscYRfmbsi0HNCI0zoC5F3lWLss0vUxHDxAGzgR0VQoPQ
grWselVkwf5kYmxk3ffuHQb/UUKRPLlWtOhSYsKLAlsuHU5nsy6Xb6CppWBiy3rNeBdZOwOdIDTv
DuLOiMi0ia8iqE233KUDjnAj6Q2tpIVLkE7zucnp3L9TPLdWb7NKw90mvWEtVXSq/6ib/qRMPT3I
cb6jeRw+cWiPMMqFBsJGzaUNUoKYFM0DZS75FhDTvna/PXn+JdfQ91iJYW5L3+TgfIooxHMv4sZ1
CN7RqgDhdH5ijKLC4Fo6+974v+2MuNjEuhhGSSiJwFyILuA3TnyocH6QAE/4L6JxllkR+ccx+eTP
O1QcgbcnWoXbp6SmMKIn2t9dZABUUd0HizLuScdRfQMHx8KR/Z6650BKAmLE0sqAxxaYM/4oVJkC
vkeGTsHqP9AT4QLp6jAPmVoOS3NOZieD14BGv946PyJiS6tCc3vKRQQ3/m4Be8iaIJgOm0u9iXDn
Kvl8mh/RK8S+g+dfdaPaOYljWBiCSfDpP9esWezjzOA3O43Bu0xywc/jZyuRm8OhmE6k7rLtuP0H
3EeL2yvJafFqn+arU27hAxnZa2WLjEMEtnCP+ax2AA93Tgez3scbfxtgg2leXOX8IXPempWJSN6V
P47RrGdMEDXDNKyx0s38Fa7Q3eK88jmFGMxfpcSKwWfufI8ZU/b/l8F2g6l5SJOc9tlsYuF98OYB
XcdqJDxfhGIPIapLR9oJIpU2z8+NfGAFplWaqsqkmPAgDC9xsaCJkj/VzsptP8IPavzQwjLD5xxp
vVDo2TvB9E/XVOh32GBdRh8PnUgtnZOR58KXTaCEELVP5OD28W9EW5vYmWTNL2pE3o/LZifyNuQ+
LECK9weXzaQ4sKtxJhgaZzMaL9e8r1X1Yp154ZTlf4xrAbufGIVlKUvE6VrFUvlzWR84uttm5mh6
pOSBKo6Q2ax0U7wZzXvnX703PFFBunLc8gUXsAsL7WMe/+ukaM/qZkGhUvPQj0WGJ1lHDJ2owO7y
yscfYkF/nyBMzVDcuyXsOdsNgvAsnfyjssBNriwBgDSVE8u0qkx78DHGcYZYCtG10F45YPNo3EoI
bV8EChxfjTMl7vKNu0M2BWdNP6M5sCWkek2Lm5U/l9DquMLjrWZhurw/bzoSOeq8DUUzO/IxhsN3
w0bptuMOY/eIwJSPRxaL3Cr8obSR42XjByDkNUaRUM+8byg6IpzhORPIavVhnYHsiiwAqSb6fFdN
uY5B8KyoqhUL4TB1U/kqPtOjKECnk0BvkX1pdU3G7sP0lW78ufoFYrpYHYzkKbhw5n/kFuqGXzf8
RgaMwAg98D3reLGyABQzASVnam4cUxCSPVCKCrlTUzNF0kdyc1NQ3bPTarvAXxDwVtZxCzVKcjHE
e6IKsYSd83H02hvesbmw6B5HCMzDpkXIgOLybLDLv2d/LJjlo+cBhunT3VSxDz0bN7WSI+dhC0Fy
+6+VZJ39+JG98F9EaFlI7VQRePMCrYphtwxd8/os7dqngY1cg/foLCGkeN5IaINvPTB6tBNlFnrb
+2H2R+SZw0mxR7YdYupbKtj+DGnyQYMuwYk52MKo2ncCMg5f2IygpGsnsn//Sb6nisoExsETlY8a
4bWapTw6jrYd1nNsLLJO0L33UdJ+FOpGQaMav1UM/GOTEuhHNXXzqK3U47ZCb088PjAnPY6Ztptz
XYqnoCPFYyP4GZRvafa0ZscL1cjMyDeczVeL7XcCn2B4agn+KqSsYot4eZxgz4gl0AbZ/aLoyB7O
ZFHahhJc4BSgoEbKNGN8LEwViTf3R6tm3hU4JCCRX+u15AuyLrZiTjL+wZ+O7QvAHU7esQwBwMvD
gwGKXz8a1T1wrG6rLTsFYCP+a8BMLQZygtOOB9+ILIDeUR+wcf9qzZZcrPbTujtPjUtaUcCWsBBN
gHcfW3BKiNbVzXq8tgeBjY1dBvFJz8W5Hq8qiv6KuqbFWg7g16JXPKkx0mcbbgn69dMRpJenf25F
xJsdxIMbTSdKukc9SKiG+QguCDyHKNlVjNa1a2HSkZ3lTRC5rQbLtU7HqjsiTJm+UnWCIzbnKhXB
6gXszGSQQdYiaW9a0X8WcbO9/Antwq56gedM+KwgwP1i6CNb7GrJZYpQcztzGz7zTY8ukpFb5060
E4+rE4rMmWFnIFgvpNCsoZjlodt5vQnDYM7elU9O1aM4YaB86ymxrS9B3Mm+Lw04in3Vk6LQ96oQ
T6Dek4Pjbn9yx8DeU2vk1CoxzREw9QBf9JoE2NkDUE+Is9q6oRbgPyYAk1iRyDKcIJcE+tzZrTHW
rgSghvY8vnpAW7ynmF8aC39PTpx/lWZYFL+oRgRhCKWoRr9TU/pinTle+I0EDbWig1ih/24ZYedL
6Z71sL1Qqmx9sPPi7Wjx6JucGg0ZS9AtaHigU73VMrJLejgS8h4ToDnNfcqu9eUh9gBmMUvTS7v8
8WDIC5d0anAD+4xCk3I8zAUBDexJuSqGZmelpNCVLyOqHmqWa4O7Y5FRGWnstgm2UTosbQF8L0W5
NJrvKZw0HsJBe9Uutc4sSvDiswbNWd3p7uuEHwj+HKwdC3gHFQ6jAeMPRJNK5HH3PO0OqLndkeW4
0aMV7gZNzmiqoxwLiuWxm0SjBYQgXlvfsUZ3Ea2XHaGhl3h8dpXHGnOgW0sTf0ETrzs1rGqcezVd
BxyQOkBFTKMeL3X1AJjUBltkXZBQd+wALrmW2TNeQFeruTEo46rHKwKUFdTI4H9rVczExsOUfkkj
/4GufSQdFdHWP3kLKnoPM6NALucMbZ54Pb1RnFDAeKBMbLgPX2RoMNcP3waTWP/NGjgyUAukcctw
8xYwzYs36ZgHtvwlcK2TzpDO3j+x9YVXaajCEcjCMfqjoTD3+q2aBJfyp/4bNye1L3I2xVeqA7P9
Salw4Y/Cw65ID9g6AFzSBcUmrB6XtUkwjaht/1nsR3LczomVj4huWBYcN5quqoy1YhYHyQuCDrg3
lRbGp9m4Wx/0y06/n1KZ6aSWyhct4uUo4ZbmPpTBYne8z2768QNR9f80g63xmPxyPK/4syzkz1om
fdBXNl4rUHerFc747wHTJp24z52fKQpfA61WwEVHgIu2Qadv9GMjO22LQl6a6OugRgBpk6v1vqNp
ZI+12ohFQHeDkgnFbikZOOohQ474BJkzfoQr3mbiaJpd2738i4Z1yaaRfErDnp4OBFwfH/+xeLnq
9K4CjnBXVX+8+MG0/wpvKdfVllo3cv2IbDeRJyhMvAtQoL4n2opf7XTJKhJuMSNrjGOsysVhrrQ+
csOV11amzXNQ1hReh1vLoyYh9o2uiKYOIW1BfkVxPlsnpEEjqXS75kOrMNsDBnLEsGS3h0lxhzH3
keDFATHtcJUhXyWacHSEdCZRn9sdxlyBHlMa3i/5r4erJ/jvNViSCjFIfUUHzLzTOv7btnNx3eDM
CN6XdDhC2+Tk732zH/jPKMzRakvyGpwR0HZzlu9dDNwzqDxvTrdJulJExCKzKQ5ozNsjsgd0rnsC
HHSyGwU7gow5tFotChvIoqpy6FEoCG87Lt8e90p3E98JohlpbihNU4SPa1lY3UKThGPi0q8bVagq
kgnobUr6iNOLaWZwnO4xKc9S5st/MMkYw7wabGFy4NnrNh0HyZVU08QQngHCaTZTz9KbTYiBLRtA
30WwHwYz28dWvDcL/kvkn/3gAJCn14rPi8wKy2MMWLkK+nynp55y8Tkd2Mt4c1d8QxkhgAHlhqd1
1dPEc+n3/cY5utAC+x/LJ/RtTXMU5FQjEjrZqzxLmfdV6jqXd+qGavTNZScs8sVdTHrWPDkW5p8o
y0pZFuB88n3UDcT9pTgPNYYTL/NbZZ9y8I6s7/NvycDq/3RD2726w5SX/zdplDpqLt0w4x3oWAg9
BH+n0zjX6VDZmO3DFNZvf+NhYKMkMPe1CK6uE7PdX/5btYSRK9/m/sgWmQj/+uQHcwKmEzVLEITb
wnswkVD4u5kgksVXaxv5uCnWemarjQzrPRVwTpy4q2T1nNPDW+r2keZsvq+BKscIIMfOGHAug2SS
8+j6vIAUmmUv2eJ4BBrYbclvqshSisFENaBga2EfjlRjAwjvuXgxwob9O1mU4iCLjk8yTUFxZUc7
fhnUiad4MPYfFkhw6xnACGQaTZo5Qxz8l6e/gcD9Foig8+ZniUHTaYEmI4DZnoslZ7r/FPUkuZ7J
eHJxBCwryWKS2eR3bj+OqeuD2Hy211tyBlZXDWsCrTnC92bB92JZu8OapR/JXPOz1V6o3aUdbdg3
r5lKil+V4Wza5InHGRrrotVoNFfBBEf8ZuEeNR+mjmunNpl4PD9Oml14riXTbsJDqQk83F2nMPit
4z58vjf3v+538QGbfH5hF5XM0CkHUhZLGayXIQmwpszCZ4sMc1JwMoVja90Rsb8ce1/nFF3Mxj7X
pbG4DJQOLkLYhZ5xtIvOTPebjn8HconVURoDFd/oJoQgkiWwKwzjzIid9+uPyrS8fktN0O2RWFBa
CD8USm6VrLur+2p2uAtEkQYKR4UcZBrs65rA07ShQBwsYUVTRWPKPUmqaGtUZND5IKRxsym7g5cv
Qyn9qfKFeH1rmplNWWi0MQAGAxG8agUtxAM3uiXtCySeA39dwIx7JCiKbzr7PeW5qH48IAoVoR27
V4047PbDPW5Hs6153mrk0qOcJYLwijPm4PrJhBVbPq9mw9zEQTFSNYOlsROd9cfI3XvBcacJwaRQ
iqzLivQMtKSeurCOrQT/zoZJmUjJh2jzlTY7ANtMc2zDF0QtoDCjMpvh9dQzPE1q4NAR5z0SaEjo
+0yhe4Q1SRgcSh/+UA6OYPHrfxYvp0OcAYpuJG/l6niZcj5VSsJN/YWRYaP349UKed/vJYJWngrH
1p6pHv6GZxo6Y1zM6u97W8F6UaMnHFj499nFQXwrH4fTLRJCuLSs22Fi6TkcCiXcq3Fvoy3ZrrgT
0UqEvYvLV84Ey9gsqQHAuJviHBWMUVIRwKRfxULfugabLMdsF6T1Uy7RmwFcmJHZAQ0x9EjTR0PQ
5eGnatn71pug/PG6EwjhPpUhpV9TMN8aeo0EVqe9BdFopoNzzUAEDWOT4vPD7aljogVBAZ+py8jP
wDHWDzaVVwqNss4JGqzw/5qv3fB5N1nrfC6Ds409nMh6aF07D57iu3X30ZTCvT12U4ivdqDmDilZ
WQvmuH5ahSbONxHTi+kMoa05PHZQztrTh+UTu72dOsWFUXVKqDHtK8Q5quPIk5L523V7BxE9mLWj
M/O7qHtQQvbHHOVsC1jnipNS5PXeMJMWfwySlpbKT8XgaFVZLfF/siGw/499HWaTAe7eNJWJxpKk
lYFS3AR/AEQvsEQWE/Np4iJU914OCb27IlG+9MtmLARFIpLJEPsjXQAszfi7FgNB8/RSz88ZMO5l
Fw1V3ImBIEgUax0tUdY/EVqTuh5t+mV4tBR1viBRLHyFn7WAo/INZp4MRTG44xPNsia/e226HKtv
May7fuT1lWO9R7SsiXdzj+fWqtffns7wb01qTVFex+cq2YmfBWD7xLYJYktByRxpbF/4gDd4efOA
inQRcj4jVkSZyD7ea23Qnq+tETbWf69J0lCLuyR2jLQ5zhF8ZfJjBsNK/hxgLXgeabB1DFIWSQkF
UyErFqUu5YSd38VzSHqLILmG/C+qBUs9ODdgU8gHnoYkP3La3oFVjvAM38rKSDvaUJRW9yY9+qe5
z0/gx7+wCr298zmWqq4DBV0aTVWlnrZOryzBiYAq+pkmFsnzA7T+eUJIKHctVPR4kmNvC4UHaTrC
COqlLW2GPq65+xZubgDbgFLfcWBrbXl8vQWI858kRpC48xFqPGJVBzD/s1Bp138gEHlkFSYbGcqB
CHc+5t9j5XbsQedd7UgHs0a+IBEf1S/2omcUQnhgIyROlL93O2zYqRM//HHlxfxLahAu6mbVjaDK
U64gHzL7BZZ0K9ZL/oSJCJd8ZnAlbqFiY82URTlWEbEFHB1p2BnqZYNVMCaxG8ieyrzFKujBmrlF
C1/B/nBJcyHsmul5Rp/UVRa7wTCLAKTgmLgk58vq83qXPR/q0Uv51wom12P2QbaxlONs4mux/6Np
hlrgVvM/Az4P0s4mM6Vc+EIJNBf+dMtCo/QLywIeGOcVg+jf87vFnrsfGBA/d2vhQD5ueGKUSzp5
xEqNyhAFE1RPt0q4dahH3hkXqqQqbE2rTSQxSF7yK3XSptF32ekTuuwr5CSyzXaL8KUG6PrEofdC
MRs4hpccGqtZDpN3jtvw3H9/gFodLy5d3aJFWsJMT2IRCsDVJq0cn8gCRTbe7A+tkM15uixm6yge
hmTk/VGv07wGF1maUDWwy2phYhqMWtKxqMw3PfySS9VXS/O5bd7cYPYDxBKmRQYZof4pZhSttFmU
I/lNKocad898OQ5WGlqBTAAd39P7tOPUA0gvYhmqmerhDEGpoAy5NS8s/AbRwOWm3TDXDMA/6Tcc
gKq0t9wOlYyG7GXWUuS4Un7v2+Bg5y0+PUrzNL+v3x+gcIlwUyz6MF6CQyXOPJoJz+SMccC7Olav
pM8bF7UdJNLfN4gcOZb5SHcDyqj+DFzL2ALjXMOH8JR3Kcb2+ZCeAFtCltLcal9Y6ZhYGdExLDk9
utBKY9zpWKhaOC9pPmHDmwf3oG+GWJkeA5mSRB2U4fVz2eMfKQ9djDOFzSJTZEyESFvqoLu8T8Y6
+4NHdsI+FRj0aEL4WdjUZ+7wF7L0/LWlSzcAZe+hn0dLTUAtptWLz7LOf96D4gLy8uLiLdlIDvtO
BmlSmmfTTc2JxI9eP0gejmwc/rRwNbYvvR6JcPJlUaSUIH+urUr0npehGRa0M4gUuB+173VCuyy3
aKfNq8tYvqXchYKMUCiQ2o+uFdMnrZ+g21W5ERlvJlpGJx+pKDHtyqdBgUGuqBAv42HcEARth+i+
JeU0taN4REvFNH6HMCTdEQt4rNoZUj5FZFU+rRynKCfQF6rV0Uji4cTwt4S7MaNyRoMcgiVAJRzY
Si4WyfQdaSq71HvN5mRAwLO9s3d8xzUfA4rxBgYeQ7snNc4vp7MRck3lyVq37VDy0MxuxCC3+a1T
PaQd8VzS7++3L1Cr2HbZBAASJmlp7c9FInFmhoGCg4Az8W7v2jMSn96qAT1Ov7a4pAUCstFKTKI1
yMBZnXAt+0lC8ABLsqNvJcopNwSliPmREXumtR/W284uv7ltkZtKkr8iTNaT27OlzqWgnUuUfrO4
sbk3w17BQUrMQ9YXGpRIdo0KtXwyCDWj48XUItqn6YqL/bP/SLd7uAOEFxZ1rS6aACvwWtMnxF8I
lf0G+hMkGQJAU69G1PiPfE9PIKQAwZIdtUHXftnHdr7xh7TkzpWfFUqZWN/t2Qt56jWUwdkSEwP9
byj0wVEE/tDS2MUpIy/oitURkVU7Iuq4rh7i66OOWLXVwQyQWl4F/++LKRBAw2oSplBVgHaoT27Y
mYguiRoFgGSHiZ5iGdw3LyzMpnUErjRTjSE1ZqhJ+alZfdkFRMHzOAxCVrcGP2sKgiAbo35x+Moi
34bq7EtcSrBe30dTSJ3Wrau7/U6jh0X1Q0KKIN4dHsVEQ+PV8eOB/1/vgeHzTVpMxreOfd5aE/Cz
GSETqMj8ym19jPymRWLE3XxnM7S55nD+x/xmEaq8NpRfv3YeUiVcpx0Iz3cH+S5qGlwi4EKTs9MO
Y0jG3gLonJPM+lfjWhV98rwYcTPKDF1VSlJ7+L6mTMlmyOmgXwdhyvu4DiTzhSBbN7+tlulcbogY
oTnVVbGon4n7Z54zRnzHXJU3MHpbS4vGCoVcL1VPL/pbmVL+sy0jsBAAL6qyIXtj8IuO2GS2pJPJ
UQ6aE7YdtU4f26BhEhwBACCdgoUKKOrxeMtoYPasHz64QhKr0J+0nTT2kC7NHml6CgH9KVfFfMf6
A0nQ3OAPHewb43TpQ2bbctPGrMq5fwrcXXFzrwJjkpyFAJA1Gu+IyR14D97k9s7szOZGKEek+Sht
LNPIwVmAVwctLjGWZxA1EEmdqYyepP3OyEDbjTIbI6+025DoKL38MIqJAOYr7pH60nDjAR+W/i2Z
ODMTWahwcR/KY7pgABn/uwuhtsmuM/13+aMaUEqU+htF1whz/1zZTWeq3gsUwApaQ1LzjKAZmcdH
H8+CYRx9ObG+dIE2u7g9DijxOF3qNwm4wmpje7mXeIL6q0H5Z0T/yzVXHixW18HVBV4H6OfXL4JJ
tsLsxnXeq7sYdKQmDb8VPOcCwYDwXVXJd2NxGxY/aGdyTkgDnyv5G7yJetjgUyEplYrus/BUXNlc
xl9I1rHMBhMLN9mJTs2lpYMAlnruAFPcmW6MsfucGnF4lGXR23YT+KvwBsHSiyAbFtp4sZ5Mmok3
mPOyqEv74X/6PSvKXakjztBjHsBeo1M5w556Cqh5sIe17PwGBIWi2VKsw105j7NB3i8zNarQe5W2
uSQB4YW8y6M9MrlfIxd9iAwbzc/XSZZshtDAmndCw8Wq0zb5ej8DYiQHQYvqSv+++wJkFaeii9NE
Pf5KnI/iSd6RC/lp6qf87ZGoF+o54kzNFEUs5D/+bk7ia/OPGtc8PSR0FMdC2d5tMfZe2OaymFtv
4hU+vb5XlA67+ptom2CT37je3/SyNwpDIGWLQKxgSqWeMxVDjyXGvTQ5tN0L2IYaB7W69obKkkGS
Yalg5ybD6U2o4T3yjXlMko8IB5VN4ser/nBprncyfO0Bv3XRhA7zwJnz3pxdQroEZ/wVps/6/nvm
ksNkhe5kNuiMqzZtpQNliqMIV1IUK0gkZLFtsScP2Gs7ipd7mDC2PsH0Ve1eD4wMzg2gFldPuDze
6dAAlutmcwTO99ARK5339ChIVd0JCewIsl20r/dVbxLjPDpczZEHZqaoL8tJTH096QZQEPDlHK4p
+vkR1qPAnrP1qEiqsEuexz2hPN6FDTo/XxbKstjzE2nC5ib6dYqE1DAZCO1dWztl5mth3zD3+Tq4
pQLo8A8U+deGH/IbTfe7KHtMlV7TrSuGwuiW3FXf8v8K65oyhHkhm+npacje/QJs4Xs0wBFGBz8B
v41XlhSu9l4JuryoFqbQRCNUGnEGTyTj8JdskxdcIvsXPxIj47HmVEQt7OJXSWboH/R1SikXphcS
tAaXCBwMN6ckRo7GsfJg+I/dO8BCTjoQv1pBQ9LD2tq7/wBzkDDrP9UJodkrRQmS6rzSWThjLjCn
Y/57ijIVi44gS7nJjQZI4DFMOVhQ50mOH2UMx8c+lQlFJZLehvJ0WXfxuQbAYjNA3wXOCNkGs8kH
xggDDFjXNvhrtgKdR5T04R9XdPfy+HOc4rVjEO3my3dTmgN385gqvypZHxHpZYuYa4RdY+1oNHr+
LYAou3/WfCd+LR760NEhoPddASai4sP4HKeYvQ89rrLHjbjySYT6L5xS1kfytLEupVy89MYz1EDM
S/shL6C04rFv5ydNYoIgIc24jX9ZBjk2Bp9aXMdAegEXr2INXcBLmq0cVyLBTqUdDUg5p1snMYqK
racKxvG3mlgJ60sKVzV5kWRFOpT7D3xsMCCoBUmaXnzIjdAKCLnnO9tFigky3t3aBTKaPec1nIMq
TEsXF4QOKT+OdXpc3mKGk30YPAqeNil/9cevsoDEWvNfiaFmoqbxnVzoS+LhAcWnCXjF8gE4mOhZ
kQxpbqX3itr+8I4+O2WGa8lLcCt4es9o9hBsI1GN6hprBh0DYvgiYvw2VcXlUoj+jAjsnqGlqPed
m8OY2/COZaxSEQITJDC2BJPsi88sMqxuqbtLtalIij4eMxplpQ+/BTYqBUgy8xaItbtxG/3Bh8Ed
WbnDa9NS0DDkNzxXVKSJpnKioXf/fgnR9T4a0yadWlaeb+AXm8L+UGzoXSxnwTqArtAGMZL6Z7Eh
aTPynR6UkL70rlVRztLSFDnd8+H9c2KQQjy92dA08p19rk6//hDJvbSzxDoKglf6U56Lgl11w5/K
lYnD9NnQl9665OEsf8NSebB02pd1wIihyxkw5C9zIIkYwhADewXIjuPh/uSkdT2S8WOoox8WVTxB
BXtI8IXmkiTljciv3vtvXaCyvSna0sAFnarm+PjXF2kpbebj36WSYezbDcrtZG9BJZwjw1Ua1eoh
gkUgQ5qPRs6N29CEgAg2X7DyiV8K12bbvZdzjqZSkZ2pWFt1J62DD67z8oA9XtoVoPL1j7ZRPsKQ
pN8Vo+ibjqtVUgghRX2vYWsTPT7SBeqnHB7mxfXL7l4C7VlPuzkIrM7ng4TU6cFtLr5DxhaSZCXH
ar9fSaxZnXca2PDb9Ep+havvxpp3CQJaYiI3ymO3jm3gb+Eo0KBmCkzQCM49WNjUDP1ea2npg053
pnsyJymWF523fdc7+mF71vXayEJnTdpwmpTOnZEy8cOoJx5ST5G/TY7xdcxJgHeGdU05I/YvZlYD
7kG0ClZVdQL12ZbQl3ADFrig0aBNyrrUo4s+bdEC8mj8u7Ygkkp7wb8Bu/oMR+f/JjrqcmAWUxW4
Q07ErxFCqHbaDilcpCFAM54vEMsIOH6GwnYCOULqgpX9h6VeBqoGalqb+uEAVo2yfZRb4sbEas++
Ec8P40Eq9WX6mNsP7RWi2N5AzOKSe1eorUwagy/zfmuWC/K5TUi4N1NRz53CW0DJFj/AdCJpUC6P
uZDzrq65bRCGNuw1jSRNDA1l3jabLuAIepZPQ0TD/4KPcel2fHl7/9z9ipBALcy8pu1cLEkKt5TR
Bh3cc4hn9UZTTKZCy8dZN01H+2y+12oXmcmXhek4D2f56wzf1fP/kANKj5y7DSS56FVG0uwb94ZN
iQUJAZMutWZ9I6R+Z84aid7pjni5Aivkc3Ls2aerqOUM5RNSJgCo/ze8UEP8K6QR7c0/ncHNaRC1
j/kfmxZW5EcBOorXDVayK31g3dfRDlBtWG6QIuZ5IxSJrXRrQMz69zJ5MSUyVl0G9hk84yr1tgqF
WzI58B8V08HltsMuTpY9wmDcDJ5Y7rk7BjNf5cMvpcGBFPoyOL1T9HzNcKtNpx/c3ZG7+Bcvo1zm
vsom0lftbqwMb0YOrxW7Z6MfzaRRt6Xlo4sEYtrczYD5u/bldojg5krLXMtLBuxu5oiIC3rxwD3E
korhwQ/H8j5a6LE64LSaeWtpt/iriPQ1mhhSObuLgqIsXNIaHjYLdZLUJzmz4hbUHepfBr1qDwZ9
1WkoEN8LDdwged16gpqMuXWQkOXPrQvr/e0SqZlBUG70wqKmJdFXw375EO+E1bpEUNMPdlwBPixc
lYrkmmiYWgaHcgC46hiQ2SHAYsrieMSWdc4B6PnWAF0Uqe2A2LA27JkmLXxnEnkjx3QeXWWAdISC
i80QmosQysC8dnGf3yeOPNm2a1p/4/R4gn6oHJAgC3vXRcBpq2W55wVebvtsbc5IlCtJA9+NU8GM
1yh7CneIKaPYvmT3vOgvhJ6TK5ocri8FxbSvVSd29CP3NxYgCk/E/7MYuppHrPp9LwZXF9/c7fEf
ahSDnVFoLcHm9YsUgCgu535s+sD258V1D93D4RJhuLsIDu0BAqg+ojKiPyH/iqYss1WhFD3LqPlp
m4mt1s1m2ZWZ4IjUZyVzYJYC2f35Wd+bccnNMp6LX+jWHHBtZ8GwVK42NYSPqGMpottFPldIQGPa
FMfKjspqitA4shvHcWSwuKY3klAqFcM1dyBeHft7ijCPHU+J5AroiiN99ZLRamgjip+dqnFcNd11
r4KLnZY7Vw/yjaG5YTweDxuKrDOu8LJhkgabM6SUYPxHu+xjLF8o7gUJffOOqpY6XgmBrXo1N2O7
g8054TOgxZJYou4A9ZSoKnOB4IDGxJMNy512h9n3obJmcEcZvMUvTcphXVXWmiYI7fmHibFI868U
SoLrQAh3Rt9651d6X7sX2zluC/jZVdxVtRu5EkcdkOEX93ShFZEZZVu92Y9Aaah0767SCiILUOWy
F/eXlcF/0B7VAv5LrLw910y7krJvK0wRuAH7eHIffr2QXOL/dAgkrGyxWw2n7KJUzX2LuaWdyvUi
Y783kCAc8n8x4VFK05z7GBMg5m27e/zZHaNlCOwKD2m22IlADtxDnmuSv0t25WRRetJE0+J2hCip
jO8u7m5QJv0ZDueq7K9wDE/bsqSbHlJ/j39zSWt5KnatCWbNGB0ILohYOKL2PBlEzx76HT+UKk52
FMRtXfC3JSvF/iQE/SgnvfbKJ1zVDcG7N1TiZ4Dd76tQcoVIxp2jMFEWZu2Cntbwhr1QmDlBYwl7
Pe69G4EoxwW/1YjzIMBkBr1DJd+1bXelpCQNmm8XegJhRbsquYdxSP0JdjUKpb8tDWpV6/058ETe
Klo90R5LiQbmfPYa3NV1ra/GNUdv1l1cbNaxzqAS2G1hZW6s+AG8pHyFH0Oau4d7zFA+8LJHum8q
O7DOj6IDJ9TmBoJy68YmyvgBhwoXg1rfbCa4/3mk5nM7H/XGzYWPKQL4Z05mXNfq0H85wRo4rlfv
q7i73rjYiceI3uEt0TMf7a60rSAle2r3C6xaB801VzJ61agNlnSlAxe447jESfOknIDP3Q7OZMEr
VMod8yOb4jdQwib7EvmvhE8DirFBgneFzJ2JQLZUGGrn0e0Z1b0JExjbNIhRypOhNa4jjVZR60da
r2TNzrI9zYQh7G8wWHIkqRm5wzRKLPWIVa9ETfThOzjG3NWwAdoZbGhskf9zIaOdtPgjDYRmNRzJ
f8HkTAoeib7QK6/3+LwZC41XWftfyZA+/Y6K7Rf4NrGJrWbcEarghww92znqnD8afBMTIYlDRNRy
cZaYhXwuP18GcDr9cSTK1LBpUrtrolJ23Y2/CbMte0uVhcsd8nU1haJAtBUKVYwbLEWqGKMISXbu
+S9P/tXg0IH8RIJKE8LIBScIgcAu+uVAAa8Bndqi9c4jq/ViE37OUAHgAxdw8Q1govd9T4bGEwCu
+gYOiRwaNjIE1+Pcw+XHHwpoZonnQc9AHtP/U0AlPBN26LOF5Jg2eVCKk+j5LQYBALU6rD3EUdsb
h/BS6kvr43I/WFe6QDa1rgjfwcpIv/Rzn/GeKE22+drVWbcI4dR1VOQ3KUBF0ptTCHx78zezZFkv
lSWNWHLzqLoXenWGYh+tQx8mCLEMbi1GOjTl1zv5/LGu4cdgMuqI4nF+Uz+B4/E7g9PxNMrTgdFa
xQPvsKMTPE1JB0+CNiQoF6jdVbx4KHayVXEtilubUxyJ74wUOPSkhS/Wb6XqYtJ7P3srgulVUSaz
FA33y6GD+IBRAHzikl1pE9GewnPPZCnakqyPGwuRmpfHhJNgXndhtboT8K6p0o7GSYr7lyYoErFi
6BMTnb5hiXfzdhDlyWFG3pInCD02jv+72Toc6/Tl1m7s6iDX4i1SLSlLP/P3ADrkZ2+0tIEHnbfR
Jk9fYH4pzufB8i5ygU2SVc42v5bQfpwCt9otEbcy5iwosG9HromKYe3eN/wJ/5+B0QdGhg/Fk+jT
IYPxtdk1sYWwyJ5c2a25s0ymgTgmRurV5WnURMynn8wl7gBWk31ngh0kQMlcU7RBtxzKbXaBpvLX
B3FWUJOs8KzkkuXqcSWN/ths9hCLtBmsNPoOORg4bh/RqjxTSoGDfNwiZrsffSDeTUj3862ki3+m
GGg4WgSBEkjX3BoRFGH5sQZN+Irvr10a9Sai0s/zNrcZGgaxjPg6Wvp1Gs894ctNexNSCKYAjj3E
3LEEfV8DwGkYgO96lCrfOKENcfkIkEyjeKb9MxhGYBHjD9D4ELAMtVIWIgrwU6ix92iuPYXEikRR
r3mhbby3cwVtHy/yKyuf0m5dBqtPrfQ6xeYKd+N8+Gzp7S+U3SZnWFMa+t6hvKiGX0ijglmb/CEw
S3inbRH59Zrzr4SAZcZHhGDkl/Jzi008NkYdRh1Vswq0y3+1fUzJUX1J8Gu0GwI+9YnmGJ4Qk86B
A83gPmNQGcGEPsRpo9VgG4c0VC3FZa8LTSw2jQWRYvOhEvlhnIIm4ZeQcW1TR2lxr4qFRYeAtrml
AcKxcGN+WWi63zX97a3SRZ8N/4U0PEzaxEFNSclLpgQB/Fo36ks+jzrIZN2WVQcJOhROnt3j7mlf
lj8D4us8W1brhF0RumAh7ahjH4EhjIdYM15pqjr018/fMOS5HVOYR2oVG0spovid5nKX1Yq63FT2
INwpQldAXcvklC4vhRZytrxHtWpitkLkP4kZ/4vFGVwdf6WG77M9UbznkbKQ5EmXCbkXRPg1pXGN
tb8uSNPMFsxMC/LPi4+VahbJjkBcTrPY8jaEcxRjBKOVW5NhMpumtg4IG2qr8dHfiI+x0C1E584I
4JXXjyxabRQSfdPIwT/hyY7kKy0S/h0MW1RIT5gZbg+H/UsaWxREMnY43k+mbbGezm+LaPP6vnRl
YyUibwg3KV48Q5iSg+aQvPeZDpByJRprip56YNyMhhHXksDskJWW25hwQuBF51A+hC5no2lJgGc1
wAmIkKG/Kq0FGH7mcoW0qRqiVMpM9iHSnZNhF+tRjE0D49Zy+VposY4qgx41dFpJv+WLmnfLvgpV
YgoBvGumC1lrDT+X0voN/cVxhYph6FYyqknu8dYSax5Kh6OfI2ek5TH5+BCxERBuUUpEsc4a5X6i
Uhxrc+8iwtuhh4SKuSqSdfm9LA6aMkuUXeCW5f35xKyMyjTNe5k+ohIj8Ief8fbOYY5IaLjz8ppN
z26HqsisZpDzVESC7v2wK8/NovzeUTKbqNXpb02WykNThsoF/EnqrBfOihRZtWyWYQJZqF9w8Ut1
qT0bMmQuLrxpgCb0ldwshq9kX4bmCgkF03vZYQxXkqu574p4XKzmxAm1OQSbtcDQ9DsNsSSn5ppS
K4Z3E+rr3L5bykmGF8pGS7qrfhLEAQCnEDo3Vx79+676QBT5jL/iv+Jo1BUjxebYxwxbbuMJfZp+
acCyDqVThSA86wDNxf1vAyT8Wvor0jg0SU4vM6/EQJ6jKYNkSVzwWgsyP9KBZQoUIiPPt1q2nKjF
9SazladJcCjpoAv+d5KzgeejVr70osIWEcgnuz7kxsU65JjhdmgAfqebgwHBCZd78DoDkilGQpQM
9js8AorM/5Of/QqmvYiYkc10fF4GBCnGNs/JbbsMZzQ2DUJ+rgBTyiqroEpV0xxX5hqUvC9PDXax
RtnPjnP/ATWPNUdDf53PS6q0zxabOK5yQ2U0/IMf3wjxz8aXwCGkL+MKaw1lRv5zY6owq0m3Z7bA
mHYdw9uUCoo2Xsz2gNW0lQ5UmRJJpcHyXiUzzXk0AkdnYTFSdTj6iAHWBHhEmyqWKhKfx9stfRgb
YBUSyzmhI6oFW0OXhlZqHAFQrmuOHjd7TN8/nBO+VtztpQZrRxPgVsew5Uk8OkxrZ77tcgJs65Os
qxLpTKnz73HCI763hhQgDfO1MrDo7ejgaO6Nx4LXgAIom86qWOwqF9Grv8z1TFwlgJZUqrDKStad
MXMDCxdJHlvKAuMpu7pw9l1WvH0xpi2B++JXVsOTJCZGY44m2Facy5p3UrmR8YoQIPsWvXbG9eXR
HhchLQaM0N421KdrqFmr9RITnCXlAvjBy/lX8YqJbBVmPcMKJURF8twwQvkREXJjK7U+cv2G0vSf
dwR9jpjd6gUjqw4Bw3qZA1ZmGEcsCTrtk1CmgN6aWqw8ClNHPz6nELXeOJtJy0dEDdTNZKRT2bjf
XMhKjgmEwpVCQAkks6LIXRo6y1rw29UJMfhj2wnH7kq2YOH7MmZFDJtK0VlcdBcY4qIybNFarPjA
Dof5yGcd0EqpNZQ7AupFTBQcUL/JxACc06KjRja6+CppzKD0oQUvvydAiuSUPjbfBomH+KKJiHra
CkGZMaCgD0GP5RYFXkx+Kls7uDAcs2HbJjLUzxb+aN/vbqvZBPcW5DZuSEq12XNFmVgTYmEHBUQf
JNjHv1ySDm1ikSrPTLXQd/b2fne/IrbCD9+OnxJhxJrmsQsO2zwdWk1k3Jy8i9lFftomjnq0k6hf
w4Z6OrGdjVOnrZU9mZbquVDOUpMyCa8ZUgcQHvleEaj1cJ6ObyUSVjNVvKTa+NPehfgE4eNfgdM8
ytPlArqtHA5K1fT6OnJpym5CAsUSf/6poKcKd/nWaS8i/xrVSvwD2+MN+xRjrwCGp9jYguy+k1ne
BMbq6p0+P5yY1D4h3F5MC15iUPwU9h2YzxLhj4vDHI/NHLbsZnjMMuuGCLLyagsPepz2c2yzv8re
u3mMrbCF51U6RlBxBiFv96Q/0Micymq+HF068/8BnqPyafyDHE5LtV7PSDt6bQi/HMN5PEWr3RPN
NymMUa1zlJTU8iLRsyzI39OfwuTdV+EdDybDMRQOMjMeUHbW59tGFgxRzPsOuuAavTH1LtRhiSKt
4lnIc27iodBJBVU8rWZeGyQumdmlIGKfijAqvIwnpMd3+iHb5Sd+jU7jRUOxRLggfW7HrDAU3DfR
P0y3zYGYu1FLxCEOyWTzYLj5wmz6gxcOzbQK72bySovNeqQuF+VJph107krAgyurZ1tYDWbjdSjS
rBsu22fUy6bDfvF/07jnSXgNTi8Fr5D1XQYzXYewnniyIvuZdm52Mhpmqh8E99m/uNFkJ3lX1E3y
EaanTmZYBZ1ITpEwrE7cHfE7SKBCqOOlobmtuhq/9T46cvfBUYl0K8xj4qbw8aK+BMOkBSsVYJyJ
W6FRG9HsPtKV2mC4tZaGzxHlo+guVp+lMIrF8+aTpVDR1+APCf5DfUvum+6RH0VTgXixsUrYqU7V
AmWy9gEqrUv7U0eXVq+4y1la7uWjKMXaSavr10+MQUekLqf8CJg9T41N+LxWxeI2rXj9U/1eeIG0
uxY0rItgLwMf8pg6q6Jvq5gZFwNIpznp2cEvCB7DWJBT1JwrPMGIAzn15CcrArbDwUQKoloE7X5J
y3CEMzZ/9PqGimInf34od4sxn2Am4LE/e4oe995prjrac/8kcttFuuNIAHvbIo0M2C1eBHtuoraA
Z+97SfRhnO6xnAEV3urS7R/0ZrLXF39eBNj5YB/YiaBMRborzkHyEugPYL3NdI2dHMzhTRIfJ1E7
hYjab96MqREytkHrbY/03KZlf6jYegWdzcCCXaB7+JYvj0wM2/BtzYeNDSFu+HFAKdZxX+S+RAmO
QRSxViEiSfa7TdkMbGmoHMZ0kzyRrT5ITlGOZwecK2M1EOUH7izq1PUELWuDWlgPnv1IG5G4CD9R
QEHZ5TwWIw6JVvyKpX0/Snm6pAXZgXUL2brN3YIbO0K1zYt/hF+tYJ6cB/IQF/2E9458iH+xON6o
Oqq1QLo3zdM5WMURcP9Pto/Pn1+S2UKQ9HGnWGJsbxB/cIhDwJdGsZEYCmO34rcFLKFxlSeFBfwr
fCJAP1vYlP18R6h6Qrx+ENmE+aA8ez5MtbtaFGwyCHK8hjK27ArGPFIwdbJl4fPC7Mql1/JZ0yCX
pwJH7Qt8jk9gPC0rpZFB5jhBZls93UnHIxqlRVsDPA0Tr4NejY/tavdDX/9mbPZj/kQWLxVBIcla
6a6xPaSESxA+Haqa7CDDjOSHqbBgzAdVAcc6FnALnuyIqcPMJ9mY2A+RnftcB2wpUYgq3kzWT/9p
b8E9IV6b8MTtLBEyOT24e450AXCtFbkvPtzLfG/sTeBJItwwVuKatgyeJE0C3BO6UwgzYLruyfAm
yOLzhmldySx7hwdhQ2p0kHvPRhHypNVA51M5SWxvZ4fY+PQch+cTs37rY/8QTuSbDj9NrJq3td3r
P1M9W+eSCIL7tMiod9gY3LVaBAHGIu4dyf68smTmXeyNYqzxshJfgkRlkEWtQBGOlFTrzv+QBqTa
iU7OQIdj6jIOVMI/pX3dHhEA1hgWL1Na2Fy5lrSDua60KN07Zf2qvNxFR6osTbaWjBJL0+Y5J/6y
uSrEa9GG+9oH9YhWmwnm+bbKpycK73n9Cq10NoSvo0X2VuzS9gKQsYJh7gw8cNJ1VCYfYrkhWN0y
xQ74haHWCg3wpTshxvh0SySLK287xRc5gR367qTSu4uA+W2IXAnCOxhc99UO570UqXQCj90mb2yf
F8VlLCWdKT9EZwZkIoFvRM8FP0AJJSP3HzrZimcYWn7DJRUpi0lC+Pss8b1UKzaDxwRGVAiqI0/H
GZolCeDacAx+/abbDV8ekgdnnb7fMAfM08GupQM5rrsa639v2DiWrB7aZRcaYZTik3s0YFWCBvC1
yop6PkNAHpXDsOT+MHQudIrlh1ZOdRMTu6/kk1hh+VSXhwNevSrH7fZLc1adA/BAzHMgcLQdjadj
8+9cNiP9/a8v4cKcC030apLlyp/gLGasf2ROHF7vGmpf5xduCSOOVZQctbZrM3OUlEzt5afdASSz
Lclxpqz8dns3M11h2FulsGe5tlyxGYLaJZC3aWSObCTL75//VKZAMZCocl2K2CKlzq1lP2SLKaNW
yCK3BNlMxBnHJpDDCcKcIRt9GvvWstbs+b5PSqJ+awzNySQVLIMQvaxSis1VGaGofIBMLuLG7xPh
VhJsQkXRBhnnlish1Rq3uNADYc6Fq9xsoTcwP4Z/+LFhv1M7kgAXK3kvdEqzPNfQF4l0a8Q1/c49
+Kb8xwvg11puiAtopJ/bJfUZ5aaLAoD2u6seLGQ+2MolB05H9AiU/kmMjTCL04IrSGqOeL7Ogtt5
zPOnkb0JSIqlba8RE+y+Kx+zRFvxYzUjBIiEVN0np0oxRdCbM6GTBFUUDgSCAlZFFmegGMsdxbhh
hZFhRFkXwxAC0FceKw+Jc2w9aWgzwd7b5C7ys3vQgb5bnDJzYxrd6UpdBC9lot1sfLuSroh1hFqK
qrWOPd23teQ0/9w0HFearcR5RzuA+ncIMLJUy/Jq3vMWk43fYmVNcfVQi+0zpbyJlFqk2cxREtIU
Zp0EoP8W3+lQhuhth6pfKml0ijG+MZpvf3bjqItV9CBXCOVhLm2xNZYTng+JD5j4MEW544nS+ch2
IEF3Ycu5Ul5NOhsKJNSk5uxAjjzDS9TsQikA6ypSCJFQcef4pt78cZ7KWAgzF8Si1aUx311W7ONh
gSLjl6vQjzZD3IXPs+i5uB2+j3k0jMD7w+bwaYPM0c3XtkgsNTN6sJUkttdcDEXehfPccXbmoygx
xqTKy6Bk/96D3PUBPrbsx4ETvD2lPBH4ENyfXhUFkNtZ8L4DitpJcTjxyt9MqsZvxUEeunoX8tof
EPV/onlpgajxfWhY5iMJ7xE2YGlUbDll45LtvEEmhcjGNV5h4e7QqWGY5fEAXgEWJkmvHSkUTZee
H8WynQ8SvSsEfhvUQrM4QA5uVGIc587HXlQgItrwHvq0BX9tEQYn85NwJR6FGEzrwtaoJynRaAO6
HxsBbQkBstIeGpqLy7F5ieqKcTyIJdeFVhzCrLhk+KsDtKMPVKb8cgKm7p7dhiwJSfbAXDViV+6A
Pntz2mpoY5bymnyt3CiloV+Ip+NwJSCG2ZFU6FceBa3QtFE0I+7cn5udqwM6PgvZd8tDoM3B1C0j
jquNR/Pf2Q7rKIS2g24M4FmghMokuGp5YMXFtv6URRFolpbVKIC2IyHkerxYV0J6D4nx/mssaEqO
FkGyFqtix+YIsFKVgyAjgnlSu9RlsF+yTLIYV9dvGmj1WrWdO0C3zTtv+8kn3gzpdmIsU5ZTCgPt
zNG4S9efMetWnwM/AcBWKmO1S5712uFilMyb+FpBAeoQ0+6h4BknSlsNlmh0EHBj5lCWubfluLxw
naqqGOBH6rXdx3pj/D642Lrz0MYKQ48iUZ0ftQoLqJvqQv+WiUhqhsnS8Jd9QdEg6X4uCu2YqCSP
GvKTciAdOiasj0DhBSbfLMspc1VcR1iHDQ7AMbTceG3liAHrCZVBTffj398Fqv8hG8gDnGS4odqQ
dIrLRxLxtqlpWax/nMJnreMaewOUxkmeg3RUsah0Rz+tFEM8G9fmyoOpOJyEMAlhhHHtC5PSkt8E
566yhChwyKiKlzs2JFy/mXBNdBPCw+mqOLrh03pkM8kGsEjV4WDrzXz5L07U5rgxgWdJlOnH+UIM
KQvL2za4J6vabIOgCsokrcn/N5PdbHPF0tBp+2o5VrtDzwW4OK/KDsplORLY3LygpomqSObFQcEG
WAEgB5W3/Tg+mj3Fk1pYGfpJPX3/53mYpaFd4uN/fNYBIEmkTs/NsoA+U6sf/QGC4X3S5XY49oYo
ksuPmRNXa2oQwfaIFXpi7p5wedRsnsBqa3Y/G7n2hOZ2AVM40F8z/E4xEf5FMzViCmTP2C6+UQPT
7JcLzE1fBWugMpqzTzXuxKxsVzEnL8Z+ZvCsR/bxYmSiem8VX2g/A+57CxvtSlKZaJWgy2MZiVNd
kggcCiaY9MeYAsYzWCWPGBoA+cyettoRGiuP3YrqOC/ij9q7Uz8Ju8N8ghiFSm9AKzQ6VOonsI/8
Ch685kyzyf4ugUhtw0ALX5C13zU8MGpF7mFOSPvEIm9TOMYZDv6fzzFKgFFLZg6fx62Fy+cXvqMy
4Up1YrRxT6lwY4zuBEVysk51AFw9ysm/bTHbROxWD6qiEqWDNPaxwRSwVcGyXJ1FAOLFM7t9DWCR
nKMtAQ6VCFxslLP7IQFtTeiVZA8wn0jQdJ43ypiJmJpZjinaUA+E2x86Th8wacy9Bkts+QRhxmUP
CStSQDLjYqCtguZBxjA30sV9W0a3mbVpEY7cfmdQZW0ZtJFpt/Rc/chYFV2QaOnJrJHaQlBhLOhg
iMqoCOEGLmgzC2i1r9PkWEIkJFwK20VX2mwg0AAnrsUWp4sfp7GRlimJR6ZFlL4EmtuxtymzEQ7v
+yX6ADSlb+K7Rhf0oEO5QrbroPWysG7E/+dm6M4Weu7XOWFSwAN17D3ysU67XUTjVxoG9uwjmljv
OYkL/ovkuiuhNdCSNX5S6cs4/8B4JYP2s29gvn6tE2uox+jDtWcgKSkz5cFsVKfdXLg8nZLVPkq+
cQ4Wia4DhGxuEs1HNI0cUHFn/rzCbbRELlIRmjlh7+jiIROefQoSE7OlhXhU07LtEtEUqRLwtfbS
R5lB2029RevFXwaDP3tVjAquhfFbzfEtsseF1rwiNnilagt6i7HLNlAUE28HynMVUXu5XM9tJSlk
KRO3jT7202EOu/jYsnb2DPJ8sLfqQmSzkuyocT1FKmxHm00poD5GQn3bit96jN0JjZxSMA105PRD
+Emuo3y2dGTPtMX1GOFs5VcTf8o8PqEj7HH9aeNBipDVpRQfXfxfuQF+XHCQKW0omW97hO49pRtd
ONIATKFiyUk1jTfLi7hDmpVzYtyYbPlRAiqQ41AtPhOUNhgXjhK4ibPBmhcTNHFMFcbfCuCKbTT5
4jgff7RDGy3rlajiwHXFOs+JOXKOV6SSZBljuQeg6Cf9l+9ISPZTgdJUvHCqu32VdhbDWs7yaIjA
N6tSzUDKNXLkT/t5y3T6mKPE4erf6vcFD+jMf8xQjtoT3u7mGKjscCZhn08mvMcgrpOfGp9HuS82
wbXaaUBJqEOcDs9QZDsQhZnGzgZ7vUSzAozYBtaG8NvZNSKZccoEOCN5HhX13fdpvUDIrrmSzzcp
Xnn+8B2hhaEjT+0MRMjs4QR8vmG6wJ1pGSsswqKOLIv0qV3M5VCKAMiuu8rjSQ9gKRig+qhrP7PZ
qba5WbHdXfnKeqiQuEzyh8eJUWe6fHBuGuSj6REikP7sOb1oUjwBbtoISJ9bmZXin6+GIGH7KhOt
JQ24tfsxsRGHt7f8tmIoxIJct5m9deSk8Uxx+E4LgYED2bYap/fJ4ni/237jFxu/CtvY1VLIrxI9
rAX5IzcQpxg2C1lOlgdzJtl0Rj+bNAQpvNgxcN/f8s+zbGLc1J+IOVdkxFl/4wjqHeckDdU/J/9x
+uIPjgoM4FnM04jPPCNJnig6TzncN8BfkWYzCc8/sFcZQWN5kZNQ/W37SOWBQTmjEv2PmEra8AdD
5KgfRcyrXcAAJCr0mBbLVXhjh7MOrHQ2CoXuDqk+hKdQBsZ+ctKsYi5Kofl/+uKfmBjUyIOLd8c4
3ZCZAI/fxwOqobdXUhyE7yDF84SHR78qdDHdU5sPFdEzVEmeeKo9XGGgmeTGUz0oWlhMhLTLmevw
T25Zx9wy+UPxh8uC/PyfaoJqytHlJqs0dqIiAgh8EI17pkiEQsQBe/appL4IJg2JLyYJXCT03S6G
wEPMUAEqNA3mOUpN5xZXNJhTB8/HkLbT26vjZj4C+dpUeNpftOHX9ez3YaPR9px4qRz3o9jIxFMO
Sw3xrOkT1oG7TNq7Kx5+Nz8/ZM9jI0pPRzvewYHCXifvZJcq7obpm2gUn5I3cKhaLMzconr9c1Oa
KAgB3vyp3Mq7unkiwpyJS2i/jn4q2bw08Bnh/MxNNKHqdWtdqpmI1tFDOr6l+AWWDjjtPEpdv65s
UljMI6sIFbWvX7pqWgB/+xY/+BehOlPx/N69beM5FBf08sqvKqqxMBirau4OxHdyXmROVISYfrbK
zDOccWzApYALTlxSP4qCAFylPTNGo5L+2V7cMNE3tr1RVlw89XsyCGUFwyrTGwB+Kx7JU411XEsS
YFwydtzIZ+uTmDo7QGGxumbM9pY4ieBOnvUMbo1jon30JdcJORONHvim9BMG3eb49SYG7//C9KtB
Inzu1Mntqj9zPsrPwAGOGnTqTE4inM9BCzQIRa+vGQMVZhc1bYwZ4K2gMps5flBAS2jMZWcnDwUi
1sDoKqFa7AxJL1nxVbGgTMShhg6FRLVsCbcnPm2nIOmmrlthua5kpL+CF1v/eqQQnsPY9scKbTLi
nr7pjn75KZCHr2iQ7+tosXlIFx0rIahh3JyqddCDniOCEE33+RXszzv6iXpg35gFhdI8qR+Tfz8a
XLQ5oYY1Hdx8NAURqgbtCvIP7CzQXSlfWjYfKTBdicxqGi2q9DwLdyOg4NxsPOQEry12KdJCbciA
rzWR7+5A/x8eFef4RwEBV2R0tLUOn+k1xJHFMyyNQ5fEG4dguRNV9b4sWar6V8v2B8cmrNe+8Xgb
dft8EBEqa27zaJUTZl7xsgRAG2OKNBMe22H23agnybEPUGqJ9b8EWgHsCidofXnYRGcgpn//EEEr
91AFON6M2AO65Itowqgsdns2/dj8Cbp49QdKM2CRoSk55QNv4/iyV6VZ1OzE8d0Rt86FpiepNblM
cLfNtnU+rs80NCIoEVILr0oZHn5b07kKBUPGPJXdf6cH9MzOSgbvjgFXlN3CWATJiIhNZU3iieEu
WJxUnZuXTk0bsqVv3GzuZXp79eJvN2QDh6uAqL+ns+QiWOAU8u0WxZ88NAAmzNsg7AzGkx5Fe/Yl
X6R72UKmNU6t7LMdIRNDF7E3SVu4ijcVst8fczZpPfajq1l0NiIJr2fuP6eRnPisYU4xlNJQ9TA9
XP5UShRZIgyjivfOWzcmSaJKKMNtw4pvVnycmK2tuPf0RP/kJd3B63dIX3i/SBYs52gqB8VwHTW0
I0+1rFv2sVZK/Cd8czoFJgmT0jGvx9dQqRqhyjrsk5TCeuAdgRY1sWNIEhgJgMCl7YgFj3BaKb1F
Ot2sggHH/DYvCZnXkrIEosg5IYwhn8kB/Plb1N0TA4a4j9PCObMR6RfW0lq8gTVlSZ3SRezJXXxm
lQPj4DgNVe6CHuAblhupWftr0VQE4XNqaucipFp5QGUjCIHxAMJoauhtK+5BKBBxpj6+9olPNOjI
PTq91WlV04axl6vtL0Pn5g80RBA6TY9QYSyxgjQp5Xa95qoU5dSGZjmpwB6Yq16aii8O/3W9lq0/
3Z9ZBQvdcM8Ll84akom7bNB/1wzjX3bCbpPFLWayqhFtVRHD41N0jW6mReu3yJKCxiKfeH9aLgnN
/4C2W/Vn4mANzqAZQkqPdQGzeoGWNQQByAib65naH7gRNErXKAUeuxIiwiUqrZaxK1V+FakVTE8c
GzIyyIxpP7pgnVd2MQJs9gGmkJt7h4QW968aNmxh14md+2rG20Ba222CC6qS2oYpyKW3bt+s9wtE
ua6am21ygCLEZdqin1z+68GZ+mZxD2TVSra+B1cUdrqU6fuC2qYDkJsTSlC/UgD40DFfn+dstOyp
rcCaZz52enU6zBi52rTxf+rlt+GpqyJgoIdOOAyIBNPo0ua/zPYGrAlo9IUvYHTUcTCGsGa1uzej
bcYTiZDg5zO2CtOX4n4o9iT4wkYiZZ09dahjJFz9B8Yb9jmNru2YD+39o1YSLIrviIdlKBnTh+6r
nJbFZJxLSwrf2UxTF1Kw0I6Zep7Sky3IgUa+YpK6Ur6rQOjIyvjktti4BzYZE9ZIW6lMMWjpJ3WT
8PikFqg/AaW1W82j8LjWLEp7s+vn+8oOKsZXqKqptFCQuN8QMH9KknOYN4b9KADmzyVEOVgAtWbG
mgPSYNM7RlX0jf2oGvZt0jNDKQx1yI3X1+2O7ELco5jntsdFOdMZEx6cF4FMh0klDCUaUboeLHo/
WVH+ml2GYsGRG7BTn7khg9T/7uhVCFRenhO92neDY3/4m4jga2847Dl48B/njslO0TTR8Vhb8baJ
olmUe2C8eIRR5zubw2dE4z9QKTIrUyrhp29SvReOWAEt3x8/2BquObb+EfWTWFCtGEnHxX7KjQQ+
yw8xn+MwZSAlIUdDKr5bjEUoF1+G92+n4UUoLhozw4QVJXl7IPaZ7WPORWRuIANs6AC+QSDfdbDl
sjKXsbFq9mtdzQfxsaBZfGQJZh7MmFcZnyrn3qm1z0ILEGc/tjM9RSpbRl6gjV23ZTlTMfODaABA
tyD83ys984Iq/m7G+7rnywS7anGuf66qMQmTGp2u+1EZqGez4Li2ep02Zu3bL41WvsDtdKe0RSrg
XEvayCfaLfj+HIpdGAQFHFaAhi8MckuuVbwXhBwCVnXwo5sIXwguBSbqRji+i/bNurCrW3IFiArf
9UdnwpC7GFFcKrLMadCchmGyl11hJYtYIvRjSoOgVt38Hh393p4KHrM3r6R4aktupXGlXfu+jVS+
u118RCyzQ4a6/mAUCoi+fXaIJlBDL0WBuaLBGEn0EXq42PGfzD2Gb/gomAiQjnUPZR+hcX9ECd2X
ShzMXipXq4W8xgpiEh1iZdHuI79xfDQJJNwhI6ofNnnD4iCWbphD58jNIo6CzxDeiT9RZIiJSunh
kj88XplYOEq5Gmd/v20NEhZxUKHDF/B/spkWIZ80GlnB0KINeAEniBjXkPfim60ZD+wzXl9jFtpR
ClGHielhFmEgJzs8Vrw1XKd9pDCh420hTb7PNl6agPw3ZH5R0/eHtiCXwQ0hfiCotg3oumvXOraz
9NxaF8zwJdSQ1TNm+kHSX0qx4vEubvXs9/udqsrIfLo1Pa3T1wF4kWBXEtZ+ATxXeUt2YzEiv0yX
vm8IF+xXFr1SngFtxxoRRirn1rcKUURPbs29I2wd4gk4yap/32f3roKxXw6iS9Lxb0so7sENiKIO
VVuDdB/Qfb1KCtc3vTblpSik8U+6qLManP0WoAx2cUyl49UnZe0aAsDX5ZNkwFHzSYLGCw8rS01u
Pe2KszXfiHqMCkJDpk/6Mnbor+BtO18Q6RF33Km5sFDYyEI3u1SKsL0/NAelOrtjOXk9ukSVCYwR
RpHgpI2MpfBm28t9c0VLafexlcs3Z9AWkF3po4b0iVsIhYQ/wQt3Ky5Kx2Q+kMk0aiTn/FAtPRa0
oq+EcpQUoYHBg9vfdY/dTnrD6tZ9KOdjs4vIbgomo8SqzCOqqUWMfzHvvniw6aUPjeW4NkFAmWz9
u/fOnRKCYaAwruGaZSnu2jkEJvqYa7+SqqrUP/z3ntdz7WL72UnCEMpNEy48kglc+d3+wgK0kHU8
hstxg+H4MVtlqQHsCdA/6AYCwAw4+P86PwmlaCAcZ6Eo15yYvsSTgA59Q8byT2c81Z3qjWNFfWQ4
f1yBL0qGeOjXBDNTpdtmfDcc+D4O2w8bdysf68Z+fIqcrDk/rA5UrkK1UfOCg5DrdD3GHgleuJe5
N4nl5Hq80vHOwrQ3i+exH0XSI8Qo+pLtzLtn76QNaf0QGuPD3ADn6prh+XUMNmUO6U8PLep27GLc
Wj8wzubqbCAyVm19wnKNc+wCu1PidEWzbbpdQQUi0DNbW1iYhwqDm+XxJDxVuoP8WtzSSpxRECcR
t67ZucfRmQBY5k/o/2ACD/KLFHBOEHHc2PXeJQi17DPsjxe9d8OUd4tv0Hz8VgK8V15k+A9adcC6
W9jUv6q1JnIhSGP8m2Z5JiOsvNDFWrbhy5ToctgP7AJG+SWXLPcl03ZtoZxvsPueJ13CKuV2Lr8C
vCUDbxpYX6ed8Ehb/aA3PEwaTLMQ7LE903Y4RoYhziwc4YdGrCuGmKpHRe/eECt5vq+uDodTvRQh
hwKdZ6Wwd8nlHXga0U9BxKAzbWfMp1eq8QBTsLe3uB+z1d4tlwbX3+0VRpEJd1tXTm4xJSZqP86Z
2Z1el3CQJDKHOgSvqRu3fniFR51Gtuqb9403WJcjXq58UOI/TA4mdOXnwXK95mm+TDVwSDdv+I9n
J07wkszJeg+MpZtAfK5eO5gadLVfT2vTBS9bUrc6UgYUchQwDYGBTvoXAKnGJ4gpkKgMfqT0PjGe
6vZZ0U9SPLkTBdOVDsx1v2xhd7l4Q2198Ntl83yP8GAJaQHGi7E85uQQoABRB1s622cBSr3hZ2g9
KjQex0YlU/dokjpexmAk3EsjPvtqKqmuYXW6dkmyeQ/OITOtaZVM/8BMCPxVhkVtmncqHzmSMj2s
vCC/4z1Fqe89orH+1oxX05sQJdI6zI0eWexLe3sl718TadWbnSxGz/3633ImVsiNRgiW1SSb1Xut
5I9g744ecxpiEWTDL5W325l2i0oxXGPQ2P7IiKWdLZxt8mJYbtIVJuPkGca4HOYuuLYLP0/UOKWA
dlC9xsVASuI/9No/uTp1mkYXxfIPSN4GNYF9wMLlQGzJs+rL+OWjMU5CYVq29MblCv1TBr5acuZ+
NlZoF21ziNALguyNPPitSv9SzHxpCuo91ENu05vbBYg3osGaztkR9AalceepGS3YfxTW22FIxrHO
+04W+1bZvsE4iSdaCot7VssbvGm19SijByJs2Hxdtm8JOlwYGkMyLqAIFBUXx0DAnj82xa24oYUn
bvO3F2ztFwS++QIJ0x4wOsgGzEGW14fMZNm2jqN0fCxbiRMXtxweMMrQF6ZfHrRAzs103aBMjUv1
E+BnmCuot8sWwZr1/2+l+MlHhWbb1KcVXTimIizs5i5lo5sOxBtn8EHtpUDCu6Wh1t67LYnzBzR+
DQFx7GoG28lnF1Rnqi36VZkDlAI9h3uceH6EzXFkykyTEELx7k0TEQOSeccldl5TPWp4mu83VRkn
udm2dvxTNEUYcaclotDCVBfxIKhNjWwOFCZ48agLyRayD982wRlAcJIW5o8W99XJ5UHvrVtOm47i
d63Im6RYj8ia601KQItQwq73viKffF3gJ+0upGq+hI47V714Ey9imyJP4Ce6H7ZT/wTL+pl3LIjp
iRJW0VVjxXDb1Or3hvbh/CHiL4sCZgYJfGh1HT1O9aXx0kpx3wrgW5Ya3YmB2tDsZS/B3dlwZEy5
t3YT/GiwUMevgv/c4BR24SFkLQxyryUndPycsxbvzoGVqycWOL7BIPI2UHL6nrWBRSVZIDJ8YTJ8
M9e1uSNdjBWDgohiklFN8K57hNg1pRjscVDjCDx6PmQ7+srlN0mS+TpiWd7SwBzBVjDF6g8ZcKnc
vQz2LeBCow42psdv5y44esZl1jYaUOU1VYp1f7BUVKySl335m/MbnHB33Owr8yHdINw8Km6KGIEd
Prau9iH+Ueia/++pV80eZZ0znTTWUj3aG+1v8jeQXOactUl1U77ingXZVm61gPwaNGVk90iDETtC
kYQjy1gUoi7H0vL+95oOhkOuELiao+fXM3QaLEUkjMkzLJ2Y29JVGnAvgCI+rEadh0HDLVycoX8S
ZX7LXPqHc6UOVSsc5qljIXDcC0cqyM4X6xi/jCUdz2A740Tp8q08a9cotjUDVayjVVr7xJvs4uat
p/upjR1rmJRJMcbxrIKtIrz8p97CecMmWICJ+CoLzzpkwxbzU2q5qEsArDRSi4gpJwXpM/IpCfpA
C5iVlYP+mAHX1vOWiv134Vwsx9U0NiajXq1XzIH2CBKBJGXa3oMRdRkVWYRT21bunbkjye1nssry
UWEqbZsw4BXLU9nfGwbvpH7UWBkTPt0uulI2KJy8FH6dFTMi4wcs5IBPNFjaPyYYE5r5qwlhipA3
+R/P+2QQIxkduMVmll9hPzYc4MlxH69mgT6iIP6ja1XnEwhERZTAmDy2M2j+yNMKARjYBXAbFdA7
TZws9misd5EFwgW27dlZqWG++o512g/pXzDejMPazluoaVYAdsY+0xvtky+jVxCT3HjK0sjFxZFv
9RgatD/+F8kl/0Fyf9I8VYKA7rkKsrp+mb1fSjJnEgEIuYdvzefR84rh4piBj6vq/3AGas2Fkjne
IzrVhcQnPD64lyjmg6/q8tRvH1rLLWjVRfDummLMAWaDS4ChcbQMJU51gBLuK1rdsrb4TwVxDkgX
ZMQ1Psj2wizD/a2xW+e7db6YTe9fz5EtlMCzvMJbafR+1isF3yEKQ2rjxPMjiRjvFvXl/dh52N16
HtOL7yZ2RwgZKsLiw29javQihSPL+mrKSg2ZD8pE+Hi13l3n/a0sTDWzUdTN9TMSU8vIXkZY5c8w
pO5svsSuiFRFVUhTX4etCmpBjAUBjnxDNxrn0RCRQQ2FditP/LWWSdpyRKN8RVYyodwmXrXdkbhz
k6+Ax/rkd3VqZKfoErz+mrqcWJwcUoRyyYp4xcHc7VkaUNy+aSW7Kk7Vk2gPyeY9dTjPbMDesE4b
evCHBLVP2iSlztWhbyGMPIlnJwPRAucaywhlZzJX4BxH0KSK1eg3hcTedoRXNOdL9R51PVld16HM
8LXjxPN3aH72j4sHpw3H5BKflyEDdIRFTXFcLKCEVkLKmpoTQdvtokq64FNPUu+jvDxlT6KKE/nZ
G38GJWcRYUqGksvmR2FOmF0/bTpArZhx02q5ic3n4kmAKmFHis6WS9+IZzGcta5Ksj1mVlCtIw7h
LNxFzyoxHTSzTOeB/KVLkwkydaNHPKkPDtZLatbPF5hf0D+5eoekku+bYUZyY5zv4zOISIDVWvy6
HJ9sq2wSrs0o8vm3NDq+Utiy6PJt0z47mlurwHues7/gCIWi70lrKz1oPU5TjtPa9bhwsdIqulKp
i8T1Di+DM9IeFB/oKPY45FzHWJnad5r6SPiafI4w6ha9xhVTICHzVDrc0XG+pC7UQxk6wCV61WNK
8oncDHCXuCUUIG8+zDVT0DP2j2YBtW6xuYAX4gJ8cHkaeV+utU9UX0jA25VRVZUHOXJyfFWztiL0
wSKwwWKft9C2nOXKpF564xTjfAfBTAxRfSaoJEiqrFb/mBhwqwolJkAZLAuEDvwJm1MhJ36I9hct
d+We772scneWRRWPSm1Zf12aq5gWCGgJrdmTlIz26+ZHj6YAciHy/CAMwfxWkvqNRXZlQhuvOfaW
w+D+I2n8j+0+MJD9H67/u+XRzs2nFYYce75r+ZKb71tppl5B+AviCWJtqlZNLeZjkWIxfVhiO5tQ
hoygsgAr0sPqXeThqhw/jRgwOON1nlurv9KuLRV5EIKB409VucXOC/G5w0/NbwlyAfJ268qTN4k+
+1CS9B36oJtC31p53+KBe4R/fHR7OhUyBa7j11E3ky4bSbHQgFsIX14LmRZn/NIAVq3DzU5kHe8+
XdjrTovaifbha7sKzpgCcSiw2/eabr+JzzcIRMoi9FyeCSXoqkXbQzTjj5uG5WKCw+Xr+QCM9i8E
Cbr9GUJk3pZHym5MLpxZcpMiS6j4Z91etcBWNWcYk3Xsht/1dhvl+o5DQqDJcXPRFd7vzxLf1LB5
4CcW5tl5J6t64ZIbdyeFratNDBQAGVtvcWQju4jqHQBaeaIS6wXxg5xcH7IqTndmIM24fe+ZZfZ/
OQFwF41UuR4IsJbpwD5FEZGLIrdvv0xO6UHrliqZEF6ir6yx7+gfR7BIZximuqvfZkJGXoI/UF/d
Ea53LetBSRsE45W8VoJAgGFjfDlgBL/ziZcWHYyUuC701z5lRFh7o2N/9R+XqXFBLnFrud394+3/
50fGU0LAFgpJ8uNt+ptj+c7ZH4xl1vxL/4QlQGQA0ux4V0ciHyA3tdBACNnYLoygwoqNFRLzlWE6
ACsu1xfNE5nqtkkBxEPdyMxF3TF4C6zq+8UX0ZJlxG1PukYhAZUkGOy3LNmTSSm02Epqsw+aw170
/VHN7tIAB+nmHMcpdEMo0gk3HsHclK2d5kPzjVVr1zPvk6tf2gzK66lK/OAWuSIyHzVrhzi5qmgv
y/GJxJL9O2LDNnOd7LQCbwF8RIMDm2b8Tx/mmCJU3pvHnKu4V6lnJFQQWY6s/BFBo+flFxoeDsUh
/t0sRVWIWNho69BJ8aAbm6e3EU1L5qU75+mWudptQY2Souzlf9EByS1aiTTqDK7H34uXMTEtZ5Dt
tD8UPERvhiEDtkGt3gt8ROb/P3t0xZs8yHr1RUSUD23sSyafj2X/mpl2A2OJNaEKuwkL6x5PrEM6
AY5xrS2hgTYUz7YZ2fEUgkdewUNZ8v5G6OX3AtTw5gWpPYmjLF0dq8mpEdT5YrfRLLeTdL1TWDN2
OaQVPHNSaXw6mr7Z/Mwi6jL92Faw6HboBT2FUBF0tVZJpCHgLG1M6nXn+a3FN6Wwj32sCc6GfRuV
eszhid7puMMR0ecnJANsRjvXgtxfqGvrJnDYoPy1MocUtZZDLWNynQRjk5EC6yVVOmrazMSxiOFG
+t1wruOiS2xXw96UkQjgDGZIW85aNq23K7ZCM1Vd2Pp4dwA5MMKU3vFpFt5df1wnNQu7FwLfz4nk
0lQCSr7GicchbOJ/BMgIlDn6n2ZYgGbur86GALM1rDRISFshtKrvOqg2uMcD0Ps8D8eq67Fam5dU
Nbmu+ta/CSdBLLlEZ9iN+1B8qrdxdmZ+EZ6E82A6aIaZoqZcXDQRpo4Y3UJT7NhCX0DMnLM21zB6
0jHo6QxftWLQ9j3Fv99w4SpevQzq2Bwms28ZwmuEDtnpjPcZM1X+DHduHT/pp1Pt/UZht9bLu3J+
DF4rODZzz6NGYh2mrqqpwcQxqYc2NZUw5todtpF7nRVGiIn2Zt7HKXmbUvKbz+1HZyufWkU4Hv8a
1J5sAQ1eLOFutIFg0IXBU7GB/UUlbQ2ImtAzoW1MHgHAVQxcOk3DXbNeE2UsREkWYNeSWAvz04AQ
zJCiFApTxISmZvnAPn46fU/2kmDnszJ0umc2FHoV2c0wogKKzD0xKKP8wsqoMoPKUQd6WT/EqXGP
U6+03h95Fc+n1GWnu+JrELBtcUh7kPznwjPuS1c1pgVXxoucWDr65hI3JYDu+i8XCdMg5pT0bWTm
cyACd/aChriTmkD+yKu3QnZKAf4Gf2b2LefIdbdwg49ecDEyy6bs6poQAVeuvvuJCoculTXGmNzf
tPAJaJZfCLjoC7qqZXfIX04aGn6wYikUwND1EhHfFu6Sao5uhaZDBf8ShRxy1HSBQsPpo5ncQTD8
+7uGEgD5RYenFWh78ubQt9H/NVdEClnUWYhgoBJS+EYz6VSmfp9GUWkUoUz06Nn7Sdmjra8Tfegx
QDDyWaCr/Zn+QHwRkYUXbkOlwCGvJ9a3ymdx1u9TfAWjEmfXd1tFPGaPydXud5Tp3nZjwpeaO/fI
kC4kjbIujmNS7s0FvvBQJzVFZOCIrhyqh6aK1Q91lTZvf65MV5GfK37K9yNhS578klmMUJKpmYBt
dO2npwwM93lT6ju0ZqlbIw474qz0qgQME06GgUbdCsxpHpnN5ja4NZliSqx7Np34HwQ3eszduYyZ
6y8TgfyF2ROLUbT2Sxaa/KFpEzCYNxHGpIK7Ao0ryioQtwXi0Ng8vHZ/bU2ouYM/2+jjTqausaV1
AJ1GAbAtmBH4z4t9TA6BQPKF20ypU1sbFTi+Z1zOG2LzrZT2TkSpSOV1lZg6ZSM4D7xn1W2+na02
rtE+MmzpsMSMLABhwWMsDnZXXio44kxmRRh6u24jVrkczSXvRZ55rxCbj+/1KDlLObdpTnbc1oCk
fjZ4cE2mkQiQwHd0htQLDilMjdxd79mj4V1X3Y+x2+niD4kQaw9sRBdAHpVDiDu24wBxXM7PCyve
5tpRH3UdQ262U1b5W6gpmoi8WblHFyKj783oTLpPxH08RlKJOD3cEtZH0NDmreMYJOgLylBrf5IL
Bf+ng+OABTt4VmnM+joZvHyialcTzvKYEknFoyC/vS1A/SnkSzk5oHzVIuvhwnNaIxQsZ/E+coB6
x5hq1MySPx20MMDwOXucGZ7FpZGsio/JFjWGGh8ZG+VLvfIEizU9e7H4VSNv0fqsLgTn4N2OoygW
385+J7x3bWgXJRlqvSBrXKz3fDz9oIE2gHan8tIBtqMauxRk+B+2T3ka9AIzSTXvR+Gn4/E3NNh/
kSKgAvYyo7As4WIu8WmDobh+GVsRgEn57LFslaHSWJSwHtQvKfD78pr90V0f8A8Zm+4tHS5PVGpQ
+6we1oCXqXuvpc2WRsjJFSwx3N5zDMBXgoCOq0VBdshPF8dBN8bAE6RQIEC17Fs9aq8KVZGTyRJY
14XEN1O6wUmunSJO+WaSv+c/EYdGk8JNhCDoGoDU2p4QJ0xXdvF62TxBtp0tsHB+asg336sTmW5D
w3BzRhePI0Nzzr1Pt/6PyTF82Hap71N3mxG8XKHUrUhcMUM94cZYs/motjZHoo8uRV9GGJCBHGIS
87XFr3rFfVL89muD4lvRDkXKdd72tNKQYfPXFWNCgls+viPiTjOwPpvA2HdRwCRBLeL4echRIovA
HUDsUC95BpeOE+zIW9ZytgoBOp3kCQ1+qY3QKikv5MULLE/d5RJDlSF7ulV5Wd82cuhuE6zvIPgs
lrW1219FuxK3FeXi2cFZ6Roe4vbRkLxVyhmVoPZ5mICJkCgVJWpxgCeEx40a7nVt84mdRExqy5WX
79L0kj1+l05nWLT7rgzBrjWXblwTwosa1ktRhrOivxystrWJHNJwCf9Ho3NdHdV0XrFLiZESzQGs
mu1mlC/vFUgYkmHEwEyHWQuh+TZu4NkzMqQY85mrYXrxXExzMeHXoNCiuMmU0LKCKffnTS7GBbXg
ngyGd3Pqkl6SOykGyi5B46xQ6wpSKzygj2Fk7s+YNq4/wbjDZ/VhP6q9sH/4Tig/QAxA7uW8vzIV
by/K+deeHYTZHXLiOCvSJ1uTDC+9cNuSy20bkO9UhJJsNB1622HIA1302Wwc0MuzGe3TkBRGHeqk
B7lBfWOi/mJ8vI6Y2gdXbYy78zBol1aJP3Rm8HxfbWlbzWB5D9EudUNi/efkUjyxVG/Huv0x5WD/
FsLgvdCPLnVdc9cVPtbn+eHbYKvgD8Ebe9S4mEbS1S1QQ2yCXY2Fvj/SiwwRZiz2RsN6tD78dboA
HU2oYLfTFD5KyyNaOwD2DRNwGISf882llK323lE1ebLp41jBgeHqmzARaPchmS585NhIgXFi9B7g
I+tZVAGNdqmcG+m5adFxFy+YmKwykKvlqRUciH1Se333HICiNyEUKXx0uekI/ySdu2pOkImQsXOq
282c/EKRYIsK/BYqMvSvVH8BNuFB6Fcj9u51m2qOofuEYX1nLWR/w7hY/4oQ7CNXzDBXiTtrTMjA
eP6a1By4PnGdUvRlaLHQPNnPOp8TOUErCaVcsdg82Bpu7p9Q2VNzLrEtR3Dgg9buZ2l21bnFopvm
u6wXi4SJ7lK6j/IKfT1QGA3t88LkhmNXnna/tLPh73iiyHabphIbykswjIpcdDf7CI743SMopJ+D
7QvJ0UefYa7I3CRmQGy7uZtD17q9IvdQq2OmfK98GfrcEDF3GqqrxSTr8cLToXPuXZsczityqYQn
dRxXzj1LuzDOi3TcxMLjUI5aHjsQHtyVjOewIW7qLYnkStqhdXl1xCiMmRRBGWQeYO6lWtM/K25y
3nF0hYDIQAa7Ozfjn1QdR4IUOOPmoX8ABQyx5G0yYVJIMORwJpKmYjTrYyeoR1cGuODkIM9cwQ4A
kOODUerETbQcpF8VrTsbotS6FzTmibriHyzpGce3dh8NtirSG6nHcxE77K4A9hygH5OGhziPr8AR
EH1sppHi6FrgAAl+5nSKGqQqGjEu2KBlAK9r5su2Gx4P0U7j5n82Vi6tzgnZyMEWIS2k1UwWYabK
qvShBtUFbr6yeswZ/b224nE0FEmxAz5gn7cnra5fCrcR+5YgBN4NQ+B45DFJLDRZTcrqeImy7/gg
C8NObkErdhnWLlgXQh3ANGXGEIxVaBSEMyAzmaFxP/4v6n2qY1w3BEI6clTZarhYPSN3as2TV+G1
gYUsan++jJezSHK9N7U2Dh7DiWzldHMp5dvsLceujME77p6q/lBZsd77s1dkFQv6Kizv6gMW3I5j
FWDwDT+AmqqRXHYI6pJfZpBhbCqf2aAMfJEFSv7tQ9f+4PJC/DeRON+GonHpJdOqIIvZwyHeicjT
NMu9OesAlKHqUQGL1WEwo9N3Qm6OwRe2UarIOypGCvUrwhiNwyAQB8xltpWSKm/F8ARJLBl6lQOa
i3M2Is5Lo14baECIpDpTmhvQp6otL9uEWbtmmoKvjO6GekcxSXPbw9ytnZNT5kCks7B7UpXTiI8s
NAtYxoejen3E9SE1Q414/EJjtAup9StVytYhzcPDwUrA3UvHqrvOem5X3p0ZpjrNT4vkZixg0xRV
y0hQY/Pe73UUSFQ4lBLyvuN0EvFZ1cwaEz/EO/eQJ4rBwE+bZk/T2NrXsGeY3ExKhi+K+0kXG86h
X0o2EFFPOkt+0BUNGczbMqoZeedCuW9IGmXmi8dx5/hxjZANGfDtyzkLOj/xqHR8Ne0Q2y2a9D+s
Fu2QX+0fT+pZDBwGSdxXEEkOGHyzWZ4XhdeISuOYk2T+CDdPHPVZMnn2ddJzPeVTP0Mtfl436cl+
FSlf0HE9qxIkBJgmT/Af7kyrYbNU2+pC5is72rBkLGsyookKd/QaehCsgRClFMUv6v4QPRpnoQds
je/Mh7oF3arSMEFaCi+c9QcqntGrxSNcMvQN5gDTFDr+DnxcCLZKjo/4LRP6axoxB+2OGXJ10694
k5A/Q/lOkH2ZTKDuFjZ6c9uOpDQhnMSg6wn/0bRGCF0a1qgxgO882mpPNyu6RbXM46J2af8DywsM
Xh4CIvCNvpSH660yXLS0JLVS4u4i1B2fOhakVGsswU+SxBTyXgyPfA/cY/mlI/tYcq8DbCQ9E5y5
ohEDzpqKoVo/L5wCiH7U9TWQbgCl1Pu5S1G+nRUJEe6y1jCk50wq+7ov0g354Tpv0wf+4M9DE0oP
+ClvurAFncTWD56YOSaS4Yh5wyX4zLnbk8Die+b/ix98Mczfh7p3VoipWUgWAmxQVgYyia5Lyioa
uWh3sRdUbPeZqx3miKFkEscjU8PizSTRB9rdFKzmQYMUxxJiVsCMiNf1hPvK5TL/Cb1goLPf06c2
CHUgMcCwZLTcIXtl78Bxy96idrpVuVPtbSda3TNieaOX9pTz2LWGt2kQTBmcw5Mr4DvZjwlIQVzt
uGBl/C+ypnwwzZjz3U8RXj7kDqhclf5mIC+YHVKClOIaxaaOCPTydAbKVI1YFOJNtAy5OmGfa2Z9
RGrP5Vd+gh9OsXZKpK4zlnW+OnBr07jDBzsJkZvCFNCw7TNwZMJbDInlf75HhE0OwsqDdNtRBq8X
AC6QQz2R1TIF4M5p8T1M/TipTkZsclbCDpxB9cUAS13wxWvq3S4WswK87Yz2C76T0J3QtQehDnP0
NwFv1YV+WdEgvwJx18SBfqRnzEADvbsHFPoVKGUfo91qlmS2xFxqFnwmaNiBRgDZXB6+0dHfLW/E
ymPfAHxZ6V3rLAwdjhWNEOtLj0eJCwmhr93ebWNDysN+jcN7LTgJ3EZNzR1P3JuTcO5liU8jdePG
HeDmPVkqdvPy9oXHB+BcAnBDqTdyarho1uRGwQtrHrG9rJ95yio0qHWiS2b6C/vm27R+v45vHlWx
zroYKqbbidCgTcZRoy/stQYlauQPEWz/pbJOkGZtLpDIbacrn+NSAwyBy9K90YSaSC6D/JLHoBQz
VPRdKPF071on7ezh0+OysQNv8FLSJrAadgCkdHLBZ2Kpm4QVTbqmGT5MUNdWBtA+RdhOMPbXL1Sw
Bz9rroFXvnxLoRYkbvJoUYicW93ZxcaibIz4ThlFVkEbRJtn/iZYRvnmatviu9ATfeL0m3iKD3ZE
AnIGrEEHWk1XkKq6d230XXrKpKEgJPjkzZnC95sGZLXiW8ZPeQe01yn0q3UtN94Cdt9m47xAKsE4
JHkn+lP2E9BCgz0Pw+zz6Jp38NViSZua0po1r+Scxz773x/EsQJF+HihzSt/V0uClhMomakIHVKe
YNvdxZlZFwS3jpnE9lPBYmH88EDwgnRgUs0KEiv1nKYz+4D8m92kfQcRPz+Hq8mOB04Ks1K1LPPN
34UYWg7rgk/znETbEoeBVLs9aD9FZ9NEHAdLGH9eO8FV2/XBIg0GCglx3zDNYO62DvJ666qe/K9b
daUO9RsTVL12W2rxtpcc0tldt8SvPNubfP/tjuFu6CqhvfOCU9CMacznfPC35cdEaOFZlDvz//qn
x0iZmXbqEwvTmtbhBB4pm8LrN3NTcqcM1cBlF6W4qULWZ/p2jqyaW9xomsUIS2pNrScSic3reugs
86T570WE4t3CcfGcrRYtkWbkPUL4R7Q+PchKYWoaZ3JnG4lkZg7TNCiAFLy5QDQml0UcjKIPxJiH
+4+7CvrqasjMFCpsEiLLg5qkDor2ClrHvICiffCx4zXDYIn5g665jvqpywmwGgUm/kG5Q3QzFNgp
HOgls+64LHhrxIcGNVcMsI/+x+58jdlWykOk+kqJ6hsje2FiKuiOrB3OnWzMYerw+awPvaNmIBV6
WxdZT1FwEpEuoe+MVNn0jiMdDSR7bEHZ/ufedgBKVSkxZd99LPMw6Pmcyy8tL4x8ZEfEoAFSydz1
dnMA1Rp2RPE2kCNkg51mQIJ1lj/eLgBXiqET8vBKxAs4hZxWsnDoXvhBD0YzWPOnpcDYqsR9nef7
k4SOgjYrmy7P7yYgeBkHCm8uoWjRrUi9Nw5LZZqaxgtoSxuSKeueOkGqvN99/vvCsPPeXBbgiVH9
96SEljYuJmOEYS/dxzoH6r6k2sj3kZJgzL7cSSDZUHsUjupOTwYYfdUDdhYDbEhjJnn4wRhyjmug
g5ulgpzxZwxIqeOrVE7X8aCfoJV7AN14ubgj1kASNl9Xv68sFG/Eiwju59CJSJV/zFB4E2+3lWin
rJ8Pz5h1l5wvR0x+Q47VomxxwNj92aLyg9yJNEjcA8pTtnUWP6DgsDiK9f2XXigRDYrTYCOi50WA
tQKs/5MsCMpas17RodZDntUkvSQSdQ9KWoVxGR6UqT33xqmna0dshoS+Ny8z7nvMy4+ACIIOEPJA
wjj7BFPthNT94WPkLCNTmXpL+bmErpY546dAQ1kh98Y237kFJzOdGMgz/m58ShIwx7LDEF4OZysP
7EYQ22IlKAaY+GR/CwHG+MOcigWdJ4J0TB6mJeQtYNqlHsTNyncfHisCEOyZCUlZFB41DK+L4Sdi
UzfEqX/YsaaVqovUr2EdeBTOIpqRlu4TBjGxVCVwKEuxtDHKw3Dt7sBeHgioLHcjjeMkT3+vrZMs
v/6rf+g26h8qJ179K1JGzfOkQHpaq8R7FbWlcnDMpV1RBEX21bOypYAUNqH08DjctvgsD8as+pL8
Wy9ey79bIkie1CXUPxF5BZZ/ga8SDBtSOb9SOmiwtLaq6X9hQa18QsGhG6ptY5tws/zQArIRdzEA
wonEE1xYBcXaOI7LlmnLy9eBZRvpiLWZ6jdlUfPsGrUpK7ZMNWtWyDfkCU8VsIytnV0cMD7RCFeA
jQtLDYT/vFYXOLBp7QBoGyIcXmmbM5GlYVLVFRz0+ozgO83Q5at8reFFxfuvXdAM1ZGbtdrIQviu
NVILxamKDACSSZGKf9J5ix4ZMUPF82Ct5b/6fSaEyocJ+t6hUhta/ujZTNU6Bvztgc/XfySvZImz
ENIKTPPmJ4wi2sQL/uVZ+OLQifuxjM+D6wD3jXWGd09tsb+1B+SmwakclTsBdvasGodE/iqJB3nL
fV7YUv1CZR3nfoU1QrjpMx8WwdJwaaG890h3pJ1NTbmmByUHHcuhPvF/JV5xPcjXo9mVBQM3jX2v
Fm/bagmMgY26HyTiToWyU1yJedmQWazBvaPEYzKaP7vM4np/ovO98WcoIHcJitJk3VNVptNwjpNR
3tJ2g/r2cv54Rxnh4yDZ1RP9Cf6e5I8IIlBocyv85w1agDFIFYzclQCChNTKJ967SXJXLfIECKP8
GwC3TXabGZyMAPWWrej7TGXciM9VVE6PUuZp5Cjj2rFBV3rWUsJcDozmme1zYfQmklNsNxdX18iK
PVpPVdnvGOsH+OJ0F/xFIOn6ttLMyg3l6nwy2kVYOIoCnDclBjBFRLsW9mtZJkexl6O8Ilaybzwy
/qyPtu/qkZBwMJCkIMgrHiPjgnV5YZG+xxl3Ci2bxKgWvHeANiTOS/v2kuIJzhZtoaCuen5jJmIg
qnO2ltvv9+PQYNh/tSTSoFGGojX1YBGQ7WD/yLCWixlXOS0LlO9vHkFlMjGocZ/AXu+I1l9KIjFK
bSwa0A4UJbMKfp1huU2NvARJUqcSG1f0qcSM6OYKcwen2eaYAcyoYhEvk6cuk4pQd07XPAYEy8Da
Ffs5f/X/LjD5ObhKq8WHn7Lpa1HZZz8mLGer6NL3y35O/240a0sC4KTgvMv3Iq6rkn1kfScatfGv
nOyqJYN2tg22WAUIeQ0BHtYHGXvDHfWaUEYibScIhIl3ki06iD1c6NJCxyBXK6MrwgFCPin58vyw
ziP4XB+/A3c5qrJ5CJjEPmJkGhIsI4lVeIZNxQW6Ob9fdbGP2d2EXzP0TRREm6CKPZeXOiNQU2mE
+n62ti29pLI+Qr0Or10pFo7ePaArylbU8RvP/lRHm9LvtsfYreLBPBYLg4YPX7LM993VY8uKypOw
7aPkBvTnme9iVdwN1TbXxwQiQW0CPGVFe/eiCnW10e752k/m3l25b3DCif5t21A8hJEOP6hJBzvV
SVCzfFa5REKzpAERqE2E5dFR69+Pg86RNXrBT2XLIujK1kqrVbbY4D+PgXPZOsdFwl2mQn/tkZxd
dYPOE2g9My/ofF7gu9OYdrWVD8t3MRPpymJvjqVucs+TUSBtwPBFIDF0Ze/YbA7g+/Lr2jbBPU9j
4t37iA2d6KDVnqt6/fSuYIgmH2aVZydDe1PJCwuSehT1DV6YcZUnE/nVDQr42cZWOnHf4fnCPVc0
sGANQE81Gl5ajISh1JBrRhbbtgsBWmO2yLY9Ika/feL/U7I24QeSQAQPEBvQy74wQ5/6xtyxrOqn
DrcdNlihhr4yGAfZ725KAlDbKXlAStefoIOdZIAGMPfVUZaf6sH3IhEARV/jrZj6Z2CsbXKhX2T0
eFh+Mq5c5u72ndT/iKf/PcaU65Sx0oanOmLoq+zP0jvxGgsbmGrRqg4pZoUkRV89mZFQdL2/h12R
B0GZyCRj+zKZT3lPlu6FAvK4c/HRbkxRTAaigQr3SraAsqD/Yh/KMoGdSlsX7ET/Dfe2+CoOpJV1
4ZExYsET7AOGrFqL0rSdcnK+DeFLIswZ1T+4mHD3kEnk9pLXmSbLx4IJHPXmCeN2aG8fGEVXxE1X
ZOpsFMBXQuI0jGfwS/CDQV5ImRxYEDZqHZzvn1MBHFmxbMfBAqDf/jo/9+x0tzB5TXRKiLIRn+21
mJMNgkMbl/Ue56zCtzdEjdcIdz0ksAQp4IvlO9Hk0xDv3zYxZIPy/M9+B0mftfTt06woquTHyO+W
oOW2b6TAAetgUxJmGxPcyi3s2fKIMX2isA1rWEVh85A+2fNRuJdEcVb3d1isY4Qz5oLy2xB2uPCT
jV4dDA79aPx57PJF7KZq6IYLIeKJC7oq5qyAzb9jFrvRVj2gReyj8RJLYhwFukZoTUyfYFX6xpex
N2cq6HssRTvDHzzUwbgK6ltajgoaqsNuHy/28Mwf8aRz1joEvz9A0N+bYyTwgh8dbNy+Z7lJ70zJ
ALwADFm7i2cSju8fM6II42cRGXQsYTRx8jMwcwNjyV0V6Myu+nBx9dBoQRZYAI+y7yKL2IegNbnl
NZfM3RxrfGWvjrJpx8a7lwNyirIGFzoDPNSxjxKLS1AEjnrzK8qyBTMB1FJdZlw+KrjjsbcMcRZq
FaiJwKvd82tG5DFh2GoxCPJYq94pyKBsEOy/RKve6URThOM7dbnVIFfggNKMhalxe1V9AsrajfsT
JfQV3Q3Y508BqZRn0X1TxqcsLZ+SyVVbEj/I5eRHemzylZh70OFp431zFrTwSRmoXlfKJ4xzelF7
jlkxMkMmgRGhSlyzk2dEVOvU4Ep8egQalfDHhOwcl7EfdKjC2twnzKpGLj1BroetXQzg+SOPBwS7
O2RjeGXot5d2dfpKCDAmsvooM0vYw4SFQt6vhb6zT792BAMWO3CHZu8WVf7SaKfH4r1aXl8/t2n8
rNA3172K8pDnlr3j1DcrzESfeY8l8NgvJsHA6jW0TiabKk+/fDwlFn+LO4QG3pD8MzD4q4f6Lqn3
kGBkz9dCspEyFXdkTD+4EYDaRsEje2cXqfRViWsPPanVdBViUle8xm/NhalhhtNTnpMaqD/X5gqc
HGTsjr4V479cHIvSGxetOEwAJg+L7wAGV3RbhXTo5W6GeFz/HIrI/iY2s5L8ijpTFT8TBeJSd6MM
ziiIExavM6Z92VtZPolHRWBxwAgEQUPE83ErA1e0H4G9D6C25znxr1hlsrxlCuYf7hGgdUWn7cQy
J9rYEVQmtMM8+kGjneXc9/M27tHihskLgedNidWPJ5UUtnAiEBR4bmvfVvd143RIvDNu7SVPZT9e
GqmXmcs7GR7rGy0CmYvjXyHvVUv4JlQDyYx3aGgxo6+U+1/FOhSgKKy/rcvC3zUygVffb1AlEfJz
Z+XW53aLQ5Lq6tVeT2TradVTGq4tAs6s8FmaCyrXiyI/hLcDXZeiZY8fVPGSIhE1qFRS74ax5YHG
JK+Nyb8YAYYa8cGc0DqhvKqTYpe2x11kKNCjC/X0jWbxe6ViXrZxX2/WGM4dk5mvXxFfrcsXA1Al
2SqnlOMDtFk1RXMb2Owy37XY7/pkshT5WhgAaVe5/9R38iAp8ccwiKaPtc0XsmyMls2HHgAN+eSa
nfKR5XOfeHpBv/oohdSrCWO8c6D3N4fuTD27PhfRKTRrG+KQN0IW4dO8SLwsayGQcmymsL920+lo
Gh9I+mReC3mnQtupLeDUz0vMPHyOx2JTOVg/znN1SR8H+z4XRWUL1qgeWE2rxzukqPx8VlTEG6ru
cv6zcxkKX30C1Hs1vOvfkGMjLSApBUlBrvByOCx7zueXFj3ZDKQizp+mj7kqQa38j2MMOXdnp5r/
obIbi5zggtUUGYmnHRDcjV7H8lugh9lKGPE+JEzC8szuCpVQx8WXsI9Rm0OU8bhd7rN2HnWmfJgc
iGVoxUy5X9hdX4/esZGaXZXuifNnkrI5y/ZxhneDIAph+iufDr4JWw24MtmKLoAvZNq/DHwsKnV1
q0IOLs8nsgNpHUPEQ6DupMmRBePVkQFtsBgiqJWSnc7rJWffQVkniTgy1SrVLHvQtqumREsS6Auu
vqQ3qYX4P42WQGapWiXMegj+vtWOm3ZNrKgkXwh3uHR+o2cMiZVvWFCtYGG0PlQPzF67M4j0SK+r
lmjGMHaIMraGIZvbhZJlnnh3tTs/zBppxp2+PpgwkihzJ7lBN8fHWFMZ3cU7N0n+/NXHd7TNfu6Q
4qChKfgvgon+Y5Ltq32a4SasQICVPuBc4YMJlm5QjlEtQRgRBkpJuINsxzYpItagXtBwgJ8O4tAo
kEhk2lyzxak00LP8SWyTxhUtaCI1YZNS8P3oUyGveXUQZrUKI0CI7Fj9Ctw8ESBgtvsFwqFiD2I4
9GkaRPysfYRmiAnsqQpuNTCt/0QiVM4EV483+SvvCqjYisYRXjVMiB42niWTgd2Q+U6TsIN/ia00
ymPVXeK1+fjbL0y/a2XVgYWsdQ0tgpDmfIXi6TZbKOuoNzSRbzj7NQqV23ld+uhjckmqfUJDs9HK
9nIda2g2tAtKRakQylcv/ygJEWjQ8wcPZCi0nX2XQTp5xel38twuaMsfYOjG3Iv9QhSdEAWM4w4B
U5toxW2qiZZ84Cx7Go3ihrEWuCRklOrVHOGyiPqZmTdw7AIwRYBF/JFvHKpNkjOpup7G1hx848+v
aKUwl8Q3hbYtRDno0ZnVtvB0v8izcI3VF2bobN93Og6Rzax3z7G+SqiEA3nku5tvAimXqJj7hKV1
tGBlZMyR1MB6f2Cu25wMba/hcYFL1p9wKIMeY5S2zsVbgkVRvWBEvDBJEZv8py9xZdc/3AFf6x+X
cMi9eRFREHlAXrwxGKvzvN7YTBCFbOArPTwXWV0gIVoOUL1jJW/9m8W+lbCI6qjRxw2Rh9xtKRbS
/0gB3Ti3NCS+3BsYSTM9MuX9Z/8E4rheaBl2ZZLRdQEJQhETV1MBOKUaOaqXn2JdVw5HMrhm/wLk
mFdOybfEfv8nCTOp8h4k/oBzO3iZEgAQkIUSegyltYbq8RdWjpHC27xMsYJ3q6tIC6BxJNpG8LI8
+cBcwF/khSSLQSQsRcniw+8ybo9FXYMh9ImUtS+DEGCv3FvT1OYYs6LH2kqNloT+RenkvmSo1PJl
c9rKaPRH5fpI/+/mCckEMxb5fi+Z3UbaFgdsAxMIEX790hg4+YgyMXsjjbCC5PfRxCqjoca3L1GK
fIA16IkfkDA4HVJ0hLsWyTNutL3T3WMj9CxvQbyQY3kNavSi5JUT1Ws/XlQGnggbg5WAPW7aLPBn
DVvuD0yxYXspvyZbUZeKM+Fc/Og8JqquXBprQV3BvTrSpTSdkyFZpvqYxAh4zjpoWcjcxKplDbRQ
RH6AlLQTxEDB8eJgAMhbMM8oj8e7ySIrO/5v6Hg3u6Po414GX7qxV7VOV7jHR9mgEl9SHnwWzfST
9J4og0oOaffI+FjOVylukun2Wwsge60jiYiIoul8Mbn9bwRY9OnN4n6lU965nZKYYRk9tC0Eg39T
YZriNXaR76nsPoDwoA+VHAxE/cbU/h1Iqz4IHWZfK2EOo4uFG0FBepwlnLe8HalOxJ/uemYOGmea
Yki1WjB/gswuwPkA7LSuXjDwVFYQfhipeYdwGuAIh6PDWTMaih1CXN4+TjoBNTaNYppzpkZKr6Ml
NWxRFnxWtcVXHmTwDCuDJfbQtqnLGnES8hk+odkHAmGBMMyerMbquCFXrkzBEt/98aJh5S0nwLmZ
+Acb7JJJA49Lqg2eURX+RfS8xyjU9+thTLR8vVx3VM3ZbC1rRp+IMmWickjJfg5BlAH6r+FBtS5/
IDgvYbowB1DRIRzPJiZYVClyBkZyIi6xIQsWiz2R8swUdehRRh++sItVZ2a04uBWX2CdPnF2r6Xb
Tc3U8zHR/SQ8fjeXfxcFrwDfEOMe3k0P37531y6LMpt3/oe2f2fZN5hKvFh9TrR+mFiIPAA4iV5X
c+xYOya2bVAXDDnnpXfmDQHrceSTpaQzj224qhB/v64+YUDZVsrr0KGQqMDH7JrTjn+NqBVvVOWD
DcNTHTxh5HTGillVkaPCFlyHdAn9bjl6lI8NgQn+fOUX2rdJVO/6K2myX27ZQL4Qih0vd29f0ga2
8YwhqTm+QzqGaxuckCuwGlc4qCCc5pdpIX2+Dzfxik1iLVdHwtBonl7a/GVJxpxwCmml9SqJWFhp
Cw0hJk1MrP5/MQ8+krjmUhUPRfJWzRazy7e9fpEuTzjyV2AkkJ+5cSpuidnrB4ZJ6iUrKXdgho+Y
uDKLtl4XK/G9m5Mrl9GKaXnAc5gqPkqWAy2S8BXFr7CRiNWupaDi0DawRHcYKczAzaRPJCFcKofH
UMgIfWHbGkiV2Gj7gMk/ASoqZtuT7u2Ai2/2T3PxJSNl0qDfvg2e3PDeuZAntDwKavcir8t1reP5
3sWP0NDOJ2awAFXYBhdqvzYzYngnhQk0rcP9nDMdp78yyJ6G2wW/NqnyBRevth4pQIaFouo9Pglg
ZxdC21atN8vUoUZsg5BCjgy2XN0KFXEplwLNks8S98z6FCGNZPKi4XUM421aa38G8RsPkR7KdWBC
oumtKYhCWHD98y1WFHSjAlaevA3YjhHB36Kxv+NkNsVbzU3Fc6DWkw+w4dNE6pntI6me8Ddpxp6/
l6FksxQV+niNCD2kUjP/s5XIzZ4HbF8MYMMKpNvSCGpuqVXB0TjfzkmGFIhTTPVzJW+P8u51+SKQ
ibcXzGh6GuasGLrgOhoMR4VDDPZtuopqaEAcgv/H73lcYZkaPDsNd52Yonc8v92GiNErj+PBsJJ2
R7UAocqFBXP9lQNpqbzbNd0n0R+BHdKcdKfTBg3JxtroCdkto4CbQwBK7dCjJjunEaWoFoUFWgL9
8j2e9JlR86ZcS5/QP+UElPr5EaULNjurBdZXp8S79gq/Q2s/Rk+YGH+l6HPFfW0tJp7ix+nmImQP
1i0VVGTx8o9uIs3g9b1cCpbxUCq1Vh3wax8/2iCeN9+LBG/KdHaxjpzB0bsTLCbnM9OeXso+goEj
tPwTrHOoKPv4TJSSoaGPd6/HQWD2wreQEMK4jIR9CNvgJhMAFSWegsu4GLCBR4jOe8RaRUD348z7
LNuneRnYu+D+FRoXx7bbvXFjMh1h6wIAhCf/MEs2Cu+orqXRpHjtFETqL6tSSiRNUvWJAs4+HhoP
1b3JeWsKzawAskuLXDLtA+Ed7gbHB3p54WysYtJGQXUv03zWv0UO1ztdXJVdzx2HnISiJqFJAcmZ
Kr3LSKpqdn4NrcTsNWj10Rw8JdSte93lBU6H5LveJZ1J8ZZDwEL64k4ygQlboEPlefeuJjbKOy7q
iCqiZ8PIfIgz5Q5Bisn3Zb1DkfnY+ebrfgkRoGeHEIiMzEXMh0M7IXrfOFxMyLJF6uHaGFS4McF/
w1D5uhvXeW4mW4R1Js71nd0XKOoc6gZUOdMpyLz7qK2W269eXjcTF1qfrFj6ghwLREvgvmSVLHmt
XD0sm29D9lD1Va/S7J/Ip/wQERJ3IlkGPu04W15yfDpMSG3L9hlRZ4WHaFjs7eoJdWacxHUpmYFS
1Wo0k6MREX774l5OiaZzNojxdQ6vny2O0MhqWGqZJ8U8Sth9Z3lN71siIFBk8G6kVEax39ol1H19
kwcAxoL64uwfhLwQe1AZ2bs5x0kvKx6ACp8XO94XRCEKK6bHD5u4aXag5BsePhoxUAq9wPr6rWov
2Nw/4OWq9bdQcss4vh9J/+bKMclBL8Bd6TsTsWMOIHO9riLfCLj77cIF1TUVHs2wREL5ToI1B4XC
tHk/X941H04w7NY/cqXfEupc5L2+2AzMoMfc7S236oys6b3FIZ23rXrJaJ6R0a6bOQ/1rOBWbVn0
5ahnC6rZY6wyIFe9LBfeaFnx6RAuOlNVRIRUWfqNjtYTFmktHJg6IhQr9gimPx4rIZAPsekV97bd
N9Z/rMKb4e5hDa6+LKiaj7nu/VZCZ3rCV07qD8Pf644SOvhHvQmkGt/BhqNrVWPTef0bypcjv+RC
5XQr6df8qnHV3qXOioFktm4gjMM24EZCn9rRo2zYR5XwWk2uPNgUWrFcnLUlkPTO6/FdwfGF/zCj
JVRNxumBpJGh4S1YHBPgEKBaLmqz9+rDye9a/a3WgWazhUyMdK/+Q0lWIvIeJ91DVw/elz/R48D9
v9hoqI/meLzRX/t4DyIHgUQEeaKEM7c+bWna0HMQkGFQ7TCMbPpTPefS7+ty4ljxhBH4kYHSTjCe
Ba94KJjKQl4FyLrj228DOLCKSpdrmiQ6akuJZFvEMs/2ros17IvSEAP/Ek+SlGUSYK3NpaZ+oNs3
8ILxjiu3FX931srIO1AHykC6BF6scQtDUrcwuqX6VrUP5kdAVGsR4Pp0hohk+CxsYqf210oag+IR
MlCLm7yW/Pmf6KB9zcDWmawbmOs4LBHml27loxN1QUzp3g89e6sa7xBBzc8iOP2DXWIaVLlafT94
IuawlK9AlP1RXllamAHpVcTz7mhzcmdDGAxbp0vcaw3rYj2qqPXaOh2aUcLAVtbkOEbbfIW9Z4F0
YaguPBEEtm/rxgz20hYn48ezdtFkKSQhbZihJtoJVai6Z5S8tEJ8ACzTsBNJuq+itraUweGSHful
F8cvSeyFz7eZNinTDQ6LY3kJllZuN4UbyZ0QZ3KjqgK40BW4+d+aHsPKZP9YSRUcS7wnfLt5KcPU
acDSwoLzdq2MICyj/iKzE3YHEfI5ib+qknrStUzxmCeqKEhAx+BbwdWTbtDKXV57as2IHp8uBf9t
0QgKzrx+TsiPZxBIBbrErnoXvwrFJXCdPZ1XSkUsVOAUcK9XGBNTglMfDNFjh5uGDpaNvb5wPDBE
wo+Ib1r93AYdSVJe69gBSK/DLEYuSZQJfmzlWCpBEcke1PLh63/rlaRe/Aook9imADXsJjcxApkU
F97hMo9ReqXzL6doOPcrTNj8oQ3CRxPs42xi6RWthM1Mjp9jOrAU/7QTGMx9+muI92mn5umCaLGY
pcxoMFbDOyWFAqnZXJzNqa4tkH14H3RpUxtilnWSeJ1ALJK+HJpCxZkZK714yiy7dwYBK59l7VF7
UnujkkRf3tmkyLyYqY0xVHdjyu/nyjpOLU8trTI4EcIPz51qacYE7V2Jg6FyDrxHKrgTDxvVrV4f
ABYtwbDNctZ1GqmT54JVwsiEOA+ZLcWmL6AFFASv+EGWdh/KkvzpCRbrwLqXOyvx8zRWoHgJD0Kw
TGHd4+D+uq9MuJxVE48KPczf/cymhSZsHWYgQh5rYGDE1ZN6Ssb/ye5mgCzusHkb/mm6QljeZQ9O
Ya16+gz5Y8qZDNACh/DF+Ab9tctLoQN2f79rVqJ4xbNYki5rx2bfsT7aeCz9iEYoy8YxzuG+5lay
9KWZnbink/e+3Se0A5AVKsgvxFr4MapAJMNJ9jWx9aeCI0FbS2t5BibIkst2CPsdYB3VC4Qy3tz1
mPS+izCR0Scg6PQ2Wa/+cGLIHWO6lAEiNvrqmlDSBr2YBtaS569pGfM6SmA1wR+wBdF4rPiBx6NE
sucp9SCSqA0mcG1E5+6ooYdoIbBIzREcN+Pos7UqisP3b2IcmBqiDDTQelmimzwvgj/G/3kJ4ei9
ea08oPaYesuW+aPzdCU8RV/2xwjV3ZllUEhxe1tC5c1WJFrVlk3OGOBvoadElph5Ly6sDs9qd8Ob
cUgqnSkMEeoRa5+ehIJNe8y9qksA8v4I3aGUqgfcroBRVLuyppnTzahe/3p8fP6GhZr7vGdFn8W6
jB922CC+ZuldIRffJLXObYuSqxXDZWarBIKRBapS0j80UxsJPmAejEMyE225HShKxXGXOcL1xV0I
56mMTDJzr2COl2g0UHS43R3HAuQBq9tk62Mv3kynUiUbHxSWSVkD/xlkxADIoAPYGWUri1IB/8oT
FjlxV3aMUg2ZJJOFSoH6XetNO2tf3WLs8z4yhiVSjhbqsThKUHN7zoM6OuHYTKCiTBXCxBp3z61R
ifULK/QQdR9FwJ3do7raASTZndeudhEwzGnyGihAVEMDWNziUa6Xfj0LMuqDLTps6o4aF0oDM7lJ
49ZR3K5rDjzmSJ+BjVFYF3CZP65QxtXCBlQZ0PHNPGwkctMNdf7NK0nUFIuT2g9vICj/+jZboNC/
rGkzHz3/wCMlluZVQhsC0dh8jgCNzk7hZO96kVUvQKtdFqvrBuN6F8aWaFsUlTyBAutDOwCz2v46
Q/6lF0YviY687u0THUA28FYYjBNnp6w5LyAme3ckKt5r2B7E6DCi1Lei87GYf4722sq+RsMMEPcv
nbez0FGTVyuV4AimYJmTuELXbhrGyyoy0/6NQ4iWZXHlTkl6g9if2QDb00BBO0JbzVXtveHr3LSv
FhDEotZqMIs4756dVoF0ZrJ0DclSLTDa/PWG728jhX8KWCeMGHoeFeNu3UFkXNGT9RzyJoq70GzZ
/6Uy4OY61RYYrrFqfikAmQL5hlVgAVgmMiKzoyslEDfUo6r8QXl6q6aE6JjRNpLVqeoANi2/vj+K
8sMEoTJrY7zKsjrNIhWVMz8T7heLAHGFlCTjReGrC8P7LuyknrUd5kkzLFWJ6lo0LOd2OBA0fl1W
wnhiL+CVE0PJ4KWXcze2ETX+PmY8Vp5H6+RYfx5VJz5HXdFkTpUQ+S1HiAuAYlr9tWlm8UgPYm+O
7Io2l3AeA8QXfF7x0IwN9mp/ZZjZkQvDkMnDE51xL4EMMXe2LaCTl+dzEdHZw4ryhzuZVU/0RBGW
MIIUDwrwzU2q6LXzsh/KBjjWIEgZrvegV9gluUU30h9UQnARP+qZTJQZSxTN2RbHpMKPMF0s0gH/
yrH2SCqw7R8S741oYeZkiiQHcNCj1vcDbPCebym68czb5lY0xOX6oaBrPzh3X7a1H4D40K+aByu8
30gl7oqIq/k3VGaBtX8f3CUg7qBOclBddIECIhC7b5/vGCkaBhpmUsrxm3jMfsTsKPnTtp6h07/P
uKmcb0X3yuokVuZ3Z0OLxaZ+7+zDsnUB9mehjFufvAE4aLDwqJeNhKtnxCJrRULsdIm4jSueXPEc
k2ixLYikd4O2apI7pALnp51xo8pwj7al7sC2LCUN+cJnYiHLSoQH1r+7rOoKqgbQgip8X0bXe8Ch
cBovaHpCPebzQtS2ZovTA30SXor2NJZ0mqEuwPwWsT1oZk7muIlR4Ezt46VTmWlnfry7ki48Mg8D
GsRdLrrFXI1n9MDWjqVuv95IddzJ9NMJ51IZm2xM0APDP9KfBAC6ia/W9HwFOHx0/OcOARLY3zJJ
44KhK8eqU35O5+ztF2XChYSnKUxjfaNNy1ap8RJRg6IJ2KGML612/8j5XdFK6x4DlgK024JnKm8x
4eWl8vHpxXmOcbwAcWyCjxfIICeESZ6pr+aJgSLdd1XnJlXvJE52JqHNNSUtEClixgTCF2/uO42B
6zXMHjv48ShW/HomYWu6Um4xphEdnd8U0kIQc6KmyQj1Hf2xVxzHNFxGMpqQQ/LoNgioLgi8j/Kk
k6yaXDE4kA3Ag5yJZacw84hMK2TXmWML6DQZ//HZqIb1zPbgIqgzS+VzFVCztNW5vrqDQRL+D5jT
GNWtk1on++tT+qNuEAVaCn6Ll/xxNKJwzx2XSEcaJ/iiPw7jTpAdXb6VdH7E5FVJ4p+tOEUyj51S
aezg0zRWInJ1e1SNVpubpptbOnjqBeQdfpl6m2rhdFGTuNofh3lX49MbGdjnh1oiH7aeuTFhs3p6
Pdd/sOr88pIFcLXLGhdCc25XE/5k0VCRW3V6nFFYYloNnsWfDX+mDsx65meUWJZMeT6hgyWSRF1v
QC8JpF0wewNric+2Y+1jPwSyYLdlZ6SNnigN3u2SMFuzQHN0d1LUvOSuwdgom5k3KHhoSmnSlkAZ
u8YWiKOg6lnQxi4lqmWVaMER1TV1GQhs4kG7Joudg6JLSc3qHs6tnqF79BQnkhULNz2VPL4EHScU
VUSIazxXH7a8yquEsE/tu0z0w+fcjg77vBpMhnxtfDS4yNXx4gKBFAkw4FVB52gwo16oox8e0Mqa
dq9mHzYG1+8cnLJcdGikZUNY2NxutwdmgyD2kBtUTIMbUcUg+cLTnlS8ntwcR/hNEUB54qlBAFiV
gOS2LXtpwYGhKWDerWoTpyXuYsx4SKDJNe79QyrEa68g6VGK4jS7Qyi5K7uU7CPa7irqbIKPllbZ
nvo1QppXcRQg7jRzlZwKlzdpy5BtPF0bERPvFxCWSHOe9ipOWXr53xW+86iRLiIXMtgr3AoEnFiR
vbEFpdlvcLHYFueTKxhBtNTB5rZ9U+ey8r1Woz8NvUnlOJDIuNE91BUq2I5Rj1xnx2Oze35Tk/r9
XgOxFmXbTeFemIv8YpCG0Y9/fa/oxA5hNzlGIwOCOnOYLEsbwtTg3Uo0Ma1GVSGRymgn2QC0NT/g
VbvMjNdw3ubU00FzMuCo+SkRRnUEKYNx6H9RdDI+vajSxjTXqGJBlRY7v7qQoKPRKpTTWdbpv77Q
sb7ZqYWPwflCN0uPXTa5ujPuvDdnp/Rtbo7BAx+J7nasePNSpVwLtOi1Pm1omLI2uVlTPrlZz9j5
D5M+qxOgUFxSaZAFUfyXEwU667gYWcqFJnZaWi6UxnpGSuSc7fMrk8n3XcdDsm30LOwZ17Tu6YGD
SCUnYeaOz5c7q769R5x7JJHeeD1qaYRa7X5m7qqgoO8ECBiQbEirOBHe45LoHGJZBIMEvZCmdeRo
bBYY0S8Zw36JAiHDxbKxAiRnO8nUx6HsJvrqQ0Q6Jqhe8xqj66nd90kMX2fN4L+kP9XD7X6Tp9Ij
BaM065Tnuy0iKUoZ/HMXI6P4k7uE8Vey2G9YHtd4WQdgMI4eKbLhWV2zUaNvXorCqPOvk4ea80pV
xADTTkOrIEHUdHvJlKjFDd+axuNoOMSHchL856SEIxv/v7xrh0UgdeIgHyrtLkQpI4hPwmzYJBAn
PHpYe46ck5dc5qBH0SqRCBp6SNAk//M5VuiKDhgP+o7rXyvn3KHTeWfQzpd4ExA+MPMJmS+SLlQT
rZgK3acNwNxTHTRWRHTiVrOY3uq8FPVLbgu69NS5TtYsQCG2ru6lmJa5QRUvL0ZUdhoY0podVCpJ
DA91icpUOtGUim6L96ckLhaK4ZAu35FRQZU++jCHuzJM+NIQPLu/QO/y6bQwAEAhntYOqHbbw7db
vDPkq+9oQKEBJILKQb7iPQlqxmUbOsZH6IcmB21SCbgNYDgoXPPdkxgCIMSovg4CkP8GEhVlKvo1
2I670R0j5O66h6tOwvZu8+BrMAPiWvu7XywKxPIvLGvhTZi7nllz6Y+5hdER3SmwKwQJPw697pCl
Z8Hn6YPtscdlqcEHLq2AzJmILjPirYHzgevcpgOSi8IurrwgBjelxDZ6NITFyxCiTnHZMFpTC/58
no/VlArxornbWaIHD4xJ5P0k6IBDdtLvbOhFcxcyQLoGyHzMym3qijxCJURuevdNuFydjG7EEOdn
Xz+cS85llfUuY1MXITdM/P7rq2Cl+R6o1KvhZcDQqrzF2RbIwUS/AFx8Sj+YtFaPJQy02Sb6Amwk
QpYuBs7S/kUrsU1aQJoS+xIceWtxrdyGQ2Y57hMG7kRGJT3FFECPgR+0N36MOYCbpRYDpQblYAy6
unapxA2CHBBr+cYLnplMoZFyrj30kMxf9MCHzhBrrGxeFK3K/lvjXART3Ci/dNGedE4QK7XNS1k4
8s97Js0kn7IcfwCMDGOG+9XHZkWnAJj4AKI+u4CcKwoQs2SNy5pmwLQ7Sb4yATFlOUTOcrVRrDTu
+oWZqYV/ysfurWSoWOq69W/b/YPbbGvZAbIF3AC/tODGf3lvxdMFTGstDZFJV8n26B1S96mFkl+Y
Dk218YWLpBakKnObipSLSYLQAs6b/44yw6awszjUDN/3iKtZtM65xa5e59Wh5hvwj7pznDuPU5jo
uCuYAOWxQQlG+bMYEXlIK+TUTe17hB8ZKDtSvN8QM6uK836+8psv0oVS1Z6/bFDeQSYP7I/Dbxlw
avyfURHO8Kzr4qi2U0sp9oHTmAr2uQAjwzkRAS+eJYqChUoLeq9TO/Y5Maxpmb3LEayDX3DGGtnO
JeiH0FpePfLOo1IH+nt+k1BCVfrIi7ABc2Yig7lgn/LRDXBODu2yLsJWtGcAuBtuxHl+iryGl8Si
cdx5rUz2oYS8hII1e+tHjCOZ3SoEUkAoiPll4aPB3ytpnyg54+8KD5BG6JC8rmOFpYTjvvGoUh6G
IJ1Gk1zoOBmZdp6L5w6nO1QikJ13JxL/O2VpnGncRblsgBKjzDMEGxJl9kAOetFCHwURbtkR6wYU
tKYwYqaNJ+amHy6NdLJ2iLX5eS60CUJK8vVA1lXc2HJEBVMg3bCjyGjGMZnVZCw3ww3XkBXRp83b
kN/JHW36kFXGGq0+67csqmZX5BCwyktAi7MtRpkVrukNi0J7K0mNQam0aIU/f4ZyxLcbhsTodnkD
d60zswbHRYbkcv5pioByNqho2H4QbKRteCz2Oa6DOiJW+lnQNojF+1z79e7Rmbi/oRfGmcM9HI5I
+uCdFleREUuLgupm2G32Ux/JJ1LsAgXSfRbpU81vZk6mfA+Sp24/jFPN3yRFZIEF5r6IBi5c5D0G
aX59oHTyA9ivVoOQ5IdjbdnlTMZaGw+7cfPYr5Fg+xb2Zro4brnFZXuo7wsGH8RaFv8BXfjbMXGi
/n+YirEkKAe/ki3NEwZmBPSiFf+Fle+G8ykhHycZm9cb5qVSsOwuMyGR+YFm5YnFYQl3cbRDlQ3g
NmMF0K8cyCuVY88s+etNJOFJb9/ExvHExRF/r8ZPxfNEr6Yulnehp52gif6k4ytBe8BuwCKj7eZI
zzuB+/3/eghBzVL/dQ5OvDnZ3URhHkwY0HaTqMuCA8qoCJ8WwTKwqM5eWh6vC8xzTPHT5bk/BG9K
XwVDz4QPe2x41x3hlSMh27hgpRaSIXCpW5XvnxfX4P0c9a/lRUj7OLbfOOLBVvyINXhhQZluS6bF
Td60HTlTl1kdUkPYyYucj/+/d0K7GHcYQtSyveJcxu3jPOblYhKMyAj3BHDrp+JSbUpGupfypVtO
iXRQVYKDU/lB/nseZ9Ur4CkUiZ+gdbFH5RkwlSXFWqZUmDpBTcx15bO5zg6ytnVHpfCL8/UWBGOX
F+DJQ0UbEGDeY1f1sSAvH7DIrMRqMjzI4bkJ0McjN9PG1pXOY/cGzA4J8P1SWHIVYzpUQQxR1Az6
cIRC3XISxJBQn4sF7FIN3wuLsii519vPVI0FTfniY5xKC4s6Qi/XKfw9lCyg3KErecOVMvDUbqra
pUZjn8G9zHMNCseTOT7RVtb21FVeNqtjZV40TZ5+ulPtxIQFu/tmPeA9o/FvvGqLMIBY0izpBn7Q
y/U+xIMqXK4LtDchJIEcRUCHoRgE0ZXxNyBCSs9p4J7cdt0DrqaUvXEQTZIKaywVl0PuW+fqpj4R
gg1wFE30DPC+J29Hv8D+x+gnMbz26jIkwD/X2mBfvT+zAM7yO1DiQIO/VpKhxr1l3p+FEpES5xlO
Y0EYOUMKMNLucNYiFsIM8+2PESIVRneCwCo47n0mk+1Oam45fY/Qu4wB8zopQDFP2QaZ9gnVR2fi
0FRKcSVA9dgJPeR6qw6F28h+1FPnYB1mebR5p7dvxgraxoUf+QedfKdmSdg/OYfsjGR0a54n8U0M
N57FqeT0ckiNsMcJgtNroZS8BqLXtRL2HUzYZV2OAo+W26TU6ARbbmNaek4B4I4m5Fpcr/z7SkwT
T0me3rMDKwJiT4oi/JaR/QfREYh3OJQUqTXnYBclhbwVq+OPu4JGAMWTWlsgZu6uLc17YeIPEEGF
ZxbY7Q5UBIHN3ob/QyWrlDGVf8Ojd1LyBUSeVkFzMHj7JJn5bm87osF9zGGU1MC24BO8SJIvvMUP
N/binLLNKEsBHuaOfCW5pgNqoZiQcGgCBQeqXx8L719tDMQ7hIRYmCeDkdXMUrJGqMmtw88C6/dg
p/71i0aBxaGqQXG+Gh7etlTW+mwP4yPNgjiEzvSzxB83BWbmmt+WVbbtWskod0YxfmiNLW3phNuo
APYSILAWkPxqt/F19k5pZu1CQsEwC2FH4mIjRqJ2Rm51iOMf2qTUQ6AwlsHkQTehBQNwbLLOQiff
kYvM45j4MXRu8aOVlTgDRE6DMU6x5+YDpCgeeubI+DT8t6LhiY6xsQ2IQJoDfJJD3qZkgaVge9xp
wgxnoArYo/kQIXwTRVTjIXCyVqE9vetq8UeZLnDto3zE+S7Z3PBANATZeKZKDu7+/aA1bpTIdIi4
fE2Iqa1UNmhLQOGfiRuuvEv9VD4r053farpia857J4YcFmH7exnrYB+xPhRLddBo/9vI8tedgsm0
Z3SE1HDYl6DW3Xmp6E76YN0Il8GCW8xotQ0x1unV/PsbFxgF38+Dc6Z73Jk+htb/RjG6xj9xvkFF
Y1T7tHlnwyQ1+eO8zS2qJOOnCdUZvyy2JdNFFcONf76D4vsIbVwxpuFKvo8Rs4Zu2B0/Iv2DD9x/
C0FcEP2our6jbr7f09929PpENCzZkERLc+cyjb8Ozmm/di9Iw71q8iRtZhFhsCNiDhBck2eGuGod
LgdwlDOHqA/qZjfWaVYqSlOowzl0TDvV9d3QFVKzbV4dy/5wy3nrLO1ct82bzUgLuk9E4OoZwhu4
qdENGB3Os8z7Otd/IKy9PzIPV7p9Y+2XEoFQyW8MOTFrZ3COHtK2jo56v8Os7e5gXzQwxnaoQE45
Kovg8X2Qc1NQC7NtM4gYTo+VG0TpCvZvlrjMdp4Uy3xMvST7U7WEpNdxiV1TB4qKfjKhUBLYTFXD
y6099Ez3unn57RzvalnpVLmbaAN49jTVOppiFj/iaAvdcH3IApoaQU+afZzKLTdkRLJsfU1cmHxZ
yhak6Dv5eyPzDdXqiA379N9EjXn4Tcf/QoBlgGBNfXUptN48n5DcexYXyrAZTLsCDwy7eQh6onWV
s2sVRZcAg19F2WxUFrBY8EqaXaOaC0jJPNXiCMsO5EfvswHiLdvlQFBBHY14+WBiawGUYWH8VL+3
CUcjxnPQ99yXN/0wqHcY2lMCm6PUdGCNrb++YiAI7dFbo4MVabozGqRnRoCu7w4+Y3ZX1qffzaWl
C5UV3/L6Txl5LAMG8XTXKfBTZHQYJSYHh2wYSYlFHRRf8RD5rI+RyK08/gVK+ZCd7zykumeiPybo
Za98SSoDpMnrTJzgdqjWWOeDgjqIhLDtE8/xIDL8bZFhYmIntVJcE7thaK+SMVO+EYHzYULFUYS8
fMng4pwsEDxU5KhQDToiXIcd9qmWkZ5igkfe32feDduCnp+Ej6vLkgsD8IY2FxNx9opfDGDs0x9X
AHLMM7rWxwTbtXV/VEMyEHDCVn412+T7dNVQIiMh+EYQOv2EbL+hFQZ2fDzjeU9mOqrVd12zRz7t
2pHpfjoLtteqxbskoUJEhFocHLj523QeabjWFCXgXVSA4ZV6IoPAh/U+l2JC3PGHwjCERwEJb7Y/
lx6FVRhA8FdPQ31wE82NXhAw8HumK6sbE3Gp+nL4q1G5RpBsBPAi+XvJ6lSVEDSUBi+CK1RU/Cza
r3fyYJrlQqEgxUhmLtL+MBknCCGRljeFNTXHwIJJtEWNQ+UDS0WEB501Um7LGkkKDrKVSUp+4Ooe
8dNFtz8k/tTIsEY0ftergBurTqkqsGJ1SXZ9aynUjxM9OatMi3KvXLANC2HeBimqmNXTE8/8cW2P
sr99DLCxN20chdZNPQlGXJGFHCI63b8way3D1qehVwOr2k4OM1/fg6JAdH+OljVyiBJLnQbVXku1
tLkzvLIG7fjV3mlBpu6Kg/lFFomFQjjBWCLjac8nRwa1xad/ydD12NOfdHaXXMlsi3MNGXMmmieb
SvRE9EOQqoeXKyBwV9Nq9rTRUDICJHqs9nHhCecXmo7n+KQOsRDZj9//Wurb1oIEGIlr0ZVSI4dT
eoZ6wwX2ezUe21hTb7KFq3wOMpb3K4Uu4LTrPjsFYkyErwYquS/7omChkDVl+e7sEKkaeNzzFPGm
dERFGoRy/NrPm6ziVcXcIADsinQB+ICBAVkTvE48irsOIOE2Lp3zUOG5VVtIBZayiUZDmvlROwfF
d/zdhx+U0Fr8nh5Jz4e4PaJAvMdL4H6neDk/76gWKGShYAsgMb09Cf+nHs/D7R2xPLWO4AC1PFtN
UezOSwT/GWxJuIQpNRRq94BtXicV4QDL8/jmqZ4M5GBlb0HAQ4QKjMH3BICC/nlyLKDJoPIXm7m1
BYWDI5UySngnlhI8+c87Xq7dErB2GemziLB1XfVkpXcR5+UqfeuCVzJ569FjbCLnwmzMXJrFqK03
dJa3l1nISmEWyHaRvZXTlpsM/sTF7WJXFBFlmCJjjcR+2vyH8JaHMLnm+Uml/E2L8PuZPjfwuW3l
gx8DxlGTRtV9JIpcuvd+WpM0Dw6qLmTc0sV7V47gFnuiGy2B1Y8gHZXRb/AtzMQ5MFoQBDY7oo/I
fRKcpOt5/M/pMR3IpyIlmXwfrPKevIItgcZogjgfCBThrEUE66WDEg2mjkR5yy7bRUHuRiRzydu/
Z3vykHRz1RceIgVHWCFH0M4Gvy+AdJ+Zy4wkFGNsza+giKC1SUl5KiB8Rcvhq1TZ8erwek6u/ogg
8hTavA98Db6Nh3BzQfJ7cwAmLznmj+8jb8S0Lq028CDV8Mv/2LMIppnGLbW8QXO1/945DnQsRmKe
1wfPGZtarunuZKjQpkfXErZeXSxfR5GQySBbj28E8vVtWrnvHY6hLX76sC3R1/GGFvn5Kat9c3wx
OYRIw8VitpxQdVHoFN0vSvEx96qaWjLH2eNRmeYYi6HjFF8UFOFyWbbEwLNLpYg9A+PjeZihwrco
kGifVkigPzgTN+N+3xdWaXVGpuseTvmVtp2YUveU2xW9wRtTF9RA6y/abwuTlX7iGPWAtD8Pz02h
xGWM33FF/wAgvtVnIyH/14FQCREsXgC0/ejVb50rnfUo4Oofy5KFGOKJGvGPJzo77tFXcfUTrhMq
LhEum5R7rIJMr7kLuVugJqpigyK4D4VOCF/j6PGcMQiqTN7L6zrxGR4a+DkRQPqFNjb/TgIojHvn
iv17LPeFtSpIUEgqfrYYbDX45bm6V4g9qbRmHpqAbvX74sYRWo2w6I2PF+lU4rzqCMHWcuXQT5sa
XAFq4qHPk8BOY9vadrbd3/9Q4jyZnRJ9Nb0gvPQ5kpa+7ukbURH9zgITSfLoSCHoyTzz6/rHDP3E
eLEDhVrqM+5x//pKL0bnGvNCzSN5PyZugTVoEqxq7bEMVz0qyQ0fpx1Ua+ctI4Rpil1X6gOeeJwf
A1guHwzFR+D3of4dvXnRBqS+JLYhTt5ZIBP0twcts5/kUv3g5mdx03SO13spTvFFfoYMFZM75f/v
NteVUcoEQSoUl8ivy2qL/6NM6ug3w5GTKQxcslU+8F2CiOVRpS0iMAhEk9Gu87Z4JBh3Zs8elGLo
puP/FAZB6SAH0EadNhNJUQhu7xvkMa7uXnU8HhMYU2YZbie8l+yLKI4oSZvqqvHUGSw90ZK8M1zJ
AJwbM33MO67d0tOBNMUymAuGLCehV097yBO44ShGTAV7MsTBpJvpIYxKjIWzbWY+Y+VWxPm2plL/
s3FeIyQ6i7pWfyfkwNZz27AZDV7zTLSMRaKPCSFdTS5Wc5Np0CmMKDOnpq85Bf2PfKQuoQreYXeB
k/I5LxvaPdGVu42Bk6t6nnH/0rUx+oJrrptKxOnhkm22LYRjDtRDKwJMKrpesi14z13EMCiysDwS
GWhu6Y93mUpnVcvofX8o3pIwzK89rUX8LtJHyzyusFwSTGWa6WxMOLT9YBiYNloMCHH35ueqJagH
b5i/aSnykf4WgKe3TR1CFTHiF0lm0REcM1mmEPnb6imj82AV95UPxe3fbagxOiwaGbX7SYXR5FmZ
R2qRkEtGaIASK0sQpqNQDMqb3prLWmY1MP/7ShN1+F6MnUi1cgRFEjtpUZAyassey/0u1qtb9whj
d5o9tpZWgblpipLo+y/yb5uWvHwy02Zu7fNt1pP6395Mp334mg8uLmBlOgw2NND3wi9qVdZOkU4i
hIavLasZQnX1yY8UHReOIHpPIthYHq/WM5cm6VXLpxrYpg/yQyT0UObEoNMjeTv52tmMDxqqi1+w
0L06+UQzInW4dzUMg6tqXIiSn/1wFWy5ySB6DBVVJyHHGGxqqAYQiHVo4QMsK0q35B+Dhlp1Rsnh
vng0AcSC87Koj+4ANbKaoz3zHQArM87vWhxbxGMaqh5y2Mit5IvxjyeVyk9SgEOKEdLMUVZ355t1
vWbKpmiNP7iBMTd1azfXMAeT+sscFOmVhhrHWGREWUn1zeURSz/SXcwAogwzsS0Zi5uVDb7bLHMw
Tw4+vigNHERyOjIzrKUXXGHOuMVxGfpY2W3WSRHSwRL5+ol6mj0WuoVmt2bhcyQY77MNfaxIhh59
BPWIiY4j/M758zaZtgwkIT876J/AIKW0Y3YGu3KWMXuPn6nYaPf+IXjrW+4G2rKyZjoJ3YERgIqn
0+JymSpbMdGxfk+om2pDauh0NxDpfJBKLeKIa5khgI6vPqV9egYr5sM8H0Fv4XgtY7TE5q+qE+Qc
xKEx0GKrSRevtXZbBSdPxV9O5TFKinOExy587b0dmEK+K7zgYUL2ftJpss8Znhm6+dNgHysdJQWG
BYO8tJG/7RFFhuIHnVmnalFnDhfW2B99xY7E9CxXjUY9YExXKf8e7Z2PQX8RjfL4l2NRxaK5x3lr
yw3pyclU0KqQ4cJh/CykLbO0S1TEMNM7xDcPHFN88WQyrqTAyIsJKPxNAmjlH3dmf9sIN+edEuJJ
ZICSS/loyuiIFTgzcLx4CvkiB80sAKBCSCZCpClgGtxpeB2rQmEpxP5K0nowVeX6qavUTR5Yaajf
WXacfZeTrXSBw9LV5Bsx6BSMnARpikV6nimBFd70w9ceGWC8XgsDp98yBbFbmXVJuSggHArYcBpS
7BRudxYuDDMwWs56+vKQfYvNXkZKFiO60nxYc4Gw0JCzDiG+RN/Dsyid7PNuZW8bcELALiCf/4xm
kDOnUBWdHsuHe2jj0KzI8JzFYXcN/t5N5ECp+f0KNOArXcxl7N49lyPjna6WiCMRWaqvI/qexhBO
sfYgw2COZba8oqKkAW9UZwdBsSFqVwNThFP/P7LTF1LFH4OxNTrY3tsHb+uOPqmZYYtGiVO+HV6s
SP+iveo4SwHZGkKqjD7OCrfMze/fJM2uVTEawApkTh5AQi3v4M0K/ETkkPgDdc55YYZIR7xp9ZqX
kd5W/1Nmv7UMXiuBJNAMBGZYqoCvb+h9olSxwY6qiAmwdpLZba2p2mPU+IumdodQ7ILX26qBTuqo
b/o4broFGnzPCcHLgWB0se5iUJ4nG5oTVdPSnGBb+Hjfocrx5m2xR7PmvPyno7XbYfpCbLuSrPyL
vNGSSUunkqak0YI07mz4jI9OKC9bvt2gPPBl4MhQA3pnOsj6V+tpSKGOg2EHC+sQ0g1Pbm+8t99K
8g4TnuyLS/WzAtyHVcxdzGjkXxGKx+k9FUbsUeODil7yilluA3+1vt6zIVTwR2KGniQtXbkwD6Nm
8Bsn8tr05cvTvGPZuReE5KcbxHwnFSf3qs34OkRuf2PN95KRhwM3CvHktXLyFpuqpRzgA9BBDmr9
sSrPV9Pz/ZyhtBU3l5Q5Cadkxz/T9e9f9wCgxj2v8ByKkGwBkCnrBmsrz1+Dcks4vsaHASCaMVno
ODwFJQAocOL8ttdYE7gjfHWgh1bYSzY+8P5I3Hqe8ldaUYrPZfsyQHK1v5p+RVBuCgoQYZU3gV5W
5IB8zyk06h6ZagRlVvNMvMv7Iohelg7PZkXJ4gzlgIBBwfhjujMz+bkyW9PTBcN+B+ANMI+9kh4C
oRAfSveFLY7hrn1WcYtETlCjwPbJzArJLoS14P2eu4XdF4WfBIqncZRGv518BLIGEkBm/uFynY9h
4Teks29511J1CRJn80q5hgSykjNRdMRFohp+z1wcQQpdOk2k6rvLq8BvQtUnr9dmAkZWJ1HoCBfj
Aa/rEVGbRKgnEN8uSNgFGDDHe2feqc19bDJVcfkaykntBMjH2vvAZPR6y9QOiaWwmij3AygoO4id
a2+VAnrGbYr0Uoh6ZWrQ0ESOQ91X1DyT8ng9zb2E3ld/S4i6E9likOflvr5WzKCFDIhZpohLhXEc
tE/NpdvZpRfMOI/rDQjx+KwICUt0utSbZVPWv5acrO1lT8e1F7SG1sBO8wKXrlFfFx5vIeeMOVFv
0VxL/2K72fVtuWmB4+KLZ9l5rNxOmlfYXx/hURNrcwDhEJ5eXWZxMe5XYOfddoaa5QZOvzRlhRoX
qRFfXQwISMcVo6ioGQ6CpzogVIepANnw3vFUxSP+Uyfrue4usEQ9YAqreVokjGJCmGunHvXNf3qY
kbaaPgzms2uLpxQ3sD9NVe23Pusz3op9DIkAJWaro6DMjlLZsDyzc9HEeYMLCVjPWos4jCthds4k
ILnEc2tGaUoL2yS6qKkzX5NwEm1CSoecqityBBLLl5cuO7VDxs96KKsxdu2rYAa8pvsm4YkcbpPt
fI+sazh8zE9RAaQMRDmyvGp41xBNzMM1sOt1cIx+jxvBjRRprJwBeGxkXUEFUMPAng66yWrF+Y4W
IYmdaGWNJAKR4CkXJWOn7QJ1DLP7i6WC5DNfECEGDkdV2mn5cwOcu2tENlpnDwwc1A9//Mj6viiI
GLVyGRH2hkmoL/8Miix/OK+ZLGRiU/QI7Irj15Akzmcak2dQyAcSxPaFfFx4rRgjmK4GwijdLYTu
Psw4bMYw394ehfEen7wyBCj1+qfEd/jtwntW8DHuBLD9GJMVgUPh4cYCCwq73hpaM+juQVigEQSg
b8R+z0Ghu0lt3DwiqcIU2bvA05puugp68Kx+SbZQlzSPsmQcWAPrgEKgxgmDi3tXJzxpZoQ4uz6M
Fm1Lxu+Y7kyIERrAycSnqQ7BwYpX8gzw2euv0AdBhgfZhzI2gHJ4znUrIGxERErqxP6Ur84vG07n
hHg0REZYVhphdlcH6muQ8XNvwrx3W7WPQ9bMWQoAe7cndioWGA9kmfAaCmWaL2dagvyfSW2eYzhs
cjg5Yti8r+GdIg1XdP9BJlgjfsWx26Mi4y8tfN7DrouerIeD4CWBDAlVvhiUnhpFmgBg8fwAVYnv
Is8108P6si+QjoHHQcPFC/ajdjm2bDMOqHtTRcu36wYH3ImiUDmOYeGHH01fZ4jJdlWWFLIQRM+q
gmKQmZHtWEhe4iz1l5jgH74mTK4j+N9SPg/wSNKbThQ9vMDy4k+WUPbDCAjE/zi+ldF+3xM7rPv4
ivGIe9Xrbteqfww0uX4pb6lXv/0vR18jdIdIgQuDCb6gB4BrhMfHbXF4MuqOZnP5Jm22ZueYrkEg
/W0ul3wseZ0L45kfmt71CynZ9jmMiJ6kYzxKntAJAl48UrYIXxYLVHvPdgr95InQZN60wYv35H/5
6iotPxBOsMtXFfuur0kVwRXwo3gFMnPWnqFx+4cRY2MT9rGYcnLIW+R4FIz+WHjKGogHpLBtEL2z
tm779aMUhb08gBN4gKaYtHvYo3EsAM0LMAc/gzBBiS0HgCqevVqtmxVjHsINomOaRmxPZH93bDwL
Mj2dFyDFMXmFkXEugj6xGeeLpcpOgrlGkd/Z9wxWVKyYzN6eMc1rnatLA59xWfcgqNYYtpkEPw9l
7/g4QFkrIFNaulfShNfuNUWwgch4DO5RJn6o3EoLqrsvP22tt+iDJgf/TGJ0K4EsRSSsnf1Aayg0
PHBWEsOALaXe66WCMLJovrW4jL3s4c2f5yMldIf2gbmxaEnSBt8KtrJMFQ21bZ1HX64nQkN5YaSz
xvhL2Ocj54RbJbo47qWvmRmx5qPQGsLksdWizld8gvPRgJNAHl92vsOO9K7Knfzp7rdaABMeUdZG
HqLud4N43SW1QNUlDlqUh/UQ8/9UCiKFeLj63T/vhieZHrrvqx3o1ltVyyDobl6xskUXpajCCU3N
fEEw3yOpgcgeDTGDGuHIwAr2JgGIxIhxc2a7/ULAjBPF6tSpn5lnQGAcV5VO23H3cat2W2QMEAyh
HsaqggJSF5VWU7sY0yGxvF/mxaCVpzYnrX+bSkX30s9sNAyiQj08gxfba4HAIl3+esR8uPoy4nB2
/UgRoxunWJVtZ7DCLqTl6VsWwwkWp2N3OMIhZH+/akLhG5ut6XzAWGT/fYHgMLboFm01/3+nlukH
tMosiSc8kD/i3DOp/XL7jP+3a4XS7wb662CtnQMHTY3y8Hq8QBx/CohBKDHzB7+1z1O+DKvBDuNb
Jw3GLwfBkaYGS30KQN7VDpTPjgjdyYs+J+lla/+qW/PwcPoR6LfXj5NxHh5mC597kL5V8GbkLM7W
+JnrORlVaZIGDmco59EH9vHOu7iiMaBCgSd3DuZ6Xc007yflDCU0TjZeR8nTzf0TWCeuh6ChIsyJ
OvERGdObU2duw+Ljr34ufVvVmFS4oVFS4j2HWwlDjFrjNUH2kqp3ytOy05SPyMUPqVz/kLoCZb9t
XdHO35tTPaB+t17kWJ7vh7vo7kckjBgA0Qk/m9cpJSTFqsOZ/mN+6RGszAbpIGTpmV6Rm8H6Bj82
BZTPA8QzEC3BKSkzjOJ9OqAM7aIS8dFl870UJpkMosrvq9tI7vLw3ckwxExm/R0VKuO2TFP2yQBj
Q1wAPZNqunbQpJPUyHuosN8bQLLdK2VTs+vxZQpx/wSQY1JFfaEBpiL1lRS5svjCWcxdPXwuOHG+
wkKQDY3/HNEz6NqUXRR3g+hnRcSPb/PtSMNiGarKcZ1ZWlANsSjpnBQoJG2NO0HIOXb0j0xh0f++
SSMJXTJ8lkwkof7hCLVyKi3H60C7vo43Nhw8eerF4jfNINpAZ2roL9Jih/BVUPcVsKE7BQfiUImm
pnVVcVsCHX7MMFRAsY3n2mnC3SgzatX8N2onXfhNQY5czr22GAMcnCNAvshS8UEXuuF2YN1ap+Rn
H8dNQ00VWqvddl+p1UHL7V0T0nzPR4XUYDQof9hBmKFgizETRc8hKyhM7gidbIZeRwRhrd20v/nZ
D0G1SDDpDsa+eWm9aLpTYKyDdl3ptDzJ+syZUHeTl+m3xruOodoPPoFY4pRYnUMM45xZuYOeVrIt
t12VEtC5ULQ+lp2R0Z+nOqmY13kWvd1yToIbU+Vg7fy8+psBBfKx5G2W2ecDPVZv1BGXJoy1bbz/
VFxplWoc+BlnW0goy5Zo9nDwbaJn2jY/kFoMUF35eO2oJaerlpdNVkYaCM+9S+1KiTn608tRYBBu
TBmleMAPfkFV0wQxucsIww50hS+hXNTP+khtkJXJjueV3PYkK3dcvapE2bsMBt+FgMSR+XBVNjrh
JR3oUAEoOmrZYXnSoSs9ccXO8BGIwRJEMMbOCJAgwPp+PTjawTaBReYfcLiuRukiXKoB5jTdmnXK
7T/xZ9/AogDQskx8/irom1Dmq4Xqa4DKU99pZJ5sdKOtxw41uWn+QZpPheAgMg0Y3lIsdoCidxc7
45Gd9qxMw6KwcHqD4BU9l0EyGcB9kMj5wGKjbVhfGs5F6rv/39VIGSAnxzATcCMsOk/xJJ5gtWvI
IPtdFlAjdnCt5XNO3jPv+MAC849u3/1ENm4Dgu7NFYOsK9H9ORT4Jk4H6kN4FJSjXZhDmxcEz+OG
ZVLkl1s5+q13/Xaj3ew7XO7V56L1o+cf8/lrtd6AF5KlDvHXjTDxjBZk65Z0bL8NnK+JktD2t/em
T8b3QLSWfYehJZd6LW+YSI/4TL9oDsgxsgP4QUuJ48Pm5AcZ/wb0eAODzLHUQX9G/x6wlO7dSg/k
mBDBs+dGljp3v+wm0XDPtu80ReMXlqbCSLnumLmjkuPWTsi0wof0vx0GVUVDkvhX7xT4d4XFznYM
k+Ir0SYAJwX/oLv0teZ1yUepX5hdMkfMlWMdpv3C99ia9vTbQPapGLBsVDdWsjCXzzjEWg/G3knA
+YtimhxdWirN/SOj4oc0g2YVSJTTTdpd834xayuyebUsV9H2FJEWi59wt/PdavuMnLCkxW//LvHU
LtSXGXNC2ihfzfA4AifZZzLsrG3xPRhCSTiLr7rIGfkiBWlFp3VidNpYfsKmUKLDEVHOi48SRhcQ
RQ43JO7wfmn+okkBf5R0siQwQpkBdg2FCmksPv92lOhmV6cT/U788L6AnH2PCIwl9Ygln7tV6S5T
83NMBekf+nNwv1JD5AiWC/pIrXgyHSAoia43Eijb/FdfzC7iexTjA+q98vdR5rFqgc0eJj+eiCTX
Y/PK6LH9acATyTd5rt1WhlyrQ5C0IbjeBXhCDN8ZDn1BHJuCv/E0tBYUcpqb34rKwoNevyOH98U4
D833xozs1E5wGQ6J3o3PYzwCLlJDpBbj14WXG7ZmaQbSX4HvHZO/1EVXRZDwHAodQ/+QjSVJq/Nj
kSIdEpJpb5vR8LuHjUlUYTCEc0s4vV5LCMsQi1PlEtFRQvqxQs1/94znQFiXToAZOwwTIPmjx1L8
QTTCjOJ/JeTlDIRbuN2saaCmtj9v3GmxvPntu9ksOUUzqtsSiRr3LuyJs0FP63J8nkN/hP6WZPK+
lIxPmJ7RVn0sdJtAoq99gTk1wkPIDNoBCpAHfPGqWs0OiE/UDfN1upgby4sOXvf9fQTtyjxpJdrh
4gBKkxFtQzwazwE8wRjlR9qNG8/AedsM472ogTiRtRivmO0epHCbTsmgx0ACIV01fmSrbKJi00SK
RlmTwtBZ1HD85oLRto45KfxQIQtM0uvexZ5BnCzPbK5jT1SXZCgZA4f974hVlHOTaiS5foSQka0s
IylOfSiKF67CWJbDBRYW1xxn0EtgNu0FObDfn1LmuuqNXqvuTS23KsOgE2VaT4lRNUxgJ6lVBAyV
Zhe8RpfYq7hNImsiMO+HWAbVSQeV5QGNRTgZeFZxg+W39sBAWS4MXp0kfptwZwTox0jNo6jZLyJ4
ryYCz+HDhioxsssJ+VXZYTcSumMdGczuVht2O16G9Cler7GqUgX0zado+U/1PNK3BPU5y81kvw6y
32d68TM+FTCGtpb3OpcyhBJBYInZh0JxZwjRLQAQ/v3VWZ/EmiMqg//2/yKBxmFO/xj0mJFdgAHn
6H2Y+cE2cO/nFIR4Hh0vTIdRM578myfEog8PW69aIdj7/ZKCIWmR0S8xtUcL6InTy5ImcUQaHYLb
ehoDhi9DmnoIekcN/gB7c7m0HBTcv/2X8F/vNSPt2yONSfgLMxg6mUP1YdzlRdV/A1KS5fHq5yRa
XXBgK0ZE8up8neq0Rz1EIoR+efQN4zpCEK6YIIq1vCTQWJ8c78KgTJwtgcFfQun+h0E80Qf9QmAc
3/i2T/YH12JbN3/uZYnq+mW1NtErikLHDhqVcPaEi4WTiSg/9V363jyHra7er9XNqwjqnzW6d/t8
GEkN2+9Qv2qqgyViYZMxzw18AhmadNgm3RIR5WppEmpABWk9QPd60bwofekbUTt0Hw5X4Ve3jnYi
aJqtXFxS1ilksKCNf6oR+IbIKucPztt9GXuRmI8mmoVA52exrgUxBS6DxizlU/0F+RhrQ89bZe74
bZaFfq8I83QpDnqsH0YSstihtcrLMfsRq3+vRgFwTQyKmA04je2bVf6VBr7Ne/qPQKXhKgkIU0Nt
3R9WFqMmRGLbhF1SOr0vM0QZsB6GVtnyou3KGrifzI3qQv27aUW20pzyjFDbHiJqJqYl7DbeCfiG
bvT/bskpMwbbC7NJvoSnX4x3KMmF268ahi7kGTRirtu7VDiKqMAJPDf73S7NE1q7FKa2CJB2AlrZ
ZwUuwuvA48dnFPSwS325ISHUMRaxPqkl5lBuCKJcoi+0Ch2wCCVncwJDsUdoJ4Kp3jV3H7ZLTFTQ
3TPXPIZu022stVC3CGUMEPL67Dv1toOziFKJNlX6OlXXtPqnaImYiw26CM34lPbYKHvHeJP/3MT2
fzWMpJZ5+a5mAC7jUBY3rl1t1YSncOYqZk8VSBf9ASq2ljPWWKDjmKt4FkBfa0k+Jv/cwumExKJ7
zVNId0JzJtO1dPQ5YGMl5QPRJks12ZoSuZmTVMcL6xlhozumA2KAEsQb2+bpwL8V7kDhhefaIpEb
BgdWR/urNfvlUJevmPmfrpml3LpAx7lDndNVrwLEfu9L5RS+ESAup4mO2n6gOCqwEqPLULzLr4Fj
PKcCW/gl6bq48w50HWu/jIktUyPRgP62v57OjH+wl+J6tfYJgmEw3i/gMqxRGef/y9xDJFxR932k
RrFxAPVjV9pnYxNs6Z9Hfj2zUNoQzikIdyLSJqsYyRqtepy1SK33cVmkKFvP8rTkiGbtQQV7XtXy
kEhhmqG153iRgP3BCCGcjomLV8Uxun1wmAc8Y65xwl0OjP2pOz4mFBmpD4ad4fqipCRk1Ba0bNgX
Y74jxuKfbrKr7rnhNgfDl8LuU9QU7xD0ae2vh42wKalS8yx0bTfx2HkUQeZaETgro2N2wCek13nF
p26TK1/IRF9ZNL0zIAT2UqCsixbhEY8U/iLP+sbV70MtAX4HPhHsi66oD+D/fknaWhHAXp3K5qg7
O9E7bogrT6dGQ3WUaaO3eNnjJaO/JdvVqeHyd6nEeHUENpUoatTt6W2mPrVB893Z6JMyXM8TpX4C
SGBSqrkWHhkL5HUafYfVi4mK6stagXEW8FijlvpCOqNNPC/ChHQKkR1komPpBkXeZu2QG9J52hbO
QRQS/eR6R2ePaDOoq1Rb/mTIAZfiptAer3I4PiE6kwNb38rwPlBiOHoOtW5992fahq9mNmrSPsv4
tSuhhv2T3XgCI28P+c6BiDszs924TIi2bGUHp0nHGtxBUE3SJAJX7tP6R2lAPRSBry/jmYNgtIqy
5AsxjAbQ0y2Qg8ymroQR5goKwv0uWq78P/LKUiQHTgpWfsySPQczxQcb0kwgmMaFwyqIREy4DjDW
p+hKbu3LG1/fdR2IJQRfnLq4wFEr4SAQZggor16wPCrxHsaFHK2imedXTrq1xv9G9rYcG46YkPlt
779M7CxZvs6WP22OdqI0StUS9yr4kEi31Zc8vdeozpMlqPUNijHFTpOzZT9s4WwAuAp/YOu8j7d8
3WEEM+u40zmS+xkrAKjNc2YNAVGUnwHZ2gdjl9qmdgPAicR23CTGVlOREle9mMtaPpuqkfo7GVjP
hIDW/cpvkUzYJ9gAxZctPVMs0KbA3RtKA8gFDBnOeuIuo/eZZA9GTwvXClSWyycTfSwABkyVRLxq
sTii9fBdqWq/yOHbFZ+/Ye/tviteXN4sfiyqfISEYLi6aN6jbSI8oH/tAkFZ0uauYu2Loupi657n
arn3kLoESXdcXjW7u2oSRcrCIpCMM6gzzS+EU9eLtPxi2gGElKPa5YQssmLamYLQsJUw/IF9dQB3
JNA7tAk+5Gjzme94HWwV6gJxiHpX0jmhSA9V6HMfk78Ny2SHed0kaRTBI02LhR0uL9otzIiOtRZ2
0FOEZvBs99tqh53LGoN5hDehjLxLFvn9Qd6b5Yy2oujJEpJQTZvBccKHVojDN+iB9yOB2Xl3PMMM
PvOq9G/y5TfQo/0PS37WdJwvb5ucF1JnXu8Bgpse1FTcH0HKcjg6sgpVllcMvpDCGB5XCLYixkKx
axz8lLWSK3GpXI1paAOArV9pkUIexTGTonWUJjIxj8F0ENLdxaYCioa48WNjxpZeTHj7swFEMmZw
Z6vnNs+yt7srQvVbYs/Cge/kD36d//zFQixMHl4bW9HJkBEwj0/qy+ttXDRxJCvjj0CJ/trYxpVa
iDrz3Y3FRRS0zbUgHiPYd6RkM6WmCYDjSKAqnjJw1wDAoTcBpSoX1cseFNP0Y98p+8KNDvmDCsn7
mWtMz9W1eA8mJSngcBKExB8/wwGLaz7MguI6ecz3z3dR47Q89vDmpOrhuc0eWWY0D17rPgkm4yBG
BeH4HUqUi2YFHbBvFFt+HLLTfx3KFmczAwMHsXuqZVNNxYA4klmt9lkJ2NZtnJayKoiwRaNpL+jp
3H1RXET4U7GVZwZzWYHgIG3nySCBW59RHK4JQs+h8RIG01TzAGkJj8GKLcWOdQSteryePcbKBHJ+
r0Fmsn7rObTiKrYTzzBW6k5DYyqAn7PG5yN46IZyOVlcvaTPUhUv17i/nFlvkg8sqGYfr/xAAy24
tzBn6kyZmX7SJ40zV2GZpE9Ua9CNWltmi4MaL1+ik01MX41h4R5W/LlKZM8ncBMqJSy1m7cbu7g2
H5sKs4h4TfLzed35Z3rH71Q6I/L6D3nKWtArSnKJc32fcN8nme/wRjT1AdDY0P/AWIwNA9EAvXgF
HZTuA/s/5s7PTBNeUJYyp/+c8bnb87vMPqam85IP9buQh5ePMx7299lD/MFLj6EPxIt5dcc24hL5
H1jnXXJacxf2FtYBj+7xaoH7hUZkf8LgT8EmECxPk24Pkpmv9yvzU5UCxu3WYBnOSqQbjioRIA+Y
q7pjzlggQ8nigTSXLcwaYBP4MWQnrJTCyfP7aD4G6PNAoGpdHE6V4AaqgNqj60aV4ibLq+6gMcAg
czyRJF1lO6YWT7xwUI1arvdI5liEM8TH16Lotrl4WT0J746yQ4B7cLBhYoVphtL6eC4KDYeOwmKt
ahb64BNRe7ZhmdJJXRuashpW2wGXkeTRtOce2IMgHAiTObNJeEkCwCpGipjJWi56mD4xJe6vxpam
+wpsUpPRyT5ASH/Tezkh5Og4L1UL0ke1zf5YikO38OJ4YHPQ8pQcjENygadAkLFi11ckMI3j1wZG
BTiOCMdcR+TmBYkNnikTqmj43PF0cXCcnRWXo0oo4mNqUGNqBc7pAh0WxUgdeZxWfX6kNeFQH6h/
pT3xFun4tdvp8PpJ+q6c2GFg0Fya7z3s++qz7viEHP1CwCdYw7XsRVEZF0Z7q2+KM5KortAR832w
q+WNa7Tty9NWZvN9aS2zzEahRkc7HwkeEjrb1ckwmxdz0ZmgIs0Hnd94jTzM1Bff5AsdBBYDrQ9F
XXa9Ef+SrS/g93mY0U8UttbYqPoN2dPaI/UbQ1JM+9IgYv3BoqM1I6z0IklmYXEW5NDHjInUDsxW
N+zWmU3Am7cKLeo5aX32osUm5Ytog2lLN9qjKkP0cUigbpPlU9bHfskYU5XKgPiW3YcP3dL5JVnR
bNB1Lhlb2+BGMnBcALjZEmlsM8kceouDGLw88MgpMCNjxixlSn9DBKT08mEbH7hlbhoHkdpk+OpY
QVuAaeL2lPKW5lfaOSpzkSo61kYmKpEtqJ9ZJjWTPwVitUy3iR8gyMp2asIGnqV7WDohPL0pnU7v
QZTi62bwFkJG+n2oZZs2lh7DjXL2rql7vyvjNqfQxQY/N9Q1WtWAvRIgJuknGdFC+AQQZu+kreGc
a3VT9Kg6hUo4zbxbJUZIT4tWv2Iw1it5G2BI+CbMjDqPvVa3leP02+10hGyxstuq4gxO31J4Zxxw
cWfAXS689DEpEohp1s8uVL+/f6emwX71BYrUOM/GK27w1UBWqc0hFe3bhCkR6Vy2FG7pVmWcetAG
AiYHyOGBo/sAuOIj/bxtvEQDptpKLTr2ZGFWTk9tw3lLvwfnBMyWp3xy3gEZv0J1PYBFfURhsbZC
7qfEuJWnFQQCmUQieTzQVZGWh0zCqUC5EZrudS7OpEhNQywL4KjcL7MktyP8/XMpkXQqbNA69pNq
biXxT4dAtynNMiTMosx4vTuSt3Si60hf1VzA23A/MTPPSlI7QUYjhECGVYxHSuWKzMUdlQj3O71j
FqTCtQI9ieS9ZPrgm+ulFBClK5zXN7/GCnDdZaRpE2TGcwzxRyPBHWpPB6JzG3/jj5R/aYttiypC
A14+gB8cEZ7G4STdLBYu+IwtZE64rMCwGUOWOh5vYfWDQ0cvT6GYy4mDXjYOSU6dTrkv/Et4pTst
83s3DPBR9MbEhXEGMm3GZoSCkkARsQRI+TxecLdP8J1OcTIAIh++pja3lClRXs1aCPYPAFxbIImV
w/aisEUhg8Oeklj7hUqy6zu0dpxKaD+KFbtFm8bR/mZQVTFJaBqfaPcEZsU+l4vWZxYCXZxsFPTu
aVOhbytv6caV2qZISTrJGtn2xEteaTIP5ZLA01LMTQ26sTGRzP6/g6nKUaLSgQQD4dkauuKDpufV
wcX/W8hcsTce2qah5PoocMzNwd/STBDOfE40xFs2TYIbTb0cpoXvng4JFRGkOsf3k+8BEXgaJPt1
FXfMdYXo0MZFzbj+Bga49oKSfXS4rthabzNKcT/GIga0PVFBtl0Yq8E5/VGJRJwihjk4D4aJ9Mls
wQQJ56TvjxNPIq+2ECVHqfXEPkGHkXGw4CrkWMQNTeNOuxdWZ8koU4m04z2vGzk71XnmbFlJGNKB
Tfpqla1ZHY5DYC7DVP8BU5whTcbrh4EhTEzphJ7QRN9ZWwvWfcx45J1kvavorjwIRKFFYttc9C6d
riI7yxdMDl6aMwKKmjAZ+iJsQEzZ0EiAJGSYao4+/kozBxrOG0Tes+JuQCeezeXNMROPxa+jULrQ
QHcg05/uZiyFdicegft2n61L4nwAO5WeesgGoGrTdhSG7r6xqWsdMdNXEybfTuDdOoU3b2VyGYrk
UIfJat3A77tEmHDotmV4FJnVBVpCgH1tW2GNvlxTYbtjJvWAmuvD3P/BbAKohrXUBzwMNqnc/oNK
/RPI+79C6zk/j3X6XoBR7ulP8s0uibuw4WKDESqehEE3vRsAZuXD1akCThu1kMX7cFyN+Th48U5f
f0cIEuzAO6jQ073XUZo4YoatLHu4TYOv9RM/FRPQterJDQCV1YTr1zDtevfxagG4HtyOYG3X6N8/
/wowBZzO21J2Pb8SWBsXFyjnWDrkBT6U76tYX2kvyfkCbfgs4PP6RDFWM0X4yoy6TD6K8w3/Zjgk
JfgvnK2xVo+mMk598FGOfJDkUE+oW4E9po0EBy5IO8Hx1zYjQRNSjWZA6px4FuMO4KBnikonjMdI
RBayXu2Ka7RJcgQpW+s18qlxXTA0Ls5HvGre5+nFq0WZlG7zUHaTC9TnUcgZDsUmZDMRPD8F5mA9
+CcZhH03/skBDGiEb0bUqOQ/ReTmGX1tbovnIuhXFkGV3/hyMphJCwnf6OzUMSaVy6B61xIAMjGJ
mGogQA2UCy+n1bFcgGyjIv96wbiN6RusL/r5WvJQeBaVAtfvXAQZ2FZB22WyZb2kgJ1CXk7lWBf/
RVe6WX4DF7tCQiqURElIb6qt9xuxlvqx3q/JeyS2xptljjlUh/32O14BIxTl2eQdiOyd5gGLcHtw
Ve7WZWxtPN4Lyecjexgwub/OZ1ntO5hdC7gGbopjyO0uOMpKCvS5cnI5dC8uEWFr4zBjXaRCzn3i
Xu0h01VuvkqOK632a5XDTw6GNkWctcb6O9Ll4PpewWMvgMFYmVH/c2+NoX3MRg5VI57LBvm1U7Sw
Nkt0VYGt27lfkoM8A8hKOpIDeIfiNx8WFnxf2+tcrE3Iach+oeFCYiX2TDd0kQL6/a1yzuxzL1ct
b2cd0CWr4JINsQzjRhU0JnVgMQ2nFqMMuX3bKJAdMbaxWBEHaCYxv/pHQWfkFzGn40fSFB6Yjyhl
7a59a6n7ZgJa7OansttBIcb6+0VVaA9bqeNDHCYULrVonrONz3N/NfBcfsf7eAa/ib3Y6Y3tlXU6
i0sbh8cNvjRAqM8IHRR/8Bq56d4OQj73unmQjptH0HoKRN2dcx9aaoiI2ugUdfwv2jeb/lIFN8s7
usQE7/n0YX1BOpBZkMP5Lt1fEQYlzOlUbhAnXnDEPr5oWfG+Y29iDLsb/wTioRHAD2r52sWvnDoc
V2MqNtbEDafebceKKemkxTKFgJm7nLOt9TQL9CiBP+I+wT7ILsvp3nwYuJpJOv11KRRPIXEhoYsA
9VpU+UfYoFm7PrARY+X6/xDBQmImowEgDGxNkXDaRZwY/BmnOlzlkFpWkhLDO+qCXRnpaQmZx4FK
YkwSK2ut4/ExUxnxb4dkAbInAqZwHdk7BKid2jqLmV1lgNfQ25fjmfeyb6ht6R4IUyTCFWe94nHj
1TEKIKGv9FOGJ2Q1lQpsXg2BpEgmi3sK300FyRKxD3Peek09cQ3sQt9u2bO+zKkeUxlphmk8Zt+X
/8wnLCOJTMtLtW+bgcgwzqhGtXAlK2fVkx67F7p2WqYWyx5G0AM3yO/5bsBTPUWR56x0I+wuzcOh
ARwUd8JVoy0EkmRdJBA7HA8ziIC5RJzkcW3LXETG74Lp5f06zEPiiHg5G0K6e4fH9+Vsar+yzJux
yZ3OxskuLnTyAMSY0cncVVHYbwXPGjWNoxMz/tGqpMPPAXMrEPXPpiz/B+O7s1q1Gzbwi+BOALRv
IsOGfpgM+0P/4Q/ZDD3zpRZUvPsBRJHLrCqGf/fORVKUWEREpB4mwnmXPntc0nPSZ4YpxJ4x6Gut
8xlfMkFbeoOvjiPc7reAEY6EMzblVdtgO5q6Zdg3q69WpgZJKARWQ7yrUSfxQnhuLdRpT/VPYLbc
Qtma0miuhzUtnv67Oc779uPR+FhMERPa1JBFecoRdHNBi1I48+2aPgiZ73eCFzUfGZSCN+7/GSVL
bjUxQu3vQ/bMQSjKw0f9jpKH5fUDEyGyaMg1QQpCoJcNCP204krJ2MEt16M2IwnGybuLsCduZQat
Bw2Y8eJ1ql7b3q+TtCd2yPmv8qDuJwTNjjcfGrwDL+sPd6OhSKcjaTjk9TTVPFCGFcEoTmNri30e
EUxR2E+155iUVZ8mdLZaeTicdLrtOCba4H4psX7n3pMKMymwhMOs+NhQ8XwQumjfe2hIDO6qoqSs
wYr2ZC4l/9jBRizHiMnWXQnmukt4gRYkJGug1g26WBjTGqJ7Qcv0dmtreggj8JP7NpD/EwRC08NH
4Uh2ZJYv3Hye8VTuCRisl3Rvjha+VtX6BdHFY+LmmtXrcgPvRjMeIvLx/tt9DTlQ08pz6lFC26hK
Qkk0kZryzDqV1UvS7btUd4YxG20r1zg/zxR0tD8+gQQZqzr0Se3oOx0gSZts9/8vfHi3YVXsWW9r
JZqPev/cx76zoLRP8oT70kONDL3kI20pdY8LpEts/Pu/LqQ+FCG+fcvp5JtMWudxriqgAhJ9Ai6p
ceEDkmRdK/PJfLYm4VYw7hFHE+HV1R4IM0aQIBD9bKxOBuISxsYdAjxbhx07hf5jOEl1CY0rIWDm
IN32c18UTRDi8HBKrXhxd4bCUL0Sgk70beM6vNcmUvh5WbCwy44hiRQy8dVZeTjDG1HrTFIb4qNz
pHnLHzpr99TtMPulFCaP1OstVoE4ao3IPsWDd2NNEEXYw9VNNpkaojVt8hMZExSIDMo1JmQDXEqD
MQDU9LUnewFqZlisqidvLVTPSbWam1Z/jcBieZKiI1/XiaoBr89tqnH8ZE5jnZejEQW12Rt3BRUi
qhfLJcu0/OQMXpdYjc6q8tk4f6Si4lPK50S9UxZcvepi3EE+EHO9ULOMo/czp98/QAtDsWDxFO0q
sOTGk89fTe7SynGHzOMk/489PQZ8NKtGr0SzDeBQIw6Uc05dp9oNB26LFGIkxDotKolVHuEoPn3I
wBiQ9qaM/UHVTrdKM/FEkGpA7ZG1H+WGvUpbYcwWP0GF2UcgO3xKyyAqzjr87WiQZ+uu5+ZOcFP3
Arq9dXRn7p6joi8tyEbhHLU65HgKHj+jR2R4zC0DLoP5Dlvks9ZrkEPr4aiP1o/PMyIch8quCxxq
yWYNx46woh+xrDWsq7VPg5Z1fDcfGnRLzpBZ0eDmM5cuuOZBRg4meIu4NZqkf4w8FFWnOkaTokw3
B+r31bd65JPGdMyABYah4f4hMe21E/ePgeTFWBpUNkfC36CM1rInmX+Ot1xgC1mRUP5iwVjX3uIw
/mz7CAzXvrZnS3Rlm4X+H5GDaepf8a05M+lNDaLAjlfHuAcU9laRrSlhAE/FrGzFrf5XHuXwVDGC
9gXCjc2CpUp/34vaLFx33rsaKQS+YJV0beVuHneMjIApy3Sj82L4GDIzXrkEPP0GdKZrvBgHlXr5
GZp3JaKkV6rzGdVrxfMW/CsBFyD9wp9KfOpM32J2fJmJXhpxWP+gtDpLjBy8qrp3YkUcp6CGCx8Q
Q9zPrjbmq5sU4PPLrAYwWOxphy7+6PC9CF/SVmsih5rlDxvaw8VuXLypvZSn04+tcf3Lpw8gBWrs
WIhFdsqMe5ZmBIXeqGvFMiXBzsx4SOLKsQ9g1Ot4XA0UUL4aOq349R8QshsVbUJaR0a0M792mAo6
lqcPVbnWEn+zaZ7tW8s84TXQau6vOR+Hahmjaofxx5qnut2RMK6eXqYee9+Tjwt+yEIuXg2g0uHB
hdihGZzCBV1uhzTIkiZqe2n5cklR7t+niqtDRj3KkfO/75X2orxWmqVmEgNbMS3JpJgYqfHvHwaV
PPpQX5x72+EXGaqb9yuTjb1oJ091CGunUDNjH2Y0USzwouPFXogO4+lVJoV/3O5O3H8VZl9Dw579
w5z5AAOqoatpOIitGwMJT+KGlRGOy0dH8oLKW/gv/PIIXRpZDSk0zrckbrYceGqec07ag3+WJqCN
AaG6497XMfmqXHmoxy8acCVv+JjhHQlKNI426Kf5d54b64/GjCScoErSsebA9OFE1kuPwpg6qqJU
Q0HMVC9YwdG8CcDOnZEhThL9JI5N+C6HS9Oxx7LgB7D9Kbkic29/0udQ/NNCkNqX8g8IVJmTSbaY
Vsdhb1Dutl6cLU7nOlyPkqgy9cu7/3f9qqwGZjaiMtvxMYG9RSR/sUhyvsgUxlTm5lK8avSsEfH2
VwpgIBQC50Rgvz3nKMFs+nzpUC/8kvSB984iYf9tyh8PSXe4WH35mPvsTVYCZ1lLIaneXCkEfofP
y1aiY39z78s8idTOEl5V6LypeiCOY0L95YQrYWLkT1F39Ooc5IWExiF9EtdLpAwTB+k6C3Hl+QWf
eVKsRG9X7hsEJvcp1nQSNL3sP3qmgaeN+nE3fUPQpif2InSbzZY+lgtEDmVNatlD/RnUKcqlh2cG
ch8L1hljxIRyUsYQTvwnInDK4BPUrOwQ01/iImVSbhR2xJREODF64vH7H7GaWYm8oU45H8uurU5V
tt5P6VAiC5Aldr2/Voj66ELnglm7+aL3MsVh6Iaw814NR1gRCXWNFnzFA/PjCRWRY+Nkwxg5xWW4
Z1stEfz05bXIpOVoJBGgLTdcClig6irh0yYxZMgrNl8Toqad26uVsSpBysxZBUajSQCZ6NjEEdDs
D5PuXdHF+Kv6ygzhr97ndpQZ3s2DNA8oVS3lsinW4QwjGvrQxIvKTB6WQD51T1v+ESaOD/U7LHwA
M98wisorSu5jkU09EB65IeqBqXHWh9Ehblc96m8UWcWMz6mjg5bdctY0wNawzwF8FacxaURd3G+M
lqjNl/d5mlvI4rGwx/Atf3rhA/SPql2STF4/LK5EWn7lc0jT2bCpPd361eJ11uyMDCjPy5e+TGyR
FI4SLPKIMB1NR5Shid3IXP8+1CGGMvMDjWWXmnjceSc7qbwHRwq6rekilICCB4UPiRmHna+2T0oW
Od73beemErKiVjb4/Gji9y2VSFiFsTMcMLWGdvmysAKkHT1c1zn/kEfzcJ4eU4fB1ShHiqAz2TNh
Rfp+IkrX6RxaDVTtnk8Dalk11H+YqKxXvQvPYf2IR0ROOjoaStGVWjSVWdGMSHlRQYjASrN2XLrP
+mDH0x3WHSUJCN2tlfUf61O/rNsfadTkgjjF8yn1AOsIJJPwKpuU+qXZBRBZVd2+xOFOvDLB7kqX
Ug7jZalHBySlIgDU/xKYryxADiSHJGcS9AzUuLf4RUqSo4U9evvPv/r7275X6fYDSGAv+mX03T43
CHwwthh8F8gLC5swRevPxbJ6DQvOyyAOcneOoQFYYEi3DeDnMSC7C0mXWBRD+C+vvh/S9fbw2uj7
ruc/nLgn9MktBbBRn0iDm1A42Qs3raa93x8zvoIPrIu1dF8M7IW30dZI2acYFAMtHYRhptnFO1u1
lnDGe7zZgrwA661z1SnR3ZSliI0YgeGVg1zdzNN9qZ8kneBvaUU/yjE4Hg/JsTMjPWM6pYM+NPXK
5a9H5Slnu+H+OMNlhq91o7CNS8TTZV3WIDr5AY/GiH3jH8WDUHrmABgaBp4pVIjcE7a20Y8/MHfj
+AKDlfr+aZqh9z5L5Cyb1oxowIGJVZnH7z4Yj99z7pXmQPzsaMHIUcqeMwQq6hy/NRWKBvzNaR97
6OtRHRcSq7aOd/QAwKMriJ1/V7JBm82k+5AbdiITbmkr+M5sHBOGhoXTszAqjT8lizNEFS22Y1Uw
7VlHoLwyaO087ITH++qjWc9hX/ADrJ07zxUuY6IO9JXzn/QLr1w89G22GDyHDLcaxj/kRfaVjwaz
T7A1NkdzP3IqZKXfo4K/2neZcp8/XiFNJ2ZGgkYTidKwunC0QbY1ThwJrm8PBF3+jJbRUS1AbSfB
qyF7cGuugCg9X+IuR6acJLP6AAzjrVdfWgHUMBb9Z3+KQSsIs9/l8j3iEx2IH+DbT9M9PEOn1JzA
jmXkHV7CzYRftMzuxoaw2+xuQffFSKxsYDqKykHVCJ+Ayv1mDxPVlRsPHcjTpWYK/K5am88Mzl/p
RM7wdhe4W2PTF/cMkrO3jLAK/IijDFyeYGAh2UctoUSbghJTRDbeWEUYgE+Ehlb6TRI95bzhszaH
L8co1fRfRmhGw5RMZnkXbCrfeNF1lP6XCNAqIql28Fd0jEv8g3UfvOMH2XKUCzTPlZJanx0mN7G2
O6V8X/SkN7cUulgGSjEDqQFHcbvAbJnGq6+xXYzJY0Nd22zRVw75cyFQI8U8uRG0Te0l91sOmakb
8P2ei1nsRPd5uHiGlds3/qKEroD2Av2q0j1pNzdGzXjUWd4DYxYliBCJzgv9zhSYkXm57SgJw/bK
Jv3KjGRI+FRSD2CxVkTXSf0BXJt88MBhsjRCoK0je+bvuJmxVg2FErUwSr28HtvWcRf1+QJJA2wt
/Qig2kn6u9pPDmGLEVXmkhya1im+NvSjQ1aS7Xm7LzSTJOX7SIqVr9p8EQLBAHLnJG49Ty5ppUZJ
tW/Bjm+PFo/HraEVNLQdLBRmvZzT/XKxZSNsI9XH7GAfs34oNfikJxnufNeiu7MV+mmetLzFjTDn
f1nr/1Sd/2iQ9jfv9hJrbC56Skvf7RoTzjzQuZP3quIuTxyJ2d/vtzumf9JPVYMHxzf7wrpHMHfb
VOp5uKe190jJSUM6UEVFVKCe6lLB+gTli35AeXyy83G0yXxQdPMOPKgJAKmNy1zxYnJILzpfPoqx
+IEwDqkFbhlAqgTwj2AI3g2AvgAq01WpUcEq9EKJEnAmvY7Z2QPt3BnokI3ByS3M0RzjH9fVPsSK
0KKOCTVomJN/iwDGOmtkJBZJU+f6fVhcoPgcwbJ7jI+WP7wU9vwYmYOpeXDReFtTyokaDlZB91dH
B5ysbZVSNu1AA2N2kLZ+56h8X1B0OcA6yXz9ppuEuXz2tSNtpS4rUrTwvQsWTTmAQ47n5ZDorn5c
ulj8auuyjQ6zYf/oWXVLUrQ+XQQ+3N8SDtClwU0Uv69i4OOYqzyaJlHrqq70Xp1uYBn+axIBm5ht
oUN9IM4NWWuEM1iDOcCL5PmNci/qte1X7KUcxv73ii0GNB9DvQZ3jaffx+bNoRtUtSx87VpGqhli
iDqENiUPwiw6i5akHnUHVDCNArjELxCouzsisyk9xIRqIsjkTmDiEhDKN5szHkr4K5l+U9f5c2wj
fW6f4E31GMcMqVJrIIx1EUm3nM/yuACFnMRSdvP6yOROBilWz2q92l/aJXmYy0TI3Unaz7MEdd4o
0Lhvaq3EZZdTj1WwDXvRWngzNBVwykaQIxgVHJLBEaph6k54C8mxfZ2gmhlZRbqIC4RYk85bX3fg
hFESawEB/g/GA3LZ87Rd6CpGsCGcBXp+PihMGyzWW7UFLiJV77nwNoAUl/rq91VvIAqDSAXDd3cg
u/k6yjC7BVranIOz7Jw/HuTeBv8F65d7LiUJlozkePnQ4f81uM0c7PMiseXRvsJXn+X2lLLgnqvi
1LjDNUsAZNx5t+TgN+P6akzgjdQjUi636d7xaHBwhcbXe9U3fqxVGq1zhIC1tM5GPdnn15DVki4p
PCtGTsTye8RvthWAI+hDfCGf3KwaZtHKbR7aJf/ZagPNNovpeFwD9H6WodQEo6OC/pr9MvRLa9VX
uSZ6XWWKIlLZnschDaTxU7AvIamM3rv3MmznCfLh4AJ7BaLAmddVD+PexZpVv0VJUyzi96u3t7JB
U1UJO9PdDrNwHA8znvr8huyhjOpJcSCIGhFTl+X7IEwA7UClyI+tfdLeRW5h6MNPySlIgloWYT/v
C7uPbS4gd0qGnuMEpBHevUfhjeb2XAcYfYdTrqh5JqGGQ8uVVEojuroot6xfzOkbs7ML0GgtzX7f
rmV67dQdT0f1ztTtZLIbHDk1ettuC9opGG72yT68nrpNBP7fsUINzXUwArnUKjJ6JSOpbusmzb69
yArRhPSI+FarEsE6dwLQ/108+S88WW/5GanOEIXn6qi2Tf1viMal8eKZTbNsWzKkeWGWCVe+Luib
sApgWT/9IkzRs0GBSZGxLm2N/HKmhaHF+YbqUgNb5xC5TdoRhtdbQvOWbl0YJCaJ6QrG8LZaSuP5
7ITlV3LBwLPShIbM62zxwF56AqgDlmj0u0dAm4Z7gaWZYUrKf22nDciJot3whoM1GZ72fhQPriju
6Fx9gGKvHkAJtPOsle2myRjAZ/tSv93DSNwT1V2yTeL2xBysWJ4iPvzoT55te7oxN9aV0Sdnwc0o
BgX5JKxwYuC/wW82embW6nLwSGK6c+oEnMZxJ2rH2GojN128DNuOWtb/fTWfI+iiBrY66hv32oqY
j70ZG6GyEFgLns2fy8UJXYYdRX5bg0F79uiznyNw4livgDkXnJvMsKi8MVAXlDEJvre68Dy0+cZq
HydFgvwR+XT9/EyaHffNlpIu0Oc0lCQ1PkfcNSXcDlDLIGEMqqIHeVZ2UtQ5OOVdMP5tOrgCDtkB
6G7RxJ4wqjMdiUFcSeeeIX495GoR6cL1z/W2DYoxGFECZEnQYKfXGEmqE+9yJv75T0s5ojw7USMr
kbb/i5uioRni3Z6iggKu9jRFlhJSQWUP1Huaq7ONtCFr8zyppUR1SeGTTX9FrFt/ZhNINJ5txPZn
biIJplpycjTNV2bf/6C9S9J3I9NQnh47fFGTCO0EzfIII4JKuYEzxwCOe2FDus3QWDgQkB4PnJpS
brifOtSF8QreT5O5xrriISx16QZqzIyk1Z/sMwokPsw7GUL7Zv5lgFfYnL0n4FYnlt042V2Ptb5f
/yZKWBO/OD7Jn8qOJ65Ce1n62vNlbpig2ItNWMObH9vBA3uB5brTRogZax/a2m8R0U/BIyIavZOQ
7JWzjILjkbLlTBSpiky5sFeZHG3W/lDBhM7vKy6j9vnLNmMyCg1GKcFaodj5WRgVjBuy4YscOFdS
cTzlMxcP6w0HYrgORcQszR/DW7iTZKvmwDylr2hAz12Llpx4gXgJDLdD8cRJKzQuKA7M6MWjBWd+
r5SlGCd2QoMWop+0RfBkUCHNR3jvHxg/vGFEOje0R4OnpXJRuMYl+eAw76BfZIBSOeIHzEE1opNT
vWfs/KHZtfpKRAEvzpn/h0u9BOuzwTO2LP1pS0pWAJcvQa1gfUnCPFHKzQN+iyFRe5qSWd+Iux9y
zPQaICjpPq8ZZzhxgiRPnx0V/4Y8kHZWU+pkI1n9qCXbAVZhn93XP4il5TZ+GzOWoBBIMImKvU9g
2WeoaLlArmm6P41mgBlhYHwXk2HqXdS9W4cUO4HBZMwOHlMvECrHQmPYWhKkKf/KF5EhGclK7kdw
ptFtQnXPPEUcHY64zEIkhIlNEa1L4tc+EDKPx46g+pXGkC4eUGaOGHlG+x8Ct1b7XVCitXMeNljp
3GkoMv4S+Hvx+74e7imdVIu+ye/R7G4cJMSRJUPE5bxrkD4ZjoYPZz0xjRpr5oByy96yJAxaQMuq
qIgKCJNex20j9iTQFM8zSv2UfSHG9OZlpfclSPN4TvHQFridKP97yQEfG2jr/NOgUvlajSWRhP6A
eRJi1yEgAfMRUEEOjTZjrTg7Rlh3tLsn8FUGwLQZwSm7hy/pPEvqbVbVnRuBayN7kF8UizFW1GUe
dDxL/U2BO2I5Gp7SZ2ZnW394nTtGOfX18EkA+hemad5PI2/GjAj+VZpRbYXKmLCyOCHHjcmOHYdO
4ezD6IO3klKWLhaWA0etin8yVH/mn141fqZBuQLxGTXQDcZ8tofvqcocVBO2+fGCxw6u5DFZnMyv
AADDJ0Uaxwb6cKbrOxFUp5ky32G1H7oS5uogtRwnvD9CnABK5PUnS7zq7G8gPt7idk+XH3aYKr+u
ETNE18ut8L7iLffOlVaicn9GxmkgGaHVJ90i744E4Wif6K9d+T8s/Hmqp/HWXbQ7KU9HpUvZhV8R
A9OMd6IMeJP+b/uMTolIItR+oH6C3J3qFUjZiBdikTeVE9Pc06Jar79LuoA74MnDOIIAtjBSuwKi
iKepgsOl595TtXEZPIprbSsnyDPbY5ZM4zAJZACowqIzywJJ6za6zyeh/pOl+hI7fkmFEjSYlMjT
AXcOj9ZkW2r2heZEw3LK3pKXE73nbXp2BwSEJJ69jVmp3Cyp7KchF0meQnPRqm7weJVExDU9jH+Q
zYPgYzRIYWHPKhaf2fMkGbN31n5v+fIOyD051EDjbUtvSv+WGoxq5Qxtfrs+wL3EHFcUFzPnXfk4
4TCg/lSCD+85vjECJV4CiPVSFvw2/hqTB7ebcQfrmZ6lw3R8mL6p/hpO5V2ptf8MZEIC3294YqHf
+9N7E37W2yMA6K0QXGWTeaZkqtVzIKwKSr+lMAgL/gBcq+W95RP3toRO6JEacnQvV0yVPADS1npj
vWnS3yOWXSbc+8DIFhlYupi9mgfvo7/iC3jif6mymT8ba66gJ4L0w+o9L7iQjpbyQ+5V26woZBOt
VVvvSFpOaDiQC2o5Qc1n2U1JTfwx8Gv8F1/cbiGmBRSAAlF7SjWjOACLTrEVMyV0WKEMooQVC9YR
kS4BxB94Hgzd8hfzBjxalgqOmpFj4cvoqsyL3HsewDM2OeFfJahJp+VxkHyHLQHwLhnEzqI9bIA2
yO6GD4Lj0yaKoPjagauruhHSzszne2N0lemAN3pW/soHP7oGe71zSLGZMhuAcQx4NeT0I1kswX7G
ziTGa+pjhKZYT7cXfpkTpyhDREnv/Yje2Ccl7hAzVC7YSEk/BPDzUIIOeHdpYl3yrz8eQVksZbnk
ALxPW+QMvbBtPEJt/WhwlaaVQqtvtnitUz4dGHeiSahehH2XwWiH9uMJm03MTFloNvFGhXMUHZYl
BM8bCcEUEYvjnoZ16dr6IPY2KD6RZwSqRbiJB9C1fzUvPMj8aA0WZasNQfhRvkiFMJGzFRdPP6vR
cYqptZokxF2RkLcKHlxyqSgjQdxoHMzc92ep8Qm7BcU0yf9yhOQc5PPuqeMJkjqiBrP9GPvaq1T1
pu4qlrkgRy/1I5FtIRC57I8fNkc6c+wTKyOpkcXgIpNQIgEOsNK1v4W11aiqL+sVIyhofgPV0OS4
fnAMzA2pKbWt9Xxg1fsOQ4T8xzQboEcP90P8IPtMSwqH12T2/4l6Gl29kED9TAHVPCTZuXAfRmhh
nz9ZY1LGMRvVVfVJPY6EOXpb1gCZ9L8Y4eCi3dO+1SzVaWqvHlJzi9Ght+FuAErNRmKtCGd7a0IN
mkLG8WJT2yKYCfaKxtP0p+7Vk28aE96HoF1cY96NtKe/mozVB4DVGL3DUuY9h6a9UyAxSNCGQqjz
P9UPOU7Dj38tsqmSxuiN7hpHDTcbxqPZEfmTnSGQrDJYWATUTlutIakL1/6DbTwJXZ5d8mSe4+tU
bj9VRwCoCN+7OMswQDeeYKYg4qTzoUPCwMNl+Jq/6EQ2ip79WIupAyw7f0MRsB9y8uMTY6WVi20b
jiQ/reugkcx74C7kfcdMrMKSKZbwst+mpYbQ+jgzlOtaJoIWnJL+i4XK7nLhtuzMjfUJ5EZHT/ql
rRNXMdxU8qhEzRseLg5CCi51OX0EJJqdqdmq/28WSZT7d/fzgNsUSQtD9wulLl95pveVQQQ1zBAM
Rsnsifa5C3Hx8rKikguFCJAPBL/y4/EJCQPScQ0qJxAo6DMXnPTP33LMb/QSS3w/I2iLqhmDQkCK
TVJkQmn1on7LqOoof4CmzHLUfFUOmNsdBjGK8Em+eDtJEVlWFxsbFCsCLchjHH/3dMxKg5p/xTF0
Zv8c5qX3xq/4ulGslI0OnxIJQy2PKfpOte8mE67ATzw/JGq4auql5xBpg+MzRI7bYsKue76n2RSr
EoGFtj43VRy7mu3SXIB///h7LU1kmxt+ayRQOpWpPslLfI0dO0/zjITBA5Z5WggOoGXz+tDVQiv+
CMtagaKz/mCt+q52RSnRq+VwIYw09xHBYFlPAGocrkF9qQZ4Ch+OwJqUJoUqAlXO6GFeKxH3fWHt
QoboW7lcbxvhciYvHmtrdH+SlxbT50xaBhpVCpB+JTRpuyNQGjJeUX81FeQxVnTcv2R6la2a04ZI
52NNlLixLQtMtqL3bJiGiUbwlGCHqnMmMm2GVIKFabzxbHuBriY2COgEAFHO0e+mMAKxbjdBUEfe
GkyWRqeTWKNVbp+AVsUIdHtqbJ1a58oG+C3JM/RkNGjqzZtTwDHdRmz5NdXIPuprnnfs59To2jfU
xlDRo7J7Oz75eZvc8WLh3hKEMYiHb+7FG/n36h18VdtTI1gjpSrtAf6WeCURMkKCH6B/k1Zgi5M6
m8RJt5OsESEBre5e9s38PEoq+enr3Jn+Z3sf7LrxtEnZyjBDU7es/Ex3l07mw9KtHj++0D75BKyl
y/Y0G1eJ0x47pZC7EO90Df+M78hRcpI8zXO8DlWgxGWn35lKPtBQ5DE9yd3yi9MG2os0eNYZS2as
wPR6rj+NjKfT+03hqeuB0q5OUwzD7AAdfR6xG/9+Ok1AsxTygC2JJN53eBFjP6QdbTu6NjcFB/rW
1V6j3zHpR8wIHExx7dJbos19d/gmdgqmT2Wwg/SCbQ4nQOZdW7nx0znGAaVYYGm7D0+YobmTgf9Z
unFhGeJkUJqF7dUSSXIev1/k/x9vrCTuIm+P9Xj3CvHfte9kvOENXRM4YcABR0pbrHn+xi/2dQ/w
AGvjNCi986mC8V76alqpf+GI8KCr7t/YZVddsHceA3kZBP8gJuQHX+W764ASRr1ofs/dIb+sifOY
otLp8rJZnOgY9ywIk1QAh+qq0/mNDVEFyYyx/McvpSB59Y3YsvVYWv6m5ABWVbQcy0oU1m7Y/ZZK
8gWIfs8LHMZGaw7GQIeXxrXJNR0CsvlGQWXHF7ua5R15N7wtuo7Fc39IBsXP6Aw31SVzxNxavXzT
zpJkCJ5M6fewx4zpsgDjZGd4xPI5ln9omKTvEopPtvZ0CNXtwvBono60yj6f3wVrBoJhIdFcnvQ7
ft3eOX1I2Z4N2lq5L1gaCRLn8KNUpOWYDVd6b9AbYu9pj2prEgt6K9/VQxbRrr2MRArsp0BO6hqP
lnzseEEYZ9GdIgUkOKHAW8LEtNhtrtBXIhXuzOfazHAGkmyJ+f1K9416qvyHw4fIIJihyG8hFjcG
TUTjGKyjhBuPIi7RXOwsBoYk7VewH4oeYQdBSBYOo2Y26ZbcZqcPWPopa04pHH1kcOBGiC+vjdjD
Vu5CUp2yk8uwcgoSfVDXFDXNiyBOtqimwjFtutv75ISjQl7d0w1e1EdKJZCEX3n2QMqFef0RONx6
MBYaDksMns5mAWM0zOQB4WgV8vD0Jl1BnrMG9s7or5Lt7ZcpsuNnReL4KWrSsH9PdODyBMB+ajvy
JB3rc3wcnvRlChOdFR9/rEyLKVq0+TRTctvU/5ypmUVjlBbA+t73+Z1SWHh/C9owMvm8eGygtX6D
CwkIiN4TE774BKMDlpzYzkVbCd/99K+HV6sQhFgd6Mu86tKWYh/R5cQHQR94cDdvKMS7st+QdGyQ
7lEeUPu6xn5V+xfCaCvxvrZ/lh5v0UEEdkigJAfdaJ/u8ycKi0SpR1bsR3PQjdojN37akGwEM49A
nr0ChEtGiMYgehQ9746paroCK0XBdqimye8iaiU89WRl75/JcTcK3u8WVl9wbE920Q1l3I6+t/eB
lGrgaQYmq3gSzdrEtf94RekRTC1jeVit72elHInrut1yktqoJc8ej+MAnSLEe6BzmXbudd97a53V
lB9noGAlkjdwccKVlSHelc1XtMGenEop1WOmbW4JFyONf7H5Q4BLoVwET9jU0AiVTqV3ajsLBoUq
PFm9xR1sDd8zN2EpoTRmey0mSM/ygCpSnYfwNqr9oam7XTvzcsSltN6m6FkHNSmEl9dzJR+WJk2W
O8vHvwQXcrDJq/0fhrWkzcm5FXTum7bTEuTyY1hHy67t50UQRYbx7tnv+OE3ws7ubXrGjKJaL0mr
fHPznbjn88fuetcJvEgeS79zSUN6bWBcWku0nyjUumfP+C/NSvE+e4y851oT2AzrcIoGmKYJhGJe
UNTbRQPuXNn+z5/mh5NyTxzkQi5ht1TVtHvZJv+hLnpIKPEudxO7AY7Zfba1EtupB7XnTfcQkOAg
ICq2kPAXqYvHB9AhLAy8Vs7DjErJT8HyfBubInIVN9Acij1keTb83D+716yI6aKUSc6MntHB4on2
JEl0mYlpfsHoZzQT5sRB7IK1FvKVGS01RfBqhIiRkgP+9XAwg5W35K9Pim+5oVFKS462UCHuyXRo
WbJUgdCHTVdAv9D31U90KwND4oaq3YYcNKjgH+ryJkNq4FcWS5NHPpfOpY43PK5AC3SMy4H3SF0D
43Sb0GfJ1jDiL44qGuP/E9rczSMLVf252imttbGU0na5/+/qzM5zsb6ZaYu+aqYz/1yrJfkwhtWE
WqEjXWt9gztGVDUy48bKyrMt/GhMQaedNEXpV5pTb1cikafcUHbPPBWsI1SDOG1SeHM44wSvtynK
CaErZcbxI0BU6DEPH1sPLewoYHTy7XgU07kkKt8hxpSTyDDeozBoyMJY6MwrggSboD6U36lYru5h
pgM9HmFagFRq01+qNhyBVDppYDYvBiBZRfpn3SUtYdMOiJLyxQbabgry9jAPl0fpXWARwR3EaDmF
DGQEspVO4V1M2ptNqrXh1fuQHweH34gdAojkb3PQRzsxTWHTyZSoMzQqW+3zKmqAgGQzwLAFSVmH
FG9UViFShIVYJ0wru0OH7DcIdrMlPaPh2pjyqxXJ5Uooo65FsHxyJFf6ZR0bMi9x5NRUHk8XyXFh
5ok0I9UnaO17RTgl4RIjMd1TWo/RpR/tBWgWPPOapnSUiI1kxnPzwrAinqYXixwPDyoQOlUdjjbl
OcvjCUU97V1Dw+E0LlZyQ+q2BEwYwkXVb9nygF27se6d1oA8cwOosSfc3H3gB1pKeG69s0bpMiUh
DegYikQVNkhoyhbTz9hglSGIKXoWt5633dtE43LEN94j/5z7fswh8+k22uD7kBn0rZ6uPirjOTIY
x32XaSN5sQfgjzaIUx1rqKC4Pf6n1Ur+mIL5GvG/qX1uGtZSYDLTIq3tQ9PyQbbLB0oZvxg+/jmd
JQEcegEGmwn23iqWspp1IcSBd+rZjZhJYMfqLCVV7/m9tQVD059eFbdQoMbnxrAeef+c80YBDF8M
IcmmJyVOJFGJYS4oz3dPnSQ8DCR2pABTy8xKSd5FHEsyaGHDMTGrNpd/Q+1TI6TScvrWu0PdBLXB
1f1YrwbdPw/QUCxw49EJ6rGM/8MEPB8+joVzrYqyMZrwRg8rdh+POfh8wrzgiMUAGDwKJezNkshl
l1HqJ/HkbGE8pNNhTV4yuBfPgHT88XKSyRA0FodYbTY7oxm83cCIL9JNvPZdZGe5S4qehlaWm2g5
PxJcTT6wyKijlz6a6kK1/l/jX4DwKvz3Jn/vteArpAMHaueluZ+vYC6pA19gMCdRohJDXN1hqxdY
cmOLc13f4xPRlW91F9mXUzagCbebcwX0HuNbITXXzS+HgUXN0P0wDrwljBu5d9/AgLjMwwkpvzke
pKW9ERawzBF+w1qBbG1ByaiVlnwgHtyZEdGomR8aOCRmK/oijlzXYMRCk6bQvc3BM31soFCxGdWO
Ey+9Cal7DltUEmRDDnsRAar46FRCLNN349Twh1eV8etG6UXLAVJnq6TCjxc0SHRltWJzL18w7uUh
KwsvCzWtqzrtktEIDbee8ljvNTQIaKVEQAUaEgitufEPIONVvWCY6nDFPHzfI0e7skk7+jioA9Qw
T9E9/g4R2Xph5PTflw1OE+KVCEp4gbKN5B7TIXVn0AzaTlh4v25RstxR9n+H5Xb27G7j4WQdI+VN
XiOO/NYds555wdA3oYu4uQNqZUb8rLEhRxjHavz1iXvTeA3aARGn2SrbxFmFyMpdP4NoSL8P0sC8
nPUxbcInWD24EAbM2+DucFFlOQYRnGytP+61OU7Ic6WcZwrSMngWHu8Gzuh1R2NOo+uM8lnDPMjW
XzwTnLgoxda7ikttV7M9rAkou3D0Um5fZltlRpPNu9pC9/3n9fXncgO/WIPQIWeSnngxZKfSbUOm
XHswSgOboOzieSULjyBdZzE/qCyUcr0aNDTdy2nV/C11dLoZ3mOUqoUpOar7vl7yKNquSrz03Gn0
1FRnuk3sfBJjU6W2JbikrlCWNMz4xhuw/U1hIFEgBlKtQ0VHxSb/20QXe+aIJMu3Wy0ot0FkbAwZ
zJKErj8kjGr64MQXyj96LyDXAhgwdAQxH+5fAQvpsh4KK8e2le0ATNNz5j6vJC/0sAaypNHK13tg
9AUKzASJRiXAErEJ/Kzcj9JVnb51XFZMxe2dz1TkagZARjhRR5h9k3cn7Ep75aS1p4bT/0A8FgsY
B6T3X4jTstSt4ehifeV6FdJNYPxzvKsRnrveBfjrwwchP25GmfZ3Gq4lO5sIwg8HxvWewivIOE60
0iqxC8kYlLfL8SfhTOCx40a0O0C+audmq+r2XCqpwcqqlbxgg28Xrwg7NjnpK8f/6nB+OBiH9zYm
0R1gnYeJhEjfGMWYdz6o+xMvIPa0Ufh5vtCGmvoAq1vpELnoXP7N6KY1Re+7mYbeUsZyydObO1dn
0nNZy2BdDOpNrRXchWWajm/el6l8GPhrB85jxmUHT21BDPM+jnM8bK8xADg2OtUJ3r3koDvc4BFu
f/aP3yJlevJcHKGv74mHFdp8Nb+zean/UA30t1+y0efNN/ke28ZnAe75eeWUiehNq8Hf51pyVl2+
7cK+RSGO7wEIX3xki/QlZlqnWFahWvx/qKUKr1xaHgz/kjnl+GZAkPJtRx940qhdmc9v75AlGDSe
+Z0AjSgLXo8/ZK9OeVDbDqcKExvx3b2IEngVBU84J6Zj+XGC5aqsBhwsoP0d80zGXLsceLRlWAbA
N8WbRysNAr5x8FehcADboUHWQSFXOKZRkxgOgM3J51LiDhtw/aZ5oOnB3OnxOJ1G8MzxNx2+gW38
FNHzvm78f+fqd2CLg07pPtWyaaWsmwf43RCK5aHCYz1a0HBtrzhJ5mOdJeEiXHd2oauhpr/KmX3H
ld40BvwrN5Iiu1LOD2TbpuwD9PXyFAQ2hm1NoV9ZwWSBHnfVWRgJ1gUxhpTSo7Bv3ymvzgC6Jsn+
1QXqQVhQ4GVOe/WEXs6plqbaMQqCNndVZYv6PF7KDkuP6dgKcILIkW/by1NIHQxtw/755J2lLnEH
dj/v+Ji+EarR5QZ4XhaACAkYpz/MZ0VXhqSFddUKsmf8IhUpKpYv4z4S9PN7MIXI6zqAHt/XvBoN
bP05ncSeFHYXzNxl9ahMBIAzrcHu6i6+4r7Wy4nCbFQqRrfIuUvH4U23EvOkXrXRdugBTtghoa4E
YV+yLEsOI/2U4lSCye+eb0pknltcVzE7FiV8pLEtf2Aa5JSuBmta0PeWkbNZI+3OtkoFN2M5Hzh2
UorrMcxrTuVOwdh5stz81fyWfi/PoJLgYav+pf2AbB0Ydc93e6eYOEYUuxjlhjgMnu6Kc8mdB35X
JSMiWRhzWr21jgEzlu/JTba6fnIXXzQQ4qPkIl8fe7Wa0Qhooj9BVejZYLLsTLDLdnsL+SrOm7Dy
PC/+CZe6GtB/KbpcERhPayLWIUXdAy1ZUNnAeo+jPiJxYNQSlFjUsY20gPAE8i/0EgN+XlDW0O8t
nO8RSAUzZal81IAJVdxTSWsQcNcT9PZfHqWs+1kWkyQaKRqXpjRoLbySkfRq5nqcU+lE+ZtRULfh
fyHRcM+fNaXsv33yEBZ79j4cx0jqX+HqodS5/6R73NdHpQd2y+EgWbe+4B7evtrMXGxHYxKhWK0z
Cw9my08CgV+DL7vDO2vUh5Ss65jPoBS95VwgpzHoXEKxURWM9qgaf9Gw4mLiYhRNs4uPeyuyLVOw
L2pU5GIOhMPTTnHZu/CKVQTSuOsnd+kO/mKROT1nzAn4wa6ml0l15Z1dpVQhj2uqw/5CrVp7ys3L
3eXVpj+8T6fuSWL+uBrwWB8u0ajkvsIcaqttxBu0Wj3AaLEFk9TsljRPumBjb6+JBoCkjfl5tiV0
KShffWN+4zh29uVmwKrO/Nnj8a5Tq5Jfm9z5YuKfQ2yH+GN3bMt844BElGzfJoBA1vLfgx1QGZiO
9fyRPBB46js+YCgmX62bFosKrUtpXH1+Ic+P+qD426Vs8S/TyhGbcfYEQJ9Mxf9VTds6ibGVr3n5
63jGi7X2HQue0TE1wNE1NvYHA5biH9wieSTUJqvon41GRCdJGBJ1Jyp32KNwfOG3BEGO5QBCRsHy
2Pn64NSLnVkgtK+7LHQAowUJz6wCPFpEZavJB4g/zN3g7hGxFiEKGrzpuXR6dpWOqqLTi7XgSqyP
+ljdeTm2uuiE9f9SVVMq6FVbxqzpDnLhaENOFJca/5DzUtAlRqIwB+7XFwylQgH/QJMSwn5j4jYh
2vtH+PqCz/vmWG+vLXS0yBlyIIhWJZ7Se4E2tX49nAPWZCimIJoyWqv56lTBJiAqqUvagoO90E8p
Ubvr21icvlfkEu+bqAltO82inoqSX54hWCkKX0PvU1uL7QXOMpb/PCgXqMfKOSP5RLQE2zuunZ59
0sdezmhtcXgfjdxG28KLCwLS8O9JOd4euJYjDeAz0I8o1ieIwonZgSnVBKpXxxXyH9lJYsbGDjHN
yE22L1gpAKFiMN+LYfgIlrwcVnHLBdfL7sDnlQFuUJhjRBliWMUnoq5BnLZf6ADg48TfTCoq9LNd
ttkP6EMfZiatOX/DHNLVtvKsPcc4Onu2ghoergJ5xgW8+s5OkpoOUdIN7BofZ+5C7WDoTk/nWDIF
fZM11V0hJE6rPQNURIZwzT/1DyBttJ+aYMuupQgtgeZe43uvrbrq+OvmKfPW9SQY5HCYqsqn3jCo
Lfu4OYeeiWdGFi8Yn2tOdFHLVMOzhH5u6SFBwYynqXdfJKsYql0sa2bAkrmh8N/mt6UEv1eH4Z+P
jm5ks8lfBzFWjfoM75M3ugagMfB8Ti5YxD/lJo5t6a63Axhr8GUxGH5lUwNQtjJ9PDGNuFHfRSIq
3tSCegrAN84TlURrEs4oOEnzP65UvXTuPQS9e46JQGzlUMu9tZAdxlGO2k4g1n9K7UyP8tum6ahn
YBrI/YllGBa45htHpos7mgWy0f6iXsECzeFoJ859oo0KAR/WAsWpakjrgnFvMD03kQulo/dolW8M
yC5wqVGl+k/ILiSmz25qI7mfuvw61EGYr/X0xQp4lyDR80z6jX/57NhvecwXNu63+uzydekv1OGu
K1mhm183EVn2L5exR5sVEUOL7wSLaEQC/pGxmUgFbGR/6ZbYJsX/gV7tygo6KP3VHMC+bzlmNXj2
9o+itxR5Nf0ZcU74UXWHE/Id3u1tBWsr0sQr8Jxubmvk6ZGwdtJunP/ytismH/ihbXXnNTDUCqEF
05VWVHeTnL+omffNpnsAsHSMuN2L/eCxtaLP0DCbUUzNKXe/tgZU+HvoiK3gV92EdfOE3yHwLDKq
+WapVbw4Rt1mVts3MaptERAo72JiQHmZz7i2Q6VZSwIqtsytyWGnuF6dLTSkmHjwI6wbTAe3Dh1t
FIkvM2kcO5xNaNXLagCfCy/UpAQ7R0vHK3r2ydqCGL3qNj7gg4JG3BbqGDcYXTkoH5PnT3zdOAhR
DmDUA1ZZD+sHt2eY+5h6hFvIk9aWWa5lgfueTfVaV9DfekFSuZoRkDGhpIWZuLNIf6txZ58r8L63
YxkFY6PXr6gA4AZXCl+nUt8hdVygylPItTyai6vnszFIid8CmZPcpihx8CChy1gbc8CSAqjQs4Dc
JDWg+oPJkQcDmJR3YdGR7wTYg86KUuXCxBwhhwnmQBXDqR/rROb+VrXpjqQSBfCHiM9OksOFn2QO
E1LVXNOjC93sK27v8yahIpg1spoONoDlv4tQrDU+QsFjxmvnADWi2nwMm5QSPjsNxReqrbh67eXk
cAFxhFslJfa4eTbMHEYy7CaJq34NeGfoCiX+ecHfRljeUfDOIOCEbGTQ4gHZUux6IuNBsDVhA3hY
ICpniz69k+wJizyDLt9vGgxLoxfNoqlb/kDJ4QhT8tUXO209Z4ovzmUhQLjSWeaKkxYJjICrCaZQ
MV63tTuStqA0JMXjfEkkrJhwfsv/ZVGmBt+0ZRfWOHy8BF7Y37O7f72Zoo665egCHtU28ezPJPaP
lsUgZRkJ6jSszDVoGhBWh1i1HR4BzLmplSjDwLQ7uQjoliZ6/Qf1bEnGc1AIwdJeQuVCxEAI8DIV
c7yRyQ4GldE3kpbbV0ygVEHSJrfoAt/+Q0XKQDrJWkPay7MLJQ6xkie9RDVKgICWh5zwOhADZDlf
BkNKMBHO3sGVt6rCdNi/0r6H39gs/ZnNoJZyDo6zIjd2w+JNej3m2b5uphJT3hVgsx569JjwVCOP
0EF3oUMLpnbB5pOwio1RfOJqHDMtO8D/cPEEi8fr3w1AsssTM5uG0G8Sm41gZxYCdY8RCGeimwP8
xbMNYdf8eLxL4AEpj2Zgi2/EuUXkK0LpAP5CkQz11CuHj8uREVEVG3qFWTwdSGKgNfZC2EJnK6/D
8fJ2BqrpwlaN5hjH65Upi5WESL1e/mQV6fwxKdw3mU177YePgqkoWiAElCXpMryD+MEIy7e2h8hK
6aymwnLhE7kQeI19USrSz0JuilOa6Dt89BVm7p9EWg4ugBtQyEBSVK38b9vM0HN0EPt+ppfk9vA3
zmyhKc0mNf9q9R7bdYPVU6ycP570iBh31ElHVi1iCMgpnsYlrXTISRTWfMpGg9yzZsnrHDeiOb90
TRcKHvnvx8uWuafs6h/SaapYPCy7E+hH635zXn+w0rgNnlTTruC0TgNoyXBlDMxVYuLqbIFw5WRw
4YsfZ0r8FdbdEW0D8O8WpXYsiqFNYLSPKL0MryNa97c6uqcM7kETjTwxi6w5l9SBKytpmJJlJT5O
BBw32ou/22lDEHLYyzXCz0iUIYM+S0pWw36zZXJXheXcWRNvTUgioXzAc40RZP69fa/TewFKHOuJ
ERQk/udEYkKKnsIs2nKMGNWQcqUXa342vX7xNVNN5uINazITKm3pItQiQQWXbCU/F38+m4wxCpC7
Rj+jL/uzVRueQU4y5R+Jajuoa+o4w6CiV1ioRqe4ddUUzrvOkHVvkSXbaxfa1YRCjnmZFflPh1V/
3/RzJDQqDCt0OMYEYgO+lHNk+ETyim/BdGip6ypI/4cm7ylymO62sRUnFhdEQJkR8TCY7oAlXoz+
1zQigpJpxIB6g3XCdtXGC4Qg3x/iwj7OM1mtYAqvGvHBpOGu3wfkAV/7VZ0FEJjyhx0s6A/hVOMd
R21zEn+ugtRYdvy1CQJUDS0wR5E4mwWbJcbkvuByx6Mh6cAJNl4jyRX6rfwywKcK7zu34afN6Xuc
m+pYf9aW9Y6yZn31IqAMiY+iypFFpRPDv8uwwMKklGcvvKBpP4OkFtwN5FIzG7FyOFNP/i6JEocC
FUQrmzfOWrv5LkHSc9phCa3Qe47UCdGGIFx6L7ZdutuONMK1DlWSuqIGwGzMY3LO26UoIZNozIPu
zcBngi10VATQe3vZbWbqO/ntvY+mmok/WRQc81KOpgyf6mfhSICOho9aZUa9uTzuzOdjxHNfvDd8
MXIFVoL4CB8fK32b2mcVuupBNcR+klOzVBMZx/tjKI88vGvyHErK2+QN+t9mZQc1Em4gI7UaXU4S
MDd7Ye8DtXk8ehX4zgt35LStzmtRW6jnZvL3MIupopwc6mUylyKmSjuTZ8V0MZJqXvqVWY8nwDfN
d9sThUKEq6zfIRObdFbTJKBNfu65erPC1y+IjOAF82LcBtMHrUetrGEq/XUhGkTP4CZjZIibYTlL
HuJRUWLDzdAsEaNjv8PO4InFfXvA8RZ7qW1hO6Qe4AgYuTPtWiNM9BRh8tZQRMOeaM5L5Jx0QGQ9
VyVLYKJerJdU2GXfy0RntsRymgMubedBkkj2pVXVEDR9MIUZfv2CToJIpVtGrrg4khns4JaA1JQH
/xJ9FM6knSoHrnzPeXiN6gAPqWgMpVwRvc50HSlniKQYRd02dNYkAPB0evXmpr61RTLibAWh96kO
ilyvMI5MASwcL/w1pKzKcdx0lVpwrIr3fX4/nMjhn8Y308Rytl9m3A/o3U5F7cRPOQ2YfpRg8nXn
SQPo3a+FWbssrK5zQobxGJUDg54BCFrY7/SY7aV4KASgqVO8uFj5ly1IT/KoiRLWrfvltyWA9Wnz
9ZboYLZuEkEjDfyCv9DkpyY9VPIhRFvMlqW7eHxKcLRnPpn6tpipilLYTtsy00BSv9pz1JMOwzvq
BJjyQVHsxWZVuVHXrjOA2sFcKsbLJ/d/MubXrazmuStSSeRE/FKy6N4G7dN36K1fIGZv+Srqshzq
XbtEN8LwUvCR6evXnRVGghaz4mRFmy659d0uVGbYNBBUAxUbF+kvVQa5ZOzYhr+1Fww1NMfgwtzq
/gcjOkoF5zJLQApWl5iPh9ODgbcZrHKfWwkf43zlxYvXhGAVyxJr4hzVWe8mPlVivZqMk7DYsyx/
B6zzOysDbLjEzKn4MXjS0S9v+weTyhmPF/ETYv9ns7E4PZg7mm0vYBdAPPxkqZkfJccAaV2ViIvi
KcPNCiYXJ+l4eEI+5aGRgHOiNsuazUk0oK2noxDkdV1eaoZ/EOxXo2fbWMA4FlS5uPDL6CtEzxrY
DwKz/Mb2nDWheKsg02XRH7a2vy2Bbh7Ng8iGy+HKfmN06mijpD+sQOKZ+5edY7ayBg8tXkUYwpwt
92ap2gWZ1LrCdZH/9bXx1yCJfA6ZNJ09p9gw6RBosyWmC2SHUB60YOazOu37J+lpCsGVxhGOV2fy
QXxebgSlgOW9gRLxlVoN5gtfZieZAWkoG6MGBIE6+Evj8NAarUeqvqMBRc7z9ZIywocfZh+YATtU
WzjxJ9Moc6h+BRnyBcr32f61OECIHqUcoICDXIJ1v0l8JNRlXPT9MSAK4yEBaYjp1Cjb6n3ui1vd
Jej9yihUFsRucsuTUUr9dfHLz9ZJb1hJhCqIovKAf7P/TJA+29z+iXs0rn1Vlt7OPaaytopppgU9
cCzOPoM3xTQK82gnI509yCNQmtsj+Z502xBfTQh5r9aOmoDwRaoRZWTAJTKwncGscGf+Eb3CnebE
7qHwQ8xh8aX0Jl7FsvHP7RvIyTGz0vAiZPpn2JOveMEHdSuzX8kVfHNLLdeSb0kFKFF2IBZdVVPI
WIyz/bLHcoM61AniSFVW4niB6XNXjxbYl33KXuMr5VfREFjdmDgEDLHoYuosDLu9+cgusb00XQ0S
SwXHHGjCwLaRvPl+xYeNhmjy37rZM/B5pEJC9I3mCKnT4FwS+E/s/tyEQS9UdYyb0E1iOyV1NnWa
rgjaHpqX892fQP4WkFFHwlenp7pgrEFhpaxzT2vHWUmxMtiKGAXJXBsqdZFYn6QM9Pyf814X8H11
QGK5XnVZt0rrLq6edviT05OeKpkx1lcDLdPeWFDVtEDrBcbJgTJTuiYGGG0YYEpq4utr3H9XcN0K
XKF9h2uO5XxdO+jN+EZJig73yA02M1eTyGLm9Wq7WKGen4jjfWbhA8cT+LpUtgV6O6rfbo0e6cfg
7a3ZkrZWDfxxJgDbF/MU8PUVtrnJHIPF88PrkgvBqFcgb+mR7YT4dEdFz+Jw00SST1bAb+/KNdIp
Kq/Nz+GLPtL4BgclW30HARHUyqGwm9reEL48JEAtci63XxqZljYWXDHbkEjZV7zJR8tiJqE9K1kN
EkYZ/3CRlcvGmoe51l7dUE02DP3KAuQd+jEBxF+nCGywo/nTi0gdbjnKMPffYmxQ7tP/EQI3QnEZ
ME5nFJ2PxJEWmprBEW92X5Loa1/kyDFhCnjUJ9xCLoUyUpJuQxk0MFaZjWxWiTb6FiM976dzOd8i
e/nBEtrcVcPUp2TiNVyzQtqPkNEo6K9WIhBqklqtZ8YxUnBKocoHblM2EX3BdYzgveQtLm5yrBtR
MzHaDp9OIb8MDO8pnEgGqhfC4m5sjV4YFDsgQioxBhTGjj39TGInMODnj2RpO8OFhMDp7yI9ZRAm
pGOr+g3ASxkZXYzCATVSj1hqpIDs/VI/NMUjJntRa643N7HDguuaNbpA5BT0sFW87cIzoc1EQeT7
GzAET2x/lYluSSzq3W9kJGQSHkziN+sL9H6QAhyiUaOLnR828eyCgZrW3/VFPCI4hegBbbd+/Sj2
YCkZ4FxL2N0TxsSP845if0wulAbouaUCNtUuwZzuR7TiFGG/nz+dff5zTCspJ3v6IFw7mxAgqqda
9Lct12Ela89RokOgWeU/wELp8dueSdw7F/8fLIyJ2Pa9MNJ0YRCXSZi6zUi0OhEOIeMWWHNP/VnY
tqQ8X1tbY8W56zXI9t7ddht/QmhDG47uplm0+ce7Y2fiQSgAT7j+jEx/2nUJMeVHtWHYgX/w6mdK
2+XioFg+z33k0RY2Bl14OXXpN5+dZi5uV+rYukNPIHXx2HBl9zwd4kLWo8fwgnpjXGb1Uvr+K0QF
lE5wWJPbMMgqs7pNmYmbauoiaGtvubACFU/FViJTpiV851PGPcQokE0LbWlOlQaiSAoSfNOgDFT5
vQ2hFZIrjqQmv4R/WFKuAI6NSr/OpNzFXukagFCIEk9cTc0rtQi8OBEs3cQjXKwrwK7FIXvuPwYW
2/AAIaQSa9XZ9QrWLwcfuqRbY9K5d925GHYSHL2sR27ISBtSscA7YfvlcHfSqzU6AatxhI3OUDiM
Zw8U/vP4syOxbMhg4PBTLzZ02cpP9/XfEFoATZ46O3dv/PYSl5pupwbkZbF+qePd4UeKtqijSiLX
JcOtuNRokFjWmUCVGbIZlmac5nWr9T6x23UG2sWTeV8Zo+9NmhUDR7P0EgAJwVQ/YPn7VPQAtpxz
T2Hh9/mEuh6APhwKggRaC1d55dOq0b0TaiTNThTtbSBf8nC9+cpMCPLZCmiAxwEPtQVMH8CZ2deT
81FFMY6pgq6jHxDP/akryn5aPSTykpqPIjiL4+r+ngcETSOCG2R3MfQox95vK4jJn01cTuC36nJn
m8I5GoeqNo+7Iid0f1NwuArrY5kSsZz+FRnz4jBv8rnn0YCdyNshyTnquV4sCWZfbemiygkU1qTF
zu0R3HU3CdLJKVN66LQGFDVUIQC39RiEng7mdtkrx/n1GfsOU/L6KCs/L85PUzSeJdG0C3VbaqVM
BJRbWS5L+xH8vnVaFGm7erPTAemOOOoGK70FOrz9sSVd57L2LaIFMA0n8je/3fK/zg5cj1K6jGFn
B2tmamELNtE111FryJ/MjFhtvDO8gLzR8i346pzTp1QpuW2Re+vzlR+8UY4/tP3nJCj2wWiqEkta
G3p4AGjFvxCJiw4SjNqDiO1lKdzPqiMMz5cH+Rid9RT/+cysErqsTLyjUfBev2R/i2Q+QKopxkNw
R0wc1Be7GYEgOCfGzb9KN/kF6Bcib71SozcesLoAPS1g3pOKOrrGMHUEykXnH8iVsH2ahsebEopb
7QatSf04ogSKw7ew6TivnHJ5CNzh4wbFYPnxv3HzPKS7kuoPzLy6tA9tacakruJyKV39524BiMWL
dsUroLHwyBKw/yXlLT1gxgal41njMrVZGLeMzPKTbabaeb26cZu6TKy3WuGwH46Zv/ivaXRokKAr
bbsxSUvg+beASFmPJSJU7FAzJhMXLkCwq94DnTUjzwxGH+tGKpHsmKbp/Yk3ZI/dbUSGG2pYAs7Z
TR+LjVfMjbHEL3IJD3PSFvqhYO+kbJjlnkJET8psDkipISJz4yomb1UQJCunAMqly3hOJ/wKz/iz
v1GQarP20Jm7G9d+3Ia3zZdrNmwLmKf/6pK4E9aa6Wjedzf4Hg4cQ5z9N5VGVvh62Jf4i7B4NQmQ
DbQs/ANIlyNkov39XRcMYp5z7tE2D+Ks9MpJqRaq53dlzP7p8DP7Qcs1+sNbfwytir8xpyxJXrNl
RxcKsCqQNMKrSMEtpDbE2iBhQI/HZO8y6vYI2gA9rhdTmNfvjM54cDBg2IpP8WKIuRzG2zCJqTXG
3ufRjMplFYr8tlLme2jZUFL6213M8WFVKxJLGZZ3ujqBgYzxQljeB6yTpLGG3K/hQnxttwZzNo9r
6u6f79PYiF22CTcBqmGYkWaD0GdFgEavNCy+Qn/FhkMqTDt/ladLEmlMSl63D475wds3mLha+mcH
el5MTB/EhLngPdleOuEdRgUUPT/o+45WdYORSHkPK/5jcGx9Br5/kRrcMspoH2zPZ40sP95Y6AOw
kXjCrAmLOEshhBlYdJIe8p7FL2hs/eqrYizVd+fgpsmcFA5t+rc4gQvZhrklJs0oYKCSBS+CVbN5
PuZaqU7VOagFD5eP/ZtSp9iREwzWff7xXrjbTm/EASnwiLQVnF+Zj9Mu/OE88SYZ36EBKsGpmf4M
yqF0coucQ7V12xUQtAc7zWk0prvIsBPL/y2CswcyMEWWtAfAH78w+X0PiKb89/WacwW+G3WEkJ+3
covNX+yFnBaMxGnrvNVJzYCwGfgqdzTSXwJa59KesYKQYVcvJoM6I0xZoGmRxODr5ILIqPHfHlCf
GtoGf1Vg/B5bQqp0M4SOf/RBkALrntUM+tHj0d6cZIxzN0ZLN82juZ6VDxA4tgvV1Ptx+cWlJ0wW
Ki/iu1432kuTpEpBfEz56WfIZWAudH4hfKf7P5s0MzzIy1EaoBW3Tqv1n/9eVTfvvc2qNvwM8Otm
TLqMCZFa+VQmVYFcwkYT1HC/JpZLvCTjGd6u0YzfFrwMtFV522B9stMTeI62zZ9Ay35SxgLrcBcu
0nJ8eIAKMAOvLqkSWcIQ8gmTf3tyE7tzlpQWkKMUfgO/HKP8UEBTaLnw+sTEB/wEgWeUpGGqNlMA
j/Rmm6no/iqMes0bygLQzRMmpYLNdN0ltuT7Tjzr1/OGihk36Zo7TOy86byUwW/sJIopLGPvb085
4272s8gqbCsJ/NC9XeUt25TAM4zOV4+qZXgtBXELErW5rgDISLy9hoFF/goryVBlXKZ3XhMutLV4
s3iFq6cHMDbk31kkS0DkUAaUruJQ5a7iM9BZiWbJ+6dmzN3r5+HKjyL2l57Xxb9RsGLM1HKv718R
SIMQ6przvyXcoaYWU482pJJ1FL32ug3DHo/i8jn33Nv3ZJqhTPDc5hrL7U8vOSVuMN1yH3KCVrzJ
ETMLzLATiegfWSAI+QIhARkFZhadMNY8oxmNCjQjHlo4bhWPqvajrEAQWnb3/Y92ODHlLTuPF5Ye
egvOlQXXxa3HJL4cS1vlzaSHEzoXdtCbVHjNhqgNsXsm/b9jhkw1GtsbcmwqFybov+HipN/8+U6i
ldJZBnzx7ES3nn/6HNMQRtrRmHf6cV9O85gH0xW73iGZS05vOJs/4kF46F0ORUfLLbvnpKpAwm5Y
yz2OeEQmQnN/NeJqY2+GbjVMC3plkDWWcJCSb6r91kSveQw4WcenE6iSWpxPnn/E8E28UcGJPO0G
HSdaaDR1Yr3gBrp4vso/7rWHD+vGfJmki1mdch35b7+79Wlk9YBArUkK3tbe6ZwaABHXvBsi4h9i
CJn6A9c8cSr/+kV+g+mHt3pyZYWB4KrtWLvCiZjXG+GX7SSOxLJPZ3o+OdBrSGNfdoPq4IJRJZMv
u9Y0eeULGs/IBEp6lHZBIba+YUJkTBEUyf6tRreoCKuIZQlomtKgcmRIwf90LzAKNt8oJMjqn/Of
ec+emDbLAzlgSzymfnHfPxJrhhEU+dyxdlz8aMB2igh1+nER3tR9Z9aKOAiS1nzPfNYsS/u5/r99
xxM+TIsOmncoxi9Kbrs7oXrimbZNpzphkbMLCQmprzijK24feYtUXxkSWnlikdrSfNVjEpcAQUF2
bIXffN71zLsyE8mL7kbBdrjSHCqwtSb9laFEGW9k5HntDg0tXkxybvMzmjIxy6UqwokcERLvLP9I
My2sStdRt9TvtBJbszajXz5LTNzSVMZj6frMw71uaevZMr1QpcD3sfeiNjelZDn0ZAdnNPfy1Rjd
3MxH5pEyXD77bcI7Bwdf2EXtQD/VL+jPROf+gZPWxruRGjRNf3H52M7g6JNsXc0MUfLQdllbduYy
BoDGo1e+KPfR8pZ4VljskA/Krb7JijeeekyEIgk7QD9Yjdy3ezIy9ij0WTsWuVgOBhkRAS8zEW4L
QZ8N+Mmw3cKP2NE2fdbuvIyRv8YRYpQRVtuXhwIKdRBe6BpNP9ZCp7HeuNzWERYGkuTLtJOnTw8C
s4jAqZeWkBM43tq0V0yupAOQHayIZfSA/W9bMuc03sjtAlIcAICRg1J3jLvTZ/GpwUU+SOFdtMm2
2csM6xAp6VFSQLh8XjXTX3/fK3xUocbB3aGbL0J7sg4ndlGtpPTSS4tn1VQCh6Nc1d8T18+FoB3Q
UHP2InLmZzwX75+t+FWlXyWCDIK6mndGYLt4oUs9NgklAOifjss+7/XMfYHwtz7dKSBIOEX30e1S
7XJZtWZPf3IY7UGd4XLBRsS4iwTO8FM3GT/x1Xcf7qkrxDdsW+zWkeWJUwDdMnNQkfEJYoY4KqfN
a2TPCn9PKvz8+XsR4mLkEcTS9ip+t04/UcAG+d8CL3dMNdCX24OmCdwk8i3Dbb2pQgAfYCgedmc1
79tbRBp00hD8waD1WWIQ6D4j7/vTN1OIjH3BkBbFsePKGPZpZ+X+BQBRSpW/NKiALYhrI4sIz1cr
6msGviVoA041o0fwNieT+HO6/+PyuASez9xoVpY1TpFbcS+k6M8BbMOCqjd/4Nx9hUuf5GomfPM5
kuV3qc98E7BaK+CnUKuo7mp4h60mB6agOBC1B05QwF1xqmKist9tJGpDvnB4oywAmzDQClkzbOY6
azoqe4i/UxuyeaC6ogsgneosKQ+vmAbJXjgj6PkL8pwOQc+KGojkjJemtFjTX+1Zv0R8d8+lHI/r
fWZ5ov7fZIt5Ejv9jcZxunkxwZAkyqgqceVR10P3LKKK2LSZulpi5W0fFDtUP+XgD8iuxS6AdeZn
1hP/QmdSK6a6LL4rgU1o9C5h64WMznI77t5FHtMj7UsJeSaN9txtIoZ3GlP8eyeoS5TwCzGci6fo
BVK1/VnjZGu4vJyuaI4ISTYCD4wDffQBmwoCzuN9E62+LeWaizXjelBpShxWXBbc0R+eXaohvlM3
H4gJ38d78MIQFSK4VuPGL9SEvYFgk0AX5BSRFXj19z+G/Ef8kzxy6jTVx3e1WXb4TqeUJDoOIGpG
/saVu0HUibZM/4NCq8viFnteir/3QhtuYr9bt3oXdgCTF6Ewgapx+BCEmJBwS23Jk4HILQdMDc7M
S3A2KbKrtg4+pLIfMPox9/mWcyK8YzE8gLWQDx2H2KOSMb7GRKwuIWe2NdGTDUJahvG4TJi+VgHq
JnvnCnXh2EHkHnkn9LRlb0s2XOR9umhG6TmZgZfyjy1xMplQTBQN4n9ynpEpzspr7M5gak8BC2kl
exrk2aaepSY1NaStffcWmDzLZZuklo9cQ3uU5oUADId3fdVYHkt0il53oC9KY9Qn/lxVc8FfPBlJ
RolwdO7uf608OpW2gpTJYE8KmyY8QLSEr14lUwj8oPsJNxhOzzpN5EtHSbKFRQHLcxHBh/V/HUO5
guT5zxNCNs7W09pxxT6psL/ZHnMiYkHAIHK7+V0Ki/0E+hbvZZE5ZqA6djj47hCwkBvydPusrV4D
x0F8kQ1jXQeLJ848vEtjafiMcYa3QVbkbwo/vMEPf8bPMXWmuDEfEyL50rYbIb0FjNpV4emgNdhS
ed17kM/B4zrRhz7hdFKoeyJRucopRa7w7mB70u5X22T23Z2iucS9wIT7orE6ecSpfAbUJ2Z1NONK
K9URtOpkp2CTk9QrWIhppM89G5vl+sSzgisN1sHbFgfICvf+SdVVxFFzzDEq6H7oyWyVRYoHGQUw
5IN6CCfbBcnhmZxiqjKBjIGIq55iYbuLp3zSS+lNdL18IESj63d+jPNUsf10AaMvTpKy4yG4OAlL
nipJvqNHuA/nCFFuveQga+XJSwob2mjkLbNUhmiJIDKD9rn2qr6eDpC9wHkMvI8fv02g4ZShqxmt
41plbIhwfFlBYUFiNUxcrEacq0s4dWJZxuOCTGtSr2TfR5QskFnNb5Fzjq/rlz4XmjioM6V9560P
avVVuEcF+Qc9jjI+Uc4VB94Ac9dxCe10QKxJjcYpJQNtKJNY+7fuY8GpkxSRhl0YYSIYHp9V3Lme
Yzvz01qnkYfO6/T1+AHWUopR/rBVA0cu2kXfFGELrzTSPCTa5XR/HWBpOIYUQ5IAUhgkJRTzDRfO
k3RGfyRlLV5mTiIaVw0NX6EIgdW8cbcajbG1lXe0+qAZGbEMpTBlit6udD1z8/zON5yB63i08rSP
4AZakusOUlXMK3nYjNi0tuuFmut5OFjDAN0+RH6AxUD5FcCkR2ijR3aXFFTsyzeYe6amUhEuvxT8
WIGurj8JcJ+hyNUXElofpEIwfeqkI6Jd7zn0YxZ0OtMie9WCsM0T8Hb/JLsc6XBiaixOjkMQ7Qf5
FqOiMp+cAUNBAbVniTsRgZajEoFAbENY6G4XyhjJgBTpT/ug9U6sWU/juAaBmeWD7PmS+fvG4jyE
sCfOZ1B3SByhE3fQQ+/R+L/IYyng0PRvb6Z2tybiWFBXqsso7kzxKKBwdaUb/xlUw3s52wh+g9cE
//dgdlmWM93eD0PBtpODAFUBBwuA8ys1ht+2w/bBjqDrjqLCnNyI1UhxUukjdr14pItFVRuZjqvo
lo35X1aZTGgOxLRABwbBLH9D/1C4ntJv4XQ12rVebNaoVqHL/SWTHFH2UJu/IgthI0ewA1Vwt+nc
uMnyS8uuNtwYEXaTKFwwDFxn4LC2lprAMQrOX13Ds49hK+VYymrm7e76pT0gQAXr19lZIpa06z57
Z/WSLwPRnIvZBDe16uBcw/6pHR0zs5I8tnrerb2JTR1KSR6MuvItcZO8OSs1iE2PVylY94PPUxcy
ozs5UksB4baAhTLUka9xo0A6O66BPevB2ec78kUgff4SnFp3ujCOFx6iQyPZ/0oAmUzI9BOaVoen
3z/jSz9SUTUBAkjyI/BDs3u93PC5s5We1Cp3vtVoEDUFWH6TyFumx+IguuCMxNw6pEL2Zf+8JFJW
oemgjGgNcweXWO8V+X7Go8uoCfifl6fZJMbPS9JTBv/E3tCXJtiEGSaGT2c65O+N9OF1ZC4YzgmK
yHAJeukZygVc888BGU1wRnVfo0vtBds7lxMzj7pVhHBwwD5X+aVOjTrwBjoU3NvSJq6UimgmMOfi
fladcLcmMejEZPhVwFe6BNzYvswWjR125JvNuT5dLvUKdW9FfmR+jERY4YzQsImll81UHZlNvTrn
uo/+I30jkqXmLwHz6LINuur6QUVeRcmQ0OaG9GjgzcZsmXGLsM6DF6UoQpZc3uNs0Gl3VVy8+SGK
EMv1ufnDGKtsXx8nFpYwnsUmt3fn+ZV2MH36cCe98iHjXuhNDqvbjELM1gqGPiEEMuJwe6yN4llD
lw7eVKfKXjgqkEjeVLmFb5FwqzbL9/ntiiqQFxwnO/qU0pNDF97s1lRpWjQNBipWHDiXpB0TQAdp
H5jnFotnfwThv2qR0a9b4KD0nt7Mc8yrqzgIQjfYZx4K2Ci8BHCECZJc7d9y6qlK7k6awpBD1502
VtVlBQJhCun1juLWIp2weEc0FLrAV+2hRB8juniSORrJXanempuDYsrX6WQ6IgZO5Zj+BnJ4Oyv/
KduZsuoKjE0qn8dxlOb0u0X3tezehGqrDjX91qHFaTvKOF3ZdbCAC/q/YdG0BVBTOsGdoQQ42dGa
bzlk+GKbL+5mFXblRdKt7m9Uk8QeWwfX5CVYdpRtQP5/Lv+C6OVrspLukGpzNf4BsHRrJ50mt1/b
rPPt0B4or3a8VRsy8KXXgDDuHjaCm+eikj3pyVrHoGQDIzMRtnWBcwCWeZRQjm4tNeptXki5NtF/
d2hTO4hvueienlCRjCGfR0MJcu+CgrCIhYuZ8tUxG6iY9mzgWUQqsGNkh1OO4+iKFq2FZ8RhN7Uq
Y4N2aOunDp/2ZtjCsIkROB5T4ljR34v0doBz4xCxer4nP/68wYLH7/GlvTiib1HYYvKCe6QkghAL
/rgYCP0wEqEd3yMYhibK46H6kxvcXT/gDu1pjYig5XPmqotHsdoZhyaaOwtgBD4sgvr9amjMENOJ
S1BscBtPQ05UFm4k2PX/U2nkOAArx4r3tNiJ665Y7fckGzmwjDKbnj56ak81b3sKwyqeRnul07Jp
lS5Y9W8QGCFGb/s8NEZ4tg2KP9ga8P7+DLDftQ6HragBamaxZSoXnhhK4nEII4AWlNm+F1J9OS/s
c6hla8doZ3nhnNmLkbvG2h8mQ0S/xgaI0I/8+Rx9UZXU/aACDZv4kf6/cxBbxsl6sUbRVZkUNnyf
RBKrHrstBe0N0Y4Z+GMaSJs0tbDcobt99oSToSxmSLm9s6Im1XUICOScZkhNkSwowYWQDjEyynPE
uGTZKSshvMWs3ijJIOtDld20Pe0vGFLOOfKAATshgRkprPPKsnrZxGqH3wnsj3wIa++Y5kzeVrHH
9YjXMIVTk4d2G1qVOWTn4RJhA9ZsUS5Es1sUamEmhpGXnBBCcX/pC3wvRlkECkMx8IKZ8d9YY88P
Uu3UTRcaZmo/dfFfahsP6CbJtaIT1ky+Qcfi6YmJgKXoT4rJXrL4AJhJ1NO77wFlzuw6+SWlloCU
ukxJpN7jpDDcDdyIFOr7/eV44NR/1AIRdSllpfpJdWJELy8lz2Y9LZM89RSsfbLdyFNRjcPA2VyX
Mv+IkrXnZP+gBP9CjtBi1Jfa4kNGwDcKJgT8moIyUmHoNxHoz7o2Rw81FiBoW7l2CcdW2jwWA4bf
EM6AaFzEdED20A6KAnNcds+2WaVwciqYEMY+ntLDilm2V50io47dT3QdZM1xndTocN6UpfZUIK0q
aKUOYES3raqyJO54/eD/qw9vOdJRpL91ltsy5LDO3fXRkHrD2ex0At5dzVTt2qOIRepkWK0hP7/V
0vp3727i7Y0ZQZh7vQKwaNm0ZNdS2609r9tP7Nk32A08+UNqKcaKzx/nfGBhPLICNNXTtfxDnSSX
asv0/LSEOD9l25ylXWBFW2TPf5F4xKqpz66+F+7GCd5bWeO3yYz8ZgTGyegqqBTr8h3iOtfhAJif
Wi3SaHPh9vSI6iJ+rsmS6223by8LDX/5fZRaXGS/TqseaHA43K+2rr5Fq+NNt5DEFx1LJciNyPwl
P0amKXZJpnnDKCu0g/qK8NWQHmhFFSV4IVUzYUoDgejTfqy0H+OVYESSyEOtCVs6MPJYNdU2TGld
JJ+q1dFJfx8oc8PB+qBedyaIWKx3mYg3KLBkyOmbXKq9ftBGUyLZqmWl7NjkZHCp8K9vuAa5nQKH
E1Cc1rFi6z60wN7b5Gl52dEp7fwosHwgCDBPVh2HMFR1sd+M+YdZ9RwYSUMeXNhAL0JYfSOnWL00
YBrW+yX+WOH85Fq2bxTcGQCQQtKI8EhVA2dXypXKoxLpN+bcnIpVy65qqw99ITByxfWavWM2SkQ5
YtmwlespCKLIMnVEpasFyDmJ1zx6CaVhzs78SfcRrpfLgnaD73x4iQV5Mbps/ZB8ONTu6CnTs6WY
etY1/FKiujlWxLettsV/Qzw5miXBMkZPJtws2HqcuNfhfUARUZhtrHsX0492eLkq+Prda0dA3UlI
mbLuccwZ6/eC+YQZ3zQ+AdVqw8me3+4ZtTb458PmlLFj5xxskf9ejy7okfLO7sc4Dp2wvAVrWtXd
dk4bhThv6C06A5EzO2243gg0TeY3FF0hAeRZjHjoW21Jh/Pej4D6Sh2GuOtcQRyvnEPB0lRLsvB8
aU/ttjUgagwraLTgth2OUQ5NAXTU3vE6NGZShng8saL2EuYdLugqnDXzqwInAqqwPaAlvezEPfwp
T5QZs9VGbScyTXYO8cU4XHJSTS+F03+FG8YoxqnoQ3ggCH1c0fw4jDkEq2MRBpOT47+j+/s7YSpO
NTZ4qrCUO8l07m+EBS/BEZiJCEpPlWv7aP66JUL1MqJ4oO6uP+hxbI9X/KYhEiPObT/A659ps39X
96DxpVW2cLlIUC+GQzn7w7Oyz4FKOZpYHHyFJahld0fx6eUsotc/m+8jGUKLhhbAgX3DyDoAJCAp
UcOk6YaM3EY2XrReHT8KWHSrXAjFXnJmCn1yCCQ5eQuBvfncYzn+fBxQBPhy67dn9drx+luaSSB6
PJ6KtpaB+h5u2xFzGL/e9wRxx1wCrAjFkloDtXIBPCOJwa+/Ti2XyD6ZfjH3UVan5h+ds/ORIwq7
Bh8U0BOS8FOh0lKkc6smoIRTSo9HmZ0j/ByjWhQ4qAGGC2qDFVLdf8+rBbs2+4Uq+SZya2lfJsBr
sE/StGfFKWly8lZZKVnAuHZSA/f5GgVkev/W+3e1Ztm2SfMKt39JsPaJoSXcIFtYNlXm83kMqAPQ
b8USxkuMf+oJMzot/GMj9Abqnl6z/Ln/74Vq03JLrEDfMeapOYuWDTRxZsXuROzUFNYYYLumes94
ICzQXQ4oMKm1tETB75deGKpmUVjhaL4xtYJ2eXsC2HwKGQ5xcXg8XNSkvYSYx54LHl1pBjeAjggL
XMpZTzW0XqahuGAHITYakyDA0woQj+MzBcm3WSQJ4m+L/K/oEhVJhRKOOrrmpjW56JYJ7IxwXPp8
TawFImdqQZxbHaU/7qMOQ2apwbalq1KFICxedfiHg5gE0tpqXlsFofsgJMd/060hzkquu+ZGD7qI
oF4zTDbVpEvGc+yVGNocScQzOiiIQ0hbY2WQXdpOCVouSsRNFKQ+hJRIZu/BqLKst83Y4AK7sNpx
GP0OegR48WhG3UB5nBZyMRGjbEa4F9zVG5waPR6PzAGaE75oxlnv7c3bBNF+gQmbvjINxKLlDI0R
djXMP2CFRwgmK8RVyvCdLRTTZr5UPl1RGFhnuNAgD0T0uqz0cTUn65GZHLKn1LmdvkmiezEt12hY
7M7mGkYKZAMiI2YqJn1Js/Mm/yJJth9NPM2G46hlrpOvxjPCRZdjH7AJpSIMiRojn7qrHE1jlQcm
w3nteoJ+M8j5Mjisr1hburCYJzSnQidKHJFVmDNfqA3ugPrGTk/dKR5oPKscJYGSR+MVQt3JIm31
GvMxkx3oUHCOAco6YsNIgYIpgwLe56/UqiIJqUJ2ghhlXPsQ2oHYvOCqqVpjlB9xPOZjWxl8dzYM
eRDdDMjFY33z1IHGJrI+5A+Tgcb44CitoFGLoTQhSedPR+QOpsZ199xB5x0Y56yMEpBJBH8oujQF
fqww654xZmUtD2HBPjP4s4mZimJtwzJsanBlKxEWHD81m48o6gg4JiTA3n6ce4OHK00hbrq9e9Mz
4zCVl0TAhs3PQCEsARbxexhVU2MneGCqUgWh/gmbE2objMFeqe9ppyUPBKv1widCD0OIIUrWlPOG
HaI0/k3MIfYtKssV0C8f/OYKAviTj03g9UXC3RDxggj3areSGSBNjgqQI5Ys4DIIshgKy69kJHGs
5FviWazWKuMYW2mRWsedxmioELYBHgwWnArTyVoP+6dBHM2cw3o/JLtAoP4z4pgILLwo24AtHXu5
Pq63fiEsr37xqmPWicTNnO3R/EJ1yRgeImqz+GFzt8vBEQ4tBvOwSjuXceNm9BJBUcM0ea1axCSV
jIDKKvFN9Oa5N4n88/htEskbPopelX3F+8wRzis7IQm/CRRURi0Qi3wtnpk7tUdfd0gdrzvdPufF
dO4kF1/hSmRbN6wNE0a8JMNHjNw7nBMZVZr40QbW3jpo9JyxGsksrn0y1n3Ns6wA9iEE4uj1lBu3
NSO5xJLcUcZCO13O2O/MmyGKOw2AllrGBp9zmpbPqbrdq/h8SwA2Ti6oTFSgVnQMpyM+hgnxA4BT
xrzhx8RRzACbP4+oLCIgiOwh8Cwgl5QwRQ4pMy4/JssEB8JL2jJkbRm2ddRDVu3v+G46jSejsG4m
g9F5+nsPAoXzad4JJRy9vL6a2X9deNGtNyWBOeOQMvn1jDFGZitw6vF6OQhw15kBXh5H/q+vofv/
XY7IKFmfKCgt8M1YwBXOf5VxzIU6xziXOmCBVLNHucVPGwYe8y3tLmEAbOytOwXAyMqSmg5F+GCS
pz893KOCLmurdVza9H7jNO8Cc7IJfTmYAVr/9STv+1RoDk6VFkorWErt6EcBfXeQ15JneJ10zBGi
8fJzvUmc8LRdrn2zchMRU2wZlxKRbNJ054CrC3Yn+oYN1Y0EKhhEwFKIqQoIBRHSoAu7Rkp/h/iy
3mJgiDBmNY3ts5U9vR7rac5wyAVQ6+FbbxCfUZIP0AthxcxXd8J2Q4/6wDN1YXmFIXOuBnZOCRzk
w9V85pFydYUly5UKLZhvSqU3WkXsqVr/cYaYRjMFe+q5b0JOkbGx076F6YK7ZUA2IqedjKsWPFdA
mcQMq/1ZZQkYqLBu6lJQJ4r0k6BL1EXY/dwRDlqm/CUMqzbvzqd8hTgcckW55FZ7I7lAc2GabzJS
l3CYL6lAD7NY8wboNkJ9V7ZweUWMEvZXXM3Ws1w6mlxslbMugHBGAozxuW9UpOlOkZjChWvPGJD6
oCtn6EUg9EMQXbrpZvb4csK7bELNg5R7sEQz5py6ue3R1A6wZj3T4wGWQN4hvENUr64AqZx2X2Dv
AMjUBoK6TE163uyCJ+7sw5btaE/TWYhZPBteic/2eqQJBMYwps04/LpgV96SQU/eYx4PqGQ2PtBp
2iNtqqItiKPDpIScED0A0AAA4323EwJVZtN9vNDgLq/6rLpsFX8vkZdJNOzWfQT5G66WIRyWl+Jd
8YU5o5WcN5SbDNr27gu/feDWMKfOqQR1xc0x4kFcZrSOiLgsRGQdbdXRayreIF9I8TiorQ1sVZ3i
vw+smC0MV2pYgE32SWfWwYOTYofx1HWRBLVIIN6jtPlzm8C6mDZhzwWiCJr4YJlHc/KxjvpDpeGL
a0Cmbm3JBWsxaXDOycC5FvPpbL7aZM65smUrXLx2PqTw5lJjb7wFf2XM2bT8hPSUJj0Evpd4escl
0vxg7Zk0xGkMK7G/3G4+Cv7+d4PM1QK946QNPVzV5TyqlaHTi9XJOm2pkuCPaLNZyL69ofhWNQmX
Vp2O0EwQXyrBNGMcYMS46cUKcG50OJiB2aJpsXK5vuGEQeG+9EGDeNm+ws0+05NZCCK8tM/pbVm8
iUD7i4w3nVH2JnWDV8dcv7nID7Eb0JvbDXE6+6qOU5gQ82X0F7LbSWBTd4c1Hnk8s2rUwQbXvPi6
XNqsClQTMf050YpJpAm8ZFUFDzUN2ZFe09V1qaUfAwcguQg4cYJRu0epw94donDzYl6QmYOrJAfn
OI1cTc337C1Hd1zka+s6Nis8Iqxf8xeohxbXqGc58Yim6q5XFYL5MseY7+MreZDrvDx8tvwpvK0G
+yOH8V7c81KU7F3O1fWzsuiJA5YejubWeN9nN37uv6d3xfM61p60K+ZLGxgf3dxvKTiyuPHzCmUA
jPrD5TS3wtsxBRwtCp+Pzez6tCALLki7A3Zcgjc1rbURSWvocfPZT9IPMotT/I1GX4mJjgkNgBPt
D2k3zAeVce8Ayv4sIXDhN0ncZWvfQUoa3CKJCzHlNDL3QMBoo5oBfzzEKArtSRIkp1mMcWAEBcCn
d1Ean0jCkE2E51fBqSDbywAfOX06iMJsPnDgKrB+eXITygS0gyCagVu0doV9AD/ytck1baQwSxcA
18TDHyhmid7QpqY0XyWA5u6AsMlwbowHfD+HFv3pYVqArcya3+F42AESbv+DRM5H8of4URTVfEid
QN8al5UQvEXR0E+l2dEXdgSkiFhk3QLKJzLPGsuLCnhb0R4dlpPUHTGRfDi//Kv+VlJm1TWgKndI
CH082WUklD2W8S+ZLXg6LG/jQaONlVEfxhNaA4xqZlAb6WEhs1Pz67noPGMiODJBw9BynBD03rre
PxohUzt2p/9F3Zb8QKmZeWAQpYugM+6EMVm3z2WDzwyS6pHcUNzAWcAFyo1bGMZvKVejEm6/CRte
8EpFLU9NhAHSqioYllBmbYCjv9kgZtUdG+87R0xpf5RvwJoa9bG10vuzly/tV9BL2gPInFGcqBTU
XM01irpB98NZUTB6/UOaCrIvrJeyR/e2uc9CgibJpIJ+Btqo6pgUcyxx5sAmtZ36EmMn5rKgGQY6
ErlJ67qKldxche9jmklTuns8O7WwcXR09f2b+LOaf8RX17ooRFlsAec8FpYFI2cFyrZ4fOop3zCY
/mmXDWGB3fZjdLxjl8iojq7uLPc5vPKfC2dDMQazqYl2qmDwFox1zim/gyf7H+nin2VzHyFeYh47
R3cfnHfVTE959mzjhh3I3Q8OpMjjCaLw7NRPFwIEp+BjvCKYT+dOYrEXY4/RCcz4tVPx96rTfi5Q
verkVZDi88WLa/DVXv7a1MP8/X7KjQANkc8cobtvzDy5B3/2qjemlnMSnhDFxKfmJRm7bdxz5QAc
/3K/T2sO6o4JX69GL6v332ZJ4V+Gddx3xEGPvatk5Zj90wGijdTkk/TG2um1/wenN5bG97BDxrv7
C7MUrb5J4VctjmkD8vrED436koCN9x+Ol7GN9okE7NxawkNEus3L3jLhB8jJ6xOX3nRGhp5JABmJ
/QQSs2hVLDpZwdlb6nMrafJxJ4+2WFwNQLqmBmsya4qkRaFOWbMhpz6aRJNW1qpnJrlRijWz0kxg
Plb5s+wLBoTm5RMoN3WFrAw86vDiJYnoP0Y782kTnd9swncNLPxYcEbMDQqx/Q7c2N4tU6K0e166
O2IAJn+DDrPNfWV4UuwtOqgHxoSwwOnVil+YIHoY6Vj8/U3tqLVIIqsrt0ols1YdyW5cEGfqqEr7
RzEtbSdSLDvA4fLtukQwc8SGy5U/oeZBShmvVPxpsfPNUHLuRH7wJiOTPxva1RbQgq2XsZIBpban
nHEQnJNywk0ZRrnkOPux0Vc7WcMnrB9RV6WpiI7fstx6fp5m3YsUH53d+MDYBfbBHztEuCr/b4xt
AXh8F5jN9z1181dRSD1vWtG1Li7ls5WCbBOcld3qT5YwC0pq1j2ESQtz4H7f38nicf0B3xYZ7OVr
wiDG2LqeV5oO2HGpaoiJxwcQfqgWz1S5uR+KPoV5WFC1tbdJggbuQcdW532ft2Va3tW/+K4KuQzM
rDnBCAvc6wZ8NCpdNymSu8UQ0nuYRLas/IBhS4IpRNYbmHq8JQsSKFbTd0QJ5UkC97fwCbjufE5H
1+02CObSLfUEWj4X0TdvD0nTs7988NMdH8IcyhHs+DOgjnlL4SzeKBf4LhIjePAXh4Wvd7hnyFpy
R8LvW6IPE6cp/OBmSE8zKIFDhkuDAdHBRV28o59mMuDRh7mtwJ/ACCoDabhcZv3KOcJUbXSUERT1
nMmJmoA1n/reM336qmZrqenSaF9WSwLo1yJS3G80ncRR24C4YZN/97gqUsa/q4FHqLSprmTMaP+t
fDPAOMlnC7f+BIcsS+cinsz1ZfUWXqrk9r2IHGu6ZJgSTTZzhYGxLkF3cLGKYRa5TFAuP7h1gunJ
HT8lGV6fBfLJ72ZTy+oGhJDGzXCuVgvVWO509UxFMp4KcvfgWpK8pBn/Zlzeiw6PtLutw1sG6d+f
GmQG2AdoQg8cOiCVB7IVh0ReTT2dmIo3dIdNng1ED432FQJeJs2r8GRJTl5k6JWUT62blNxRbYUE
hnoPn3byf4NnQeFIf6r7k4JuSFnJFiyh3MiyiE5NQ9d1mRuu2n60kPpoSFE+Q4i88XXAa4U1XR6Z
ipxtUUGFxZpZaBTBu5bXyS3LG8xKYn0Oysp3yI5c4jV/OSMsJLxWhX8KAKRuDS1JAekXThty/NkG
yMg3lGsc5tC4+iuvQA3BwxaMUkf8JDfhP9/dzPpyC5eyH9rbIsl7y8fzO33rs6otix3ue2q510HE
3+TOKlK5o/cwl7VcDHmtCd/wz7UNMATLQPi+maovZCNOcuvsskxUT6SUPqa585KzxyKgvVw4w/fB
FEHrhSJ5x0cVb8rinjxZBC0Ub1ClII8xP5r6mzrm6LwEGm5mPa9GODcIfnMFU4OKX6ynPa2WfiaI
OmPfpVep9Ox+Hjz1I6UEPXzTEHM9h6ZDABanPv/U04CyaKRrDMbHoD3TJjm5Boo6RTiMuD25U7Tn
nYlGPMKPaRboY3rQK6zmRv+BuUbzquOQcaD1n/KxtZBNoa4hOcSULW0I/WXu0UqRB5Dzqeqg/Kax
3JwUlEHj8d5o6hJoxuAhV5Lfy3TWWPvgdyI0VGSVwchJLAB8B13DUaFk6tU+MJrOMAGrHiYYlOmr
L9l34MHUN1JIrbqCXHEwB+9+GGTcwoDeibv8lYIJ2yurdMULk5VNJfdiCXXE5W8TaJ94iEiocquM
ZHCiAaSiXKUmENqxAm+uTUJjBkwhzU+RAeP4nkHq9cYx1GHbpYU0dR9edIkCVYd84X35UMZqRn4S
aJdzWEbwVgSNHlNynUPujRrsongab6cs6c9orC7ULdS5lAvEserpt8JrcoYU52xQs6/oV8AGuN4C
LmsFWG7f5Akhlxn9IEd0px8gmQ83AXB4bHKUQzfXoR0W8Y25tKKJ8k60Eb+d/mkj77yyxsT3zqOc
R9YvG8/0Ea+aFbekXhrctkwPscK0vPUOY/4K5Ml0R8VWMpPCH193ZwPwKcW722KF85IVXa/s/VjC
VQkdbzphT+Mfmcaz6JC2xEpgql9nVf4jAK8DealMKQUF+sEKzvrVh2FoliiEb9CPs+4NHkqAesLs
sdXnlqJKQHQR/0QNk4O6a2Z1Eko7RYIUYMVTCz0kV24CzZPehNcDG1Yp+NFJ7igI27qg7qfhS56l
/pq90WqzUS40e7U/N/ydg9CciKqJr0p9GerxXw201a4BNt3zP34aOQmRZenofUx/sI5cDr4nwvtB
F6+1zMxEDO41W0lYRTgEjF8B47GF544U2lC5YK8aaZpjmuXgbiU/9S161y74ODItprbhIzdwDc2C
BumBdcdoLyfbb5dxuKahcFjQECZXGmWVM3TCOfylRvMOV/qM/6HpvCz1wyiBw+PZy5vDxwI7Cjm3
cyRpA9tS06W5Xou7weil52kI8KephQRhNZrC6DZjzuV3gYrGjrdhlmhjxNEyjLlbU9prg6ZCiDb7
jpcD22cBshnV2E27p5SU/HBvCLyHvGBdFkoEBfBkrgLZXzvppINQt0rIufjqxYnfeGgH+p/Y/A4p
NnVnNNNRP79ElprBCarF7y9yXObhAOWtqWnLSlZRmle7f5NM8+Ec4uIunRCTvkTswAvIRVJxjoeQ
ygulSrJx/m3AyMSaU+yEKgXTbghkikr0VHzHKuuEDM9IpGZ6yF8GmadHnba5qZQ6cgy1b5RMBIw4
cELFfYe09p0xhLyenbBJjC8IRSvozO9tLph2Qsdpg2QEQB+HsY7YwzXxu+7FN4mRwp/dxeNULPcs
Ec0n3NhpcGpLaLD+DB753zrlD7El+722DnHC5RLfOp//z/E90xNqVt/d/QeqlslpMEdUsrY9nF1G
k+Q3jEkqMaO12499w0/InUWcacKPzFMOEuyBfNXIIJKL8FdcLJ6Wxb+Q8s6RnjKKCJZc49H+RHZE
9tUXrFYBpT7Pi8SpYNoqw5GS55HNORbYrX3sx/sVMtZOOvi3f8dI5lKhiI93XsxsSQ5IgipmdBKY
sJKtq4c+VL5bbmJnnPS2VTw3EWLmDozmg+1rF1HRAozL+wV8NQhuGDVWpgTpPXrenJMshIvEZU1i
3w1Pd0zQynwkGqYX2wffwNvkt7KO25UdXHLOeEUkfIH4/1LNeq+zF32DrfHscGnyE8O4o8U5DV8i
tMX5yiSxSMhTqN/eCsep8xPuU0VBjNapZI8bY/0xxhVHq4rpjDD6MGL1BksZA1NmUxEXpQsVMAZz
Gt9g7MJmWoppDdyiWO4q3UF82/5vX2bDyOp0G4SUpdEdb7jb6O5OW8p7tXIDtiHeSXeyImRtR6cy
4xALLEbHvj/IZ6gQjEXV2jRV6Fx5/UgFIwFbAVpsrYs2mL6odGdxSWmEOR1yhB/b/JKsHdw9v9Zg
O0y+7/C5K3ts7DPzTeUFw0pP+GKY7pbEHSJITVKhpGNAdZVI8a7yL+fccyyEJX/DfRVpaqD7x2un
IT5PBmxkJt5qYslPcPgHGxE+QqLbqsAWhT99Odkr3PoOEb8KHKRGXWR6u4lNaKBWxQvbo+2uFDQj
WBTvzyfMLktMVU7BDl9NLA60XiQjp6m1y1/qTXTc19v+ieYCLZdFh3EYnZqel9H1UO3u5hUiY+ll
BIJTJmUCW5zMffnBkSJReuv4c4pF8t/866YxYdjW1ZQGsz3fV7jDvY8S2ef3B3+vQrsRMNQyJWIQ
+1KdRdi3+aXRJtg2YI/9++b3Qf10HJI1P9B8sUOiNimxFBr7VH77popdwSRHUXa4wTAcpsKP2ybN
d/ky3Bsr86RSvgQab8DncGePRHkS+2BzIAdZca3Ukc7+TAHqG5yH/xWWBDCnW18su9N1Oh+l3wEr
oDXs0luX6Z4655xCKMBdNHSZ9Y2smsPasCJrfJHpuSusumg+FBkrJAKBWCPQpBgRY+2n3h5m2bL2
Oq9TllUjWShuQMmpq/GEOjigtvWagFcrfNkygi6KtD5QGbPvogVV17bLPBz7duhoAGtOwKc1NBs9
hZcwChDdvPFpVSl9H+C+jrzAJAdPh7lyKPf22k8gamDiALUdEH4m61fYR1us7MLZd/3gL5IUX8gQ
iVp++Y6CYjZoWeEokzCLXYRQC3aWbZph4Yv/av88TB6D1dwxn3FzOHdzGAKRQQuzrD9jiENlkH/A
ZH/0GFiT4+K1s3myONtukMnSqOIPpVttQ/i+ZMsruJiRcgpkwubT/TCStU+Q3Nzaft10vv9ClZss
4OHm6MY7er7KSyAtJ20lxwQKGAIrCDDy70LAnkrVCrRkTVGeFvNtFHKbkmkRe13Rgd7yKnxGcpcE
VIZckXdYdcZI8uwWDT5fVBe4Eg3ak8K2s2olEIFzfFOtHUIoukfOWyYQ9Z9z0hZ18zxNHJzw7RH1
qSNnNkZBO6/T7xoa7UXUdWDqp+A8hOoOo9j3jZiUQEHxRxzZNwV4xBRpZfi4pYAuPt+E9j+Fw+KS
xGwsEIY19HnEqxJKLGFnfnJXnk9I9BkQQNw6qLMO65I/97ppDvpE/OBYBBUmtcuZft7XIVCuLUgu
7c8tGLXOCyI33NeMMhH4rXNcZnMPPUdbc3qq0GUsevVXyNp4yzcv/5BiboBr+TqEo/sOCyqQhBUA
qUoQINwDiHKEGlgw7AzR9H37kMit69Nx9PkgJWhsLHFQ4cqXziNMA17rFaBhK9y5yfxLJ0IIZxg2
l4JsL63EQaotv1F+ryQTWvJr9kjz8H9Ke5ZmP4tR029UAHKzPha38jCZV37MEgoiGc5EITAot6g2
Xj466WvGcEbHUKSFXc6ObGql2UMCn0sz6FzBcptqJfTrCx7KaMNIP2CgsTj+ZUfPwtji0ZXjtG4w
8avFCkncj9ca6Mn64NnG416ZCVv7O8CbnJUbl8IPnOj+/KRQ98AAWTg0gUjsezgURBU0ymtm+PCh
Vh53kvygDUrvOqnx8DkItyxwlZ2aAUHxC4B8Pi1E5XQgqY0bHmaHnLhMt0npiClUyRGL6XdvRm93
H6fQkJNOfFDsAEPXECpXfPQFGahBARfJuWYG2xOrqiK2Avng+7qqHzWuU4WxeNOo62BiPUXqH+bT
dMJQhzeeFlbYtwas3KFdAY9IU8vG2PFtjpawIqY4YGLJUOta9kkOFr4Mgj3rnIIFlgWOeex67Gri
YP5DFswYpRU7izMD7SqqAqPfk48Os7IsLMqN0oN0r5v9AHrr5oMTpAt/2F339VbD+V7/Gq+T7bi8
bDGpjN5jo6WrJKfyiy8qWCx3DYZ0ig8eYcnEJgDOuxyo4qIGULcHK/3joYRzd8kx0FXFRSml40e/
GMVA7GZbbjwkmmptpGyhlN5VsFkeWyZ3FAsfvMbPN+hLvxs3n6qNvy+xrBMN+pH/eIgVcYExui0F
BfyDakM2sBNusVAhbdTWc4vnjkQjgx1j4q5AO0nXXFK+RDPHw9mu7xFVK261NakZiiOeC4DPiBd6
+rW/bkVJ+fbnKuMQ97fDJu+QDJzZjvnigMDtobZ7PQl6h1tXxFz60B8/e1GoVoGJDQebtBVSmn+f
MtcnzYCbqIevZ/UDno/JxyXtPdIw+W2y8/s299F304cdA7O/OOBgP9PhuYUXsuFOKhXIp17W9Kqr
wCtH3/CiwYCutF9h+TfgBqWpBEFZpMPuVej7Z9L8e5e92VaN4vY5ZWO9qCZHWBxhVFgaXeVEVkZS
HI1aU9F2rMj8zaZesJnERCiDR37FiXdBFzF7ZjqZvPUTgT37ywtE4F+Jpdam9Jl9JVBvwQP6/yIA
yQuHhalrKSgCwdad8yG+OWumlkths/nUNo1hRosc4g8fvNtPdHPoKbnln3fnfkt/9RUzNmf9waQk
v/SKsXNJUrlrxhN0hZp1/McTwthyFcZ2p3EcuHeW1NhEsOSyt9ojubRA5CazCXFX7HgRhYZ5NJsF
OlSxoR24IFBUY348HmBj3t2EcuOfKJ+IZfLM7kFSyg3zsSAMqxzUAUhL/IRufBbuGV9FLnBhMDC3
1wf/NHdM1JKnatNfkIpKqAwRKZkevbfOp4MkMd4TSZ7ys+9VLHqgTHSmKnoPz4z4zeZ1IttkHKaE
rIlxNRER+GzSfa9J9LphUMf8RQEsV+NTvoaU0uZdwm1h4q8v6iqxF3ODWlwVOnis2YPCA3Xbienc
TvlrbkqFYBkdP1/X9+XT1NTOC2JkpJ3atUD4D5qVF8h7azluxa3CPW3ZmLS2iQ0w/EtR8lCdIYEp
1GjdT5k42g7RGbtrwTmxCdr0cfirF6m8doer2phxWiVXUlUuqPSyZpvpQENifMLxlHYYz5PKksJ0
AaKtd8nA35OLj2ZFu/i+14jnoShnIce+tdEZA+Dzwo0Bdo8n/LZc69128jtoZdux7p00Hf/2o3xU
sB/WMqdZoBmhBzOHCICm9jyXBFNsMkyCpE0e8M41PEpvWFEXUnTv12EzISPrOlvcDvlIyAZ9wQw8
t6JhB7wD+KeQKhpsu7ZAZTMgV11mCD9ReRT6D3Z6+U/TgFROp0xmIyK9cOthVNfbI48no8m93bRS
MJlkb6R9isiRDH2u/9w703+8hl2Q4QqglCSI/FAFzjfu0QnJWXRmoO1rNeoWlpk8jBlwzxlCunMw
22MSOrNg5m1GaxQhfvGG8P5zGbm3ZDQucwk9H+OL1cKR/or9XcRol6MVmPB9GCCsMzpW8ssC6oEz
bDRXza5XGKCLfKhh738VFavLkT2/D7fDqyM04Ss+4L5UIvJOS3p5tdZ450QZdt6ZzOOXSqCnfD1U
uSCHnT0dfRySxDwMyuuzEnvfaEbMODdLp7Lx5gAXfVXc59id8NChxgrerRoU3r3N4qIxPPejwZLo
HJbyFI08cSTobl7kQGhj1E2yg0Ad89IIrGqz7c5bcRHB2grs/WzbIKDFnlC0riMFQ7JvXLRgrhwc
EOZ3SQlQrCsK/G+ZoU68a92RR0Aik1Zg54XQ7p2nc1egI2526K4RG+k86Yr/CHjm/GBvE14Y6/8A
Fp84XXCeWgDNDrYBg4vP3sAHk+eUxbz6rBNafcFfXiiolhDxDOkaWF50AXuP+6Jcrzj9KA1BhlEC
J+nCSa0ExzcNxzPBoNPPlwd1IWLlaGB88i3UDV+AhZ3OdM0MgmRe7gtpV67fp3erGmNwuz/do1rG
PmqqFFUvXFOc9QsH0neduqhZFg0vihXDBG9CW1Zx77qTiAkgqLZG6rikYisttXcRwZmpW/vWinug
6pUc0hwBk3MfDndU9kLcNMa/nmdR/LtEzfwLm8+QgDIjykuxcpeI+jxVUv47zT5vulBA/hWoHBIs
wgA2S67NkMHu8QXKU/dBJROSY+jFF02N8r1IhuwQmTHuEnaEdF4IG/O0CDeTedDGw4bHobYfnxOS
i2/g/pkkNxXB+CDG90I1Lme8FnS0BjuvlfQFedya9umLp7F01xAsfpkn+a1iCsMLXmqXmDcF1c+d
+KnRMyY2DwhrkSYpVe828P8I0jH62HiZlKzODaPrbcZH8pKACYeRJqsS/q7Xl8g3SJXUoed0RvdZ
zqix6OiEn1YK9tmGiF3r1Co90SQWsH0TzgvqRyOlgBXeiJyAjBI2WILI304bi1nNPMxFF/3TOf4D
6j7rfOaiDFsgnYYve90ImfmS9y56u7x6pJJW4z35PnZBzSMBjAcC+UdCJTIg4Gan7/q53nwcf3Ba
QUMd48Qa3sYWekCdh9vrXD5JDXfnaUOr6jifXV7hOlrgiJrJGrXHqQvadrqgA500UPQww2Su//dF
wMHLTuUvW7uM+9FoR1aVN4rNfMdpGX1ZO/s8JKMdDrQuw0b3Rw5h1WVcrb3bpzj0LNcHdrRwsz0A
ObzPuWchVYzEdHRy/oYRuFrz8qs5OgkU7C1k/WanaW31kt8ksNOtnNXDDkq7XekgZwFLLXoWHNoK
TbQG3UigC+OJMx6t/KIM0fKgT52lmVwSbCw7T3kq6QdyGpHKvITf/4bl+v/oGvNi+i0mCkSrkKbC
DcVe8/xhzlHMYvYfi6H2+ThZooXClh2gyLCwG24JvTVs02lzWJVZ9InPLxYeAES1RfC0W0BSkcRS
uGn3l+BeZrHuSdrpfRcqcGhXgwH0VAL+mlgIz/uAcApkEFFhEoCBclgU4pNHSlM+LiTDlXMx1HkS
SK3biqvL/R9lCja4RCJLGgpwFDgmKKYA0QDp4vh0OlIdmmz/tD6/Hb8e1C8Dqaz3UY7MjPillSwq
qqlDWrn5tk45I3NsbGJV1E6/cz+MGYLTw1646zaoakPa1sZEFpPbEA0wX+fQLzylgJ3NiK1LGz2K
0djvQUdMKzwKJnMomSoaZIjZwKGbmcZ0TuslGygemSdncDZtQAT9Oq1clc5uKyXa4c6qzMRWBm11
tdyyALYKVctgfn4mNH2TBYVez7ngv7xd8hApFIGEZZPRgqgU3iQlr+dencTbFjF7uPBf4d3zImQO
RNsJnbaZNMFvLgZQ+1Kc5V3KgPAY7q3c13UhBy2HnrQvPSew9g3T4bkM60zjS7gVrpZXbKeTq9A/
ZXwoZZAhx/IzdqiikERqTjGt/j2qYvDSM6qhtPelSppdXv/bn0tw64T+oSiCqHPWFPWfqXcI2kHD
lvnx2cP0F1hPfKA3XxXjJYq8jrituoS2nfbZnelYy4/FnqocBWAI8GHVfXZl3tw1RMJXBkkSVHcV
GzagxlM3RYoi3ucWvwk/IQ9iUuaVwl6kESquARu2/L2z8stGaiiOsRQidWJob1uqvp7VwItojk6t
3adpqx4k+DawsEjAy2BJVgNsF9a/YaH3fVKsu7gJQdvmjoHByMkrl0NqETfBZbwaITfM6+J/i/XI
7qurTC9Mrhuv0XvHwn2C3XRsh08qjAUxI5dItejPuKrlQ4+ZHNp9bo56K/U3uD9vT9Mydc5HRtBi
HHFfQkMKXzr2pMHAnb9DFQabe65K1qhzxfBD4WwpUbjLZIVec2ngun03bVsxBfLzVd1K3elHBRJH
EKimF6k+5L5nU94EwXe1sQgw9sCD+/2ALDtYxRWE1lPJAssB/BSjTI5AnF6B5IJXH2C6U0ykLpwY
Ad+kTOfE4HuQvjQYN2U2RN6w92qH8sit9vlU+S7NEmzplIwji5FZuswwEE1mt9DQcJr9QI9WD7+L
qqGD1GSc9qoUJ2akJjHJzPW0irN2ykBX5MOjUza1r32qtgPMtcPHLnqm7LoBSpzohbWgd78ccaIw
4qlUDkcbvLdSUrpU9Bg5qMjoUptitJEIpNYkC4oVJTDLNBX0slHYyzNApqDFdDh5mOQNrKU/hLIz
Cs3PjyLdPIn5qfOFKYd0lI/wcgJMUvSESGTOZLo2ebwyEEeWNF5YeOfQdH+p0hFojrvqczs5tu0u
hYX7LwMngYT2sAGMgmeZbD+s73fcN9kEpgaiBIpYft0JgXgPGZZWWlUH6UUIzYiza4l76Uy3fJ2U
bSYlI+K2BSDjMATmJWNHdNwcg1zKBFVrbVIcUmsW7p104dbX3h0RBcEV75SoUNP6Q0pHJtBJibhd
3BBsFD2IlxRRTlX7B+veOn4VPAWrc9LxUlXzzVBjS0d/cTSUcvEkuL+/58NTxEjmMMhiN2fX9sUl
nJa49Ngx/J1pWIRwm7zSnOz4fKpYjnD80j8Lv875XlwVf4QnkXqBFySsaBTmCEFBMvHWNcdIGgaw
8cm3o3gyoWIoy/S9QCqNqJyiLmzs9Pmkl1zk/fdfhiwV042r+dgwdaynVpqeqcUqlKevkfmHjUh3
TGfNd4dUMTmjAph1dB9sxkXZ1Wi6yN1RZrQlKNd+wS7FJNhvAlpMbIIUhgIfn8FSdfCEOpapfuI0
WY+xaCpnV3JmDom0B7WgbnilG333PbODBYCdUsnJO749d5NJODQcxNnpiATnbtncn8/0tak0hWBg
ygR4+99vOdxgnwZZz7A9zd+Siav8s5dPYgMBkAbhwL1RHmqWYcNxLiR7UegT0n0Rf00rZ6qbufcM
OTYF7VAI4qWCF3vkYQD2fVp/JhgZrXIU1/8c0uuJGBcaZJqMxyVt/EitWTMPnUKB2TtRNwCoZCop
jbrXqTtczxYaQIgw3xX1vPocp3/8Tc+lNdZ+RKx0ELEK4ZpXbiqMhz2ijaUBhq/KURsIyTylWIBG
1jLocMWAOa/XygTMhstuG+HpHnGlL/HveLR/bC8n8kHXyjBUYAmpsaa4r+nTCJPHIWwAYKaXY3Hz
9iUs8j+yPBxNZhnO1TFz3dT/MU9d9KnOu3r18JN3xnOl5irmx5YzakokN9nIf6gtMMCwO03NvX5y
TI4FZSYPbOAhX2DWnrPsELmi09ml4xMyI2NrYuDxZsitJ61ZbcVCrFbmoiPvAzDdJgdamrKHMKAu
+LAl/queUfj1LfqQsv3fC8/3EIY4WlBabHtOgzmNuLHPNEisyavuG7SDG9DGsxqKiMGEsmyNS65G
Wd0IrlEVKKsMCe1c7g7NPlsVH3zoJ+AOQH78hauHPqRWTt4LcufV1Ris8JTgAmD46sBGQio5+07d
QOeyNiNdjP2HoyLV/jSKTsuXLp81FOpNpKynxEjnNFcB9iwd2AgDEMNStXrnfmklB7pJIcpAMrzx
wQ13C/9jBdOD+8fxOoA+RfWBhYVL8nRoIVbB/J2OqrjdA81KoS77yjZFci8P6UCHbRmHmw1dW9vQ
B4hm7YqC5k9++LPExpb75ULMdVTmKQvc8Xi94rKBIESlgbN58o6poXSZePoQSg8m3uvetHFT0xzb
5kuPod7T7kgWtKafk4xtUn7F17TwkYgoH2QM3CjIKI4kwyJxtm8aJfvYEGn3ZFhY6iwA7Ezbp9Kb
375s2cnLRHyAA2ri+qk7G1ytTchFO8Bb8BqU20Gz56l2T4Z24K1tyBPiX4xqv2OVSUwqarOFRYQ8
i+2XbmR4K6dRAWj8V01jJEmdCcuc9IVKQQeqmBNj5WbebV3IhgkrN4gkvo9j8UJgSf0nnrCTn9Y4
jOD8gQopjz39hts0p5OdM6+RxZnncuIRFhHbMQu9xY+mZnmjR/lbKdmfvnae0qcYfj+HErPn3a1n
01DKrS6Wvzrs6MfiEb8CABGIyreSWuAhKu/VMwcT1exHJWV0u5YKgGsmr4myyDJRIxLLA4pp6Icl
nST4Dw++PXjwyHmx9Wl2+tghKTPOE1gaYK1bX9gn/zw0xYtdofr7NHQniCA49Q37bwEDi9N0DWlE
ExnLjZD0dFUgxAKgChHSx+BjDxjMhxi1aACVPTRpNdqPs+F4vAjHZmSm/3gvxbf5pn1XoEsRSNUP
tdj5NrhRZ62DIo3jblkPr4d8jBsHnrSqU3cRcI/zJFxf52UtqZZ+oSMYUdpk3kA+NDhuq40SsW12
x0X27CMrTaGVYNZe41EOT8rp9CbW81mftLdGH96QZKw/JNUfGdmxFe53if19lRBBDSYdCFPF0j2y
Be9ExERq4tEqdIcflYTyamLlA7xowvgPIZDrsjHPXc/cKQ6MdF2ibUDlMP5ckvLSmt9aJpPAQ6WM
L7D8fJKhQHDA3Ecb6YR6vv+aq2AP4nI8vGgodtHBb4FyMMQ5zyDpzW1qbMMnpJBPM6C7z0em+ve+
9FHsQfKPdv7dlen55bz1zQDkHWS4dAobKTxHVkQsxC9LIotXRXo6J4k+wWg9FlnZ/eyQvwfrnBtz
rmQN+Wa+Cxpcraryu8JQh81vOxyQr4CX4gcLL30eZB0KcMp5S7xLzuV5b+z6Tshb2HJtYEDB6yKG
qnQUcQf8Txsge2yCQdCpR2NuprBTQNrRQ0joBR3z6fjRxN9UEMe8VxEMqcse5a4sowD5Nn5pmbxl
UXwAr1qWbDrcXoZheNCCGfNoGJcnwCBwxAuen6E0gyhrBqZIouKhmjtH0B1SW9QLuuble/J/OUr0
UKaaOQ2+a9f/DzP/Ea3WL0D5UPszv5iYY9zrWKT74bFm395XCBzUko9aBe5Ato8tLKz1GSqpSo4f
m8/CFoWJs3La93INVKSDiMpJcBizCYBNJFG47mqOw9ZBxihfHNqZrO8iJrq1TcdoMbvtohcxkPf7
mCcZU0XDohd0FEKU2g3P+bLD8cN1n4kOHjmzwiQDDmAhgx/NxXJUyLy2ks5mcSZkmLdfxw5d49jb
ApgVxTExiHATo7bJTgN2KgSSE5Y+VOXOid8Osm5qtxPoPfLjw6o/DA8zB/SRxMQY9cJZwuxSr4/A
A8lGXMfw/tq8NW3oizcBDnynvMmTsBymhUKl5FSnAvOT+x6/N6X298fL/lbBm88LoG7IQgRnZrwU
hcLWduGNjIYrh/gNYMncZtwHawK3TRUm9qZy+opbFoPCPHIwUiIGUepAubQRSFp/0tioTQc7Zf74
6MlhI+ioaxprpQFa6L2YV1y9i2vQVCppXRDENY7qGHJ1P1xJDgDp7ZUgEkctHDl8Py7bL0khUvPP
xiS+9F0nFiEyN/Lh3WFGWOL/7MnKxNl0F3MxKU+H+QJ9xzQMByuwWiJAMRfyCP4vHHpjh0uXI3UC
yFL2B8g+agw0su+bU8yZCJABfoqIrwysFTeA0obV11u2SLDlWmQ6HsoOgDnkLS7nN4TtEPncoIeL
44am87pNYRAeb/skGlWdxuYEFnSqT9iA4x/k034kC83J6yj9m0ZQA2vktMbYyImaVE3AwaphxE5r
OuU0Fgv48V8FEGnNqjSMY4jo5paFJ0SaLijxgwHR1OKscA9s42vWbV0ZsYMQ8Vzw1RqewQE0opTm
1RQ9bGFPNgBA6r/DakVofXER+hNr12/mJ78c6pYLH2uPK6AwnYEleCMLsvDKPFt/xm4l7gpZOf6t
nAYDIQZiStNNbAGD6RJq5FOVKH8dBcxN11PgOhxPLOF/NnTsPW7R5CX7qSqf+UeWRFFvkcsUUJe7
iH5eBnRvaeo18hUIvceqyuo09cdXmA78Caq0dn9bPOhaon0bebLVlnJj+1FMDWG7ghKKPksYDv9y
OPSUCaAuj9dQu9YxO5MRQ9y7AQj9WT5kuwFxjDYfd2bE04qCigdNEBf6FP9j9dPbBqS9qGinGrYk
lLaKYRN/lORxC16DkDJeUC66XYsCDqkQZeyzt91p0PpCRFCvqCLVidqjKE52cM4gqK6XWHxT0mcZ
n32WUXviuzogpm6q3D7bHrnIKsxJ/wvxffMixZcqzX3er7J6FnYpPz8G9++UxRTXSdqSkMF8J90M
zEQE+FkzHxVTBIxS/oemxPqdRZUo6z3Jbq6Cdky88Sq98jE304p0NqGwrG6N5cIQIH1UE7S/jDjj
DVGXGKV5Y/Tc11FsjK1elsURT9bVWxQtviDSTKYlR651XRmAIAZadN4PP7fzE4/j8deAnrna7fyO
4imQUQs562WsS48NL4atcAGRgI9lQ1bPEbbNnv5QSV8G2lojKHRuHquZIoL69BogKbIspAa6iSgk
Byr5MxUZQFh6AQj7mtXelau7A4bVX5h2VT7xMq0o1uQZthmlR2y+5fmChtMkoA7Kth6dd24YWgqn
+BmwbKTjPKT9jsbBdQNR1zHEgsJNt/saFlQ+WSBYyxatp60S02D0Rc2318ycXHI/nzoPSkLX5nbb
y14B1Zr8vpFhpVCqocPK8R/ZXoPLj/MtN6EEy7KI5g0Otu2GS4ubK/ybaqbAfq8NkLx7OFIpJ+zr
ncayYP4N80fONzi75kg4nE1CNUhLbANKA50GQ9F1+sWAWDx51z3GEfCNeTZc8oHfWXEQlhvnihuW
/iW7aE0q5k2soLqq3Q5x62L0iU9fZTjU1rSvj0g8eRH9M98oKLSwmAEZF0MF2bTSRXGq/UAWkNFy
FHz3uqaUVJZegfL3wmvqfIqRH3OOTHTGEtHdfQdFOlt7T3pDzBaHLlCEP/onPrg4armav44hzVm2
ILkwfozaL+yswkeCQlTTYiI1cALBtCA5W3RwBKWiTtygrrhM12MNAklOZRbaFa5WYbQ0TJ96yH0e
U3Mc74TgNRLCmZMrNI+DTtXJFWz7GeMNyKv1LtDbBdnTc6F5QDFDlQdsxlQV0+8GlS3+Xnm3M7rd
3+KstFErvOtogYFXon+sDX6/YDBMXL1gQktqvBCFt3vkk3vpqbbIVFGNzLkjwnAFK2w3LtXiMdwq
NZIUmZr5JHm9C4JZVcZZABImmZ7Cdz7dr3pcqSC51Bh1sc0fnPaSiik7c4QRQXbnwJopgagHDRQI
osgER9VhrhSOhjxlY9qqspx7anDZpk6QvEV9xdUJX4LLe7qJVDHK3xdqYPce4CJrIsGawupXTguY
8lR8GtE5QYQTONvBHut9N9cmQvz0HhG3dTsIvuOolwCA47K22UF1RdtaYq0fDQQz58nD4cxr6vKp
QtoDZ21eYtKDd3ok8eWdsGRnCoDUW7V7AAQcwIpYKjU1++R7A1/U+u+M8ojmCkLU23G7hxzAJsTD
k0CaLkfNicf+ooJn6maWirn44Kg8Ri56JdPkEHEBKDB25OWn+Ia1OMB8Ujgc5SPmdgCg9eIVaYJ/
Q0/OPh45aXXatOMdoFp+c/ENAGpix0sJTtY/DiH7zg1/9w7+S8xTDeLRtqKs2xU1n7fWmT6lsICU
IDwvuh2r6zHLkUlgUUUpX53OT3dOPxdUM+/+KPKXiniW1KAnjUoQfIxqHdDL6ZbhUeMx7QsfVoGt
3lM2kJB2YlZcmviDe1yfDFVJoFPC/zLM+pYbqqd0u/HkuN+6SV+6RXmU/lJpAXBrAv+z5H5fEuFt
yvDSN/lN5ulExOcz+T7fklrWyrL5TX21b61widen5u33gQz6OdwFPNLwXxMdL9J90cPr1t6H7hLY
NNk/AnGZhn4lV0lLj3vrYgm5zkOcr+JoGuMajsR+I3HI/V0GxzQZCCeQ+nB5X74vxQeGYi+glHKu
sY+R+iSAV6U1YPrQ+r7xYwoh6IibwPuUCSOnHje3tRn4uLHtMQKXpzTLljWNWxXAoECKsXZuY7xg
ZhusXkNZ/t2oIsoRfmHzLKAILzUcVqemjooeWL9DBcKfhIx/tcp6po55gbQeWT3h+aAHdjfdCumR
xzFmMUbRXWjQ6+TlIDni0rP+9Yps+W5uyDDx0XleVpNhj50w75kasIaokQmPQjKKpZWYuMb3cBS7
0AB9Zyk+CFkpYQFymr6sMFJ7R/ikXlwwlGQkdiOVAKFyRd1dC2M8G0YJ1XCFaL9qeNa62sPYjT99
7zRaVIyUWg09lGHV1Z9ejBFyAqOKpUitXvmKMU3KXFRv2/q586qZchefs5SI18bOLkqNY/48PDFb
BUjRJQxpT68HxViMI+OG6paiHy46ME6SxMcFBwu4NF5Xm3fHdGTyV+1vMnfKHVO9dQ1j93PONyQ7
eWYnkU5bQiMfll4BV0UuC+bfdok86cJmqhkKM06Rz2nzsyuhIZBvEngsVn+zqt3F39+GAxE83Z2d
A5DSJB97MvK346VSyEiV5RCEz0n6f9GqigpupbUO4en30a06zBm7S4BLINVEmbqX7CJjUf8+eRlj
k+QDUmkdqc1hH5UoTQ6PBDKcrsAvbakACBYQ3obAufAqWdlAxiSOvqclcc+7aGJdXHvLhb601dcD
OCFFesCi3cQSKAc+69iOTaO56efPygc1fhkDqMANOiE1kO1LARsP+MAFciCiepO7AACWb1ddt9MY
0VI4BfYJk85F0dnQPyBOsjpxwvPKc0PGQ9WQ6Jh7W00KJtIumqielyFGrNQ3+5dVlZSRulh7OGax
rcUhByWG2qUdKave7SS3mRCeBJtUZl/ch/Bxw7CeYdy0+Fgeh1OS0Tnxnka3V0L+C+Zxgiz/FumM
va6IjLLldJ1zQ0rf8lYobZzGrZGbxwuMXEUysUj/OhbbMKkX/hqomVKchhnck7uabQ8wTJTkPhrF
RjDaMqpoJQxvPUGUTi0NcvEmpiF+kfHP7kUM/gVuPudVjInrnIafjdC8kDr+euw6GISMHoAABXr4
QcwvtGzbaIM43v9AoSWGyVjKn+devslMv0kTCPjtlxQkz4ifc9jaIxDP9U3FOSv/asVYJmbtbCjy
8/gzJroF5CB90g7Tp4NuTI31daCE5ofG/I7OKDt3QpCTsZrBfmEkS0oeihrncXUeiathdj7ZWO1G
dtg4yh04X13cmcdYp/6RZJQVOwCOSzYqQjJvENvF6lyfgiNFB/oQx0wrQ7+dLfq9fdHtstNsm4ZD
+fPtcPj/GOtJ5pFlUv42xo/UGj26QJLpoBm3NCi649TLgElhOVJUaIRpmX6AcD4NqJv9daj930g2
aMJ45zDGH5SVkhejme327BK0UIXDpwWmgr9ijFa3CrqI8GQxWBxJBJlWoTRYb3Xz4DgonqO7UtBv
J55JJ+Bz1C4p2vXQBt0NXwSbEdMDN9qcAuTRQqSOh1bdwp29g1NhHxBpiyCOSGmx+VCft7lak1Rv
na7+dJeRyFBa94N89+NQWKt3/Rs8/XbmH+sUJw4I4PO14OGngpYh5aeHV1ESeAA3IrbjxwjbfvrI
MczwyuRUff6Fm1QvBobA4HjFajAf6NGZSCEUug7GQ3NtIsYc/ohUM4c8+Vypma8P0wdlkOJ1QRE3
z0WITHx8RAQwf+wwpitIwI2HDM+fRkFiMwA0bWVF2LTy3MTxYb45EqrmMueC2Rsw9M5lutRZzkjn
EIk9zDxpDYGQXuyadJAXzHitpny39HlczJOgdLgbFiKt0spKWG0Fj8KYw6rFaGLQVyNm7jxmN+Wi
PHjJV3XXJkwa8EDLYTHqI/i3Z2urpOw1KjZUPFVUwPFy3tpNmAX6iKCVZgxtkwP26wKivO85ckFB
JcoHdnVVuVqomJckeUjPgGnjO0u5uQnEnAVgN8wpWBjNJAC2VYKrX4Ac3hkW5dV8c9JMyC70larP
3Oymsl+x1ZPDz0KnHxbLLapx6qdiT2BTVBDplmgAQk/TJCjUGC8JOxeAM8XE/gxuFDlviXjSvAzx
X/de7wwyudGTdctNOGtXObwiH2STEZUso6EAzJCVvi3RL0bta8MEVJ7KRXj+cvFsogRO1ZxxPUuy
QqkwRVQI0LjOQHJxG2+0wqX3FMk9kU1sjKTU97MpsIcS9SWqk0gNiYYNEtRsIxHEtRB3KvexRXUt
mFwjy7ni1faPirPZPay55S99NgWs1V9zXwrOfH7BKqHc4/rYK+vRzFmEObeRhZKTsDWYaWum6Slf
9/bWN9ExmhPNjYRZu+Sw4mGEwaaDbvpGzXj4Z0XVlRn0IjbvJGe2YGcSAnoE1ZmgiAYV/6GHS9iR
yZI1N5D8Ei7/kuuzwMi05a1E1CtTp0pbg40BtV/ybu+h1U1TLm6UC4Z4dD01gPaiZMwSE09R92Eu
rFB7tvn2oHmrK0FVY1BALGIF9XMmDzZ/dIZhq6AoO1sLQH8Wqr6xNvzO5C4ZPKkgLIcvNSUgvtUK
Y6ZREvMb8KbZMRou9WcIdjogQbAFgZ0SeKisBg/dSwkKZZrYScszIhwJrMfErVI5bYYOrgBQQOy7
nnjlmLOT+p7vjekp5Mls2Mwk6Rbv8bvameicO6oj+JwX5IYmOyXqOIt3wEKVPR/km3RY/dtDCsOp
xAxCyJt+pt0gr6aAvd1cMu4WgyKlYBrcGYs5f5DN3wj77vnSEMGcB5seOVTau3EAbilvWA29I58v
AAHJI+Ai/0TcNpvOf2VcMXu+z49JtPfsGy/X9562RPXK7vR7DTCYijZuHfsJHeQc4DEMKRUn5qAW
j865E7GposupHsCTALbhkHQ7Zs9hpl76IBbwKpj+ggYqezWL86cRjumhBHY1P1PT4QXsWfCxCZ9I
r2uV2LIdaNyisB1kIZWmKPuDO3R7YdyFiy1Oq35gcKwZbq1jw2vWRmkv1k76yFBD9UFxPyX/8/Kh
eu/LGv2UWlP16+83ibVYjG1JOWibuMk/6xG5OSJVk/yFgVyppctjzcfGjpc/0gyHZw4PfwjeVThp
vt16LnrO+rTS/Ty4ahi+5Ejls34J13+Jmn/MuxCDIxwcPoKKf3yIzteqtDpTiEQAtDAMapircbvU
nvZ0J4oaYhBerimPV43QABNSODhK2pBVLfcY9YNVLSnbzd4Cj0vDkHROKMEN4YvsWLzJu9cinylY
ZINRsl4ChG+4h41ymJyFRIB/RZb4SUqq5NhXsJhYHGUGVOaZIqLByhBSpWWafvU+4EWlfhx4AjBY
yNxffjro9Us/Jqskly3u/BV4McPsSZoMW79x51sw7sHiADLKsNo7oH+YC7m43T97KqsK/OLbDDNZ
+ubPL2qD11g5YMvpbC4ZT9mUExpRHhDPgdlEAPG/jsV3pvUTy3WX6Yeu4McECTGutkvZL2k4wX/+
cS5zZG1khEu9Fcf2oFkBxPgefeQOCnZbHziIgXA1/PXnY02xdijNWiapYpVT0cbmqTHQKQ9xu/cM
VECvhwzPnHYEjPUP0ofpH7hOEZCODZTfNL1ACeatnwMWVI8WuHVmvrk2F4tQTOGf+2fs6IF1RKyX
Nk6vMkpbF6VTSLtxtc+sYoO6wbskajGRX9NhpLaozmRAT6Zcmjo3S1OUZxhanE342cjH/cqGtioG
jilT1raFh3zp+Wh9zI1E2BuPqL2CttJP0U/B1y/BSyyr7X0r/idstYBDhAGKTBpmRMwC7/v0j9Wp
/0bpoB56dcx+8e0oZFS6VTfPg38LCBFhvyQdItE5RPWYKt8F4FeJsFdkSvvWMRatILi+yPQgirX5
Co9QBZrxg5KIkKIhgg5IVpLFk98s31W1g0F4a65bFsAhgfCugEcHu6wsDQI2h1SNUFJOkCAAHsqU
gJ9qheYzTCpAE5a9Sj0z77hpOAvwsIJ0rHgTHrteRrVbgKHu7Ccpu+rmPZoy8oJet012xSvZmPhT
EoQayiQBU6oZeEi6o4pHJH0xiUMdhkKhBoF6HFcUZpajwi8r8IHj3LIaADlKPUdB420ifFIinxo6
+WeDSd7WuNcAUEtYaD8ul7aKQHuLWdyDmqYga6GDY3t4vrlrxoSBmCGwNjxcboHXjDjuLpdzYtoV
tm2VPzhOUYmeBHjXlxpZMlCEhTjQXaFeyB5VuKSbkweBK0zblw9CUG2xdiWxyx4PRbTP4cI7S9R/
Qf6GvLWg4VM2lZRhAWX/dzvi0ojGSPtegUPgdqyGPaNV97FIQYd+GmCAfAtfU0GWRyO+NuWSNKBn
2d+PW0VG9/DSipCxj0r43JosxvqS9Fr4QEaaR1+kxmGhpL4Esa2la6bZYlTJwW+kmRoQiMnaRels
8Fdh4lvmNx+MnvGoaYfaE2DwUQ6M0STCinaO2EPORl7tpt8aLnWEW5n6JnCwC0bgq+fxaq+1m6ao
gytDOrYwvhuhPmOf4ginHIeCkTj425OagDLM8ue5fqB2yDem1G3aKAeF9pIv0GslP4tTThOuvB4M
Qi5QReBo4ct5GbQY9Gr6C7X+9qOl4n9H4o8rnuCNXJ7RzMGbc2rjqNISYEOPbWRtApo4NUPJo8Zx
xXUqgT5Ch55ZQsIZASopN+JyBBTGcpSYy7w5v+XLbQjkeGxTuy13ElysQSpuhvy3stDJYM/RlHjM
bFjOrBIC5emSicMFubO1ah/2qDrlWd/fA5/s+1RLes2oB9aqtxVx+rcky3SnTAs4dueqvca03XQ5
BkDmo8mqkTUEYrZ1N44V/n+XLj0n/1YD+qSRgXJZAhjx0yrii58T6PT7baoxPGKevG+CYYGpB9IF
l73SdRSLs8eHimny9WyCd49iOHSQK8PUj62l5EEzogeeDEEnJrKmoJE78tjh/U+j1qjyXOO4W+iL
1vWJkMw/YeqoP9HX5TOUIt8klWObId5cF6RFgzPU7t+FSoFjCQWWYQM4WL3KlZ3cANvxzI85WQlr
7gwK3t5vpy5Ti+lxzhcL5yYzRFWzI2qkjLa7IquHnqarXdztIHykqhfG1hVl27ukJyjwhtCW6rpS
hcB17EJnSGWwfbI611evm+1PlaqDyWCrg76pBEpnEEyqXX3WOBwn99s6dwksJ7f0ce4q+mIyBlYV
LLayy52WMnO/W06qQbl0GY7TySuFbt3LabfK+HUvCkKNgSH4BAH9PzoM2w95L3maAr0Ga2kOssuN
vmufmlXnzUktXggwHqMASvH7uBPMNAOJR3GbUsxLZUydpkuvQUa5hk7IQThqusRQPCNRKWcvUDFn
GEPKZ2ptlhpLmpDtZIb5BEj7lFxku5Eve/UBdVr99eoyd94GJeesj2Pyf+EZ8jUC61qYpJUGbVU+
ZJnaj0fzNBBTnPhhArnjLJh3HAPOKnkoEEI+5nP9o6BNvcGd5lqW1HyOLLe17zlef7cg5+BVdWvW
yqR99obH6jGcJnfCE4h4vFhGQ9++aBW8XunX+qpXtD+bNvZmkGiuZg1hemigO2W3SeD2mfbg5PsM
adc1PM9/7DtSGQ9Hq60PXIwXpCE22N4eIAaPqRs5Y+UlOyxZ/RuU8rpQZan5LTF3wYkeQ7HdwVX1
secHdYvx1qJKylqCn400xP/wPRHBuoe5rJb5skQjnvBFJfQsE8lOT9bUXCyCH3macOITAEy/erfz
Dr89micHJt0KyupdDN9+ICUPDpuwRbczyrehVZoHdsqlS25yq/7qYo+Q9xxQqBWBH8Ff8XU/iCf+
uESa3qi4ibLS+hZQE8uLQPO9DT205ZOcHZIU0/bVwB/499KL7m0L62zbACgo0H/+aIZtkRzjhsZd
1irLTe3Jz+Zg+kZ5vFJu8jg0E5rinSlaIX3jt1tzuKWkSeElrlU2DSAK5MA52yXlIAXwcm5Z0cV1
LqHFCFGYrkfNwvyY/WYGg6jC7OWsLhC/lUGWalW0KNv4BYUNfa51IYr58LYmdg+7StzSV3eAXGrq
nLf4qgqtNveno5W+ULYlCuq+xe9bmP0MRzM3jeTJbS5ae2ZKf5SKB6ibd3MrlUuw+PgK47Qlwp6c
XCL3X9uCY064DU1iVMh42xHyRs8AxCvhAz222L11pERn03TVQjkEPLT/59o4EiKE7YE8ULQxttEX
6cS89r8Tf+inVi7Xj+c9MGN2OHlGpmuOHxYokncvpsfiZuYprIWOze6tKiLeXhuTE4y7mx9VVDeO
TnKcz2/zdgYc/DIzA2Tm99zVY/DtZZdXsVvL89IvGzXyuHMh3pZnXVztO9yOhG90Fx7XnZozOSL3
ljB7P7DxznseJC6XnJU5aae3djTByO+mpg+sIYqG536xnW7ffUC4/vYbXDcFZ/yEQKY6kfCZ+1tk
P+0eRWp2s2/sC58aQNNsm6Slay7A/yMYsmXLHabWMcsEYXH72SgZOl+vnaFckt7YJjGqF0fLY9DO
JNCHxyq5Zx8AhIWSV03f35UvYNluTqP2fGLki/2M7ggU8MYYYDOHyNbu8YjiS7UXzdbWkZ9+HmZN
5i37WJjbjwRxHkGqAKqLTBDyfZnS0RiIqHQPur/sq4TrKYc1DoSOiwAAw7kCMDKjSl5BbMms7t82
KUzeUnm14kuwTq2aQh80Rv+4UkmNRLiAiRZ+r2uxOSVCFHMs/qQL/zoU3UPDYDpUc+FgqD9zXfCb
UxpS9oDG/U0uoFl88iG+wAYQHW5AsXKK/W8p0F/7i9CSe/RfInUb+Lg4pItxqazmoj5Wk0NICQE+
+gHpS5kGS8pUaJXyUx5AZs7ovHBjvaNRpz7LwczmM4Z4v7TPx+nrurLZlsYR7XJ9RyNAwJfCY19C
ajcnSqhLV1ImWYmWfDc7BAJxVKeejYTNdrujt+5LiCXNIwdr6PL9GGaBxLBW6ZqPfzqWD22MoDC+
S96HcUKbZkh8zKEm5e6vh0sX0qUOxNFr6upegkeQqt6qs/UrNJhbr0amf+tDwKJADyG31IV8netU
UBWJfI8q4gUh3jc3b2DfqBKKaHzceTEH+QBkn3sakht5zaepLx8iqDTdvcg8OdnZZEWKftLasCpm
vMZnNTQp+M+a9NCEt/U+92qEZwhViXzGFbKIZBFOvnc/emFWHhLhUcIDAtLAXMUtuV2ftriaMvvo
vKfEOyEWhGRFLgHw7xmrO5NsKsog0op+ustOk/ZlPCZrI+Of5D71+wQo3bNtdxg56L+FULogwoje
LPh3hPdpveluSmbEizuqyJKrjeRJDPEwtxnSKu0LbUuD3IRhsfdHiWKENGy1kgYIKLmpOY6LhClM
rYz+7+3n8BvvzRzvk29vQNboLQaJy7JBuHpl7pnEJ8YJn9MFhr+6SWh4olBt8gZmEAED1yP4ZKyQ
gJAzX9V5Pfl+nCYesBSPDT21Klj5YJQ0D8f+n5GpIHUc/ag/lDorKOl07p+z+8cFvvdGdKebg32K
VsKRanSeBPF6Dyy0sS03Povjpb+ywCtFXljd9TO5mTrVE/llOB36Ss0Fn8FXJVrKVP1e7kVknsoy
W4AJXDCwyFicW7s4ey44A997IRFIzBPm9fzNiwQEbRsk6D48CQuMgrcKVPDKTJp1eN0J0f+P7V5t
UTvrsiKBeBNb6ZD8dzwtY3aVF/gJzXWHgTrS6ESi8f6TPodfKRO4hBUKkq2ui9TN3Fk+wIC9SlGd
pz2+iKvbNXh3Gt/e2ItZ4NmehDZxSgCKpeLcW4JMgUSLo7Wjg3/v9PNwH/IjsctGV2TzrqaC+GWm
fYW/8XlhJjlR10yaYhFIRGF63VCc9TCd4znEBX2E2KALcvcbcpNg2GdMN7Fh63bJ+fJn458LwKZg
jkessRwfPpBCWWnKCmUBERUa8eRpy8kwurbP7W9a+M2OG33I8k85f4D2N2zvvko7NYW97TSg57Ty
ueHGqpQ6EXfNwy4nY4oS0RWumtIXF27AHZI/OrjjX1UeHiXC4cneysysg3/bAJm4uWswgGlQ4In5
OoK/Ox57h/44qdsspyttsbdruAAs7ZG5tE3CDLp+fgyMhL7CMIRe/QN86ShaZC1zG8VysGhapW+o
iQM8PR/dDxNBOwc2qlsvkzyRWn53WauKloMbZ64yRcp4OVrA6FB0ypTT8fO1camYpGVgmVA/M57t
QaB7d/8PXsALG2SDTA1c2ygDhRUIQGfEI33PaNaz0ZzyFd00YkBnIOa1H4PLcYF574Q3yJD2DVWg
i+c5f2kUKdUutKieT74QWKn+iC/20OM22sNOvhL7CAPFU5Zu7q0smWOIW64yQpz2Sl5W8j47C1Em
GfFjJGlC6RgPB/bBlfu6HhLz2lFF/oXwketNLzZZTAbD+O4utIZlHB35yWjGZDhcZBlIZsqnNRwS
KrGyY6/gbcru4MPbG1ki2Icm7KSF/zhEGSyppLOlt+CiRhkFQLg8I/yu/szFPKpzxrE//6tXaty6
1SbDDflZ7lXyuSAprFfBtqUHzDFWh0LBw515NwQaVk1ayOQ6x99AMgTjJUe0sLahlGkyawJGf3cA
9nmvFsWnbe5gYg8p5tgRRBtVt4cljkmfpcnHaU8BxkC14RZYSazNUkhBydXwZ697lO/YpoysZt9q
TFBTs/Z31RHyuSMd9T/+nRXJzNbflscTLZtEcsylS0+Fd2aPSSDlbe4SczXfQ9TP6NOrqPFnIH0B
sP+vHLP6tzHKAA2Clq+H2JnSKo7fmDfLojdt0IyTxDLIdyeAPWtuFsjYLWHmTIjguQzoyAxr0h8S
Z4ka14ubgc5U8L3GC6eH2865HaqINWdu/rDJVBxZuCO8Q6CBOMPBU5i8qOTe9wI7ZB+qwbltFgCq
FVNoNONzG+E97+F5eJYCoUYBM+iggb1Bqp+GlelQbUwpuOnVY6INSe6Aww7jVWnZSfnKOkgk8Jws
e+VQFsrIGnL+ahQavyuCM9MFVVjCkkszQLSkclXppB7UA8DIUGgPr8pW3nMER230fTJ96PW+DAz0
joZtP3z9pEXjk0vmPE1b/JN41ajcY9t0vA1h/QmrRorZRuHffFoXWFAVdyGaJwJBXG0XZVrZM25z
FMxj1EAwV3FOjzRjSBl3G/7UYw19JDwjNV8ymhRsQtMuVNFFgtSlWZZGuC2u6tjGYX7EIhv9Iu+W
xfLJZQUtMnBwjDK9t2OAyllfcr6xeQZ66CTqlHlWqnUeLpHuLs8Uw75CX37XNqGEUvvhzbGxq01M
cbcxQqK30HlFNhrt3d/50lgcgNriI+Dv6WZvCeBPWyG8gUGKNJg+IRzftU/WdzChs4gG+0N9ozB7
2cUdqfLWs8XScbs4+r7ZjevUErUvHnG2oojZGmqfMSS/8EYwlsssf0DXUOBSOtBligrcwgeev8Ta
HqRZNni/N+MpYoIWpL68zApjGvm5rfBF0lQfrxDtmztBFDoknadiCPsKRW0HNgZwADm6H2NfKy3w
7PxvjyK0AaiDIx74ep0aEBipqRopQv3w4DT2lVvxJ/oMhhCE5G7QYtkugyBONssvCIhIkeR/tFCg
KuFDytTfI0B7A4b3+WUqADUIflEWaMohHNQ6hwSD9J+39DP6mLE2rNO0/i90on1J0t1DGlYdR8aE
yh0nNaJdy2zUc229QoTHWnCaAgSqu6D45JoHaGOIaB4ASupBxHV8N5rwzL1AsWcdaZz+XzvdZM7H
DfCETB2B4yUl60DJgu8Bt/uHdNQoZOB1m0Gvnq638wyPKF7l82dXEFJyDP18CPs4Rx8rleOO6xUf
13SKHodKen9wP60075SNDS1R5crz8xef2gshH2fS1yrasT2U6ZD0VRqwWVJ8ukVSn8651TZC4Bvl
rmX3l13eyvPZAoSK9ZfpB7w606r5mqqoNMIH6XkuGqqgQNWfYK6BWKSpfPVVYQ6qh8+pV9JrHjYH
84Cb/m9lGxyX+M7QfRads32bzql2R6fOebBhH5WipBcqUWl6pehTEvOSlsyRxgck9XUxB4TAvE9+
/BN84e2UhmbMi1zqhVIx4UlnDv7E7Yw/iha43kn/d0cEc7iha/VeA3wxSMTxAnEf3EF8cSrPIbjN
DeQvvdMyB9Cet/8ZWuoF6Da9grO+cOXKMojz0J2xgcvFGtu2TOjHhfpbFdn2YtNdPYhvH6Gl0O3f
lJOTeDLgsIDFiGVBqzGgqDpnS5228vt0/K0IW04P+Aj0DWDiPUycJrkKVHCuVIhuJzS1fS1QA3rc
X8+du3/cIiRCgJZImXlMAcrCWV/kX5tWJSyWmflJXDXPIvT5PwUjdEnlGH/5/uYVC41pzfk1Dviw
C3RzY2dTX+QNvVjkivnsQkYzx5vq2lbQD29Iw5DypI2MXjgYYBrRuu8laqQh92BnNeAb1VC9hr2Z
es3HCWDkGiaLIrd5vmdvG8eDX/iM4prJNIb+hwEkYubUpS09CHwmrmsI7TB02HWJThH+ROK0hrny
oQM5zl9jPBzWYQQCQST110bx49yyK95PjxqCYQWUNgzFG6Kx5QH6rCdnN2TDurK7roEVkHR0Llbb
ZEXflfokobea2nUMfC4wLYV2FhoLDwbF8sXdH+UZSYHXmYYu+20lca61EVDHyuxMnujdoRptvzed
pEPNl1Hm2nWkPeU40zeKZyYnOh9rzl/w7qRUed53EpFjPwZmJnxjsH2PPaIenETCDVxwjg1z9Hqh
K5vz/60ijmClVnKRk5AbFd6mxG9Ow/7UwwSRCyDhgDd7EGBU6kQInePS3XB47glj7keq8o7Io8+n
9mkKiraEXDFh43OkBPHGnMiMYC2NF+YSERz5z7hA9ZxOvKsxGrCwKURNabf1rlZ4nO1g/IoTD0nN
sdJ1D/V1aUrTaqXUAQ4gyEf39EuIDpcXzZDkXBkCnRW1xmXEvFK9MmX84fFoeBuDxbSc8uEYH3I/
o6h1xsh1N9mKs26OnzBqEwHgXgbkTz8ZXf8z+1jnamIyoIbKxTACvfXadY/YBYT91PkTY9NkRR7+
U9Vm3fMIbTpmsaZcByI9ZpIuCZBBkyEoQfmx9LT2oCgaiPSw26a5gr37to0luVUY5g+/kLYzghzd
5fTr5IH8clLCSH7WJCv8B5CWMy6n9lGy4cHJzXsEJJ+LsES+YMRLDbMWIAdyRVZdVRtCpBxlVvbZ
yVY+Wschvty+h2pBTL/1R0TnRM2FrzRtlHsLnRqdwBIXXUqCf84D3uNJQ5gzyf66Ez2BlNJu4jab
naoBHo00WPKJVcn3Q33fK6U47I6BWFRF0qEK8S1nxG5tkk6EH56xhfog/PlIW00Mtrq8uHHYizXa
uQ57EeZ8zOJllid1Txl3qe9dP0ZEagoPIjAugS90FRerJvrtD0kW/wRfmd/KXC+Kz7bWcu6iLaCy
fB5CH6k284I5WjMzwJ3EoEQBpoukqbUjVVci1ZBjMe6lZbtaJunDTpJheQjpks93pivV6BitK9Q0
BPNN7gkS56ka6R3wfONw0Dy8wtqYPcfR3EVYmW+kufNWwZ5skgsaO2Ol6ePYcO6c4fLb+CfBG59y
ns7ksq8kyAmTH6kGsFfCsRhzWb1Q4zj5GbvaG08b//+eoVsQWdtIhuHeSmFAUudkE2WrNmTXGrjh
un4ZVTzsriHOtpEEOqzLPG+e2/N+clxfZMryVwAXwmZz3eTVDCy4oYtgM65tEosjfesppH1CTKeI
CONMMKgnD56jER+E1rCuEDvgDpfQMrcGfSVSsa11GCqDU8qTLFHbVMGjO+bG6UOv2MzFCPFK3VBY
uABoG1za15ae+Ev4K3VUmLHRPRAflfU7BYf4og57TeihV6SeyINesUPFIdASyE2xpW9ikJgr8L7a
y113ejfMinAB1za53Ls+cYDWG7ADEbmnSFTcLY0T1onxNVOnGeh7v8VKXJDc2CK90weEot22No6g
totvPT42jPMG8cVx/9nqpLzPsWQvQz8ob3XhRFq0/+yureAIYHuEG+LXsCc4+Cos2VAtBdAUKBz9
FFD8cUt7HuZOGJutcacsxiPoqHwP0+BRxuCL9971YIZrIUChTO2Px2buVFsqwJed+8hDzWZdqa2O
NL1JoOfphr5VSVqSqTIUlJ4BdzULDZ/8laiH9Wj7vnFsMUkGiykqK7qgcAPYkDrZ+IcthKOz/BHo
uBQZXhZHY6DFK6shSIanE4wvvKaKie7uw5NXVQ12YuhfcZNhRnTWG9WQQN9Ku82UhdXUmPPGO1W/
Ufla+atkrOtS5D+m8xeAR8jWFoJdG8EPGlkOCkvdyO/0DwBEC0sdh9/SYHYcBt9WWLld0hGuCqKX
DC5aQ8K/CoMTW98F9Q1kd49lgoVLfZgDFl63YY/yZ9v/TnIgov0uk7TcVskdo98niyjfkphutHxl
94UxSTW3rSKb5XH1O7FUcj5+Kq0g/F0zB8lWPYdyfDcpCDWK9gvTp0oNw45qjHrtwTvvz9YEUoHk
ftW4HltOBKCY+lgUUFsB+dc0F6MCPIFUdetAHrzK67wj77yai5Ku0JXKDxPlKY+WpXOC19+4v8yr
NzbiF4ORE3XEHcKe+ukdjrhDnreUYLdZnNTYTHTXi88SayCe7UwxQJfcXI7zpI9rfDAXG1Fs9Bgi
5226fnCI/yklMsB7lMv3qC3eE4JZ2AvRWS8UGmTJbbJBBmuRP1KdaBxd9V1IQN3eCvmAoWmfW+JD
HPsWT53i1GwenrdHihqLdj+nv/dX9stHZQFC/88ZOyDuBFdyE1GRrB1lVQkwPB2NXtHeXKQj0D7s
cbj9kwZ0saPNGtGPYwXKlPcx9zx3ongzOW+WK4t0JzzyBB42MwDm5FtgtNg+1F8L5zNchOkmBLQe
TCl6gRtNh6emibh1NsB9riZifah8xgTAbskXEi6FBghuFfg8VWcbJXTI044pK/WcSpnVfyhzMQTg
qQJFPnvPb6raQ3vl9mYNK64f56g5EsHBlS9OYnsaFWKwPgH7IeSc1mShViOyS/PWI5Qcgb/eUbJx
hOC/AQGJrYTa5k5haTq4bAwGrOOervS4O+A9U6n5JcARgDQW4mo8cqFLy8ErRxRsH8wLEerlFT+w
Z56wmmNQlz8Z+5VMfxpnt34lZhXs++HA2FNDfvBt6PB89E1MVXIDQx1pahMkWmjwq7q4T2Gyom1X
Q1Clc3Bw4qTcLnrHtVrPCHaJo47NQaYpdV5KBDdyWEvPS6YCaseaI20VyojWRyg8udEIBYDAlIRJ
ZPvoQGhs/2KRiHZJKLMl1QYVps/B6j+YHIRq104D49YFXnx3G6GMBEdfQgdyc0hKk0WkpylW4m7z
lPJ8E1d9jTzF+cW51/ANN8T+FKUAgMHW2x5zwYELFqBpLdCyMBRXJdqLfTkcR3PeM9/kbQ/nMWAi
R+opscNZL+ZHKPMIiTUALZOtDhKvvQgzEZH15hP06crOiUzzL1AMP6/eQmMCZfnpooZV+kuL6RTT
K/tlLPOIVF0Od9gPoqWSVQz5YLzsCCvA7D33js+c0FkTpDD2r9OVArPJ2NULPMhzbYwVDHVleaOY
ruDrFCW3IovFxaKoZsOzf1wyQf40TErVgIQ38DgvUJiKAcmdgjrGh8QQPDOqbUnq6UIbORErCIT8
mCKcgogrkY+pxfZzdboXp1F81RiwkBNWiMudHAOgoidsZ8YYhdFiM9SDtsj6TH/Iu7fNATZpR+mU
8IeKGPiQddxWuayf4L2FIEb8H2eql+oKVhAQv010jKXXnn8HznpWMy+0G+9Pbz0cLQhk/pOjxHMB
Fz650vKp5Se1cHFJiH0/lDgjyeRN1bSwLcobIdJ23GVcfCEIB3szjhoTsPgWcAEQawGmCY6aZ6pT
Z33044Ka9m9HRXVO6vVNNxsNLFT7HioSJiWViDueKgVSkC76QBn/MBjySu9CVwHVBAO9lBcv3Wxb
vdIqaeaqNYlMC3TyS4RdXDIiWW5KppuaSR3MDX7bKJ2Qz3Hx62uifhYCGasomck+7q7iLXiAW/CR
uyKrSaCnbUvv5gYocAo2y4B70MUkm6S1cUkKmDRTS1oxbaXw1KE3oRcAoG69lyavlYGqHxl5q0kN
vIOmyvO0CUIS02rJOD1lKB8AFSS1Xq0akP1vjQqK2MAfys6Vac0EGL0WBQDmSWYR2ATWYNy6bu3a
e+zj2B1Wo/2EvMNNX1gv2YUj3j5zoqyWMC4vSmhAnNq6b6zSmGaQzm9iRNUl9XlBaXoc7ChVLaX4
y7t/Kvue+WDag4A4sJKFJMSfbs+vj3hUejJ1N/XFO3ITRUZhGlq8uTMWuTVE4B8W4HZnlBmKucNS
oTR1scKD0mNDTf3rThmu+sNcx9ELm7XG32vF19uY6FD77uUfXe+UPNbtKiRTjw1RuZMPVgFKuVpG
7Wo+vJ3P85CcnFgxd7ZoqNrethcG69hYGPoOyFAJUd8uMY0emNO45GJJClKTTvfy+v0p3NF9D2HE
nwDmLDAKhVMiEbFHQ1QXTe20bri6IL2AR3Tykc4dzaciHWZcNQ/5wBERV4Cor5j3E2pXaW/K3EAL
jwmwQ8DiA+DXSkJUKml2pIcRroyd26bGNtKvMO+BDagc5mR2nSwgAScapUWhKqNYNZbXvo/Gti0J
p0nUYRmAS9M7+xHmxFlpgYb44pqEz2XGW3Vjsp3quf9OCUhM9Thd1kkeIUYJCzrZgZPa6r3rBAnW
FeUHFgidUlgdKDKzYoR1SZa1v2OSpb/fMMQgPCBwFMk7YxecNlJvhMuZ6E5IGNgz5iNA3QFMVr+h
918+yk7PyAzJQDyPzcxZdTZsFkhh/D+KoVOErYV3u9shIP0ey2BWMbb71R2dOlgeKyQJdshbXLkm
hAi/B8xaO4HDRiQYW9Rzy/iiGLb4pjUBZOAhm/o+aDYQNgswZBQxrsmhKU2snlF2YfR3HsVckVdj
dYw7/mKdIc+bzfM9vztyfVkc+EldNbK1Jljw9WCYLid8eHsDv0OtTe74zJbhaWXeYJ9bYbw3yFDO
Ex3vzhIOX/6WeqgCTe608VBTIDbfftHCxkj2UQXNKnX0Ixn8CbmKy2fMHlQClO+OmwqhaBTzLMKN
ie4fHCmmmDl6xb5GvnPP9b+kamyuJqyBQEFZY9hIXtLDYCQ8QXS++rHgYY8Pshe/t95O0XGNew3S
N+rCXnMkwuBMli7lYEMev7zghnmBAkyy+5lLIXCnsYwwYlKZ7gm+zwvXAJz6n35E7Xs9d8tt3YfM
y3JPJ5XgUz+ZXcaidilraouXuQsudfx6V6iQXtwumYiofOUpf0XOyew+3B0dpQGwhGNw7cpBFBn6
+0O7nU9UsGokHeLwzzddDJ3NbrPiwCRtz15QWvkW+cPTdS1aMlVdx8RXrn5rUzs5gwqDOLQs5+vb
Ri2E7cW+9IkawyqPKXbfAnX0AHMl7ss4JiCm667z2NCXbXJehO2oa8rGOxRNwLtUnIZkry99iPyu
am8nxtP2CZK0eBET1vrzhYtp+uARWpxiipEbqxBQAJC2+9yv9mDEUfM0avXeDie2P7zQvqnP6XYe
BLxhNdOek7p5QgyCqg6Nfoh87lBCIWTQrdz7i+lk+CeZLxJfTATesskAvHKdpCahkT5i/Pa68+6C
Nb9uc+Xr4w19JRANUuWXzI8+lokQF3di/w5O9O8je9CisYRAsPIHBHtKPrp9DGUK9Vb0VVFrQW8C
5DatwI4QgqAohFoJgo52pbd/Z8SXeu4bl4yOEKaP8+ik316n9kLtaAip/nuQRI4XTmQKi02QDpF0
6zHmp+5zRWoQNIe9uBNVw2bIgZIye0kiZMeRTaKFXx09ymHU42B33ngOEksG152YnWQFbrbhkWoU
x+3nLji2lXB4fszlPtvDvClcLC73a8W+INJMIOWTeNY+yAbRFZBu3Q74eJO0/ym5VqxB1ZrAVsBf
yMCePFgexfKKMzsl3vvPz08/l1GyZT5gMs3aC/t5/PF+Lzk9QiyVBWDhNZy/+47biLv6dnTLzcaB
CmdSjw5CQQErSMiprVBna3VO4PHZvv/tAvzlfY1Cys2FgTf3lJx8JaosiBfTPbbRoJI43WOfH8Ai
HLkakfyzWyLJf9i8P2i3W0O5gu79zJw5iK28LbA6Rg0q19yNwed80jw6hS6RcKuNoVKZLen7KKHK
DqQ/eNRw51mxv13S6QFAGFdMJmm8X9KU8rb86UvIxW3lQUCIzYodtlfLQi+shpKp6B4aCRj5x/3q
uuBlLbEFIQ8wILy41YKUqHu/Ro6YyYoxjueViI/Ft8HiX0AMvyDmi7LpBF/abf0QQVtr2BuUUNbL
D22LZsrKRxkmCd7oY3gyqnD4n0j4tTnxXuPt3U3h/4pDF7jlFw4d9m5XMi1NDtueT3jlnQr9jnZa
GQScNQqKOc8+TpxGUKcQSXX5MT6cKAhG0IrP9DP76AKjkRiTvXmnzO4pbjl7DEqWwsjsGWdjBMLl
KtnYCsJtqGWhsRHs89vfeAWADRaEDGHWMpjWx8ZSBlWZFNg8OwyB2DTYvi2iGv0589p/7KIm9s+7
ZTIJ8o+NMFydW/4gF2Ax24LSwyWBnwF8wtRDXooa/DNIKxFShxpIqgtkkH53uuNVpjWZXdYbEzHP
N3A18xtHjVusCYVYmHgLPRyPIQgMeSg8kzTAfQzpgpVSFjkiHjWg+JTSMdHQuNiEtK6s/8TH41U2
4BezEn0ZjyoHzVGCgO8raM7fcxqKc3PFLmHHATdJWj8Pw2qL/egbfIVN2e0427F4QD8+dOjjSRHm
9+5wvQ2DdWGDrV2xwxjq9xyTDbE/xDm9QXVkwteE5fEdoU/XNFsERPLvF2ppRoMgr4Hh93D5hIU1
dFnLhp99YhNfZxNAp+vIRob3p6Zoe/PkDehiPqwbq5GyQqW7NBzRZuzjxovbOw2fZpuVJUCPxSPv
909CRyrSkvU3S1e6shtIKKbjpn1/2vvMuyrK9vtl6OkX7n9JMD5vTG0me06zgUic3uAPvzJL/T4F
Y3BOzn76aIATLpjdKEmEaRuk8qc8ASvMty1a6K9W+yYukstqvStClj36xD/1trvE3vGZtrjIe77K
6BbBK0vZPkbLdP8Ew1aYyO4QAqgqdqo1wgxdzrCkV/ZqYzomdrXF8++qPAxEtOij/9FYRZkv+Ekq
E8DeaoQpJnOXEES6oXJ/ztK3kLDYhHRUCIAeo0IluCiSH1UhZ2esi93xWKp2igiQyrp+rpjK9wdW
wkmcZGh0y89UkbupzgX675nnSSzjrghTyBfwKjvBQ7UCD8fbY4ZqGtYc9CdUokc31BB1JIKY3Ubk
L9QWPx1BHtOKOuW9A45TbpZ274V/MtG6nA6KF9e2N8E2xLKNMXa/lPsS2NaYt2U1QNwkqTza3s/a
8cRilYYYQEzeG1Y/fePHK+0nKrYDpmkXlUdgsv69RWEyxN3lwg5zkmQql9oTmbQiEWwEZtSSDFMt
wJPHqzNlOPB0cF+rLe5xv7rQYs5LlfceGz4HO4KEmFOOtRaZb6ZSNVvonhbPSAzEEucl6KmvxtmX
WqWGdOzB35moorbCO0GYOg/NQVoB7KOUmO2D5Nf6cA9lC+raayPc/lt1PksndG21OcPdsoXqEHpD
ZNX6Xe3gYTmDtC0hXM5flRaUbsnhqqLSQwzG0z+lTrvMtynkRYXhiizkFm5bAzvSyGxFzGhIt0kD
dfaRlc+aoMqztwRVhpOoZGlsYXCQ3DSRx6cF89d8D6yU0wf3mKTq16EZSQxMA+zvasaUGjorNx0R
dwknL+FWAg3p6dHTfqYJhXrq3+KYf29odGHhMUHMT8vf5EtA/5qXVtaBuEivIZATHHsACf1CzPB4
K9DtEY2ufrZuLCTFyNs6OdlPh7syhWNeOTD+NjP7uB8B6IOfe4LWOlrjx90u8ljHgdATRBRNvecW
UuTBi3tii/+DPmXXN6fHT8c/LGCWgzLon9gOtRz1CAhE6TjxEG9308VOA58Lt/Jk9Lw+5ZD44wLg
t92aR0SSx+fQLI6ucNAXvSMBOHSHD/cY1mtOna6RWgd3SjeRBbyq9HREkQ3NHX1613jek5vDmDlm
6PPkFfRSGlDfM9jHfWChZuoPWvKCXVH8Z0mPisws5VO21xozzC38ensWZmGq674py2vkSaMgKQRN
uCjDs7U1ktOMEhnKWw5bMD5X6GB2IyhH0k55z7DIuzEOPCQJM6bpwX1gf6B95C6HqzSshDOjsKDo
cVH4o+n29VWCRFsmjkYHH/Fs1aN/wv7+9sWD9VQtXuls0j8OHUZNINkC9K5hZGJ77plgTWlWMdpe
5oiU5dcyXIGSHefLkFxYVSXxvnXaDaaOaK+rnVL0igsQgy0bl/v3EM4OzS91RqaHkpz8/FNS7Iji
YDioLMaUgFWXYsFGNlNi/Kz4ne0Rlqm5tkbTtv0tQSIOZ3FZ9Ry+c/XcfUifzoynLVveThFIfUQ+
ys+cn2mo9pDIgdycl4gdufe+JKOZABIRUxVcP1nLWkVxDQHgBc/TPvLFjK/eUMfbh0Dbh90uyDgF
Cb1CPjH8hAlcnSCy/BBwQ48Vk4SBl2C59eTADOx2ssjtoNYHLC7Yom5UxYTnrzYbx3PNzkKA5bi7
ttF83Otp8nlk9BenxRQQ46cObyQg8NpUfDEmT1BWOGq+vn9XDD524TVQCYeikvuxltKYRoP33ld0
xNV1PgythJvwzFmJ6Dd8NhFC0ekZ+e3Qr7sz+IMO6z0D3tfrXbAJA9fXcJMlEe9mqrE7pYC75tpt
Xe1ong9rd7oHQe+Le7XBFAp3UjK/nGkwIW3BIfegx5quKiLk1NC1FZsNHDXVKcnFK3GByZiAy1sX
Nm7JNAPuw9NH0O68EnUVrqAXRrFVZNHnxsI5eoMFehYKDBaX5/+pkMjXCnJoCGDFCWA1e1LZcT1B
mous7A49rw8qZpjp8CKArNTq/Dhro+HsOuyrxpk2mO2yZrZmOAGPeVNsPQSIXIdnA0llfLSfQDkq
lfJzIPKNfDYMLPu23F6IxNrVYzC7kVxxfBRctCUH19XRYVOmEyeBJuARzoD3jWoEGDrKmt8cLsqc
BS/c9Ry81QqF8heqd884cHn4uRtsr7FoA9gYTDdzP4dlauGOC/jnDYWt83A9Zf3wsYGPm57ocSGZ
iQ6hX+5SzRgMcpWiLoWaZUj42I4wz2HsvmhO8wdnrUIdgDgAu1LxBL5ENKaJ06+be5XxDCUBMJF1
lf1l3OlCt3d8VRrh/cA5y6QEjzgPqRz0UvSdrT8DYgMlRcwuIImImS7Lrc9p8XzvvWmPQn06YGY/
bpJBo4KDhELgB39WBfOAM5tWhS002NuI8bDNZRFm1mLNi5X9QkzLNzjOwoqYQXZJQw/sGMRX5Sdr
T8NEMDJNjGNvvSyJ0O6H0D+60VwXvU4xwkuoJLm7sXkkaM3DZLRR/FeNzvlXzLA6cUc3jn2gwdb4
E6TqAt2xYBnmjhSjS2MXUqfPodBXKdRU4PwauW1RF76OHwFpcf1uha8FzdJnb+lgmDCQiJcsCg2y
wkcJvgB5W98w064aKV7wHfe7FsfaiY8hC1DgghLsFQ1RGEpaq6wZ0ZcNLx6A6zDRxH04/BksGYUu
kJ5NxElMuYaZUIlL2fQW9uf0Q/Bj9AP58Wq9zuNzvepCwdw2Mx+pgaWe/5K5chFHw4AwxT605acy
pjroYEGW1h9jhZt/IPYLw75JGy1IGJcsTqDp3jmxenS3zlbaK3RZc8T/pFYJ0VInMXgkz+9lvUkK
6facdmde9G6/d6G49H9UI/EkwqS3Qggkw6YV1gG/e5k1NsdFd/UD98VyLb6HDViLvY2o5wKzS7MP
HFwdoECASbwBN43t84HPgJK/5WKinHxP9RF2NRKRdDb54Blz8u8XT8x2jqVyyUDxYcKs2noyD5UZ
RyArRjiA4qCFZarzjHfplsY0rOSsiUZujqedYuPT9qOX2QAB5/KoXTO5O+eISMS9ZDnJkmxvIBIM
INXY7dYmhxTydSqX6bB7Hklsb1FhKp+R1UlEoUR4E3u5Ss3NQ0srQsVMvuB2wBMISWPGZuBEMJ7Q
JNnxiqZkUT7U+clVb4T90K+VdVPTbz2eumkKrZVnSFwDHLd4+OFqr2lSSNVqTEyw55+8nGGfl6lw
OeXGGVGJyfqDNGh3NlZRhMUqDGHuZy85iNHzFXwHdZQzmaAvJ1sHXTTbmaw1dPeQ/kmi4fPAgxqF
DUKw2Eo4fDgCxBHC1LBWGW6A7o36iDxdruCt4BmssjMSGqA+apPifZmUzCf8EVL4eOs9S53WVPiH
wd51AEPqcBuLK7cav2hngk1NGQz/Ncmajzf4wT4H48fyhrR5V01FDpGsPNmGR+fDj5/eH/94iiAI
o7FEJ2YrGEq15eTQ068gj6kLL4FZqm8QiWHQotJIahP65FZ6ovIkojEfnQUuUHbM8EtiZcE4HFzB
JAmUJSaMBR4rcOovJZ5CKN0ZppnFQjwBn+1C4kvrLlPm8edw4CNHS/Em+1sZ5cX7j+maS3Nyq8Iq
I1bNjMGyNZo4DWVtccrH/a236KU7mWnkJ3POjXk9L4/Z47Zeur0ani7SK/SepXYUPPxd1DKnQDQh
bNWAC2vrXqrfqH3SirxegTTe3GMgYtv0OwjYJ+Yl0nyzArtVjic+QUFgErFXJNX1KU9hd4S6BmrW
SqkQP3vyS/rKKBjZDdbWdRp/SonPzy1ydpZUxuQtQB7QEzbs/ECRfyKn2abProLp4fSNRf5f8Y3y
mUU0F4pMHjpodOOM8k+FRMSjD/PBcutmnCfzl4VMCbKqsaMzgjv/tPJipnzrM71O47GEwlA4PJ7i
NdRWVpn+IHPu3X9akFt2zQ5s5hpMXzVp8ZobTkIH7L50FBrUDXLE262ZWb8+Vxh9AZgK6eRw9vrL
mEnVamaFzQgh/2TlpBhCSoF1tQL79/B21hcJKWk67hoP9P42kQUC/4J4vOBXn2DNRntLmG96raGP
vtrI26gTOfybQr6fsdNLr9tPtBbU5gQPDOWl/lZQtMRtTgCIUDt1agnn273lVvy7ddVBjIH1Fj3Q
FxmyDIXuLtbyMhEuqZKEpuwv+2e/gPlujlTdz6Zv/tBGD59EGHL9xuIphAGqmOa7rUVOt5pYktlt
VHvPFhzWgjBLzf2n+8OeTLOwgkJhskeksNanm0DSxQ5XJbfDT1JUwZaBYl+6R3jyMntnqErON1re
5q+98LEU9/GCw6QEtbIDJS5NYPtUhROjgMic3k95PPicSZq33F3SoN1yESO8K8/WOwDr5kmfhfGp
K5bfm01iv39lRVKz9GhnJng2IlLdro23Gf/mJ0sv4Mqd8KCXcLLhc4emMsd2azQt/h2q8iyXKtR0
YEsrSIUb9s/EKaEFD2rK1vVeuh5PiTyyszhc94rbuy2T0FzN/ZizLOUpXt+n9h3ltcAW7dTFINJ1
ta261knZvQcSBm/jvG5nBGNuRd+T4f6yZ9DuzbFfssnYohyyUMn4eF9gMUY3GA2g7c3IPk0us7YI
AJ0Q+MOiUMPJ0GPNGJF+/WQ/QqEIjw5SQP8ohQy2gWseBdJGFeTip8MUnFqs79hIqVUOpvpa+Z84
xCyalduAUJK3y9n3GDbzw4EMyOMerdrqg2tLk77ZRu2GuQRNMBmkClT9Wg0qvE0RSuw7qci3W9n0
7K6Hdw5TnUQIAl+CJw+B1wR1HQiKIuQs20Rx/srNQ9sXDCDtxnCSc2bQyc0HPogg1qGfmF8lvdco
i6HP6lYJmOXUt66eNQIYlOaJkqjwuFCCk/8g06ysxvlSwxjdHUzUGu1qfUKR9euVLe0mmXIZMJF6
efwpwdoDVMqrG4lq7kNALupGA4bImElBBsAVPnta60FesdgtUCZbkWr7fZPP5PM5hHKtE7FyOTTq
ttAQCP8WqzEzt4v6wPC8AvPDvaHXu9No08jh79S+JcvmH6f6wdOot9rjpgA0nHheLDzikh3W/i/F
uPelcGfuiXudN6gdawuRgSg9Efud3t+fipuNdOd8JlhS36YoTpkXmr3rKvlt6onGUGexDStk534y
qE+zIYVlLsBcFM+CU2hAzxuof2UJnf6nD/uOyOuMO98509QZIB13h94PDWU78r9VLb1K+iZgGjJO
CtgnPB9bXPNA1EpWQkGIgVSWY5S4mejZy/iQAQswr8UEiGeUXQIX/CU0U+yPCtNfP7V0r7crGIVb
3KwiAvNWKl4DSEzhud5gy9pTrEbkV5gkivQ579+aHQrn2xfBRlrl5c+XT5h9fmwHNJ0vYdj4cML6
K+zLDm5DYdLY0JC5AAktM/kCFKxqFyVD+euM+3oKUnm/Ea+F58/QtElznl71BNXNSwYHe2wryASY
gywZpDwy4cXTTSEG+FvTdyoJgiD0cIas28FWOyfl7aJ6yrcUj15zyIwxkhyku7ebKYTHcjm+S9yH
GluV5uinzLPguJj6Fdyxd4iC2XhET12qEldqidddLtrQVRp+MTbE6wLerQC4waPxQuXGmqTLOJL9
QWGPMb2/qxfMmQo+Bvuvkp2Q7s4L6niQnymQWDETJdc4xgQXBfB4graylucedKW62Kv/LW2R2hKZ
R5yRVDT4e8ZYZNRiGEF9p23/26c4dkf8m8GEsrBb+64u0AM/8dgsw7Dxar1ykfwAH2EgNteVP/0M
LZQfHd2AQOslD+RdWF97MEv4l8lDcG7RCAjR3SAC2QX1jOiYHmqLJY9X18jaax3V7Z1mZpZGyhlQ
2Mo69g/raLsC6qJJbL7tzEVkL1OuD8l48YtXU2Nwyny7M6rlR9oumnzFavnN0415grpjJX2XZ4gj
mv2TJ6MXdrJZ81HpaG+IDRXDZ35dBqv/gz2VKSSPh1BE9zcRRhtTgyuRkh+UN6q00HLtwcW4kQ9k
KtGEo/tGu42+ryggiAbLs8L+GnPg+YQN+5wsAh9xxRSYHEunej5dc5aqVg2jOAOFko3foFB/iWiG
gQq59g8DohLfgnl2YBib1rTeZzKcs2t0IH1ZfNYumzgP38Pj6wB2as4pq3Ak5kwpwqiBr5FuecNu
daSfLAQBqcIVd7HTyqgwvB2jhcWtYX69GZTyyhoj4s/T8Q0EcnsAOmctah5P7TfSk9cRchLMrIG6
OiMSidXM2c26oZtcmlItlMAGweul6T5joN0iZ0E5dhfD+1ugUbQ6dl3Qy/ePpgVHDQ/VmMKrGK/F
jtELm9Bv+liMzztlT1m6g0vSsRnXvbFhYV5MlXYoiTy+1U18b9wrce2egsAod8fl3Od4Yx6gI9fo
73LFoaU4YJErFpu4Oi7VZWDRnDLdpbTyDuCTKiChmO/yZh/c+bKn+O6TLDAGfis8891jGWDD1+mY
FFypsNrfuT7yIq/9Tmc1cb6SFkEu5W0mcqo/bDMLaIzV2DBsJ3T5M6O7DPyNHuj9x0L9wAmdxRwj
h66XhEZbXmBtTnsZKvtGLFDP8zVIWSNbkTubIvvRH1DHGZVj9JIcUTIjS3Gbfd1SMrot1Gq6RKgd
p+7+bULn5mT22DKqYWOwTu8nzFgFamAWStixTdIVZoSbLVESNb5u/BsSiYsQdEIDyoU8pLqF9jBF
0TfgqBnyoRLyQ86thmsPh3TTvKcn6sdHwYtcCYTKyl4uEC1iFwcKvCozwOHb/hewsaYElqZXyvFj
ZKegkZKkU5+M3KCHhWUsBoERQiSWyVilXRLGWlVFbcqgm/szIpWrLoYb/fNpkllCxEn/SwWglrP2
xtPHxByTYLz9tynim7P/pNz73ueViRGTdC2jBkrP5ft1bUXh8scqlfJL3fxBPUAuwNTIom3K12zE
5wO0NM1kWn4jvUx4HqSt5TaqMMKhup4uV13rCMklBro6IXiQQMDzFGb/Tu8NhVPIywhwd5IAytL4
KaCFVCZdVQcE82y4w5gHjRu1penKoWebUa/ycraknFv5qsdRHJpvFJ3jIWLjkSSz7cy4JK511mr1
dJJRrl2mAxJrues1eaizVi8ZlNGHIN05u9zj2S+r+OTtexRZzPUXHs7ANTsJ9e+VvKYCUJ+q5Cvi
/2R/yOt69uHsQzxaamcIPT2KxcdyokcLIJwtCBW8bPiPYWJilIIlteWlisba1RPxjVTmXyvcoMCn
BhXs/suKnis6JJrQoFckJ8OBdb1W+3C6KkokL3LD5/Yjni2/+rOGsWK39tfhdj/RAqnkH3zhAvO0
TDixMZnzlx2beSoFzn07h3dduA+Mb9sJeU5hXpsn+pF/3erMFYqmp40gIYIhoYDOz/KoXbL90FsN
lOl3oh09Wem3SR8P9DV3ycpBWI4o/auCzWQwYbeM7k3skcG37A7HB7piDx8P/5XamHGmByY0EYyE
WdACaO+o/YT4iljX+27P8OJRQLE3pBANfdURhIELmQbUUSk2YC5NcED18ZMERHF6kAJnEJANq+vV
Re+XlXanRtgV7inVbNbetCzeHob3vav+nA07FElkJExVPRFXGDmu4+RqG4ggA8AeXDEx3C2QbOZQ
dVETojsiVDcY92CIX/7ZTsGocxjUlQXXftB9JZYhGhGInGaRcw3f0WHKf/LSQ9k7gjW5Vf8xuMAC
8+t53b4sXAIW1fdBTfj0f4smfGYpBbKcHYqeumze2u44rZWMJ7Hn17aeUDKA96Tfs+9mI+JI/Pvx
MyDcbMeSpjasnYbDxeToc2SdPXqZ/LGya9fAmqYnFWR41XwbTGMtDMchqFeMetd64N8Yqqhg+Fll
9bq0dR+l2ODhTJF0bD1SAOEcapuTmH9ESm3KNb4rej/AYDAy/k6mVOU4vBxYiP7C2vyIqijp0HIl
IySrTF6jdf3Juks9V3NmJKLitzM2XeiV1KpDZ2rK4MmXYEmGUnur7VhIW6i6T/G6DeXK0dgX8lkI
Ymi2y9pVyxqmJq1jW8sI2UjDfPfPm113h+kAnPzIVOVHXC0prsKqUvl8rXQfb2babkUiWEXSx4vk
VjpuMn6c/7cK4+bFM+ZG9sHD/th+951ShAVQDSDJX1REGD3jScAgcZ5KBoP+TkaOZU98dS2PVQHw
xuxjl+zudPZ5tEcWX5+zv8B2V9//QBbp2g5z43dJChEx/42xpMU4mNEnf+vW+lSX5TVfbdzGSS+C
UNkKap0IgDr2u5eRO28h4yaLXvLDzQd1bVJTnGmnRLjKgsYQ9GuwPrTqc7bSm8ktaZV5+F54IVXT
X5XXURAYhLA6NxTgBxEs01UYJXeeknUm9v/Emvay48gKJ7fbufnkcGgZ2LicCkRxg6sCewwFhOfk
+isLH/YCpvMsZVq2FHjaGHUITHF/1uC/uWE9hFrv/i1VOB818LQ6Dj+ET/YpphRsKbT0HMVXwguh
yeEks9tiOp0V8yY6CFmkhWYpm1J+x0huhcvQ0k/VVOqY8MrQ6WqWN6N0nd3SR0AGMjr/UfC1dSqY
1wSEAzgYDp1aK5guOLABl/QkDTJ/s2zxA5udAXek5hQInEOrbuYUT7TBsYlPhZBe8shg1oRpqVdS
pZzYHz8cc6NilLfbACg6E9EhyL9h92Hk1nSYBPs8Qa13/jclU8cy7pCDVBL5988aSacWNvrh/9wh
DIORVdfhZ7IPGUTE28GXiS9+UA4oGiaXrsof3TGdWnlZx0kOTFHIACQcCg3TIx+h9PiHuI42Funp
Fcjr+8vHtoqt2+a6dqY73Y6vYOQMvaHheq+3zu2LhJKohROH81cOWVfEChR12SjWoFwr8fagF5gG
P0t2PED0Tol0Jqbgc4M2F4SregwkFljLVkGi3PS5acXODq0r+oTNsnqQBlaNAOtj5oHHF896H/6M
BkXYpDSdJxV+e1Hj0q/2otXue3luVUxy3+rIv+8/XeCtrIWM9FpVEt6dF1+aeKAsn2SEbD9gmKQk
MBMmaR2Icg+1JZFe0iBl21lAmT1G8ZjSoXv5rWX6Yu8YNt1xs4r+4Y4+6ZrkqnkdhCkUPfwXL5ka
hC71nTzt5E0tIHdhlQFEBl91DTfrF+nsq+XGbGGqKaYUrLKl/1aZd2wqcu7b+aFOOY2kmkFz+y8A
kvl+WmD5io2PbfqUSfsSRxAZPzItTSnrWzj+qDUwfHFSAWGMUF1pI3CHoUrw6yWJbEpWWJt/bVrF
USpRPb3R5oTGcLeKtalJ1mq0gxRJnEMnoJnPMM2WIg9NLMcoUMjPNn72W5+MtWrqBh5lMPDtM4wZ
FhXeI83ITbPVcT9rVxWIDMthZaIsuGB+buwlEb+ql8sa+J71lGfJ8mM0DvuqlkV65tmqqLrq/BZg
GYz57hefUlWHGccqly14/kyPSKZbw9Z/+JPLIbiNwiR4Ah6Z6IbAd9qQe/JrjnZDLXJVJFAtlJJE
kOgm28cwwpN/8iXS+co0HeOdTz6MDdw2d9DdMysREu4YqqhzP3/vrzzSdUK354/6cFCzUKGoI6XD
44OpabBQL2dQnm4FMYfhQmfi1xYgVnLmBclNWp3hLjgr/JKzeQGCxMwg3FPczPVvFvgvU1UYArhh
4UH/7J1k9d8ygrdtgO2SIsy+xPsygXdfyBvTebha4cvbe3mx7pEcZibxlaWCywtwIkPhkhsBEcq+
kY6CawUwMRXWl0YxGTt/j+kcQM2EYX4/D9Xecvgh2xVm4RshVvyasv+I28G6Z8i7zpSPNSUE5EGP
HL9YV9kC9qRT4+1jXgsACXF2EMIEUfw814IDEPpNU+Rp8MnY67Rn6R4S7JvN+Q/84i+ltijQBRdO
AiOJ6AnvLyV/i1SXM8n6IJXyGHkcMPIIekewYxHJKwhdPue3kWz/Nk0t8njWY3/NsH92WhMaXS8+
VYlwxKm2+EO6yWt4mqJthv0UrCqgu95vhTSyPVkhhu7SGs7DhbAFOSNsUytbOFcYHVdFkq4BlRR0
4+zQngWvgt368cfVzt9tl9RqbL7xXBKZj80JBnHijdgZMEHIcbODI2Z0Pdbnzc6G2FiUiJRvDnUO
ifI0yoeMc4Viuyj0PAfU2jfZFJBc/1fgEOHfREThbjhtceiNkrlrQqbelpGxA5wggz8bA5yzWDIO
DcX3UqKwqKdN4nQWJQUmj0RLEVXcT8oG4OVMPWEZkvI1O560/ZSdDXkXbLLlNfwQk1ZKly6FMlNL
vyCgRc1y4jXPETdUVF/1tP846IPFlzfH4uIbvuFG6Mt3SDNGrNuaZ3CkGhRrhSDnOXYeSfrUmVM2
6MEx9igSWBcLnm/WPTCcwijbRrUkgVovzFEP6125SYgBBkvz7cfcAOSAOb31OoYV2MxciMiop2/L
R58qgNxfjblTV63lhB589IhxU1nitZnFCJwGao/0OlypSXKXvCxoAt2B8PXgjlndLrYd/KPjSax9
gOX1Pd454xNrnTRkHtaq864Heff3kUsgevSTmMSftheWldVo5JUGNas66EdIj+25cB1PZP10LCPg
cTMM3ei2y2la1vP73tWhsTCU8h2f55McDC9ImLoah4obD7DQkbYY9jGvSukIAQ7l58c7/On8ICfB
JxanpXIaGJzmEcT2edN5xN/LaQK6+UJE9oAUId36bqsbVsOGMoRFNWUMN3DWJ9qe/skYBmrIriP9
J3VpuSIRRLy3zCxQMKn1xzWwwxkFC1yoi2xFAgPzmmBmtKG7nvknGmA/lJD3i743jyWyd24+W1rL
RqkxmrCUz+p14ymwB4qKBQ5cHOkyXgoEYXlOTQqPvX3SupLAybdTcuGScHSgHMby7vDz0m5LrxzB
jIgT+hXT0b/r4YNTZEqMhVPuaYhmlyASMb1ZKGoyrDNVHvlm+fvntfBYdYC4ilF7OdHwByneu7ZJ
7AEyOMMeqUL55zbLAyW828eszBfevgbLRRDkRNQgvUST0KrBByyOorDlfhmbPCH+mWglJMw7p6L6
9lF9MbJKV9QcAIdlfIsYb3fSYs0lIHU4Ih6YtCmx1Tk4rHcLg9vhNU2L2/7O9Vlidhc18uUz5iyj
yVbeZt21S7AsszrPBKy2CWnvqyncT7AmFATLDzZyhvznPkA4coleVWz661SF5or/HEv7T5/HzsA7
zyUe/3oV+BQ4429J5DWeW2Y1nZx3MziSuo+rDlxFNE5ORNmToEah5h1ccLKnORYo19Z2W5Ao0xj2
pkDKYgPym/gPSpAA/pWjThB8sbriIGlYeIgVkN0NX+qCgIjLw/Xyt4N8ZN4HUVRaywMKtWfIE294
eoXN4dUZMAXF6/6fYNwND0F8lAewnrhit99WvzEF6GEAmG79GkLPLjn7kG4M/i/4txghnSfe/Gvj
6/U0VmGAW9t47WRrBUCH83iYb9XWeCr4Va4wLqdACZs/TL+0OwOdgfbfFAXjYdYoDfQbQOlbH3ZJ
XYrLvVWZaYdVzCVb5KREHMao8yWJBLJ27FXt2K+W7RLchmcWHB9QdcpppUdEfGA/seZvaRW0+pFl
3tDQs77+5I7PiIw1VZ+IDBP4/+gkNk+OsNoF/FWzb13xte/0xv6gvcd0rr5s/nYNscjE5N8O7zK4
nA64Hcqk2JuXN5cROxfV7vE6xvhOpXGvq5qk+yxiPyUMN7fsfQaUKr/+Cksixifcsfd7hlUGAd+r
RV649mDoyYxtYKO/b1CJUhX5eA4asvGCE+Tv/gen4k59wPyP+fY7Go5QqrEjrSLuwMtN9plD6ENd
rimg1084zTeRyp6nnAZK/FIn7c6GHJZ24XSlEhB3e2Jt9YmFJ6wgAQp+ZY9eG4ZmRT+hcsf2Qr4P
86jRRGCBTcr37Oe5CMVNdnRd4YsjwHTl95DuLD0W1Xeun5McpSrTggpcMlEeLmEKadxaU8mEmwU5
qLtQkWiKrKFM7/e8s44bEcwQ0WhvTjKZwJUBiCuuNErmpnaKVQXMzQ0z8n3AIUEEe8lfl2TP/xbD
LgF00w2kOhssxzvVwmaun4iKHT5FfGQ/JBhKcaH3yFu1hhCKN8qzc9YYnaE/dAq6YQN2PTzNIc4w
oF+yhQYAy0u2i1x6ZtxTpD4aeb0oshE6rDKc22zPPvcmANcYzkTdaoleYMDdcJ0CgnIHi6R4s8g3
vp2yxVdOCrx+FM3gM5nL3vjXZzWx7Obo3a5zhEazgLt8jcH8nH7fhpBEBPbPeSMM2hI16O3ixN3g
iT9M7vXNyUI9gIqichSSQphGlGxst22j6nugCj5fSIDm+2acqm2bSGo5wnMsFkEnQ0y6sbsnL6GD
rXLtq29XDQHIOEiK6znsvJz9TNBIN14IuhhG58lBkzFj3w5NAaHzSUv9X8zG6b5fDDyhI+yG78lX
1AivCuLdSowOODPKICWjja/NZ2+K4h300iIqnsvJhSdF2iXm2HdATj854sN2J2wUWmiHzQUeuTUy
Yth/MFPbtM44AzTvAm0r0vep5Gw1j4ifo1nRKzYeX93At+pUg6lTBkM0kigBrCgfhsQTX+pEcmor
mSTeBg2dl/dpR8vjYftnCtVsZJSaSm/eP8UHqwrp+7Dm+OayCAxG/OmaxTPmJyQQxaRiFhz+y1yd
Dsi/Z1WEsvjOwEn90GS2RAD9xv0uA3CghoBVfAGQ7mkepgynr9JZACyJe3FGwxuORIEKXFLWOGW9
KSFk/2Jgmgj4s1lgWrp7nYDd0LRF+JqZdM99h5u2AWHw3IIZTUm7qwm6HkGkmGPV8HPzWbZ8j4iC
3MYYI6HDH9G+xJVtXR2OFfswj2M4hcx1qgDVg3bj/pUho0NP9c/ZfhMzgG7tckNxxj15vqW9zP7P
0ExfBx5WvjPimc71ah5wnxm5dr/eaBnI6CaOw1wNiWjfJKol2M4OnlS8WnUYzUUd67lEHejXG+NP
dc26m91sfn0LepGGnwfZ9EWghTxL0hscZqP5nd03MZl9QS2AS/7CJ2ap9LqAZycyJuprWdNnEn+w
/S1Iy4vZpC5KMKXYXZyT8SmB5EBZVIxMu7CJwhMzMXZfKOYk94nXlUi9bn7spoDHu6wh2xjqe8yD
yX1X6fyoNBewrkPMlGr+VyyCYa4AaxpYeoiDZYjqIW5HaG7tGlzW01Tn8AOinNuwAtV29FHKpsi4
eBYivEegDeEbx2gjCKAP+OP++U2Qysjraz89rlqyWhCcMa1Hl5eq5bL+pOYlmZfy5os3mARjOmwh
AhkDOHTHX8hb+XZg/rectKNkaIPNX97a6c139CN+kkHlgZi7wigLfRPKh3I52zwrD0i+wM4V2aYD
yAQdIlJ18HfEem9zlwSQ3mFwy5sWJGVZdPnnU+v7Bv+w0AGUUwgH3OM7JG+IWkF5yqmneclBMnW+
OUdb6cvPjeADDXUWWLnUMHw13PO2fJxDYiuYPV457phtqNHvlAcguSSzoJFEnfswT7cmHdFsyPsf
8M/GRrmtbqkJMtyqjd31mGbrs3kapKHGGcMu3ek9dtyWRbTp/181uOX8hYb0tl38KuVWvmKqzJ1Y
IJ+GGbhUWsuEZjj99ee7MPYEe0vzTZnM/FIpV289CGAdNvvk1YFOZ/LgA+LbQwJu1EdLvphcW1Sx
UTe4canA+LCQ4AxMQVLWn845xoXuq0pmFTcaG/QdrVSsquXeL+jUKtFJIomMN8P9ufmuLWs5m3gi
08BpVEdt0tR7Zbj/c9pKMdMMdPyz+DzyMGbIKo914mIw0Xyl4yYSHbpBLjYNbdT6J9o6H/54GMHj
72Lrw8B4EnjIBUfFB/oMXqzxBWa1lTGlVIdTrA/9IVOKEZ7rUm4xuaeOsbL806ns1R71O6KbkEXj
QWLyvi3QlF+K0LUg6gpImXaRSCFb4fl1OGOnfWFOPQJWjIGg4YhD6Fcl24B1KcEpsZ2qkBhLwZ2z
0CfCroyQVBVSeEcIN5JMi9NduamotYb+MWvIyoN2QQ9elC8fwHd5bWiBOCFUlX6cflglhomSrZAL
soVupsOy99WVHN9Pf70F4ZMH782WLkbdn5HISf6hn3Vrrr3D8DM5KmY+Kxj8YW6RIN/vZt01YgdZ
CmS5KmcFRW6g70aTcHGUEvOsW6FSvo29gGdmP3Vrcgt/7Y/utFUkBRbO3205nTSDFb4toy4m2JTW
Uv41b3t6prUcV2beKlQxHUqeM7IDtE8OD3Zic3yBUrGwd9x4gXalLV/E0gzHVvOv3V7q99ej1/Sf
MhDrXhmm7s7adxhlAKdiw/eZ95A4QszLnGlE1EiHx1jTJhaatUkJA7VImd9Wp2GgIibKOYrv4XGA
Mwx5vH4JCKjaPTBwGg32x8Um4SCjxVI0efVEKsxMtZLio+InBuPguFO2srDhOhXAiaIdv+o5w40r
j2idZrk2AO7Y7KvuQyuSJuZmQtrUiiM/naHTbUjk01MG4YXjYGrz8CBksEMltNpXak0nqE/kRQLi
LFlgSDRvne6nXSkoWVedEaBkbP/qUDxl/8x+rs7ipvcd7DvCbB/6ok6k/GEXPHwv8NELpj2dIKEL
Pw0nSE7eoYm8cyEN3dFRthtKBjzV8HfnBeWXRIQEMKfz/WJaH/AbjD+FuaaxLk834mI8x8yBHCbN
B53EAeKK6kvfL8UzC+1yqHVHgBUAmzqGm2PAkED+qoFyyEf8A6j33qn2kCVgGl60LWLKnkjCCnKI
NMHisXl+HGMM/NSQN7iOVrkQoGDL5KZnlmoyklAezUrlSF6BiVNLPt0cfMpEsgSHPGH3CeX85GDW
MBRIrHi1fduAhE4H7syq3GaWbFx/ZD081L9D+rk67uvaUTKafM90YFVE5Ngy/Prb7G/8QYAcdz+2
YE5pNwqRk1g8Fv1E211e4LC/L5SH4MhXvcp5Q8id1/ltqlwfULoY5MrBiwmDxftawzoSCaPqciWY
TjKvxYXg3FVZxQB9vNZbX48qZSzqdS5tVLht1eq0K6/5m7yRDK7yw1+Jfo7GczQOB4a71/eUA9xw
PCMZtJCmZ1BwcEe7Mus4a2FhURdbhw5Se32SHUVoOV55enf+Pj1Rx0wzXuWEi4VRccOL9iP1/om4
kD2lfQHSwNsDN+W1nvTEpf+VV3pVGHfLEOLR/gP9fHyZDFs9JKPsiDf4+0MWBw+7OF9Er+76ltgB
5Pk83WTiSBRE03Y2hgZWQhu1yBUemvFI2/cL72FETbDJx++j5L7CXYNIFChzBbVlO1mRhshNDTS3
QBAqsm427AyL5YZ54EQi8Hc6/6dEKdXM0YRiaXowIvSBQfom3A/S3clyn9+xwZz2thhYIrbXcrDj
PH765AO1J24SltuS+dm4emNc2+KxPJg9GFPwjgvSMz7B+0scjO4PSikFxtZ4k2Kk9t09ctd0sZ19
d3BFNgCbbr/611cAc9wQdkEulYsrqyEXsg4edziwnZbVZHviO5H/aS555lvuHjMwLgKqmf0DZXTA
zNHk9oSZL0z1rOd29fKPQxvXZlf9EqNbWDK2vY0ExvYJFRoLHBvwK/5G2gi11x5E3mXINXE1ls/g
trCjUe3ZUEsepEELFGpwvPj6zZ/mbEffJnc1RaCRtEAI+OVliRac73OZETk980Tdc++nCBgJT7dp
t76H31VMwuxcxgqV4kPaIo/ZMCxV/SbV0royAmcY2mdl3aTjtO7F2H73BGwb9g8+i4DqtwV3ajrV
dr6PiXs23q0DkwFoW5RR2SQDKSnZDvFMzbkLydwQK92rh4hWAsqID/FIQipZAEfnu9KpHfQAXi3L
hJKNT60UpsEiQ56jug3uRjftNgrqZ1skHyp5ZnplRtYY942cJhpAiqQ+5IMGrB+bJFoAOHPpjN2O
/QwvWTqENocFWThlPa1gzs2DlzdjjzzTfHli+MVHIoyPEhkvZtuwndwb2yXPf/euh/GDUZ7FVo9t
yCkKpa3SRlwxqiynjOCRyUevXBpw0ML0hF2D1wlttZvUjw/AMas0Ow8gckAf+gRJtVmgXGrTfaFL
BFmV6jSuCVcJndtiF70NvqFPWYo1x8LLrKqkwfrXzSjfzMEkEF6ijwzCa0Tzp/yupOAditG14BSB
CB25u5KGrJeZcQR0GpWF0/zFIOc746HTS5gDkPn/FCtBfDh8gX93/3sNxnq+v7z0MBpq8od+1Pkn
7CQEvYXKkn0NKroHUNML3/HnphFvyEgOZz7MBxwuLcnJbABf8SQuJnGwo4RPPu2Vo1AHMxr/a94W
rcqPZELRiCZJOPk5/N8K92ogGhj1J4RXSvcl/OAIz+2/25l/u58ReqUBf2R1UqGg0pHiMoPH6NV5
xQUv+PQ8DDCfLRHchDyJUsfZ8ThgOaRAmnJHQ3YmgAgYMCgC2flj3m0FvaiVsjfmzEVEpcoxzpb7
n0kiOq94IOElD6ttKH9j55HI8bkGgTagYkE+uy43NQ/gmGpc2AGhLp3+7jdSPn9uuggJmSqhh+k8
6mqrGoZpMzC/nLXcxDrJHcO0WHwRd1M80+XXmiHB5Rz9A6uvouxFyHhg2UPTIgrK+hQtpwoN/N38
LnLk70nN6f2YBp7+Tav2DU/jSX81fWDXg9cYlTlllhPKZ4gHojHjcHHD/TceIeQ5Od8qxHxjdRsW
TsTOHqyDayEbN61sSh8i8Mv3wYKu2Z+JxsogPNooRi3LBI6Hv8AjhpvZviWLa393oVAqVGt5Pde/
I8l/vqy2yB4VFd+HVEQo1my+0RRTeSBik6BRIZiiwBM94Da/5by4kX0nbXckqhiZ3gVfEneZ3v26
MNf/90o8x7P9Ko4t7rJLe43LlhNOiA7ysWaXG7KSmdJVRlivKBQ9eX9nnaUSljhJozi2VBM+2v1X
QdaiYkJgJWDsSb5i6mAYdxajjNK7NPoCklNiyZaNiNzWA1knaCTV+IizfajAL/vY00Maxg3oWwbm
iaWhMKofbqVbybRcX2RjYdtBgj+YiMnnWWb6Glk4xccTSG+owoS/k4+VCs0YKLNEuMaV3P7RaQii
K6AIw/aIwerniGvbSD/Z9KYJvwTxBqmGBaQawew4WIvh31NALPHzsztc5Dg7Cc/90FE22URN4cG7
AQ+aJ4JlwxTZA7Qci0ogMCy6L8L1dGJDNfbf/kLcwGdJrKse1Z4WXIBjr6swsOsD3C19E6nPR6KX
23fUhAHIUvvHa2uOF13MsQgZbTBvg1sciPTOaP8/bmaQsJP3dWpKc9e1BGUDXcGzr52U/FDnkLHW
FQY++NBCtuHi5KJFFTJUj+AyjsXul5OIsbOUAls1wXSLMbBoTpR2cDzussjBtlEt5QGaZ3yVJCOg
7d5+emRtE/cCot6Dirwqq3xQJ3a0DzeL34J+TH9qZOfeccFD2lr04outaTMyEHfYGAD0cEQrfrRW
di8AZO9nM596zA9nHFBR22C71HALn2E7KB47RrV7SDaR3d/1YF4jriqk0PcXG3PjLD+75OnDvLL0
f1r8ZyanrZ7zsY91b4KiDfkztnMk+mZ9xGefKwY48NbGqqXUeoUpg0JqoYmhalJwjYaKBjsHdtap
lA+WmX7IEe2lHnr1bzY7DH/mFx00U0e7UOunNMCgFViwVzkdZNc1xjR2VvPwkPMcr5ZTMgeNkqlD
yG8+zXSz6gprYekvUd0GwdxIYLwSwPjm9LQ+vZApwtR4aoSXbRzcUCbfMqDlghb+eOseYpyA4RaY
EkNqfflvkhoK7ewx1On13rxp/FNC+YxeKOUe1Ufh6ylZpAZAA0wva9sTjfcK1vFRIawvShyVvSvb
Iv25gpy88mCdU20HPrKgbLJHV975ojfTVi7Ymbzi41uk8IvkrzDVhe3kPKXObiOnOtb2pNJceNEP
CvdT1+3AaCor4hr5nV+0SG4Bty7urOGVKtxVOcnM32kkMeQj7z7AF2GDwom7JvbTZVK2DyZ0etuo
HlemelFyxhKNiFkSJw9YTKTBC3XBDvfGxkzC7oH8rE5G5Mb++reSklkIlxTOxP8do0gaqErCOa4W
ZW4eCHsfTF9aCMsqGnAJSZqK9HzMz9WTCfCixkg3dVEcwhfnXBEeZut70yYw8VZ7n1fy/sphaWXt
xOyRFFYVRQkkQz+twk4FbDrLCGIzkm4SuVZNNErm2gcujPoNenV6YrgLYm5iUvMoLb5yAJzsNjXW
XL5lZ8v8zUthepndhBRkSNL3zPTv3VVFet36NwrufX9Os+dofWleuN8JK/liHz5G81eLZuIbVMDL
ocTYoSZ+zNbHhZ/JPaXEAfPBYf/8djM+NZWqW/UKwmwO5eBgKadcVKzdqgBfVuH9jZf++dE5OdxL
xNJlE2croI0ddRTkC07ZMTKpX6DiTSe1hd/Ma9xl1OUB0toK2Luj0T2zLe+V0oRVG2z2NCuJY8AT
z63N4HrYtfQv/9/HxBp28VKYfVjUs/7nqr/Cz+7mpqFzLlZr9J+jFN9UvO9FgPftibICmVClizhZ
HQhKhnVZVqqRMbEffymA1XmI3Vxf/j6SGde4m9mDK2CKXmbLcu3qo8l/Ynqs1+z6vf5B0d68itTp
U818Dl9rLW74hSaHI04wN1V/E5C1d3br0hAzaccAzRKRsRYE2JLIvzCkz60E5998rXT09ikHrAAG
3g8LPsgqGHZYmGaEeBVmq75wdo7lcKC7sNiKZpKgGfzB2e2aJ1vhqjn4htVAh7eO7uxPJla0A7NX
79kLO0zWDN7fRd7iWiZbM0YHMa6g4Gv4KX+msk3fpGJXs/G1FupBHd0h7krCrix5H95+A/o6rxKu
GekxPmT4jX7/kqcRUGJta0IgklXP2sab+/DzuD0FCoXXBlP59wqcy31o7RlkrVnvAAxcBbycRSbX
6L/8lDGf1iifW2Vc1wcSfJHIeP8UxvpAOyxTUWZUWjNsBISlXtkoU3Q/s+J5loSfwdY8QtAsT9Cp
9L+Y0cV2DyDO6zKnZzr0gMlPQ/gNQKPnMGxWRAhlgcoQAxnxDDiFlaN86ueonZLi/BiMMfZMDQ9N
A7DHAsaeRYHmhAel0og7EW4spIfpC4FQFIkw/i8uS+2LG0lOLtOy17RQozGnsQ5SeaP2kwrzsYaj
6zKfb8aR/qaJeOYqaQXBXaJp+K0NTTa8MnfRqxI4EnyE2y6c5rpcIenE1uRgfoOwlqV+Sg15Q6Xt
in9P4CmFgqSq4ioH26x7sZ7VzAAEt/tY6jC42SN4frLWiMY7pH4r7uIIDLHU39RwfUJKzIwioVY3
tz4NHl73Djcfzxhk5n+CNE2eWJsXPhhTOglwcY4XL4M2ZU2HvXDA7MtRjb0nmsVdnI7RKZ+IwYBE
A1fPjja4iY0WfHJsB6ClT9S/b4MtktD4koZJO9cc9CqlhCOZxI1GlCCnbannugycs74H+L+5XVFF
FqKGQNKid80iUUWdmXNrHJrvZtZb38kYvOFwMW2izDJfcHNClwKNUtRykcCkeduVZv24umCbNo0Q
exQsT6YW5iHl+S6S7NTnCbwN2nZOyXYI3V6ae80fu5/FkVhkl4/WL2uPdQMsaArxssycewWzks2Q
AP5Qherfx6tj7JD1yOxMx57C1vq8ODo9nNrDRuh6BzDNIvCfpCk+E1lPxPKoL5ytJg4HgErY0t6/
XedfSIw83EdSAAYQu8fv4scZ1Vywu8Rtg5RZ598oEBfY9dthgcFfmeRWwbC0Q4deD7GdQ8YbLDA/
aSguZGUzJrdahAE8af+rVB8fPfgcsSBYJO+20EHUCTKB4dcXOr/2jHxvYVAj2LcEQ6jnaeaYxiLi
cJIbys8d4/PPSssnUr5YgPLLZLtzAqpo/4kbobTmr/jTHGJCNKCBgJx/SYlFd2cIZ2LtWzD/VzVf
akvlUGc0XQz4b1Up6LiUgbyQk9YJJee7DPqtqJOvA3d/MT02Zx5ccyYEw2rVOYV2CIrMa46pmJ1w
5eZrFEiUkfarV5bTWqML52Fvugd2r5Ml8Iv09p6Oiar71lbnkpmMq5X3nuxtYjiDgDRxJq6lYgvi
mKCIyRy8DrU6ol/lJ9CZ6gkPqh/8wnvqX9VAqqawKKTh5bMTqupR5e8dKWk6y3JKQRhRaZdTWKAK
1zJKpmUbbE7aOcnBNJu+nQTk9XhSZiOeFJQvpfLyja4bxQMyogTzaRsBZvJSpNBybZrOfFqMr9Ej
3soi1f3ayZIFbfxeqNP7tX2O6foxFhE82pgIXvqZRj/fk9YFWKNLDlIgklvaX2zyKDeM8E1hsiyf
P1v1d5LAshGzE/samGjlMgQC7X3nzMiqKxIgv1Eu4yXtMm0bob3FD5HDUdiFmeuVigDn5TWwNmwN
LWmEyy+Mp2MJ2VhdeeOiBg9E35IXWfw0B7zrYshykrkTncuAaQ7H78cGsbY3RgaKH06+Xi8GL2b8
26zAiNIcr+Q2xbi/QBpdBHntfHsSFQDfAhK9PjnrnjfY76ErEtLwS1Snw7V7LiBWSY+LnoVx89Xj
qqC6DWwOS9uGn2nZgibpWibOzdPQ2ZWvdVQqtkMdW0eUQZyb8HIJMRtw7pAbN29ibQNu+RzW+Qyj
B0LcogCwtBhPMtuf7qyOMCFTLDuJrG+plAL3qMEmXhvS9uW9qNybfg7PAjcW/2K3F/QhrAG8F0jI
9Nlv1OVU5zgbeIJwPzou2GT5tM27/PT59nTgVf4I2UqErXxlATnmuAK0PLtoUG1aa9oBfkg2cbVV
AJ0atRG7KO6a5UY35pqn0WEElRgPol7EVkL/+IW2zDkAiEuhPRy+OKEgLvcLdH5u9FTrsFORhDCB
941ZgfqQZ7X8nVEw8MKunB5odOcvh/fA8zlNpWopAb5AMkeDoipo4zl8Syohett2ioXB0gWbHhz5
90wlgpEjamBNtwyyth7IdfTxBsxDA/GB6nPWY2m8++b4MSEE8oYjueovOLQMzQgGgP9U+puixTwa
7Rwx3BWhAsSdPisRO4qDgO2s5HnmB7YO+OALtQmtKlbQKmgVCX8iBawMWOdt2WA/jfX6Ocf0U1Rn
x5BMCaZZNiZfiw3wrDNhp9NpBKFExktUscoQmwfO/ZceIvIVaZ+JM067mta+9YD+pjzS0wNxSqvZ
tPHLrDHhCVqE3FfCf9IjgCdUVuiMlWzWWHQ5977xYyn1s5NpttcJHWMFiGD+EVEhhCy8onyhwnRW
FvVgEcY4WbyhfpaDfGx5JuVebiX3RhRa2qjM3yRVGEPb7b5f/ITfBh8XIs8sckAYoYKIrgYZj0p9
mrYIaW9aIwQS9lf55QNhaKYVgx/9DMWB8vG7thSpn64xm3x+ctESorA3M4usXzm/3Df83S9eQmxh
ochzwibeRWY7bFRoeLQQ+XiANas2aBLIL/kQu/6WaMuUS4sRuXaNhuJYSvT0irUZHqPJA1oYbpZx
BrQPa0tOOCrjqcNZXkn75bcNTEIj0aZTIFESMB9+RfQLJwYyml+QWPdRT81xm85sbGX0Jmg9s/5a
oBsoLZUV2GeGIu9iU6J9l0/x1QqMMJgcHiRGa8INMra1yDSxo2s9M1dob4Ul+SXpiUbs5qSbQc1d
+qPtegc8TKga7myQxa5eugXxYAwEEBP9vknVTkmQUh1EiCM4g8yEuMGotoS3xXA25keRmlHiBJdI
fFWJm0nAZMThvHuSNnypCRBpNcRhWgJSyrblXubL+3han3D3KVZgdZiaCPZruew2FEymgLTAkF51
5EKPV4maWk14ERY8p+GUt7cKGhunn8NEHtUcDYx/qYWhnxj5mAmUi5/z360/aHtt2X127gZPhC1b
OVL1qmsTxNEzDP9JGTOi+mnwI7gYAJVSHhTIrjGBCtjgyz+5HkCk+LcApu5frx3GiDPu69FtkHJ2
Narty9Eezd52OfMYogFTZhtQ6z49hz4xdpzYekvtMFe8CkjPW2Cloo6yKnZm8G7tHZGT55KQEX+E
iq+8B+bm7F/jqgvdIk0aKjqMlIsAOoJd9TmbUUV98UxQ9BHljZ76X46w0swtoSJEVrxyOg4KYXjh
pG/wteM08Zb2HiFGQWysDIeufOtO9P02W7tYXfTr1mJNWTIxCqUg6UIG8dYl3TVg5Ilos0sLub9G
adJgmKFnLy/smWC8tRGE5NGvZem0UtM2bwJ+SrMKd3AiBpEyikZSg/ITuMFPz33joZ9e0s6umJza
Q78yOhy+kMsApQX3FgEVkaf4f/zPbrBv33U3361z7npBQwYGJ4y6I7Sk9f66drdgJiEIC3Zpdfkh
fyweoLA7l/VcGpHIVGgOEWieSGbnXu7cT5nhVTlEZG3CsOgLYnQsnxiLmxjjd3FIYObKS7HkOyoq
pKNNqrOh8z2B/AZkMrAdtsT/mY+pRBs5F6izI/P8XWgRL52Gg6HMmjc57eayWJSarVandCyEVPkw
bV6IheNgBUiNUigh1EOAIj2bfhOK4rM0gyfccr2nSY0Lu9ciP0EePMthqONea+oreOkD5UepwQ+5
FgUYiJBa3WYtCEFM+e5pyu2yQ2Ratc9+MTs9+p/2MN0JxL+EJVAKXBwvEPm17XKp99DI1PZAKTZ0
7UWLo9kZdHKoXN8UtE22JA3Par5ZghL5e28naoRcquZ0VfdVRptwUF/TotD/zat4obhItukspQ5E
vRuTDQpqM0ftNsY8yCtUYMefwf/S9fbzeXmUVkQDn2GNo8CwKr7K3wmNeMiMqDs/ZkHOMCadccj9
zN/c501ptLhQ0mjfayV885xnjiFFE5NEURNrsiZ6BArNaKu/qI6JWB1nJVcjPnyG9yOPhjaIaKlW
7WpXz6vVXHMTTncuH1cmSF5lAmY7vPD6Kb0eUNenJnudu161UxppBtlFvOrn6VeqEQ8Aejs4ZDtN
el41Q82Oe3AltIFeJyuCoeoaAknVQQfzYfx09PF1MzNdkp5peO1LLOnXO9PYydqqwz2UU9LThjBn
1ClYvMTCnD5tU138DS3umc3Y//5aprZqiqbGs0KYgiiLrK27d/D5Lv2j5/VBIWGaz+hcjPXQwaS5
nKut8va/AOuF50J3yIPrOiprhSs5/DNSKdyXaqjQ5GV1/TO0f9OUS/IAQiHpm211IOhB1tBwcuFK
QjF1wtVW4u1qYGDj6z7dJUIh/AcerSYBsu5+t/hakxmEMHEyC0yhh0MRiuKqsNshXzDKhTiWg4q7
rhnY9hFNes9w1wMclRqUn7vEIiow0drAH+TNBmFrntcBPrMoLzJTH9Py/w4Xfizsd+MMwJkwhz5e
cDYgE8j5JevZ2zsURuYosWyeWdiwVze2R4E+qmt00r/GDWwVWyVo0A1bb8v4y5FFx+VIQ16DKDBI
erDM23IxPKOTSV33FbfuhrBaDQVsTJRRZ62eLdDx0pttNOpQ1tYZVKeF2qj8ziLqNp055rB5pXjC
QTqccv0RmUDgzfYp++6qvOHiXzvkX4NhVtwO9Vqk3cll1THNgTIFJhJjRmeYmYdebxS8XAqMd7NS
MueoHFzTWFuFBQnc6ecXCcXpTbUlbryfdg2fFq3XBZvOZwnGlIKSExj8B6rvbtJNCv/EHGaLlfsj
gsXcHce4UNlLFmwNWJR0ItnJPHE179433KYlXT8QUdN18JCBJWe53lU3F37M7YGUxdJ7JHfHnRyJ
OXnVsrYojNMhd2PXaSW8E5ATLs88VUWxCWTlpBfEbcdOc1FvZNCL7YKR7xkuhOU2uXpclnjndGFP
8B42u3How3h3gkalw40hwlnW3w5CU0IKMevLvv5Zk97wiIxAbpYxUMVbPVxg34w4Jh+tAXDsj//G
TqOuzzUty/U++dagZC7Cdv53MR/6x0rcPTnWyy2F0ButvFhaPXnUt+gi/46WHzNRid6KU+L5LsHe
uIdIwYNkmYugVu5l2CYpha3r4Ke3ACTy4N26HK/Vp61e70HvygIAYPP8nnIA+A97JvCyyxk05n1v
4eXpinrw5kO+vShNeQ3jvoakXSkUiUg8WIkhaoFUQk3umqyQOhLI/7y6V9BvTHGRQSWYCCCbsxli
6zPgXt2qAanM6KcF79rUaSO0VVlSEuhJhv3uTQRx8eXt1DUkYWQocEHNziaz4vBQRtl6XljeoLEc
kaZhtZMOjLvhFOXNFLKYNhq6oO+9dsZXUrjeYH/cH9mmZp/ckUV5CeRAV2tEh18xkQn+dMGhbUu0
Tc68AFJzQK0rs8iTaVubVecBQD+0Yf9R4O1fDM/UZCxtFR+1S1dzSuTLc4ocxt+KrL00PO/UzlJA
5XmRmNHjNPt+H11/7FDYLWW8kknnbkKNrjzZx9nIdM+NtN9i3CLVJQ1AiDp3ZQHSOd7mKR2FzYhT
/QbM7hQc9vKs6/5Fh/s3rFF+k14IRC2uq88laiweELqZCUd0iPluJ3t/6AU4rUeFP5rKezpEEHYt
is0jucJBncEZeWZ9QWkHz0LE9iNrqg0YNdimrTBMvsC9YDon4TyP9rTuS7uLAOTm0xMxiJ688AiL
8KcNCjJx9YrCawxEFnVPwzUpEEabM8vx5KJiFmMJH7BEWQNXc0Cn7BZ9Ks8d86uqF8f/0kh/jWDo
lICJ9m4u18ZsQzU9gN+vAjfirrIKQIeJIs46i1OnSpLKvOENEQcxlhtr61JaaJOLfnEKf0PzQSB3
e0YI4agfgyNn32THp9E7m/5QaAv1KUSc/g24n0+K/3CmWs3OpOePiMU8CnoN+kzgTnj9xMO14Try
iSe9qJOioGLvChWCR9JEhEHMjtcJJPeES06HLHs5/4vh5YyFX6t/3u+Gvawms0OUtNGa8xkDz36K
QyDeag7Mg5yfqolpoJJj+e15bEHHyiBzAUC0VQd7082o7YgKMt/IWZk2jrcNgKDsg1EdOZjdxExs
Pz+hT9UXMERnH8maMZYz9koW2oon8nVLcszyPHlmqi2qn9VRqhGZmEIMXArFKAhz2Tg7M9W6J1PT
T3+ou4DXVPJSD9kTjjfH4/ZGRsMq3A2GD1n3fOk0DqysXMTTWwHUgm1mIoAa775xdm9OZ8HqmvjQ
77PbrDsZukCWRxk5iLWYX2ccGDCvFlnlvQkGUm+fgQzaD0kieYi1VcLML9kcufH+F8dENvPnKT/U
3QkDGQlABxwfAnapnQvKK5Hfhm2A6NFhQCz2JD2cuHNgUpaTqxN1D6NFioUtvAFMIsQG9r+ex6yO
eUgKDed8QUQcuF/TYsE26oup07PGQJubBXDzAY99kxN8VKkojTjbMKI2+983iYdfvqw2GEDQU59Q
SdrPF2nVgJK1gFyDrhafPuzdoWdiIepuNYdjaKZ4Y+xk/vvvFLmLizP46O7a0Icx4E+5KDlPzU7t
5cy/yqBEt2jb7jlfXC1B6lU6Pt9YtXYAbx+aULh/ZK2vP9B3FijjmKzBjRNB+TK0MABgQxX+Z6Ln
T2RNLlhk/9GlSmtMz0kI/gqfMaUxhhoeDkaRiHtTrUClkNDQFFqdk8TRll+NTTyZi8AId0YifKKR
CqmfZuzSA5a4qir22LBMqV1LCmJQNboaTJJf3hTVvEMGQAbTz/m1Z4E1nDzK0JaGJlgSPRfsNwyA
M7q62rpdsOiu9kSTjBecXjIakkpHanaxBvmOvubOW14AciE3UGY1POx0h1AUrTRKYxMnDJrqkFMi
wkMQ6RQRmP8daM9mrmJ9/ofIqVaa0rrhPik9crjwKOm/EN/n1aEWjTP7lnMltQlCW1GXdN03nJT2
BfydxrQcjvs6oBddxMtJILdgBjjiKbU6f8kPcABNzG1hm8KW8FeQQbVbw/A2fG6X9xhsexP5DBX1
zoK/1s5fMWDfRdOBQacLocMqzznjQuyhV6VqMXAqbMfQKtECy7OhsicZOQ+p890QG2628YcMh6op
PxKZz0fSF7eOgMaxVbR3Mi/3S8tHEIQIZK8mlsGKr3T9N1y9yI6hLpQBCifKTOWXZ7TNwBLrRLZM
OVCC0fl8Asrvq2KP4zVn4WynAIY9BPSrQB3PLr0SN4AQ5IEp0bPg9YlRK3wv+IzmxaMwM7FCPmui
loG+RZLLNB+FwJHC4TarilJ2ucM/9Nm0veTvqopviVqFb9WSNuQ+BOvKO+Z4XdKP4qZPk/7jfu/p
yI40KayR7XPkZDKUnxZtTMOQ9eD2+Cud21vff8Ib+6uPHXP4us5B8DnqaCNq+jkBd9O0aDyqw0ua
ryIABOm0Svm9Mq8EDmCtO2OzBa0WqgmJnhK0zg66HdcTl9Orir2LtKlWteJuVSnHoExsjD9Glqh3
WqlheLgv4q8oaWcrt49a3Nc5stYci/gW9MP7X8QSzvFoBntl4rAPNrdWE14fUxCjsFpaVYBJitrZ
vqAnkez5be1KixPhNg9DraGtXcXde/Em0IuW7xLGMBJd+HaLwErI9r9VX7b/0MqyofpVj16u0Czx
Nz4Tm8Wmv+2mKH0XeEO8T2tIWunaFl7G3kpmTyikJdGSGFc/7G/SJIJPwHTFHK3Sf5BJQvpGZ0ud
/I6h9eW20H/ep1QWVITFrs+UuFOVN2GmuY//GBb6WihSOJTxGyBfx2Tw6K3do7VTQJNhco3TK8WU
qjTxIjPZ6XiUAXXTD2Rhvcsq0MxEm/zxIH1zA3AOTjdlKFAlNf06KGarxe80G0akYGbs0/ldHEW3
iqoFY7VXZyDcdkbX1VWpaOjqUHF2hlZKkUfNUdhRSfiqh1h+nuPsdiXKG5PB0z6iUD5X8oLhwPUk
7A8vtCpquUyeKEVIWOPdbS4F2anZ6LCs7bAVV+b/QSUb8zwnFtocDXWauqtBeKnixmblJZdhRf+d
xuLN8EnUZt0oiiawtr2GWz9ST20GWh9MMFwztptJoZCHNDlj41Pz3mYQSzsRB/8ABIELGqRmdhOG
TTZygpzpgwHN/qESSU9/QxiqZIEdXnIf5j/754s5qegWJ1gB1NbWJLgMO8mQsNfB2U/8HZdB3oKB
vM+jVBArha5u+m1o+L65UErCxHSz+iO6V/2PydSNgQP5yVkBteSJ1Ms+hj5VXbZb8GNf4290sUVt
ARlb3w76RK4pXdiFOetYqn8tRn/wgKtwjakPC2oSdpYFOwtNLwpPwYZ3YYxnmTYrO49XoeM28MLz
iFMmIZGBaRMh0GxnAarWH+0qpaNjSKfGyyerZWmTxvO9Dc56A32/0hl1sifn1WIsqocck6gDa36O
uvR7KTCq9ourvMLswG7UJ+cakRf5OSuyAz+DioVUWgKYKOraAavYavakmLMfTd4qT1n92/QjVYpy
GpXAaPpqutagGKGjoWmiUUE2mwEDeqFwe0wENJbGhOjqIxXKxkjMFhHbaahCyDR+HiCfyvbXDIcB
TRfJUtMz3wp0J86u9cXLWz3pEPsy4GkyUrbvmRJyJzewG/RbuOYht3+ItfiarYjKhaJmI6SMjCTA
Orvp23SRq3PuAvU5ggg0gtCh5YmALdx8JHo+cEcMIaPziJqwK9fvk5QXae4Z/n9DWdNxdoO18Ctt
6Vb3m+A6xSNU5LnREjzXrPbQMZz2YUql/HMPq4UScnqeGHkymk0Vnj3/dIAcubNXuhq4ihPjvZAh
yrBltfdKX/0nK+40ll+zPASQKryPaFJecl1RqxNlJ1sfPYmtyYmgS/Z9dzklxaVTY5VR00kl3uB/
XKWjWxIfiC5rEGmbZg7MrgqKBaK9C9k4mWRTeKU/CS9WXZHRNXGoTpSmwXl6W8mtmekbU4/Y6CGC
vJ0kEFY+NBDDHpNdfP/ExeTkO8CYlE1tK2P4IrHPbx97BxJG7zta7TVzBq1/3M0ndzYLP5gCVWN/
q99QeW+Y+tOnmTDjgSVBjb5oEvqlT6ATva0Tck+b5h+qqXwwHSJrtb9w7F/1qjjjgJmqyDsrAyAu
WUZzwF1PvOlYMBkOYu0oTkGFc8Cv16CnqmeIgRaNeeeatBa2Zkv8uv8ADDBCaeyOvvVgAaAijyCM
two4Esh7+O8K9+ySEBkZlP2DZ+Y+ti2qjXPKxqYUbmhVcjigx0Uywpw20mrgCCwteSb1ApNYwCIc
nXAqxYs7wZscqneueygiCvd4OxTkrtZOmYoJoPOo/4Kc5eqk7rNQyslM7ZHVIMixGb7aARvr2tx3
zyYm9W4QB4eYkGf07DHHI7HfMRw47mU4ClqDjyWUCgsvlTefVw+GeF28t8C76KVD0aJwbdqGc1FC
GgB7rcEKe67tuC6aNbYZfbo+tKt6umfH9ldtRq6dN81dNIVrxq3Mc72wkEKUr4KCyXjCfvOV/oLF
pb3uNsRpM1mT9wUL3WWPwKxVY7n8qBdzxVvIYu2S9ruGHXtAndCUG9pCHgBIpCSxYu3OFoeogpVO
CEgZxw7sTN9d+nkCrcqpBGYe/qapVbXwv27poWpifDDhEiLi68+3v5L/a3G3I03zkZNoQPvWxBfj
TJ+xprVpFkE4ePpCf+K65GCqkksCFC62/6OviLbBBlocyrOqEebLEXKb/LzfGLjVpstgtrwopPV+
w8dEpFAd4Cq41u9BBZtBxOLEWnwetBJCI78VubmOkGSsWlDyz4gPrEGUPVvB2k05LTXxtbzCzWfp
QKeQdP1aDL1XPEJEsLwhRFlIm0h9iwxAXfn//KkD03Clq4vJwguT/PppW9gocYXpHkETnO45x94x
UIAMVZC9oX7WataYalCd7RurWrMCzBD7AbBIZQFX56S7Tv44kk2vi35i+PP/6EPZYbl2dwtEbSib
+Zt0LsgSVfIU+8sjY8nJtrqpr8jEaulDIu4TcA6bzqkP6MEg/GhDu6thUFtIHGIrHUrf+3LDZVEj
cSZ8tVLDOJmcr4KR4B7S0SGUOc3drlR+G5CFQqqACJdnv6E0TAgJheSnsD7EbzPUAjRLx+iafAra
Ee7M2ktxGgtPYjRYb/ors/oBh1HzsfYJRqvf3g/xSLrt/7Q7cODnpV5PkMOCGxrro3rbQRwT1MPb
fEBn0UQPimnrEQz297I/t4lRXQR/YDHyJTk9uBxD7hffk9gmojoqKFyvb5fnW1DFvXsL97Jn7kFJ
qLu8/4PfZjcslfWzZivC42DNMUt5T7GOE+57GO6L2JEeUOkjKlVFNlEj09Tp4yz8EvQyriNbCLZP
qSn1An0oUxZeqDz2OtBLELZ5pYZ+2T/kVmGofe60HJkw0nUhhfmTY9Wd4VI+8cYLs7lmzbQAzEbn
doRvfmhnIredrH7+TYhsxgrHOYMX+S1aW1TN6YIZTjnk8aRXwhgkKltE+0r8eaFYXaQeRiomM6S+
0wQk7nacIxWrkAMkQCrq6MgxOEiT52cG8MQLc2Hok1Z/8SkXQ6d1/4s7v5Wy4897a2w2eVdhF4Mb
7/gFcuF4E6LvE2X5gw1qTo//GyLJ6ao5cq6glC2ACG4R+lEyz9Ap3k5uBlvOuKbjC1QAVHrBE0fn
xmz2YHlwVY8onSJpEFgFFUogbpXG4EKKupVkz+I1Qzq5/pzDf984DAO0bJUAVnB/Z7MKl2hBn8Bc
JLtgcKZj9l7PpHkjfcbykJVKejaFMApCy7eTQAMUBoFfsKcG1+5/RTasxmXq2FfeylQKpZe/nHfN
BifcASiKI0g886/Mlq0CJ/2TR1tycF6nsfNbBT/P1xx7hCK8ykXsDEF+uQZmxwkNPrrL4SOWe2cY
9f8GgNm+11W9Jg9zHOEsuTEWUndQPqhwQ4cAw8o5QiLXYLkwmKfwenseVnTrqf8QrwklnBpVloXQ
qrgQZlLaGxla10ZXgQ6eY+tmB2dj72y5O4N+jiFkcQFBmXwLUMpXkQQ6lyTW2TdisXNdObja7CcN
3iczYyt4KVVkaFTED77nYum+fSDewj6A6mDJcXZN92svCWETBD3Gb2C7d0AqjCyfly5/mRelRVOj
esb/L8TcP7RzBv3TaOgq47Dx3D51+WGRyIoX+GzOSVB8m4SibGsd98vao6RbB01jRIb/mjedVjiF
d6/GG9y4YEJoBLPn4HorAVGSI8KQPThkFJjHJRbOIYE3yf/2cxXLd4JEPnxMiVKmC1UDJNMzH0Bo
9RzGqwufpxW+dwEkojeQ+ZaxO6TjeNAJmH3YQi5AxeoL2w/gIRA0PwqtY+VYeLAOmg4lbXd9TRys
Y21YtQcTU7sSwWJNOEQWtdj6geoMX1YL0OFMcbXUwXMs4lawEtnuN/x4vyEB+Fv4oQv+clI1ssHX
hc6a3DOlqAfqCvzhQPHCHwn1oq3BzkjzmFwh5pXpk8PzpoMW2XxmmMl06LzyViYCITctNPPL6L4S
KmRZP6aY+ZEdlHS01ka9Xl99sDQeVjor907Ndv0Z1DQkuH5qAx0tTOA0tuCWG1zPhhYwMMc+Gn6a
BLNOov2736q81NFzUUhM+CACE/PUgDZH7WiX2zjHiM1Y2AWRWkGHG4/SjRnsokS2ZgOy/IbGcNzl
2HTjkjuf1EIug3hGWR66lMVOkS8uUNEPfx+Z2fBSFVxTnUG8FMqi6Q4BwNeaV0tFjhMqgWKZhb6f
zTgFjaKQz+l/hnM3PkP9ypv4+9+545CcgXhvGqIUChnMK0DoJdurR2jUjFncIzhfpCBKOreSMXXv
Z6iCGGY4DEjd+MrdhbPa3AyR3vqeCo2bIG/nmoLjo6yyZMmeJ6+MOYAQuNwifqbPPRC9rcEc8PjB
0DHT/FpQ1CtTTBwC5eUkdj3cFWppB4KFQ5hP4y8NNSN3GM4XDf9IBbthh/ti7Kam4jonE/ntKkbz
Hu9cUmcwgyuZwld1Ttv10u44D22ZVTZSjKmK8K/8JfxuZuJ5r7N7+lKB3FEpXhhWmFmYolTjDQgt
h4nmeBRM37vohdIVw8YZ0Pvmgdsh7cmniZMlO5J0Idd0Wr/UqF/S1l5WDX3eJM4dSlQBTx9a9p9R
OT8WGeIx96A8xpiHdxByNPfh14F5nCVb8+xyoL0WeUIyaQKpIhz3yu5Lb5TgzMXEiY1Z+bcKF9fZ
Pyxg7aT4GflgKmb8hpS0YGXJYMh2ALcjZ1bRg3gYjflk0Tah7c/hDLQ8BZkcdJlz7Yf4ofxRCqBJ
JHkuDX+JH4cSznU3xyA/gOe+P9GOhahdL72aApdS76j0zeJiwY8JJd4GLtFAfUIQKHawZprUwbv3
WQjKCxzn1ZxzypxRrl7MSVirG0vhxYJ/UMI/Vp8JYvy+j/AO0JaHEIOJZw7S4snmCYWD4VhHbb4L
1By3YWnQR9Z+7uvNEAheNua4CTu2CXf4atts/64EXylm8zPV/GnXm1m5PkpEQPDcozTFC6Rnp/Uu
gX4U0mJzPKW811AT5eD0TWtKzGB0TetBHH2WUuBfJB5aN3oIs4UTj5p23osBkkQlb0fZ5auaNHpG
+fAJmHplUeKrmWJ+82v45qEa6jvJ4rJtJrGDQGmnRYF0CuatuqtSCZuNVL0WYqjj5h2BQSPybjso
FGA/SnFPcWjdP61tHgib9uJzoYl70V86Z4S1FXj68wOab+garecNmCM6CJyqELYOxAot+JNKigTg
1RN3DHM5X7D+FvFHYvH1RKE5Q51X4O710ermLV5y364xyZNNZLudajV5mjBRjZDXlTyS27SrsVbr
NQ91CMFLyDF9EYos6lVXNjPVocLXLKhGTu383y6suG0lL18vvGBba4L1edeoYpmKz8LE/OR9+GAr
JCJpBbGjCndYMdwe+KWDSh+UCj4f7rLyPmAebGzJReBCgGdk6COQrwxEhhm1pCkG6cuFH9xFRVkZ
FQ/Awg6F0q7pnhwVM+LX3QXc5fQS0NYXLSgEfBPwyCdRGaeVoxDOoywdQi5/GcLdB0wvEnw3qRkN
P+2YLN6UGoZf+x0rT58O3yzOn2XdVCgGRQA2Oow+i95VzoflL9q4ch1+luo/MAwUEdl78FqJbPkv
p9cjGkmu6w26idkWvK08A9Y6DAZDlST5Z3lh0ieRqHaOPxNqhXA3NbRTqfR2JKFT2r1vtJ0xsHB/
/2Ef+uNkW0T1oUAz5rn2MNAYadgQtsdusmh8lY7R8OCy54fmME7vJJY5EJnpJ+cLNJZqDh6RYZvi
dTohwPP8Y2Pk5GA4c1+5ufNrkJyvOMJrvYZoXVQvMuEdRhukDunc0TNIrmXiqrOheRvKMB+pKufM
Vy7tjtlifyn5gs2TpwH37U+cRQVj9iWEqWLpLTGzIISJCT/JxKye9HE1CAMg0o1A9+9I6WX897Jh
QB4s+qAARNdnssrYY0gGVbE0GYhLNgAbrG6iyHrXhwM+HQS43tB74+bVBsOw0qJOKbTEz0Hvmiry
rwh8iYCXwswV0UUSVgblDSXv71toz7EuHrXS+eSxeB57XFLSdxX8snW9UFnDgueaRjLtySsxpB8t
0PXANH1uMuCKO7vpQ56AYaS2K/mwmQhRROeJflS0FoP3NMxAq2x2zXDBjQBWjn4bdUwcCKTirDt+
JuWo0Prs0gv90a+ef2d0+oO/HDoXwYl2Duf+cpU1qx6Q80q/Jf6vZN37lXplqsxQQsEAfFWexJXb
aVAamUSKaImWRvv77hMlsnmCNwypZLzc6MmaC7SU7IJDw80IvnCSElWmIOrZdwaicsDUimBw0pxr
hIaOrAfLDDgEjFVaG8MKkKw4HlDguwDvRnb3hdshWhuLGKIhIJNYk6YC4evis+v1v38xvK6H8aPh
lrJvoAX2fzDswJrry6IiiwI4AwF3qonIXjydJa1AIZwAD0UAzVpGkCdCczOgxp7GwwzW9wH1H+H6
8/Rsa4vh7Ccb3KLn79z5toLQdiiNcwa/Mdorce/R3MiY7SN7dnrRuQD+n/UszpqnRwnsKquED553
iAwIPOlramglWVaBt66s6j0FHc8ZFjEdkETkIyTJ1QYcELsjuubYF2xg/0oqCOcyweGDJy4PdPxd
1QQVl/OW2Z+fmSVi8HOmWTyVNnGW8a4s/FlPdjrruGwElZMsGsGGGW6Q4cWatBC1LTnEcB5mOIiB
S7imQ+r8KzwrYTDPMP/etZtKvMk3SIayxvjdUpLNEMDW8hb06p5TksZhEZC7UjgD1CDY9bUXOtEA
AdpKNJxGNlDZrvsS2CWEv04NtLVxrKF+lVyaR28OGVCxVeKDrRp/E6gczAA7Z+Hp524LJy55gEyP
i5/jmtQQ1jwidTsrIxdnLe/qE1F0dpSXr3XUeVmqxPdzTDqDiSfsxmwOyRKEhU3RcgtjjBZFkLsq
TndEkEGeYNdTWiGTd6Du0Goij/roXyNV0rsVp3gWJmEy1GrdvLZpv0LuQrl/hj44xRmv+TdS63KV
vbCTRBinSH7oeF2/u3CHoZTD0upgMGMRn59VeBY5MI1KVqqqpCNRpvdV/k6k6RFILzYmFF1LfgBG
E/txV/UnVhFBz2HU+DytEaLauKJEecIO27zaufxpmcbeI7fpo4SF41ElY4ZMFaJQvdhFuVW11rWn
5ugxKy4KfLxM6sU1ty+XtU/Q1EZ0Us/8sabw4FUeFQ2r2wUobKcDgDN1YatznLF/3/vYPYaNDyLW
w1xdjikkwn/Bhhfk59rAbbPTJoCQjS5bKloSNSQMP2OYU8gPfV15mtB1nQ6DR98Hqff1KMoIr6ha
/ggq85d2rTPRF9JzgieSBdhUt1GsYe41G8btTm0LPtfC2n+TnuYHFlPyaIWheRjIg/HpW4VqDjky
NeesNefiq8k+HKO/TbJAdvvBY3O9IdDXcoojZVr03UDpcpm8mMHy046E4DboKaYzz1kKi89SsKDF
wiW5lhd2NEGA2YHlS9+yvYEgp6JB9/dsRDi09ig3Z+IIt5EXhzdgEa8/RuXeB2878QrcgyM6NhCO
BZq3yg6NkgYRXc4z9t+LMF/ohQdB2ytrAqn+4fV1jZUFTRbkWnEHC35lQZqk35v8Y6PIs/wyl5Kd
5Ntip0qUmEifi4soswYeMikYA/NNMUoFW1lcVkXYaESk5n8oGLup3qNXFWRK2dDB3cY75+AaDcA/
6rbdIvrQ7OaOk/YvrnlpV4OTQsZjLol7w1bZt5JMhyywnxt/cARzQESvrtmeeD+KWS+GZbJIntdr
n/mVmrnoGw8oE2fm1IU2T9V80XDw9SZT80saiRdT4fQX+IoVxOkkrKWCMMD4+0ekkovy7XjR1mdH
kfnv6+Em4FbpJNCTUjw3sr/0rvHxbG0khbZChjK/rR4aJ+v3EaUdOA/fe9fbZf2ZDR+juI4pVnIV
Zjrwjh8AXME7F0q8Z6y+hVahH3u0l3NJizA2LIf6PE1RyCjBxUXZbtv19yhFK/0VQcHjSJePKc3c
ErDQooHIA40J18pF0kVVE93CMOPsyqregeuX3qSnLbD8EUWf+otfCbOrmSVYct1/LJrX+mDWR6rY
WD14pUNpIWSus550LFhVRaHpWYEIiacjq1r9UThLZhxhGNNC9aZrgAYNSSAE/96vSC65kTTiPRqz
kMAhx7p23jVKM6B3z+2FBFxLTN+xOTTBiLlr+bJ4kgj7Q3Q35fu5I+WdxDtdVnT61PAgQGLhY4S3
N6frZv88YACQN+hM/HcJNO8x7v+Hq6BVZ2Ig2g113viWkUOZS9uGJi84/80gqqveVX3zupbSS4gu
U3MQ7W0SmEz2z2DpaPD9agDHaMs5aL+OiD0uzIDKCk6S/mlQOEt0bcSGSmZYuNA4rmr8GyYMi2xv
+xMD6u8lc8azxA1mRQ0h4dFE4dY7OxRjc/c9M1MReNOU97jGRHrNS8u2AFeGABbDyvZfsgGXQzA+
kTYXdcRDSxb/q4/I5jFCP1nNWXzA4xbi/k8HVQ0ohAfaHhUgE2OAAtxQwt7aOpTe8wqXc9eeclR3
LgR1wZn3MK/6wLs/KsLc4+tAKj8zzw7DFxxIJNG+q43np9jdcVBcVpS9Hejgf/CX9JLxDrSLE1HZ
idRMQWdvyhGaH+cpACxFb1E0kvkzNTdDUVZK+K4mRWLyln+gadH4iJQtqBDqWobl5w27vqEd+TEH
CJ3/7dfcl1Dl21jIqJ6bNTFq0WMS7A8kWDxLYh9zQOKunuY0Dy8m1mK86YsvSpXMZivwOmEq+y8R
haXGd6XAxTE+bl/cRwnrLguR25PnHtLaBeGYePuEazH7e9cQRh8UBtuM1uAHnReS4g/7IfhBoi1u
2UgkH3AntvMh66iCQq/2KQXq5KBKQjZss/LFY31imPRCDpAcRiqAR+E7M/fQm1WkffxtKFfGH8V6
L+gNCpWi0SVh7WJ6p8wanNVQqrSgMmkWn55WbwHevav3U2dRNou7fidl2XIBRUQEzvF1fkdrDHlp
rw0HO0WOhIsE9dOjpn5How0RtuJJwK3DztdnrUFMH5Fs5Hu7r6T8q4YGaGoGmkB1LIdlr54ccpe4
M3I6pQug0Czlh2RZAxfTKETN+9yRg0Y2XJAzMVgr3GL8UwpteTNC9f9r2qBbn0RL6cO+MXq5il9F
z8u/6u54wZj8mci6kSWef953SbPanUWX2RCrYSYm01xnw3K+SG/ljXp1xR345qGx166mSvEoiQQW
ZvFeiMbxZWPg7XgPSjKb410wS8gd0PIRhTPZ45Nw+Oi5adipLDyqXAARhgHtg08ogMYL0GvNDcYQ
JFwuBFmgXLyqF5wRNqIpy+U7IiIYvimc/rP64w3IexplAVmt60/nsYMt8MTpP+SGJ5lJjiO9Kbu9
lbxPLzEkSJPULwKoyb652eFeBTjezpuwIoIwZ4zn6Ru8XOB6cW/abKbQwZq7vpwGLzqkbv9mXYGw
gPUtIaJuq4zHx9Q8C1HknAd6W5PYQif7IlGYDj3bGK/OCa4Hoe1b15ZDmJ/5dm8RtZYsDSFPv4d0
arkZI8j557hUO98tlfh3eR4tFPwZ/R5N+xFfHovymJFDnsJSBTl9vr9XNkaxA1dibHz26t/4osI1
iBZEZJB3PDzc3AvhaeRIq7WU5gKXCfQZgKu+7v5TId1fLPd2jMi29vXZOyO+9zdVoI5dfG8LnYU4
rCS/B2bgpWSzIm8hQK6G+xGpFFPiu/wnROM2sYs2R3RQu2kx9hN7UwoDO8ar4S1RusqmLn3WJee0
BkYs28fpaVnACTlLoiinyq3HBeFm+3AtMAco9XANkEToamwexTTfDuu0SAjZ/SFTgyCNK2il1PHH
BywalCfaCIynX6dLHZ5UozDkeGo+c9GnSNdO0r58aqaWap/c9FNVOZ8cVRC+bWN5+Ftk8REI8kpk
ohPpKVpuUUPLCbJbs/5nnxft68I9Rz6Tl2saZEDv1bxjBlE4GvFNFOa/iCbFw61IPF8YAvvEMpNe
Lax1GL+UptJUsI/n071VRe0iCcPP4Hyx4+fxO5bFgK6COdDcrQbgl72ps2VCfu2jBMIbjaUjpR7r
k89ESWpWNB2aZglCa9+Kj0sN5Ld8pQ+SmPre5iLaGPamkwSXB3NhvJGyT6XOD6R6VHU7CuwWu13x
Tb+3ZOyl510dvPPJUmaWAvLCtYH7CXBLYfuQktHoWcue3QUhkT29Jy8VhRztmPhHn3e6vlcGGH8W
XeL3h71fHAH56d2OsHzXYzcnQl/SaKqHrQrEbg+4NrhNbGNG1krHaJBhCvYUl0nhMVwQ4GkGY3Kf
ciZQQnw55p4lF96pB5MEeMIsOZuTQtRPP9D5J95VBn0Abc1uP3alZlCgiimf5mTmhG6UXyquX8sL
GcEEeEOrHGOzGtGEAvfPH5lrCltf7LDOzcM6K0+n8P1Hvdjxds99SiNEw8vfore7xLqbAJ+eaNyX
ZXbjGUW/kyoeIvyBIYI0WWGj+uYm8HKAO++NNc8Si0tiLvh/JWRg8eT9ioGRnCnKGwWz5fR5/Yiu
f9zzvhYY6P2EBpOzDzOlV79XDrzkXjEuVTsAFyC7Vz3OFV6fnazJDbs3vsC1oPtEbqjtv1XBbShK
RdQ7ShCnjpfsI/w6gLjUBH5umiSEgiyw6Gf7iK+s9LrunLQ4v0ojXEl28egqH/DycxQlHoboSCXu
b7LdSSaum7avo1TbSqvSmCqHfIa44y4hEfR3XDYVZCTSHweczaUeB5qi0z8LxeH2wVBF4vdvDbDk
Fmw6YS2rbpf0RmgsgIVEytGlgvg44n9OCNmiYfTcN5C1LgkFh/R11XAXyxEesttegud30m1oD/UX
k6f5g/wbBcHtyLsu/FQmfPFR/D03Vpgr+TMyxZ5H7jCDIHpEXhbiwdVl6ev2aNtzNAOKstpUQlUc
eyiwWLrXHik0DBYH9X7gzV7X2IyHabmQBf4AnfcVh0Y7rn5hnvnT6H3hC4IvGm1+ZIuNutlStst1
ZlAgYcDyHMmb1cvuB3PVM7SC4dtdN6FRZi6sTfxiM8tPq1d/4uAHFbFBFnmMtafTBray/CBG5xCw
Q7FBcnsPsCyS+InFgEp2dSzSB1xuXmB/KYuZ0qHhB91DjJYMV5DQqco7AmxZBi1KihV8FfF2mTNX
BzdIyjSl4ekN7MvyUQlN/MO1gpnZNtH8XihyIx0I+IjTnq0kBD2THwxMKy5XZnnapVRo2wku27tg
qlivsNyUgvugnyPbhKxgxycBhI0qLS2DQdRaObkaNbs5vwCIvzflSTKtn7u0HQb49RW9eXvfBGcR
TTCq5gRD3RaD+jR2c76cjBmN+BURNiiQ12TevsznZG/JdhdLW4Hi82Wf0bKAKmdkM21qWZ/GrbxQ
n3TEexpiqfgX1lNmvEBqlhPx9yCSNM+f5v2f0rWXAFYtgGi29nOZiT5b+BK+BgK8zpFNX4Ef2Mbn
wtROh58hw+BNPgf6dkxeLGAPIo3wodqncfHIlfYFO9S+29WWCQlvw5e1nggEasJ1PF9A+flkyJ/A
tL+3VSOvfNAeEtzTlyaryyfZTfFeeiAD+nRYmdQ/vH8sawSyT2dLOzvZmBw1Uaepa8eMA2MxrG75
CvM6hRhw+GnIMoIz/zjGq02a66DVUgQXqKpDGajAEWcMM/EtrN3cnbkoXPCNRot8X9/dX7XY9+w6
K5iRPrT1tgNYPZ9ZqFDCf8CdZ/t9drbNzuOFTtwQGGdTHCxAHtzopGIsXK/RxozixJzAiNmH7cNZ
6B0uG8u5wDc8HLTogskvGOtD7RRaoXbBPpdZdr/bU0PN6zDrj5j/o0/CZSiBzD1JTPS+RXgY8qxj
fb35aIqUcIgwmwSppb/1ikupHReNl3a1cRvWEHj5rd5/hmhana6UPfdIWYbtU3BpE3xUlft4vD1Y
8BJbdEY39oUJIemrj8CSA6SWFTT1QE8/hb6j272NN/C6wzN94U/uxS+m9vghVcSeMOoNqYREXBEv
0UL2SOoAYgKK8r87xQk+sdQpIa75OwSLp9Qcs6YDQnXX/wnKGMLP5RFpZZyPviVPPvyNCCZlPrwz
XiR8pGA5gXBdvx2K/ilO1Gsbz/NT8ChwkwhVSYqb08s+2yQyJo0cmCCR1pt2FYNt2UWLwuIuxKXT
qNIBYJhbb6UmHKOXjOZLrax0ZXqCIcACJ/ob+Vb8lVAL2GkocR7EzEV8mH4T9AToxnAemKzRbKFv
2Fpw/rCzqK3SOapTWttqCA+Puwfw9xADxwLvKDKYr2wxJ6sWN6xBlipiwWIbe/ipT28IfkOFOq9x
XE9ut30m5EksDQoXd1cDtVmsrrPjXduOChJuObWQi/ijd4sRvmHZv+khyIzvvFIOxVZZ0+ib1l8X
gSfQ13/6dQQiZsSW/nCbOLFlFCIwpPCsK66zR+xVrKnzvVTq1iGVprjAZtaHFi/G78zXd13+ns0G
H+l94CFbTRUpGkhHoWfmPRfbRpJdHhV+BY3UKJIm52fX+yAOzAn7wtqTVCOeKP+pF1mt+7gfmWSc
zCFjaieTCwJW7ERGiHExhNZPpe3TYEU4SavgdL03Xj2yUKCUHhjuqMNmpXKz3PUop+V9HLRq9O9N
LpDeahu30lGlZ3sWfo9rrBw6owecMYE6NM8MMbstgAwSn5J8vI8aaKwCh4gejXT9Fqb41rRogUoO
oE5lw+vNs8wwU4m9nBjpxzOomlzPWtOzOGJhApjPHWfB0Olu0xJky171EHXs9v8wPIpf9RO/d2ky
AArFyOazMK/ePYox0rXespl0V+OeKSq2gxFWR5zpLix1GDnx1jQAbWi5xi8ilwLzj/5NaS4/yJeY
Yo3QScg6X9FMvBxQvC2zafEb1sojSjBsmD97JuJEkxa2oy2Sqp1JGAcCEehX4xoW+6n6zux9Lskw
Xvx4PFJAGvhSUMwhiyw3ML2kPJeEZQfPJfV4FkHNARBIkkn7vDx5KMgZyd/MENLZQ4fSUeKOH2bg
ihkyC0SfOh0hFe8uviSzThiqLsNGgFXtArC6AzxRD7FK8tjnpVO/W1IXYR6LVrPfInB6QmHk0V/S
ml4ldwf7EzJoUF29hkJ3krTlRRsRLrS8VfF1EUM55beMcqxRcV2XGBF7xPHVme4OCmYUYfWE4pwi
9dYLdmILHQO3RI+Keecr8FRK/GXmfnNVpcv54LisFQGmFcicbQVnM2J8sPfyuuTw3/HdWTxqbOro
+NHV/wpzlc7RqQPE5gRYxDEJ8elrwyPL8TptmDpdm7vEL6c5H9SwicNfJCHpZRIKc4ozwjvkYND8
wfSSMltZCc7Ms1rHcGmuvfxacrIfj3p3TJyWg2qcg7WlBnixMtAKwHHYsXKhQhKAWg6Ef54UFBkv
xf95+XudqB96601JuyVXzQEXaW4zRAclrUu1DfOArU3lFSU0DjbONLoOFdF1JQGgunHGL4SjOsm3
s5RxaEHombuqY7oUoFfgjsUksHI0sAt+Gs+FgLYSH85p514nyNPnf0mcUBvaar3vZOcmRYn+GRjt
9LS6H/sy3Ihkn1ib9kgcN8wvn150iyFbUqkiY0zTRxUBhNJZS9DiaMMMm7khGJ6u8fw37fPJdBnb
eiA867chKaDCJEqs5priIIfp4ICDfSxbhGMly2L+FSa+c4KDoG0YS49nPRxtzO8wqrwJ9MEbkJ31
udKHTkDUOorW8QfmVBBmhW7rNojQbtK6KXCSELss+v9qAdUaOyKhIuljB/vWrR3qDqEvYDcmSiYf
+aHJuDdjsDCiYYnU+EsTrL08yZfFvwtaobjsvAmJj2GkcNFbKdmJDyy1pXpO73tuJHAzX+q79Z7d
H8RkQLfvwb1jF9KtXCcEIYBUavufj9rynUCJ8mrirl9EmC3YWmzXK7q3B5Qq4h8yNDriQg2xbcep
9R4YrT6lV5sWMPmxLg8mOwK0c8n6pPHg9KFr13zN1MXPrHtJVrVJl/dgxdctLGGtGaSojiL3TOTx
oQ0y4mwFZXkNgUwgRrgcWhu9xpeZBVWWe+dJLAjv7/5z01kuLjI1uzQrg4o/l9OuG+HVUSGKOKaO
6quriJWM15IY6lMBN8c09CfwPYyUvcBlAX2m5O/Y0dNCgLVq9/bwMAgLSj9TKxriwNnUZYC2bWtX
kgEKCjnz/I3ftuLYtQZ0unddCbLP52wWISeReaX1ly0DYfQiCuS+Ua8xju7pTwb0oQKfruZCzMMe
Wxp6ssXX6IYOBI8VbJe8F1xrwFr+c1Q6WiAV6DiIiX4WP3LR5MDwQp7h6YGqCFoZUG+L5/XRduzo
Bp0wyAbzIe0IYRCi8MHmp8n3nIoSzzAPQ4uk6o36KkZVwS0+NdG5Q+AJvjbcbNVmHxzCPApY85fw
BmeW668iM/UYCHUr6HAacyjbHhNkqfAIlmfiPTjFViNjdlwtirPWqQq4MKRpDd3cHybcmf0fQwro
lq3Ua/SJUUS+HmAvg77ps6HDNreeCmR74AXKs7FxIP7k2+Ep7MKFcSAKwzgHJSJIQPnO2NOW0KZu
RJssLdrNZ/CCJH2/jJMH8OugZh7D6ShtrDlFAKE3RxPdAeP7a8VKVeBkVH/1ie66ZaTRexawiU/O
5+M+RfMrB8TgcyboNsYuhzeeM0NUyDgcGuOtCTyJGDfHilvfARq7XZQVWG+Rbqvsefp/VSnAWq0s
WlMMQmq3npsaQ2zrFLDobPYXiqwJwqnGjthCjzAI2e0xAEDU5R+2qQn2k9rACdpq3HeztoxUlyiy
brZnd5VoZc8dxrS+s992Y3gB59zJ9Hviy1rKLVRvEfLIQ/m5ZgVm57wjJu8ybWcbL8r90Na9MRWY
3wm5cFGIC36vcn91euLtqc1alvX1Lsand3ovAEY6buB/8LvfKQ/GmWrK+3cm0f7g5cY+Uk+zIf/T
Y986UCo1mejm0xIEnGkyk+2rbQzkas9qJ/MsbZcYPhRjL4IIJrgyDP/XCL8z/DDGX+gC+Yx+//Uk
eR/HebQ5Uocx/qz4FYQwLdJ7fbPMAbzXANGmK+am153jMsdCudErLT9eCDfRlpbeULYBefMXRn/D
TzlB5ix5IkpN89qgaa5nPALLlWb+yrsCftlQL8EC5myIvaAo2Svlz15tKtdG43rLT1gEFxoN+590
7Uz8SxklUg/MvO1ZQ79oWYCKLUbVCyruWwhYq8kLqQPmbFbcKw3a82cX5nEpDSkOr7n5O51luKJ+
FoU32JcRGaWArt8RY6aNQTLIifv6vmk4LbSBpORaaprhjFJb1ps8kfkg/Hmgw0D01nmtyBroKPk6
gOtDGLD+nvRh5khTzM6BiFJwvjasl4vp0HN7dS69kLp+rUGoMDVu7DLDOulJlojp1R7pqFBMqOX9
y+XMpKh3E9Cq7xdDGzO0qdwLQRaGOraYRDMq4t3u3Xxh6ejmpsTQuEmatYnbC6RU/Wb+nhEv1OlH
ov712YG/OOime5VptLJ4xgnnECpOI9XI6TrnPjl66AhVskFwpx5hTLsqRfWth1pqc/K2Qssr2fcU
oboud4s7WkaDzI2EOOrq4JmZVJCOHRqZHk9E8EBkmjgOftezjLnSeiK4HLswtOpwaCh59LrcDnSX
MCQgBZ/+8hwvZhTzy/IbszpbQ/H13bv3H0kbt9azp8y1sHXVxHT5n8m6GQJQ2LgooWd5Jt9qn4m0
ffHVrG+pk065i7NoEkRElCA5YS8bbqaFt1P6dNSGTK7tMafq6wTpMD44Z40puR55a4VyoxpOZNDh
at9CWo2s8jmHACm86P7w8d4urSpxrg95kNAIzkhGj006jAY3W6iLOnGPRYfjfouE9eDYb8Hk1DNy
5lxxBQ6DHuj1DGBNOMghcvXYOuJyGepInrz/mB+IUFCNFkLeLaqCksfuHPxC7YTsdT4d7odO8bcZ
vgI6jIqNmWd5r0NywaVoQjPcbnc2zOmkwGNqbvJBj4GzO7PdtRZbHUtQRj5ZSBO1dEMNs36tAz2Z
NJf0wU/SeBEWyHLPgQAabV6dVKtNkyENKE8qrHUDz74x0NvvXyjg4KHKSeuWe80emtAztTJQXhwH
8IwT3QDExEFALGyP0vkKuGVoa9n80nrnBlAOHcOgbgyUr4z50a1l77hLaVtortL+3dU6k+CBhadj
xJLrDVyAu8nSfB+p4yBE97kcaj2CZ4+xwogqj9UlcYJb/d1xvNp722lZOxZ0JWaWVOQl8cH0Btcj
5d8UGudL9xuh4J8hpJ3U5wPtXekTMcU5C44b7Vv+bJfeSmYr5m7rncfQ3W0t+v2F3tqR/rtGgdkr
oBnQg7hh7Nmrar+UJCnxkx6RTbMWq5b0qQfBbq3rnEGDxHiLdaazDNOmj/LTQDzloqKY25tmIv00
9lYF6Qe7Wg8UvZtv9Z/WJqY73EAO7ZsTt6mZUKHUm8bQmx4JJLX+Sj6TPt+1jTB3DoGecDBi46a5
dJdMV6h8/J7E9w47pJCSvdzLctBbX5V7SjYb5qSfQnc83J1eFhli2kk1dWEnCKUovaAB9WAhr/Mo
K85yVpq3YGZWoLD0bSqVMDGxy5gX9s1soAKVT7/NuF7pqS6lhji5wt3e/+p3eV4HwmloQW+D+PXr
EqMocuiS4xJcmq8HSTJERRKIb+epBb3ud52rj5jNYFZIz87G/6UGjXOM++1PGt8eKVEkVw1z6Vs0
mDt1H6Db7DjFPGKqu3TGtPd7dD0rYIoafsAtymahBfxWcNHkHCWH9eWcL0oJjLCL2QF1QvFQZ5jz
YC4ZVDB4lHEIcfM8YO1sO7USGTMPnVTbuLQaz4ljGdEoJMmuA+p2hMaBbibWSgJADyDqspxfia7V
RKeLAu6bQIQMZNpbe6EjauyO1YVKb6vkcCSD6EDzGlnsdUbbFaJJJDjVnXS1LfYrASotOmRXYlQ/
o9dhbs/4Ym1MyTA8KeLXV/OTzQ4dLXV037zyBhTyhKgaygblrO2QdX8Gc7S3MkjMtgy3uu820nvd
egePo4RQUHC+VvDlch+mO+zPVgNBiWxn2T4502fLHAMtUlgA0N3/AdwB87MP45KJikM5p7m61MYR
lksHzE5zOF5JFsX/2ZrZ0WBbwY4epjoXc7Rx0iSjuR6rIbA311VzZAlOP7p7IpUIOQgrhRGOaqY4
QUFlyhoseYzD2942a4MZnFw/pSFDY5VxsLAEmYYnHnFwOXx6MLmIo4ziwQZ/x9gxOqQ+tHzLr+l4
Ht8MwHrdnJC9V+3XKs8TIMYrGFjTA2xl73BnwSp4Kujh9ktXonBo1W9gjbzvKyDKlSPQqY0fY4+s
qTZ7orUY5nSc4YEuserv1tW8eZ2fcKJswJmi91GupdxM84IaQ9sZmMkc8Whpr2sSsdOvc3RPsU6C
jnArs+r3mQT5P+3RsNVUXgpFNLpmKlOjc3KzPELQlDmid8yTdIZboftEY+NY3vGpB2IC6n6oJT2O
I6G6EjWduI/9xCWF3pJgFPezc2aZpaQ3NZfoiEn2lD+ojHPi6m6bLEGFyVvJaWvLaQRHH+rrmO6Z
gcy62VhpBmKVjFEt5kSow1Yaq43Rioh8IE+qFjXsc+OjgO6Tdl+RwpntYcYrTmLDCA5qk6IU72Z0
8YsJJibNWHt/IxpArExXGubcoLaynia9s6YUZ13ii4vW5GXVKCh6gnaYqXLHJeCe5YLswh3hNFSI
yfQFxPxbPR6Ltv8TTQRIY1DFot3gRhZocodawXLG3w9b+nA5v5fMDrivaGhVFxktaKOWRlQoG3tP
jJ5WPoGEgqH4Jr6A5amhdDPyUXQVcwoLwnc6prpIELNvDT/cuv1oQfUoSNd3QJ1cAZXhuY0FHTyy
2aQVQUZSxTjzOPY78zhFsz3534AutRS2zlQ6Vil+0HS1XxHJGTtXYijAgRjSi7hMo17966ZyTfPg
wuZhDZqm840ebs9jY1r4GNA8AdZPSR6ldi724z2GE4gOTE0mLXr+CGKBABD8bHKmAB8uzzBfBWfZ
NY+dH5Z+QMlxXWl4CoquU1QE1B5ESILfur1LSqWRINiONn5peMNIwhfKOLPQCRJItePjuxGH1gas
paWPP9PU8p9VJPi8gWtJm8uKp3NG5m/GdKgfwAoJIRWIA11yRXIGq9chYoss6cNJ4ks37JPRb6Kl
audIZD9+0Ct8u5wSWjdyFMT6MPciFUI38dKEu1mD6CxelYEpfmrjWTBawf2GvnPGsRJamksH7VQB
KEPWNEKVcpAAp5T20rAgjbfeNHKu502WUzDOC7YYGkyIFpPw1e2lgwotDHI3F0gKUQs9dH3doEJH
JQWe/Y29qkDUnD9yg+5ms24tgPsOICFcsuRFqFoT3V8sHqYE8UDVRo7kyiZ6lnYURfhCIHJRGOic
PgrYOHOj1qCW0eAzFu89OCAoAiz+RCGkjQxfRusFFZDRMBtVNACrhkv8XSmtp+ENRVY3BrlTtaYO
97+ZnFjixrZnzS5FUwYKK8eawsDpR8z1iMMhFLKtJ+eArYgaz1itme/40SI5yWhrcuV909jOw/YL
rhLWykf04xKaOIeZyVrWi0DsND6gpADg98uDBpDGygt371yxe/KEAUXKPva+5FiFvqP96AQiT12x
dLx0APIz66i9Jp0O8GqnwO27r6r0BEur/XGLLYPJTWWi2So5DidaQjFyXEHe6kNCBRGyZM6iHVWD
jABbTQXLXp9GVmiHyM35UgIWER2+c60/229VfsD7l9s3gg5ZQpFeccYl20X4t3BDJZrmDpyH+weC
utC/C0NJNbulH7fkaXoBYpbCtVU4WaVbGxHK0rSQqMXoXwhciyV9E2xYh9L1ocN6WJjIYhOmgfh1
3WnxqqN38ZqkfTw5mOOGKgTCe/9MiPLD2wV1xGObDsZzt8PIJaKRwxqfI2FWxT1+Dvld/3mwqn5q
dQO6/qp7KVNESusT/NPIoPRQagjMU5uIF1OYDHyYravHsOihzLgTRYPWg/IcsYhr3LRiG5O7Lwrn
wbAltaLWRRCb6cuh958Rh/1vMAMeKS0KhMefltIV/gAVApiEgez7bNq5ztsDlj4tvQXmaBPIZ6fu
2E50KW34Hgw319lt+tFqM6XGjR/qi/KPjMMY1mhURAhduhCq31M/9ygly8vhhoWUJjivQOUgYE0A
ek7Faujssdkvb5SHuf1ZTiw7w+zDDXGIko1ficZbMHcIhQb+JROd054FPMJRh3/CxpbK1AGb0oy6
7fKq1kqHJ9R6WYmCSyL55TAJnBhOmNVOTCpK38VVkHBi4LwA5gYyxDV4PVYMAiO9tuKQiJ2vpJ7U
ZCqIsU4YUNFfLfF7p1AxGUxMODtTEBIl1oCrLzVekP5VL8gEh3fQ7tehsrq2FsRMZwlgMfJnLhHj
Ooe+yRSMVNkqdJ47lps5p06jDp8BSdbf44DXSfycIvJEewP5X0C1kQML+roHAasFDVoziZGFWxQx
FGwtpEkQLgRV37IYZG+KjfoSOxppUZjN6M9zVn5v+jPJ5L2ifMDh3gLkLtcAS+jW2+INpXgphZqP
aFDB2ueq012wJZ+3zFF34S6hnuYq24S69rLQQkA8vWYWHRc7aeaIVV+1cOM3JGzKOFKrVELsfL16
4BCYabqZlXWUJ1muBGR+u4I7IXsnrwVDVV0ir4T+dOXjq4Z6noPwgzafvYvCtKa5v6ws2Vc69aOb
lzFvJNOcDCH2ig+iJc4LQDnlR2+8+xgEPhKKSrH5kt1ToBGLHL43IwJwaqtTAwQfyo2tvA+s5fqf
g1WxosVPejUtJ0KHYa9rmjzX7iDcecxvJaKiSyzwadGnTdOfgjl59KyC8QDTU1ndagkvy9RP7hOz
84hCUoPRN4nwIZ+RHRGPvYgcGni587bpJc4QrZkXZt8Gw/22C5YbUa03BtfmNsoSxrwyVzLXZoFD
nS8t/G96hnVZo/IhgJCEVsUV5AC2OCxc2MWeS1VgPLJjkFLUle16vUfKC1OzodmhPu4u8mibIwkX
xJ9G/2M2jCKreLmp1KRq23a+dH86iS6Uafi9+BgXOm5uv1gipyBpxhlod0uPZ5I/xxUsji6YkAOy
+Kakzks6eM7/QHw4kGVMoe5F4eMsc0bSQ8UimyN9UYQhHWg6Phms2AKitykOxcnKoE5i3ZzxpgBV
cLrTMvp5iJcvQiAb4RZlMeQ1a1S7rSmzOUTFGt8qYX54Kkgjz4ce/LGJUtEQFcKo1ECHTmMuL6d6
EHOCQnDL0RiKcmy1K/B5Vn4QRmu8bDK1nFoWaG8dlCXYtV2Ad4w3i3Y1fXFA068ieWZ3j0v2uSn6
GFOMcjFCHHlXqxtZ/Jwdywz5Uz+GPfcv/yUMRj2WZr6lHaiXgVJdPGJPZTEctGX2wa0HIXoOLgPg
Z+ZdOyPGfUIUxhOwXbSmJqMPMpH4FAzxCBjZ2vswzbcR10luFNy4GQ6g2jyBqaGESkEBbm8D2c8s
qs1QAWzT3AKxbsgeVpXsUTKCi1EeGi8WgC35KDTB05I2L/U/VQgQwpGvV24Bu3FZcr/ZbJWNKRX6
OqPwRYymW5MB8cYpQ7hbX7ZBcETpeX+dbMKUabNdo5bFucq9bvttnPB70n76P6DHZs7390p7GDQ1
dREE9pnqpqQqQFTiuBSE6DJVOQ8obEB2XHte1mFtZK0GuDridqHWxdbjaVjMHGs7cb7SOgi2jti7
I3J2waRbgsxGBd7ZXfe0QALxxUR5xNrfBCAURbFYZO8Th7aNkcIgEk+93okdloyvFOgtqh7XgXdw
lZNmRE0KM0dPUUQwcVf+s+KIS0l5RZkW20YW0ULF8T+FYNWVFrkWck05NZ11YiHI7ZRUOKEoSC5y
3hFSm5rbUcjL0CWiu1F6SpwROmBRMBH6+k5ni2PY8fuZewHiwyqarkCHDW24/x73EkcWZnMvHIF+
hGbUJ7w49GAa8I/Zqg0jnzJEFW5wiP5eVfRiVeY1PetcwtSx8J8OfcimqxduTanSyyqbfOfBqU5M
rv3H/XxrP2Wz11qKw6jWZjrGHtJtKQK3PW8uqeN3FHHWZKEDmdvv3dzPnPTlppLgLoJnL/EVim+F
b7i1k5rimVgiJTCq8Dm4GE8fRAlRxh/Srz9A5nxEPpxnXsHxOaAMPkGpIuaZrh2aQshZwnkjJBv8
NWGIH3nwf9ZnTIAwvcUwpzmsOR6f/rkDxlRAjq//+76VfCl8KQKL8nTXkDgeEsWuQDG8OiUTLLWk
O4D+g6Z44f8RJAOnauYuyWXBperEOjXv6mP2dAe8i0Gfmrr8aAhDGsewAejTYMDgSsRz8FpP5DeH
etIhhUhG0mibwhPUYNVp4FgKnyqQ2o4DObzuuEfIMZU7tz1VjA/J4aeKPpI8cb236uonWabJ7OMG
d6tY7DPGpQYP3zrmP3RwoElwPTHz5WBlVq1eO3RQpp48aKL4caHXHADj/WenNSaf0XNgc//Zv1Q4
qSSj0ns6CQGKxCXCNs2W0U12N/TNmwuBsdBGtN+AyRdidmPN0SV22KSszo+pPJomuYqMqfFNMOgD
0RFlNMDXj3+XwJvNjXsRdwD8knjhRkSze4jn9oc6+bfWEDM4Nc+sjNgxFEE77qSwMxQAIwH26+yQ
NjhSzJ58yo4Hg2QJlcdbJzUaptOfLDPLVDTHIsLr+XZgkA70dYJrxTsIlwlgIBUyMB4tsBcXNfVZ
I6SvnbltS+wcnrsq42DRBaZNSblsWaYYyt2OoAPATUvRh9HGzL+7Sr28V3EoG7HP/ms3akS4KuH8
neDbq4k0zREQ+GMNL8Dq58usBnp8Gl3z1buoB8e3rQiaN6f2A7oND1SiXRux/pgEV7elH9E8ygef
AlAglNsFx9VufuswyfVtaVl8s94iZjVQiWvjI13Dqi4Nl7gWX3ce58M3otzrsMkZSdsPSJskMT3G
pyoOeBc0Vl2f8EBv46X2ubwBBHNCtAZ+kk8HiCPw+XWkzsmU/XuV6zaDYSh70K0dEidpzHvw2Dru
rykU6HVuYX/T/e7J8fU8t6hn7T09BFQzkZQ/cRvFcECDmbtOWkq/0+xyhJogF/m0nr35CjvcXS8s
yep64Fgf9SNB6sn5G3fMBYSvdcQcIHx5F4I8lbVExx/wbizv+I6rmxQYj4SsABXDKIiKbg53hkGZ
j5yYKR2lDDYwR1B+/mF8I8/bCwpvaZqTGaFJrzoiHRW6g/KFvXujTyeN2mQKOvAEzFxOkMJDyJ04
p9IFDKDP9nwvxDLhMB5CnOZ39g7emY+ey4A9OertifTSyEES0ZIN+BJybS4K0HcAI0EixbzmsB6q
1WbmUeOeVvwvA3CnjSvQHMw8o5LBTWaWR5P+4uPlsNTJB1sRpyzPTzN6XciIXnrPscG1uNOZmgY0
MddQian1PNVdWwZcIkk1vaILMmx8NpMUb09NudTTJkyYnVJ0MNdNnd1F55WUPfuFB3JG6PcnOo6c
SbHckH1HnvHS3zkCC2UVrG37N7G3gyhgU837G5cMo9xUcRo2Kc1jRK5BurHHfP7qb8x0ayPPPpQC
QDX/nD6ZJIzojxRGZztnOAEaPa1JQfeKDLwYPEjtLaM38dSWvtIirmKloUi/Oz+TImmAjb3HEC96
1mHTGcnA+LXxmoCivCdiqFvqeK/9mjKpyCLjhk8o52o4RKXEkLtC+vEtDAPjUyLgyBju32Hdx9wC
ciwysYWcJE4hvdxjshZjlu+Qs6Xqa844K9N0L0Y9QN5NvkfprYHLNGNBA/USTnbGAE1QDsmWDi2R
S+d1R/eEMXCiP7JFBX9Au2aMXaFNFHpH3Cswz8bnsvKQqGTMxDnDpnyadB6T97Ou9PvxnmB6ImKr
OnwwDoSAHe8XJC2xVWuOXcncG38RJwCTVmos2cS05D2/0h2/02UlaekiJc2+G4qM3Nb6WmnlhMX0
Um3tNJ4MuRtobLHjfmNQM3sqyfaFggLihH3BH278e7RTU7f1iD96aBABNt270d+V+8BbP+Gtl+Yt
rNOsLKUpC/ENM8WW09FF0NIPP/8tlRHaKqkCT2xz7ohCii3toxwibJt1fcdtH+ymaUjom47KTCf8
yy3PfLPdIZSKHdqk3d3DQn8bbQxm8iO7/m9nOMhdYeX5e/QJAXOARSlAKbS83ffauSMpXM/e1Gbs
3a3nPXwQGnBemacjqEz1bNFMJhBx7toIiTx4D0mnvtz1i/42NJSUaighmgDxUX7TCuchTZv5MM9+
d7GN7MCnh7fsiZGRNdHz4rm/UxyGrDmI5nXkvAVfhQw+QyO2GdFvF+qAQTkaSFj9WirJJnGl8KrK
QqoWqEg1LIj7lNeGaW6lW2/zwf96OoJAmdJ08Db8/zSHcWzA9iQK+Sd4tWta+9oJJdGc5llrJqpb
k3piAhy8DTdyZ3SHR+frDx9OgsZksgoLAGRgJNUfM88/F9pET2pA5O/ihKPWxwtwCrWxt1asZ3mh
tMcnS4A9wzCipu+nOYkjy9uyDszTlWyrFSys0S1QN88acuL30qg7P/lY+LvMY7WS4RJOgLXvj54T
y7eQ98usv8j4Ch/0tOWPxgn/ShkvkNl32bTLHltTzuUgTlMk5TcKOpZqgSjPwhzqZINDfCO3xLQX
2iFozntUM2UdmrGl3DEaMpXLnYXQ//+4OC+cUFy6qkOoGIDnj0/2LCnhrQ33tRSCUxjrTO94WBeS
taQdItrdD1C6W/YchW32x67vKWBiQZAJBONpkxrOPk79YvBb3MyF46+DWMu43UkHd0Vpnmep2UJg
++yDX0e43N5hK/7+3bbtwmT8dIEzsD4/Uo5CplG63r3YBl0IuANcbgMeTGXOI1KPyCHo0i6/Su+b
tpsJeKZO5XWiA4RyjfK05WWKkt0SKyzu0ap4mH8DXLkt11Tpdthh5TDvS0R0hYk//vTf703+bUsl
nsNqM7FuMLlrMBtY27COR0c5lkzAfRbujl/oSFs6rbER3xqKHXtvh24eojlg76m5LWnK7QG2cE/a
H2cUAdQ9/W3KBZ0ARlVw8NhkliF3vIGnFD/9lQuALOFnb1u4B/FIOcfXkJ5TAbyfTlT5Nm37EiUM
Y/oyys/BPXCXpftPg9myolLXMyHz3ynRqsBiNAzwjh4lGqw5tar4PdV8pDY23a2JtefrjiAq8gNi
68Bt4fRDKZi8AdbaJvm9Sb1DXbPheo2uhos/I+7lgM5lbFv2BGnjUGDMQm5lzRM7nzxzTWeW3Lv1
2MS4P8M8sByt6/+PZcfifDL5zEFRGcP+IwRIcqFHsXTpHrTQIOqtUyBcZGFq+FmA/Yt+g/ZY1Opq
4ErRdelngfDIP1X3Kp60HoVpvbtOX7Zp5itLbn0DZeq8MmvtC0EKU5g1Zkg7cFyTVSGh4t/X58TQ
7KDEque7/trCpVSMpjeq9M4J3QjhVs52H0E7hhWoLqFmHYux7D7D++OJ2ycrFRpy/LG0WB4yIWnO
oC0O3r6BOvK7aopXCTEX2FR54DWuoJHQnvBG8VzWPo6upZXhhegoXnLDPvwewV0xf31B8iebTlIY
nhKO40DjBc0cgmdDWqLVMpMUcDlbObD9A0jPvzaWUjO8fGWq3ekYVd5JYm7I6jpUE32iXT+anBWU
OUf2F55OLYIjJaJViNWSznyHHYvFolvTrL5Wzoam7wCfgb6Mj3tITo21EGhsbN+unoreaUYNr3aY
m8Zs7HzJ8HoVGfBgXAZYM+5jDoJM6sGhx94V3OpIYA4RfJRr6uJSoQEKTyBA1nNV4UDpSLxhImFJ
q+uCTrlh2ET45+GAgWkbT+soohLcynn73oGhytdJuYa0SgKoAUzqk72b65glqLlnN4XBb9chB+eS
1R7vGYqLjE1bPypwJoAyL2N6+3aJVvCf5irTJu76rojH3wuew3oazYcoVzhgnSUzKse1RntTgrEi
blnoqiZauz9CRC1CizonoT9e/GS0QSJuo6GqwAtvj4J/Y4ezqO4ompgz7whA3sK/Fga2+SzpwKe3
A/V6c5Z/Q9eM3cDmoD5RiPIqhxCy0e2L6hYXphTARK0rl7V2MbLbbWScJ2uw4C0TGnYkBqUi1jIS
vSinqh7340eXqONFTZYSzfVBxWisLMJcuAiP7oxtZI+XfKa79PX8KtQsPejlrFeVFCIiMr39Q3ho
AX28haDKcV6NtalvIhhRYAfynTvn0STv1sY9nWqQYjGbKECUQtQdEhikV+03X+9rjvnPFmAIjWbR
piHF0279+YixNE6TZiICVxhxySfGjnHDkHzrsC0C5ewH9l6puKH8atbi1AoObOXCtUM2voLvYxbQ
qKNMBu8HnXWd2smg/TM4vYxce2MzB48nvjrpKfOWUniZhhZGTXUQAtz+gj5zOurTYyUPIFNJFyT2
VV+Yx9izHMtblwzBVeeruSEDB9uXoUnQV7dXukkH7Ebr3j8tvqFXPdZJAZF1moMaYV9cl7UOfI35
vWTInl78Q0GEUs1gGHsmY1rrgFnd6jFzunllzqNKwX0dC8Wo2na8mTTxsiWIBH0YJIY1Qjn+lx5o
zyEy+yZhJlNx+yFVm+RriJszxB4FnZEKCld7uYfdqo8W7hyX/EvMrNaQMagV23S0TQdCI8xNUKvO
9ryE6BuFxMiWqNkBlkix0bRb2hemuHuALDI6SZ5xJgFNNnTQC3gTSMvqsxzJlhOsp8XDlxxbU4zd
pyXbZgy/LbmpIWDzWPjAr86af9ML4+cFQoxfckEtLKTTmqz2plcLBJdkL/7eriN7GXFOvdsS1bhA
yStBSUXpEpanNqro6YkL050NZfDYnvmbhoQVoGevt3PInt9F5U6ueXpok3yyaVtwKNKJ6AWEEmD+
tleoI+eSFUYUnO5Yf7vyYiSCf5y8KG2H+r7Vv/kkXqPKSALldIi6yfh589X8BO5kxbI4K4rsRYow
EhTlVpc8A3yHtuzYR2PxzUAv7g7ibigcGDcOtCKoiapJYINHw+tIbBXsav+xXql6OYc8L/mLxgxT
MRGFlLrV8tCj573ptxxfMsy4jIz+12YZ7PpyrwcntkH5/TTId8sqmsN7T4Kt8N1NvX+HHnhaAwaG
ZzqjSK/+fB8X1svDETls170d+u9BQ7znV13tDTLxMhH6JYPSQDGRCvo3amXtfgCwsD5aLSlpV+cD
xsUb66c/gj9lBWUbJOXxMMUHfieC2bnb4AXkgrFwMQIu+BpM9WAMzFdLctJ/kZEXEyil1gDqCdWA
pwqAVEklEeybOLb+oZ1LYPapPtXDZ7PbXdeCL5e85Kw2PGB1wTVRrOrKgmZbsIB3hQePsHxnYsCp
Mt4BBGBHocyT/BYZdVNTflEYpauperQzFm0I+8VbRganfFqvboZPqYbzsPFFjkGf/qirNWnU+o+v
+aavTuPtsXKzs3mh4D16LEjgnS392GqGy5V3YYzuh1dOkfNnRshNznQ8jxXI3vW0tO02ImNzNAU4
piZOZySCiLIDHKXnqcJTvvPKmhHQ3azaD4pLJYSAOSIUNkFflrxN8TX8HhrZQOR/nGWyPjEOJV3Z
NTric0Km8gPhRPigAhWhdDnqbqIukrmcmOz72uYcG9HTvxBMuSsLs52ddyyY0mi+/8WUfs9ImwCJ
vFxsudyqoKWeTiPipKlsrQXe4ql2JMO30V2XmGcAqJTtr6k+UdI9d/O6BZBR1wsudo4pkK6y9ups
nlOVj3Vu/hcs8IPHwHGLUe3D+vNS4TrtDlbGU5Oa4e2f98iFBkvcmnFyqSPSqN5TmqZuAW2YaMh5
B7tiAOyGRhiIw0odeLFrC1xcaZ0Mqxf+hzLEkJ690unxaYaGvAaDcJQOolj1EZiUHJp5AFEGTylb
3W7iWuqT605eQ2BPBz8wb8puZ/55RmT4VQgOeyd2jIUMPp+HMuQ0AsZd8EQ7ymIUdN7W5WLp1xnM
JMT72voiUL5ZMQ3iI4KbazmmV1DeOddFCmbnvVBKYI6egVoadFHZ79ORwYaJEN3p7B8Ye0BCDm6u
QlBkjynnHmwSKYAZ2oDk+GKHf5qLfUTIbogkldim4o4qEx9hY7Nn4QUlnzP+7Ck2g+TlEqgKwS0c
MDL5bM1s9pjdBwNEoEsEZRug4tsorDn2QdIWvlGhgYi1kEE9CMeT6PXEReOYbKM/qhsmW0dMXp5G
SV5uDACTHGyBzfhhrYbmrzEt8oG+UtENHynsX164Hpk6TLap7V2PsNTO3O0P6ChwAKTArcO/+ikc
Ez7Dfa7/VtGNMRwPgG9WkPDByAjFX5afOSRTXKMBl/+TiblBqkTmz3Rw8sxIUxXK3UumFLbKZCn9
jk5lYjtrslniHN7RbdfT1lfbo9F6fcR8lM1c+Oj6Vp7Hp6N/BF7O7y6i+fiSxAc+HKMRmtCpknMi
s3XFZ3RD9/iQ2kjTVtYd41Mk7ONnpX3ciaEo2rcsYn/QIg4FNVpa+LWslXI4dFBktIyIOaRy6nyi
F6k0PGae3OTqKyiIHY6YzEOXKjum+FCOHR1yAoA+q973KD2aEu6TcyWoXrKHbmNODQZNO5S2IRXJ
7fE76fS5svoVzM//A3H1m73AzWZ0MMw+PzJUgL06vP95QUIJLcxi3O6Jg4Zw5emMx9zSlUYG8O3J
8Mdhh8W16gX0gqyB/cAiEqRhdQsv7hlplvI44vmbH6+F3XnvKw5XHm0wKnmQ2cYWZoqNvUtBVXJu
cZpohiT1NWKYAz4G+3yUBwFIfqmWagtzFqm1wpeWIY9QSOlstOgiL7haDAAP0MdEyoLrF/En1mjI
NLdv6PHZVGhB3k4l9/0nirxmV+nk6nB/fR7SbP5hT4sDIc2jGS9l7NXKMDk98Y/Eic2Q5I4PwQxo
q9cQo0qRPF4j3pukKPk8+SHNaSLjHVi3sNCa5AWN5i05MHl6EkvGfxUIl0Jsr00xHhF8ZmdtA830
0+Tlg16iCOef1UKb2SWZd2+lndWYZGz+nps+8Bv1gDjyOpRKHI3kZJDJwc7X3yqWootLSn2bmizD
0KVZRH87CF1EyDjSZrRGaOFB7TTDwfKrjGt7xO89wUEg3KqNPd4UfmNiUvDCeOvKus15oMBtlxbj
xLJe7LS1J4ylvIrGnpD8aF7c9+IbnQzAaNLJaowqC/CKiHhZuW1sHF8TWY4ZKl4Gy7K4cwV2LEPI
uLqX5LQV80Jkfo0PAlMf/MmTnTw0Ak0CVzQtHOeuqUMcLIJKlvnUdaO+X3ukemGiOfKNu9ZH1BqG
WNLcWiDAaMFWrNmafYqwG3DrBCl0G9c/Vz0ZziOzZbwN4pv+QVe0WzaAOAWUE4o7KBFQIiBh8vr0
bhlN3kQeJOI0cxkCarfDZU8aeX8kNyjwTWFOmMfVb3dSXSAK6BE3ULofCzE9ayVbZdOgMu5zNMgf
10zmawQDiyXuu2d7gtvb+C4L2PzgPVEoGjpOw6QKQXYIs45X0TAaVkma4Qn0dWxhY1X2hus616/S
X9TQIiNgiOSRJcsaWrOUvKOo3vEKnpaVxzoWjgsDE0VKZF1mhlx6WJWU0RBVyS+H7dyEfTRDeJLl
lKPhtgjj9JxO02o2rF5ar0m0RIIBOnfH9q1QpUCeiEYychfxV/h36Q9ckCVyt7O5n/md1yhKlujq
SauvmvLQDUDYpEMkuRMIs5OxClLoBHL8h3DiLbRJFdtY7Tpno6Pim3KLT6U0T89cTVzuPakcAufT
tk1mwuhDoK/j0FMlYsPNzgtvE817Pc26Qj9coLDjoo5GkVxAIIvF0OG9a4z4oHVH7xQPYEyMIYIW
kVw+eCF4UOP3eGsitokcuCXZEtQGpeYAsRJI2bH9OQJ/JraQImigYgjw4a5rh7X15zIWsqJ5E/qC
I09mkjkU/bZbMSn1Dz1X+FyFyODjzg904WNF31y5nKURj9nhuSvg+aQaXM8E8OQHtdIzLicXuRdR
Jl0IC58xZG1Asokdn4rh+vqDJbH+QwVsrFrscXq7EEObbYwcZTd3Y40FfXFes9hPjOE20mAs2t0D
Z/A1IYOcVlmRXWVfadA0cwinbixmTKwPUVWEjXTsbNRS5MIQxwAHLjgmR4MxwlTwAByav7Orlum4
vrkhDu5ayQScphWxXx8SavWzCRmiLwYY0FqCX06B+LI13j77QZKYhwS7S5q53b9gmwduS/Lzv8gq
V3JG8uVc4w/ehu5tDDJiUSoX76diJIqXSZLiNrQ8P8GkeQf7qLkNxJ7c9GPyp0RZgWWjT5tUu4CU
K/V808oFsMfFoUteVsBPxqGq8RnftG7DEfH4Oja13yLMnai01PAXq5SS3Q4DxNqGrbdAhbMqLaLO
qtzeb/LZKPU4FUDbhDRVucWvSe6EbCZQP1q2/QqVej2LEw93DEXv65erSNXJLOz/d+euY3s2AULw
AW/OXs3sJS1bnP3WdIZkhlCxuxuOAcX3PrpwB8O/uDjcjedbSq7sft/pDKY4nt12e51zbOnc6z3C
4zQn9EgHy54DvfRTMFa3Yc2814jqSBf1ifHLt/CimU+eLi+5aYN6j8v6XPuWfQObsr0N99jNyTXZ
q3V8Uobo68O6MMUdCCzMztHz0MshK3qlIdNuiAYE/VMH5pA07xRvTkjUOgoW8jF0G73rDihPYKlI
bYJJw0Gidcn//J27v1/w5czUntwuMGeEPtwb0uHM8Fhr3FRQVxdgrXKeoPnQulHRtMImNASguJFU
4Uaxp3RRMFd3k4QCdwenrLvSyv3NIP88H90HLNCT2Poyg+bySnFTZLW0NKvymzaxgSJLkQyZofRT
FbYw4TxbSX/SuqTjNmAcEOJNO1LUfXmXuGmK7iby9hz1LpOc6Q0L81SMGXCYT7P4djVE9pC5uGum
BsoCbZ+3piCCK1vNIaoCRo75tW3cEHKXX/K0KAfo5eUHhWk/H9rYwZzL2M0vTQX6MZREkVmijfLM
SzSlx+mjn8Sdhmt1+NJOynM4rahKQni3Djvy6b6Lt4TPS3RWqlJ4e+OKBdY+2+Mf5Rv69lYuF/t9
VnEYxiONA+Xhmw6OQ+p1gUe75Zgbwvh8BXResk3BS9lA7xW3E8vVu2L1qJ94cKt7HiFBwZJefOPb
OgDPCnug/JPCb77XYgHadsZqzYGkCBwbq/VbJCRdYcNGfQjNkB8jwzu8ywusF5dS49Sje8N5eCF1
S0UYoOgIKP/dtUKBLd9l4WVp+HzCs1TBxJZqUc7B85y+nNH9fgDujHkZbj1s6+C3VHSSdaRd6Gcs
jWCnnz1UaOxcZKkcOrv1BVU44TfuyjL3AhFqjE0nLVkB8vHpI9EKwuUU0bEpAVMgOhqGvv+0xfRi
X9NSs3jHTD3ZVKfJUe6dDrVhly9bp5Zc+d9+ppnNZjgz9M8ignZ3atlKt+SZdS3mszfOXzxduQKO
Z/+DVTE4SpeO5NfYYJY1bm2CD4hC5oUxvQgN8R4qPr5xrgwcT1TVIxP4h+MFc6Vb5Es67aCtHbSA
Kh+YoF9MuETv66r1fvCg9xGYMuHecTfRfHbJRooybtw/1t+KfyUUu4tEfNTEzsYBMIKlUaj4dltu
oV/gCPJnih8NyO4OhYqfIO5hnav02FuwUsU3JWtHp9QI2n+UtfmvuPxBVEThCbeIajARTIR/sSDz
YcODWRMRVmnSe67IPkDUWXVn+bFZJqjJSVFOwZo7DwwyA8HhyR9bCWOrp5c8a7BAx6CnNxjZ/UO5
6zji5eBJ82dkzWf+R2dvN83sI5tDowz3ZGmvczWpvAG6XBBFzVS3Vfp2mh9xM0Ng4SP5cucmzsMO
M5VKZHxQHEzu1QShx1OOxMt9Qqoe7X74aS8/RnNvG6ku/BCfcjbcHSFB5RYGl+hFOReILRbKiUd9
5c7ngCn2hB/oJKh+Tn6GFCtRipj3flFwzsNrhXkRebJ341s9a1vVYdbZcSxrc+D4E3nVuRQ5mBJq
JTMQzn3BWlMN6skYvE6r+MNPWQReNX4g/baAkVzY4OOUTz5y3zmDG175v6Z9uHozP1DkSzusagSC
2+bSmZ1oFNiFp/AY3oIq3ilRXWe+jOZlQxtlwdZn1xtsiN/A6NUVfiQboepfX3VSBSQY3LUA1/MV
RL2k/RbTd4glrsBRbuXxogJKVTCRxn/lf0e7Ebl/OMVkWpEcQ9VhMbGeG11c+CFToQKb9BAq+DK3
livSh81n2daUcmFnDgkrAUxZ8hoQ0or752w8gflaW/8ISxDMTC6W61xlgCD4v8kP9Yb7zzE855hd
ULgXu7H7FZCpajhpc8OwkcN1Mvh0bDIaaNEMCCS4wLu/OS/gRm/oshydgS/M7/g8fFs6RTZfmqwv
pRjnE+1I5aDBNbaZXncWkQHBYnEPN7ULgpTjwcJ+XosBdFP0+Ajbm5XD7nTG+Wa9XsgXR8a0SjvI
wQXSTi6PQhzl9g1zN1tf/5bt8jpe+7P4hXzINu3OQJ49T1gIT8LOewEf9xeFipAAA7ODTfuWsggr
SPjhVQCAj2qPVWSp0P0VgrcQ2P+p/Lp7IWfZYXuYc+FWi6AqWif8/bslhKSx9qOW1Rbtc6Z5vYjf
wxSpwIxOYgFKtaj/pz/m5nt6qe66Jjt0iyoZ70edJK9hP9ooNIUZ/qqS9nuC3zpv2epBWwBdKIDO
aApOZJABrZIgYjnU5W0Aw7ggUNPFqzuZ5lgXNQwzOFnPfUcwW+lPL2aYY420KvtCcuL23Bu1+AOW
tZwIb9TbzAWAvvUH+SQUt2DQ4YXw0zBQJUPKr0H9oWl0clhHKI326WGBqLyVHe/ap8BfwWVPCwg7
dITfLKnxlr78mrIarvgEDCR/z67zJ93BeW2+mW49garaTY0zK8z3n5gsMjRSR3FGO4M5Dxc7879f
aGcdZNDCNcXfbpkWxe7A8zHNwjSthwlIWhSDjlKCP2fEDJa70Q9iVYHI/7w4rkuPhIkei52hhqxi
+ArF6QuwWzQwgZwGxTeRK5r3jBCd+aFVXYjEjxeE2M98NmBoDaYYdXuwMeAfTO2boZsB1msfGTJa
EqZQNwydJgI12GIgY7Lz5ryXtCubcBAoXotXborVp7Im9b6jIS2RkXWmcJCizh6huW4Ih3aJwlcu
KnCzmG7DwbYxo/0rWZD3TVHydhu6vQzYK67oUjyJG60bhfwMXxqquNP2916i4/2829j2NFaXDKvA
e4nhzbpCN+SK/Y6rdhdruB9vOBrD7cqxaKPlH1MrD4n3HHFJPiaj1lBBnKjU1ZelZccYamfxaGFY
d7ZkdTLSfeofxoT6yzHtR6uheqmltcjPhulaBVTsMiF2XgWLZE0pYR/gPPBQJhpnR/Tkl2C5tWiZ
rg53+3ZzrN6KMudJd5Iv+WpNedngmzobRkftigbAlNSuTJp8j5jHAtorw226j9hR0gi9Uk/Y/nDr
7/H0WvJZOA1ywGCOqf5bKe+hJFVy54fgdUy+McnNeRudIeKhcFG1dh8X3E3Icyjz7t1cgxTUxFSj
CbnYzU8jz5VmxkIielHCoWF4ow1ElNTmTlS0B+jsTH9e8TPNDgFfk7qW+Bhs/vuQXPWMH7A3+XbQ
qv9if+fJtahOK8vZ7WbL96TcTluiO9KEOG1d0aRIYqvSUCj8t4ASPrKjenmNP6ANn0DyNOIQc+K+
gOHJIGgkwITZ9LvI3ZX74Nkg5N8PyZgY1FoATMpUEpl7ICLOJPKZxx3xdkzVAOFxE8ipyptoP9CC
EEebnPDWgo9OJAlWUH/RAKdq56Z6Kryx10uUaxlmwwiwtppni9GjwaHuEoaPOFnkHN7x2E1xEv8L
PZ2rSkGJ7sFjgdjXwthFSczrRAOYJWkMFh9cXrQOGqRkGTyFiSjOeUjykJIiOcLUYI56FJIFqLAa
jcCdK+BkwY9+MyH4aTu20YbUc+jgPWNit6KJlaBNdMeH+UwcrUVzuDxDtwe7aYvEdR0fAX/eBYOf
ZaSkmaZ4UBEOxOdvUNU+ZDlAjnwExF420vdU4YSj3k8Z7jBLegBCBdOCdT2p3Wvy6pw0dUMBhVCk
Z2YUOxNuT0WdJNtKjqvirZBFMO8iTiemDhCTvOBuapP6lXxCEP32Nr4ylniOZmawKqbnL/Gzkdvs
UjsfEEfV1h9dOtrQSF+lvOSu2TAO7CuKgwTy1u+twaxOQk4ocGSPWbcKanEwsXRL+ZdVheLD/kmF
scpc5FjqEnxEYlOGMXyFMVb3w2RSPFJjWPsQFI9D4LUr2A+Y38Z4Jd3eIvlAkGtHCU/xgUjV5QYP
G23M3MYHEr5IOxB0dY1Mu3WzL+cXzy6D8dCMKvGKjW8i9k+wTGQQUJAKIHexN4kvi8kUGRj9E9F9
rnFc8OWLJ3V9ymLnmkgOQbt5VOoCGYu24+KRv2BFgBDmSFEmt4BrzpZnhcCdv4ZX/WSPUrV+NAUh
QPu6y1Y7bVIMZczYy8rdAdo33uTUM/GLRU8tPNXc/ktQiUfMMExPx/LhCkhAMPDW7qDC/0NqZNQ5
xecfhQPpiHNEhG7aMwqsGlZVNBU2lHr+Tt2rgHiMH1GhpMGAfynUZCPqkgqWzj/IPR6Y8g9HmItA
uZIQoVAE5g9W84rAcoVd9a1ce9rZDtvA0uyFbhX+JJ44qc+gSG5Xrp1QhL2tWZLFAXbcr8dXrIGe
DlKXfOUXcsA3rOzv9fuGYRKSfvGnumzcQLhD6t7i06JfxrcqjPCwVieXnGpcZkqvolGjOKi7+aP3
LMx7piOoGbDFqb0JMFvJ0ExybVPQhMPnO/fv/6+ksxQxKawnYZglCKMVEZ32N4t57X8neel2tvR3
7QWDgl5CZOEwgu1PpvHr3yaJKFY45b2IpRScsFLV4xNHjMJn9PQIyaOEC3un2hgwYpPLLjdApoqu
xe8I4nr8BKaOhoPAggIaoN2sW+1ZfJA8yNex4edQvUqIrpi6nstF0tlR9d2KkFh7wgTLByPfY7YY
bjWZVy5kBiSUN8GCNoMVNsLVEcntXa/h9lAeettcWN820DdRwPkbtnR/k3Fvp4Ls9JluJvT6N/8i
VgPGizYe9mud7db5aLI7/DO4cLR+oFZafL7vhj24OwmbFEJ+ZnQoQQTY3m5Kxq6SlQuBIDgGodyZ
oXlGjLuF6rkILZQv0G0RqJ9LBMPzNdFxTALZcsrpM4eTmGnjLD3c3ngLqeVMa8PzSjzijAQXJ5+A
giiJfyNfwTnHWzZTlafM9LAKw3rYGdmHvIOXd1cdJBnVmR3RtNDAMmmvNQ+X24vcr/40TPsdlg+W
rtrHZTWqXYGXk4cxzN3ovIpXqVxXRrk0qGrSy2K+6FRCz+e3GCz16i2SLrcuIXKbj5xjtRie0KZc
p0aIOEU1j9Krik3yB6oiKSUyC2PzsSRB0UDz8O05z2U5QKL/xd394bmtOvfqh/sF4RNphufdkISF
8VLP8bSXQ1NZMCprqki5lpinHOitVqPEFoCUuCif3wTt9VxL7BeuOu3Bbip3BsXI9D2MG3lp7nMO
kJPaeWswuXjsBnXImp4jagcQPhAEE8Q69IbieCRrVw3H8gvrgBxpVfGgFDJGa9WaXHvqeFV2KUzt
M6hRLzydKqxo17ThVDshY+AcYdmGDFcGYQZitSXyei6E8ZwGOx6o9yhcipiPzVyrTZrBfySOCNDP
RmNZcKQ0/1563MWaf4EXOfSwK0ioGb83ZmjfyjgxgntpcSJNf3DcwDgWsoNgQwtV3Xn2eac2ljUQ
CAgaOD5WWoLKHpTJrH6DDLxVo0GQ/MvCZZOzcuLe5zj7qAsv1rNw+n1TJ4IRnh6NFLT1X8NYXpAd
Ev8jT77cJdh7ge+WgGIm4XVX58DHcrgC6zV3v6WiiY74nzTocpITSiSyuaLySulwjaj1ZbTvp1zm
5gV0XOB85OqC1hMQHisGn7S20FeEXR2IhDnINE+dHwHUbj9RBXKVHvHJvyoocPfjrKCIXx2QYsBq
4bwtFnjXxmBnVsevnIMUP9ofyLZ1tdTfTtyQBt/qYCvntPP5rrvK9i7AskuC/aeSQmQYI3RL+GJp
A+l8pX47/hE0Pjqxixel88TrXzU2L34QTL5Xs+AkHIQCvxFkGCRITFCfGsQMfQGr5X+UWvwt6e2g
SY6o09vBtgVyQULKOuVk1vXWQV3FpHvxjoZyHIk9zG3TDzJ0IPc/1Iykx9P7vhmSljlYfKnKg7yx
11PJpJMSHg2CwwCNeNlWAs8dDPcZAGQHSGxSqbyf/l/8vcL6kp4bfITJEYMQt8JEynDOFR9kFcJf
JrHCCCB7kSU+kajZdgGfP/5mq1IUBOxagbWTGs+kIYGyVjS2jo+qNcsq2MMRTw++Nj01Qkqarf2r
+IaE/fr6qLQoLn6FsuTi7hxQdGT1Bn5BJUgCDGtrpcN+7zgyJOyK4hVjFwNMMO2RkE/x05RTyixO
Deb4hEJ2YZI1Qd9MHyCPu3QUolSAwSKggiQ19Znx8ytBp1C4eVJbMXQUpKJk2QswZFhWoZXTr2W4
A/bEmB3eVBHs+/ITOMazPSMOreDCiZWX9x8GpUjWiWnyceJvRLf3KTN5HV1XewC23QehCIoe5A0o
0sCiOvVUAJ66qaedgHjfxISYnGErumnyY66VN9PSUrQto2p7WiyGBLq+P7aYM1SVFtpLhO8zfb6/
hKGH8x31ddlSJ4uPvcJvrUIG3NXDKyIp9ylyH7g4ByX7pgIDWiQlK6ed6Vvs5sfuHXeis8ao6i1W
2UxyAi2xv5Yae7TShIG6j0+YGRVu8FEPVvhp+BxSAUSRhoZoxPT9TZT6BFOp1BeGOjnoZwf6EWv0
UVmS3cCXjJiHWkGO55v3o+C7KTWkxXJ/zQA+TfTCLt3Yzz6N4YT9Pc+TJrtptzLGKClwclmKpcvp
H7UK1mW0gA7Qw9/gohh2D4iti/EGz2f8hEthsedFYEXTW0lrfxea1SzJysA0dIA9tCfzJVFaFLv6
n0xRXsUS+yX3H/CFC2jd+TJ0JDDUopqueWMLXDJIErFnyBRfghl2NnfMJYTD9f6XSNVVrZa3X6a5
f6knpS9Ld6c4Ahm0CF1D9+f33vICs+pllcVYEPCl0x8h6waNGns2NNXBTMCkzWoGKgwIskVqeHdN
6M2veZYCmhLb9xGbgNCUfWYyHuVRjA4gqbrFkMlji5FX3i5HhTfoHTUPNGyYgVUrNdj13Ixq11b4
jqmE6C2nV74dZ7Z3QmNHRtOmrtOED96FGGpp3Dy0O4ELCbEdXS8V5PGTFnfAJTTRxeSsv4TKORZp
HGianpYAUAtUIUIYMNpdzzkgi0lJPeQ1pfJ1jMX6LHv4G+Z82b7ZHn+qEdLP8ZBfjzwJeHLQRb/3
QY0vHPuZdNfQPOX2ogp2SVNUI8sP/wh6oKtD+tzw1oAaPQbt79Gp8xl/TASvYUr4Xj0CICZvcaQh
btM7nIHSL/APS1gGCHedyqbkcqV+oi2GqJ+Y40I2MIqbfUjy8gCzt+rLSV2DpWdHcAs5MBSHv8ou
xE+r9zHESWHRhu1pIOZU459iWaL7kGKQZgJPv9s6hGguBxEqSNFq7QXx1fxn+atT0zhLpkgMdsKg
/GgNwly3Ip0Fmr3R6VjZTZu21wWU4wFHpfn+kvsS5Jncytg4m56DMtazECvHcZME5BCf0Bc+VUku
vQNY41GohH5aJAH/3OQZbL23lRXvLSrN3p/PXVNWypxd5zoQaCk9DkngT36ij7eL2vLHaEx6Epsy
f6U9EqbWT/VFJ+cS5kuJc0zUGSoRo7Gw5Y4m4S5dDUYtKQU8nVK/pZZsfqP47BV3CDoh1xlXZvc5
/HiwS+dZSfbaVUa7uk4b0rfTgMyl+5EtaC6LL050/b/FeV4R6rJHFkuoyRyayiHjpMivvzWAfapB
RbbpCTUHum59AzRsf2YGb6epZIjf+mFX0bIKbQWkETnBXOjjuh9/DWKs7GCDCmevYHX8PbPRAGc2
z+wpYxjm7jvelG41Xy/R6DZMnSJkKYW1OloY7tc0z8fmdPtuVHxyWyEqO1P0PNZrh9+vhlpHmDWU
q4KCd4tPPxvn9A630jgllhdgDEqtwpprHTHIyInn+p0FCp2luYJb/du34dlX+jnsXt38bv1MzuMB
h/8nicwhF6uogevexiAfItB6ugPeDQTbh8046JkvuFwlvErFxKhD3MNymSGJ8pyRZVSNbu9D1v8a
wL29VW0pEjobhMfSrsGn9HUph2nsT+uTruw+6TKWB8XUu1ej4wYRtOEb7ynuFO04x1IXtUv8YZAj
Lk84IgGHny11CfAnNbCYclGmRB0oYDLbXTnu8c9f/UWTBxl+xOToG059AgBE+1ygq1zzsXn8ZaqC
L5lJ8tf5Z4X/P4EbGxpl6KdWc19ZpNeKpyNyfgyXiir+NyHiioUcCSBG5/qjfiJXPn0gTtJsPUyj
6IdHVhwhNEvWAf5/icTSx61edaoeaixS9UdtcdH9mXhg/7ytGnOJ/580wt5oVnIWPuoVarnWVOr9
uzJae/n7IF3f2dOJPFdyoZYLaNwRcIhG+Tq+cA3vo9ImD8L3ecVoI4N1WKIJRjiqvNplXnc81yPL
YPsPk67BKguhNKC6GVAtzKpIQsqwXMkqksoBkQm+ffBMwHmuxWrr+RqyTSJDFq1BeEoIjOSZwdjI
vw2UY1noRnbbOHd6paHgZ/G7UDbRfcg9Hoyi/RSQcI3GYcB73ZZvRWMGW4q7m9E5cM7uK3ATMxQx
ZKfrbLlOKUBqDBMv9WXo42F2PgI9tKy6aU4SOLkMI2oHW5yiwHZvzMRz7p4bXb0q2RSFQY8Dl1qF
vb7/4Uke+cwPdz7/dUsFwNWn0gOaMsWi72dH9KPdxFzOCsc3SO7zKSN9Axoxu5sVWcvnXlSF850e
igE55cmEHwSgKZ+OWxxjsEJPeNvgtkbZH21pbYQV7TJwOap24CMdqfS+9BCa2gA3bJ9nt6IfLge4
F9wFDCRudNisD3quE1HOPhYE5mLPuN12YHziydIBsqPng6QeFsGnBCrtaXVCAM/XjAP+Ia4kVMGM
nFzvfn+XYqbVHoGaV+dB0o/d7+ronqEBYa2rIoUceifS67uj0hz30+9rza0haHTETSDOl1WdpnrP
IpiClhNhLADfdYu16rwaNptg9xDA9OCseF5SExqTKjr0Ep0aMsYoiYUt+tpkJsnip3YK8gCSoHQk
8FRtDbkqf8kz5BemA2Up5iUqhU/nrPECx/Ka3tRoHxXU9VMh2sUzxAr6Xrr90DhADDeWh8/zi8pI
M1izFWqN9p78V39nnFPY2AUpMYXTshLcydx+1Kd5GLBye3lrTI71pZWJ/NEKGaRp1hEwwnYx4oI/
NTecLowc6E/Tnx+p6CsuvuqE1Gs6U36UdP9H+UXYHVDbiqfa0xah5JZ3GZKrhJflJ6Py7XfZ9zYG
0SP1wQFT6zDilzZWz/5ZfGj21mVvDPlY47JaLQU7Ebsp+l+SdiP8kniSWpikg/R28BNOu+5asxbq
bf5xpyip11/Nyn5IfTNRLDfYkACMsFOk6LVP/moJ17fqAd29ckVAlXorX1cw6rzvQLonlJpCKGNq
q+NiEmz5UuDi/KpPqwRvjnJHJzxHuBeBFn+hAWsVtZ1qc7/O01JFOA0odf/rgpaKmKMBy22t6aB5
sXgCS8UK346/mA0Fmc9hciwosL91Q9fTYkriDaQH0oYKODAEz9IbW88snpvSpnvhrbCy1FssM0J4
wXTc/BkkjKWRbN33q/IYvyVzDPgTe5/oXo60crUCAdK8jhC5JLfKEhyLGljmoEEjkI9Q3AqURIfC
qioXoW6IxmHgJEDo6xNLssXXxay6iOrS9up4aBmoNeDgNbg00d0qhCm7XPGZw7gXbwqZjUkOpkov
bByXcTLpTEGPOC09ft9SpBoALcb3BKzLwkSNHbP4PZK2TTCiOs4HJdDqCybhLEycoM+WrLCrh8js
obaLuXT1HnWFlapaH5KyfOwpi4SVuxjcypCz3ReMjEFvLBOPkEKtMqfXVJIOVcJcoTx2iv5Lt7qQ
tbjnszLR8aF6VCIMAmvcVZiZMMAdZzG+mNDB6qmKwLuMUejYlfcZSE/5yl2fidmOTPEn3NZSQy0L
tkTHyvIqWLJVoz4mLhZjWgb76OWZd+ORgsrcphdYHAdulmNeses1evNNlXl2QY9EunvNMKfnCdud
ry1o5VEuEJfap+j8jK5fKYbmQTPK6SXlihv+bL5uCbNkyd1d+kLE524lIjoyx7No/MFTFY/no3Af
fO1wHMiOLzObLDF/FakvtCmC6y/sIj0lZVTrzRC9iOHLkVdHV1MQAzoQMISPdpKCBwGOmkF9fR0M
gQTb7MDgxSEToYISvE3Wj9n8BV+f4PRq/2LObry+ioHqua14fY249GzeVjmS7b5HdurHrcbu95z3
VOUK35+Wh3lcZ75Cz+uMBR9nFvz19WBV2BnoT4vJI/7FOrg5+TDuakL3nm9bCqEB8DuPWU6JGkYw
Q3S6p35WYVr7Kg292qS1G5IE3Y+geMiqVRH5+19D+lAYwtgI5NMgqp+2J8kMRPGVJjhs7tRZUqiy
RGsoKsgMHxmGy9ZJ53MbCGZL3w9KmRpnyO0vY5LdUKVrEd+qcJEd/IuYFXtD6Nlht/xXCRiklKDz
JBFd2hI6TNEU6o/lGz0NgacQXmsmVB7ws2Wl4Rsoq1NSzf/Of4F9AsKY0ZtjcvnGS9mXYuwSz5jW
fr89NA60sj0ltGto7N7IcUx2mLjxnrfDJnvSKXUMrtZ/pDpmU9r+YJOBMNHd4yjnO+PSPluzxiPZ
Xb/rydRsG5uzLgwbU2hnsbSp3Qwq3oa+8qp9nUwJkghSrZlbS35BXalswdUZO43GEegD0aXPKVXJ
pUbdGz9Hpv/9nIFLCjgliR48boxAtQPJVv3qmqSafAtkXRpn41HvQdvXTUuNgkXGBe/zktNvCbng
X1aEH2nDQRqOXIJ5hLD+3PlB0HVOv7XRfC5IkI7A3FgD5G7/Q9BYLdpi/3+VI3MOfHpG7JrtQEmy
3K7afnb2Ei8KG75ySyaGXhs7INEtDrZKsSxPHDvZwTVwdE7JYO8zR8PpDjNRRtM0Tu2s9GFoPKGd
rAR0g8UVaTPHptLtJQvPao6q2O4ALNWeCGUMNmQDK8GYP+y/y9TSXy1FVnC7/j7Kud6C+60k974r
XjHzJeg8MfkCaR/pEb5/kPABfaFKou3Uq0qeTbmJBr+UVZcOuaGpiqQDFwb8Co8PICrm+yjFgKXv
almqQL8TXVptGoz+ukxo1jdqD6L9w0DuWMtmhyK00Q5nRIbVorTHUz65U+3LwPyWl6adekM/8fqi
SfPtsMmBtDouOZtTTp7MFiuOROwJe8QsX+6Y6p6jino7j9dui97qv2cs9iwYPht/NWRbXvl5npDr
jf4brlo1++zS6fzRhgCMcFbXrAaA3hDz7aVUnolCHjlnkvX83YP0lQr7W9bN3gQRZD+Rn9ERISRy
RDxksB0UGGlt2NG6xqQVDo+/NrBHQ3FUmUwtX1YdTuUPsjb/M5NNiu3mQda+6dWJ8AuK/LLip/tu
0i9jZkJCIHvdvCM6WAxnd76cnjqhoRvcx/lLD1ghUaIM/iBnahZXVfbK+JbgP8BsSYK2680E/JCU
7zf8WiN78Oqfy0Lt+bse0/3jguE3lBpTSt5fsryN29R92z10O6GYwPSSDho2fVZcKtD2u4f/3SY3
dV0b+BVw4cEnktnnNottXIgj1gvzZcJwNzkLpHViMb6ezqXviTwoT9E+Kr75BKF7d2WESGzPHVtv
+YYBhlEeo5uYc+m5qv9OZqHM7pZAEsnGWb+Xt1DwBgkcoH4UTWPyEBatHTnqcaW7J2Y6TGn+XrWR
+CiildMqe28/vzCe0yFvrPx7yKq+LRJ/RLSftenyQ+vqUh2RFiGe1C8bRkVwOOgb2crewgV0Nm6g
3+mA7rOqyQ9oxiB159phZHYzBgwITBOTbvmIeKHMqS9jfHxmgaHLGrfbAMFqvlgO2YKboE6tZ3Af
wo8xk1hPqNIm8H3qNJEYHalFhzhhaJlnsqyQZJvNy64EivD6zNbQgeJSnKhH/eLNrlpPgmTCQRL9
KNYNu8niqT5ZdKPSMTsEn8NQVBgl7vWlPVZ0JbJl/ipGnGW32jzhsYiCWZlIr8h/YECr38VoryWq
eueyjrJudtJRqDoWSeBlnnQc1v4rt07p+SinuFuX0zYfdl4gf+mTowrZwQ3VpLTena0o8Ds4bTlA
6PmAN/n9ggxj0MpLz+1YB2G4oPHAJ2cb1+ZsIf+GXwZyzmh3idsw72pParfMwt+y4uEZYWDWZhlX
yDQhM5F0d0nM0yY6Qzr9dO+huK660neotm5PtwzTSO6ri33QT+Nq6JNavsTJ5S5nNIIjRWaiM0y3
wdZxcjhwkjazwUAyn8P9DkkMaqvVl73m6JtNX15IBIpQBDntZMPZWmba9DOhGMf1G7e1BGilCccf
0HSv9a///+PMiDXknGOWx33neIMJIloVLqp3vApjMBhPEscVkUgqzesGdBMngeHIp8wZdGrztG4O
31G6r4BTRGUiLO6xLiXDgnEptaq/X1KgI4E5/DRbYK2Iip71he/u5E2BZ1lq/NH//SMZPokr6tes
BUy9+n9F3Z/XbSgpITsKe5DzPjT616vXlSrzw4cH9Ub69VAyVfPeJWQFVKXDS1JoVSsB5KK19fdl
8F6SmLHrPmdD/0uoKXS2JveCf5gc7ewjREMJ5xEuoCMVEp+/oV8TCQ0GTYShO0WuuhWfqhPYKDlq
ZVE0e25a6sMn9fghXuD/XYuJXKs1pucLQBgGh5biolDx+/WtabK9JIhpp2RZFnVZ3TAocSpMQsE/
4WCogV5+KpnHd4hGh5l0nz8SvQqS11L0QHi5lEkjNkajTP3YRt8CYuR+IUoaEw9gsddHcfuw7jhV
5zvkG8WIZD2AtttfHxE23MWz9iSOYMwJaqliqq3GJ7BgKlEhkplqqHASTMED/77lwOrDO52r8Ee2
YElF2jqhDYTo5tXFftgcuGnRRe4sXBgB+9ir9JATTvMExtuw1FBRZc7de1FCOEyWbi7wYqYtPx/U
YNwbWpBuR9uEb8L/YqSg3/l96VZXR3vr73mqDxphVHFKD5Xe2NgNJH9FMuX+MyYcFYws0By06ivQ
x0H+d0gjEcHTWrUPK3D9QCXnwYidtJMC3O9C2UCoHPQtHTx12sUje4cRxCKq7G+PPT7VkgK25IDj
GdZyhukEkMlMFvqmCNeflkMj0fpzKQmJtCnnKzDx5zrpwVe6ML70H8DLU9Jwo+ecz9hA+xUOwpwd
yZ8KQbMKqc2gYmL+PEBJqcigiv1OT+6mYpagnosK2zB3ohremiHZK8/trjBJ1GaH6R6tgPSi0TI8
CgE6lwg9IAAzRYknusYD2v50xOb3fHC1FYH4g66NFOT/oc/Ncbp+In4ht+6QsO/SePoWp3iInvhi
VOGMjvkzbEM1nEsuhZwIJ4crAZVJszMf5kBP+YJSkRpMvWD3ugw7cFLssSjxw/DJ6oAhK5WU6CRL
YgS3zL2307Q5x2Zum4J6+FzEBRIYH7oB9SYjm9sulHzgzo0rERFntkXQn55Qw0eDuxSGaHeFQm7p
QSzbPfO9utDtrIRa6lJfLC7qxNZLFGZepPCguCiNp4phfC8qFWqLvrKXedcKqVPOtFBRLOaQo8R2
2c7RgRmdaHVG3Zr41qhDNV8/wG/Yg8MnYq7O+0OTVsLl7OnjME9k+wEPzZsdnMDcMb2kphRLHeMS
XUXA8e0qn90WdJgY7ILCkS7ihoVc2x2ClC1pK+gy7ukXEtQC9E5hR9Lx+FAtRsSZJRtlgCoHi+Jt
sfKcfaWcJc/ML1sBpDKPHRS02E9td/x3yzkWlb1OzRuX+x4biXA35l+1/j0Vak7SDyeQR+odWBC6
Znd9aOQ4ScxQZwHIQ7vSe3n5ubyD15RI+3xVS2UIha9gmlKyXRsI45Eh7bbgKbPwZ0UQU9TAPEE+
hc9ZsqkByg8MJaCnfcylfcXaMEXesnKabd+6ixvFGpQOwkZx+Y34QD12ZPAhdZMsSSYUqhCHNjVP
u04f77WnX0+g2CBNnbE3X7UNLjme6RSvI1HCZK5jXLLtsFaZib2uc9g6JrGxZDfTTRdspwDCzYws
AA6rU/JJj1/qmd/eTwEIK6KOQdTjwVGJ43BxXRiyJk1Ca76QHJI0lXudMIjWUdlEGOLp8iH7JTAf
DzO/AdGubLaN6kk+8k68KUmjdf2FCkUKq9mYR9zUNlUK74zktY6I03ESnVCGuP/7Y/UgbdoW7Que
cAQ5nOd+LDQLgPd7+FMClfxUthYIFtyhCccdlMATAcnzB5M86y8qkO9aRCp9hsBpv6tD8IGCIM/D
5v2Z0bER5CxAcRMs5NCxGtOpfwCxbm1PbxQHnUtUeW3cF5BLngnxQb9H054ih6mGtQJ95xuwNLNz
tOWjOXs/jFuWWL8el1FaRf4RiX2P1s3apbAP6o9e9FgnBckgXZ9I3oahTLG6POLXc0lr1ChsRBYZ
uqaKQ+Qi14anQhFAsuz9LZES0FHocqcsZMsyzLA4kfIZEnOjyFBHrGgigAvr/CAuaB2NEz5q12B2
LdI3vil/1CJg7YMrxyGfdzdxV124Ct459kOA4LjNSXeBnkB3PhREk03wxUiGNToUqqUpRXa2uFfj
qdNLOXLIYshoE4XT9mbKW2m9YXS1KADDfNvuJe76gihKE9Jo8KmIUOpkEIawSXxOFACmtzU6+Q9j
IX0SlTJy5tkcpMJL49+3sBnmwbVAFujQyipBdv4U3kJxP51wJno5xj7KoLzH61kwqW1tbGaskDf5
n7bwtkZbcI7mhjwj1LOakbArxNK6Ineo7omejnIkukDESsGs+ZLm10DPeH3THZ4KPazgxQ1nmRX+
OdQT7akNHmtPyyE2Eep8Kb0tHnAQ9fvlJ97tjO4HkuhqViZuv5fzopJOWZ7o+ZUbDT4Z4tJHNpOz
60YIfIxZGAryWxC9U5xVzfmUzA2G95C1gg8JYRrjPLJjeNEtwS5T5fB+Njzn+0QnQun2rmP6evJF
Nd3NgaxeLXxvy6AkVTVMkFh+VfI9K+ykBXBszXjkmlglJdGf8TyTsVDKO0qVz0uY1cyK70nIj1v9
cRsPe/rNyw0BnfVmSZW4q1TnhKWoV+ai/29M2VW0ld8yL8IFhrqw6pJx+NiCtNhpbLoK7iQVfVx4
xCrdA1UJPmLJ4pf57ZERn9C34FA7+eSw99G1agZETv9XKQ7H9NDwXNf+MfqV9pK0Bc1/mPe/l3Wf
RNI+ppX1m2dKMz19B6R34vGndpqhSgTLYAKSXgxYT4xflwW6cV6qsMzrq4iLiO9dnAlGQdr8iX0e
z1IRNfFJoKXhEh3Ui7lTAqTusYGaetmGd2P6ca/nFlbo5limEdWrZMUqoKSQ+9lqm6Ou+krpBFbd
qJaE3aT+r6JIG4ly+85lm0LFzxUWZ5LfE1SkKIojxgw6GKopFT2fFmQPlslPV57cyHdfhF9Fa7iS
tWanFPZSgKwbXhb8vIb72M6HtrXuy9aUn9K3jaA4iJDvB8rULDJA+ZOYxFPb5kN5XxXQ73YDVF/Y
OY8yepN2Q/9ljkML1aytpTBpTtCkTqdme+6sd5uQ2zTDYG44zfu+ACF8/IxUszQIy0DF2URZTH4m
gH5v0NAoKJE7kTDqVder+SVYUDoTeTZsvFZlBg8RQx2Xco7BJTDERn8hYZO81FzxnP0sGaiNZE6Q
PyNd05JGkP38WWJZHM7Ye1gyiwzOi8cPCUF5tuI13kJYeWkR1C53m3g2fk8h899vSZZ0D+rCyhFG
CeJDfncLBKUpGtdkSQEH4LKZryffXvpn0JZUBXP/qEzMyn5rbVYf2W6Fr+TJn0tmgyRn3Szhj/AU
VUdz6OialvM+YKb2HBixUVAPAlC927xw93r6d9ih+7UTpejTDZ0eNOVrl16Ndx0jHbG38+elCyyE
kUI9dLssur6Z1Vy1u1qiQQFIJbNZoDewMWawxmOPB3EXmtlUZxMMOMmeKVRi4CeNVnwB3Yv81mug
J8jsS+A1ZDBVu8+Yw9lmN9f+l79UzNrbvfyGxLDkvGW2T4hPJ9tqHCkqhmqgljlBLuCn28erOr3f
jB1Ri2HJ2tW3rA7wW6SqsCK3iTENwg+x9zz3RT4etfpihuOQvGIYqW5P/KiGNsEaD2V0ebpUvMzJ
2KAVaOsFchBJlT38j6UO+f8deXO6AvpsCwkkhzDpOkc/M4+d8Vq60tuQb4CCqJkWIJ4X8x4s5wHy
3Ee1uN62bYrsWvCz7ZnFt4bb6MGW1zk3guonFovuVHF6FU6VR03S97azhhwwoWnlb9q2jxBADRoi
8rAIVBtmelsx6Tl/g00uhyIPRs4vlLh6dzuTjJKFopfQR5nAMjL6xB8DsMmWxkay5DZI1seQgBm9
klkswhXylZxPs9pBj1NL+KibFaKBJ38VX88QJ8YGQMs8/9tJpezu5McFqq3rI/RUioD9pNCMPpoz
u2OPOcGPj/IadI078OnccDApzG75Ze6kGLmOnWA1w+nEuFxs72x51yUChA2tuEXrOx4nodhD7L92
GahPfBKC2AlJW95oJtk/Ox9oYBL0Oe3eIQa8I2HsZozgSSUfy6UI4ZX/FEcjIlmkRAdjdpr9xEsA
Kz2pdb94RuJjVUfjHhhMH8Ceycviz/YyC7B5izuAvu3UBKmAYPDJ6oLhq7WghyWgrqPleDgcsGo6
e110abJvdBHmCCMtiMjvS4d3OxaNzhTtW8u0be/w2uXSwXb17hOp9+khRqa1/JcY2ezvyVjznp9t
o01bu3VRODbMD8BTSSTpGm20krpUbun4SAsXT4BRv0xXoqyRvlxKotGjw5tIwy/q6KSqLYTpiWTY
QESimHHAAT8woeJnDhB40km8lepDnwZGWaNQGV/DbOaBs2PeWbe4xsLlvsOnX61A9YIH343TCO1h
o064hvabUACDdcebq67RowPOmz7HG4u5/y2pwuCJl2UMe4TWQXss0/aW45/JyKwjnRhW1DT0HkR4
QhU1EnzJzgvk8TH74KxoA/Yb0dAKTAHOtRhdkVW5s1+sFA9hwqQ1reNZKdeXv2VzwwhzIQ8kfWTx
1ilQOZJozfGa5YzAB43CsN19N2dvIF+7rxZ0+wmUcFrZPia+jg152wr/Akp5xWtZI09A/juHRnWg
b/uRaEgqS8k9YFw8iNvZWWy2KiZocvmh65Cs+n3cWk/yAFMbfOFXl4Wu1EQXPQaRs9G57r9LcQPD
XH0tBQ4pf6jLedD9nSxwM7CRMpbXwcXbOhQO80dZlljj07+HLb/LMZ0Kyd1/D9EpXOPCHNbUz76O
qEgX2ezEBYjWzQqOEkbX6u2XhUzvq6SFiBEV5Tmb4TYa9pm1bUzjc3t2z7FSlUctXOdwezaQMSgn
z8VSOvfwjUFnqqvYcC86pu6zh32xIT4yoyrPd/wfpxD2U09dbtjM6RF7b5EDqXvARbDoB5xGHP2j
WndfEGSVGAx6TGTbkTiG9LlFyLQJwijVjkAc8WHPbeITwe1mry3xFqDefZpBfk1k203CSO7HBbyC
LqFqJt414IQIth1D8GXcwygwsit21QCZ7rQW+H5nlHvwNhkOMV3+t13FDz0CqFZLShnOjmwauyDZ
iP+3QDx4T1jIITyMYUrpVQdsox0lT59nObWjHy8atvyuzufWApcdmWP9qQ6i4omjJPbBXaQVDvuX
/ZkVWgd1y2Ooz2IcnDE1mm9qwb6K9kTqmv85qoLPtPTrmRkq/akSyFAWheJMDQOJC1jFL6/Hwsrv
4/N9iTLUIR9jkb7RSDVhFOZ6842FkvUNfDZjxWleNgWfwJJ3Lizm5YgzjX50eWBHHd2cPb3MOIus
lSrBX0MBMx4uU96UBECmtpbJ20iK0Jd9W3C18h9Iacf/oaxzZk+5ZCpOfCkxKqz9X5vwLphEr8N2
fuKLADUAuQWw9b/aSoolB++D45MBPHjTegQaN+H+puOE59g+7ahwI72tmhcnHhtkRvUzdeDJah0F
QNwin5f50+Ks+6MzNB+0k+x6AdB2XHmK0dr7pS0tnrmj/kvW8qMJ39WAtEnJXs9NKZPFkP/vZqo3
7NE98m8aEI9MIk0S0m/x4lOxstIFsuQ+Z15+QWIzM8529CteNrZkWwVMUTsb+YFqEN+VXlTA5L2c
A+44JmLUM8acS3teWxohddAlqEfzpJTCL8zyzNL/i0mtmwqzK2DYjL/sSbjQV5UvLH50QQlW2mz3
ExPqwHBNRNCmiKDBTIK/FiPcMsKPo4E78HVnuR3Bz5RGFFlm9Tqn1QXOkmASTx1w+7lI133gY/Ht
UYLu+qZHhDKmHIBbf5hcoWk6fQJ9F67oy0xJLov6d+TvTaQojq2Fd2kfGKHEW7ONtNw7P0LnYxQn
tcuQIbqjVk7T2ff+dvBp44oRoUs6mIt8oZ6pZSL8rYYNArnJA60mNzu16BR2q0xJNMy571rpL4VL
kG6U3z7F+EIt3g90eyfY+8Fi50Uncg9Gn1ywMZzQlYjoHgh8JmfEJyoIu4gk3sd7mK+koTXUyMy6
9TxBx2csR35GDo77+86chXuB9aILGrLQXcP1zh0jxeRzw1/F/2XSbiS5fDGWklSMb3fNjIvouqji
uzZkOTdDVN6XZSuSYkbhxZ1gAL1Ffa3hBPm5DAAuJ+LCbFWi7C7CRVkI89lDxPy+5FBKtpm+Ljtn
v6T2pycxU64PDqyEjHeDOxMXMV9urX99CgoGveOnbGTXu/Z5kIuLA2zW1C9Vb/Fg5QHzSuP9MZHq
D07hHH9dPfR71iAO9zxeRMut5V17kUXzlODD4X5gFgJm+jQxo+Z6pKUZRsNtBoelhd3psEEpFsXB
V3pK/qHQIL7oiKi7C5W4AoYSLJzE3DJQhZIihs6Dg5TQrAAgAA5E3eBbMo0vj8UIe2Zqg6xrRmcO
rMAjB8bfmwYI5VxFfoS+Q+bJoE/MfIH66G00PckOhRGPpFyz0HMbDAs8Pf6c3gSEYJEefM+W/pys
0p//uXQLIupSinIw1dN98NFcc3JnJMb2fg5XGs0+aJHIXH2JCBFs7/d+lag8ZMt113bS57JX5//R
8hGO/Bsoe2KV/pMAJ3EeXKV0bf+Xd8EpCMer1rzykd1c84WueMCNz0ZsH51hEJwbDt00mAaKFMh2
lpMHkis9R+UwBmLvi3oZ9rOA/Y7w/Q7RtunN1UdWJDZ/fu577y+7jSekFBRuTUjVwRP5W8b395gr
iP5d6tOzN9qdK4NeRqT6ATwillwMJd00VTqLT4AZTCk+HsZsAyllbGlWOFP+0pVxKarzc3Jaa8LT
rfAfHHri7MQlTgpnQ2UxcKbVhsB38dIAgrgvgwrssjYyag4VP4nkWRiPwSIdXXbs+Aa1BU8ikvrG
3CS6EvGU2aqc96VqVAjqc8PQQbQ+Xftaj1rB3TcMwgkIa1LKj6/U1UhhbVlpJx3sETG727Y/LJKS
OIKgMwBb/9O6Rxg1fSOksUdy1L0WY8106iPs/CMOw4ykgaUh9Q5bLm9JW4XTVEl/7q8DMRhQFgvn
aaQlLYodaH68wSNDFpGClyMWt1F8jT3bklzPAXhJ8kC0dDvZCL2y57QkeqS3jVEpmoxqjSZxJRyq
f2yJiZhNofJgzGN4l3rqFr8JuHsrzIuMFLQ0nt5rwgc6Q0GPfCsL1Z2OTE1K3PC1MWOojNnV9dgP
Uj7dY2k41Yv33S1LIp7Qn0lKDJC/fR5isECx4RjwT993XVRYUieIGG6fcdjsB/26B5io+2dJqBGJ
aVYnOPemGCbQT2STmyJpLMQ6E6yfLz2osmcWxqZ+umavwtalNF44q8A93PLe2fWZ1FT3Aqti1XYa
kDAaYqwUsrNt0iYHpQ4j1xsakxl1RcteZ7EiXM9JXkMsNSi6fDUVAjJ32zVSBdfPr4L/9pEQ2fk3
V35Bjnm3Xcy3vg82bVqnHKFRq1E/BFoXA6hidH89+owUazq1yukIPPic8bYnno5qAJC8y3N/2s7M
7xJJcJJtA7NHDWdcpMaSKGTJq4/lIk4WAwkpDm/4Oqt7vVBamt2xqh4pu3rKbSQVtIHXSq6psK5T
i8L0b4aeIVaSvDrRFVngSmteFnjvOxqeMr/sJpQK+CpivVt0KAJXG1wT2XQ9czCCGjuzJcf9bkXS
pJh0MGR41kxpaKegEnMBLFvWeInsSGo8UjemzJwzG17qOisHC4u0ggsh2qweSDfL8phUX8sJIvVI
h3MjVcH26FWiYfRPCtA8C13b9D7FXHU6yTct+eH4+pzX8tx5WQ7nbZ3xNmGXhpkjG0HQ7IGFCuIV
lKT/v7pFo+q47lb3yWY2FToOlfB5urSUzobBI+oTxmXYRb6kGWetO/VQbpnCEw8K9sOKTSa9OmLz
UIzVnhUqqpQJnovAu/md4nBhaq/fWcu9p/4txqOP2A/NiAoFYbCjKKH1thx8Ns/7Ig1MSqbGx696
64S2XPfg/caczYYLLJpuj/5qkRoq1qBMf1ZjmREihSw1RKy99m+F8XiO9DfSGjO0L7aqZfcmmNcQ
VloHiXWRSqynjNCP3iWdGriuagAN8Vo1iDOCz3TwHq+nmMMhP09XNlg+xaegS8V1HBhg1A79ks0K
0qklmbeB9RU6FnZmGYFV9vTzHmBQO84DzkyOYhqZjyeO3Bx2gKvivGQZQT5MaVZuiPRpXcCzHdC7
Hi93BWdhw+hbKvJJ3wmgAn5JgpY7H6WTaaYkoN0FoHWsBafcda7+nULkwb+JwkDG3wmmptcUyjCd
cGmk6VO6QVXeaKMva6eZ4Qge3OCWcu2JpzupQE93/fGZ2VJbbFf99PNailluf+Bgh6NUwZZWXiQ1
hGr7oWr8ddc/kkGS9FMGXLLInFsdGnAsLyQ+XzU4DCC6Ld7EmHZooBLpWBBnV1asywbxjaFXVrrt
m1U8E/3UVpm6UcSUf4f08e0LOFleSPVnp4zLEHYZCdAA3geUWhONE9J7Fk/56R5HiG/EpHIaqzya
Fn2avZdWN/S2hZXe2kZYccsn+Y/aoRaXcqOOFOJBvCgirZGo4BPw5znuN8er+NS7qhcVsc5JaqN5
R9TM0Fh5kLFEy/5Q50wMdTyaFbi1al81XX5ytUgCPC3is1Ro2aU6KXMcAK6JocxXsHAfgWSH9qne
4e7bBNS1QCUNcfFS5e+Y1NC45+B437mHsYQrmdBkRxDdBz7a7qb7lGMfB3uAm+pkzGcKqqmFUBlp
TzBOCHPWAP6b22hssH+JkcirJRsrJamlZnP9k+MwzqWS8KMa4BW/qa0RDEiVMMZgsyc2Mma/g9T3
G9OdRRdanygoOR4fnnzZtLk+ey6xRqHxUeoWJQc2EIzIJE3YKRmAN7WC+LCba+pqSpJsBh9Px2OP
HctmWb5kAbQRR5CHxRrHye7lyQEJZNPs5MaIz3rHcU1ZVc/0Y9ZVBC2snGflAhxogHkBpO7Q1kHh
kRXAOj9b3muFfhfl2dlGyIe2EkIAiINYmvCd2sJJr7iFwcB8P0BitM4U1CjMQqu1DAtX6dCEO9jp
Mf/RSE15VB7YKyjVIOvrVdiHioHtAckGkpCkXcotw0J9UtgqFJHADic8TkFyxFkKptnfAlwvi8HL
bwWanW/fDKuKaeZYdjvuuM7+7K1Pmu/eo+1lPN9lpKTfIwCqvh2PQRLG9ljw0Ppx/ooVFUHVjvCo
yDmvAIgiIxkA1DxHrUItEAAgcnGDP+j8vFVDYOculjO62gpfyDD9lVrIj+OIZ/EWGP/F2Vjlumak
YfZamMFRlIHmmp4HUgZW5FjXiuAk5W2LAxE/Pqjej9hb/VBVSjc6X/3IgdbUWyycSVj54pRZ5Uo3
tP2YuA44s6mIvbvlTRro64FiSUIZHh+jjMaDs81NCmvMpH48Z7y5Q+e1jDTLG2oNnWMZyp0CRMv/
XjNjF8posPgnJ9fWDmY5+moHhMxF/u5DwQernkx6qxgpRT18e6+37DOoctQRllEjzLYHtGJuiYdY
3pbaKgTFQSlt8sqpEq++PsMD2Sn3it3pyH4ZhypTeskx170HqFDfKsseXwqyS/VjONGO+GIHqnLH
oYDG14HKi3GThw5T7QEDbq0rb1fT/IGbE/dZ+65X1ieascjpykbl1N0hyc4D8Iw5YM3HZln3+n1a
2J7uLGwqyyd40vR+rtetx3oVOPcbs1BdBGHUcygPObVrM62DMjPZojPPeiFDotaRDihArd4qE6Vj
acmTMvKX7z0CKHM6fx5TNEXv9IQrDzbg6xfstckJ+rKhz8OmO+HiRfoUW/4YVqHgDhdAtPBF6RbE
by4V2XDVSt+0ZIDzbR6q+ojWk6rDPObdD970jODDHmdW1J0+5+2L6Hrz+zcfTLuZIE8ueXSzeP7r
AuTCrNbVlOkvGHmSl1xqV89l5hRSXdgPdJ9YJIWfjkC3hzeyWwgw9Lfm0vxWQ/uth/8LVuEXBZSw
Rvetx8YL0EucYOQRIIoZx9Zhquo1zvE3L40e+ozmOw4XQWGpZa6RtyeWhJp+TSC+OB+A4wsc5Tdq
lJPKJ5R6RKNsuSGBhFWk95nROWlvSDU0E9GW19eTcAb/qiWnygUOqgJcYedIciV1CE3eQU2AejRr
FP1o9dx2P95LgIqhHbdimn3A/lg4AbBuxqcDBJTWpVnQ02m4VXaZC4AUngJv6fOn/i7b1olpFOg0
U6M1uzTpAwReeTXtFwNub915VygDwmm4W25KKAzmN4ThLeZ5x2FfUxkpD6lgoMqiDj2WAfk2kHbj
Jt9x8Rj/ZNBkE0TwZIh2saXO3MlKDUQn+P3mczjf0sMgecGBan+pNO4exPHLiwu2TmEjNM1DJaLM
uL+MYXSpLpBcAc4WGnvkRN7S0Gwy/5QbhHSFWY+RSyNwLR55RonMpgn4WOBx3/v6ix+QTytFUV47
I/27F6SBNPEXc4aNMF/7sVyKi5tJP8Hv9S4T3XMpWJN7o7tQqzYFIYTtmFE318tlbBuaWPil712G
YjAKT2TB5/vKNVqvQ2BYC6+wGNoG17aPr82az9/WLkEAPeVPC2MB1/LcnjlwfHcuB3EaLYQL+Uzc
ZtnboPP4R6uO7voVoSitFs2Ib+jaVDT2zELPq+XqrS/0sexD4pme0LBFanV0g4iQrOSbKgcHM39i
6+Y7BhLlkYW2G09qYfBmoxuYN7kOjiEzRCbArAIhQAv64eZejO3Nh+Ks7giQntlmLOVWAT8yYzqT
xOgLMk1DfXf7ezlCgxQaWC22t9Hc+InEjjdKMAY40InXFc6iLFanxAomoc5P0BKDCvRiLkk21k9E
8oOXxVu+Rvv/Jh+sPumMcarppekOOfHXMOCbVQ61LPUVyG4iIPz7sN01qKosTSHqMadmU2dty0JR
xu5bNL9DwDYlwSPc7pcYD9ja4ECIc2h+OMsrM4v2Us+m4WkeRFIBodVq03RFuUMWGsmPDCyVtvBT
5cbG/I7IdEWRCBUfYRwrdLET1TrZjgahveK734fMaNIii+Q2iemZ5kU0vhg2XI7RKNUfJK2bFjr/
BxzAaxhtkwbDEHF3XxLCmMcU/YcwyY1Z8A13o1kZt68a2fSc4OepFhmVE/7OGkAHd75K3k9AimyR
7vmTyRdaaqWO+Yp98PKXT5UBzd7eYRDoOCeMbuoeeL4tah5vJF86+wU2Abj54wb4Jq3KPWJqXOJw
bUsgB6ghJnvhmrBXZLY6FC0guIe/nmhA+leN0mdU/WB6YAHV69enx7LdfSdY9kYNhYolFNwnBbXO
LHZey6dAcgWawy5bFIraPAo2tbtggRfh76lu2V1cuiez1H79BbAfdcWb2IG7s4yslIlZGXn0CY0V
K2xnegMZ3pMaf2x52zv2to3kw52Qw0mCtwSi3xwHo3m9vTbM7+o545IX9tXZTnrJm203PQLKfadk
P0YJG6+JJZ4q7uEUdDyVcrmcWFybqkHM9qnivb7W0BSGJD/ylNNOC72vwRWX5YsLWUH9v0sJaBqU
R+AKfyWHNdNwRu/EHxyqXurNaIlD0k60It+VtGpLXbvFazxdvI4auVFjbWQVhyjRlXgNfTri3NJH
FpVPpjt5nYJuw2rtoP9/hJ1Koo+YEp6Src+IpEFjagSljhuTJ233bmz004kPzC5BD6z6xJm94iGI
1QL+9toPxWcd3ADGPClIouwNXXZ1QMkmNN6SDUeEvcEfJbBh/dIqd0LmrMoPLl7e+3eQq7fDdbez
mxBKT2+K/2nvNlm35iqRojwFZdknXqf4t79w4pmay3CAF8zK+HVqYw++bY0osF5taHLmMjQWVp1Z
jACTOM1gCe+vD/KI2R0lOkpm7y6Mqo9HGcrWwn5RrIpeY5GL++w2iBHzQU3EfrxqnLdoJkD/mO9w
dPLvvwwsrpY0djihp6TMefXqHTDsgDPxTJ8IMJj4pnwcU8CZNqqdjTWlS48K6c91w0eG3b70bHzS
TYCBb6EejQeLRT+2mCxsHHgLJSzbyl68xoOPi0YwC09WEpNulPRcV0/qT7LPCgaO+dOWQLlKlOCw
ZmbfuziKByKWOln60z3T9tNwnZGnMDanScnVlntqCaa16P4oz6blkaAaDOi3zt8l6/2seXoJvonR
yJuE0EpQuqRcnGFUuGmGYmNPnXsk4zss3alBpikgsoLuDp8LyzsHaKXqVoUnFN4p8FHM0/DU06n8
oC4VD99WRqh824dMXt5hBsSowgXjNH4hzLkhoCF/BXranpOx05I1OxGghasia46BZ4fI+cPjxmXy
lxNss20REfbG1WcfQPPz3vZEdAgMy1i/miTQbJ11SiiqMgs6FIm+nLEAaNckiew88mqDQrIEVJ9S
iRNbFZYkKEQN+S3min2MUMrqekDvqPF4treXe+JMb0GMT9dks+2Ebw8tDwMUKKBrAdhBddtWvqTY
qH9Uk63W5xN6BF0rOxEpkJ/z4UKo79GNkd/53SahkfUjW1Qd9UEW4Yh+HNznLlTsWEGBbZqYP5EE
XCC6pIOMD/botdw5hFmR6yFa37c+/F6yUnzpjRxf9yLBXR32uYuQC1sRb4DDFr03WP9sbRgoyvqt
Jnovei6b5+OrsIczLKHmqnBnGm7z70Kw67sRSV3TOtMy8I0DxMPd8705lo5opW+EGl/T/WZZzpsf
DUWDxckfvuB3tGzZM+b4qCeO6ZxyOsZ6ol2zitUi3/hMBPz2AE6d+dWudFLH/NH70NIIt5ZCxovO
K36tL/iIdF31CXU4lelvyJTzyzdgie+HrSJhgSRhOHbW0IDDyNMhWUn6zlQA5kBSNs27CvFVKWiN
6+1CZjG3mCexhCPjVlTViguH5mlw3sq+tK+oIrq2IuR6RJmIn/lkepe7oz3pVXRwXo3pqkuyx/60
pyDolbWxFv1njCiG6d1stxNspVRA79Milksq+2PeE7gOnaf5OWk0kYDGgC/Qfoh+mPRCv7uV/k5N
D4LFWr2s+XQ3wQgoxWGq9AiEH0nFBFiQ4R/xGZtNzOTLIP4he2dnI3Z0H8t/KIgShmuPn8hG5gcC
I+C6gtZkCZRnw3Qwvtwi8SIRIuNQadYqinp4JpyzvwsFicfbBskzy2eNov6Khk3i+fqYSIYj9rP3
2IBK2eVhJ6UQ0+P2DJEyFTIqw5snxD9sXEFlmWAbx3j11M8D6FiniCd7uSB4LQnJCiK+M+lJfIAs
SUWdVCxg59l/rr2OXZVcs32GMKM62fKkf7bG4NlWrCyFqAWbmTpuRSFdmHPRnbWmAeYZTpo5318R
/miM9V1FaGkUBKkdAF2GBqVgE118QCD7vp6r93YD9i6A5Hp/uNYCtnTaJ5i12/mAsIkF1JjNSIzQ
y6Ko/7TDbD4ehWiCmm4cemtLrB2Apnoe8v2fNnzcN7lHVY68fJEnSoCmwF5Qs8MylUJj0UwEsMdY
uSVs/0NordmwecQW61Ps5NbIFF4Rrip24adKlHeIbFNIZSRfA4sJoTon74izKYPdNBhlb3eFz2Ki
hea2lhpW0SniAssN9s/GecVhqe4oIRWq/uyLhGtS7JZ+vaXSCBvBsFfpHRTx1CExFWpeJ3XDX7Hy
PwRvjGR97UZpGJytKGFLBq5CgfJfJ2sqPz82BQtAB4bJDOvcCDkFvEJrOWKo//8fy6aj0+368ELI
vFA8qIluv/2XNI6Wt5oa/Q3hklKPcjU0wdubrOWztL0v0zC9+REqoZ81o5uOfXmaphhNLlob8+OM
fYmsExSmyT8jECfNgWmArs7MSwkpIjZBR4HU3NrK+43+ar3Zk1sTYP148EbFpHaSydNlQGY9IG9z
4IYCOjtfawf70B0UQCdrlvJWS+B2m8iHM9o/Hs1l6lnj4kAbWZyLkeOxPqb1eJy4HidNRFSVSDWc
J2nzEWxiRRTFoyR/5wzscmK2gyH0zOK0l2WIX5VGFaQKaEpriZ6CsFSJzL9m9marzPxoXohB0E14
Jt2/P6Wssrvx54V/G/2/tWCCS11HUjTssF4xD2fGMGa0qX4OGRJrvvZsZOqFgLAy8ayQUbRG2xK2
QNEf9uJI4xVdsbhR4t+lcNXNFpv7iANAAMWoJW61+rpHPhGzSqFoopILEBX3J9mBEQ6diq1H2K5+
airGLuBHBzIma5F3UD4InYPVuvioPBhispZZq/GIBpczSIkb66sx3LyzNA0hZCZnOBfUFMlLHn9Q
fSxH0UwGmyU/SZv5aF0lFzAdusKrJx4TmoW874oDGZ6dRdp+SXGSihZmGyvtlwBHmoufDhOCcMwP
wMuZJrZ1nQuWS2Z8U+IVip6uMF+6sxENATF9IpLuFUivEVP+RDSgjFrS/B+DZkuINFJuCB634hSr
qepbIUJJhsRhbqCAZGaJ6KAhMpMl+0Qnv0XV7DGTYhFIuRQohGc8mB2GB+Ls+syq8JLuph2DXhlA
LCScilz1ocrOU8JlRsC/J/DfftVbq4bEasbaMG+LGQoj1ndQZyS7G0LtJy/3InNAk/wn9v0CfYWQ
zIgLa1SH+4BB/AKd9AO6h39sqU5vJtUc+aHh9pSpdbry1EqIkFM0MzZiW5vl6lRlFuLDsckNl3tL
om9VBjDfc7/HAIwMJc3LpQbtHSLx8gzInrLrkrs7esQLkznlPCjcU5vGM/1jt2ByrshBoYZQD50B
eEIOe0th3Qfl1eAy3jCWxTnmVQ+JY5dB3hbG6jtuDAt52YKXN9S4u7obzXz5PZtsywMyu7j/mWQR
qneFCDS2ZSy8o5otvaSYC/UNRxW8jkerJUF9L7dfSQYDCU4NCJ4X7dX8+PMgm7rwEBeSiGKitIky
xPvIULbKgkDx+fS4NsOsVgJ/2+KRvAEfLzSFsDAtzqTn/QsJ7fpKt0pWyqXXn0DsHjd3cpeNdxXt
yaWvbH0HZ+WktqfeZdMBPCEEtF8FOxFBnycpSfbB4DxzVM2YpCwsVpjSLzXfDG3nO1c4hrSUK3lL
kthIyXl11mgtKya1i6jH2YKlz6ktg8L7s7Rw+DgsaSKCGCsIpa+50nAALG4WqNttpfCzkuAh4aTd
5658Gw4+6OiKwRsuXbnzxVavRCLRRgYj89NPDkKHIVzXy5jqY89OQYwezVp3fMqdkIocKCJYMeD+
ZJ4SjHAbcDRZeQcTuQziD4Wev4Mt0WO1g3J1wzd71guqx7mtBnl+yJuzeogoDLHPG91bdF/L/SWX
7sgpbuDjpq5cU/QUy0J/XcxsmUgdVxX5GeuuHtFOtJqis5hMy5oTqTSnLlNjL7zpndPGLtKlksQi
k+F5kD4CZobadB4nw4y3tCZ77k2jLWOF1QPAAN0hdsOIOlS0ipBXA0a/FtvLvjHYzmdkoU1MXcEj
Jm3xDyP9ui4yBkkj24hFdjGHX3d/vjTbJFWT+PFowuwTFXN+p1zJDrktZMxz/qyme6Q6RdCQRTXc
i/Al2A1jBaEx9m+soEnMJbZbmPrWD9IK/pZmhkkmNEqZOC+0cvEKMalajRxPTq/8DQIqwxaYCQF+
G9K6GMoLieRoJ7v4ob/DTWm4KYHQ31RndZSLtMMocbxddu3wb6iacykmCQVELcwRK1MuExUjvS8W
LNDJv68U1Xbb6RWmLSg+n8U7D6V+1tFJ3Dyxb8J8ccA2QbG7knCbDq0Z0I5UuQAPdrv9TVnY1lT9
pu/0eyazSlwImz3uzIEz533DIGBJkqrQYrCDTllnEZ1bt5+xiemIusY5+YQ55l9TkDwJhKB7kvDf
VsjiSRPIcAjQrZ1igS8UsY6KJYwYz0iNG7h4LQ3jelsKoI/rP2+JHc7VeFA5hmCGdV0Eqwk9R7Sf
qkc/kEKgGuEtYCxh43Ot4EBshodakbFTN+uY8aMTuCkVKc/92gGrCzN6SIAI0i/2K+WgiOVJhMkj
Bvwi1OYb6YMXDf5rM4PgeXLCXwlP2dkiNmfTBdDnl01a2xbdzCN+VQiiQz9135T1lNMohYYvHIxh
BlOfSLG82b5Sqn+4izQVc2XuphXVtkCPPhI2zLmkh/lgj+rdQI7EbYHS7LuxcPQY3hHaq2V4BcDL
pkQcvVfRiRuWyjJ7pe3AOCiQH+PbqX/SS9Z9T5ftaItGG44KVB+YXsV1zg/cY0lAqIk1nBjYQzfm
JldXIU2TlB5Y2NLwykZ9hqpR8ObUjxD3RZAVgvSpe6KazfMOLUtpBh45RONksjx6TyKxsvRXd6Tk
0UEsXJL1U06CgWwFWTqTXIbkG5IwK0Rexr0gEdxSa3N1myfXuow8S/gP4Toj+YnwP5iGqjQbN7s9
m0oVO+EfnRRNZzlnXejavfnEyABXlb3j5s0YhsTc9ETmaruzwR1J9rpvEenm36sUhxYfFdJQJoRt
GrF5jWhPhCNyV4vOaMRRgETpmZTlu0HccuBjAQsvf0mZk4ZdjBGpCbZrNus58vkzlNZqPoB2i1PY
GOpsfThtyKDQtnuIUu2UZe7/tjtlH0ewr6SWLuzTWQiF0i1RjGpgiiZdrnftPEtN6JKGa+1beqmD
xVeanVoofrhKaoIV6yaorZlnb0gT62sBRocFDP1GW4GmmHX/musPpLM8x5WjTNdWB/sTvkL8Uo1V
qReVUmHJuS04sslfxqGRD/+ILhkjkUa8G7BBlgF0jUAEF7pkNoYKrAswbQkZWgrMcH1YHT7691eq
fm2jAUBE+A9jNXbqaEhucmny8o+h0eYiZ3LMcEVk9mxcgfW6jtJbRnVq/QOzTAWhSgDNfUiL0d+s
bpc6jWUW2cn4x3jZ2i3G0WCjhX/8jlC/iuU/MihCn90yS43fFzAyYPqz8f/Jf+yZK81tpzHJBjN+
wtmaPzYgpyfj4zFmKOY/z7z0+rrrz2jnPgnyqbaKV2ZV1MRWwlNQKn7Udzleo4JGGTMQoAENq8va
apLdEkk6teV0asFg4zFT2b375gUIWz5qqBkTpUK/EGT0lKoBjOveY0oxxSiNH61EWYBjUbRu+H06
8KXQ5qvEVIo5q4TQgZLPT79EIp/fXISCKOg4vdhmaj0BdqnmlEcvjnIDkFiLcHh8bwnF6+gkm7iS
baqPoUl5+F4pTs9Eb+5Xv42Ey2nTONfDKMI5C3Sb8qLvcNQSF3iQ9HS0Y8MEK1r0vt5ztmoM8++s
S6wX3/j0PjCdJka1PbN7BD//XZsf7c9r2jxNqBLslf0ybKbrT49VJB5jRntvo7P5G2zoGIbF69pN
I9oLxmd1/35rI+97Rt/ajXFBD7w35ewFd0gPMb+sF59dJPHuxpQRJSZfHDoRkouQeyYV6nlBII4j
vm688Vt9TmMW6LG1URAjZdNLhG00vwDD202RHD+gWySKSdhCxTYYqR/jYEZF0+ME06vf0ddwH4s3
R6dV0zpOmPfvwEx4KL0Hb8YLMQkuHB3ALmjsF4Rvm+OIip/7onDMugquso2m12JJ5KHXfzpfNDOe
5lZo6D6RrnTTG5rx8+imo/QJFEFlvzoowprMHHqpzYo/6e5CW9pTSKhZm2wYPDEtFFcwJvPdB/v2
l0Pzc1D5Scn4CuneJT5ZwO1QwFIGzGQKgkpOlMYMdm2qpA+Dz3icwrDmC5/AVvT3R3pve0b7Qi2r
osRZOT5koACy3Ha38EgPszfbUYWsBu36P5JhXFmElVUZ5CVnkimvBmfewsjMl2gsEB78sFhC9EqI
YPzF2C+i/syDWz/YW1rTGHO9fU7dSpty9EejJfi/VOZzXCKvftgL/i4xAZmfxIMtim44M8duNPbF
OE5O9MHZq2sdJtlTJx5S71+qAOjR11HJCeZ3/juQoPoiWYqj/z9oF0LeOU4Xb5ohmGntqqovj4v8
bUZrz9EMLhfgLmFXFDK+70PYWpBvZ3zy91x8jbRV/sK7QPkYnL8HAb393Ym6GwVkNvDUXYBLe4OW
2cDw+RFfc9fRH7MRIaNpGL564nnknNEr4pDmNDv2nx0RlGbdP85OOtVAe3vbEziblwquHMZO02K1
+2uNKDubkhKSdLN+xBJ5DplUTPpH/ryO6A5cwXcaz9WNh+2NPDiUR4//H+szEnBKT8L+1V27Udxs
ESesmbm6Z8lsJovu67RUkrO2Qx1O3xMKvoLfNCTofuKcLJi2VjAcqeTlKUQui1P01FHX6/QqTsEZ
lTm8rLXWtR4ZNJV6Jm3zjUP1+Pb4YlOdh86CB92p8U2M0Zf8I3pYQlKSrtsWCRekQpvrFEiciqC3
q1BXJGcHyCsbsWbQ1yFUTzpsbUuKuNC9JeWgF+ezYjhyHtctNnHofIIdeYLHAkwQBMs0a0y+f5IR
2nmtBE9tN5VcrNL8gZOi068HxJcFmVWD5S1rAvShHz7I9aflen0+MYkF7WaX6NlBdVIiJ16bfgXT
sE+jOYieyoS4oolwACo7p+nuPDH5aAvBuo6tqhwrXaVtP1Glf+9I15WT7dAFDWXUlh7dlRfsPx+P
/OqGyt/CITH1B7IzlKlgV29ix9yAjpdifkAH+QPPxUim7JWd2Z9ul7VY5LoyZuDfiAo6f9aEqqHr
Zwh7vGs0djRGlQYh685knYRvM9Sy71NC9151aTKXrkf8mwcLGaftyX6UzClFNPgiRnVSddONoip4
Rid2ViHpXRys5uRD7TP5Ub/Lqi1rpXfijqaK3a09TyjYyDEt4Dp9/5/JhYPVJ/ts6OSZ3XlIrOll
C9vqZ6MemlBj4nVay3UdFvEvriMblf5QgQXSODib2rYMEpuCZ2Oi2ggP9IUMVtAbvegL0MKuxWuG
A1lyVEjnEH5dwsuLw8piFQou7G3xwdmU1yYI+PaqHJ3DfkdoXmzVEQG05JMbx1sa/oZwN9vcEwEX
dfWWmhSJ0UYrj0zXAdJ8UXqFt/5Ievqt4EFbYCYlyvx9/Pd7cVgqh3X0KvK0x3s1Dgqvgk5R0uWR
/6mizMrz//LtwOufvovIpELzMe4yh7kZA4AmS1rJeZqTnHGSpWq3Itp8WszCVK2ej8Qa58ZepAi2
LvBjF5a+4pynxH/5VWdmDe/MnhcApaD724mF6HrqCcKHWOx+NlPwwrkOGykQEIIT0NSPa7rD8ouY
1TBuqCaPFfEbCYvBy2HyfRn7jzKY38h/IS1Asb1F4H9wnvcgpOchclkjj0K8Da1Kvz3K1reSO1Sp
jZak0XvVL9XBbYj9EipSe7TvN+TI8B2hZAnDC69VxzO9Z67uBuwJD/3XrejJYsHfgiv/MIFxfoMO
s7LS4kdlxkPJSe11gt+Op7aN7GCl7BIV6UJ3Jrl6kxgnaha5n2zJSkzTIb3V+sbH/5D3MSEBKw0Q
pWwK7j3JuFJ5MGWgPmjaZllAd60vUYpBfxbUEGw1A+9BCsPbmIwXM2prIrfTicGgyzv5yGloDe/A
J+L1wL6Wni6GHXCCEUyYurgv8nyqL+eFNHily9c6VSrojrVWD+f8ZWp34Rio3WMJILRDzmdAnhgK
Bva+ZKAtS6KuYzr4GNq2D08DzjfC5c6XnVJaO96COnICHzrVzF/1lZySrv44fYYnhq4SwWh6fD7a
cQgTiIriPQv88cxX/omkjFMP1TqBHrMp4ZUunXVRtjdSYWACBsip7fqqvGoYPda0J/kq8JgT7yPg
dSSe8tgduF2KyJnXOcL9UmHEc4ns2izYLL9hD6N3eBmW/idulWWGreGYOFIfwQcZ5yIf4bCTCiTo
HKoN4qPi53p74/via0ovr/HQ1xbiRHiU37vu9Q4w5cm7/bsNYlqOMn9xvtBqW8aNPpgpvVTc890w
2CeBKB4tNi5XnfKs5cwe4xcUU9NpUUyuoujh9rQcKZxinE49HW6Ivuwi6yD24WWrMriYxpqf+sLH
oa00YfGRNSwbx3zWk9yh/nc9Z0p/ovS/kguisXw0rZnzY+YM7VCWRgbu8PFNR91AZnQGtZ2Qwcuc
ZUnDndDvsq8TXbqpdi4GXzWh6zp71zX60baklVXHKIklS6z2+gch3C+/3ZyRnjy5F0cIXQn6psLL
ycOULZQXL5jwSX0kGxE0kRPFb94vLVSzGLpa/2wpZTRrgzm5EaD9lGrpqJIJlCCMslmKN2SYrdXB
HYcdzEDt+6dPglUa/pY8UAYYSByFwFGO4NJJ92hqRIAjAOgYFg8R6x0dyeq1U4/YJZheGfcX8d+c
WWswWKhScdmblvLT5iTCStBU3/TeC4MLLgc9ohcZrHbU6N+56y0Zp2ly/bNJw2Z1PL6i/01I9jyC
Tlh6V5m5XjYv1kUMJ8oJMSrESL/c5l0gLinP9iSpMStqIkgCjpRg19qvIEXiewoE4BkU8l1r09ns
zIBoNUepCtpm3JvOvXrb+DK+d2Wf8WdazpIsPOE5kH8TaBDGqfRbK8ErEuL93AVyrT+8HmHYrgw8
ZTulhFgX6GPSLEJ+bQZwDKgayCmPKcNfoIlAENxE4A5VUSmNf+2oeuKRqDOYJkcpFAMaMM4L6Qhm
GQJIR8D50sJf9NIt5nOtcAWN2p0g4pFI9J15/kYKhLuW0WWoi4IfDqhiUZVtOTnb4PCtfcNZPpvP
hQOWA1XiywN8tiXPXbFG9PyzKohdctdssBbDEa8Z1yOflVOpKF/t51T/+dyYfm8LidtcgN5JmKkN
VJDIKnUte2R58AIGWWqJjvnKkZNu4kt2bAZhLePa94g6C6yvpmKjD+syxPwbHH7Qy85ePV8MKMVn
WwaZPVTPTUetfxPEbm4kS8Osh+qh+BHuZyOUK4aHmMU1tzPBli+94TEFX/GI+eyB5WlmjTrUI4iV
woLLjdS35V557lyFh1XJM4dq3skvQbZC2pVyBj4nKEsoGftIyuLgr6s+dAOmGDsEQjNZ/aypo14n
7fnIeh+b+zt/guYGk3hwD/mGltlGBmsqi26uimuKhMc0ii2aQ2d3CXYYxLVFdS2x+/pvt6bnS8Ah
Le0TgYNviaSweWxytzbM7PJZjjyUQtt5Oi/izuWfLHkXlNGdFCnafx/wXU40rxMRFW8dnxeVEKau
fbyueXueZZEqLiHsZU1olxD84hdZkNx1YzLtzcmqJpYuhVOmSYtKSXQz9PY0rJoGg9HnC2DyS9d1
V+98w4mpR6rCTm1XKwvMkMuBa+uwZhLvbVFx6zIhktKQiRZ05YwStcM1dxpK+Lmdxx3PKeaQo7oN
IGRRpjM+f8+31TmIA4vSknsq1gJSw69a7LpBEzvFJpAKKyVXwyeIMfCHElIxboPrLDNGHDGsScsL
N7I/Y+q/NUAZOvPUzFcT2FR2XEMWnggJ3cDR+xLHcylRXOV8FgYT2qaAqAIA+G1p3GUOrtJl2fYy
HIxAlWD4TMTGNzKJyKRUh9Q/IpOkki5tcSY+k2/VYkvDVlvKkpcHjwt35HIEfFVfED8jtLjr0So0
w45daKGOdJxjNd5aqJMsbAT6Efq3iTrhMUr4ij88+MlfoEqZ7XqpZAJpzCF3JSCKxUImuk0mShp/
Bp7UFem7LVt/rSKWinMx5Uxbn0Ey0YRwSG5PMwKE2oSzhV++BokYR6iWOgLgIQine+569DCyhlmU
aogKMaqTGJRit1qwRDoEwoNfvqvgKG/RjbhfiiZ8Jnrsv8Bmdxa3Gm6qfUDC6B/iCDnCQgbaqzTP
qPi+S9GzySgH/ph7VEHqWcILr85Gvd1GFfBy1wPkl35QHMZvsD8v7MgICHMux8kkO8fNp1KbSQ0r
Z/brG4rjcRDqZW9A2MoPEU5Lm7kCwr4BuQN8cOJyuNATJjXafcdiPNLdG2mL//xaTIYR5U7NkdcF
x/QzYJG6b2W9oWEKEf4BjMiqnj1DTaXJBSh+AiMvK+Qk8xV7wxlKRPNmf8sIIzw+KSPPl051xstT
wY3gfKivY9WMenK+Dzl6VqtNfs7EeShcXm3691coPSJZUfCFZ6II9iZKSIN/qlST3lNt3CVVZzHz
6mR3uvPQaMAQxr73QarR4MCDdaeCyiH36N1UdUPFcDIMovBW5pluewp5/DKL89y9lI1oAaJN8Ufm
zYTwCuk/OyYz267i/46+e4usPNb3EYgJpq7Es6QVkIJLjv327GPc8WHwWavltu4J6UsiDlbJgNZI
Jysv67KKjBAKXybRH8vANK/RP+c7a/g5e4CPoW+msvBkTtU3RnISq53HBP5ZFzeU0QS1t5zYEGFG
8Qb7SeM4H4edDmTS5jcUfQRmarC4pGWI82Yl3udMWHH/DasKg3xTyVtniyUU4irDIR7cZJUQyINX
YAPN6rrfpYrONfahMiXwMSvU8KhASytQdjLxTf41nmNrhYlPQXvHG1lFimLXpJ06UkV8o0qbnNkA
VrcmgkdFgcTQjXOVZZPVhO5OHp+0bUM97kewQlg5YZ3Z/xgL5NOCxr9UvJXacbS3MjAABAHkcO6W
nLAP1/Jp5N3MVTYNq1Z/QHmBkieF/B+6fXixLvHwXZKCGCG7BmlSYz1BCwGuLkOq2PTrcL3FsVV8
s/mEv/7eKi6GkhHpUjqdQQJWixqyZRx4vxnWB43SP2Wb+soWhYawwQlhxsr1lwTtfCAhAwZySP3Z
qZt5iqh+V7gn3wPSVEiT09S6GHusbxGOdN9nMrzG0xvcQZyiYi1LjmqNIvEfQyrh+FBGtKDN7E+g
QGdjGrIf83IZVFhzj+UmH/7veN+RniHrWi6rtSKTGIGyPDzXef0lAQmBa1zaG8L1jjS7Ybc6kaHi
fHE9YcGrwIp6RsQsFxWvlRKMTZykhhwIuiXQjr5sUOErT0xYIgzHVlipRXnQw1ncBx7Pu0iHYrti
n8vGOfdzKkyD56sz7HleOUkNnQcgakx1sZg2fQ76Me1gWBqXXWS1j7UjCgbxlijMhhQ07RnawI8A
HWtIwyH8b/VPdb5x5HdPuV7Zu44C67pPwxdg2ywdwv5qEDOaHxrqgozBxoGz4X4nceGV8NR3hzXw
InxJYKAovjcokQgTaR0nC4KFPplJXma6Y4lGxXPrnpMgXultkwb8RLzMQA2Xfkf7sfrU00+/iTPg
fDrqu/dBwqx6htDVB061MzbocVNgkMK65qb0OIZIH5CPS7+lCIB20nIHVC/iQUPD6mipwIqEIefH
Rzr/7Z4w+P7Dj0PJUIQXftuGr6+cFo9yXA9OS77DXNndE33tgkM3KpbvexeZDaAOlDcDAI3270fD
MxoUArr+Za+Y9AamyTeaWFLkCgQO9TJi5SiXdOOuZ1j6xUVjoQPjrl8kjx+0yir2DK44mYlj45TP
iFpRto5z3H3d5O3dFnLdkK7vIfSoCMLS4Tn7mMUjFgmNOu/iNZMPmp5vBbIWmDoJc/Hs9DMZV2so
6ft2elsUpUGREaHzQ7AQ9NRTugrW2RFhwmzWlEWluLcYS3blEMk3y1XSMHNSpQKN2UYuwYa10VQt
OqVKz5IfN1pOwgaQge98xX7MtKjvyObSlCdE3ZqDnpYXze5rdPEY6PydZknihHkI5hJ53sfP3T75
VtM36m4Q9wxSntbr//xXEIZ8WWERJoJy7ujj9eqZ9RoykJ7OT3FxfrN2FrCURvC7gsOObCuebasJ
qXwkglouN3/F6w8LgABA9jgcrwbqe348loV1o2NcEDAKdiP7X6ATd/E/wvYu5mv0U4MV6xmRPA6b
+Rtb/pnJSKR0kEe6CRcwYekKpklJ/rIQIXmJs/H4Olr6c0Xl3ms/tN8To38N5EPPTge7gdgifYRf
75KXLj43+syheDNl5PVuk9U9jzJBfeuDEkQcBm44Be9GYpBsIJtvhcaSHXisgxD0Ba4aMOlvATeo
3P0T4yv/fjIZKI9YwcdY3EC46LfBZtB6HHlK/lYpZtbUuS7Qc2c6DOdUL8cYNTga12/I4HLtxI8f
6J+JvsbTRbvjSSfCWD5bXarZHMYb0P9DfD/DA6ckhKBoHezzNlsy0hDAkARJ2c9H5cHAnvzH0ARf
hacyVy3W31qwMYhYtke6iOHHqqOxe64G+3me2LrbwguhswMSG6hpyXIFw/hcicqoydl3tqC3IK9p
mCQKZz5Fpyifkd112C9i1yiSoayYLIZ5gBMFk5JAHXbS/81pe2wtcnRtqzU8jKZq4+9iXYoHmPKx
Yh3mmSRUneL/odcWOYh2qaNeHriBAQd7hyIhuEs6arS1sk/qrKw8xfBZpjbj7u0CPfUBWH6MBZ6D
aZWLkr7z0zq5utLCZEHxYotUUkihz6L11OJuuJKHBRquGmg/LxF0EGg7lrC4pBd2CqomBZJ1T4mV
cmrEV3RGeq/J7tkCdGdd54R7FeY+/qHMTkv2payiJOJ7LiGKr6KJNMI3Bgz1GjYgK6+Kn67KUxKk
NNoxkezl6Ga+08rG/EZdpm7co2BUlypBveAgXN2ZPxhM44Axhb3C7Yf4S3NW1eK4Hti4fp8rTxTu
I3WJRZmRgXnoRX5ocm4fUieMgecmc93ZVeNpJJknxUQ+yKXHFouFuz4jiSKjQo5IoxGPCSx2s5+M
Td2u9ezb79LQuv03x4GOL35UaCWFF+9cEZFa6VPyz7f62qczIQ14LbGVH2M05Siv7hi6SpfuLfFQ
q3YWIr0yiMXySVOGeKYMrRpc85TQ5LAQe+gQ1pZRzRK0gCsY9ncPT7f5+qyJyqzFYFl7hGnuef2u
j4uYQED5mu/JAQIlRNKyHdMhMq5oGpBac8qOuf12K0JgrxUJesZy7999c8YNUYI4rBTuGwr3A8Ge
BZ6kIfFggO8Lpf2UB0uWNIBkUUjwcYmLTrhAx8pEalT0kzjA21yl8+kaPExG6wzimsns+KnHdFal
Z2ryylNkCHMh8lQYCrtnLpXMhKflDMWoyow7goz+jhBLcPo6KFFuAOOKCX9Bo2FN5bpZt1M0Qtfz
7oclL5NhPgtRbydmHjFqautYoeOQpcKnHlb5QBNJROH8IHtbOEKA4rAq3hF38zbRoRhwuGrhuLt6
qQjkOug5a8Qb2LuzVB8E5XA39zhc1FMQZWShibn7ULrVdifEfoSGWkyyL4VaCm6ES/+2HWAymQ/a
mtIIx6Q83iZ/WKspS8JCqirs9+YNVY7y2jeATyU8qdTgx4qmMM08sPVcqLYh+bh6ZJoX5a/ZXDmb
qtNldRKjMk01bNJnElwAjjDChPher4pTQ9UEp/fnu7qY3XWVv6QznTXjRImK6C2HWpso/6sfgeVE
aNSYWZAGAlwLmxa2NAezhsGmU2E23K8dBMVmZ0w5KdeWVwLRDbH/zrSvdTyQdXxTI9IQuN6l8HQu
u5DAbW+4lNtEzvEydBVHlOqTKbykPLp/7pJ7BBjHCVS97tAvy/uY675RayaWIHBrgwuTb0ArcVqF
eQX9uDZM4arccSWZdWgci0Z2r9//rdmoWqYr68+cXUbFlKfJAb6xp9HBwurDzL5DzeoHUSUzovdS
xhUzQZblI1p09D9SAJhwMVmVpoipP9LPQH9QSODU8fSxTZ1F+pbxcBFwAwKA5yWU/BCIEWEfv44d
Jzhyd6ST4wDNi0sS4An6GgdTU0PHOT2ZX+xGRRNDpPa3VSOjTbhfZmmzlaFaGA3nSEyJ3VDm6eS7
UFdao3AQlNyUsGBfLTdR0o2Iok9UeJAIEH8Apza2ZnY7137fqMqtc1Turq9RyL2vWmsWOGGBwGjg
3NvFFcy9YIRgwKC74JSYr2JlsEXRhyqfTv9jJf/FvsQwPm1WblIkvjZ6RNXjpISzMLq+qaRYvajI
DcT6uyf4mKPynk1XscXjsGE5RBxNlNwTxzoxa8Y5vWuNbfFuNjN4qvzBbgZ8MlGYgybhPY2AVY9X
KDP49t0KWsm/tUGlww2JMh9LHSnu2MBCSPBtMm7r+Xh1lkFfG4Bi7DxkG/ExCAa9u/tym0bMD1Pp
Y9mOsTqkdXTI/ZN+XDMoUutWzid24788GVgHR1NvkkOa5qlKgox62SBS1415X7yUhZ/6OgdpILOv
S4JOUGUPakcwEJCSY4M9jUWAZzYisaGP8Q7m5uBCrEpFsrxpSPPOHVhK8x5T8Wd2eqcuKvJI+Rgn
dlV8I8GOmnMjZUiXlzzn9/pVf1q8qV7Bvpw25UasSdeRZcaq37D8E4b1MxiplK6Ez8jv9gylbhc0
zuII1CjI1nLWDVufCw7B0zP8EpxcAWgNIVj0P/bJcxcENWkdmsNkhueEUsEcmO0vEg1b8HZBF88t
VjXS0C7tq8Q06kV9jqRDLIndXgWslsJuc1l9F7tnXdf8lUBBWQFllmXcsyjRHLAmq/fxJ7aBqE7g
KzfbGeWsYngFXKhsdPe+eqBkR+S9Z6jDcUHmnm68Q25Rk7Uf+/lQxeA0yU5+zYx6UXuFBakyfdg2
9w0tkIl6boBUCmplN01IxxHXSijHR0ZIjmiP5rqMWMURpViFZsRxuuo5AseitZ9tirjFb+eSH/Bh
+VYCV1MxSfFgOtPnbA2fwG3yOp/Y15/wokxNhyunPbYLOqAtDB6s85XhrhcCwE0PLM5/aZZRWuZf
l89Nwlpp7zQ6CIXxDHHYourDvlCdYbMfc0B2mk+SKY4nIJNrvyVWJTjKPlpEKlKrQzpEdsbB1UQf
zytJalVU7tfPHmPzBB5fmxmeODKYj1zOlS5XEcY57hestpn2JiqZw07R9H0c9BUmPsfe5J0/Jwtv
vAeAW3CDBqGnBDBC5tJIrO8ko4hxG7I2MEkchqhR1taddXjGcEDL9Sko6k6/0EVuHWy6m8c/waZS
AT59IqkHBMpS//DnMld7/qIxqxA37CzwlhuYj4u/NciuRZ2IA7yDF2UIyBIRYW1//uq8YrngbwVR
S0VZs5I2ZBK589n3hHtd33AjEuzPpgfXaNFQ27Ex4TOYqp/6vL1sxwHpr2CzeHbkLtjSirLTgFyN
y8PVrlI69CVi4YYA5fAU6L55ECtEbAE4p2lh6FHtTRva6XP9mbfKdXTSbjycS5vYYxlqwJRa9APQ
9Zh192u8MXdbctMKkiXHdINtG3NtzoD53NIXHsdMKyPj0rI+H+WwbkW5ybQSsaV4wuMLLSYzawK+
dxZkrECYXZI2kGf6la+AinxA+k9ytah8H2WhweC2ywVZXk1Ae3qgtmI3TxSoScWORx/baEQ7oRG4
2Sei5O1lTDKW0fWqgLTEzeYsAy/m3CLMWFzOJbY8OcxbNbvPbYVpVscLJnzN44GDwBeM+0cg4RC3
KJXZUXR1Cm4Bca0vRhMxfLMD4Afe/Eety7gVr9kygAMlhTmIRayqWI23XEosAA0+vrWTf9lZ/5yj
XM52kYSkVGc5L71O4rxskigapVPwkdhss/bjERuj0PQ3KWR1yJ9xneVJ7KtgHFU+0mAdWKTOQbof
6hCNi/RmxEx19X715GFIOmFkwqPVMxqjpC3M3syMzgCoznu4mVerjhKceZpEFjIgem4Ot/JSEzPe
b8z2KFagi3f5Xf5vt4/bhJPrAG8hzSrgFvw6zmQ4eG3PAhI+J1x9xvjFFtYuMT/2IshGvt4kS4B8
1t4mn5xfe2As2BoKWR1DyEjf33K0HW+pnJ1SyT259kB+PRA+QBMQK2of/gU7JU2msr88/3wzH6g+
ecAmBsvHSs9bR0qe3TS2zkJnnMEN/IrnbyEByLMlpdFGIWm1WmLHrGrLXhPgxFGtyjPxSDn6LsYL
1EnAXmQtp+sBzJsxC8+TgliQXxTf9vIgqqs+E/rCcVQEqYIDGh7AaA8S7UVQqxdYy+6ptu3aB59a
UFQxK+meWz12ge7umZhc3jhUOhZImq0PVqQXIQxQLlLDkcfpb8CaLnm95JWEE/aVcjvwJRkG8PDt
Qvv4UzArI1Br/VccUdd3MiM4y8PhERfEvzQyNF4KbCQjiabXFg3SxrCx4yYPfnuI8umgw9L7tHQ4
hq32F1rnccDwCCMhnGxs/lwJ/BPJdgnoCyUxjOZfcrVLpNZCtXc0h8Pu8CpelFsVSxM78UcZ5evK
PzZti1ksbJmGMNajUGERCPUYRUvR8wkMr+eePWFVfE9By4DeZd61IJiU7a5R34eXwlkT+hvYMBE3
2lCdSZm2pA5CRakO0COVff0TIn3a8XAmjRrrIVytMebNNOO7ZymUqwesLCuXklyrOAJLe1XpqUv3
5fR2WcnGvbXSCmb4tPPYDc6s5xGvleUSc7pUoA7HXJtaGVWZyrPD99i6zUrZHYjgPtdExjHnQfcG
C+7uI18x1mKsM6NKRA4f6o5isNSciWTmERTKvul6W27ZJJwjW2xc3zmk653UDLZElvVSkKYYJsBa
cjAW1tQmhwSMlYZ+GFrIiDnfgEAwi4zmpjBmHC4HYXHRp6ydJkEX5rx+GOIcNXZLhH1yTPKSoQQZ
ETJBsuGgPu3und7MA2vvgSrZQxi7neUeKJnXWDGH2/+KNFhuTr9FKXiE8oDOj+arqZPCXzrszJzR
xaGyvDO2Tza2icV9gOOp1Y9fRt8coR9DxEISp0jl0Ja8J9KFvbeLwBrEb5SCGYWAJ1h5wyKPL9Lx
szZxMlJJWJpc46T7sX/bqY98c6Px5qvjEdJGYLLWzV1TvkR6YZjzNKyrVH9RVTpXTC0PCRw7C5vj
2OMwFeRqGM6+7y0CcB9FDoyeK2HxXwrCWFZ3bpqukUY8EElkrJ/QGUZfGo3nzTEhGNehcTWa4CsD
VT8tOdTzszINHxq/4z00JMJfqm5KxShDBg0wdkIZbBG0VLJ26CjeGUQNqVMvr3mVuoSjgaYgo2Qn
g8MwpiccJrZMEXdU2e6g0rZLbnCy9gQ5MADQ59rZYURPTUDCDm9EhkDoCKniQTgqEzclFODNMtSx
r9RasH8cVheOv7eOlp4SeOgJ4o+/iXKDIfqWrMF7PiTWzVLPl5/9n63YlpCqyIMWAs7Q6Jl38vg4
eqFg+wIocsYGPmlu24TrVABSAUOBICd0SWNCyOgf50WCJDREkh2xOY8DCmdI2ZuI2Nuy71Ab/6Oj
jwmOw4Vndn7tKR/UO3GuiFcsngWB8+NdoAfBIXeGemVc2+IuGF//aqArgYSkpmVqO9/wjd+UT4fn
n+92a7HgbzYE519ShYK/6o3nPzmYyNS19pNgjQA+YdevrMl09PtBD8ci408/d86+/9HslYJsyMzU
WX01Vp8pjG5XbcZf0jeVs43RSRfs74M5zoJ++UdUwfQ9DbQlhTdN3wsuUz850HQBSlt5MddbWhwP
LOWd+raCEf+tGbvSjrJfc1dAdq6ysv66LGZsYV8N19CluhSD8i083T6L47/CQTDJtjZztoGCh3Uq
x25Mak9L6sSq/Ctok0jiMnseVPipb4keWyFGtfTyC4UVz/FBU9Jb1Xjt2ODy8ypo4ryXo0jJu/xT
VGsDq+r9a7kqzPitJPUSCCtsyI6TTrHTXf6ErbJAvE5B0bo8cKUUtOpYYzY7R8fFqjjSg/Ojptli
5ebgwi5JeMqoUscGfINJIT60BQC8yvPZUV4ld/19ixDUK9NG7TJTE2Xn/oi/AUBKp3nocTCeX499
z4S6Xuit9xxKoBo4g2SD4rzuaitRTAdmXzeNWwC0fWmAwazHuQsSlT8K1HbHpMsBuBXQa4HamGhI
cnnuLZxiMBhol2hIc9hhzG7WSxQ810flUV6rQtZvKUzXkHhlxaQn9bFiH2GzASJXjCcY6vKuRXqF
JvJCmjn+ogj7YXyjqkdPP7b9qrVqL9SsH3KMALouLuwVqPtBCmTcl8UbTlIgdd7+rZH5C6FMhljE
LqhHqdkcrYdcPjcJ9kjGE3SdgKfZLaFMM/K+Jzx7t/VG3G1tOyNHTeybA0Cn4B6oRUA+n7SJvTeF
TxPUMU3PNLBmuG9/bbMF9WudBqmKTUktuI5eOJ3CHrLGqRAfAMQU279VCsl1BjDRruv9S3GjuUsf
Mt6te3WtDbKNLl6a7YmM3Qr8/P7xupgAaQ/J3xgFASDVfL+8zDIoWWS8xfcZizaZyoUE5MBC5fzO
QzNC2xAjYYeKsS4PEr24tWP8LL8NVWW9WBl4nDKtjA2LiqgUA2K6AEiV8lMe4V+IheU6MyVROzq2
dl6RdXmYps9g5v16fmc8XqGTS7WodbYFyYLgRqEQelzZfmbzWWJCbq1mLqLIq125WbB0mr+n0W0k
tYvgGRCIc2MjR9eUEnFGs15jy+Room4zNUVKIKz/dnTHSv6IA9w/2aT5U3Eafl+jKsQO/ygRgKJe
+m54z0Gg8m1NnuJcWULFf1UUfbaARf3vIRe0K/9J3CAcBpYshXY9unbQPgDIEslobmq8YOKF2n9x
rVUS+QZmzX3rfpR6CVczaSU64kYkcFG1COBv8UO74kFdIUJeOR4+LjVW7bYJ8k4QpXgC//y47BPH
1ZgdMZOWPQWnDIA9wNL5und0EoRLY42ysLDSkiJN2Y+8I3CXbaSAAD704ptmQAzwf2c1BYCDH0fn
VSV7331VHQY8ZXFp8kf2CilJKmhhEeYi/BHVde5BoUMMTvYgtfPiFGggWLGYdoNt68XW8G2wINlU
enk2KKNN+Kyr++a+fqlWh2Cqf5BwXtdYT1tvY1y+M0TsJJLMf3sM8gjQA32pzdCMj3vIvawNhJKM
oggF3WA4HWihW7LIEo0ZLx7+etjPTbNfh+5+Vkscv7QL6aRp2l7zGaVbKDGldKgpNSeCHC/ozuJe
GgGzHhVrWxZ0/kzlrM13QR5HLplYjMU9wFlndvHjQJAqgsYam9dg2I89VUZVP48zZqn2KGOBFB5k
3XlyYhVqpAIRo/DwBxU6hnV4sethwBkUgR9H5OnYKnZ3JbR6stg7tGlg3EcrEf4+mCg++E8nyPQp
fXDyiJfEx3IS0mfTJzyu9+WNgOs2Cnh2xEvJjnP0ySSIpNgpCdNL3rnzSYm8Gs286KU69c1RHOVV
d4QsB6ldBnTlMwI1lWfvJWx7cTRQ9zTGtr3mgXngYpC2yvQv+zDBcIe79jyUofl/eK6ucedflDQ4
Mh7ejuyoIfBoedlJSdBSYbs9oQQKJ41RfDmjPVyB3HUvD/F34BBFk24jJO2lNsiurN1omWKx/sHF
daM8jIRXDEduMQ3/GWlswrIOw3EpCZp8ZejCiGosZ4QaTlsKyks7bVzWs3SyGkkndzYX5rB1OW8w
qR1vjgNGWrBTUXsrf/n6nKhJr4nnC01njWG71AsxR+8Ym7La2bgg5pRnrs5B7Tc+Bp38+QcJhU3c
Lng3wxBz+/HQEYQk92n+beGFDgi2eSMPkdpVn000ezQD+/WOVe7x6ihGr2xgO3KUrHYPPWK2JcY3
RP8ZfJd1QaYPDqYq/3VQge3a5W8TY0Y8cd2S2uf0x7IagsMr6Lgknt19mVfvmdAwHx91IS4klWMy
pJ4nd1LJdSngkoEh7yNwP9kgMRQ1JgLX5bHIMAgZSg2aRw7OCMcpQ511aPLz0sgA5CZrqNbx7OwY
i2KgAq6ZsX6VfffIRncVFyHa2CnXyAhLKbpMXUPKLb+A5GAbd2Ho5LLXeh0IWqKPYrSyipMJG3VQ
mzdL5bbbYKwhftxGOnawAYLd8yRrK1wDPLfy3pM481MWvN5jQVOVE5eJH+V2+lmhV7qcHBstxd2F
/NAvU7hkN+NVUVV9yBLlW8CyYiDfzICkzMXNnEgOlyZUAEeX7BLbuHmv47lOtZniI4KZCvrN3e6n
cSmvplA2EbbfBkkILGkHJaZl8lAR4rdoQLtli5mOwLLDyIJ0Brw5/psDo/M0NnT6ZgKdaG/VVL7+
pYdI9P99P22DoU3hfgjB79DT1vcYNFPGFF3F2EIYGEbrNdKDOjjgtdne2JX4nn+HT8McBN+SHt1X
gGJTN/3EeScy3cJLAzF3ue+SBAY7NwUmsA7ooevIHPnaV9JVB4Nxgg2qnKx7kRn8+1wW41p1Qrhp
D3mEonYRRy0yGTDaPAdMwX3fB8LEC63Bzx1Lakn7gaJQeeOkkK3e8r/M/NVaUsYm7jaMJVbVxuQn
RhwX4kakUYhasTK4TAdymxG9Pz8kllsxBsJT9u4FCTSXTt0gE7fEQY0/pme9UxI9xaX35Owiv9t5
e78mEdf17ws6uv4f38cW+3sot+PWlaVGHW+8sLghq8xKiIGu5RAbDM/PJGvHwUZga+xMkzdjNwCe
WLoO/Dn6g7+VX3p/oxwlVokRCT6zuQD1kX8C9TKFdeqTg/0lBFVp8mtQWLfP3ROkB2oJVjeDBf8j
RUFgOLv9/65/RhHgOYwLDVoD/+FdiK91t605PthwGBLN3C+miFAKCORteHd842kmvgau3v6kqi64
IptAOw9yqCOH7oV6jt8YSbQhiKszEUCCymP6ASbv7ykXaH0k17KAtkOY2d41hyQi4meTVgP3z1j1
zwTWUjJXAyZQEWNQ0Zbz5SR19s9bW3f+qePD5U9Ro4npASL1nWhFeVJ5XFsTl5XVXzIGUq6FpnfM
MSMRoRj81FvaYtkvsW606NR2qIQ7x7UldcyCbtV2UajyosUGLcgWeCmoOX2L8Kxbqm7HtQOrxMKN
gSdeSBXdTN7DrMuKp/WefrwMciro9NJblunGC63p6MzWGHWL3dVFcT4STOWFLsnNmYovJoy0hltf
/TvMOchLA+MA4S2Si3n6MDErZEyvxoWT3Fv6CdrMMObou8CxZb6kJdDkD/YmNCGSOlbQ0nfLM2UP
FuegP5CGdBq5QMWwLmyB60y46kZANctLpC8TvG1Y2C+bNey0tGp9b92ZL4rQMGiUTlIR8mwdfnC6
yXyrIsBbXZfniNAb/ZXDeCwVkIuYN3yR9yCCSH3AjJ3STu88P/6X+5eIII1kwwA0BayFtYhhQ6E8
E1ehvL1t1/qFey8uELFlNoZPz40xEnc1ohbu1vzPD6gwcPUg7XhYwisMM9TstwhvNO9kAKb3YJX3
fyjjj9PiJaCrs4L+s0CBWEhOenNY966aYBsljXrELBRF1h/7AQiV1AVDtKXj2YUgP3T3iqav0BvR
0NFGXWrKuZ+hUnnzWXGQ/uy2UgTCLvg76F5XWzQn/npwl889x1zFxPlE70w/HXguIHReSEUHZilD
l1lbPz7ttLz16S5P7EIa8mBwujPs85LsLvjXCCqvdT3FlcutgPiIdhaJbhL+gXRzruwtEBYodz/0
6cVkREYBlF9/e/M6i0N3XVAwMvdlTjU+81+W9P7THsgmbVYIYoWnMskCKd+dxR0o2LRhBgWwfBdK
AauSblItDGG0+07pBIPLCLwLHsHH+HqpktGnnQqWtL0nE2qGbCpTXEhixO7YQScMCpP+J1kwnxwn
hyu9+JNYIw4illYtLTdeQn/1tOGAiT/dJlJZ+Di98vauyY66tXXnsZW7bCD0Qcu2Qorp6F3S1lwT
5NQhUvZ50LS6kQfnRgYX3BSLhZiKU/rR/bRrpr86wENo/k2whJhzOte2b3mIYh+TOeqpP9woYirk
TeRNr4p9tnJqNtMf6BqbgNflG3CTXrJSaNdwHe90kW1JwMPmHzWh7Q0mrL0/8GtSf009KCkVvCoB
1IvLVBQdqgf5AqAWkZ481u3lFtVuHOg1gNsX7qXanKmw/aEGkDHLu4Az8kRRvbUi+B3k5Fr6sP++
GTv1L3q1R20WHFMIIVQlIqGTdVPh1dBArLQy07xeLFdV+jy+XQzGjJjgrw1eQFh9W4CudUdpCGsZ
irAnbP7GrSOpMjCPfXnlOiQTTVSlHsO/9LNPMn933vPBkc4jm1zQixdMnCJL8hF9waNHWoq0nqri
OUQWJtOuURPIyIvKT60365m2K5/Yo9cCe6DQnF9ROcIvBzWuVWBwEx9Nc7DQki3zBgkXoQJPk0W7
8BhXx//wJVCZkq3Fmkkre/CTyMRkJFFFl8UaA+iYf8GrztyFoVVRz4qHfj6gaAIBiWz7v3qRPAK9
fqNKAXAJVcvsfgp45MqacbRmrg35p16ZrE9P+iDe9qchCJDBgkxEKE/NfZJTJB6Gz5Lgyezmgipz
MuRrtsqkhJd3Dn2YDd9pyKdSYhUNggTaqZsv2cqnHIbQzpQbOCmNPguF8ONDWK32M4QA9C87PUoL
i/YKEGWXjhRI/qAAakkHTiBr1NJLPEJ07iKQtz04dSVQU9i6vI+v807tgawaN6gt0IuCFlVK6jmc
bW6hkh0oPxnEN8egRJCOkO/7tOE6+UWLdojYGSqDuv5NJZH4JlNmcNLfpIkNYgk6CEuo3GPjPRI9
4nI+OsSXEZgpsp62ak9HB6xCeY4hW98BNKKBZIHAPb+HoYvPRF8TTo1SKsMbFcWVRk6+q7MpSnrk
sM/JDTZPaE4oqRx6suMcGhmFSEF+ysT0trarSthFf8leST58DelNr1jajDQ5tvztXXBsSaf0v0D0
EwVokdysd1e6CQsaUrcFmod10GFm5jG1tkW5AMMCjNPDlguRbeF/3Y4uT7uLosvLLN3/zFkdpZ1t
qbYikfuV7skQ/5S0t/VOZVk2i/3Hwb/iKqMmYcMD7dLOWZp2ZZcjdQ/gpJ9wTq2FclVcVh9CUWgU
4USjqMpgpWVj2qS8DlOeMv2HF/5Cc4O9Xrjb8r9wS4UXqpCWM/hi/01E3cj2ujeSX55KHmHWuZVT
7Frsx1tc6hvv6a+X9K0tL1XPw/kOUvW6Hi0/2JvheLr2Jt0y0nOclUoShCm3ouBe2KsdGMznWwrZ
uTc08ZzvTSlyCQRXrBiUfEt/bhpMZUquashZQPSC4ZHYb4f3ORe/UK7KZlJkNLKTq3R3P53nfhhK
tg8/mTzf+kCcEeqfoQVZumxsdBko372vR2SmpK2w/i41Wn+wBxQinWPY25TbTzTDCEPj/EM5q4WP
f+uQaH1wkdPdP+q8yLB1S7wtGVRlt/iTPAoRLsZlKyJ1EgJ9TRtnIXRSsXwp60mu0DaOjYByJnIL
dFhNhS7RSMF/o1f1fQcbl5dLoMSU6PK6B83y1ZVVnOhuSecU5gb6DeCdL6CJxjA6+RnxejT+Z1Lj
paV2W126+PELGQxP61+52l75KyI2ueLzRRBZO3fkY26CNKwpnBAAVYjDtaTFyTl/CBIYYhpJraVc
8ArlLidqKjj28zVJ3HUGiFMZ84OrlcT1hX5ZZbl+rDrqx/fD9ztMsqIX+pA0Rq7BtQud/+DPzyH9
zFDV92lEHzYC4ztBoTA2TwN6ZhnXjZpK5mxygF2bUQdy1U4WAL5e4lTXPIyhh73NXNkxMxTmXj9U
404oxeQfYb/SLgs7kvs02nAcBJlOpjwNzqu1a/nIZEHvTDaZq34avFYbzWigSmtjLtYhdDhkqFga
hxt9DEawOWiX9ZwMkBrDNI/ljy/dzrvCrUgr9QlmufOv7XWwZlqCHqJXVkFvT4/SVeA5SC9F7g3i
XrqNwbm+3FQg/w/yfhIYqdwxsoaMm9+r0+gCdd3eturYds1P/7F0CVl3w91KbMxqf/cy2x8390BX
IWvj0vjt6m7kNVy4kZuDfF6ESsHmhI0c2K6x5yIEcQk2g8BOlFuv7OecMdu0lV4xF9dSJn3zi7/z
Q3Nj4bPlVk8XkqucwBqVjPeMjfvLFZ3zFrLfs091sbn/OenwTpneDXLHRlzEfVgLOQ4nCWnjYGOn
wJvcUE2YhXZ7ih+u2K9FDh82iQRB9k7va9NelT6KPXDbeB3qovXBo3tzwsTvMqoObLeEdmDuqt0N
JS3GzDT6Kq4uJM4Uh04WFnzirFlXFs00JqwuGkOJOI2c4WD067pOSgPhBB59Syr3S2BTdRNqeXJM
OIM9dfYg+7jh3jhoS+GMC966JV4GN1YB1vskefofdSVQcxql1cdZ0jbWsuAtKa8XRuVig3QG4Ejf
GclOPJ7hjebubOVU6M91olT2waQ3zNNd9cUXGuO4sgyy3aJR/jzAs2wrsJyNSUYdH6FUH+0Qmw5+
Y9mWyhzs+ktEOqeNYElUkzK/OLfqD6cap1Pvz7rP8sLPhhIhT+lw41VOvt110aBzI/dEdKWvmSqe
gT2WFDEVxUTgKQ2OK9Xo/758/VFWpx60KeEa5KUkg2FbNwHJr9nFdNT/G11gFtvZ0UnFFsaJb55G
tpn6XNDzj9KqAeki1JYmPPxcZsi08NNcaGs0Sx4m3/0EBToXbsttarGdTrkQhM3xNVa+PoOhFDXN
BS8QwmA3U8nqrYoW9KSqbtUfx0Zxsyj438VzQEQ4V7LIIu0jhj856NmvTfFHVEeqIP8v3bn50rlq
TY4s7doeS//npTkn15Tzr/qZPoTI02ZQ/w7mQA27j9RnM9gKH3vNn4kwOHdi4xCeBNvBOHDeUKn9
EZ8hRxk+JLj9Rgy1I+iOxD61odm/iNf4uZ/pveSkpC3tSemtSkhAd7f9tXZLOB1joMsIY2tWdnLi
wEAfe04LXONmj5MWUGVccqvexNzOKpnjbBKpLTX1JH87wILKiI3gM9blmfwN/IBQHmT7nvKWJnpX
KdFJ4woLXFGCCx6yrU4aXpD7+7CfBvn/h4oyUtLPuXyyVz2JLRni2Ohf470fb8w+7B7rSDgmHc0K
m5FvnhI7UI6AzKspFCIsqEBSD/7NLEqH5Fxg+fQbuZU2lAwRRfCWl2ASRlE9XAtUgTgVywUbrffm
HKcLYdGRkqduSBWHYnbPsbRRCiZXHjLZ8/NqbmZvRr8TMrwh2DhDbNO18w0/QgdPksjssBIKTOLy
7utByO2HQdtmNoddmzLAlMQ2ywNcssjy3hQ2FK9hSaZs8P4TRwIWNK23WngFe/3vbxbuMamep4tb
Gay/YiLLyjNMxZlNBAoxkkKa+SzVnpaZ2qsjKsev+Ji6gJDzT9EBkhnKPccgSyNMbYBLMUzlGqL/
MZsTYGCmrIzxGm+QE6++FgHr22b4FGQWbzXbHBbz0ZnAIpNtaki8/G4c0LLKo375AhdBI1La/aDA
dDD43AywosY5vWt02N16xrEyUVvr4c6Z4csFY+Nqmsu/+8mKyizwznI+YEnywHwNiuHFUXxfIVvJ
I75sje9PAHK0RHQ0BqferawM0yD5KvadFS13bACMsTXruQNGNIneK2A4PLFcCIEOgnXIxwm+K5kE
EuXZM5vECd48pyhydL+BXNK3/7fNC81LWh/oatgg+TLs83q+ZINaYg1rbRqDQGPsCzlaUeP9PS/w
WdVOVDDCYP6eTEpjPfX+e1///57XgdbiLhcFcQV6Uhc6M/R2YirVPN32uVW9X13Ayac7Dm3fpjGH
vu5FQADmr1wJBb8D1vsQyJUhqmObiYI1r4sir1ONecvwTY2hHABYJhoDQ9Js3VOjKM3sOPLBmIvu
p7/8owqP+t0cyp6xPskdWldtqxAjE1uf/hy5smJk/IzFCcvw9NmignfPF4CRCEPgXIL1SlOEn8YF
E62TE5SLhz7HaeJoUJp0XRvTH1HC3AjBGwp+PeHLgWZ4TGTO5U1FbYD3sfdQAv8Ecg2ep/9ruVoD
t2T/FYwrO4s8n8bdpOhTAQ62EPXNtXN+PV18gzASO23Ck+tL39jwrA8JnPVVk4kJodvibdKiogBL
X3FSFHbkuc2R0gJ+HKSHIoZ02I0H0dByU1McNPi4cLi3i5kgwopG/kuuAVQI6We43dtchorhZYO7
14ZL5VMRY7k/+kGQMrxnR8Ewv8AlUz+9Uh5aPCIlQHXH8ByS5g/iV79p0xyKxyMVIAC9UdPAl0Nd
I1rxW/7MTd11Xw8B5EmeZoUt5r/YQgQYaM2UvXc2xGv4ZJdBVlAQ0prH1e5TPWs0wcbTsFPZtff/
qXiCPOaYEZMgg6kBWpw3hMtfjF2TbsMNu/SzeSAu3oa1xZg83J7pDoqN+NECkwdhR2zRXJMBH5cO
Y5jkuDabks844cmIE9ZknC+pYHQE4ybFEjVUKGtE8ZYayoAUgEu+hXg4/94D+oZwewCd2Zva0Zff
0K+OIJxvZepCqBuzehDobCziMWHoFCNK/t6fSlHVD+uxSGsquOGO8VZaW+cC/OAUSCfQPOHZ/+I8
NHeoSiXzmk5siMgnGLR+Ud+7zi/srAn4A301WCDHT+y8+LgEOJ+w+3sxnqy5sT70/jmPaXdI4gT3
Yny+Sba3dJst5+DQSTGm+n6kHKiuxxiHG+KxSK48XdjqeLxMsqKrljfFLVzCU3waBQ/hK1x4lx2D
8YTspaC80+dy6UWJqNITnkt8BqrNH4bH2bVphiycCKAcZGmd5K8meUI7N1KOBBDZBbrt3nz/BRm/
zVkRIMTWQn4/Tmhc36Jz42paPKail1eGN+ihBvicrqLybhHlbelhC7o/j9Igo6wuMAwrfw9lfEPw
LWlA62tmTYCpQSJE9j86Q0HMijFh2hIweKlUil0YqM6eyKxdiAdtVkxEZM5ecJp2e83Zuip0Oz2Z
A79kF+qDh35MuVWR56wI78SgKYXfDE0bPEC87IGguzmmp1Ant6VpL3SuWlKlaa1586nSdfDGjicU
rpioyLvMz5fKdRzsTDshjxa8WZkpJuwJXsWhoT1aXnaUEP1grmOKM3ZjtGKEWJoEAbMiWFNuOqrT
H+kEaeM/RoaL3G3w691XvsyQ0DJ1YM7oMQSLUTxAtByEbrvPabLq2adqDbwPgtL2o47vTZ5UKmS0
8WtiuHx5A9+m18oLwY95fXSqStbs0VVIQCwIu4Z6+1C0E+XslfhBgUowsC24ztwmOJHhzHx+Uya4
PLPRe4WYS/uSKLrDwT31IlrtyJA0Am9ketTNH0+1u7CWjr1g/LXyjTmKQHAVnndyMxQ9vxjjfdjJ
WVwbk3/EYpsmhVaxeZ/UEGE59/G/Aa1YOjLFePVdAnfRxXQYUCDfFmebVwEnMJh3LvrZXn4uTheL
izcpM02Rj0QiD6locNYU1pHUiZHNchKHjiaUVTQTFZqLN5q6pSXxBLliAMyicRZp1BV6hZSJghON
TAqTzDtlXJQOh9ZxtJjkobHskd7OkvEim+DJyNqCzdHkEJor2b6ejKPFqNlkFoClg+vTXT4SgOlo
TzCbxv+NAim2qFrTKra9+nxbbEQSG8xK4xNLniTf2gtnoVkkWeXQS2eu2sQADtm6fmjK32oblnF7
PPj4VFi7rVC8LLgrhK+70uLYnnoyYoezzczdH1e1UqqFvb+9Z+6+vimTLgJyrNTryCgoVbeYTduz
dXHqxnVHUyIIy7cDX+i6bnQM3y0HGd4Za6AXqBeLWNMhxtP5ZtQN7sdEqFR0qu5Tz9GDCtAy0RLl
pJrUUeVNdpq86BHo7gIaeI9YxTc5ROojVGkZdTAbkFbiwU2nshvK47BDb/3corICCYSswcMe64w1
xDfA+8iR+TOH6kTMq/CUh/tLiS7sfCp0jkqzo42UkejDja36/TF+ojJ3X3xLWmjClQpHjOer+J6j
geZ+lRJUhV159PY0olPn97r9ldTSJ1SfVPtMjHSiUNUyI7D2x0WjEi6xTc96JZ4unqbVkPnj/pm4
Uoi9XUkiikAgeB1xZ01VIrdvZ3EgU1PgtQyVLSslTdgcEp65+NRN5Ropx/iOQGMLtZL/rcGzYqE3
XRenTC/YRm9p6UohK5ucsdfZelKZu/yS2KdPxTuZ/02r4/ypAFmFsUhxVn0jePt5ImObctBGRVJR
5BaWKP14cbWvE+D+OEHiBPu4PoUlyoT1966Bd68Pjc2VuIMBYB5nidBTKe2pCxPXZ3+lFJrTe8/v
ZA/HqHkQKHCj6nEBl++JfwiELHPbJnvJKFRQ4nrOF6xjQIDI8eopnPMmAHqQ3K2F8mc2LFK/Iljq
sGzMbNWF2lPS6wwpaejA4JpWghMf7Sn+jFBMtl+qJ2Nl1R6YocyZGeiuNFmK8VaCwmIWWiNMuY+u
/ewH17+gB6b6zIaICdOdaDmTu6yEh1CTjil58+jsd4g6iNeLnAC9va27QAJAGizvgBNeHWIxBhcG
h1EcbXHPxfG4BJJKOgLG/R5JRFvX1kxZUWxgaT4gTaVJt3WA9NuwV6sGcC8qndAhbyp0oYv48CLa
W/EHSu7w+iAmOY8d7YUTnyjDx+TsscS9afnwhRTkJlwPVEoKR7c3QMHAvPeDN81Os5W5jiIBEMrI
0pPv3yls9OCU3x8CXDW33OnTyj3H9lClDjOVqKO8F3XMMqvofqNJbKIbAZfIeRllda8Yg5Z8h2z+
xJu3D2+o3y7YPmcI1dZMNXu1xWqIjH7AgUCTg2wfWs8+fLBTCkZyr1N8HhELMUwxSQvvcd+GjKtj
ZHbpBz7GLPd7id7X10yEYkzT1KZ+Uf191Ve+Zbl7LTM+D0DnPTfzB3PSMWI8ni37R/CnWQV62891
ZNFt+wM/1O2sgT5JEfxu6R2rcpyBYV9pn3P2ALN1G91wbunNXlDM1Ja/yISgj2a79dse3SnUGZIK
pWqpJRe1EKpPyb+37zJxCyfscyyUQq5DpaHaUqHwXtAXrBd7jkJ5jdSnyXCCjdxwNPpQKv9wQ/8a
bLoFeqhiPYxPXmx7SQVZ0aEV2W8KgPMV8Vg6VSCWILHIj4yae/L2hZD4GP5Di+qcXwTj+JvL3mWR
PugQFBbK+TQ929FsblukfYYob5Z7ddTqeAGAJ6166gGSt60uB/jZTkOKzu6ZfFurV2YEkJq+lFlO
k68A90lA1BZbB0WptYmSqO58dQ+ywyJVJmrQldYC/QEkiIVuv/OX366NJsRh49RAy7RHMaL2exX7
qmli/LyM0hoX4eEyFpBsqMvT6vDocw/Qm2CAbqKMMZvhNTmOIzy2B/drQpF6JMuT6fl9D7Q9UkYY
YH/JzhFeKClv41RxypohLXhoTfSJVXkmcYtCH/Efu66YunBfFAVej+C/knynBS1CwYWG3OScjhxK
+DF6rH8LRHbvSAAlBmldxW+a6vJOwIyJQBt/yoYPe8MqVNQ77lvOENt2tl2rjLwzws2WLAQme0GZ
U0Dc+mrmRSBb5rQGf9OLJEeiT9y6pHSa7iasFOojluNGSfFSsT0Ob/X+1y0S5A7h7wfJ858cVBb5
7u7tpjYRDE1UtwRLtWe5pQ+MAlpFho/fo5oKGO/OIqtOjjOlb886GZW7aQ7fIftghf6YTbx2fDoR
gbV+jTirtQ0nR3iDKpnAkr8t7Np15rDi5jNnZaeBqsChHMkoeuaplLnZXYnmvvXMKfDy9Gr7cJbq
rX8SHsEmOfYWYmaeB+Y/URVdpV2ZGQlw8frzVbjwzr//AjKRA3G1KkbIiL+EjXy4PDKC/Xrs1zQJ
NrVks4dCvcL/XlC/skm9O2MjPILGSdTkqKYjlURXHsAEgVDfMn3kGhN5TEQZSyA6cUQWdTnOAgPk
KLDL5Yuph1SIfQ1YVB2oVP41BmmPt6OKVTU4ShMQ97dqx7WeHJww9PljaRaJti0cWEmfIqVoLmdO
o/hHbUzPDXckknbThwDILMImPSLnsbR151osU+pEc5ogNtkHSkGZaHhSWEpGBLVHILBAEE7UNR97
3eAgQE8glg3gAkPghYHbqArUffcAGlPvimvExpcWDnt9TvGpAHdRBn5GD5neKaU/Hs/nK6g5UXqk
PKo0/pHdw9n33lmAL/MZs2BT/LpMp8rlKgE4jZuqv/d62HWYyrurU7fsV/+o+wutOi2prpMIeerh
iGFF54wYNlY6GFHUF5y75X/lACwWBvegUW0PJJHFPOt7/yad2wIoQIOU9thK2hn5DGTjangZn2RH
DFIlZFJlnJzI235MiBTXj4xMNOjhFnx2FI9477zeUc6Q2vryF4dqTlUpckLJHZiC7u/0yttAerPp
S5qJPGBx+vHWIBkaV5ulubCCeU46Awpg9vYVxqQ2OXla0CAWvnz2Y/ndCFMerhiJNfGcmI8YNj0h
7GCtWp6d1mHw4eu1Yld+yVpBEKYUWXAvaoAkpLS8JqwN/gRO/nLCKl4ygeLyTMk0pWpcwehZuqgG
45SGHZ8mAMwdBpUKKbH13ZoV+tXPt/jiZJUwtlaQgpvCsW7ia4Hii1SEloGLT+gNw24VWrOszH2T
RVUw5MO/BHL2U1/g9HJ3MnsfgWjFpb1AJ1Nc+OcFNYVewRryTmJuhSOhT0CNV54nth/BpuXZhwZY
FubJdg1+5J9GSuiWPxR471RwayIBPjqPRaRMBLbscUjGf8V2jXiR5ywPpGIsL2HUo9rtC8z4rlm/
strhwWzfABpOvdneCILhYN/1+IU14Thg8MFChce51iXqwVuJTjEeXjmAUUJQN8NmTOSda75N15Hf
ZDrKFsNPMwFZAA8qAEz9bFkZaJ/ZeT5Y4Isj2Q4WMf6LhhaBDAbQ4gwtBKZ/aMSVm58nPfrMh2s4
n+5Xw1BxCBVA/im9iNna9mQEbfpkkbYPCSwURtYPvcBIlVCRknRBiMUSLCxNem0vNnrz2MibfAMN
uneZw1tgrNifeLVTSyyi0zGPBwxwb6Ve7iLUJtbEBRcVGMQyXn+6j5uAwRRe724tmHt97mN9psuc
DbVBaTuZRR8ThJKU59UhMWiu9/rLbsMHE6YX2xVRbSyi0Qo/PLo5R4gF8j4GGOzibyFAueAtGYGM
k5QMx0vcH1HX0O7LiJwxBoTsGzILf3Uyyep3Zzt4cXQKGPpkUhHno+r7b9R+GEvep+CxOb/x7W4v
NQk7ep7PmBFUcwFP24HvXfvSB913pzhRHTvFlV0gAYEqpHmT8dcqtmJE2M+ZMowIMaHV0s0Kdw1m
9b2zY4GyeuYv1Zr8V/E2hJQUI4+iLK19/2ZESNzYznkRw3lhjC9BMFqWVPp5x99ZGZ4zet1BiInB
JG+yo4/+J0+VofFU3Qgo4AUm+vW6a0/XIkNCfc//1N7cD+KvV8rRb+Sg3JhTe5d3Kact28BUuZ3u
59p6j7ylHsKfJjfFynAxSn0lDLwr5IhnK/f3sj44r7LW/aVnsx9aVZwWdcAZKw5ps2hhdRBqp23e
6zwAK6SVafHLV7kpqmBn6m2g67jTd3Q85UNimij8gnZJSSN3ah3rsecN+XnK/FI0E+U57va6jSUg
TgS8IN+6S3QwUS+T590xMbEe0cJ1yBiB1z5o8q6A7QEhmWVWMsstpCIcG/tQ3GqzIoYNax/tIeM0
LhaWIiJdRhqoc/FJ/a2sR+1drr7rEeuZ94eEz1bEZdyaMGHkVgAZ+R5LW/P2vHdnqq7Gk57K+43J
L16+Kjloida9jZivAzWD7XmhF236F/4pE0h9wanF7nj+nTgoZwhqLj4vA+0/B//r3rWV6Oc8U5MV
5khCUsyH1ALre7xgbIU171VP18KqMz+gcnQOYwVt7ZqTCcB4fKMiaTPj4voW1lf6hyvlj6EsHlbX
P6UI3/s0bFAOmZe9tcSt6N5YoKTbf4uVAtDfH4A1Z7sPSw+/6aJ90lB8gToEWs4m/dz0lM8ciztJ
8v2/2lsdSXP3hmipCjI8LBlu5mVSIKj2ND8tQutoXmjWCaISeRh1w4DsPdCghEd5usI++AkhiSzF
BgVkuklT2EcaEMOFkyF+p5PEAuWxmdit5q5BbQSTw7JHuYuiDSyfn3LDCBawldoa0rQ/RruJKkyP
t7cjB+6hkq41q0J2we8fO4+R+WQ3gbW2/sT4YwFgJv0gniTv7kDOojtKY9G+/oRlPmZxWkO1uFgA
s25AH9oW+o4UwZsIArozBsYF/OCGg2dIGIKw0yAxfYMC7Ma9nzNgNAU8A3/CTMfJlDVGgsCYk6ty
3TOF0vm5LOpvk7hDtWbCmm4wIDLymzPj601a3Nfb3WHFMuPQhJvGnnVSKdzYihwUPkoCxYiQMlrE
bE5N1ctaju4L4dtNl60MdOnZ/VqQeQU3t+cJ6rWdP6UiAlfBR4FiCRL2dlTG5WhCtGS810n9VGE9
+I6M4mlLgD9rJlhh1pbpyymDELjghM+SCjzlPRsrWhJAfkXezlwhRvdNYVYDyClRJwEr+O7YnzRF
3ipJ/lvn/hfT1W/7W+vwsMy90uAaV8a3BUS9RDSZl8Tz9Ygb6ocngoZiA7w77jjj7QAyHYe5+2Qj
fh2NBnq4ywE6qJUgFrnBSOnaT86t0klaJHXf85PRITFrig6Wa9uIRruUWdrvaxOWCMs0MhGWiKwU
RAzqfgMhSdXg5n48RItRw+YelGXDRmHn9rlcueyfy+QIApk10Hcc0brfMSiuc0T5fllTQGwq6A43
LkyvHxxzu0mFC0mvXygfJmfYitSzScWP7NhicAhHer9VqtRk7xOkfwOuOEKzxbJiZhKioYUhMjN3
HZWNk9V63ovhW5iZeFv5YFlosgEoqx/rkCARtjAp8GMTfgWryVOnxqgcowoAitMMajobLgsxJ97B
SIh5LgItUTyDIIUDmBQl1cCUBaOdTiuLr1zxnAiMcA+XdLsbF+8zQ338ty7ONXePi41zPVp1G+Ip
3WwdKs3Qf58jVkCKwNW1jXz8mH0X/aHeZrXSI3ymVmyDsdlcrwpALM1DKL0AMuT49jvxMYpUOsjn
kpxBLXVoo7XUKRONqYS0y0l8N7K6KcDd5TiejWKeREdPRSCeb7mO4XeqLSH9Ywy8ZzVPzia7Tb3a
JYODrhoWTIwBeXOqfWU5X/gBTanAtJ3nG7tMra1D+1xJ981PZlmtvwvgGDizRpfF0OPUASrJJpzr
LBQ/tXVYcVadBXNQhNc2uK1fOPE9IEiHzSsjxVxqkR60Q7/XyO5cPUOkJf2G+szw1LX/JoHbAuge
Jl7EoUDwLRAExb3lBVk1TjIy+H5mbKm8OmWouO8w4C2pazjScnEoldvjXyTsD8spG3Y9HeIgp2le
dCkidaWhe+LI2ICVbZE+UqMEQcHCYly2xPK6QFfuLqWJif5JLPGgVdsXgVVWIWLy0w0soMMvpQzN
ZJ5ZQ0r5WBWdOLxPMFEpYNcfHGULN0ybyo4RwXQk+YM1CWsxBuFEuTLZNJ0npwbKNuoNH3hhiEUr
j3mVAQZOiZv8kZ+8gj+71xXo4069jnKUbSqusD8DhKMmcOdq97GTobtRFt4os1qAJoVAs0gUdtMX
uGRP6ytxEb53eg9rks9ICGRtOvuAV3p6c6qznunmPk+eft2Ay7dzrblCZ22HeMEniS2EQ45d3TnQ
yNG5Tsl4LHYZzgIlcMy9RyyM6SYQL8KPs1LNVFyESbnVkowEI5MGxOk8UEPHpsFnmfRGsykjqnfE
i/6fvx4KSh9n63ESOWydzXHc7K9C+Ky5PsGI7zn5njXpJC7G+hcGW81HYmE+2Npkmc4qr8691azC
x3c7ZU2aa51miRiL9MzDzvxljgXFy2O69hO68Mh6KSKhjVFmo+WqV2R4Dwklt+9/Boq8dbopCw/b
Bpf+TkbviZkVY1GIGnFu83E2ISSdp0b8Qg1nclATUy+O+CvTZckPqNZeNuZ06+CQgJg2LXCrR857
+iSAg0dNMrCWAyF228Lisi1ifpkPqbqqq+VaP0jALhHq9OprQqPlisMSyi51j1SO4V+wlzx9rG0T
hwgw91x6mOVdNur3a77kR83r2jTOWTUo/5P57ZlRRInRSuo3o99zPqDAYDEocZ6O90zN3BOYh7+6
H0uPMjtS+PdOGT9QMo47+aqy/xTXbCK1BHPoteY2EzF/CZPkiQ/vlqC4L+b/NIbPiQYmESwC4R8m
EFKvJHKCRQyyu+BAtUa3xaMN9ihFc3ZjsIu10e94Tj7qs1GtcpDF2gHbmTtr+Ybk3V9cEchIaODW
uaDhg7EilmAlhpnWr8Kwq2J2M5AjBZ8oH+Nsv1oP6XQWFsnR64+sPwAGwOAhpmEA+GyYuXprug7P
09kwJ2s4JGkpQBrMTxxPTwT9cyoi0enTGN/sCKJ8hZueNMg8d/sf4eTwuupH9NssSBbajc2AxCBU
TD2INb818uZpMCuzTBXnW7sgIWjaEmDfg+eEocJbFJyp2AaFoobwacL8UmX27nNbJsqoEeKZfJmm
ilRl9LITR28uWDbIv9j7TSpbuYt+/lsjsSBHckXzOglJimQoD3Xv7BLiu7wyZRt7UUUMsOowT7H5
a6p3oODhrKBa8Ymtm6A5HOUTG9tLWHqdEObNVB06PZqwyxuoy9RZTyfJkyqkBHuvRpWJmtyE9hOk
sAv0ZzhOBotsOZhtid0LEKTToHxm/r+DiQnK+GVn5qqwgwEwLYXwewBgu/1eGfYbV9xhn6qRKx9m
bNtgbPJfGn6iyJTP+lpHhV9Jp+6TgF2vSf/+uiYoOhAqGRW6Xd925EV1fj1RHueiQNCHOldjt7nW
sHtXCc5nB6W0f68LKQXgjVvc15p8h6f4+leKMTONPCzK4pK0gsAj9ATShGITaYLH67uQdsEIIoTA
xyk7jqyz1sUsYBDsDKjaHhVmhUM49d510Pu43rhLSn5qJ1fAjdk8QEAm02yFVmSiw+AHMQ0eez8n
Xs+B7dn47w7GtmRqmDYZHRJDrpMLK4n1OruUr/yk3Uqv+MJge82xEaiKUWEEcWItELTXgQNTKVnj
ujLYsDPh8ZkRsJdcpMFfa4xSP6KNq1alYG9OYzfa+kGChfjCOaSw9NLEydCMwoKPtpmOa8lFRpzY
ly4ukzVsrYMdPijvsVMz5uAYSPsNFFjZwQLYiCx+f8+xbILLPWxTT2o13Awj+cQYHT81AFuRo3G0
GB9XKL3Tk+wHIhIb87GoccTjHQEs9iYczqpxXoSS9ELPjqFQfsF2KdvK9nlk7xlQdNxVTPjfEQxq
GFkPMqV9djdWHfP3C5ouszPi8Cr7jFUTowf4hdFQEW2VsWdQqTftdE9NpoL3kkB5LuR2Ks4yqo5N
y6tSLtMOanl8PESio9TpbJWQZAwNki9AqZfbqjb92KuwQeqgY3vDPbpi6OtSJr2MA+Wyvwakq9iy
9t5sGzTBk5VTQWIx/IGHR1ySRWX9w676RVWy0+eCg2+rhQ2B1zlOONU7rq80HGA+veX8K5JKAvq1
30aw/q83FHdKZpXhg/KwgAN79dMyhvLmxYU4Yz50QAQUO7jaaTv+DxpayPQ97GKBZq0uTIkTkIyO
gyCzvQy62SBnTCvqoz+NmolLigXGOLHun88BSUWbwC4/Dvas7xdT1RsGHKlX3UN3FnsU87xwoqlQ
X43iYOvVwAKzAzyxwYCG20uMcMQaf3qhiqzc2BwLAaPAul5ejslTMf7V8wsTXPd7KFuSglenFk9a
XWGPGGtdRUOIcMmnkJ2T0ZXPZ8Mj/1HU6CC/9Xwbv8jpB20hMUheye7UJ0gIA6QhlzoWumAS0p9u
Q1qrCqBe7gaSr8DY5vd9r6STBTSog08dZ0kTrFKbWH51n1MV8PTUqrDl+O9iTysznSvpZhh2Xkc9
htH4LJR87uClG260l15citlV+u9oQl31ibLEg+w8SP2QUzJQh8U4OyEQCkJEbV7ci6YQ4mcgI0Oe
3t+uauKi8JYHKNrFSOiKJbhZeYhvnb4aY7pF+ekHbmgHP+7+ZuHI/8PYLtC1lR6i8yvtZx5OTZr5
joCRmKaR2wREAAhWW5UxC45Qt0kB/hlv/iwp+4mTHO8wu16aW6NXxNr3RLW1TSsDFGZrIE9BOuTt
lsBsWZomJ+7ViPrEpo6uBLAHAxucMMzSckZ/AtWuzTdtNz/Kp2HTO3Yw2jApOoRCYZ6fVM4Rvl2k
SXvlTTohgm295HjFZXwhUV0oDdq2KEIhR8O/0TXzOvR9M/Jn/PDo75jlz4ssP7v2fLQhHQ2rW49w
8+az8zn9YWC+hFBxuyDsigNXy8DUx9R1J1RiPdqxUHEc99QsbZcPDBWuumhymQRXuhqAb9dV36+V
SrKi9iucWgMEYj8YvbH7WTzoqaFaKsSGPQMtfuSYoLzmgFAtL46eiY7stidT+Z0dsrYHsYlJAPHb
HiZJChmf9x7mN8BoH0aBbzGKosaljYRLL78VsuxOnYM7WjkmgQVcKwmx80DEC3RQK/IvX0PjGrRH
RFCoGeeA3lFipU4WnCGAYVmIDK48mTM0aO1EXelgEna9tW8DWkBmN2ChvMVGpYtIY22b3+m4YoaL
91TRq2AshK47D8YpN7LoaaAL2guBrTqvcZsFGNpWitzfyqyNoUjTYiF+DVrInQNqgQx/TPZQeTCf
KZOlxrixJ/JJaV2C8lXzpaqqzD9MF23MP6gQh211FVNk7lOqUnngkSXSg5liwFZ67aBIb6PkZjSO
EuDkpY4JVYfBpM3l3Bt9RN24ipKbzDO4RXnVuG3v9MwA3IWk5geluXeC2cwKxNcB2B2wmA1icM7p
M1HcvtDCnEFyjUMBjqmsVE9/Mlfkyr5ZnjH3nks9wbzZR6RaJ6uPNl1bn1doDrLFSbZnP//5AlEq
LHpCZYHMYegTKxyrd7TzVxATcN4Ezzq7K318YJS/O5rdUcX8XTAnf8L6I2c7raWFaFjRz2qk1Mto
EosFXqTVLJwZxxx6aE9sudQZl6qja0jRZVJYASAJ4H5I1aBHOiuBgBC3Goyt9plrg/9ApWNARVVv
MuTsqwACuGPI4jfqT5VgJM8h+6ZnEUtU6zxLhPEXBR6aF1hScIVJRORPYYUoZ6GdFcu2RjsY80Qi
x7+jPi8PakfXIWcihVNwWTDR/L1/8XhZbjgvjkhEA/4m7iOHw9+HT/pRVLRZenPGwr566cdHwvCj
5ZzXHeRI6BfR+GC6fKc7lN1U44uAmarWscvzMOvsjfY2buHWkOvNRz9GPrU8ENQeIxCOJzW4zK2V
V9AEG2e7hJRbpSFt4lhwO64JNRTtLLYJjHfbyCpN7Nk5IHQsRWf+4mjAgikKL4B3tz0Wb3YVYoq3
R0cqH8rDZF1ZuiRXqPn2Kbgr/wnguzJ0QGubR8gJkpm7EjKhpVLPsiUSZXlG2y4LgA56bxXTDPFW
vHwcZn6p3cSTAZ869CEnFQmXl131P4t8NReNm4/2BGpyX6HPAawlW3z9Ou1YqMEbXxHdngH814Il
AUT/L3YqleT1hULT9WP1QFf+ekAOrKR4VIDODEm3NbuKXgpNTk270AGmObHq1CXftZozEDJE15Xb
5ASpcN2g2uyC9f7M1/+3VBNVoBLZT8j14QXz7iDuOb0+D+/UInqd6PNhHti5t1iMuCvKIs5iNlPw
BAZyeXXyDpXPWo06iiGipWkhM6HTLfCynDri367vSMOHaFKVdZqXBcIX5DF+g8vVZpkIrJ+g6tPl
gvu8gstBz7vMuwEWT8ZP5KRfwgyBTmaQGh2Sq74xFlno6L/5LJR3KY98L6Psy+lZ7ouacV1AQrt0
M4blbew9gYeJCbySVn74dzTc7NaR8bPRMGCQHWl05k3EMMnXAODF6avYoBbo95riTKlX7vUNoiqn
brerAJhI/IAVJEBD1fXznI5WhzY6SfNlELDg8Biio9XV8foRGrNQxxwfj3X70vnxDwIRbkql8m1U
E/6gEg8+sFQ3jC9EzTkd+17cppxpTu5pzP3C4PWfqcrx0NClJYxEcE56Zc+uuwhH3+33zcotjIPJ
liZudTctzVzXuneGC76UycimGp/E5kAAfr1/prwgm75cCPbuEkq2HtCQIuBn62f8pcrKjbqRBVbM
yNcQQdYqRldQtNSDAOR2SDQRyhhILdymQ6doJVp4PKLimTk4BvBoUZjNjpImCA/agq1o3Dm2gNTJ
cTPfvfVT2xoXXL626jc9QzajM9SzrnL9bvLtQMrDobU50HvDCHyKMWsJRoDLxG7nkkRfHFvMFiC4
tcSEhLquhjG/9WgS4Y8TafT/uWXqwDyPhA4MPvh2P03Ds0tGFUwNLLlpZXuchGI4j7pDmcF+5DB5
4OvNFb1w1rcU714xpT+0g/IVM7eJwDieVKg5oqWJrr8BB5jn5JakAGI/NTBSmfYZ8EXtRPGZ7e/B
/nWi3Vsde5IXQqpFpzyquiwunmjE9119JPjj3a2D29Sa9QiLgB2PXEStMNs4SL5KcpSUtoCNsk7X
xqnfVMP3Puy+gYmfh3yImX+1Ox6fmPXzbBNJ6dgbDGBDkCeiESLwz09vOxNwjKJPT7AfShi5L0NG
n03MT9FwKLMF6mdJGkyqrRx3Rkw3xgqpS7ogvnZz6zCa0ZAGlWDrD4Mfc8K0Ix+v86hNgM24L0RG
/78D4G2wYu9FDQT505mfWukeN8W4R8q05qVnKfktaHhiU3lwjej8b5NX8kE6r99nvGAR6A2aoXFh
0AclTs8wSX9qODncj6GDYqHxjAuHWsmdXEOCbDGbzFRELl6qDy14uZKoq2zCEdHxQzSnCx5Wjru/
M0/69juh11tRk3cboXe5F1NXS0tNVSDDHhooU0OlgYEfKhGsEFKZh1vgxoM3PLvcY7Qnmiqhhi2h
36vPjUlmnu21h1H4ixAkpypbYJye+s7EA3xq2E8HFQEXJGOuxkhHd2UvJ19ndasswaMMO0W8M+xG
wTZK89RLHLiSJ6o60wohtdouvrk3LaFEyYwex3obEcPazAi/VG7QjcnMaO1Gy+BR7n4xh53bjMjd
tBgjQH1DLbARNpYits/7zykHzx0Qr8oZo0OfbETNKTSZnhEj487ENoOliSH6gO1oDnBnanV8Pik/
gd/4gUDjN2JH9yiQb7WZBZC1yjEXQA4MXtuh1eL0oHIGbePnRLmwEna9YAD+Skm47xCPkKONGJL4
JlyLKAG3edUkDXdoD4fe045BBppT4exedSkiSMJ7HwilNDi4MPMuliiwfz1Up8Kl/cNQOJJzJqxn
gtrJgtvPNHqONWxh9ynnUcuymZbygMOyW/FkRH892n/2y5+Kdbi/7+vM5OuQLaP0VvmRC6SoD8vx
uqW6/Zrv/R5bzRQVOalcHKj+t1Xmy4rBHx13Emev7V6cCal3/5v7w1M5y7yVRBjtiVazPW8tr7cB
cJgoiVT6lUYyWTMDmPkbxfnhkTczKPRM449+frKV9UOttovM+B34GG6/muum4OMN1KJb9wye4Vo2
JWHYUlhk5DviZbqqf9ocCws306cQU2Rlufdg+VzR1N9pm75hLwsn/5eVPaG7TITtMRqgKr5azE93
kLDaX78OpHv46F1M2xEIB4GDw4qG7JskV990KIUjydbd+PwXr18gAQsEuBoWUO7+XKgO1+TtHhyi
UKyJ/9VZMSBG76VPA8WfUQhR/+2A2hAZTI1MyEtPJMr3G9jwnkbSW+giPHhvsRtopUosY8hep5lk
wsFORYv0e+uD+55LtyF38ENBaur0cX8jkq/ZB88x3iomKKUPudhOBk6T3dYgx70jlYOZOeziTWk0
0YImUTMUjPnc22TBOegcTMndMCgKKt09xY6Tr1Y9POF35TsuaPotP8GLs8XpX4qg6yOsk/dcBZuV
1leOG/wU/dZ1C1hn4ZJBTN+3OBwWNwKBVo6kjeZ9pAfMvCEh+2mEf5HJczz0RkoIELfvI0yt3q18
k7fuGPPlv3WdbaW7wsKzU7a8P4V8BlAPVkdiJkijebgDU5xVEkFoYGXCvdrsv7qfVj1Pq5D8B4f0
O9ZSzuae1Vd9c7afeTgrdBZaB603aRpR9XID0eDjXQKojqIT1bLyQTguTNr7YZ0XQKMAp4EyC/93
N+x3WkAdHFsKsUHpkOYqxY9kgodE/So2FjRoGx9YfIP/72VoM8OY2TugZeX8cDr3HSFVOhxfucQM
8piWy/DAy7r9++vTuw119jXdKmIqF5UwgkkPJyfMsvsRqgM5xyZFzOJUTuVQvBnug8N6+5+cGtaE
IOCemW3ZgsuU11T6w/uHRREIOjN7ZW5VjYJqirL4+OnwlERPDBF4CIMkNwJ8iskYTGP4BWqv4u/H
8aNc3Mn/WjYTBgSINW7C81BjPUCBEhD4PJ9gBWdeptaH3p6j20v+fbSSjJMkit06f30TFot7QA76
sJyOYu+ZkHeqn28WUKN+ctWvsi/0IlIX6nijPLIXLLl7daPI4b8jr2AT+xsiq8Qsspv/f8bd7y1S
OTiEftj+hEtQbBVbI4wj5EzF2PDniO0NkjouiT6bQQAM0sYSyZzFBUxGVkN53+qDUm7B4foVxPJ6
d410Qh3K6rQtIkydmc69Yt7YpJn6l9di5X0pzTfVei27QJ5xz3eojEkj09x00e1vhNf/a2wKwhsC
YziLv58DfgWEzGoUNm4NCuKhtmMFmKarCUp1of4Y3DYh9II1k2M8J63wU1h5NwvryH6yxqcJDocm
Vl9iwW1Yj8L8FbNlt0tAFdF4vV55Ql+vqhgMf4KEWiRQfKsCJLa8kFe25G4toHs8OoKyqV3jJrn4
Ihgq4kYLIXxtlavpLrbeC/ESsY3D47JV6zKR/hlp8zvHz47W3AWPwyVhnHsKHOa2ztgCpiERu/bb
7/Qg9U9cWGms1Ep9sbymFY8GrW1Mf8jU8hRG+D/DN/b+GncCz7lbZgN/KPMyjPjg0i5699q+4kxi
Jg16LZxFmZM9Hq4zl0toR+q5y+dLwSTw0eoFUokqV7w54bg0LXgIwZIKKYH3GufrluveY46qy/bX
LdAQdmKY7Fg5gNPx0e+WJkU4XagKolf54VsObooiYNecgcUzNBBsKwsF5U/DhWRD3tW/wOumFFB5
yP3YEs9skiZrj32bon9BzG7M+9EfEdXl2kTfrPTuJ0oDT6a18Y7Mu96Qjk5YUfEEHudH4oNRh/BQ
F/IPWQFJqFyMwzAoeZmrTg8qZo8/pGj6UtkJEBIJB3t82st15wz2X74InZ0TC7e9Y4wmzPkcui5s
ho7x6LGy5xJHYBa5muDj9RANdzEKjCLVooSBV7NtHzoqqP/xqRmYAAbrJSLHbpysbHS0aTROm4W1
AfeaHjts2P2F/VCsonnXZStFi9j/4fvVaTp1b9myrW4KylMoq2pU27GPIWaj2m4P1oFz2pWRwIAF
OUSDFOjssoyHYHbJUlRwv1u4DTR158sPR2ASjvfMFVZE76s+M9r7or8sLjqLBV4DRcvNdFuBKlvU
daLZOEYjx55bD/97SKY4lyYXas5AnF4zqzxsCvzSDkf0ZNXk6TMC3KG4ggKDMiAAxgxx2DDkb1IE
VnhbX5QYSlpuu1g2sMISSJK7RCVP4waShtnDs6zP5LRtWwSd2wmB8s95dpU7CTtDNSgOff+zN/Nj
LAsoKdERV3VhO3ePozW6M8V3Y23R3QMflDJzpMCbLYVlW65qLDWVZPUgIuhMdI0V6Zb4hJku4T2i
K3T/RH2K9nQYIKZibYi8klWC/PsUANjYF2sZrGp5VMRxLzZ5OIMHINEt3E6sHeQQlXzxHfTmwTzK
lOMJ9eBxxU6si4Wp+OEXty6esgJMWw8cHT9W/sq6GDy275sGkJOR9ZxPPM563QLASSDF4QtoYFTk
n3OlCrpQez0zPdEyFVgx/4CUjwu8THBJ1tycpW41siW1P7CuLBQV46zhRWEKqW9BfE8QCgQcfkeo
pjq1JUvq85ZAnD1AnLNaA+dKy3yGCC6yqitQY/MqmOMxRFi5tCdE/W7wz1X4nD7yHAcups1jfbFm
KpiD+RmHy1dSO3OJmlQk/6LySiIgL6OFpUCQMEB+ma180VTM7eCjHvqfjRjRNTi1Usc6Gvg6j+VV
UMD5v3nAOUf2YQ5T5Wn7Vg2vjsosrLluwtPN2imXk6r39Qa1yHKKWw37wfJId8eL7ZZ1EoPVDVfK
92GUYLbxrs4dZZeaDsHsoMivgEszN3pL2I6ol7EOYzkQtg6MMAgEE+pfNasZfDtyXqcrkIOTBeS+
YUdkIwMpAzhboyNHLMBw5+rS+oSZdmwWPaHGqvIopF9q1nTPYhymd8jJg8CrbYDRhpsK0LTu6tkF
P/gPSiMA+eqUbeJTG4bH/xi3IU9xXLKlWXKBfuTBNvLH+5JZOLeuvIOIKJEnNcSuh8sGN6GViGs2
JDLmqU9y1TrYGmiFL/M+dahvSeB6JDbm/XO1NghpXYmtQGuDU6SPRPUgeR+MRyTfjRSCZF7JMXCT
9nCynVGrfxFPwCblhWBNCpy5qdJW1hAMmpmEFacPW681J4m4zMf+iJ5OMbYES83Z2PdPCgyJGvLd
c6yf6pEIg9VfUmn8r6sY0qRD+Ims7VOesdI2jISawRO5Q1ETQB1EH/f77JOCkj9gklhF6FoNCyJM
d2uX6u4V3C7N2QydDNWKFmh3d96iWUiC2szs0ujirhKy6X89EJlaPBXHIRJfn/k0tMMGQ1/96Dc4
D6YHcnG4LMXNIERubVMbE99+HGwqiLuROjZLlgnqd8Mks+ej6G60Ck+oXHobnHgUOLF1N1oqz7to
7bcrujlKnhmnhq2j4jPT8wDL5tjTSNcykZv4TW8mR4PYU6eCP+ptD5IGuvKyT4KMvvBZwvRhHbww
rA63kKqvfvBE8ahH7WGPCwM2xbjnYAPX65/TSsPJkqsx+krYFcJaD3+SYDltabxhs9m35PsFg01F
j3NzLwpGcmCP4SVuS4IBixn+tkc3MSwl9z6/YxSreS9k8D6A9q5+RTOrCrxugjHmFqkeeLQ39CkN
xPZYrXAD3gqS6pfFHcETaI0UjLxML9n3lFLfWB2DzPOZ+N3F3NZOGt1NG8wYsFH9/MBqIKT2rofQ
s3p7iLPvZImHZ5bl6/HkBhyr6sC+L6m7hxvNYNP7A9r+BuOenzwB7Z9U1g594V/MS7Sn3yBJ41G1
b6lj/Nyma7mL6CbtRbUW47omJFCsmo8dEb7i1+1jwsPClebXzX05p2Vyd2VUq/ZqP6T/4El/eMQz
fGsax5ud5zxc3Ry6VT439Db0TRmYOeVzJlUw38cur9BSE2GDlSfJqmdO920D/+lraOGWGZReH7ZQ
dXhfHVpKIKqCpIO+d3YOfcs4Dz1AsRp2+4MWkm+pHDPlOr6bmcTxHXz9CiUuEuQWfSDH6/Hyti7M
2AkTUzOvEtaI1W5AxChEvybrlugWMmKgsXc9Yk+DlQQFno90Ie61kwVyAZUYV+kjdAKy302eW5gb
3OmmYgOhPziV73yXR3Z+p8gmyaHMHfyuCejRwf4fRjcYGVEpM1E0MHZENvDeiRwb2BCrKmOj/+fi
EVfIfgiw0CiuvT99ZRPGVwOokmTr19OwuSdld9fnNFUe3ZI+CloHlZCgtX95P7Rym7BQ+6Mh06Nk
di8s9nPkXusm1PMYf7vujWuEVVJlFoulCIIbZLa+xEHzY+PZaIIW06CSl17BVDOltQ3cBx6eb4VX
3OyvJgSGYssqSvJLRum0AF08mxS+v+K/xDpbcMOVmNksXQxze0wKMmDV/M9B+t+dBChzqJ9jiBtR
yizkhywxbMnk0t8wqcdPcll5rA1e4d3x8yl1Y84/NKES7Ml6RnoRJ/UcCLtXubJnH1LsExO7J9X2
Eh1lOomB2zWP2hHYpLskTcmoCaM7yNYHVmf2FoPcvgPeUZtqy+6vrPs/w1UwJUxqO97X2hQM8NLf
gh4HjJImwMjwG/ZoztDUDMXrz2ogPLrfighoQeyjB9tYyghg1ey+hCyMwDl2rxJXVtNTTt3ab80o
oxSVgXddbkgOE8IxTuHXAl99/q8yggT0CC0FUn/vvoAQx5qmLeky8nbK8dnJgw7n5BripKtd/pTQ
2X6B3YGk/ZfQrVp4pruPwD8BM0ReWbALsGMEZJCL2qP9OOda9qJsu+XKoSFclfjZ+YUUc7O7amAG
prOUU/ggDsoNjMMMBH7yHuA1PwgCTSbpqfZLCeW9fHi6KS6wf0MFnMcAINnMevAy3y6uxPnQ+Yaa
6+X3UQdSIlAWkcN5heM1U6JWF35pjoQmq6Zikwt1ZY0+4Qmp4T8k6ioQRRMWLSUK/2bT8l69gvrJ
W4ppjqBvm2qpvZg5SuH0h17s6Gc1cRE4KF9vrU3eaaDXASIpAklgofVs0A6PXtCgLGk4emj/t86X
Fkfivp4jI8NmuN3F7B+KvBittrpJjQ5beebA4gbJvp65sVdsGacejbcZgCEF3GSuP+6SB5rXs0hc
T/BssIJ5iTK//HwZ10llCvOArHzM/U4t+55vEb//xE3IPINMxxcgFaWk5pILTP/rb0Xh0RjrZ0wk
jGraL2965C3Y2d563eg1ErymSM+uLwSAVTYti3D4B+FsC3xKXqlazRJxhofgTFjIt9xnMZWDOHiX
wOo/OJMqEOkiwosy5skO+OSYJJqe+dSujQfePDKyTQ7mmrT8I3n/xOa29wO0edSsNdLsyrDwLRMZ
X4niI01MRudlikBsrYdVZt8T4CSOjYsTqXjoXi0UJhE1z8PqY/fWR+HJDIvhm4bbu7g10eFFOUP0
imgd6q+jiOawDQDlZagYE9bRUmKgPKq34pZ5sf0PeoR2+qyPaG4R3QicmRgwFhEsCHt9OSh+HgXH
Qp6ZAXwGWwA0QZ1hErLfe86MkAvDlwE0gshUYpQmZSUmSsTCR0eS86R9QrmcDTN5EJVXnMVd/KVS
mv+RO5Vrm2nUt0f6ZBCjAvHd/Ea/P44rC1jn06w0/nEK3mAI29fADr5NvoH0+mRzsErBBK5Rdj8q
Zld2way5myJuAdG9+etX6BgPVqwFiLGp+GcOQum8PrJZDHIFFb5ZgTDtV/J+E7xVK7+lo7esyeS2
HXvf0nrnUH8jTgrjJBDw3jSTqO49bfDuSzintPbY6tbUrwUn7zg9Mw2yUrxGSJtiau0NyvUf8Uq1
0/UorrMhPrsWybj8ZQi0VHGlpbtYEZpzi3HqHj3nedYmNvq61jnz0ToypbWHvPCiiSAoXoXpSkVL
zamFzxDhcavb8KiQh/E/kYrJMzeg5AD0CkWQpGZzQQmO/Hj7zoyHep+/uRBAWbU6tJFw4acs2ATa
7AdIsbYetRbxC3W0lFmgkKvzL/KD/yOKmcuP74ZL5/ZYUecR/CygR+hMh5i5Qa/MV+XOjOpGgaUx
uZyD1J3nB6kDYyUzcDsxMkSfGfBUJlONE9ANEY2aXJ8dadKGUQBZLMuh7EqmMeRSeyCSN7H8M17e
hNqrfRzAkwcyg7Q71Prhl9hVTlOmXjwDnTcRy6mQc3E9NBMc8s2CT2v/+BUUKRaimd7YSrmPNzjO
k8SZRDxJDIRpOA2uIlq9+gxa8UuprdAr1zKOFGTtCv/RLy9iICf8JqEv4TMDEt/96Goj0AREG2vt
EBGzdP2QCcZRqksn2bC31ucaVVQZIKJpxNaOihFMfGqYM0gZ3Lg9Nb9v3sN8g974j9gdENhAOGPt
qox98Ee7uQhhOZhEZ4px7IFMWktTtAZ6MQlnKBI8UVyW6F+9XK411mh6XOQFUuSrPCEuW0SNqGZT
Y1lJ6do04wnmIHCmsMlwShqShaW/OIsLrMM2ceO0Ye4vGygneSt3lUOG3aQM032RWq1qxRsxJE+B
TOy/umqm6Bu65wklPM0GRXWOc7JTZfJ5tN0yJDNNahlwbnvVo8Oc18QwQkb75K18s/ShWl1OTUIY
/ZAEBPXfStSrvjCAHNS/4Rnz9ztg+TmNwrje9eFklD9Gbsw9m/wy2LytenG7gGOLo05hS1cgiQL0
kmyxsJgxDUstTP5zOM+JwEXU9F1Z7NUKr1evCCttuKjykD8uHpwqOamzahCxUzg+XhPDOa9dqHaK
JLOGVqkPcMtRxPhbpZL83/d2Vevmch2Sw6/vaP+mYL6BvqbKxdkdZ1QHojZkCAdCuOVDtsH1B7tp
Kz+vVIHyIFMBIcHj/1ATwx0y+1KcT/6EkU4Mz6FLLNJO13h+N3XdBi7DdvsdaDr7FJw58IK9VeRr
4B+xu+vigvPVVusH2s2l5wlhCmsNWu6QgePwTCSB3uN6b0yZoZ6zLjwEZpOVC7YIxuyRtveGsp50
zl0hu5Wv4olBO391M3WeEChELH8UIJGIlhLJFgM9uhbN2OWiTmfmsIhepkeXyYYGfStSDkufgEu7
0jkEagN70pwHZrU/u+0a5/t1GHmg/S+7FcX6IaSaY7seTJwI7c3QOasUTiPKGy32kwVGnwVyMmaU
MXk3yVqDXfSoSWg56pPl+4SX99cFzT6Y7IdRoHeXfAFGTNO6DqRsmb6iaMVI7mpeZCivmb+wrItX
pQMp+4GrQf3e5NlzYopVKxXTRKIIJXAxcwkgH1soNXQjGLq6k7vusv7/xORKvKxdX3kOZzY+/5Yl
rhgC/PhqFYfFdh2+CHW4nWQxp+ZbGqm04JuIQYlD9ay2gGp5LR/oLND0yCz7j1OutYkkDIi8CHS4
YJvmcfGiLZEvqVt7ryctdN+Z1AGQsWsMTFDyAJ1SRhwOvkInV1fsSOLu5rYz5gti29kiaIdM2Egy
xk4Zfubd2SgYfs3fwGrh9hEoHPxCoIJ9PJmhm+9t6KmEasiyP1pbFfyLXMwrZ6aUdG61zjyh2ONr
dZpPkr0lb1CAbdK0mMN7CL630g8iCuyg9vIooJiXeERrKuHIk4ySked8ognjBkkBTxH3p7lMH/3m
9gM4OG15qh++0iR3PjUVQZhmVFb6Wo+82AgmOAQKdjZGAw7WKKoaz97VGXec+YxRP3mcVXMMjMbM
h2TRcHr2+m+0pOr7/dmq2vzBh+DZsRi7MoaxVi642bHY9f3WIe/oq7cUZ1COdBmZfM1iFXehltqP
+X0oFE9PbLhZizC/XaaoAnu9TxcFaRfn/V3aS2LY2xhk/XNJfy8UEXjDtiuGNu96O3k7K8w5S2fS
KaOS2AItwkDO+sT0G/hPmc/Fz7p8kwdugYsnSdVtLcAyhMvGprA3uEdZ6Tylyo54nKsSI29vzxsJ
8gM6CRJWJj9OJXf5K1+8xI7+8I9MQpDfz/ImE8XlzmTMVvmd3WjsVdUfvAn9IScKb6gfe6ughukb
a4z8CIj/cKr/E/sChORQf8F2nj7SA3QRaorvvdvVxZ809FWqrBg2YOsr7INxbrrfUHy1X8sk7ChM
COHEewBku6MlGTm09RPElEUe+sLFKT7FymOzBimfAuXEnSPTLI+I0szVbqVbg5Y9UcFFtkc+KtDe
gnORcY3QvqDS0dpykeJJMIsy237Qa8hszXSDLgjhMrYaPY3cpydV43giVnhnjNI5YLIAAhBzgYYa
yU/GKzyaCWBM+f+fns4/J0f+5uo3ojbTx4e1l82OaygUADgGBCgxBVfVlG+EdbHCyYuM57SRhjOm
S1ILYnn60pnIZTksojPI8Re10oyPjsiFFyV6SnOkjotef9eoWnsmh9+ZLhkoMBvGUrbi1P/4+MsX
VEoDdiicaBtzLAXXzBct9UN1TerfVgepqUjLg73mymnjQAVWtLZZPFvG3LoBqo4bXcLGp2k8HQ0z
+1pEoNVkerKkcYxLJ5/qI5ch7DP70J9IzTBBpxSv6qfe2DG+HeoEToWR8zmeJNALddqHdp7fe2DF
GTcyqJLwRXFuWu02p7kioSnCQOJ+qMDih90jp4LW+jS82vOt+A2kmkbk5oAp/xM1IT8KQenDukJo
ZcymBe9X3SdxkURPEbYl97PlyhPRMKfKJQhmAAh/Ivo+WYdMn7RqYHTgpXsulZBapoDRsTCs5gwJ
t91RBismTTHJ+KT56SoE6gx2obuUzgiG7Lxy6umSOIq2TIuWrhNkZnbYFst8Tf2df+iciL8BZUmC
k4vE/ymdLNHFPaeovqJp4YaQyi5dj8ib6cLKj/byPakCwxiAIcY9iz6YwbEaLsIxp+yR7uVqzryk
QCGMJxhtmT88bBg9QWFyoMCSijymlHSFRMgLBrd4Th1mC3mwxKwBcLyByADws+t3x9k8bMe4aOGV
cVq9B6fR0LcZgwowTOro5vFhzOnPtK5Ox9LB3vZ2ls5X93PqxYdciejx736Awb7QNPp68wxtDkrr
heOuTE5nOYpc++g7Pnv9Fafc5dC/ti9IGAcRJ3k6Uc3wwFW/HMsRmRlojfKyOR5H2NFniXK9q8Ab
HXsKVOn9gVAVXS0XOs17LZEUa7N0zyiGVFmuNfOdr/Z81PTEgJniWUoVxUaPTsB2XEXE8yhTyFFh
0wscK2ZfRksh3A7YX+QXHfntdMjqsjRscHZOSAP64H2Ls0XxOhs2CkMGnWqCzHt6JEivGFBiZC6S
hhp9M9viDPaqoYr32Vjm/UXh+pk4D4zAUfoTfLIimGIv8ALSvRLRTZfgdKRRHypjp830gKHHZCJM
58HSx7bjzHvHNWSNjM6R/+jscn5hlcCH3A48CgEIDczWv21Vq7rHqINRYWC1zZ0eSJ2s76JdOcL1
Ovg0FriPOG4aA+k+D7bB8WPcKLd7QFgHbpCPCk8ZfI2YAeUbquiMbfYvInZjv+f2XIXsz9fKjvTF
tDMuS53wIFnoyLwys9X+w8O5XPwB9wEdd+a8soEf5ckRlwtWlh8utILYUP1Nys6119nJYjg4/F8S
cd7NUYzxuSYDSa+TGxiiYNLHo8zTQrbMPuFFvpaJwFS+gGyf7gXWvbQM8WydI8zF58oSIwJfaepP
Cdx9MPOeArOTFjO7/Qpc41vR4nsL6HLbZ2DUJ0d9QCOSlXjwjSWEKD8XArh+g9Wf/OeGtcdpqqOF
unSio2E19GJFxXhj+bcUI1+UBbe+uvbV3NzmwtzbyfbnhSe01oIQhDexg9B7S08YeWCixZplz2WU
aNDxI2QdLS0uCgiL8+kVPyrEyoKyYQixXXD0WUEFsq/A6SsThwr3KTcsJzdM6KXPMyBqvMA+NxiP
LMl/s7JVKpslt+bWvJX0tEIw4oYQk+1zNIdVsBGn6LR0+l/fnpwgIFX11St4vjl0kYCeViR627rJ
OvDYCH9LrjGO93uLTGq5QXjE8qA93NAI1S5zls7Ml0uYAoN9XhP3/F22xEITwmaAGpcHJTkJuoLQ
efQQLapMhpkPoi9cNmSJ7vbWl6f6JOQqrUfZpcElzHRVrINq5hxGEHY7fIJj0y7OJTS/oBttHVs8
VwrzV4nROqZAHDTeAMzRyVWB/DxhcRpgBIbmCrznArXn1epLfoeQ7R4BCLqk2f9mpRSW4bWs+o0e
v9sNrhZ7mrCrQFmLlWXAetT/d4bBG3jB/OMP5MKuMr+7KBOTEY1TroT3MHAMCVT9Vmft0i0LZ6WN
2plN/uay83ONPfqnaZhq4Qa0jPdzoArAu3YH0WCFKBRrMGSU/Ilyp9U9tdtfYMrC1vRlAPwfGbXA
Hn/Yz4Gu5rLoDQStmB1nq14BY2kUHTjfRjyqxNhcrWTR+BOdsiqzPIoxzPJDgRpcgFcTryTVKgyv
8JDr73yp44naIBD78JWeRzumJtHi7c2JDYjt0dTw6LRfu8uCZGx3tqOzX7921ONEXKl6F1Y/CUDd
J/XcHbPYWWnLNf9U36tY1RobuQ+6/4P6Uq6jk8XZdkDLiI1wsYL3ESkbV19FTWKB4ytGLFXO5NMA
qTuAqKwc5L+4UIX1cbfXNvtReXXcsUALc5I9U6WUoP8x5r5oaCHY/ySDwx0Dy6XrhgSgm+k62zDc
MfZ5tNC0HS1IbrdEi6YgJGPFa/Ej0I7AHwP5yIxpM8lcLbmCtvv9bH+2HX06b/XZzEaYM9QzYo05
Xr1r7WG99W+CqclAI1nmisw0b0yPLQGVOAdmtur0CGl5fWKP1Hxb/PMwmdZMUY/xblT2MsIqR0VH
nXrYewFOZTsFpmYygSGOB3WNVQ0vx5PmjPMRf8q96CBPsBAc8q5GI4Ki3MSd8fNDfTqshPnLTtYm
kqvP3889PNPo8pkovwEh92DS56IVPxmwzBDrEpS6zsKquBYURpMo82KqQXjyoZGK2fx2OTgrcCTM
mLRYN0ccWijiCrNNl9fNCVNpJ9ddoTvDmqb4dIMwcIqAx0jj1v6utwlcFbk+AO/eYegJEtuCCSef
pKm3zKllPfFeLGgs1Cg4df48FiU7l7fQ6OIFngtRLDirUDAufWZNOZnikQpUbKVANhlviE6TggDD
vtItHFaXFnu4EXgDfQYzCqwgWTSUignRP3k1IG4UxRvPU8YYLaq1XJDv1QI3iCa56GwVO7qZDjk5
3Bd9J8o0QhSDM8EOBi8yF6fYZ4j5TLnVGL64VDsmsTSNUcsPp/1xHhvidh5bGRHup8/nt6/WvWdd
qhKDDXNM8t2SVDFJvwEWZcBxVNlGXsLFbyzUm6IMy8yHVwikzy7bJDJUIl5kB8XfM3o3EqzkR+7V
6KvD2DO1VEnIyuPOccyLf9fKZRl1s3lsoRHFZ710sxcOF7ylv0WlJ6I0kpHPN0YLCnqzpl/aPoaz
iRliXD9PvedjTla8F/p6IorNaOXBK+vNhf7+6z846u2+cvQNHpKCnCrz07UqCtPZ67N+dDDvBiuf
RNBuovbxzcoYL/lAlPMsgdu4RoNBaQQeeR+encocSR9cfZhg+afv3y410aTpf7sQQjj6wT+gPl81
eKRJcIdUDZc7lOKl7uGUipiup7N2zppzSkcxRoftd3L3I4OIC7TdQfb4ZDrAcNhJ3nk6n77MIKWt
h7r0afi7yJMzvVEMeqs2Y1iisWCeMa6+tWXeqLmgP29PmstbTu4LgaN59TR+OI8Cfi4hM2qQaEMP
UIfEzRzYYfMWXv0nNIqnEgz+XAv0S8L9v+kRjv18ZlXmaZ/ya2PJtpgzF7vEh/XPE5bN9r1+inHh
Qs5/ciWpjFZJ8UJK0W+k9irLRu1wzFyz06JYfmZqGexkzE0mVG55ALUUixi2YiYZHoWmeBOXjso4
fpiWwJDyAgKUrc5/znjh0fpDzAzNE5I0R9tmVkc38+WO7nS5lBMvFmaFZmlYNQNIC5Rx4wthyRpy
rDjKALPCHRyjalmMwO8snUnALVANtF0ZBQ1HYKqdwEmVKLuYpEBu7Y8y7UaMThR0riGFn1sz6nxt
hdZsCnV60dUUx5808szPay9m5mgnpMNeuLrDFJNHcIxidnoH9qb8/NMC70+bS5HvAnpn5ygRXVhj
uz4WE8kAMBzqcpKlZNScHCVhGd6HGcsbG+hhOVPb5v8SegcBhY4MF8+JBAYxpJl08xN6c5f2ZZu4
spAK7NExrMakpPmLYK/Ls1ZTkNswnVU0bKCnCnmPVmD+wMLkUXA0qyOAB/InAzhLPHRucp26gWPY
wlW2eXQPWN2uW8MOg8ZVeNNsrjRtPmYWxJfduCaj4qmLllH06aM55l4DoBwdO9xFjSJa68znL0+x
GCakK7fj92HgFobLJ1G0SzvBJZbXJfxMbEneYzvwdjJh0Fm95D4YpQKLc0e9WAAMyMT6WoYrlC7Y
xIKzU8iMTuQXiea7Zy7aSBoAdPlwxCMtE8d4Suytx/+WjrY+DHxBC7X3zBdgH+bZgNhTKcBEOu7R
fNC8lQKh2YzsDp1lWyJOym3azo3XVpPS4SUBzDsBuDK3IrIy5Tm3gRIk7oKSOSxfSCtwfAO/n8F0
8wViWbwy077Fj+mMHWDXUTAffvRAVRDb6cnXDgqoQi9MXmh7X+CCMuEuXyDX5Hyx1/G6pr+p3bsR
Ey09Vw/uKUZb3BzLVfT87gEt5gcqdAPPcG3cGZj5yfpClNOfGucOFekjVOjEgVgizr1w2BlYGN1V
gcMRH2cv3fCQBAk2HSly1wDAPMkbocwxmfbptYr6NtwEGhBUusHHf5MoesIByTdVx/empK8JrGdH
f1+CrEzaBSMm2G4hvg1Pkk5+qTWrEwsb94ISWki+NfurWQDuhvPRl7H3+FnGtkRGIi5JRPnivgai
Z4GYzqJ9R5uuEzsi98r5J5GoiDXAigyCDolOjaoNuvNsHd5r9bs37LitmUgoaHFPCh6QaWaERqV2
BOxZ9fX0A6AtTy/YMzW/XHBEahHRzzLmbenlcudoEvmTnInt5weT6Qz9NJq99gC0JoHgJU8jhzWo
hdsb24a3SAKZAhijonfG8tkAFgTcLXBqF10rs2tSNorcmltxiW9dgUMPDzgq0NEHYFTtukPpfttS
KZRpfDB0KBz3IzkvS1vAN9EONIdbxuYqNsjD2awuCUKrzo784VIc77prWK/YsIiQYFnj6O+2I/qY
9bu0ahbFLy9GJW+cWVOMm3mbFFvzmzY7V4o2aLvmDiZ4o1n6XzoZSAbUG3ntr6Fvo230BtH+KOCq
mXfP72U1J5GLtQwEW56I5LCM3Q3Ueh3ZA8/77YiC7sa0RacBa0GfjfI8MqOSXNSeL0sGEMy+tauI
nuNqqI0BT3qLpeAIkTHjudgjEfkO1iONC4vzArgBjF7KpRFLSv5ez3YqNFbRI4CpK7KTezRLhAi5
2FQ6FQUNbzqh/Ku+5eC77YUcbjYmJO01lJd7ejlvYDotr+gRrFtDI1wua+PGbJ7QKvwmfmSgBKhD
7iuUJBpMVv304sKFsr8s8lzyV5orOOpE9WoaS9qz3FJDeHwZbMXsUF5J13IFHTt4/dVtjaBvpHOG
1IiONke9U0JU5bPoieqbGKtL2r2FLoB/W/02RwiwSMlpc4GCxxIk4vN7ABscdBlAw6SyO5MyY4jY
TEDOKxOl3AesRG+4vcxTHTNtY/lXqZX3fKBX7bp92dJ0QtjMVZuQIfFV4NiBxNeKPOHWSInjwK4K
PO55RIxAX+cLgbCRnel2QOPEMAEjtHkmhVY18eswqwRPYffB4WRVyKE8BbCLEK1UpCIuohqdPrdD
ZhTXVZaQZjGdPPSnEFlcrL5mlH5qVbHivq7c3BwQ+Z9EV2fn/46Zs3MmO+5vybNsURAQ9LYSQloL
BRgKePf9YKlaW8QEqAx8aaWcF0WzrU2L2TSIS/9SiTfMuFlfD2mmmq3g9y4h67mfh0HUUDogeB6f
UCumn5+TR3qi5847Cae0+6jacdQDSkdnLiemvNNmAK0dgVuaZ6qy7wN+DP6vV+BbfFsJq01LEKaK
lvHlNJcSU9HuZ5iw60xdulqvlGiRwPqrd06Vac8kSbFydmbhBEmyyRluJiurbTscOmJH7/q/Ldyz
C0MpDbt6ypd6LHRGzRH2sOlyhNY9vKFMFQ9/arn7OT2lOrIZtC6dQC4PxzcfyadtCmoF9TlKqGaP
G9vg7dfFWEgo4kHwKyyQcCurbrcGzdYdvRE+jlqUzuzgdMeBQ+HlSB9xVkqWtMcwzpHX8Wyj5EKN
UtPtydz1hyRmz0e0wmFgZOH4YjfjfnSmrTzEpVysuZ7FDuVTcfrmfmvqL/YyDUMBBEJEGL4OXFeg
Jtdn4juIq44KpWmY0l0dUhIn/lkbL6iuiNBhMo1gMTrZisaI5QAnyy103qTcljQxb87CIgRFK+84
K8v6pTJOMy5JY2xz9/7O8Rwq+Eqsa3XN2+/of66xIhtyGI14xnaaIUGoWGh06MqTrAGd3BLMCWqC
OPXEruANndBA78wdunxdpgy3ZWUc3HhacghadPPV05MY9pimrD9MlYjj044lSsSZ6WS9i2SkV4AC
ywYvGXA/1XCXpSFlmFY/xoBzq9t1TaZVK/r4nw5EqRqLfKFQO6QCE1vaQ41PScy3UxwxKjpTzfpN
tJUQZ90HqlcT7PBWigWU08DTQWPxC3unn+6Cy1MWNeNvqTPdL1IHFRuLaD7jClSeVqMTZuDkLx3T
m1R4qvkUIAU2eX39I4SS5PxbHtO3LkVjrUnr+ts7vKKJocV875dFVIJLo8IA3v0GmPt3m51TaqcW
gYR1NPkBxB6Nr3dbJKnpkQnzFoH5irC8pDV5ds4tVRmRAlkumt6Cm3sGYku2t1fOXZiKibnu5j2Y
NqQ41r11Lu1bd0iqbTfzqhD9RsD+V0MT8RYzIBIam7lrctT4AZaFCtKgXe3t4QBox4PlFsreZ3Go
GjSynhIbtCgBjElMPPa8D65JevIHEVxJXZXJ53dXVFlVZA9HfoKMmJBM/xY75cd3Vl7cB/jUTEwg
8h13YoMBxNZZK9hMyU3/PUvi5jXvRWYU3loG4CWmY/BMbW0FSFPeWfYPiKiF4aQ7rd2YkM0YnYFW
+vijZeSA3+Kd9bngS/1pAvNvrhLJ99OajKfD1B7X3GnuNQgoi3ADMeu2hoIo7ahaS92k0L1u7cJ9
O8bmrCfbU8n9vQ3SbAPyh0oSymL0qqwG/4th3+NOzE9Ki19XoqhWLthOmpbY254wMEVQPfmKkXrm
WQHP2hvoDz8WYF1UzqMIsb3iP0AnIyOTLGbMLEqeUp5QPhvGtF7JVdNbF5r0Bba3GDUAeHpnQHC2
vXI55LKGYiWw49EzUn7Ax9w/n8//poeZ6Tq0OjdxiKluGeBYyW002+wYQqvziYqrpyFdwKO24TqB
mUNxOg/CHagAP2J+7JErAt+u304ikLHQ8nXNtA2ltl1WpGnLj2gXiXFl4KnPDnLnazLDUkezKzOe
W90/JWUzq7VCCYLKQdM2Q21TujvFO+BgTY3nQu4q+HI7O9PAuEG84vEE0y5Z49PEfI8tejFouqVX
3VLHALDFAnhnPZTPNz6hAiE3MvuWSWWRFoKQ1dC4RmC2NMjCw4zebszAb9AaSO8x19X8mRPUAv3E
vH9tliILORWeeoD+SndGLpgUJKWn+sZTrVrxgCFO21Vfujj5G+1QDf/U4Ga8c3YHQSBYhUs00y2c
D2kGPQwndsqdSWcXcvHII0v/vYMs0c0L1yE7vpG5E2NJs58NuvJDEANJh+qv2bcH79Ec5oRVGcXT
IebJwxT2qrHJFBguDuGaOFNtHVzJH4rzrucX2v4Omwcze2GxP4wq0fYFq+AjxBfV0MAjLFa+b5LO
MTF9oepeZ1eARtffeuBA9HzqBENUu/JWctzQbZE3gSgWHaRyHY6PQmJFC1mkRkc2OwhwDZMuNA+6
imTUn2h6P840OF3bN0YWUm/CmLEZRlNdDP5lTKW31qPS5jtUnV/OpqqBe1N6SLy1sDMW0E9BOuNC
J3LYHaLIh2Gw9y2VCcD7GobCHoYbzodIj56v37ybWAUgpqhMfb12xM62d5mEXCUzg8hw5dtRyNwa
WEQvI0o8Kv7ddeJMuSYe4WHM7U8zf/CTade3Ot819mzuKbz0qb6V3CC0wE4xozgHvjWA0zRiLSrr
KB7AQd2+36EpIR/cFz/naE0DruI8/MGQjKuphDhHM1e4+4U8FCu55QRkcqDk3N0i635CdpFDmW2e
WYCwQnT78m5WZrGfvprurDMzvGZoCvwQdTOU1uVb6ZRG2UlxZ5wAoBz99wDOLbLmK/fDlP+CGU4C
+DgGrbM04Nt0dVjXUn6aXPbrZ/nq0ScCSe70d4TvpaUspPFwwkphxaD+eLPoNNpzKGlom1a19kr+
zlgyNIxG4mRzwRii1+gv/COwOzMuYtUfEzbGH0YX2En1+x/9KooQ8IXYzThLmBqfagakceQ/u6oN
1cFkZdSkqa+ROuYh124bKpVDiXJlSGejRdfq4khpEWYh0tsyp36vv1sJ4B5DSp9UzH66UgjRLa8J
TEmEyJUAMwJsI18GggfPhQK+70AzBS7SoeCs0xWaVPmc17dS/+e7zqk6Fyg5E3SAnaNRl5kyp0+6
uZv3gocWtWbB3KtamsPzKKl99kfzLG5iYYoULtAjQBm4NnGW5Wao+0NuN5CUNvCqukORA1MOUkl2
evHlq0ilpMcyIr2wAVynTiZ4fjqtYdF6O/7Zbcs0ASz0wzyWTGygi1zKmjkORocToyEB9GgpF99w
44fwadgzLnrRXYJXqkrmtAZnwugkjaUHB9FH+ULr1R7KNSOwHMOLhMghHs13HS/h13vQ4OLjYz5g
p5vyXtmb9B3X7TS894CoMGPceWuzIL+LhkCF5cdhDWwrvhNSicuLQfZozZ30DifUyDQ5Hemt3r5e
lQ673mIlF4IKkikrLgvZbuaWrZ0MwBpqi2wIjoK7941Uotk/auVq9bGPkPXLdz783UY2Flo7ETiW
V6Z8ygv7qmCyzvqo30ICO3OYT5MXfILpoBncXpvVKo1qQ0+KTx8geuDAgeTrfcXkDzeXV4bfcmD2
AhKL7AOu84ls79yjNhNzKS2Y01aqNxPz5/fLoJpxic0ceI0ZOkzhw5Wnxm2FADP0zNv73rSYmIFK
onl/wxipOfjkp+wVnDZnQYRAaW50k17cLs5aw1zosxwRl8KOUvh6B0ln8M+nL9QMDjsrcGHuAgvy
BfbE15ll74OQqTTdgY9nAWsuB2JZnCw9wVyAfj5qNtINUoW7ZN0+JSX8oWjlb6oeAnG285keyafY
CjbuGAKE4W6Q8eVoxhjT3saS+rn3X7sxs/D9/ZQKMr3iHCZX05CkKgVnXa6PXhMRPnwGzru2BgTU
4I3PeDsc9DYEaF6a+ylOqvvfXR2TkAcadiDftd4v7CeaXOgJDabiwbq/+Z7H9LRscUog5yTokF8C
VCTmXnnra6WJ58vdUJAzcTS9HGutIabYK/N2WrDScuvVpxuT79WYpf5GQoDOB87xAXogMZkBp3LK
O5H3T7bntofROqD//picgFbvUlFNW1ePGYDjX4UNIUI77ZGIjpMEVjyvjRhVmy4NmUqf07vj3ZYQ
XChIqKWn7Cv5tyv4EqRgc1udplJ+07cX67t/84aViavZqeDiVQcZQae1MSuzdh66k6F+4K+c/4OP
FVQJKfLFZRCaKBr364lA963vazgcLumnvRrEn+aFGoKAtVFPcyz7IR8nTMn40vxHQMtS2IAMSHVk
sF+ocitbsk63gIPDcAEGkEUkyXalL+JindWmIdT5fd/7xe2zykYEpDyyWyFJhYJT9/c51QH8azrP
AZPCR6i5XgGmyMZy4z5LdSkgrpPd566Oq4Gu9ZxIjtBKmn+cyLxwS9bBzdPXMr6AGq68Z1prQ3iz
wkb8z4n1OVaYOciXBjqkQdUuZzDInis3VXMpi2vhuwI1wuWqU1YLY+ildffn01zWhLNY+Zdq0MH2
wzsr/YCl8HL1mBgmFoS1inxGwKqRv/9IAroPzvpW8oBCPlW6f2TRsrRlZuJ4J8GVwwFWIedLYdhx
t4f3HRjps+J3ChvtPW9lGRtTDv8/U6aPDazwLTh2ytXzx3USk7L6qZqRc1XyWbZOoGv/u/zty4D5
1GJF/eREjaum3CjLgCyktoR3Sv84hbkMeP9O3LDMLML65Ao50a7mOP49R8dq0uoOc0boqvVizrle
vc/g/645M6fAn0pidVVHst1AzLwCipfmhE56yMbIsDLPp2VSAkrdhFLkDI2IN5FHSVvA3YOhZzGi
//Oms2Vu7t40YxLYWwUCPP0E/Mw5G0Iy1pNNYl/hy9O0dPibxZw8Cd/MxoxUdlZr9Kk9ntPsOvb7
iqIBf8qR0d3qZEk/mQRGLHL7afIzWHZWDKTauLEyVX5v/An3N3i+ZEfMrg/hxl12Q33xLKEwdzA+
/btfdelgMOuJOy0HAZL4jPHtAm40r/a+K+VaNsD2qSYI8YU0Ez4wTDd5yy6PbpPzOhGyuhdnsj63
/mIpz4O9kAagTaS+o0LAxJmzDD4rybPFvR3dt0IDcE082URzC2YIhpdPd2zWprBu6KzjNEou2Lxu
Re7P4OZ/U2u14UVfym6ykKUKXII1LiAzaHzVvaAbsN6MM+JB8mQERLh3Yx26ZbBa3qsglsYaBfpd
P9yyMDKKYsI00tx2nbYLjmvpRjJRaL6juiPrNm4Uo3uSkebtn7+QaC1LhTn6FKjl4mhlW753JBq1
AKlohxdlV2++wsG3KZslEiZeat2OR+lzWtyHlwVJylimuQZChSYDnGwhoKsjjhbYDqDdtvItlya4
kEw+wvF0vna+XkTq3reuNal6VxIAsXPnqMkxMuSmveQB5ekKrM/2AT6DdBwQ9cAZRgdj6BguH7ce
8M4CzP03E8w49F53aJxwUVlvfDwAbuGhu/yVM5u4XurJUPvSUq5uXgbGNlVwzBaH0NgmZ1OuGS6f
JnOSER8JlIXip4PELr8RQGSCjMCrQJz3/jts31D9p50+caWwYQFZW+Wl/dwdr4tjp3kHk97NC379
jcdcFAaY99rs+MReDmbZUyRP/GwDIyumfke8LwrhUZ0r8MMb4idTwpBaL+RKc/xXhc2T3Y0sH4No
c7IAGn3dY23/VoSftBEhoShPECEdueDUhnlvrgK5XMYeLYZ57R8qoKlGxDF1QzCNCqHyr2Tq78zt
0/qqIwb9sUu13xRMtpAv6bR/8t5S0efWp0DkXKQ/Gi7KSrNxOfFg776RhpC/rs2wS06u8Uunngdl
kyuJtjsWrQDYlS37PTHRFjxvYa7z/Vftbq3+7eS9XcXPRbdsPSKc4F0m1PHl31L7q6moyO2SdRYJ
1zofSLk0u87HGujt0OnUO3N9WaolNBgpbZsRbMYwhJp2mGrbuLiM+8st829ed3s2+jco0jcwvE95
agURsKuW0YCEdCXh4KCpHHCPneGU6qqDO2EDGDlDrwvpGxWBlUBJX8N9d5OsNpRd6PI27N5fT3oe
48xIn87SgdiyuWzHgAMvT4/vcd1UmSF47IPutDMq8hTf8N6AXGN6uItXOuiMhcR9X9VuYA6uvNCQ
fIVZfiK3jzjQ+LvX6zT/KtBqrkY8o5hWVLc+Q6rDd6JsbMeWZ2yu2+REJnBA1WeNO4FhqGt3xov7
4QPTsO+zDWM394TVHmrZiGKhY1jC9XOC1/Wnthx8ECimBWQd5bdCiKVKae7T0hlAXRllOCE07lsP
X3L5UV9qHIF4i7BlN+1TAFTZ6Xejd6+yAexPI5RF2s1oi9kcZgMUHK2R99EKUb6jCS24Am5il+Wf
lVeYq+b9A5Cb7i0cxiHxW+SaTKWQ5jU/6/cLXBx/BdTnzzCLfixgKpU+tjXHuPmCsIrdYiSXAC6j
aEn4q/5fVKdasz5R1OT81bSuva5A7KkWDtQunfYKssEe7dhPR/LWfwuiAlrgqXKkb7LNq4fodNJn
UDap/pcozi78XcDBALIK2tEm4jjyxW/W7yE6XXkmG9MV6H9w9vb0rhUv7hbh8qVBwZvA3eGiPryP
KnCfqXrCtMqSGLcO4vlwqWgS+HHH824CUdz3fZrP6MyQ0JNqlwFmFFr1JxEK+tTk/rzURVL2XFer
Bhgf0vb9PvYSW0VhxCHszV/ew3ARMOE2iZPhmO5Lxfz1w3pVJHzvBUMYwV10nm6SyAl4phMcEsTO
O+P4eBdMJLp60g6TPHkW+4AV/jcsOT8cMINBL0qZEFk1y734U5tIs/lPUXMNeMZ7ux9zXkxjhU+1
IwUI6wJDB+LHDM3RSjPNkIHKsr53LV0h8gK+Ze+cmGxIO+ExP7t5FVRw6ET0oeQVuwb4j5UDUW1q
s2Re0uZkhLv+KDpKXe3KSnuvXbAZT5iv/5StpnLeCRkEjAvkX76MUUY1fbLEXmpZ3sN0pg6MlnFK
RfdyQrODQ3cy/MHjkxCHuHtPzj65TGwMEL1IX+DtisikAkjmWxFBk3Y9uAM1LwiEumkSndtTqRCE
/6nB6zYAA93LHlDJLUT2zPLbwr21B5hLuKqu6t9miNDyqK9Zau9wInEet9MbBupqfPisLcsWOUr4
Zn9eyMChnRQrp+gXHieUdnrAy6jwdhHzWAGjiXnGuCggdsoalZSv349z3P2e9mk/jmbhnUvaq+rh
XOpWXhSDV6/tmR6UPqbL+MiSOEeczhbuOA5JGxlmH5FEPiEdsUnKqZGpcLGkWJsYXbpfeDXlK3T8
r0CCU53V/CT3w36sDFQh65jsNc4hD5KVXVk627+zwljPCUUOKZlTZunIItPtmZ570XTLD/OrH1Z/
B7/17vdN2O661TLG/1t1c4p/CS3W5smMGqsjEdMqT8inMI70+TYUuTxsH/iM7hxS2XFA19qGAwd9
Hp91ASL4ADKTfpJa+hLzTG8voIJE/SZ7APyCA1wOW3RoZsRvVBItzXuoqZ3KKTtxY40sVzisr/ad
p9oSwe69djnUKbmMEzQJu8Y8ryCwECnL8D1gFqCtdppWdtMc0egj1C2cfEMyI5pFNAZcJHmntEYK
pLROAlHj4S/0bhzrE4OnDHnrkc+Nl6wiVKJwq0jTUayo6mHopL5s9tQrOsXXGENh6cksnRFsTglo
rhUIPW9D/7oAqJ72jVcy0FzBsBt1Rh/no8lAx5qK1VoXZszlvbJXY64r6LJTB5r02k9Xm5H6DcO9
1VXrfys+TgLlaoXE+oawPbBU4ZS4n0hFre9TroDcTbhpomRfRIN0rm55mW8qXAjsV/D4Sqpw5KvU
sE+tWcd7aaNUyftP9vv8zBWdNSXM/FAYcmCgPCG5QKN+n+DfWmrNrEkS+RptYW03eBhJ+wj7n+jG
EAvLyKhhxLo3Hok0YzDnuSSfMVzWo8J52GbeG2xcFUxRwSBzd2MernWc0ebvoRLpz+yMfjsjIrXR
oqcJY7UHqQiHnLHD++8WuzLdU+vjCxpBcALl3tZL/VzC805BWbSJJIWi+jLBUYVhKaJ3VlAIiirF
HVuwqCjJ9SpxVTX0ItgMZ+yehbPJkAMNvEwr84w+D/s+WCem6GVZnNbZh3ui/EN4XhLhuaHCoDWe
OdjNsC1/pBxR8BjN5TK4kEY2GFEmlK/cFwgS8fCXReJMon60BPeJOe8zvlA2fNN2cBRvaTMckMuS
MOy/mfN9pRgmrJlW+4qC7i7Wivj/rZLik3Ob/kc0lLsJRVWcakBhfq0jctwIKdLj6qS3Iuu5lsIM
F5oh78qmC2PDsttt0TdnASW9jc+jg+njw48hx8RGmTaSX1eKFH2k/6xW97bXExMEzQBbhPdJqRgo
wTZ2wEEmfJBUHy0Z21XHgUQ+9yDpTNRbC4nKHHjs2Yb9xwAHgZ5JwJNqkUmyGr2ns38ZYI0jP6iR
8VsmL1+lP5XRloI23VPt0uqdO6UUna8lo1iI9JqU68sQf7bpnMvKORAueEFQ4JTIXqhe6mXlnRdZ
kSa4iMI5JWr6dll+UYmYiCPL/nY4l1DLpiJco0K3uRYUX4FXpQkWIuDhTlY4EQVVOq+aZk8RAD7L
qJEQ/pl40NgE0erHQzeEliTUyjBZWMfp5cpH/H1TBIccUHKyJ0dhq6ROmEkZ8Zftau3+YjD7qzLo
hm04cqNYySbrKTmrICEf/34rivjpxcVSkysY0UJhPPwSk89iu6ulBj0nC5QKtcU8QB8cQavIeFEf
qN6Jmx0EwYE+K78se4TfRDIXwh9eLuayde0zZOQ+EDwpMwX3oaJcq8ihjgNIFItYBstrZYdFeP8Z
K+h+SPMXm3uG1RwdIshPu+wGdkML+asvv3preWMWprPMrMDYX4kbWQ7+Owrodqs03GgxRCVSwmTF
b+YvXsRHxAochISTBh1Ji7MKmrrRZwtMJBLPudULW7Zv56nnKXqczDgsVtsZvEw+jq1irnx3fIJt
ksOHTxxjdnjd/G2crXymBmuxaJw+g65dBdhoVTw7auhStzgjNjLD60NSgyMr6fymXRhKpy2zg9RS
FSU9Fdj6EJY77B5rfMxRbjegDk2TsuTGxm9JZynjaSXFgtlv3GiZkrpQtpVQKHzosvOdgql61u6X
MgCB6BUCCTcec0HO1vD8t/fylzxE8o66f1VVkR9NifmVVenM7CeNhkqkyWVtyerfmA4uVltk5yGA
0W+KoHsOkiVrAfi6JdVWNJXTfMEjwMc5somvCJyvlhWXdInLVdIcWA2hRsBA92pwf82Ei3m7pxku
NmqZJNpe+n/f5WePGPzaGK+GkhNEwBGQU81HOtevIBEYegOY9I43RGVd7HZGjxzZzgBSBjZRazJl
ZToXlNRdWSIdAC9b41Z93DlfBMX7M/g2OyBuSlpVitBbtC54NsfobIlUNq2FEkitlC+hm6dfhyhE
wzPXS2YyvJev7z0kblYi0w2A4rGB5ZJVQPLoAkCoKRB2I9svJda+DawtQebNvXXq2WL+NW8TA9d/
Sv1oKJl862Fj1vf5JbvrUK+88OuTH+/CaHexOQDp29DysAPzhaAEG6kfxdofyZ3Ui9okfHS3qNNU
4splTSANbDNiNcl8VGTsa9LitMrqPdmIZaKQboLAURomUukLHVDGPeOHiIV5eK3CRqqr31IKOxvO
sGnKncLdJwtYqN9dPstUOan9JkUrUiIk3fcIObE6tMSZ3mAUAX9OUgez4LUlE9uV8X+LN34GjBud
NDlPF9luBubyg3co7kpCQ1/uQ0+mTpuBHJEOyHIC/+6cpAYnialfebYhFbKVJhLjHAkw9GLWRj60
ahOxItNFWeS3U7E/thPgkxm4WBpkxb1FFRc0BaR+XteFX3usw8JQRN4VYw1ApUPOmDPEftc3J1RL
oek39I325Zo/+CQ6NVtAGVR/UMaJi9mRW4Faa9uUzyvxOlO2HRsgdx3xWYWvrcziWYXPvNXHunBF
0R0X0qT3/kDxo5jDi/LseVaU8Jf1jbz3tQkCUKnbXp3+3TPY+M1iYzod3oixqz4zLw3l6QiyeeZ5
UfOPh1787Gt23xc2cBfpLl0pC5uDQbhPCRklDecbqdAeE9gDdl4/kiBedEi3l2nmXnHvUh7Oi7tb
uYVjOMWtPMoMcdnJTaU3KsNPjZFyNmIsEGFrF8cwHPUH8jqkdimT+/TtAP36CsRHCfnWAiYszQEn
i6WrC0SkznjUljxNVwGtSDRsjTf2aLnIcgiqQC0jar5q1bdBlFm+QsVUBH9TLagxyq5wAtrGkWYG
u4LAFu0BYjEtfDM7XHoDOGwb5QzKgtvAMoZbtsoXN7GdHpd6qq1ugGj6chp6yMzCyNUJ4JflpXZw
mfGl5Aa1+NO8ClkoAZES1MrKRmRLOZrO/MGwlvXEKZfUP+fM2mlIu+mquMX3D8KDszETDqrNknOn
m97q7qxXHQUiKl8TqXt+FsfeLx47/CD7rPVEhfgtQj5wiWcQVZ9Aq62FDxc8haq0/tRi7m9VMSJ5
Nm6zx3cPFMUdeyZLIKTY5Y6hR/gq8TfJ3OkM71rQENYWzRAZhqmg2YSy6MU4hrE2JuScl/Eaa1k7
1H1PjoJhbZ87028POSxJ10qNjpb6XTJbAH05Gq04CbqLJKKcs5C2z2qInKmQtdotzIDGMif4zqTw
Cl475Z2PiYQh1M65O/xDPWbAXCaWVNuGCvqLveiyFNowEHnd8kopEdaN5RalGFM2ejeRdfqQ0pTw
RRzAnj8N4i4pxy1hNeKe6iYZY8SrcIGKkxhTtLR5Mp6tUAGnsa6N+zBRx0jxPAF0WGaGJJEZ0ytL
OFeIy5Y6bDaZD9+Nyxgxwhr+z5FPKq7vyQPGLZ++bhl1TWIV5hya8deQq2e/t3nCqVI+oSBExdBZ
sRjfapE6vx73mvGrxfNpbfa6lhYt71O3MFMESylxlc8v+YLOpWThtYujkcSsH4yY8f/TgXDVyO2W
TrgQO7QEWZ4ql1Gu07DgwqG/FYbVW/3AX1Ap5Z+BNnwlbargdRMfdyzSEFZIvTaUAZmpgqOyyBOB
r2uqncThNSLItaQK9lp+Zrzi6hVSZZsGfq62SJ837Thji5dRl28Y1wxd9aGipQAEaoiCndHzG553
qZqvEoHUkT/4ce/U5MIrQQeoSQXg/prAXdMSjlWZIuMc7jaG5rBVQ/uDDXAD/v/02IQd+j8qrfLD
zWj71SLeafBBW6y4WX5YxwEIxZ0+rrYcaL780wVtwip7dN1u/icvzZ6t0ZhNKe2PwsMzPMxaawfU
jeNNBSh5r42Oaf19ZCIwMGD7QlQu6OdLI8xKJcm2RCreG0NyNaiuxfHU+7xfnVyPPL08xgXIU4y7
2MujEkxrjevw4d5v6LjFVyWcPlMIv0wuijGgRahStLuD3YXhVgDiPMOjYkA7WaqnLUNDmbtqphqa
+vyBRkGod01j7j0FrOPwrarGSXH/2lq/jSseQVPYkn1jCSpt7QNvBHWutv38MxcxRnt2Z7+w/sbU
P46BtIhdqbjgPdmbk8QXol5XPHHgiLsszQSlKiecRvXaoOePYdU3vt19PFvjMj5GCL0nuyQJE5TQ
e05W1JfB4UGi8SiINfBffIBz7UAwu+wl3nBVtml1VmwZYNOhVKC0/998HnJ1TYSK74p2bzpe21bm
MPEtnGxw2DQO8Cj3a5oA8KP7mPf7sOZSn8ebxKFxrANdlBiFcvT5Bcjf4guOD28ML+4CLtR9/Ngq
auE/sPeYlUrg8T+Q9cgivK4ZEKWyFUnqm23sVNoBBoOLpJMx/4j4KjwBj0ScFX7ak7j6KdmM2HjX
y4RfNew6YdTQqJHetCxL2IfYvIiBSDdYGWZPl36zY710URaWv3coHymRjfAjfiSKK0nGRBjuTw5b
OFSH9jWIpblPbKIGuGwTIshKQPnqL0AP5cbllrtu0mGdBbvewkTPyXQDAwNdmPCqwJCXojSbbb5J
y4SvwFG9BTHeaBPj9RRRVvj5MXGvEO+VfbVyxesV7fjb49Gepo/2xe1ivMTYlSEBrS49Vtv6K8X4
oZwva0cUTsKgkKUdhl6ycdXR/ii9T8OttENqYVLuarcheWadSQUCMVT0nxULEpJB5HEWXtbUIIiW
QfCeoeVINTczIwpzfaDBjdIu18PyfMM5RfU1BffOSfB+voZNSYqt5NxWMQuNBy6goN7ONQENwfuF
1cERNKsJlyWQKq+o79l7hAaee7/WJOCchQwKuQsO2n3wYbrEm6jWJtyMcX9sVhw5Np7BoPNf/NyJ
ilnIIMJlG9LEFMQvnexctutHmTsAHYonleYu/77geC/ELRP4n8Kwu+A920Fu4MrGpnHKFaSyZF0f
jW9BuSN7mhggc//UcbJ4hw4xWgZ9mfpqMXexPidLYP6PX39XuDLUkHyWNeCDFvIOrsLwKPM9zIAV
umMejbkMP6+eWbZPa82hqZkmudbGFkjj1uiRZ0BWdZA51H532KueIV5PKHZHG0RpSVNuAIIxwjrV
36cJRNxHElTgQ9BMMlWp6nNFNnlCrBRjTGrDonccbjKIgqP48866KYO5revsQ5Pd+oCKaq+luQ26
b22Fm1BvvCKImkIHcAK364z4BBbmqXEBQa16uXyx1rfPGGL4C+CFRsY2s2+p/tfh8okK2H4GmR8F
iGpJ1+Y0Umfpa7yydluIE+tXLs1DtnoGxVftBx3kLl4BU/b+hoEKpJa41zNNjEOhQx1UxQr9fTX0
wWPcKQXcCTU15r9A8JJgF31pZ2LhP9Mv56oc6EuQSkwTQwgO1ZmHVbV7VtMvkOD6U+RpxVLar7e9
8dFILxw31T7WhGT+qNHeEgi8HKlwJpLtrUNKUZ7ctudKvk4+MtsWNpKqTT8F1VT7lI1k2HWw3Ezm
6KtqJ9wA8fuBcCiskHqnv+yBXvNRkK6RT4TxO+osErMXfBxJo1SM43o15mHBvl5t8ksdZEJDUPfP
BXtDjvhY3Ycwx/NfF3phJfoznKDNTnHnyMOcID4zGpT+4PHd1aT+7BeFsLrhxHAaNudPeEiI1QuY
flnbXX5VDjcVDVukqhaJRg0ANEy7HSY1+OkzQ+xYqn9PA5XiI92Ydlbbz5wp08QjAGuIcPPwQD2g
UP3g9VEkouQeDWDxco02fbW4CZfMnFwJZzaKoen7P906YVff8Hsdzo8z72oINniqkCTod+yntvz9
L4nkZeVjrKEnNvdZCeXQtUemLdhub3y9IR1gPkd/JVhobgkft0MaJ5bD2QWGBF0ZdEai3vYg9/qu
a3rJgvJiERDqebO1QvvC8wPBI89SUOHkz7AJ7H3NbgHoh+IS//qz0+U0Dbr+O/0jc46d8j0TZDk7
Jxs5orET2APd2gh9x25D7MHqp4UvXAc9tPlo2F/rBN8Q/SMGQWFBx6qBUoXFPNizBX23gyku9MP/
F1X1mP0UwpDfICcyhVbLED+vEHqiWK7FWJvL7O6bZ0IBiLwF+AaCv2A/ggxb7ZQM9P+mdpFuaT1l
oGHeGPv+JD1fkT4x8gGWbxteWKvteOfQY1YF5+mq3r6JwgXZxVW2/Ewl7zHsfUUJCcr2POESKipK
Wv6pJbTtCozUKJbMClyybfDVMIS5FUR2UBRBFWddo3rv4qHCw4MUSNqp6T+hdyga2II/DtU6xMGn
JmP4cXlSTRNb/dcj7WkKBaju/UTRZS1vbEoxTwBKT4H5LSn7k1KLVD7nlZGRlA1pLf04pD4Ng1SQ
+uCvfyGAf2y+XqW4W+WXNTj/8aG5Aw8fIGdXfAl9ANp2L5wwp53Ey3hpNtRspmXCUP9aGvhEL9zO
Rjmge37kJ+px8JwcNUlksfm3m9+bBPkyFHokf/FnIhyKlJxsfGVCJ3vpU2AYjmZYIyGLx2XRzoYX
SBM0d8jm4LAe6+jyWyHt7IXuYioZ9mZizHY+1tKIauRd71A4szlpQvvsNkMk/kQ59r0X7g+fBn6N
LhMRiQm4q+VPXRLUnchKvFyZNc3/egDTXMwhrVmF6TvI//z+uwpomUylzsqEljk0GGcf3ExKDohx
VJqVwlMbcFN30wAToDNXtBuG2+Cl9dEOyKNcMtRDwWfpr5McvPS8Bl1cROO/i4+2EBrLqBDox1Al
pXqWgLzlwUuZzFkcB9ogXdxLvjInRL3qrWADr5dq7fN2lmvi6MXTvT9baJYpv83S7Gvw7laGAzki
a8Q1pkuBqE7av+btuN0UxonMY4cOvLRo1tw+OSM6GMWm6uqUMujfsiSHWI01xe+vtKfqNqV2okW3
D3Rvuxk3ePBg+shVvWD/Fj3gpBFOmeMYYLli+wCwMPSqPEcUUH1aCvcK8rVMf7y6+WkFCS+F34YM
58dw8uyWbZ89Oq+94h5YTlYHM3yylR78ST1vEXlw5J4gfTAKgS8oJxkMBbf0cfc4yvC9+r3DHyzQ
cvOmm/YHszLmOP5SFpMmS5j0zjgX6SylRG+78aiEBsHVJPSuTrZAZfPW5EkQAeeDtoRjWqVH1tXk
I5EQvorsFS2oUE9KhImmaLILzYBOG6m+E/Z0k6Mi3gTZwEaSL9svvxAijnC1Ll8ZPqm+WKJMmcZL
ii28HLMkztICSxtOYMKcbibMnXkcp4G+89hO8NusG6RDsg/D2p1U101fd7sfWrFnWqQ2TMwH8gXn
3sMnSRfrLRT2uZ6K8mCvQ+WVKuJ/1ffkS7VEjj9/sKJA3anhw48IUbchg1u95nCzyD1omAMANtJl
C7XVEvR3o9LYP9zGLKgBuvOKGm0HAADXyLDgvcG3OXwJEilBQRobS2JjsZTjGP5LwUboOOzE3ZHu
8Oy5fEHtUODzSJCZ+lYy+HZRIFdwOeIrxHtWN+sCUCwyoD4MbstmJT9lBdEJIaTFFBl5SHA1/A4Z
eFxjMmrDcfUyhmBQh1/FZCGTJBWznB2SeNZloVB5vsMS7RqLu5RtPWVWF9Ny1Z8cPGNz5mAOJCrT
cDQeyJgoCwt+/2JmFzug0WgDkmzCTGoWGlcCJHkvJQB1kCDk4nmm9WlbLgWhM2p1r+GrzG/IPyu/
qBOxjkv1b2vPWS/VvFNR0INx6d6OnrYfjcizi4vd0WbOQB8RWuFypHjfzVYQE3yPJWW1agSXhiaZ
KUF3VzTYelfd53x1IzpDydAhHn4coYjq8J0oUQoe+zjMnZs0lLTZZbaC2Zl4my41PQSnXSYkVjMS
LWhf2TxOVljMQPb5Mph8FgfF+wEBPrw8spGMauYKtgQnDMw1y6i0CGbnqHTMKwg14vTquUKB9Kol
9cF5zX2Sp/wtB3JXom7Fg0aKEztZiYuHlD6VQ7jha1X8gx6bKqEGk1WRTccqUqu+zlns9cPECP/c
9ZgcS5I1ixpj1hmbCrQmR7cl6J0f2lBBMNdEhy1FoowW3yG/f254pn59+tqKdtpEvv/+RnsY8bRr
ETjnBCxX86XsKuh3C7MBpL+Pv3EdC4cVL1QIRy1eNUR9Q4JSXqQKY19Z12jUxcryuNdC1WsTd4vk
d232arPuRrPuprXyWdjypd+mSYe46sAHiwGZtnwqnnbE3KSVIcrnlqzr45f5iSxRgo9bULx8+ef5
gWYSH6sCbm2l7a+dFut3VkJLgCQlgW3rxdUHzt28+yiocJud91Jnqh0sq6QIjK1k91Blm5rBRbyB
NoQH1Eu/jmVp1/59KKS/dGmEuNC+IqOBlTXidNb3l7f2mi01bCBPR/LLfA85A2Ldn3Cmfnz3SfLE
k96OKwA/uAHf6XJMcX1F612nfbnVrUsZqoRWWy74BzIFjPbAza4LORQSXt5C9yuQbNA4RnzyTZ4E
zWFgCUNjFXx4R4eQOgNmkYCheiqiOkszFHl3LvMbuOJrkmXaSSVT131D89+TW27gocsVa4+vUS0E
9gOWTxfuIoHErn7hsrxj+dp+cDBiZWjmyAooW4nFXY7E7nDozDDW6pU7/0ubaokF0ueOBVG6/pIy
qYvH/FkKJjviQMhLinmxOhMBYt5zpizOk5KwAWf+lO/muWqCJB6FzfVY6U5rSq9hKkUeLmZ3YVNE
eqN/TpwderZlACj6S0Fw/dxC0iUwn3gJ8Vrkk1Fo4kBhk34zCbXxBOacu3h0qe7cAHQ/QY/wCUF3
FUQoru5+MJj+8rfUw0s9J6gGm9LwCIVwLP65Pq8aEiWwilhwZ6nNDfwTbSwvnT9Gj6Jq2+rCcs+B
tU96Dta1gbL9W32/TZ/diKz1ftPZ/XuW1N7DoUB+LIZOo7BUmqHlsgn1DZW/3tgkaRSRi8z1EagZ
g7Pkp2bsOyJLo6LY86p0T8lBHc336dN9qU/pTs+thc3i/M7NDSOiiuFuPz3DXauFdVo3dwYu856b
69R2z2LSAbGQ4aC9NrqnAYfE6yLFP6rlj/MnC1ZZMDnY91sd7pyGTRgpuwJeVcp6Hqex4MXt0z7A
COlqrxCotRPJqeSkk7mNLdtFQkGD3Oy8eS+dwFxK2FHKAZa8DFSt5EW2Cn2M7mQ2PGbT34aOdPDT
0rC6tTn4fjo9rF4BYzBgeR0yS+zHQeW/oylCBExQbt3fLEp9DasgB5T/Z2KeaMKMugsntuv1KPqw
Y0boQxcnmMjKxaSePzYvZjimatNgVzG790HM+aat4kDI+Rfp20LEPvby7LjuUOeldyiY4M80Yizc
KQiHO0TDDQFexz60WKXuSkrHw9Ryb5PsmvjStANtHjm4bnwj8Pfz8I1UwlX8sscjVHcyYTqpRsQR
TItacVbJ+sQmYNZokeYqF8cKgLEPp9An46MLZCmc3l/5FUxsPRcLZLfaOGeYdB3EaeSr4TB6EVuG
1li19kg26UM5gCSFFkERE6qMiotppn488+CcBVV9638n5e8PtTHt5b4+tJtIDrz2OoI/xAYePUnu
juBSgw2E1asvz+uITOdVEHgRDS5+DuuUR16KwzROhRa3H+pIc74RY4DVVdPKdkJy+K4WbiCaoDNb
cvRd2CqOzbuXpcBIkIvRbr8VfiIki3ua1gYt2zSCh/OSBlvNUoinH3wz9KSXteQKhD9/f873RNzj
0wkyevNh9TLgscSMsv3xo/kEqkzK7zYGD1xk5gkA3WqYAkXxMg30SjCsa0fVDMNzYgEXQEFkA/VT
tGgEei/O4S5Cdm8BzVW0uJVPvDF5h5KE8GGEryuRjFJdMV7eNGhocdXPKt6B0vceaboHMiN9tI5T
SJpd1VukdGswmVl1IxLIXR5KDh7ZjqLbjWNBlWvg9I+mIyfMNxosWtHvu5+IkgldywiSxR63UcCa
BEpkNLH/xkOKkzZu92wsYMGmkBmRzB3OIUh5DhNf904h4sIvswqZZCboVznMERcOPuvkyvcDo8gA
8DKfHNKKGDY3L8Hd0ft+/9BGa0OYbRqnZWlq/Y37xEbx2e+tou0WInU91WMivPU6fGTDpeIVHs+c
vrOZ6jRt4qhR0x16jy32QRpoESITJoftIdBGnlwk840cG8zofOcOnEy3JPnEKTeXJbPqGfYUQZoS
idgyadeRMgvDFBXjFRxFsZsiQ7z15TU1J7JSBvxmt6fDYSoaaDZvYN7mD6j7rKWpwU/harTxoGRi
7zOq0ZEZlv7tjeyJPzy0E7XktaagjI8jJoRUNJZx/4NTPzngv7ZIiGaPNGf9xObMfOdXRZXzc0cr
GcdYNWHj1tCnx/UntGubyP6p7opj9+L6r5REdZuZXdLpSfmou869/vmWQ6Hp+XZTllxRCBnR1RNj
NH9hcR/Jq22VkKeVEnXWRBFCwgCuzXBNoMLUI2PHhlhLbn1a1BwSJHF1pJ5pBZEbFutzoyX1fEDO
z+lUOBuwLxT4BoYT3q8cL70054pK0+MVFsgUY8aQfI2ryiNiuh3w6YXetQPBl7d0SUy/8e+fF87M
LHiALkhwR0INMWCrpGxoxRQ6/bNXT1WC0XcdXA4WA7EacaOwG7EUTkGKLxREGP5J/4kyyWXDzuYm
p+IWpi+j9fKesEYbGW0hIfH2b/BhEOCR0wrkaSmL+3gs+mI7+QgFYwQFzY75R3ODFMRJPqq2iRSH
DgoZAp/ovfwCzIwwkoAnOGcQlFbCTYFr6jxGJ+6FoaAHlxDrwq73PdN/VaWTnNNnj63KN37K97/0
FTtBsRJlcK+Ck+ydQWbE9uLZOhjZdThDHGfR9nPeUxXc1LAtksQzMtUb6P8I20LNs+Yntj6wgs3C
qEPyeqb7vcjN/oAB66IE/SKXLvDJC7YCh9fQUHVN5I50Ux1a7Igpp4tSLuPLT7/FSKzjB3mkVNnf
ZeUFDdbHgUaku12mveD6nRWbxTOjhhS/L/aV44CdlIiyvdJw4rM3Q8JNj2cRgc7zG0H06l9daMKG
mosYQOQcCOfk7vHCM/zxOXwDtiVy6lIHj3sZz7s+xw4sYHWVnrdx6TYuZ9GjnDVVvXXQUexeMBMB
T+I634QTXVqcEab6ixeU3l9G21rBClDLU/tXj+stiQ8CJuhNdy6RO35Dp2F4fyPAVxanDMvvafK7
PM11svM6EgCzPMFRIWxSMa7HTWnnoINStKEoQWlEBFKP1J2jDC7rx17X8LU8bLW9y7zDeao8yx+s
6s60RGKG5t/nfTLPKShpyoJA3QGRa/+pGfNMHkgUiTwjKZbfl4EoAOK86v0KLv/UICZrqhkl0hFe
EJwKGx6jaCaz3g4yg6+aoC2aROG6doQDdRcae6N8T8WWohFxarmxUKFIL2IZJj3GciLf12zlPV3Q
s8b3x4l3nEMTxNUeoNTP4LW50wk1ZfBWs4MrqCQCfXT1EobYpujQFRfAIo6lM+OG1pecBuCeWv5i
FnCOEi2seCO4ocoDDPdN7h0ZIaMcDqGRG1PYjzIAUc/6fa9fqrjgjxI+g0AWLhCg+3vRZKDN8Ccl
I5b9ArVYcCOmiSbk3PKTYc8fE+WKlD0d9TU2ynoOrhTtWgLl9nDWgbJfOcGRJy1IB4ff1en+3Wkj
EWIOEMIPWYlYySZ/YBqZhTX12CnqJKydJlVxVcwvDh7inYSiPM2SoAGaDWfSL0jLbioq5YWMvG6L
o6gjxRmlZYle4m4nawYE/Cl1UA7I5l4HORdPDJMU0+vBWWFepsWmU0LNOVC1nWQ7sYPSmoUgJs0f
/YfPnLgMCKu4wirWrIs3oOp+tHDQ5O/9l5xZ8B7AJXWlFYUk74+bAcAoH1ZbtOWsiwdaB03jFbbb
TamovN2XtkOxk9/GOac3McG+jTk83C1HPVueWvt26RLtQ03fvbdU68lyFd8AglQZrn5CIH8ZhpMx
Hoz7DjwmgJILiEGjV2WYNKTEF0sO47Ao3hn6sZ1hrRS4Ijk7r+TZcPYtn03rkgJsw7lXvadeGbHj
NRZgmJpFmgzBvMoBEgjT3vTzwl2wAmlnw1KKhpO2xnU8TmPjX9tl01I49FZJEAZuqmqcr3WIZNjz
gao+QbHVoCvU/PksRFDOpRHbaibahlG5X/T2Bk2ED6BBk75y+Z8RVSoOqLql3RvseHSXgjDDHKZF
RI27kYIwyAlVJRVs32UvUySyJnTrug5K2VqlfGrqBsvheEhrpREstm9G9beNrwg6/v+oNRtp9tFN
P0hXy/FuYWsQdsejRpxQAiyEgpGSpG3l3Q+DfXFL0lswlE8rIWYqfwB8OvreKCRoZiokFo+pZfmN
aXEetjLc8e2eCL0fi05C0X+HHMHLWq1R9xLjpBL0H/0S3z2cxMOxbmldVt87hYfy6C6xb7YLdfvg
tP+YZSi9a5mK/1DkSRlOItXQ6yfC8TSf9jGfWnDQBsQQt35cnJ2XISYigC0YuS3BYfSSQvq65vrw
8xUORGnIRmyCVAoWu9ugjGsahNpwwYUhWYakSXetdfBAkiFDJ+NGyP4HRy4S8tmtnfh3IBE0+uDs
TvgUEqDMsier4hfw13TlC+ItWvwsYiNt7EcJyZ+FE56IJITzKw0KPeWs98h80CP9Qi3xOLNRkFA+
BO/cDGgnxewDpXOY2Gl458t/+A1cBU+NDK7UkyzoSBDqIe0Rbp/5rSgF+2DdQgR88OL7pqUidJlO
b40PQEGhDCZCphcqh/8pBqruIPBsT7sCOF3zQVVk4loCZ+4l1+i21JY/sPKvK6CfiDVi0L67jCAo
etowFwOW2+bap6T3gMPayYz1ZjjlBzVNpyvWmc5DlSxz2IEmVuIspKnn1MuvByqlc7voIFDqpR9T
Bb2OGntaca4O0frJFw87ymyyHVEx82hbyfBzgTSI8+bxpoSq8KhFwMaLC2OHpnIm0m8twruVSGjB
HAOrwZFf4iHFfd9kE+/gjp16Y4NGIORb9OEqpxCyvwAYYbvQXE2PGbnrBGAeQqSpeI7hnWlkH0HX
skZg5/cdpKL1cymDsaoyhorqAmZ0eGc4puubwT6LrUs7dX+BHjHvNSfk/HU/+KoF90oosxdQAnfe
ibToV7+JxXvLT6psWYz2mQV25Yzt0aRO/nA10ljq3zmNE+965W1CO0Q6634rcq8TI7+0PoZfjlJl
YVdmORZjZQJQrZmBdvxcWe1xCYv43/LoguX4Whk1uLSMfU2BvQNmUW1boqIKIJPmNW08HIrioRBf
Vk5IP68zz81l9ThGwnvVYXnyoFZzIucf2Xwh5ul5bGF2AMXsNVqdJROEWBGoM/JijxXbw069fN6G
TaStXIimVIrqHr+ASoAQT+ISmGnLBx0z14WdRwgLUvE8Tpk2wi9YM3Sp+gk+rGMPkmknjhIqnHoV
Fu15ATnEkelpsBNPv9A3+PirWAGin5Co2Hy8S/Qbdgul+4QkI0BQxesbys+kGNsp3Y2vzdUshMRF
QKZQiHcCRHsV0xH9TNCIlKtCUOirSNImJMbPBsdh3YHFDKiZO76Ns7c1K5o8PCZaezSknnPi50xF
GLcm40/7OX10/Kc61qg98ZeBX76gj9ABYwN3vJb1DzOY+DSVg/gpPBKdYJvPZ/t0dWxtSeB3gOgD
pXrAZlm11AVJHL5h+eby80jJAYtpf3TUumm/oobC6UoCEpK+PsEwsgDQG8MUMWgd/xbCrY3C3vuJ
1yVPsFtbe5DC+O7j+qFA9wBThgF16wm9ISgiwxkBWWAHvZ8lEHDpkzz1kyqr6WwXaHfbOR5BrQYH
FnsTIldxy1SeHkMlojDyEpGL7He2b4UBazy07nAkijLzrpb70yOmGFY0PLvMmADIC/C5mEDpFc9V
P9SIDqP2LWhARIHEsN6MY/w88WwzJ8g9lz13hNltKGTZjL7550sCKHX3gqy8oyI7x7zZ13E2u0kV
HSu4ER1N5srVLTvOlG7dQJlnuInOOplt2YXWxAvlT8Fi8toGQoJ+0c2KMS/X8P1lbLn97aTnD2rQ
6ECIjLX6zsHv21ZZ/KK7Dk9TVSIFEP7wkbzHmDQOcnjyC0RQrjvWKOrD8hFymK9UNp8+z7XkYdBM
8HL3Im3GnuqV7amOppGJqrIUo0p7ScR0Fnevjlx5tvRaWy1/y58uG2PV1uQ0y5uEtc/fWQgFsTIO
wLW36GgoE1JwDkO+4kT0f4w98eqWPnXnXbyzcqwnjiR4gO1iTyCI8xzmG6B0ed8KxurV2fT/OgTg
n5G9TlcAeIu4QRhY1Px0yh0TFXFRuiN2kLE/bSDHndyOzjFPFWHZFmg8PiZZ+CUS3G98zVMHXRQ+
PnkS0sLplUAiIr7sx+4VEL9asHqFDw8b7sXsibsUGFeJ2qQNMDmLZC3mKXsfcdwXeW/nrBxg5wKH
kJSVBS1UOSiIWNI9jtRtWgvFSIIwzwtrCnqLN3gAdRfGjClUGbYij+IfkTVWYuOvxOEieo68OKa3
Xl4AqozT9kbZD9W8BjKIOWImjJ/B9fsylBV+WHCA5m6Vh1qrQKzGk10+UDDvDfqGNHbrXLmx9KOc
uBdZeeIGiIsGbXBoPU4j2pCjERIFiB7JorLTbAJSWxiicBxiuEMzgIOo2zGvpTgS5C47TpO4KMH6
fEm2jhWezwy73BZ9qbAfWH5t/cl5h4cTsmV//X9KW8SabU9dwa6Sw9YzxPeTcvXkr+usdQnqOA9X
2OBOp7R706oKAcQjO7w/Z651tjVe3x6PRmHvSohlrfd9nRrmkEi30znKonjUT9qhbMFOobuXxP+h
TKvI0hX/FvR+c5PjSCND0aC8U9TQHkj2E8UmcDRSAfuqghNsWuD6N69jICoXXYLJXNJzbyiYfyi8
Q4MUTsVUezMqPEhMpBYXEYSHdLw09RNr3CDyQssX8u7/zcEuQ08ksBGgbsDyRopxFQ5ErwjNu7VA
RJnK6w8FSSGDe6/41bMh/+Z2CU2mtBKSyYyQf1+zTeoJvg8Frc29wOr76euS04n9q6T2ucTLGwbB
YxSZnUmcXoCEIz3iN7A7CXVdfGFVcSEMpbrQH2rvVIUxFSXKYbHOgYp/ev2+cRW5hMyP/A3vExmC
QujpTofmk/GJYROxuQfxMrpdgo0CNWG588T/Sv7zYBAao1sQ7cXXwuKce2qN2Ug+MfbIBDEXIRtH
DPbCqrzZwty2XRmE37md9spNDRfRRfOJLxxxB1giMxg1khUHrZVCaOBUCp3eyEVW/5sFEexF97JK
BZcoFBQxrJGQm9ZphyytvcFB/H4OgHPBWtR/dBpYN1lExrljKLNR6kNO/gwM/c6SHUPxDX9RBu8I
WWlT6Rx/65RVrphPobFdJYKE+gGtG6oSaCYlcz/2wDQ7tPL9/Gl2f+Nk5rVVPyHna6MfIIEwm4pa
SehJU364AdwIlYMA+X8POR7XJBqldcAxA3ZkliwBZSlWva3dcDxeVuOwdhOWDUyQ8wV4KaQZOQ5I
8VSSV0q6BhiFA2NY/tENUSEwqgyEmsRekQwpNZ6jXxPN4PIYNzXgW3hVaaSe4MNHmQKfw1QNSjmn
zFryKCEk0VJRm6C1Dal6VFQsoX2c1/trujJ2fEc+/CwcPzbTAGHAgDBCQvSzeFdDwHL2pHnP2VaH
JIkM2UYdT6TPtO+4gm5n77pi50I2/Fi2uwRB1dRDOL60MxBjyLmg3SJWVtId7ZlT/VDDI/tvjNMo
SM+D8jt7zwXU/Osug6QWcql7EgqOw8vzHfdOAXXMx+5awnufzNmIQ+tZbRvmC51RqFACDmowFmY6
LZYXnUlJjybpVWLL02GSxqjoSJVZq+Wa3w6JbkcBUw4clAS60n+vhaBfhnCssIvlZYf+LdiMdLgx
BLWmSgfLOEt1Y5UIIh5Wc5QZoow6QTQ8c52AdycH0UgWADGvf+aulTWEQFf/13/gfSiIEZDOzoQp
zFSHwuq9hp5XomUvcpCxCPEJX9xHZscpt/lL1cOYcKb6MirfSHjtsyZNVjiEgZkfPp9PukwtNf9K
e4QaNZLTHY7KWrbB0iTtKNomazLEa+TdGQIgx6QYiACOS4WGqJmQiJLh/lMpRpNa5MyIpEeuX9nk
DejZokwCmKjasHicgi5Nk7GrQRvqEjl7TCzp30pxfPh9JTUxxkOfi3BGKZryBlT5Ge+Ikqx4NL9k
dKEpSg0RsiIbpGHNbPHZCeiXjQru7fF3Ytu2k+U5lyD3Ph7Ibn09YCKPp0i5JmyuGOun64bnEP1W
M0hymtq0nuO5CPUU2zRZ6htVSM/p9qkstXlBAdYkDy2K+mj7kFO1x3fNKjKGqV/KV5BO3v64nKjo
WW/dYfWwKTzx7JkHj/dut/Az9mTJsO9fS+Ih8hhbNygoIyWD3tRobMFfxly2pkKHgMZy9KC6ot84
E9rWjwCJ7Y3JyJajlL01533kWdWBdLSTJYGdTtXB3ZbsWYAj4Ib5Jq6gbKcX8d0MFhRujo208Ew0
Z+YLsHLA35XsZhBh7+IEpij4a572VlqZaw92U3WX9FdJJbQhjhhv3kFitVJNfMA/Szdp6whfQ0Az
tcp24d4PQtavA3VqhOLlfHyUB6hHzQARNb+TqBw7jaq+XoRLaWbWYzUpSNldFrQG9sSeCEwtpIhu
JpZv5aCe6rbG8+ansI2CP8TYArvG7jGQrrjKzg2YnFzZO8tIL0bAF9XgHAl2tUF929bSyGjxFSYV
TwzF0Lyk53PxvYjf4LnqjSlFvde7grndEX+E56NKUioG76UJm+rSC5vXjcpk3yxeAZRAtkxXsbTN
F1tsqTPKMNz0AM208A+7OLyRXuIUyKHsq0Fa0NbqVEX0bNru3ilZGiS6QvYdGFsPNu1NaedVd0me
ZKu07cq6N14gfzzco+PCuc96HaXQ63myUhBQojxVEkR5FKN5Nr54hXgOMSgnFlBf9ID9AnZjAxaE
AR6KA/rOIPyCCQwLY+rdH6Ud9GxwyhHX+5Mk3+47WZ7vkri5eiR+j7UjfqbMCWtkya6n8dQvU4vb
J1QxO/eoN4Ys7qIrNrNAWre/zK1wywsFopJFJce8cPz5CcnefH6SzW6ATJzNLImE9kCUjQfm4jww
sxn+WUc28RxlzIzzTPLSG7Fb9xZ8Gx+jYo7b7F/nQPLePEIzD4iACN5sH4gD30CgbV6xwX7HJsMq
LziupXA2O2W2R4imddOMCuXVHtlV3LNZHFeK65WQI3YHsjFRgT6VeesYimV+jMPPh8UV5a/KYNHs
cFXdf6OsCYgCFAFGO4++fiTocsYUMa5o4YrtfN7iocF1E2rBS8Vdomt2N7tlYrd4modKuZUOI+8w
XebKarTbOVr+ZYe0bj1t007IERkaVS/NK0aE5+zlCW8TpOHVYyiJcL5A1isyKttG7uyEvuheVdM3
+tqzSoy/LA079gyWqbbhCH9MX5YRe/z7uKvxNyAfN5TzdSaeJvmBSYWW4miZYIz5x2zSFnpxlJQH
9mvwsolQuwFliK8Yi/0fLsX6iqqV0JJNzxte7mfWtl3UUP5K/Q/TrGHZnyvrEXi9DoJUVzgBYJD3
OfHoVGh0Pin2t9pZFcGWmkvW+/PfSalV4jFp2+NOn6ONpr/RvPDHAn0Hpi2nOLyw0Qfux/oc04ir
yOG/cnsMnQtLKXZ4/6sSJ8wElyc/A1L1IH+9m5H1nJjszwHLWoQDj6jYDyq6P2akq5zOxhShrAGE
WSryC9t+LtsxpPqtYjNI9Q4z+GMEdZcNiZdgDzW2jSL2XvmlGPS/BIOhhU+dwwGBn0WIBcjwBrnk
LwUg1GPdfI1G8v47i2agYGDQGBxNWYe2x8E/aDXQZ5xES7bGJ+K/E00pJemk+U0m3HVubkqkxP4a
IUHD7reShLPx0gF7A0FrDg9/t9pU3OCChuRgnUyG3Ax+1GsYmn76FEwHyIDMBHQstHiXktegRIi0
NUDKuMyZJrxo9n90l7orBftms1g9quE6RvirMnCZRL7DaFUK2Ghi7IrvBNGyeVl5+oMk3n5/VFdu
HHtxDyjJ8CPka+FRh1AMwYUX5psX109hLniBl9oX0aAyJkSGTwkNaxO6mVA+1Y0UFjptVul2FoEt
kAI3NB6/O1PxstFXWE6eUliaRmQZvv8Cgnq1PGRAb1/ovBeJNbXFaeyfVUAXVtb1F46FvKkze6d2
XcEEo0Ukw+t07X1y6TYwtCmYu/XpYFVNrPhDFVaLtWa3Gq2bkN+i1neTD9WdtNbnkxvf5Rc9u+dH
1CiK4z3y+kDgAWokJNWFkBR4nxstF9rHOY1gvw60L+cfTKjPFcm+nRvZkDNooTNoAMMMkj7Aealg
C+vsGQUd1xrPhQKDK22hf6EynI7++Yx6QJaBZudk9gU8u6AodQL/H0yHvQKq+yojFvq/+5G01fZy
kY5qlZHp29Q1GbikCmjXi7O9Zq7PtJSRnKCfmgIQKcVk/kBxT3SIxAH2H0iM4Li6xxjUwMt5Ib7l
2L8ODOke8Tq4V9t/CAjkKFHOLu7MI5HxcxsgZRXjrXJ+ixPbh3yJU7Azs0IKBJAFH2+6pb+QalFP
fHVLeO+Zlz1edulWsIow45n4FZg0wPUHtzAwOdNrTMA8HABvVPBoEt8w4jcoaEWyGWMgtQ+XiDss
1thCPeVTKIfAKJBycU8KZzCD4VJMFzrGBY8sFY+QFuGI+LNXOqqRTby7pYcCbDKCHjsn4HOtzu4C
gBo0DIgbsKpmrfCfovFyzHxUVtNRBBVD6w5rEvB+936y3UFLOS7J0AZu6lBb/ys2rlZ1fYuNrc37
Y1i/rbO7xQrEeerBJAoRKnN15Bk6mIxSkb/zJxBRZnYXmf8FvzkjRVMSmyftGS4I/gModayUnTOa
sSCHJqziOGbEEWlkxuAMJ6HPtO1vRxKRTyNwTnMhigCvlaQNMIHJqgWG7Nb+9lXKSNEj8qJmcFXN
MsQc3a0zQRo69CJw0Ldm/rNutZrRl9WmNAagzqf28TQUhvQM68kRwpUcUCyPwqxJJuX8No5ilVJZ
HK2yl4un93cC6ZAn6xmJ+xGL/iZ0bAEeuxjDDfAt6mYaPpL5LgU5Bc5i4GY433pqlp5YCBRT1yFH
1TNJZ/t7rLnIRM1IqmwpJdZf5+HmjKgbwlHVOCfavV/1JyNL0VZ4GrgAyIgtjEmJ4v2ww7E0AeIN
3iNhPBlxTj/hcgp18vtQEJ/F/7q/uJbSz5gq6e4Y9cyUiVFs6HAgvHpcJStyLRnE/OYogbbDh8KW
4hAaacspGzRCRTJ42cevS2PDNpoKPg2x+K+ACvJsem/30yjbdATmQZVeXFaIZGiszSPNULvAOt7T
c/SOSfydOZ4oKyuCn50+asYbQ7Q6GFl6gUWJrr241BosBHZJqopuSgJhLSyZDKQUhiREJpYhKZ5G
qb8lOnRBzjVIlxBzmrw+a4/WJyYSk/QWLJDv1C+0SrW14ltsEEx3G6v8y1uXkGSUXifdA6f11cDS
KZw+oX26EVQXHn5aA+v3eIFMcFoSI9tkyXE64yc/282MK/Zsask+8XwpsH/rDzc7G0UthqIg31XY
4j82LV0RZkiGPzMilkIoL0lW4+9jNft0DV41/UPtqTJN7PNCh4kx/jg7qHcXHehfhdOm8DY23kxP
JL8tVyP3+ebUakZLmVrMLbkhY8ZWYrIhFqDFT5DqTPg629y6x71TM0ai7ay6hUH15TA43I8QAhx7
E6FMp6p0wot9xbWntYTlnIgFbv8z3uE7NCTkwKw18GJDsqkK+eD8iT6w3S06grlxFMR4cRUBorB6
XVzzzUPrL9X7bqze6CP6leie1iArQMSv3ZjKCNlCuQZOFP8b3jiW5aN86VPaBzRZYugA8aPixo02
KGOVAj+EHCmfrlmdZ/9tCsVhYvxjPs+hOjUPP4QXkqYD1hJUoNSTzJWzxoSKji9JIaSmXeEz6RTy
yeMd+ot3pnsvsmBM7IVJWMfsM3Dacjt+8AU9GgAsqR9a2W1y1ZWd9VLnCDlTr+c5AWnflJW7ewXZ
VIyvEi6kutzob6FNEyOKPbBu2YhZq8Y7KDV4Adj6Lc4oLz0FvU4XeWIq/ljAhG9GHL9m46GgSYjm
SeyoiUfmwoNoThmCny1ygvUAdcSfWlC76CgCFJBTQtrHSf4rmXvyH0TSJO3pwI1doNSX5fwP9i2D
+sPMSgKG+JOM53RPRlXwO/h0nGTpnvGL4UuCll7L3uceej3f7MScUdwWBIapNzF2la8Amm84KicN
vQLLuGmqYaAp8OjETaA8oN1KRnJDJl6F3s0fi5leOqeL7hNRsY0388Xrnte72716DzEVsAANVaA1
6qd63gkF+a1zjNovvbyROs+Owor+vzbOxIZobqEQ58h8qpjokACl0I6Bp4arCC8gLeQj19kAFGa4
lXUTQIBfRuh3OIOdY58MF2AiayRiEWK3NJU0Z7mGoBGpAMOmcaju1HmYOi99wPgHlubalSvAZ0Q+
qGEu/WNzFWICHFRYuZlRyYdXuC0gQeA4jzLNUvUpuxhFPK5c+e3XfKX3t/teVtvIzc/y7X9nlp6/
iiVM6k9sUM4lCvk7xYHMYZ6LwkXJtrvmIc2NcJA3TBdVP1xjlLIPuMdZT6akudPcM1Kw0ASZZ1NG
DqHgHm7XIJzbCbGT7ORuJz++j7LrgFV6Pn+/qIa2suCaTF6J+9U2rDHuzrsFPy2odjMOHmxdnyHq
bRsdyHlc4EXUG0WcXvdu2/85uMdbyeXaSFDZzVa2MzOCJNLDSdE0oJzwI/tJMRXkiJTeq1Hi7wi4
9pfM6XnVkETVwjMhYo11Ic2k+7jffFC5kax87mcgHwA529nx4UvmnclFpfI7Y4OmG8hQcDeneYRv
XlUZVyaDbNziIAWKvkXlLdfktUItKCct2k1vvAbPvVONzzqIBK1lowpGavJ2FdF8xRfhw25N2Pwz
biW8kFxOtRlkQylxISvWvPCrCL21v+WkW/3uRvuAnfDiIZEbjvWIgT1yxwMJvo0yKQue82h+0xnP
nF5IqG3ajvNBVdHA5iz79X+nY9h5Zld3NXZwE5qdJASZYOw74hclQ5AN5B8Ami3C0cMHjGeJUcNH
1ToyEpAxieHetwSPEdXRXBehgJ6LfXEAs0zmsTO1au2Pe81N1N/lI4lwEN7iNYNv14583OuQPdWB
r4TvzSokRXPDxMAkK3LfT1eOB+4wxyqVIhUM3e5TZc4GsKGSkLCUiWcR7RBFx7lTJjJLZsyMZzQu
fkfdK5YL62bmvzhU7C+hmCCZdn1QyrtdiK379uYLdqNFURM6r+CsH6OAU1Dw4Nk/o8KMz9uNh7RP
UtJGmOFtAe2wE1Fc+8+upy+aqSD67o60I3tnmaW6Tu9Sj5vKHIo+UbXwmJUb/11eT845hkO8Ppcb
f90kY+fza2tUvn2l5xLG4wcYuDOmtCfQR2gNnMxsO/DBTRdhumT470F/ZF75RuH7/Zn72zfIhOjX
MvK1XZoClIn/dDSK6U8c7ths7iksn3uZIizkh/0Q6GVzaS/14/8MqYqDeqRWbxbmaMbtBp+iyhQX
Nko0WgD5x08FSlqNzvVJEsxLpnYVsF5ncYul4HFgkKbRNcrurhZ7FtbHLVuMMs9jWTypIqvc3EoZ
ivwCXgtD7hc4UCzqgPClZgbyRt2vZF0m0EHsF/swXFKW71RuUYfhXP9+hcGxV/9KY14ScvWgPbXB
tC8NOsoErsNO7XNI3+qHOjcXd7KOmKBvgf2jxcGPYLD/p7YlhrOeuuBELFfjjlGLtPqK3f/UvhDJ
d4BTWCeDh21DA2WKd70dtUguYm/A9uvK2klfYO0eCnaxpORqWgKZ8D2Qlg7aJm6C4KIfJogLcNSF
qeLzY5L4uhoHfOKLzXDHfkSqNBuCEymYdtxQx8XPGdrNpEz65GCBSYCvsiJr7fbXMASqSM0ZHC+F
rLOGJ6kJHqgWkgl+vAHAzC1TOw5WucIsY4yA7NQW1MAdr2cir8TzNeovs2FFjo9DmD1oJMy4J4Su
OxUIJGb8mjdJxF3dt3Ia/j0Lwz11lvzCStcLIw2hJ94hQECpVJmkKtX9AGZOQRC83aP674/z3E7W
yaKFW47vkruFOBKVghoupworMek434g+QfkP8MoD4ctO5dyJk3e8Hed7S9lPq7+jqTzNsuwod8JQ
wHX0iFugAsQbXMInJcQOlF8VqRFtG9f++Tl7OrVJck98SNQiMQeV7qM3nTrjiTiBVaoRKusAHPGx
fQNo/4U6QTrFT85RJJ3sS2irxOy5q7NwcwWdqhG/ST4owCy61+5WZaWqkWq00qJ8oF3wUTU7Yn+X
SJjkXQUu+GdbgDGbCjodBOU8o3feKjoQz+w5oE2JzeuU8Jj+4V/0pRMA5Izo+6MFoO2KwVgfWGDE
zsIKZ1OIhdNj7SD3Zrk5y9mxu2L55Ric5MxtjHiuAdQpvImAUw0xsxevvbO+nWbXnnp+mIkTfjy3
SgI61XlyU/rgSXeAYetQIL5CaSKzK9J1VeWXBvkokMgxXZtrkiQ/t4ev79D6apnC1VpSTXtXoQWg
XjJUrLMtyk8KNO4hTuWk+VOaUTf04AZZjV0thEC7HyC1dBd1CDLHEe19Se++MzpHXDdikYR2xCBq
8ZG5cDbhPTSlNadB8smWdI/6ua38JmRSAf45himx/gsNKd4oR3IzC1yrDT7/P4byAg2SLgCLmLB1
6oiixSCZNZBIIHNiNM0rzieUnNWh2WtWQLssNhTo5mPFMVksPdryxbQpReMyf0BINOo+WEqsbqQ5
rO9Pxp+oFzeAbI4cK+FA0+/RnhB+qNG9873aF8FEdOkC7fitymyjqbiNG3jou+K6+hAl0xn/LDs0
/sZnunyQ/7E5suuER/1D5Z3Jx2/BbuiesV+3akj833/8Fkufh1dome5nBFdL8n/jbDdIITxMrXLl
amoY1UAuXtB/uf/OWjnYjIdX2RSouSDZ6TKhoUIHdjdw7Se7RI85XmfccR6Ax24foNNWLGw8a9sl
FABwqio1EiG+Uw7p/jcO76M4FwGrqIDevpAbHcJSOYw3I9hXgFP9AUgAbIoSRK9DatZSfSWd+WhB
KFIdatkUUA8EctfHPjnyPh6+DbpkHXnhIPUEG4N2Rgd29Qi6Qn/QUD1e6fJ98womoGfCVUuFfhcZ
waMS3evetqXcSVkogxhj+Zcg/n0OteLUmOQlgTFFSut3+bU6pa4z72EKjNavh9vLuFEdvLyJE/en
YV9zp2SI66nkhBAfrjjKdy9EGOjyDNcoSHIr4wS75LcBSCbgo35K90NcQmPYLmc7rWJgRP72eM/Q
dNtHZWTHyoQFVgaEq6eA/L/3FmDPX/QksxhKqAmqz4tP+GYU7mWTajaQw9NiGopP8tEzyX7hYEG8
vzPEnt3uM6fZ37FGimb9RonGuEp3lGRM9q3Wno5Nh8Z15IITWWQ+SYo8jCjfXb+kIUqEIuvbA3/Q
sbfJWgd2E865ZDInbNhQeKktM7os1Sbv2HyEEPfduMWu9ZhPVMXzHDPvhFKsVU50GzKUlx+ml/Qw
mScqQnB2yWC/IiztouEEZl8hUwNb+1t5lyn/jJ4wtEr5XHMI25186iISin+LeOCmsyU61lCobCQ4
xc+g7ktEy1EY6PfATqHWeT8vFJLDnGplmRbvsWQ2w1kfa1LbawYkDxCdOQVd8JbjqdOZ+OWxnYU2
biD83QQdq2WV2/Y8hoJQ9I3pw9zJRg2saqqlGaacUCwfZCXC7KSlWraJmF1sUkGXllKnx9mdPF4l
6MYWKLoJAfuKiacgscSNEeQf5v5VfVAVLeVJWPZs8fkvknqaYv6ApvDI0Zq2wYumVLUqpCfoopcL
3IMBUxo7BEpUrhln/qvraxMVUrJRJ3QCP5wTjyWtW4X0PtfV9tTf9ECB9aoPYijp0Exv+5p2++pE
QuFCX9JkYPJohE1dP+lVcoaVch6AgkIZcqRp/YP5tptmmVUTXdXoxUar1Bhq+Zh1/DlOSUP/T3sJ
CFx8+IBA0Yn7PjmLljUfNoafiYOa50Yh7PhKukgJ+i7jgJN2JtnFGHMFPCFWmdd6Mq6d+ZdkA9DZ
jgdHO1uMkhStjE8VYmZklN1PzHK9SljmVoPeMLNhokaPYl6HecyB7QKudJ6TMXM5CqOGRfzMGrco
Yior5l98pLyImYW2P13sK28WkZIZtj2kAT7VmuJZo+wAb3OkAg9alKPftZjlp7sS8ECbWn/DAfsq
jejR9dY7LW/WH4Vn0AQOas7l/OfHpZnwTQmXolKTbHx8vdxHlqfsEMuqB8UdsMJOx9W6wKOWFTTg
uuruyWQZ4TBWwUOiWjVsTI5msH90mgBJ9lNHRyXh/mDHNrS4QVhpwNlRALhLTvEotioYf8c173eb
vjfpnckSY20Ejb/CeJpSV4x0zZJVSGtGnWh+6/3jxTGaiAH2KbyAbVJ+eLjQtnKKGFPWiVBFRbtn
ZN64WDEDWtJZ2ZMzMMmWKgLP/IFfgoYM/yIMx0qU9B5+T3tfCz7pGLOpiIqHGcXS0mzCqU6O7cVE
QW/IWcltKeYxThUlk66J2KSX5Klq5wNIw2HBLq2+XMy/K7jPcWzkkX4HehyZXzCp0fsy/H+VqCba
b4PRGWmbKdiJPC4146AFVWedUZ6/NsDVfOIfp0wNQZHU6tRfB0MySNEck/72qsibgPscTydp8/Ye
fTpORGPmkS4jdjIgaYU7r/QKW9eCHPRpzOlR5saTNQ7dZ4vFZ+Bb0xHaewswpWPmFDVtZbNSn8VR
kMyNVI8VMNxD8y7daT4sE2arqex6xkmAFj09X3AywtwvrdXCjRsDY88dJ7WAfdrfMZDMkG0tbUjT
KrVgM5plbsKn73n37iHMcTwPPlWiGL8EnplSaJGg8eJYJpiwHsUDhNs4yuWy+4+8BuRni9gt5e1m
7bKFHbDp042DlLSdbfbW3CbzZRchDQoYkUe4j2tCSiUKG27pNTw7LEplPaCi6Jjlphvb4LDkvI3U
P27FjJzpn5EhZQyM5ZsvKLLzJb2Bw5A4sPFR9byCuebvA3WXUF047If8zwjIEboi5IBjIoHPvVuH
3LpmxOYey0oxwFyeeKgIOCEavMUvjxwuwhPKLOqz6WHf/adY5BXrjTZkd9mflDxnnz9zDuxuci6V
ANoFOF/u0c7GD0X9k0mciyhEOtMSxEWC9uOtxx0fThMg/KOvk9EATaObe1paM9+ZPcQnHCcrpkg+
TSiKqKrBUJRbXIgqUkB5/6sZ6Y6I/KNa8OI5OQFTemLqHN5NsqdbRujewJqilWU6gm12KC2NgJ1Q
lQ9iznV0PsEoD/q9Kcqa6eRd0hRGblfnesROItuXDbeHxDxU9iB1K04psSzNQBuFa3JGKrhq0thM
x2/uwMBOlBMofJc4DC3p+BioTkFEXaojPnziKGEPkZrm1haWLPhxb+yialKYOyid8JwvthY48KWv
IWVNrMGOJCdk8efDGjZc8ONVCEWdusAQr3eq3A2WBabO4tHTTV1xPataDJEbjf/gHwTTqxIJaR3a
RzpBsQKMUNOM3TwWKrPDMDstBfpYZYW+yDwVF7mDhdhJMTmWD/uLH/KlitHb50Ud8AhpH990Rpex
WGhPPU70gz3k7F/Jz5CftSctWDVwTVhTJDqU/yktIbfSh1bOaxU07FRLoeho+ST6ACPMeWbYPuxO
umicMKUFLWXlpiinMDBqrxy1Xa5uGK+AOORqzk1D2X+nJCQFMDoLijEUGU+mAbun9geWmNfIUVTY
Exeq7VG4Gzt2CiqVI82hrC9Fgj6r3L/CgSQx2cUo4aJunXWiRruHY89+rFbVjxh5qloBfTWHljwt
EYL/0pIZt3FSiYDbnJZX2raksjcBvotxTIODIm85iz6tSZBhcfrkA6Eqohm3bMdq4Cyj1y4Tjs5x
qAqORG/Hc8AlC8QxYkrle9/1OjVBuLMipJnNw7irJgxYQXkMbrpKRP4cP4VHEwOB/ECoMz3NdXdM
qNNPPYD7vm9WZobizA0ibKoJEdpgQI+UBN+KLuqgNtQvjoCb0VmdA9Jijos81HHZwVfy3D8b4amk
DGMGin+ePJFwc34PlpdB0i9J53DL7nSh3PjWAiCO9TFcZnRl7GZ/QQil3TOiNYpASMaok4PvFj84
Zmnz9WG+Qs4aglr8cPN57CFDm2aZRYO33RQsKf3+NWtxD1qkBCfTLm75VSfhPZMdkvCjHF3/dJKn
aIygwHaYai1lS+2/lRomKEsHFsWtvBNWGOGPvltZVwHhLhlUVhEGhobygtx8qhAbSZodk0YWRzFU
XlJMf+ZIJBRvrun0j86wOQAYxSC+eij2j2XW6BvtTR7+cnSk5fiUhQw5HzmbBc7FG1FhDaL0DlGu
td1dsrm4YVT4RAvg+TwUM0Tq9M72X5XgJebT4rYWSNVg+GJCpn+IQo07PRd+l9b/bR8Nt2TrX67x
zg/hMQXPGd/KyOAUNrfa8W9KiL0o2krCxkk2mxKYJzpIsqhQDfZRKM//5lgAkrMdOLVT/Bb7M6ZG
La8CPhDd79NeQGjJHQrAsjA/SWLxmhwhQqI2apY7B6LbMULapaSsPzuM4mhMwMk0LERnsbVrdK8V
cREk74OYeu3ZalnaboHGD8Dq/Qz6YVf9j63Ms9ozSq1aK/R0Lfv6M/BQ52PW8Kv5Jyj0Qn+T686D
G8mTyFBJmydERBEQc10Crp9ynvaE3D8EkD29C5hsKWgD8RTjdvMbfWoVNZAUrR94A3JMRHT0z1KB
+IR/H4cstNr23hv1orDrG6HmJbFT7elz859i8Yjg4pHTEelcy9KJ6Kb84mEMuxmT3zthW7EHtNIZ
Kp+32puq59Q/tB5NdDtQjNs51ikPFvrkRJC061HDeE9Rd/AuPrVlgCxmlu/MTiChSuCDGrjXUMMN
HsG1xG434xeeyk3yOTRQarBmazaD93bFTEleZ/hvdVw/Bfizybf3s64N0iUVmsKONh+qZ/dmUQoX
rsOseiUM0q6DKsnriW7IRPzHOV/xUvhm4Z41nA+ujCUC20/zt4kK+Go+oBlsEDbPE41fRJ8ezZLr
P9SW4RiA0+0tVl2pDh7YdWe/3BNy7NMUG9lOA3S3Z4p4qr7CNXC5BYUO2IUU2VlQx4OFpQjd+72F
UizteJKJGIf8F3AnP8E3XsR7S9IaQrqCTWWFySPY2MtMSFror+Tc/PVe2YNM5HtO2MGn/tX/8RmI
TCJfWp9KOuZZS3BtaR5VDin210imtqYXydayEo5ZDVG+2kIf7o4Ar+2nwc/qS4Fh1G115WjTMIF6
1AWJbpWeLNPeWqJb9Pj89tTZ2iB22IexS80t7/HlzpGJ4Bjdc0eY86KC2ol5+kZDL8dUIF69DkLf
iVJC0ZyE1X8eQBMPRyOsaUJ9Cv34xMCFoQYX1RuZLK2zWJUu998LCaW4A9Csv60JRBFxIXJyCwvw
pQf13//Hh5GlSVofsa+vjbDrurwF5LiDGk/cYb0f1Va6YbDECgOuXfv+lIEns1726DdM/ednMbWx
8lcQ56LkaCne2g9CTOwrCXDyqrGlG496/TGolY51auM9v5xb+6oy0Yc5HFkfKx408GOksXpZqjDN
T5QcV1h08gAb0YnmNGZMbaqaQI2dnMPeijSx90oQNEEcMgQNM6DwgN13QKhXnWzQMZ0d9dAPx7C+
avlQalK4HGgvTiysq9g02RQ+jF+HOee0eIenB8Z5xPFQXgqg2mSW1h4FDBODEu2/qBlBt5S/4SGk
gNDTGDL5m0wAijBqK9A9OgN8cZIA3tvOJ4HxDrqa9ljekRc025To6YyzdLJ13i4w16WS+MMUst5i
gOXkU8QKsf81zpT0Td2+NDbSCkikvZtyY3NBIGEl3aL9g2cawQDzQjVepql87VIjCx+5LFSBGwLg
PJl88747x6t4+S5O/hKcdpIqP7jx+FbO81NTdgTI3KAuhIksmM3nyEDK+zliMkEGt8ap2WQmopo3
CCzSAq9I7MbhBqHUYHRt+TsYRlDMRBIrFBTD+VCY0WD37CWXADvavHXnxE3+7+yK5hkRPQfqm4OP
0ciqhrg7J9YC7oqrkuXb4WrV60JVBFEOaTnQSJ24AP9dsb5Q33wp/GylBSNe0x6t6ADVtUDOu6Z6
F1icBz4RA21vFMm0orzbuoUH9szILHfUzb6ymKj16exQXJXa1byNdd+W8SoNHxFWZ1X/OaIG9Zdu
VeRDbXOWMd6GWHQRNJmA2En+cMaS2mv8hD4jXG/oVsNCX4LMKNLByp8XlXCj01WD1lsMa7ntX6c+
jwdmolm/JVpmQQsHLkmGh3uUHnrfjK2ZITnEGvWkyV06/VcQhzUY6GlgeuCg+WPKCQwCSArX3xRk
+Rhh8n5YCxlMjNIRHPVdfJh9LP0ffSa5rITWgnBLojEopZf6R271x9/YpqaIDEG9wyIHej9yo8w+
rvpnDUl9LCoB+qoeYT5+1dQAU17OAc4RnAMDVp3ZpPvExw5JHNC4i0q7azldSeF9GksQ7V314BFV
pkG52Md0WWsHqSGOKgb9PcdvO7Cck4+SLeYfPjKR+WWkwDXJ22T3N8MpTbQaffaKw0gy3wna1pXa
9uRWTHRWnnJkZ4lfTpdxuYutsXxnl4YTeI0Xk3BaO0zuS27sLmxfcT7E7ZJGBkrrkvAhdwC3NraA
gNlgqNoaXBP7rLSslkdP4YK3Dn2pm6VhwhjiQ0szIgoZQHRSpr8ZarzPEVgAkw+qN/GezSRxwtGa
rGHDHka3DbUpQ4BBIM0XVLUc3cbYctGgv8tTDV5CVwKnKjSzrtN8n+qhGXC+iyIMlckHgQyHhMfq
1HtcNPywDEaCRoILH+112I4edqEmHu0Mr74hqFIhorOkwo45CbewNmEOcMLmmcwE6tY+60HJ8YTL
5OPKbHiXUmrGamSxxShWXw/6PHOK1TvHXFtO6MbraniyeDkcChwQC8Ve/cQAHjT5mAJvPxePGhlh
zGfkrdwFC2wIq3I3NjdspEj9qBfrtM+tZx5uUh0NSL7PfPXObLOe8jCH/MRz3ZUhF7a1tvIoHxMy
V3PLjDP/oU/HW0bXtRjOjXyR5wgg4mTW9B1Hj/QJMiDeqKTYK8QT+vybEdwlxa1j6G+uy8HibJAu
Bxt0crTQVvrrD0cC/bhYsJqWFH1mI45pfNTy9jcel32QT9d9bUHwH5oxrE5GXTCKpckXVvugIWnh
BNvcPIxKvhZ315J4kg9opdCEIcLKcWasM1zG3hKaCWFbLfJA172wYti5QjRcb2exIputXeFPpbHU
bHoWffj8LLCJNnAvMlQ5XoVfWfFiglV46WVcTdDEb6cV6M6Ix4nuG7k8qBApwWZqpyGJlJZSynfa
quJpQlYcrbwXaHYNGRsJVZPjebY6mMA+RMj4lTmKnE0LsC52/BHmbFhMVBAkww0jaEjl1o0HFrr3
3yNjo5cV7u+a7nrATY/CiS12jumdZtrYDzlKYVUZb4vBLDogb3FE8Qg6jf88cTP7l5wqwvH410uT
zT1Qz1sP0kQaBsHzEKuJnP93iX/vLdjc+YHP6s2yWwnzITYt3vr4WHETtHKeyIItxljSYaKtzOmy
auOlOGYVpOU8SACP9bXvvChTxbBBc49oYW/xt+acgFPOU/2U4VD5yn0asxj7lRq16wCpjU8CDpS1
lo56sAB4G2kKBwLX0qVFlI2ewJcoQDAL3Edh7IzR16L9rkrYjvIAYQEH7x5aW+7lePbCtwCJZq1k
Pjggo6pPt3PfgXGMdMt/CLOwGfAaGXeQXDydWhe4tf/sH8SmR9zLOvfD36+VC9ONcMqMvDZosO7C
A6AXU1H8GyeuzL+6aSwwFOA5he5r2OiFA1z/oyBxHbc2b049ueIiMityjpDPjzK79YJJzDgqp//9
G40uRtWzY5Fac+/zBwuATYo8KV1BDApgSvRvxlusc9RmWiKJ0Kx31BkmhCoEmF33bvxMeScaYTv6
0+gZzOOdOkWhVogzuy3UEAVSj9b+9QqQcYOerC0uMtAUbAM0QKlvYz18NMZ3IVP45xIPSdAdGDz+
BdYoewpnDq20//lWB+ysuWwi+ZzZYHN+DEHmFDekAVYC+dGqQRYOylWzqM5u1JFhiGiGAWzpORM+
9PYXgFEN/rvj1QF8LvDrrM+l0JcytmMbA4bMRZwo1QFl6o8EURkDPHZ2a1SyI45O++I7b38A93jk
W/XO8xvzrqND5P8EomoIZ3waA/jqjoq6zwpP1IZBeW0nS+XC87bfongfb5k/R4dNlcPKuxD4auq8
79ns0CHIYFrppK0/GRdiGJvjKK6KQiB+tN30o7kCBDRvehU1FWX8H+hoUsbSBUL74lMSRE58oFS0
zc35iAyeDJYXUFuxSTNIbGrr/jMAicBba4DLdWYuYtF6ExIs6drVtLTAr21kMwyfPa7Wo657GWhI
OUrBYrco/enFCSz8jyT3RnXeVWqFmmT+tQ6eBTC53f6F+uehZlleW/DPPN6ton/2nOQvXT/w15sY
2R3BcRM4iAGWk27XJmL1xFLsjD4f/GFNMxU1VqGYdnyBpHL76hY0mvtU24Gvbp2G1rtzUMUbjhBm
5hUr3+ZrVmipb5HvYTM5aDw/L8Ydjg+BCfpJzESIDFWCu+nXy+ZLC+hV0hGB2PS7bNq+zqHhmnKQ
QmKiFS/u5YnNJ19NihMZfjjk5odurXOpm7WEUqsUymMspHOOJUnu0W/9rpKCxpxix7Wn7NvulgwV
VtzWiiZ/THWrPaVKI2rsqtUhDbhxRjKexaRkLJZiRzNgX2Auv0cNZEuUwQgl5wX17esg/Ew6dwXi
c9qUraX4KZttvz8UnaGJZwvwq7PvdCowENh4elXXriPwhvRwaKJnnS9FprYoXFFAfIR9Xw92bJjW
hsOGWBd3uDUzIPR/iFqygvbCjtgIK13BXB6qSmNPLhmS24C4OCQs6XyNEjUIkkx84j5ie6PDJlte
kNaot1W9XiZtxQyz7DEmwPwX5KKGhqeOcaRs3jgNuGop0Lz0vBcu66BpRIzSUHzKAAMV4wcKam7n
N/O/gLbL0MM2WnCC0dFvSuIYCqHG3YG8myWfcZ4fy2FMuvshXnEq4mk/nqtmLiI+COxykojZz0/K
DdDDYcsKEk1sTP3IgoYUQgucEq4geEsvVp1Q2yXYw1dJDl/wmpI4CQHEvforLJonVEZZwlA/sU06
PblMqP42OFnj6kk1NAUVZpOSc061nijWLSXfPUnHCFiaL3MPOQsLKMAVtJVLSoMH8ySRthWXO3Wa
/2ErP1djEu9SKFx3dg56UFj3sm36ZimScrsadwmXXFVhCmvAFSA0X25HcWytx4Y8Jvvsc0kJOTAA
EUU7SINSvNtk9KDidHqJPi8EeKxNAv1dX63Bu2oZjaNhGpdSaQsaHlG4Nd+eHVZIzcgcw2pQApk0
79Cn5ZlPsybm7PoziQco0cQ+68OpKmIuFOuTjq76FRpJJH1exko7ogaLM9mLvmesPboP9jyhdIko
LVImJOU6YwYaUhnNVd/G4HnBXiL7L5myqwjRFG7XpSoYOuME/y8qIrlBhNYUMwH3fyRZ2lAKUHlg
imQQr0kPSflyZcu42heH2fxJkxiS68xSQBM/pLvcGPwcTaloj1YFKUpwIfL+b9VgFK83vxtd/XW9
ARrjlTTYFa3Kjn+P7aAGp6XCiCi4/tH5ChhyoW+OVoz7fPxpShOA5hoEB4YQf03XivgibAXE0jWb
kRd33zCiufGBCoQ5+gYDYECacx48Su6i/ljPRKfzJ8aWky7w/iHn1UyZnaC7I5iczwd5+Gis2g39
jIrX32ImvPYPH8N1xpMMHXkwcVqzrG9bsAsrnC57IMChTO5XeooceLN1/a6J7v1H0Vgzxto7iBhd
yr32jbZiHTDbc+F5Tm4qByVtIJtXiKG566p+CvWrE38Vm0CzXuMSyWXem8WExBgVGa4OiHdwLIlz
B+TcuJkv+t56ToemqTORRUyQtVC+J9mcESl4ZIeu0JYECjOcMmlR8Ga5fkTqg+AgDiKeaVCLhtkR
byBl9aNqtl2TtoERpA9kz712dmUK2gPhD3RIQIX4xQ27vwJ6eLi7YRqZyrPSyvTp3l9YiIpq0kO9
BqhfviVjyBJaRSgK3UQa6zuMj0G4EaWyok9PX/P+ryoydvYTSOUQsdX3/Ien0yNTrBsgjs+MnqWV
EMy2nUxZ5MT64MXgaXn9X5uKgfBFC1M9UJDRSXCOgcnLv5xhcOUFUO64JeynMXu0jIXH30kS7M+W
0RMd59Rw0wINPtjfZKZYiRCTw/sqR3LbTmFOZ4h61ERVRFlPIj5RZ684+7MUN18R+BPeBecVzeV3
9YQ7mOehHnQ8Xkd0elPtt4YAYc7QzuYg6+K1IGk1h2uY7pokedfzbVihyDW2CClc10O7qo6ASnw3
dtSKBFRvMVp5nVJIYLnqRiovEXzPB2YCOsUVCnakSKXPENp+qHqCiZuup9ytB7WqNuHbGs1dHffT
UqlmSir3JCfwlhgmXGI4RD9kSi+SnJAw/dCjwT3Ghlw3bxF0xRkMyL/iiwyFlJJ/lojB1XAYOYQb
OkSwfd6wTqQsa+8qE0o8CF/nmmajHRjP7OreMMY4x1EY97g0LFkhQWRV976y0BDaWFqrCBsuq4a8
TheFOX5m8kaKq0J5FhLNz7YWk8Be7HJmuXVsk4ISftkW7z/z3FeWkRTSISG5nDLQrNjmN2+xeWyK
zIkcTdDVdjCI9xpRXQNRXAHYUKDbpL+q3VmJSSEvzDT0yhZ3wexdeekxZ7FzEqsdTWxkKSeTQSl+
B/d7i+/Pf6y1wNp3rsWAumVDmuHqJljHaOlm7htjgMUIN8x+1DCtd3PbFvMzCHanfm3o+uNtUS/K
FIC0DR5GzuDV7pGta6DpEa8Yw5SWbqutP1bOX58QfYgnc4xT9gpd8Lbzx/YGGaIZkk7ZRG+sbY1Q
mBWm7JoEhd1HFIs6+it59SLhGkLrEa5xFomKemO3m/J0JdcAk8SVrWpHucb5NFsauThdbdaezwmU
aaz4jUUXEVJw/LnimKM7tKJYNWwf+Ttghh5r1vqKwmzehFjEmUm7VxEnb6PTVpBwHndDzat0B2iO
nCRxa5OhbaBKNsDmoGl6NX563DsBJ6SV2t7hF1z4k0oRkT+XocMzNYw8vKI6NIKbpfqnBwSTtvMz
RtU/3FGIZTSj1YL8k/MPl393RThjacvxQWpSGZJk0s9T3m+lsub751uCgvSv+IthDZNzl6fynCdU
SIrPyhHG7R5Bte7CHm4OS3grZdGdhSHL4l9TuJ8j4r7mjt43ZniMHanDUH9XEqnv0rpL4bX7xt+x
bejTqzV0Oe8GyB47z6D7jpSPK4LHX2LirhtRA9a7NAKtLHExBhX9QEEhUDYw42pTDXr/uE+iaeV7
uzl3bvDZgCbNyiDufnzhVnQy+lMa9OGEOCL8tj/0/B2iL6aivvx9b58QbzuiVF9ezx2PHQQA5vfq
m4U8f1wKe6DK92m2EIYRCyVl6D5+ZHpIO8G0j2rt6CctSXrMM8h7+1XetcqQAevHWOx7wIMQEP/d
WQMQlZ8otIpK8euMRvHT4D2pwePRxWkRhP69kLFSo4sJKEiU1FMKNy3kger7NafgFNDHj+BPbb0U
ZFHtIpFj1Wnx85o+SMAn6LNFnfZhKwUTunabHLLBP4Ae2sQkmt6oqpuFzEEJX4Vt+RvA2rnEzojJ
1iVNB06EQJgLt4rYM5i6JRM6NgkU2GtYePr+GtuwV765ZIDEqEX4YhqS7d3rmT814t1ogSc7wNsr
INH8wUERpzWUTGObt0ZotBPuDmfpJLYYuqs0ZAKdFrqfdX8Fl7nd5wH7J9JclETB6Adgy6zxtp+x
jHD4+cMtfzDrqmDK7l0B/4jaT73ZakGxUHMYafWoyFEz99XfgMQUP9Ml4+ZOTo2AFJEPCBkFK2wJ
d4d6nCt9e4jclUi7MGXUEkvxxyKFCLVBain6jxgq8qRVKyyXipQr8BgWFw/sBmGxsVKe7w9aNugq
4u/XUBadg+Zw6RNa+J5KDcAibiC+C5kYlDSCoJJwXc3yVvQ179HzT0ZdjxtMefRqeghoS/ErvVoE
scKwWJCA/XtnZiVWKYvswG8JLMldmYuNx1edV4yBMG17dCGyFY2a56SbVoi1IjRrmMxWKpGPAJi3
mOlk1KWQpGHzzsDTRgPD4dN7WJyKTxgyyPtrCJu6dxxEMj8hexdjxlM1rTEnTAgiuwHUs5xoE1uk
a4rUOxDTe1hJG+DhahitW708fqTBq6rBowRd2p4IsBXxV844S550T+aGYfshzpFGC+UxdV/QVfFV
NxUYvvcj324EdMlKJgPl0PkAuqA0BxVNzrMU2VsQ/JkApbUr1CgwZMBVIbODk5+CeB+veyG7KwlK
BGutnbM6NQKx8U2wScSUPdBJSaNPFtMVCPumm9KIc0/lcbXdmkOy/7Jpr0X7fBxS1n+OCKmCdV/b
hDRpWArvjzlyDuLQKzbu2eSvGSDpJNG7bkRZiiZFc+wkpha9a/sbkX3kZXxdzN2Eo54AbkncAfEO
FIn6070m3Edr2ZAlVPOmm0ZWr7iNs8YzwSMgsdIkZLHCOKaJ4sFjD9p1YvhwQgfdpU6642voiX55
DI/viMADihEEGIb/yzp4qW95zA2M3t/LFRkROxG7w+y2jUG8XiaEx2878sbJu21NMs1q74J7Vj4Z
ldCawxH1OComatFUFCpXLKmrJUNjaJazh9W+XrI0QdfunWCQBRlAhidksfOEUSewXe9WPS7Bhold
H5jMny+VT6pkjv+t5k5BTtde3CAaAo2wh06dTzAUyvEVc9cUUqwThJ0f5lyknan95K2yuKAYMAbu
WrFxS9w0wnRCoYUKVjBu3Vm/k7dFfS4Bbw1sSd33jfeH380L3vel2GnltxvZ+AY+bph1XyFmVEP2
V5raeDgqYwbaCoeB4wt3d1ZsGOpoVgRde0Cq3Cg1eKq46rNrNH+EcAgl88tPdvt9JtxvBdaACbbl
k8YuuGYroIRhPe/pL0asu5yJkU1bhFa33Rig1I1MXHxcbhdGH3kraTyUkrciUgUbrvGU+9cgs686
8FxFkUmGLFH+poBJfQSfuN9nl5kjv2PpSevQECeJaKNoRvDcM/xLXj9emJC12yWZh3pBYxUBJJKR
dd2+Zb5pG5Pa6EXMRSO2dyCC7t92BVL/Z08RaZg669ZIG/j3fj1KJVwh6zL+pcksxKxCkTibaucj
TC0NN8aY8ekZJMjBOBO12+LqOZWnAmKU39tZfigMEIBXavlpVu8f5wU7taXjtqpWyqqJeE486JVv
t8trP6j/BYRlxUNYm2LddF/OhlZ6QjwRXvfOjY8NmaY3Pjzl6+nrmHbCHgJcVXe8Weh1HF2L4ipM
GGGkluvqTxeHowg42ZEbHisITQVwj2NrucnTT0aJlQC3nsK+OJR1JxjojCGE9iCcpMEUk9zE9hML
Fm+Pww4SSmRzjQ9hxG0pHC8UjGMNsqMLXFrPenGctLlBvi0cMBC7cOoRVYvEXvWcF/GUUuCA5piO
/gwx+J2tc0YXnF4ovZj+JScgEN/e19ls6g8EjrxErYx3Ep0ssU/psDprR8pamFN3AITrTwNHtrfM
DvCvbbfr52Y0fsYBa6gUhVjlhjdiLoOdrnmmgpWDw/iKlgTiriXgeQVws5p33Ri3jV6MihmAsY+r
zrt7eXCjvB7mhgCxdPqOA/qsQnvbxcQFZTCTly95xwLfEmk7mO2y5HLE23cWNWfYfs8TB67kxJWt
lP/ZWSEUjQgdEpnOnd16eOp55ktR/TNv4nBz4Ovl9Adauf1MabfZ/rDWyTL3r+vxg/MZXxsI0mDC
7HogIXED6BwUA70etcJZiNIDBEoXEejxr39gyGq4KDpZvONJKmIFpP3wjjJTKBu96XvPNndWcb7c
tWXBQGzSQvBVuCjb3GhGiY2hWWZeBLAE6VBgU01VOFNv4FB/57XqqvXOFOechANASQZNN8fZ3Kad
glSp/fHKJIHPRdOxLA1/GzlEh3BVCfiDDRhaNX5qsFv8W7T5ZJJx4FJUtDIbPFQgbKMnnTdWUhMR
Cg+COE1AGRtFuyE2tn9MBMLvWl7f+/Y9QA4Zx5sKbHOIkkV77e5cyLj1hS+2WXOKNaIK1cD7CJE6
ZAGidQZIkWvC14nT0L3EbbCLDE5dYqBaxYRI+oh4OsVZT7LX2yTUkKwm1OLtfdMYOI6IOb3vadBH
dOOBajB/s97oMTP0OrTESsEosnpKGoFV7mV2slwWC3z48HJC9coZjlRgUjPiw6xuMEm9yFGFHAHH
VLgQmNclN5O7ybv48MQ/ZU90IC/mDUT4IeJnedLz9HJrHjQRMVqXY9gNZRPRxkTLM4WEqmKia+2I
2FVfxMj5y31HqATVSyXUW2y44NC06+8fgBAMwNULCuXy/1c2q6UnUqt/uaQ1fCExBmvUWLE15NEc
g7JIYH8CVKWQNmIJVuvCmjd8lGyEz5X/hziN2l375r9B8iMITvk8Q/ba7rXCTCRPnZk7ChqaR6ea
oxQJPrRsMIE7UZVntya5by4TyTpIEjOIKOqztOjKoHSe59ygWBFLqPDNS+V2y5EmVyo5kqSV73zj
1yYPqndpVpErmizJZDWZ+C1MVKglBjbhx+tFrwDU3Zdbr6jv5aCj2DU0BQzcd0hjus3NY3jcKLDh
DqWtWKg4fNaIGrAXsUWcQT+VP3g66rUTuLwazbYPk7N2lptUdMq73vlGwTaI8o9r2YV6MgZcwVT0
pVNZ0BTCXwKOxa1wsvAtBkDSNZ4u3VGVLq+U4Pfq6XSscnIQFeHRj7z0+arb4DpCSS2tJWoDVog6
OURldzN/jjZGp3NNpjSbdC8hhhut9MbfloJf6mRd6UQ2HzP+4h3adqRm9yQCyL44+XJG0gCoISQE
Ins4B1VAgI73XcNxfoDJtTDhlQsnTKHTOGHa/Cm/K2zL9x3zIWbc9HUjuTVVB0RdP6S3s5OaE1MW
JzB+V5Lx/982UoK/y98NOTi5WKJeVHGiJwRspYkmTl826HxM0A+oA78a00wR+OReII5col16s1UC
wbm+jqWmdwP9EzagK53JineNOVoqOitgPY2/uUaMx2MJWMdp3rXY+Ro2okV8OQFfA5NpapJIrLMJ
DiO9HTtBhkerM3Z9Lksh5GOigN21MtZQTim5l7Z0WQ8hI/ELAbuhq6wAi/6uxD6h7p31CSMEHwNA
VRhqXzCn8BpR2fdnI44Y3IYrPnkYuin0j8eXnbsLm7EdAlLrLpWvYXYL9nJbLcCeWJIzbGoiwtWn
XDYxluUctlHII08v5h5Zd/BA5OPuu1bLIaSjcXXEYrIOULyVzu90kQHVvyd2aH/s0VuRbz6gGGGX
7JRSFOK+CjNkhbCOXCgWJs5NPPuiQOScpEyBaEvrEAv2dYI5bjs2h7DXySmkllMheVVi4QAcD3Lb
T4Wx++Yx4QlVXS9qzcDrGDTu6UnodGSA/mi9k0tMINCgcFtuBdHzDY7O/LrnH85N0C934GgCZ9iV
EOEiwr67O+7OgJ5DJOxVZKFGdYf6cxA+iobvCjzvSLTcTqB+M7AwwWqmKsJzdOeZnMCUHSbBtbjx
lhALo0QirBwuU5uhIcOre3h8/Y2hRrUITaxbEz2wIhVdrr0Vgc4m2feUXpM6fKjQGKFL2/EOBqRZ
8LqlgcwPLWFo9Jax7oV/wfVc3KpSHIXy24yJT/6Nfp8DqpC86+uroED+oqMpjx+CKqhMgFNc6ghr
PCDHtoWpoXd/S95yRABH6vvnHNQZ3H7lLHWhSZFDn6MMHkXcnpjlgIHa4xgWjioo5hSni/HT1SJc
W7pH0Ir5F6TceOZzX4jvU8EHkxdjue4FnJZN8FfoT6ONbjSr7d5knVf5X/au/HOY46BtM9uvXMOU
5ULV4o5qlJop67MOzcp81ZTyvl+SgSo02a3SOFaZdkNSwB1bl5WP/NGO+KPn/kWpuMNMn4jz+XRd
FIJ4SSE8Opo71w5ZHc5lMaoEjWGnT9QMrUrt7buphIr5NoD/RrZeIEbqTUK54cnzNPy0hZto7y7h
ld7NivKqmOjjNkYmLvFL16Gu+F/zFXvFWT0wMoItQHH/77PNnXxjOjP5VcSm1haULmjFUtTTRz0B
I8dsRYkezjKYKc5YJDRy8ArLEzewA3D70VIl+8q+OkFiZxA4uA3Iq7UuJrqh3F4SpjGEnVFiF7C4
M+5ES8S33mKsf0jDziSQi/FDdUhrKoFzQRNl9du0D97T/OpNZ+3nNjA9tleg+YM/8JMas7hfLUmr
sO78kqp4KR+m460p4sH+3thfMUJHG2So1xaKK4qNDcpcedPUYQ2LSzIVADjX4QyMTRyTC71WkjN2
aXVPiFtbKaPb0nD4RQtNFVfGyKqhXuxH3kYjIZ5gDMpM2Gegxs7lFGPZif/YYgK8sKWXdrj1fyj4
j0UcA1h16uBkL+4tEtbtrrinRWJ5gfh3A+S0ZpnWCQV5M4+3JNCrJMdsOADh6PbXlUpERZtE7/BP
DI7zeJj9XZ8aeTAwwiAXS1+68nSMPtiQkQtmRELlfmtZQ3TNF6nPtR0RMGZVzbbBdKogHm2Llbdx
dEfhSKl1HoO97hPF+pxR731IthWQeRqYsQVrnN8w1lYwtlayg1mSwevOMgCokhJ2s1Mt9LTPWkBw
40tMtOBdOh7IwVYDmYh30Ke++5Lw2gNVjqTLtUuA3VLURYlR69fv5V7O6vAr0f4nzRQIh5cOYqyc
7JvtUylQteaSYIZboHhUw/LgQ8Sh3UoRHvIWiN5AvWBLbwehDTky9MCv+CTE+j/urhFRy6/7yiuu
Hz9j1JhM9LzFi9rU9E5wZO4k78Ld27o8Zofcxzpwl1x65fOAuck5o7Rua445ztuodtTwL27Q2+Rn
dyU95vqZUMMwUEpWZOdAN+eF6IlmOXjyRNTFmnoRBQsKv24BKR99w9fi3WIuStspOIvOgPqm+jqB
Wvmz9yLtjPjw+0pyfkihAw22F+M6E5xZchRyH6EjOil8J2Xz+95gPrTSB3I+U/T0tVkEYIU0gLzG
lIlmZRkFaikklrvM93MJlf6f+tk7s2E2zN1T9I5CQWM7UIYKFm4d9aWJzgpll44T7lQwG2Eh4Yl6
FgpgTYCKVDiyzvzOGzTSrb1TKuLkQfTJGLTl4J/nr99Vex2XayVDUPtbnJcYILpL1B/j6AVXXH+V
N6PIUNDCLRstDYWbI3DeCHgQDukqestZrTa2dxFHCeN5+Xp7BZHwmU7SOdjpPto6d6RgVt7/1UdT
ITQn3aEbdVPAlg6TAVAuN3ecKBsoyg+gMVPK3253dfUQv+z1juYgw3CH3OYrYqWorwv7OAM7prls
xAq05XpN/lSrIF9MaNugvbVFsD8FN+4dmA7An9ocjGPtsCAQMvugWIINTdVnhCop+vGo10Sx521g
56OJvGqTm9kK5gYPJwUt8+SiLZykbVvk27nXPg/O9PDWXxSRiJxvE4Xi+4i05SiIdyNDu5CkHRXJ
+Usc4HWIL1ycdeWVaY6zVQ/zyBM8K5Zi9v/cMpfr1V42jznSQFNfpK2hwtWSpv2Ae0UFyYpYtooa
NlfF0R7+3Pw+8DtXqzKrc6YVtwgKRLBtbQ4FVPRhA09JGUa63xldT8KJyuLlkGnU07nue0fsX0vB
qKiN8XzmHOOV/YcRGRLMC++8Wo85Sw+af7/BGXGfkB7so91Oh1ijFmzjvK31Io91MMPgie4SMfhO
tMdw3bD+dYlvqSi99aIGPOIhUAX6qZ7aAP8+MXr584iBZFnquHNB6HV0+SKbhhjFGFbZfnbl93Md
tiPbUm6TGaLPSeFgBqKw6DnIwVdWaeDJcJwmR354Rt3Jfhix3iu1mJ6Xh617oHpgPg4YoyK+VAyx
HTUQNOQ5tD0RjgTJgEaGQlzvHFD8mAKRxGUTc07lrrCvoPZ7ksRCJEeQpUYdGymAbqOyDLyDV1rd
cwd/nyX5iqEDTOFC67Vqr+aGShP3BD5ZW5ZcQ3GT9ihrKhgPyjObb7RlNKKhKWo/YqokYzNEdaVq
DGCvxeCRq6k/BLgs0kjLQchE/IthPFbBEwiDq3bhIiiWiFXD6AAoGPlSuGLQMM4jjOti6EVWJNm7
zASOo+IbWIEowyzkfE1YtTAUkrjDCmG4A54NB6FJz4VLQxyrzd6EtHolKVC+mEgJUUCBnAvbLRLL
bDVl+IQcqert9RTxHBG+mOrBvoLrB41E/yrx+J+EVM3mD0JsnD8D8muX08BZmcQrf0TbhIgabEBc
TJv55HwmMGBrIcGpeD2H7DvZ2sljS7+AciJFdDmeH1eDZrj70+4uwFuIWL9feZVmuT86bFYJ86HE
+KSV+eICpFVhrqVUPDrH4/0V9S6CNYR5a7MOVDPf6d0h2wo5nHoh51gu0YDM0spHKSgXJZBPKU56
3iASCDp/G8ZE9zsormg+n4KxnmOIY5Gn3QAs1l4DI456gHarxSgZGcX0GB6bot/CdiUh3F+XTreH
IId1wJ+HxSAYTb8dawlq5mOWSTiAhi1y9HpArKpBZtZl6wVsFrL+WQRaS5iGJUgi6EkuTqGxXqqj
NhWU6Kv3iSK00phEMxhGdtgLlhOumCTLazQkieQt/LXnSLAy43A3sdz9A8b+DowYIlhdAdE5jy5k
GS8Ni8jtqZV74NfrjQFzfVB9s+8qz1N2LtJebw9zVcG5CFugSZlyV+MM92yPteZc7hz2Q2Scefu6
GMl2Fewlh5N3mLUpRfW8woIZPTT21yl5wvaupFVJ3qiJPLtMHB54MqjqopaadJLEQPs2HLr91Htu
VmFIvtHQ0GyQ+0TThQVc3RbiuaMxxDJtHzaPveZ0w4L1z+QhBju9S4C4VxG29RRrQKr4PCfJJfi6
etVxhG1VPiYc8qFb/Mqw7PF1MAU+a9lGpiyxOngog2rxM1UYzJuN7sENas5Cro8hiG/5Tz0MXKzD
NIr5XHCEitda+tU60+KSng9p1aldWNDBTR58PdM2SNp8lGUx2BxNJbuCHDWnBNbhEbDMb+wT1DKy
8B7+cv9MmU6AXkY/mxO6Jb9zdjPMYQDEbaG2MxEQiw0EXDVecdwvajIjkj/zAa4erPNLqfArEij6
THUMRJFzLL2HgJlm8YwJS8QeMtm/nzK9DK5OgdnbfGRP9KNZpSliCzR9Y2khVuuTePEfhGvjOGLK
yk+l0wXinhbuGs00s35jt/vugS1Vqp6aPdGiGJg4fNNbEw2Cp+Y55uIjLog7T16lZXqn5JBtMpwD
z2r0VnaAMPL2si+1q9VJm6z3ZTLlwzOvoDgMe26c67LxBGwvqW+tDLk4zDP1Pn+KB2XrBTZvyFnE
r8oWn6HwAR3Vdme9M8rbyv9UhjBmDUdPEw5zFE4fEY5TaZiM+y6E237xvgxPPfn8wJ9QfaxIY8ue
tppPCbL58HRn35GpZJyZZgt8DUMsj2D2HglOz2ovRVLs494o+slLf4yqGelIKRc6X4zXMsHeNnb1
6DzMFHnr3N6MZLn/oUM3miM8TZ2pdlwlhw8n2jbr9WLg2DxdrH4HXw7mCR59QyuhVerPZWs3NrYS
IgfDu7QrLqMYY4okeojaUDD3MXRpY2bkxVZiLSoz7XKLtprikU52IfQA9uajZTj7SMsHGgT78VSX
GUu9b+Ttl+m7gFqF+Hj5gzLusdesjJO4fCe/gC0PMNdRAorb5iWy83vcJcyKEdh6UvEHSg2IWT7U
WO+p9+4q9FnbaEAPA9vIvkn1SC7AblYw1jiiAzuuIVjDaegVXt8B5hNRB4wTzjdqnamMTH02KMJP
rKPLu/qpMg5iHaJ5hbT3g2DaII0SbQCInE+Cvtsg4Mr/5P6n+2rIdw3MR+OXeB8clFYaX2P2heXC
oLEQwxOGDS3eo/O9ySsog590OoLA08nv6Q8H/9Ex6TeEcreF7/Hicjm2JjHpgNb1rBhLGUw16n3k
dVUwO5zKL2vJlt6CoxxsCI2+pMyb/nohgtsadYsYAsC3dZggdNtiCgn0i7Mhx5n6VIZex89CqKqf
/JedBLHWniP4H1EAWIzHe+IpSmGqYB6wW6+DwL/qBNPiiaTEAEMD+NeOvSIVI+dOJvwRUaj6NaVk
9j4+i+lvQdjr7clfy6siYYhrbVYYOUWtvt7opBm0tvFdRxsZWHExJiGlFmaUfh+k5YbkumxTrAUB
u1JIFxs4GNDrk8+nxoyHB26uwSS/3yf077Z7CPimtKQ2Dcqomu/BoZ7W0uByoXV04HeO9Fo73StV
XELTCeEvis1wDmOSgmcvPTy+RhEmP9qpLsS/RpSlAsvJMAcMCvk5IvfmQpel/CNKbcb29ADcFW+n
+uvUQyxVFMO3He1yckpks3f556t+9ag73TlPzsdMYN9MrXEmXemvEzwpm0dEc29HM/jXdTxzO8yW
oThhVViUjjvMV8NJcowxKbbJMEntfWnK3eI+Sk8qURkckIU0N3Qi5pKUWW7mJTYWM7q2cjstZUKQ
gEU5BTyflVCAxOD8Dm9G6L3HhVWL41K5R+prW+Z1En1s/xQPE4xrihP4PiXRdKsmDawoTCuNyk/S
fGR4CAy7x+ErWjt9z5jCN1yE/GCOMiLzPnGeubJkI08myOIwIUzCmI0juP4R1KbQ7BbdoEv5xEaa
T50dO0YEB5Hum/FC8Jf5/IVI/HyzglsUiz8BrBH78p50F0UlSOn30rNt13gouqqY1VB43WRW1S97
DvC49T1V+moIne8jjyuhv0RT42pobSrvOfskPBdne8tzawNUDtPNuhUJO+ve6RtGm60Ca4rJwk3G
XE5dNuL7Sf2qn65lg9wouInOBTOVc8P0B7YiukNvAlOz226AcrTaMJhM4EnLKkkrNa8/hJj2ZkDk
2U101fpSP6L+1aVgVpXeSgzxEpzQIkoGokoZFJfOHlEpViK/HmbE9BNHSKbjlE22BmZiN4RmvP7h
76dB3yND1vj1YpgAtSZus11oKmcDYZ7kq3WQ+w63OA3Ish7y8TZ6BLtJi88v/ZJw9Sly1OlKyp9u
6mHeVA/9oJNG5d/VxCySTadQ1cZm6sGHN7e6b24ksqVO3P3wMMzorzm1ByY/Q70tQE0IR5QjcpcK
Xk/J7dtdUAEw9Z2Rhi4uUGT47vS7kh7CfIOUmxyNsawSsE93I7RiCguiJVRarRrhVQCeRLLz+bdH
aJTgNlubjN3LIRZAepmT0KNuAmhn9LEjih9iXR52yp/klRqraDLYLCCFN0FUjRmExYbCB7GHt4sP
rmG8oL//gblibL6juuiUqvrs9CEjp3CU0CzzN4Ld7Ig6HvLR+EZslGaBqt/uMLPeDf+xMbhzWF1t
IjOcHAli1mdbklfBQYuhimfHPu3e1r2yKEdJk8QuonrX1Mnfrje8pZxAusDOrsUybRPQ0wgjrRZK
rg5FEK1QGdSmHb68xB+mF3zEN2vKqseQmhF4Y2wpFbGD8Le1asjWtHZl69uP6AB3amotcsi5vvx7
62ZWw4ixGPXRXILWHwgnf1nInCCsbxIrLpCqX9t+ASbm722ivzfI5U5ZNe/6KmaM4Zdw3HY5NQa4
K6BeFigB+iMqy4MCYua8Ch0o3blJs9LY+UFR5TmHR33e0xk3WKsaGIL8MCNUjJdEL7kjOTEVNTOX
gtn9I4UbWqILKsi80PhKfG7/J+EGX+VOGVQmPysBSicnGGq7rXK97ndVhJxMeUDfOD5DA6+ptus/
fmQDyagdLhuGD8ZgomxbLEF4iDtePth1ieeQFbi19xrw/FAMTbD+9QIUsWPZGCRvvw0nwmOgh9iX
/cGuNou9nLR1LDQpWUnLw+xIA3h5hle8fHLjMwRKioA/o0qPlOaIuS1z7UrnGQWH2VhpDZ3quzTs
WWw7b4S9+32gnJaR20r1CSfTwRZ2XzsSQk0RnJiSZ0IX9u0Qev9n1yTU92G53Bn+QVR2ES3pEGen
7TuL367wgmHxbGDW+uFwWtjXF8Dvalrxi7UiDKnrpChYhSan5gJi6wJxQCQyzQe7EZB/OzlipwsH
SGSUgjzPz7V+VgQM6ABMSPFL+5K2UjWkhaWGpZAszgfHEGtcchxoXsj7ODEbWgMHZcJeO4uqX/d/
oPs/BfZG6wTh7G+WLDnUJ+sqDPkmKn7AtRr74qpGDYGUPSkewtd765gXWJFBESLL4nbguAvuPsD5
qsy2FqYG1NZE165W0bEFZW5jxskkpXxt+FGvpf8Shie0RRU1bN9VqtvvmhP68CSbhVJWDHtbPr6b
PESAU+LPZpt9tnbmNBNCqfaEMF33DuQnYNSl5SSDOTfo7ZsIEfnTCCWg33pvRcQXD8b4Utx/QPY7
vFyDi9/t4qV3GMtXeNYI/tlbHjamFYGTRV7DZe+abaWahKF7ZBH1t8cI4Jpk3vOpewzYZHUob025
9ZBWhhuVqkK6/9Cy17/fhFruAYJqeSsxDIZ3yzKLWSg25acY0ONM0ysC8lyc4XEPeYCAMVtk+0M4
2WlfSltmUMtDpzKrGVgPzjyAVxDPeywB45DmCitbCyklK0MngP1j7N6tMI9Qojz0xyv+Lg/lSSvk
e3xzBXbhFBUUDTkRCwGyw/oMMN0Aq+01T5tIQe7HtfrtDbXmu6wWPKiLHHWUHy+RwFTXkUopchNk
ttefq15c7mxPtoBDkdWt/wk9kv0r6ORRTMbBj94mGCA0wBS9R0A4AIV9ha94FNOkRse6aDKteW17
pGZ10flR0PutbqJyg70NNZ6fpSCAiSR3uXXiaDn50GWwLDBLjlHTJQOI4eCqlSiqWKyL0v2I15B2
T+KXSzrjcSMc0F3fsqiL+93eeKCvFdpdXwA8PHeEoNEg3MNQSMLKG+X0fkqPyImXO/3i9lqK/ZRK
OtMdYjVgRBjeWPVaNG5jWuXmcD5n9ZBKJmF+IfvqNvI2e5eLmSW+4Zp/gr3dHhixy/vK1nCWyl3U
uKWb/NYALNgKpt/fso3eJ4jIwWN/1Mpp+fcTcw/aSIvhp/s+aLDmXMkTXSTNoHKzWLl9QkHjNYR4
6ocal/pg4xnJfR5q+L1T1gFPq+Sr8k8q8uqCeXesQbHQMgicrJwQxcjJbN7CUI+KSFRiEtDb0x87
n+1KlT+yX6Rqlg7jlK+yb8A76dpDQiP9wHQo1w4j4E/ScbddOc9MUOBbrqOgpjXaT+Fift+ArhBG
bypyRYNgggtMlXHSWKVif5POPMUtZIc/QL9BeQoN/Inm6OoddHVL0hQMh1qwJL91GpSyivOETSr5
jz06qo6aTcPpXEa80455zySkmGLNNZdInr/zzyRk96oMkolJxgw+D+5i4hWFXmZmnUfCuRXYgqL0
doB69alFO0iaIFLfHvajz8IeXiXMIkbnVtKNwaOYjxwuLkrRz6+MwYqy0y1ROTcHk7UNN8I2gYo2
w7HPrk2gHOolJ30dU798Ow6hLFH3788hb7jXgulb5mkDR6LI01xpnRAJbnm2pgofccPwPpHSP49R
3d6kCKpuvaQQa85VFkl7bm2szI/g7jPSjj2vFaCsDi+GuzQog3tS+pxaZr1cC5ItGEzgnAU1h/BY
YQuz0dRYSnW5h9+c/jKAQFxfgnJ2B49nGYbINNy3vzLVH1McLvQejWpOXE13hDAGgtfhru+fCqnQ
C2a7IiYDDC68iwUkiRr53MGaRk09kuvOYirF/STXUfEi1ER6L4KtLIVjEBTdcerRH/CNsmtglev4
awFhGJW+Rvxq8nEilc1T3OCYoMxtXIW+/R2zFlfz/MdSsB8omfuxm6kW4ZRSz4qSSnTkEIP1YXjj
i4o+xm4U+77XhdOGIS+GM1tfWsiNqlIjqSoLtFoJflWnvOc6gyifTyw8qIlpmgKd0N+u2UNK8DJj
sRI9s/emiI7eHOAq9hgKEfKrkHtqD6/CwJPrg49JciuncD6gId0+G3huJHB3WxBiv+Nt/4Egvg0j
Uxh1QLbB/ruq0m6MKtAdcsg0sy3eTdi2KWwkP9j17yf4oegRpuKIOohs2oEohwyMJKuFmdVGko/2
lQnZmw0rkZUsqh65eQnuFf2wmhVQdOjknkK6jTB/ve4ISpH48Puvvu42mJxaqULKo27eUy8GJASK
esaQYq3Qa5rP/tTiOM+BHaz88tIvm1bi3vCcK67NsHH4iArz/cbjISYODC/380mdwt+qZ/wXwqjw
YiKJiDW64bXJOLBG/26pqObN1W5Z4nqQG655xCToADCGZ+7AQSaf5sLAwQyF980hvS/dhp+gv17N
5yq94DV7gMmig/4xVz/L7iYQvHBpNxvqUB98yIwniQh2GPFDXX53z/4i9q2WiRTmvaQPvZt1JFrL
pFIG6z2ORuAnabtJaYX9m02LIbBLzDB5ynTbxXZ9J1hBJ60O7xFR925IQDRZK+RgsK/iLHBmGg7I
Meed2E32SNZO7aItam/c6PY+N4E3GOv6Y51kWJGgYu4wLrqwISWvuXh1GHq64svNCRX99Wxf3tSq
HU0Tr5ITvSpZS9QvxZvuSEZNrAIS0Z8xA8D7Cf3kD9yAZt1zNIVSI05TLl2ipvyyZZ6Xtbl6TZuZ
7CcTvPCVQd62RinnhRTWkqQdoW9ct7VwsxsZZHrzR2GJJ+Roscu3s7LYdebSx0qEjZspnRG14COv
uDdplmUuRivTj39omVh+ebxWuqDo8z1Hoy8BmqlfdU4UnLZJRnfyH/Z0dw5ouitp8whRb0RB99SV
MjekqyJuGbsauPRnG++H3lIdMxbfLPN2gAC0Dd01GQHn6wB2lJwGWhhTlHrKW1DqWoYzxC8+YE7n
AXPZbEHVfSavlE0faS38ZM99dxMNBX/Mb1raYqbtLdMk0hAJ2Wuj1vStueIM4xigFaRT/734k5vM
b3+ZnKkeKfLCJh50SIgIiYXBJkMAY4RIDUyFobW2ySnFbOOK9lYrk+Fkx2I0EJ9Z8+Mgk38pQZTA
jYq/lef1JlQ6CGN0QqfrmvvdTPOyz2Up441CJ+3BlPA6WJKFROrjF1CanuNGUdtnqBLV/dcmJ21m
+YmtZnV+NxbGdBvLmk4MlL9oqqXjNYivyY2F0sPWzLEE5yVLwkYqf13aKvw6WqKmZGlPP1GsjEKG
uQ9xQf/dwy9WcSVaqRGNeQeCQ/v6AGvL1C75c8/1KYGR+6wutk1eQ3o2UMeiWXu/7c3/+DsdDhuS
aosu/2OFoPE6N8Q18Qr+lseAj4lk7DUHLGthH0DiwLvWyVj/UduzlwZqp8kepk4myKip8eewhUaO
QLl5/c3rE3Z/jbKCTQi6iIDMmMyftlC+ZGKHxXf4O6lha3ol7SGTzUWUGFauEN3FIiuT3YpfIs+o
5DWDaJdX8vlKCR9UJ+nDNcqI+YgwaF+velW4EeUVVYGdF9HHwxxVajvJpAiH/Cbu71dxb/TrebvJ
57BNQQ3fkW5ldKlDMNa/ZfiYW5S6VIlsx/FfvRJN8B0t4eQZVLnX7B7oQYVdv9oCXCfamfcqY9Ey
yKwixIj8Uhwn2Wyf0MGnk6cJYG0t7J4CAea/DcrtomJfZKVyI5DHoQJH5Huv3/2SKi/Sa/vdcs0Z
LSxyj3Al5UZRv37tDJLv5RjHQRGCMnh9uQsMJuZeqUnjROkLiBbHXOEnknHylqdiPCkdEMRYSRQc
U7fZ6MpJt3gSEk5SC19yIl9uQBK00prEIbedsUk4FjAprqIblsWxbG1OmjiGYskY+7qbMbYe0b2L
XKJhzKxVwv5dRWrTUHUhN52Lb+/i/B0vU2+lcNjzdbtafkpH5TO9P9w+7fNehOqGQWDZyhTnYw7J
+6jrWQDltYfdHpAN0Mh1N4amfY2VjtHZP9zz+2TU/SLyMRMDYBomYNPpL8DDvZCotuyII7yrurZA
6m5Aff/LBvech3zU52gTEZhH+eRCjs7IxOctTw7AeQeNwaDju4zBCwNV2ic4LV0Gs7mhwevQFeUy
9NQfiyV8CN71pLipEmuFv033AiJoPEYNRMQv5LznFGoMAS6WaADuXk038+D3OJOGrypndi9+eyLQ
2AQ67mDMrtxk8C8OqqWcRQd1elp/Sp1+G4j3Em3SYqIju1ioseV/ezofNuFphYygwjomgSktsR2d
kdwSVFbyEaDWs5WJ+PT6HA8QsjFTUoSsw2axnkhUY595xUD1DXa52TmOemc152TRUwZLBSdmT1Ns
K19/WApHlUfV/ENpBwtKYInWr7WuVe2kPIjX+B/ljrOhoglRFM6OijsRnf25+lrxgP6Yo+Jnk1c8
LVZQCGGmDLCYNc8n3pJ9XsCUxf14Ue84/CM9P8R6i7KabEBViqqs5q6SUj//Mf0lFUzoL9fYvmKm
QWDxFxaZQLQd0/xjGkY4t8gB9xP1w7fOgNk8oCVUEYDCzpJCo6wjd9GFP6C7y4myYNyjOuc6f2kl
MxlnYLAST5AErVV9sRI5V0MgC2z0FqHXLISFzeOoB2i4n+QhnI83rBYSG1HhD6eWuVd/gJ0+kq+A
ud1wWoYXLHH/GUMNm01wxStZ/JDNMUH9GTD7HgHSvzejTkRzNo+a7gR/KAKBgBkbvLAqR/ZBrEGx
Ay8sQAw/x7ReEkAie+jsMX4tpmAmZnbvuLBrEzPWP+iakEuF/D8bOXeZEnIhZjmj14cTROlX7yFr
El8n49t3VHCiaKt95BZcj5As6fMun6/iw577AR2kyFS4vYYm7macXmLszXiSOyVx2iChMdVPFOyl
URHDCL7iBcpLqeVHGQWPZR4q2DTvnkXAGVhkNkbvmC1kUZ9oBLN6897Ld1rtXgnOnnDHCpp3okqk
qqEMSt2+MpYVHZ4a+NgJIa0uFlp5I4LYBZBdxJeEm9YMrrbetcZXAh3I6Vwmz0AloUOL4ffCVHiG
MbwY5eLC6Jk/JwaiDJBtlX6w9xQeT8meAVaqE6mwX2uY+NP32BCMxp5i0suBn0g1Pyqs/nLpwRox
602icaoriz4+q1YxhzofcE/NtROU3CwMWwxj3QPx3TJvKse1g6KU4yBCiH5mAOehUJtZk5HThxmb
KhqkzuP/D5SqpxljR6HsJ3Fg6maV1pvMf994Sem29yTDFvWxNYx+/Tp3KAluENTqlF8fBaCuJwZ3
Tm98ruYQCPt4IInYHYdZKotFr4Naqh42nwXZEjKtuoGA8QK8J1wbY11Yo3zFtEAdcgPXjdWjcs5e
8u3j4SQN+p2S9JAZooXmyKuJ4c5iUFC6CUHYRH008AN1/M46bumjJ1yX68VKbTi3uHmeyh+k/FY9
49HPfArbOdIcBKCEobWrSFOTaMCZtVmF+2fqnKwpB3auU9v+aWHKKp/zBLkvjpdYSIzsfDYNcR1e
97obfX+By5fAd4M5l6TpXpgq8nt9zQll0u9kqCGlMcR//90Zn9C3YsPI4V0FGQFm0PN+zS588Ia1
OLChd7KKY44KndUm29n+2GKajISxrMUE9lduUSW/2NcXcOIJCVVP5QTi5gx+lAFcA+l6mg212mUF
jAYoHosFt1Os9Jh2CUQdC6n1MhGPECiB/d53ReaHCL0wIlEDOfYVZajZV6kwdIDTZz+vhoX9te8u
Ggh4rJIzV57qK/xwOiwFhKEwjW39WzrJ/c0fHW4HcnDs7WHk+GLoecwHkDL/jOL8SxDBq13yjYt6
7AKsac/Svl+d6ke4zX8Wp8VJWiEKe81//LNJpugsCSBOGyEteZ5tAlom0+/epabgLdnlKTNFojK8
yEhdSsmCEc30Oj3g7TB7hbDt+uI+6PGKSv4vJpgzcUK210s/8mAhRvF0DXWxRyADZLgs14ofgwc4
i0GS60WErEEg+WK96mGbnZEYBUCOvGfAlTNb/33B8NR/oYvm5uffJ2Ie2mlvnPWqVdBLgNOFtf66
spm5siIZJHG/nS8DutWnfI7P2je3zO/ETVdiIK5oaCw4rDXS3G/yNxcxzrvfS6lCfh5k3B4OTRif
2TFsjBaHIpFqMiqBtkhYDOh6XOyZJYEjMnF2KoEuuqS5TX9tOM4+/McotXZqFqhSCP5eRTOoCtU2
t5ZFyl0Fu/ShoUIMBwCH018RMEkOE+E8dqtPBbprexcno1PitdRRFN1KPt+dHcpLk5+fcEo39MDM
ZoDWCHVrw38n+v15vQF3zqyWYg6m1ldtmXnblR5Let6qxzZAYYWV+Ytxzju+BdHI7T/YeAPwHD8i
hKJUUpf1aSAlOjW/amKe+6L3twpFivxlQ+CzpSgeQtpdLIryqPMAyif5hm/uAvN6EmX26vCvCgw5
UH/gemEy4KpIERhHgo6y/8JZN3c6agpZxY0bTfasWhApszpawVfN/EdhZCfgbYYCOdTJ6w7FdGnc
Wx3e9SIq+MkIBgeX+BIaE0H9mYpHnHij+Sk2yaO29X8xX5ATNdS4gmOvC5V2tDRb1YcUjJxCvzeG
++xrqHAET6+t/5YXSioZAFL2S2Ku4rrgyplV947VmvoPpnmNpWecZc/EyHm+KstzPOQYmIMBokcd
zV8o2KXS5FWC3wfOZL/vYfOQ4Ru8JqCXtquWUvXtHFDPhJzK0gZPE+AFeXtqoLaOa2ni1ALl1HbN
oiHGRdHM4UhiYjZO9kvPibaKzeDwPiB1DauNavQnHTisHNjtTcvY7nk8ufaEM5epWHU1e/6jry8t
vLwg5xsutcLIgjFzgUFuJICSliakPz8zjZIoohpPIgCubWjfqKk4kPiWrYau+vt2UYGuK/HpJNDt
RAZ9WBBqK4I1TXpSKwNYvXSQXdP5JnxkyxPftFjAl5Cmpg51s1dBzaCr+lbOS1YNd3CaU4EaHIKS
JZDIYyIECgv44Jct23FiLruh7KhNN9IrnF6SJ1Qqe8u925/zYTGWOiPkFUfz0kzGDKrM8ER3b9H6
/ZVOMOhrzdlXGI71XUrR+HyzsXWuWGl1yt7y1s9t0zRFn0E3GzV5YQNY+pA5VtPa6n0k2hpP/+z2
S0vq5dxzbPIo39X6Ih3+mBZ5aqWhEASrG0MK9z9IokvacDwt2tQb8o2ph3ppOEdXCpE71FupmGwD
pAiHPpSU9brr11t1h4b5sThMjG6ysrNgafmk8EZjsS/NaEihxvvJnpCtzZiqCdrhpHB1wH56yqoM
OM8i28mALw1EEyQwhZ8Lde6siPLfqUGTGLGSuXapdJArejmUTYcIxldbaQG9JklBXmWBpCpPJcGx
OWAxQmy6HYG0BHG1d/HJcywSiFkdtppsRLuIGZJ3k0LwczhBxB7g1iZH2FDlu/EQ0cEnb17g5P/J
Cf9EoZQzFU7iy6wszQzbf5aOM5ah6HyCEcoP5ulqxbyopQlOY5Tum+7sVApDGTR1HONa2Q2+ZiKE
sjLyntpc52jyBrUENlzErY3wuJbLROx16aNXnYYlJBOVwwjHLLza1VaorhGk+DZhU8HxgnEpmKBo
BRi2M2EcKp4Gwnz0Ple6IwQLweRlMy/O1o8FMVxX9nXIy1/TgE1kTbniMrIEvdf8Ua2rLCK5psFp
L+QQFZzE5Wp5/WlsxNA57ZKzp49Vx6P6nL8SIBZ6GnI6/raP0D0ld6zlhjn8r7hptI3Rh9n5InL5
yVmM9y7gYSlkepFFclGGIoJ9G5wLWVALII5XM/y8sxLLkRP6uOufiOoRBqmai7h9C0FNmBPxheUN
IffhFJybgnEFg7OPOL8MyzV7E2J+OU1NKvK8vbjkWkNrnlXE+Pk3VEyJR1VIqokeeUOddOqz5KT8
FUu1GigEVpX30oKddSROEtli3eWxe7j/EjC7pUSe8UN0qbeMJ0i60g5afPZZ5NIsSFDAw9rCrG10
jffEzsR49ijzMQQwfBdgwfUDfWNNUwTKNH7YMgf/1VQz7riCVJiHro1BVf+BVDwdgVXSlA7p12i8
+fIDpXOukvzNapvM/7r8Meh3x4ZuxysuTuSqFKlm42QhMu+f5M0yYqnh6dFLnQ5yohBT5dDS8dqE
L5OL0R42pXn7hgZDeIamuy1TMXZQ72LJ1M5SvKZNuYs79o3oP2YBighmsyluK/mizR81sGFLv5bB
MP0QbZNkvq/f6kYShW9nMySbcgqAbBhpecpHeucf2W7yojnDD8rQ0kK17LAw76jO4C+N8Hrbw+o6
K3fGk3cNydSv3algaH+hXgf4xx+dgQB3avGa/x4Cyu17RUVfsoPAd6Qb7vt4UJCFVpClW+5ttW3B
2ysw2QyYvXvyQ0lAvitdkYrfuDB6nHmRU76J40MRmxt+gRQIxWHaLMMzg/Esftwf8K/JkyqP5qgx
On3s0xsuB97tDq3AZKWtFj2IMhCJDurs7jyFsnyP93oRF1YdS09dwBHcoogg5WWMr4Z1ZDuO1vBu
xWLi6/42SkUkowpS7YbxywoUQZZCcfcl1Pn3lFcKD5AzaJFvLXn6vQBljXeuAgcIWcb7Zp8sSOe6
38v1wz3s7NUozi2O/rFvIWF8Mguo0wscxl4bCJmjIAaGgjvx6lZUgicCrfk0gZoUgpb6rKKg1PuZ
JYvq79Kt8ydSIFjw+yzsyGvxR1/SQXTq/PGtCfhJ89eV8ioi9mYHoDoV+tjvzAIRv/nrflLNxZ44
OJlfolVmD1RFWJB4iLLcqumbmRmRSJeQwUl0t+vhYcH/KOhZh88LMzJSrN/frrM8EMer26kpkFgR
JJi3oQqm2RHrdmhNrCnRLc3Ko/cJ/okjvniTdh9wwUf1bIkBE8BlwFsmMxXw4rl5K7/rGfCNu/hl
OC+zEaWcYShIpmXV/Yo2WF8Ws3/lrHOcjdZFJtzjg/cIOPkxY1OG/ApRgePMKZEp7+e1nAe7fOmA
EgaBrOcTunngjTOcYsCS3Jvra9vlTAsvC6iuHC4Vyii3TLCwMxM1j5eDW8fvN3BaCzREnX7tZ4I4
TLpzzbR0lb7XVOXk0K5ZP7cvu1C1dYAMPlQnkow+R2bxbjUTs1Nq4nqadR5Z6v4v6zZofWSZZQmu
3C/V26umzkt30palHGzvGgEveMslxBuxfdSGNI2DLh6mnbIAv3Wv/yI07PhPm5Ka/6qsEoc/2hpz
E1MORBp+NWpMbgnSUgvXCY31bhkzXlquSvMSIsmGiZwN/rCLWvFxoaIxWeLYYs+fWNaSUg1pBq69
5VTxlppvZ9sdK0AW52DeCT9VNhXi4+s766A22L9iA6QzCcBwOuFgHH6sD0wIKZLDdle+6y1+fpVM
+yZQgi8NqqKCNt30mmPtVzUPAx3mwK7YK0MvBGd9k6KEzEKwuneBml2vavDuYDkmYx7RGti/qSRJ
L7Pe0Oz/0ppHMLR4xnBqimNXDE2LBbpx7ppd+yi7lumFwAWMNmjgR1YfR3hWSix79mbhKee26G3N
MsorKLV7OKHKHGbPNRY6RMc9dO1xjHMG+UhjDVK8600RtOq061GYqIA9PWETehIukIQzKV81V4Iv
d243KkgJrGwVtf8VI//wJQrBrfZDBmDjxmP/ubu/EQ9i+LZC7WOqTA3cVW7EUG+98+PjWvFVW94x
OHbHE72D8kSmX5Vf4Z3e2iwDVcP8Yg9mjgEXQYommoe9jbKHAUwtTup51MoVNNpLdE8pNZoBExIT
200S4uak1bjBJk6+P+5Tr3IoemnEzslzt+7Z8U0I5FFkibouF26ChUxaZQ4AtBSzwGiddhDfDqaS
oTAer2uyVJPTN6ltpq7M9gq26zzw8XUw9Z7Yd2ocPoguJ/izQS0/2jfT30/77n8gG+Hh8fvC9LVe
FjNkZ7zalI1YpO2+3exxs4K+MKWkee7Z0sHT20Q5JQOUfb87M1h2fSuORH8jzO4pCfL5JKY6obB3
qN9D64ng8yh6tJWxJEB0UOy1K1hlpKE9ZyH2UsqNmLLw6XtBL5Ipn4ZLrJ5ru2xGvRjwwJhj3UjT
KnlDBfJ2pEBy9oAGWJRUgfvWERCIWwCDZn3niPZBumm/actaedMsWrE8wHZx3ldzxjarFjTgP2ud
dIIFk9rmZEUFaN3XmOToc3cuI2DjcuLXIL928AtJnjkqYXr/RxyLiumTKihBKyiI5H+TgI32SdeM
E6JHE3nHN/VOvTuICisRletuUaIvPbPkJ9kcEwwvBI5MPGQS+kZGfPNTzyxeJLqbOISq2lCrT27P
pb8/dUlO1GqJRLv0/vparJeZa7u4EHho5KNbX6/j3tj3vABvRFPG4eFS3zxnhEcCSdWChRbPVDkE
zNw7GIS+hpI85rA/xNgHHS8vFBJOKK5Dg15zeMNM9dRRf9gsi5dlOdgFk9uQpj+nIQw1udIkqBN4
zkBzFMpxt7/m51VLXJh76pbiyP9sUYwnKvOrrFAs8oGE2JO+3E/ctkArhYt7BE+VF91/Cnw6R8w1
tlcw6WMJp7B+AFjRH+UvVxJp/8/E+Wb2gn5/AFvM8cft3Q5L7OTH97k1a+c314tEW8PELXvQ2Fol
7mrpRaFf001J/EYGPie4x3VqDboJYl9zKr/Wol4jtpIro/NeZGcR/3r+z+UcsU1Yw92+c5pcaQp8
4xlinJxchrULteoaWHiDOR0WqMcIeaGhP+m1R7KpiF+SPzOJ8xik5Y4Nk38NFZPV+WqrAaQrpLUX
rfw5n54b8kJKm9c7bT+4dIDcXd2vHJrzebumB9AUakwOJQeBZ87uG9kHkDrm2NglqAR/9uBLLRbH
famoljeltyXsrW+67GsHELGZdchxy6nHJSk+mza6yI9v4v8iK7xbfwgwoFuXKkR84FB73K8N8l7c
S2wdKg1BuK+UA4IXKdYu9RCR2XdHh0qHdYNJ+xfID8dqYkFPr2c9kU3i+Rqh5m8bPo3ERBBMCYkO
hNn5xHRzEf0z6jGhU8c1fFXwmThfOMb1X/t+AGTXgohR/F6ac/5n8x8GpBv4B2j/vfCGlW60NI2u
bpuA8SUuGqjKSC6UBo1fWQQbWASP/HGmxadEeLnAb7bNrWGi45KjjVGpNRknlsRiIe0M+Y+rIZTw
1mJc71ulSO5uYXLXmV/HqRBRUv4qq8EpWbeNM2jxe3o5fFjUjp9/cAmKnHGzSTZ5Ic52LGCIbdIz
xCuqKETSLxYJVCwWCeNCrCxyu5bSFkYQ05wXHKhsKSxlsU5hsVym6jiUgvoDxtmmRkOxYZAKOdNs
RNkNOaDiJ16d+Z7+VeJsHI2gN/xDqOGGvkqIrD3zIVB9cbUW3MU/SHDbSVFReR5AQG9azdkRToQC
z9cG+XJMpd//3bjizRh5OGs86/PPmG85cuioxRac7VeeHF0jgHmgJvcAOhSf3XKwigXKkKzNZeLP
5eop4CyorX2vkRQ17b9zEEfNM7ZM/cDAhXYQ/p8Ra3jDbFTd04tzbYLBJuLkoJcw1elr4/JrLwr9
HyAz6oLJuwlkqNK9vUlIi6bkCDLafi5ThKzGeeEjwcO/ZNvbiXWiH8i5scEAGlY595RoAG++N6V8
ZpfpKCFsiwC7wG+462xsROKvHssNGekbV+YWMmh2zOYRwiFhwVYX07tIqBQJuF4Ykx4RMIiQYPOX
9sa1C+FebJhNs6MRlrYu5kg3DvxWSNlFGDn2AqDk4rX/VOWwzll+xG7Fcka3xsdAg0V+hBZ+HQE8
b91eCrFLoGRTEQbRmPxh6bmpZtGPOwwKTykx7iYDTFsfE4hwyw7o3VYwvyOLAldMTLDUsXmsRqy8
BwbB8nqr0ZqQzSfllVh0sU4/do0pFvXeSIveC617/VvUfQxWx8eQEcwxCIaaGoW0Ea7O3TBXGr2K
h0GowEAc3Iz95GIfaLJRskiDCeFpdHDPUSUwpGvvUok8EFnCINh+6aPzTO3qtyFHNxKbNqaOK8Q/
4mspGFxUGO5Epir3wUsAwJIfQuF1P048cqMKKK/7q7WLcCbPbBGk6TZ6XIwNwQ9LEvDdyr0XYXG1
Sm1mKpMmKXGekDgo2dgSPiCxhPyoSGs9aB0zB+WwxHPi16mBMTezId0iPNhunxVxnxKbE2c7jUHn
rec5MewPEq+yVAypNOttU9wnagEavnFu3rGydSevboRWuYijpHskd5Mm6wHpEPBg3Ozxf2qERNvB
NymQMks11dChoiJDddFfaa9OqJQEKNANY8MxDc/5DckwETY3P/1MdHGl4UAuGmUiB0zs1wGCxM2U
q1UKQM5qxU0aUkeJBGpt59I1hLm6TgmHXvRnPyYImyZ9EOsksVftBUPQ6LBIL97eGxACo/jtRZHt
q8LN4iTB2ugVnsCpdCzM9y0O4c8KmMEIUTpdCBV5UXGxkxWQ08lB4LaSW+TpPaFOxbnzaiNtWMMa
gIpdhhokLkvsctEf2XkIEd669rtKU96b24Ph7Zc2JenXT9rR2nIhI9Bkxcnt06YN1ttJ34YYmrvE
aYa0wpDCARC2Y00HFek0CmtFNLFhq9ihy0jnMaH00gqz92vj+LgSVJmUl86XZIbpEGpjRgo1WlzC
No1ehEMz41fIgr6SZIU8rsgDYxCs+KRT2zJMfo3REopjCuRpCtZ6O+eYpiUB+Qq0/KpBGovbLP4F
6301WELbS8A/6M/oJSICT1U6U/dPh254AY9Sihg3notzYXXEUrYOuWgbTuCmoGtt6ojbyjh2/3Ls
kUOacgaEL0EAPB13B+eAoiuC+Vb45u8AYxqoT2f30yR0P1v45Agyp/oMSH4NLQMg2srB161461DP
6qX6HZXlfdGqF8CvyE5D/eSKEsBtQqy2PPE5oLj5i/2Iq2JQkLIUQgngURsb03z/NrFjl2PnFyZb
uGSQoIFfshGONFikrN2Nq7MeynAFBo4d1PL673sJUcDNk06lp38MDJpI8B+CKfKqptMA9M7Tsc7N
haqvq5PUB1zhep1CEKgGiBavTEA767LeOLJGK9+FF3JV1F6gZyyOeztv7shFsZiQviyeNqYprjYr
p4stxpTqDyFbgze4L+zNmz2JkoC0I1OFWOBMUNqHrjsDT45ffyJmUDjKM0OpjkPXhzFXP6n0DRfU
8tGBpX5Xh2NHZV1QCzjKxYL0NYE0pNK25CSZUj0r/SoQi0TJgJSqm0qhsT0Uw102N0NXSf8oytnj
EnWmPHABLyDhMim+K0LSlnViqD4XABzisKolzkgcpa/OBAxp4Gt0mF/ufLxy4s0vg96EWmdPTced
bTT1lkutVXWjyJpaCVWM6eP4XOteH61A/kzu5PQ3radJ6x5NgX9mZUT5foxcHVy7LRx3nHVjfIFs
6qccm9ckVDBWjf5hHbWb+gd7kFjmsbqeJH/MO67/gx81Ftpq45R829iXmtNFO39iFbRGd3H9Hxc3
QBi+uyXpwzSN50mLkJpcriDukhYTsNIU/K66o+7QtHtmxbnNRpPwKVKwjUpSgscbkVCjaP0yZaMY
ibDBQ8SISxRq2uxQe8IbvhQIXzZVlahCbz9vjy3IkKQZWUNwm0+3xR6atAnIbaY7Ha2IVsUhgdFq
MvuL7NdY2nBGCYQofzdTluxu5UyStro9aFF4urfiZjAx+Z/pVtzsrYh0LVXEAKwZ/MMZa+NcGyN/
ophd/CW4doD6Px+vQItxHkZNEWlCw6fdeuQcCZXdawHMoeHC502ps3ss5enF7QK72B8yNFzrdB7n
11KrlG4S4PIY7Y4m//2sBQEncBNdoI918uhSOCFanH+2EGDxq7MrRic8NJSAec33y/mekKhFg9pQ
PCU9ZkPDwnfp8MDZVKnPtWTl+v67NUwxmlHiyH1CLa9KVLUxkCMRq60kAQtottBfrp117JctcZJT
7w8/H69dROptHLlTbF60/DTSqFUZCBhg3AEToFElKlHVCxlbsKZS5ojtpv3HaI0mcsmoGnZKKikW
olkAMlqPSuOn2b7J4XL01YJ2g4mtbWKj+WmlLuZGSuRDPfqGDftg0ybqE5ULDIlLdXhUV2YJD0LL
V04yDpeFa9jgItbbQ6/6ooYoyFL4njRxQAXznmlubScTyXZnsH4ZOOzL/R66z778slGeyUFuWdFO
FduNjI64/TaEjkRoduIkMUUp8QizEnrPmmqZ15hOUxhapuX66kjcHqXKwpb1nnK7gvTUlgI2OJUW
s9jfJLsH0p3g91y/z9tVeMgdwrmAVuxMTrD1jrMGE0i6rc0IibhGk3/PcnaaJPklH2POGIP7JX7R
srQ0FAcwQKUXA3NOuycJtrPKpg58ORE12INfauqth+bnqOqNlSGCr/TgSvyxQpluLh3nMHujPxwg
LoEzRF4ls1vzx47q3BH2gi9+uQ/bcl6BVHf4IcYXwOJwSMMESBpCCXeoWz1KsVg2GDLgiOCkC08u
BrgYQBitWLkwIa8e106kLQ0SY6kAl18WphBsUGyjWF7tEGzxk280Ikijz+2muZ9euh8nXSS8Au5M
4GLGqmbCh0wJ1WCQkxUI9+FIfmnDVInGciLd+yyscYAYg6KenMe7flrHXttO7TeczLrddFNi/ZJE
Eumbq8/pr6GpiNJxzPoG7pJGHZ55P7g8FTplbpNORBVAoFmPuSAPF42LAZtv1b1Q2nTFY7rVzes7
ycGiRJcF9NDlyUsDvo4c+pvtyHjSTTN/yaLBXj0RbMOBijdMswPeHwTrX533X69e6rjVV7q9qAJl
0K1/LIjGU3tReA1GndVcbX43tuu/PI6ngDmYyEfMGOckrOyJ6AbWpCNzxl5ZuIbuHPdVsN6EJQpb
441wK0qmWmPRi6CPIHc8uxE4noS3CSGkioP3wU+MMcyOWKnqOY0C6gF0TZ2X57/Yu7ceBA0ukcpZ
1byMm06A/ohZfPiw2l1ZasWie1xXtLiVEvuy10MOUYFURyb2Hz+Zh1x6tJUv90Tm5mi8/B5auciw
Xd+D1B5FlTrvo/G7nsWEHJTAuIr0JSolvoSuunCQVGvZ0Dnupo8LF1zYtblxE0TxCLeSyEs8L28b
HrORDwk3rmfkip6Gn+KxTKz2E1Lim6W9xqF38wTNaoHf/7JIXLY3VRW1iRdfhyS2MxKWdaccDoxP
On0M8OTl8brw8PWAfQqfwK67UpwYzFBTo7Pq5lRAk4hpKhwqq4MlqjkG3JZtH5XTuTYEK+ajTZcq
cUqwVemK1Ma4U1Bmv8rRSsRUsixfb7zUZWf7CM4k9AWznRsaQaAhfWLu+VL93iJJpyiAXy2Sv5xn
w8n0hwlhUzlbjQyiFAvjSeOPmrOf0RFo67lh36M1UobSKZ6FYE3zSl+jUPD8ZCh/KwGD99Gj7CkY
9VKQZpj1hcyn/PvKzm8adjznEDb3HsNphZGCap6BdVQ5WyDOFIJTUEIVoXky7gSTgjbQIZ3RKinK
UGY9nZFlGkJpL+Di2uQEysouHfE0yuNJ1Rptc9oNLjQWSqyhgvAKoSIVYrCb0MZtZ1KEA2Gb+ZXv
u9VI+QQeOEkaBCDopHV0y0h2p6zvHbeBwKnYp0jP2cS2+AJm9GvLm4aW4LZ+7IhLHLibyXoJ4O12
l3dWtqUBqxRvmWPZhL+KlQWRlbT4jpHd6fcwc/vZIOWAAgQXkfyS5yKD9tQjeTgt0Cd+cvvpFDQt
fSEyfctV+KdXXdKQdj9pw/uCaH/4cf0i+S8No+qQ8Zpil0VtpW+/puGKUJbmj70aPgDWLOp8s8Iz
xidLuEhvUT4n/DlLQ+/sDDttYV3PbiTQunqc3+zy//Crnvs5266uqSxDUrqKrGA+wkkLxVA2nQsK
q/P/qo1Mzjs3PJPveqypfJ5Zy4k+71FVpPXW64rqXzcGUtTi8Uk/iK2DzzZY1Q2mc7R2qnzGIRW8
k8VPuVgdndpTdHDF1WlSd7ShMlEn+8jvRVmDnLBXcrNBSllLt+cqGjdp6MaI8AWr22gaWWEIVKtm
oQcZz4v/OgsdZbaZCTylOoy9wvS06YE7dUUvJkv5M553CEeC8C3HuVWp35OCYuQGMaOHOq7YARWv
VkZ70xpqA6aEv4DBWYeAZocNymjgihBg9mLgtCDhQFKMHGGLh41WAGI61JeTTQ3RzD9WBehLbEFf
xO6wXtrzGEADHd1IAclBBcId7xQ0/ntc4NGJvqVuQL5hv0DyzuAJk6GcHpnOE6Ln+yGWSKhFzNeY
XvF2BnXHZSinCO8DVE5iMvzChC7ZUsdOre3djgF8AyVt3+67z7e6tOoPPBqajqCdEZ0rCLMLVNcA
NsD/xeu2HnmvgmJNTHP9zq7iju6mcF2h02/QrGKDvA8vRmpSyATnzOG1GqRxRq9nzZWIG6vqeOu/
cNsAX3bu+mQkKaeg5Bjs7QnU5+xFupagCXab7P1VPeVelP1VBdBnjo6hH0/jqZDtya6HVAAJfMKP
3ftPXnFJPzpK/Q8PPerflpTHSZoff+SuegT6Kin3sFihR2yza7RbuXazAGetyOGpAnG+10M2K9YA
QrtsoOStza90flIzKm5u/ioH0AJEVWV3O+Dv1lyUQkc4DWIAd9Q/Iu9iyY0mtaOzmVkqYZmL5vcB
alkTIzuLSTOssvYp0jfHeIj0v6yoZZS5/21zvCmUY56Z4JoGcZKUC4Ax9WJ5IU4Pc/slC5m82NvC
66blJShvdTxpuEoMiFhM/xCT3Fj1J+Jxczb6qrM47Wd9TILx9KzpRFHfxrlYus2T9xpK9VBh7YkL
4IvaLi0qr+kNO/u0Eofn7P4xjlV9+eqZUA4DX6mXocPHpiwNNDioTU6iZ+JH3gznXHMgKqa1JPKt
55+5m0bP5lbhcZBSs1fCx1D6MrKRGcSxMtYQVb4cSaHTaliRfrwE69Nu1oGPZC1M/911Ghxhnq3h
dRHgPwTtotpzxlFCFemsUhmpz6WTkZk2CVgZzjxY/sEq0t1+B7tuaiMSDcPWVwpwPBqNp0+Jn1vb
oYukmXFo7OKbdA1hDfdcU4YgbPFMwpJxTHoWu2LVYVkWyk0+RordJZWKhrm8SoDlJzbe5QrQczZL
WbIBf3AMIcDQHM+DCtm8z52WItlI7dIuzzcd0a2PWEmYN6nm4noAAwNUyMyEDKksPblsarclldeU
p8KMXca+tOrs45XWlXyw3mlkh0TpoC8g3vrtaL1nQisD+s85+AWI4/zcmX+igzgiaFPgT/XepDP3
BfjwPPKP7xhwlxBV8/Af0Mmop3xmPmyooaq9cn4yJpbFnSmGRMAR6Ukye0DTgvHd8DMYq/2EXJGV
U8OOzT01NZhlKxP8vSFSXLDiWTm6KvfxpPqIpdtbxzodVBKIAcrfK3u0sDZX/7MLCcwZkr9HD4yh
8zt9Fc8ZesFKNysNGQBAmVh3CN4B18giPrMVrz+cMTBL9DSMYSntFsYYfaiOlGaY/N8dZUEGd7Lk
++TaqysWhOLuBlG8Esj0NQlrBwWR8FI494UZb7z5ediyLJ5OnkeE20zAK1tVSdsRrP1u6dehMipX
Igk8KfuLL8wSFqrNYZhmvBadkt354XQhtUTIxDx8DRZw3D7E/18qEgU4cJS9ojc6GlHGHuXELBAd
pALRVkr2LgonO+GbxkpGpwRd2v9cxu3olKA40G9wfPuH2rAeJUznaybeMED+tYu6prasK/rlRbEP
TwovshzPxtAIP/sgBI6/RjAotQgvF7Iv8DnYiILUo8DeGzFUNIWwqE1X4mTnwEkbEuevBcgneKBR
sR6m6CGCK5VbeHcIdtodAq7veZnffCUFc/w7tR9YIA47PcPbzZpD/QbGuulenlP9sBlJ4DmLOesE
l16uGgQR8pnWF12kSFjm8BwKZH8YprbDbABtvDEg4FAlQ0MC2S85pu/5Q+5ev1Z3k45xPGMGxB3M
KIrvnHj1N7X/lLYPReZK/ejI7xwSTLWpQcjVO4qcOpdPyo11+iPofUfjSVFUmve+pU7ETwPel/VF
k4G/+n3nZPTRgomIKa2Xx+P1x3BcmwCn+8TTYXLmgENZ7WbRUDTiKXYRVQcbB+AdAusOIdSOvEL8
tSOT5jT574S2qlP5Xpm8wNhraXoO8r7VdxEiTBm+kAWSCz3W5PdRL74gs6YDBWpNSz5XKb5cCz7+
oIqo9cNPjncFCvoh2WkMvVXnn/P2p1iFD65sn9vbLWWDN2CSZ2cEfnuP20TbEOhprjCv58kr1AKu
7Q8yMzLqYEaFDBBK19Nk64b4dEGH8KfRoXBq1gfk7F4XrjLWIeHM0xsbM/VKYoucsE0bcJfGb9O3
uiPO+3HBH+yrcH1KAEqtQLDxZ+xhFsUyBdaT7//meIzYQ8aR85pd4NLxfmFDQDJTxwnD4fSActqX
pAGHFFTJZRDI3SGNwv/X+FuUKd9KPdI1vtrr2X8szP6fJeFJowQ+eRqJnmmPNKN/8NSdRbLU9I6D
+ECohFlNf7Nnb11+2XYhM7e7lvbrIAAfn15z1ViZc6861OZ9GprBAdAOgA2JuEi6HzGLEZIJ37Rw
WWaRu39htxtM6reU5AxrwfHvke+hFHCxUXb5eD20xpCS5vZdQUJ6ibqTmM3qMPmnccLT2wkZNqm0
GhLIYdPks0PE2zhmD99OymcdNqdAtzAQ7b3lebjOaZwKQdbdLDIdx3yL4Fra5PbJFr0w29Fr7bSF
CJOxm5HI3Mt+WHpKM3BR1d9hhUOhoma5MZUu948EEG2aKrsrtJ+SGW/HUOC3DEaBqixJvO6d7rJW
jfoqZsCTu8wS9jL5FZXJOrSREBk+/xpZ5cXXFGknilfL96fqCCPdQhSZ5ISzqxtIq9GPYfxvkrwi
spo+MYigHPb8NgjVNk99KytYzpHioCIX0Xuzk5PhVKx9p5aRBwsYAryz1xFx7bdlbrWV6h6viJji
lmossne1SmlbNQDOoCXMhU3Ih0/AqO7y+/7ExFOhy1l5K13QN9em/BvU/h7Mpe2LVsxcMsAmIuJa
3Z1ZBtBm4dwHtXn86oM8/nUiYaV4w8ifSRISgcQmL156QnHZ26LnDF3Q7WpjSJ4ezuTIfjJziw2/
6GQCn/amHLgxciRbHrUUGjGR+Q0GmI4Sg9N5vLTRKvMDUc10Md9lkTDI+pDVH9lvfDZum2uwjC46
jkuuOzat3fjH4MyevZM+9dRv7VLI5VaGlK2tTlTbbAljunRkX+Y7R4Fgb0BPiLJOOh+9D8zBoYht
A4P82zvUNVAmE/74HZapgnAgLZLjPi18fuD3jLbntemXadyzMu2Q+Js/2vjT0YjiwolpzbFMOrSL
QVCfMNfEE+0AMRpNjjkJfY+ylIcbxZ1ANBiZ7BLyoFx7ju3scJ/92QGLm/D+zOOgjEureCBG0AIC
HBG6z0H5KxhOnHYquy124WlMSBXDF3EsZZVGH+l3bUnoHh54SZA4ydWkeQXWECxh2EEAqper9dCj
bIPZxBgHRVk668GON89if3TF+hycyg/p++5/9a7tMuWeGzpPez7ivGXbAyp8veKIq2dZvOsKykeA
jVUTHsi5hi27oBWNilgqHaWhtDvZOfxsO3KEf5IQVgt8ifX0l2K5/Kw1zqiY68ITVSSCV76w0DQ+
86hz3nxjejBVeMsdzncwM7YXk1vit/VUkz+AsHibYwKlb0Qa2PqbgXkZbaacvBc2qD14jYe5nee8
P/bUmruVqHXcEQol0bVum0iNHBh7lVzc/MjsD6Ho9u3daogzMJI66HNVaeb1SlZNG2mugSWXU+Ea
Y2GF4ylMM0vGM9E/Czvv80Ya7iolj3YEyDLA3PtFm69xXNe1p8VS5mXQbdGfj3ImETqOOMLcqgd+
keIx8XrGa3/zvstFNqAbqoMckU7VwiryiC8RF4vGgXthsKMSpOwI+kqDygQFmiq7/4ELxkt6TMUR
59be08LysA4La8nFvQ0kAOCUMIvhx79YOQwYa3Ql5uMek93qrkibgKYZDyDaZSTvbALOeMhSAU8g
G/jLHs8+ZLTvn1tTlh7ghVw7Ev7eCr/6X5P2CfrZPZwDrxaxBKJj6TiqghRsLZATe7iavEt+CTKK
vhAuQa9awPpkzJ2/hnK45ZcqKqmsO6hAkOIRdhnQHiPCa0rqDE3GHfp2aVoo0R/Q5Lm4+Cm2LFkA
w5t2QBhOLEAZLZ/ZQcLzyPdXjNLm46GB9/5dmFHAQ4FGDAqM46Af0YJ2irfIsOOpB7klC4QZSxYn
61ImrW5jpHZtRSeb0stWG/EHlW69PFThxA65bDx1/0deRHqglTcn5i0vebFpopK/7FmUcz7+C5uq
W9rqr3uWssD+Sp6+AlCZXT6bCPXK5NDAAsoLl/GbYslaSSjjuRGhgWojt7ouyyOHwv1QjaVo52qg
0dce+obUNncyxhMwTDTqNSqhjCKz58wSyafSxjbR30Sz2Ii3HeBFgxoKg9Cze9G3tnokwM+cKwWB
73qSqasw+isnrQq7tRTdR8xz5iGDnXKNAp5U4Ca5pzslqiop8+XcZx1tz6uLBpDP3RSgXqYogZJ2
YsUP+N1Rb+Kxqb23o/CQlKSe+K3PdrwJCWbzI+lUokribUfE0PyY9vFcKKVktkyrDj4V9Op/W1vs
MmCh0OihNdE2D7QtHpfEgei7oN949erGWz062AcncZrpvvwA1rO0QqnvN9r5Z/b0kMuFbzWKBfhS
0f6I5Jc52AfaDNRqBnMhn19j+0dQtMy+nEeFBw2gmh6/uxpd1O72YFwRATXvhb2gva4te5uYC8MD
+UQ/GQfzkAPSUkxsHokCqWzoxi3QMy5fnWdfm0cRdm5cyPFfVcvCP79M13jeQTIfJrBiymAHKlCW
lcw+/zRP5NnVkeWzKxJSvIpFSxU7ugkRKyNL7byqqsCnY6jChq8kpTGxC+yczDO3iAwRnrmr/389
EUA81wNH5N1o28rT8hdA1/eRzDvQAN8miKPzdE4D6SOKROHh0sa8gCqZPV81nuKRXK6yGXCfszMz
cg08aplM+igBCjAMF5fBAr5pta0jUjUXdpFOagdErON1xl+ltaWUY+dyRTc6OLGyrnsdLye4rZzN
2N5d0+jv3hE3Ck+mfB7Zl4wLWSA076AzzPfF9eKv7u7Vv2ZYKtTwoeWVOXUfriVpzQJaYZq/Aw76
rsDjv9apcDCxpHXREE8J24lY5EIurgopYtoh5MbtmBGY4Tli7HPEED2eN1dibsraOS48+cqeau0h
UgskHf2Y/bFyMe82Xk48zdLNKoEpzhY+cRZKG4iwV2Rc15JoCUGUCzcQfUHOdJRPZQqVnJQlqzo5
b2S3beC6l5XKwUS3TPO866uhBfPZ+jWpJaJIuoUTKjYCE/4qP+mPzxrMTt8reUZ45c19psNYDLMf
KzQzSpMCZlTl7NnqQ0h9v9eH7H7SslZLL3yqJ+ZodEe8dSuH/Bg4ZP8mO2GG+iqalfDTbrXMRe/s
M0OwSFcS1kFNNTJSFymD08q2iFwkRP6KQRUxg3itx03xeFJPvns0ZysMR4h1wlX1DkBLWhCI6Uei
2BkmsH6OQC6fZk5ODrg/xXv+7kP7J3ZyTynObfoA6jIP7i55Tl72ySuW2e1AOx2YWjaNK6B6zgqO
my7t5BNjG5hEsrJw5Z49dDUcUN1dCyLxalHhfVOepUqsnzrgtTv679fUAyPCgpwte81fx5GGAinb
JVwIb63WTQdGMu2V/iRCiRIZMt5A4uzHgcV4LeKiS0whwD1Z+0hE7MFl04wWmjjAEtKBWFTAu7Me
rNNgK3GlIZ5zt6Ayr/J40/aheaLbqJD+cSeEwINDSkOyR9HOaDaZvQO4odO6td4hpB5dKnjvVJJm
Mhi1JxjdBzT+PXjvnDRfa2MgMGXixMgxsBoWezSw1IEeakx429gO4K/rVA6xBfLwoFYLUmRG3z53
iLIk4UsXle40m/sq3iFJhPSI/hE+Cti+Eok0qMiVJrSuW8+d9rgGKPMnreyO9JdGlFNMRAbW9tXZ
D9G6lwYf1ZyXAySGI99WvkqzzZfyg8FovWbfsflFBG5YVA1aYq+qD4/Sj21VyMa8LNcRcCe+2e9n
vkE+h+xzzTazB2W1TYMJ9qYCLKDXLDNuh5YNbeh+XPsL0RsZo45t67wfmAx7HilXr2Oj6i00QeiJ
e6I3Vazd61orvqvObwhel5mg9T0ZLo5ae9tB3cdHxD+8mYT5neHRklXguM2fuWbcmudTzuLaN68o
sL8GvzsGsVCnistfgf6aBXK8q/rc8D9nPa3wHLb2CURHQDH2vzsqspic1T+hgL3o43pwriX8RLbn
t6SKsgxEMrqdbnlQBwnT2sZBatAhOJkUsnSG7PO76WgMO2ujmDDhmq33w6l+CC9UO/hoQA9J7uD5
iZITtDbSEPlaXvX130j1kfANROg9DBFdHHwB5WYkfN7O1IY3M76GZZ2iVD3bcwf7Ro56hEKiamNF
Secfg94gkhiT9kZC7Bq4XqY4tX3eWPBdO8JXdPUMuqxbgcg6TOfYYUfjPe0tfFwgmiCfoOJcBJCt
ZhCisQsiZl7SIvy4QWc/9YVLqe1dgCSduezu4vO8OJuOKs9dXiY4kNybQfFwZbc10Bpi13cxKMzp
qF1gG0fl44HA8xmuIvGgQ8pTLC0TpAaGPA5TBiSXKFFIUFTb1YZ00fgOoqGLezZpQa1nW8DXIH+X
OveWn4JenDfzdRlZ+3iqF1bvxDu2Uzs6E/22dYS3B31GB1KbuDWgm3nZR0hHGNaaA1O/lsyJ4Jif
SJvxUYVQdmvatKQ1BXhtmjy6FwUhlMU2sbuGVpVb+no7wRF0Obuk3kPiPjbKLQ6rTKhIGT6vrtJ5
VYQraCZuO7Dh5dXwEPXmKoSyzSWQLQV5NOyaLPjO8rongSbNdeVQcN3z6aeXczezEQF1pSYgFSGE
22Lr+1ZtiDm3Jh9TNe5YgcT17BZLxNqhFlyyuqjmN4EuwrpnenHm6fU/iml9mnFd/37+a8M8ft6y
NasjVYmuFbvj7B2l6CD56Dlw6yAq9pe8nxLzUe6+6sRfkn4vyQaRqzbiQ0ymtrtWzb1did0PYl/V
/ojdRc8SbXYthAs7hJ9RkD9XQzofIgxo8aH8wnviITV1n57KwLtuvwzEcS1xrE7vE1LfvOT6kD51
pJZJUkOVCZlYmKuFKkOqxCxD1wuaeW+jTGoqwbkbfpjuuAo5cio1sHhVeEpK413p9PkW/rM6O0PK
EHKkCzCMAqfBbIpptgtPde+ugB3qBD4oW0hDzwMLEd6lWJ4z56Esx2NkqTdl30I8PYch00tXI3S1
qaCGbeMcUcwis8m4XjiofiSLBjW0kyuFBlc8kpyaUlCgKBiS2SvcMrHCAfAIQ2JMn6kW3oubJv92
IHu4QrKWt+lN79psJpzI9E57GlF2LGzksqU4/KuRXeMcOha/N604XyoC+wfKIQFbfqyXtXpBnMP6
ihBw362B6/MnofqMb06bi0Sw4axAofhwYwaBFpcJ5TGlu53w9QVK5gqE9I1iXcBp0/e+SvWtu3ov
SdODmbFuIVXVcIRSrnWDlrcuLW73OQClmZbDUUjfauw8GoTmgSPfMncL8KxMlD/tMmX2FofioPMC
wepvDO1UNUJmENIy0J8hr6c6DTVBf4EjTX6rkpuWoX+iuwbVV+4+Iecx0iZThMeAO1B+pteFG3et
Bx//gyzX48u05gIDit7wwhPtSEAuO8dB8XciilgX579lBRq8W/13WKVa3IzuItlV4V4BhKDZp+M9
2ATvpRF7DnXyd2Mx0RCJKh2/QKw7tJXC+F6Z6HMAvrPVUVFoRUX7tenF70cUjo8aBLbXrFWJOCK2
yuQgOUIIE1/n/qFZRadMwADPIP04sNr8BFscBivP4m1k3tVt4GjIqr8FxPxsyd3hhyhYxTQv+RJE
XG7e39LBFDS12pWYF7JQssQcFFM20rw5kNDcevWNTs+kG9ZW1eBtNB75OJh2rY/hXyoWwKgx9Y7W
1/ntn2qJAFTmptV3X2M1VQe4K49zGRzbyhiCY414S4MKHlNp6LsS8BnaZyVEfCbm+8QhnG54UxHN
hk1/WkqcGSzBtoirNlDg6m2gQ+bFq8VpuLQuQvipzAlQdUeW8/u5W4XVPzx19S1ow6ckgQl8veTO
pByIQIUaPv2X5yU4p7cXTqAd6s1jH/IGVABBEn+vVz61nvkRAc++KyaPx1Ts9LxsjLxJt3rUxqi3
VnMrSHlTJ26P6P+xURrMVE4l7qNC9R+ijZPHkORgeuyDAe/Umixn1rFiWNKr9EbugtweM4+kFS5N
OtO+du1NiqUiuNI+sK5+Rvivdtu8s1UFzRkSBB7BRuj/kG3QO9LwtN1DbwcUKFzD90hch+uMTjhW
YiRXVPSAX6ZlPsFRhrrzOZS3e0kKoYdTFTDriar1kYWrjlN3SEMDqeaosFCmrLBV2j4mL5K0UMfK
GU0WSTlp4JZL2bKzgt1beuxS7kSJr5QJglRndglOVrl2j6VGdI4HrXF3jrMKcHSFMDkUuxzZufqe
wwZ0NTRujKAxhhwpXBn43kgmpz9Tp1/VnLnRe9GCM59PMj8ddvQzvu31/IVe6uHOV3iPVZwdWn4m
Qp75A6+p+XAYPfbGyCp4UYeo6UH04QaFLJbayI5Jf39gIwJqeeuCM29EcgVmXRLhIQDbc0E0Y9ct
N8hrQvB2qN9BUfvtrzamwu32vlFwuDVtB9jHG/RT4EkJdevDX/j7jsPenRkPpGK/aNmBNWEaQodl
/1R5tw5EDhim3InvPCDylEMR4QCmvJ13zvO5loRoIgYImJU86njhsrDqCgsjXjSfR5HPPF+TKk+R
22QnvsDaZJwpo85+XSzlgBO4ykyRkjVmqDhSj4258h9zksHlTNlJdt8VKx66RYpMcmGAx54rUGGM
AzV5wuqCxhc6Zg/CzD4R4AsEDPzDkV2y6hlcngCwURNed8UwMWqDv/AqjddFEqgjxC6wye4cH/xp
ArVInKM6gzHlb5ygYLwziZgBZCiYKAR6BwkBadstp+Duy6thpgphjVxmYuzNikU9ogd39bpnu9Ws
ee3FVYns0AsKf7XXiYH5W36BcAD5P5re1cM0I5X81Bqwe6c7WSkx/PATagNI/szG+7gqtRVj4yre
G2JnSwmJxGREFyr1tpTJdOAERZO94qBtEKvM0K5UPZLTDCVQFOWNRAZH2KXrokCT5fm/4pfksYiu
H/vuZOz89Itre4wAHPehFzCKH6AqxQX7NVW7IZeBt984kISe74bZmwEt9cqZRQ593TnBxVjK30OJ
E2oyVXaP9wl98jiiX9JNEstMeTGmRTcX3uo+Y9qTg2HrIrDmKJEMQLzNQDO1QHIxGGUcb2649TMx
QDofpbuVx5L2dT6AVdo+BbiM6RZQF2Yn4ivVdZFtEk4RdaQFFReUuztakk5I8122UMU44AmuVcnJ
3g6NoyeHxGLXvkshYFV6uTWEjmWbhcIbb3c2h6q/AlcQqBMLMkOeviYKNRPBanDMqff8snC6+mbq
bXYnWQStYCKtq8aTlqQIdZxfMk3gLGTaoyYyHSfMA9WtsxFrOS+H0vsqQiW5GiDzqL038UIYZvBd
u9+P1vGKWi9YQ6qrh7l+Dos+f/XVfbg4J5PJrS2oxShwpUSRNSlKjXUQR8C2JcAQc+Tloi28gKyj
2C3Wc5/OeAx7jXjv9kWU/btqwBE82KXPdRGxs6vokUUdksTA2ZKfEGCg168L74Or5vFZgmGBWfX/
tBfUiUY2wAVvUKqJgWtIUyKH9U/19ZW3F+0VsFLbMldbaGf6B8IqJc7cn2SOug+bJRjiTw6QW0zd
Abq+559hMhH9b5cuC5ZMLEyKl9GfQgiYck112jkrqFBD702fntwjOuLJ2WS47JUH4tv79Gv0PMUy
GDfWRc7RyDExs413quOe6mom0qzqZ+TuIjxnUzOEUiGCKz2hvBoUJjmpmE2oIGTCSIgxbRvUWNL3
FOZLvjglf0OoVXnfgranKha6GMzXqt/9+1SfKDCIT+T/NVdbqXvBSsTgebXdVKBz9DmfG4bLvxZf
0bfZIgkw+EsvoPUG8Ks1yZUp5NmgoR0wuG01G9ihCO1mFYJAIOARa6UuC+0dczW12Z9s1tGoKSDX
YPz6Ke8LrsTpP/cPesd0qnt/6UpGCWIks2zeEW3Qz14PfbdSzVMGwkXtDkO1LncyBxx/cshCaRyC
7dPvCpZtSj6nBrpXHUgueOSunWXvdrmgYoA2uphYq9s6ke9/zhdLO/TEAgHGOMsLS0PiqmgzJm7f
Ktt9PgvXutjkjo49AYbxMX0wM5TRv+v7wJAwjlZBfE8ogl6ks5cHlpJX+Cx98qo+k3Gr7IswDpe4
e7GxBJe7x/Oa/rKbZdYtQc/EqccBdUWqLde51TmeeJvoVwaJPF9X1Gk5Fm7F8K5TSW4AfPn2JEuz
JCJSL5E5rDzX8+qKcswD+H+cl9dd7cu3LdI3hen9BIX1+xIXBmT40XIakKc0Ae3SXH1dfqXKpzhC
aFMf3AdUOUUt6s/UoB/NwMMlUNVBIPhOXT5YurL0yBv5GpXW5xuJ9VH50acUcN3qO9h0wUpil0Ye
pcb2olN9JslDnHEFtbqSTRl7ycEsqhGx1/eRlFGx/rEv8KHRBLovl5guinee6EhbF5/XIw7tWiDO
BVfrQz+wzzHaoA4F9rvSZHW5SoFdJSIq2aKvWlfGzwt60td9TZyh6eu5Cpp2LPpNW2sa/IJfjG9H
aQFKLMSlgod6+8/wmdFN1UQFxLKJy/CleC9t9liZ/Hx6FWZehbbRoqZIIiL/U1LNuIeCcDUGECgL
ioDrM0hd3PzJeLxlqsdKV8COe9U2ABNeCO4D0Rwtq4cJhvJtYb5CNw/rTVbquvrUV6P39gzioUjh
wEDtz19r41oGEmZRstdA063anjS10TFZlyLgmFw5GqMmCmkiuy7CDuHAzxvWu9/8w6hnG3iskNxK
7DhnH+t0USRVNsFhxijsoV3qZht2un01Y2rn+Z5VeyfIJzfIIlMiSj8toEIYVMvJYA7eXwTDx4tG
h5gH4wbtcqxapgzGVjwBRH3BANgLXYJEmZzWc1xiAC9Chop1HItkd9HNPEr0RpeYqqA5Ixz0yXo3
eGv+hGl2e6y4JU9Anai1SXL+OAXrIpuVplfnGt/rC0DEo9lgkr+69V4F9Y0CKQ58Cb5X1UobrhUk
9qdepvH9M44+GXe7DO4r9+itbZtu1RTWrNKy1cJTk3G4cdPVjTQnqlD7ny2/Ba/HLyXJGRHDZugO
PpsaRDHR9Qg1+Xtoe4G8PMjhRKFAGRbUWKQh/hRk4hDYFq1AYoeymvUNUGPYOD31FC/EcrlqhE7l
esC+uLzaKT//V0d+GrtRgSuAtKbR7EouLybHMrpN5vySrjcs+yPDEJ5Gj8H6h8K2XeKvmJUWot2g
t1gwhnngM+zgH9sAXvk1VdSlTTYRfkalCSR90XHe6lr3Okh1lPAJNqY/6Osbvl9i+PfnpTSNXqqC
08MI1epbIZBkwPNBGlZHsoCxIeAypLLlNwUJwcoF8Qa3dZz/w0532ZPB8YAroaYGnb1ipyG0Dubw
xLr+6riCIrZGXwo8RBftoQVS2bfR5cA9hGzNAA+vT9T0mTPqYQK0szGkbJT9mQIJbMjftvYIcSyv
ISDu+dgEeH3TtcFJ879GiNabx0aKcmevJtx8C+dx/Og3fItGcQWvopyTq1/FD2L/4zOHM6Wj84DZ
l3b/XeFVtfQuMVQuyxKxh6rKIwDQWIlOVm0dJDa2qNLT/AGZU7vv6PuHJQx18IoK9u1p9aRB24zq
Yb94947wmWHT+MsTRn6mp2YlJYAqSut3zG/jxUGVo8sgMxFdlo0h8Xth7y38atR6WQa9GMyOz4zs
MfgUdTTM7hBK5l2DKZgJCl9R5x05gDvRZVFyJwQHTlVOblNSzHIJnl7J2/f+qmDuiqOBgDG5FYmY
djtSDed5cNSzTW/EiiSH7pYLsB4HNd2qInpQlVLz/QMvT2uXgvozYeqsoGsYrBrL9uluvr2BNl5/
i765CSNpcxBgfEJGxj+gd64a0SW/vdptu/WfW9gvtYc5r6MAVDGHE3dWsslRp1c95xpY7l/Ub7nF
j15XMF+QK1Sj16eBn1xL+d5m9ArOmZCgsP0SrTHxVu9f34GomBR65CyqHF2CQJv7UQHHg0XQ1ETM
YMVIQn08JPN8CBB0w6IEInNjjkPjzKA8IjzqgQ5TqbNW8wE+YHzoFSRqw83LbKdfks1guJRK7hef
XyiazmHrmu4BfA9+ffw/DRpiGBQLKsN3THyvIidRyliAfzAegS+LvuqZ/Wmhy4WGKixJXUc0VLMN
zlXuoh9HIdKQqG446RxGF4KNZoh+ytoDJYt8V0f+Avjy+Qdm1NTeJ896y5TUutqGfvb3B2BNsMJ8
uZz7SxzA9WVt0TBJ5l36FqI3DBUVCcJyTKhn3r3kfCWqX3xCEVlkDE1pwDSGXHnKgqoySzVdoD2y
Swu16Jo2HzvOaVX3u2Dza9E/bH5DBrl6PSBDVPnvr95Z8PQeKXvlikDCgaCmIF+UeQdiHa8MzQi9
Vlc2LXVr7J4bksc56uDSDpG3jzZxnIR4VCq+YotT6HO1Nt+I2ALPa5jiHXtLG2A3T0J8u5MLau9h
uZB7YXb9aWCs76VhKYSIvE9GQhCLZrh2qtwWSjqwv2+zbHTh++Osz2EYTabs3wIo3AcZKexhf7mE
8HAbwRRQrsr4NzFjnFG4ThJJR8z528YY8/Sm9AJvRxvVggxROOk2fwZKeeluG3ew+CeiClvx/mOj
FBPSuld9wtAEPiehdKlNjIwGxgkYBtKlEn4mCzhzUngY7fhDDAn5p/HuypZy1+JqXu7RAN+HRQ3t
luxKoMkXBZHBtS3kOrcXHSXcCh71wWTJtfkE5UiDic6pG5+uafjFry9d9xmgWezFY+eTXx88+Iof
nIB0qUJP1cegnkHjzvEdAh9BzwR9eaWv5ln++k5AQYvTp3lH6hEHG8etpjbGWlRJMFyYpZyiNDre
RFN3uFLhgz/yH1zBSR8jXhd98MOsjIeudqcdKBdBItUz/Mi0/wnZ6fTdpcFo27WfnqE5nkq/K1SE
iNSFaE9s67CTIwgtaP6otSqwQaq5DaBOaaI+9ignDm4wN2elq7cP0yQx/D1GduQsX0XjJbYkqGLW
r9mDH4uaYGDhZw5NV/D4oraKuT4GhZF7HLISPe17NSgmdhX3WkX4mAyP0/U4vzNtGA99QaF3B0P7
Xc+pg+vZnbE8TytYryN9jOPIUwOokIOZxQrvw3GVvDCqBsn5Rn0sP5yuxPBPDDu1O/3Gb1uqgOI2
XBulZuu7+WUSI5Rj5Ipnqp3F0htLWtgLs7xHbP4Hw5cwvj2ik996RrZjpUd9NDsYO+3e/M2QgG2U
I6wPjl66jyWcGc1tstMkVobsbzR1skgnGX5s8yw5F9JfAWjRg1ewFINBwjLlVDo1mIs9ZGD2lkMg
J6jSn9jAkQ2iSVfrDHFwx4V60JZeys6GD0//PvVgDnqPQn1DtZUFX8yFAWyc1tLS2hmEUEbLqtMX
6m9tI6mC49fPk1TzRXBSR2w61oZd8KpsWwyzAeW7oft1tz5op4H6DL8qKQ30l5WHB708sUjvwkGE
f9gh8Aeg8dd92QVm6dr1XDnYwutNqvLUDupyOrxpf9ounO/T3MASoqPJAdzTCQYRjOcHHf21ee9u
YcX5utudBdk5JGiKYqCqq/bksfWJo7UDb8x+f5NoGcr4i0HNHZocIzHSzAEMcBmQLNHl9ViGDzHG
894D0l2b7itdt6Wob8Umh6DpZR47b7zeNIJEizIhScV7XbWUF6WeAWHcflQapNBFwmMu7pQdvqwf
KPRBN5VvxLXZofGEoMOQ4iqyRMcFFf5BWfNkclJ3l4F4QEyHcDzncIEtq9WuEg4bWFWEXgIejaoq
vN+4gvMaMRt764vG03am2TNYYlcqvjYNKADVa1zpeBmRCZze6oI8ImCfkQvLw5UtZXmrc2c71obg
ZW2Dqt92YUquReTNIBKwGwHs+N9BF1nmRaXQgtuE6/5Uh71aAOcftfZMZyh7aXnORfx9vMNP1C9x
nzUJBWkiNK0Y5SNkrsffWaPpiK8PHdn8AKkWxF0nb4j+yUwaxoJO7TxTlLXCCxDycjos9vULBIDu
PP48L2pSsb9sDjLtq/bkCs/HgB8rnv0hAtPd7iHMQ+RSzsfba6zwFWgTYMpjHXQlb6bVD6f2VQ9Q
lZxg2unt4Ucs6stLetePkt96TonB+gCrnXklz9smWSlWSh2RDgpYTNR7h5FTMVRdal7S0yEimIDV
ZpjQ5tXgs62naWgzgXFrNKD05fO7IaonyShFP1xannw71hRfXYZc3wYNDqU7jyveSDKLJltB+wIX
S6P6EY5hjikdq5c2WS9lKefl6hqKcNrCdiE7HxSwrplNZZ0xmyHJqPhRUW3lPt01MZ1lIDNzo9EE
5nLuhmqQwFyuzDSjodpYoTpYgYSoRGFksAQDBqPgKP2Fhe5qMwmrHYjGpYQR4cBfMPSsMXFcFha/
Td20vJQNGonDHG45mgSJc9/x8LUdlGLGKbzfcUezQFzjT7WqEkfPTZnAWypdYwB0NP9g4sGNAJo5
sjNMPsIf9rqZWXP5xWo++0RQXZ4KSVCy9xsP0x/sbpdOwtJ/Ijf6ONPFMnq8K2mYf9dCz1Wlc3sc
68UX+SqEy5dQP6zJBblJC/gwvw0Pgl5aXEH3LLdc3Z+EVbjzl/7nZeg6GK14f3zC9GHJdp6aUilQ
ew6RTDjPonO5nDfC8YlO2TUgrdXfrgVYNyrxUQS1A/UsQ7JWyPcxBP9Ll6/eGJL73IakeUOilptG
kooAOIrgQFBfCuk9TANayHK9WT0zmpiIvKyw5GfpgNZvx6Gjn2poDrTFOJVwLO6t/xC+IhQk4y/h
kCx5muFK5sOA6Wq4wbNFLfYcE7bOLiHYbIravTivWaSQFZijeIRqvECarynR4PGOGhJVxvYYPA+C
xyOY7UdIDqCOigklcktqnG3BdB8+lXxgepkdqjLe1dPVr2zA517XXZJK1p9lielZlm0nnDaS6P4s
3Do6CWlSIQRlgJHuJqr/3ji0IIDGJrykbmoj+wf0EojvOxKJV8JgGIEyMYG5XSRfk/APn05URseC
PomJbrxwA2ec+mIsLnhfYGKoFy+Da3Uy6ysN8/46Ww74MgZ7RKWQwf4GNqJQZbaqmc0Ub7+wXNyq
PD1Co/nulifmH4T6hud0PXCaM7ZtalwfDv63Lv+w3Amz8e1HC2RrLHb67qSLUNVj2fNmr618TVY4
vSNuELoy8YlKhzXlmvAm3wlFmk7fPtMFXKhbbqT3bpsb0OrEdSX+1WOZ6VkS9c7XMuyp9P2v9Gdy
KgPpKNPvmfvgo3X4JAnwYUp8qmMQpjeWPxDu0c+l51LHl1LnGNRh+hggmH0fwrhZNXa5d9V5Kv8Q
Xxjzck6eKFnDSo/3eWw0VFb2PwAqb/vyndW5FGOfiyRefTIoeyfIBURDAtNrsyBUQZzqtcvQtTZz
2jJd5Hkep2R6owc9rmy5u7ZNh7miNQVtpT5wmXpcuvXL8b8HNF4Aq3p4J+HFC/6xK0XJhI8iYgFl
U44foc6NA1W9J6/cUvA6MTk6DtjLRXrSsJN6VkI0SWRXhEWLsGIbm/4ZxKlqaLkGWYVqDNoqvJn3
9iUffzjEKcjiFvxM8YXHwlypC5yKaNSCJfMmRJ0sq7JYkUtYxMk9DoVHfoRA60UOuYVffZem9IYo
SlRiWAiRVyvz8CB0iKtYVOiMbSUt4WAA1FKoRWuutH/fHYjIt7+nTidvkbNBLp1x/K+kopw/f6aL
Rn7l1jE+RyUF8rcQtZcBATf3wtBw6idWDUzAsCpGjm7fCGqBK6DiHpiZIBl2zsELbpN+ur3AJTLD
Ww0ucZnqRtpTtnqlUstZOTfHTnm26UwCBesRM3pPg1rREmgqsS9VnW+V2lf1RK0cuojtCVvlXagI
/Mz9Uqz5p8NaYgkny4yxqX9l2fyQzIclwZmLIAzW/bJ66KSIS8IzdTf21V9cBY4YkdUcqrqg7unH
bCt5gGzrI7cCpNKah5KionJ1iIddQpO31I51Ia/kvVP7MNtZJR6v30zvbd0Jql5m+XZVEia73Vdm
cOLO4N/lTeKuxB7ChoMRRs26LcvgcDJ0Z0k7ZOEdT9DSzO/myZSRFJ3gZtzAbDPCLADkEqrpKsnl
fqG+ajFUgzb/pwuAIz88u3R8PgROB2iJVEc0eGVmpjOiEuI3wFVaquzJNsTisOhCp5G+A7abNCfN
SvrW1pDrp1KkELvx0AnVvLWQR9L/989bmrnxIvZaGowPtYiyQSM4c9mkSbb5ZeVlFhJNoYdExTEa
5gIJVaF8R6tbQWNz37g+3YwYY1pHjm+A6YHuwG75I0fQLsH+7lNlYIVHPhbdGCRpFDXP87P1hliL
jIrEVdOJPd4EV1zuTWU5lVlJuOVhLYaD2zQu7BNDPBdmah22DJ+fs4WghAf34dwkM57A97YCgfr9
mOGWllXOm1vmuf6snWkxpFVDWLQdYOmGK5BQ2u4lvHxOsLda8cyscJUMN1igqMYyITCly6jZ2LAs
3asHUv6W/0a9YeFHfATDvuwsb3jGCclppKkAwGNaPHZppTG8iv/m5f3wbyJjvY7bdGGDsVuxuDVe
7KmFZLik+Y6Z+iRpyA7ZTkrvD6qH3P6bpm3ql6UJBF/ctHpFAra6j4PcNK88Su63UwHaDcRcnrcj
Ha7vS/b/DgdC93o21egpD6tDUI3OwCeQMMIulOAj15EzpvRlkQHVHq/hScrO4Y6cNHuJhD5OHMDY
93nFyqtYGF6H0du7/9K9U8x2+SqD4FxyzT2AixyKMBisshtNMGEIxNTQEQBj9mFy7pqkgfGsflUz
Kw6Q6n76UDb+gzdvBr+lkjBm9ryjhNZA3FWMt9/DTQdGHNzHTYg0Wsayi3WdA7Ap+eXZaXYxNaAX
miHs388TgADhCxkyqUk8D7bkKMrX3iFC4stt9wCEaPVMi5uXhheSaFmG/rICwF2PvWDkdU13O1V7
BJbbsxcLyl9XicalAi/ZueszCNQUYvwy5bwBvDus1pXXEslhTMEeblsuxGHBSCTRyIEmX0nbro2f
QY+FJPCthVomDoG+dg4r9IZ7B4r5zbtf8uMfQb9GkdCDcxtwvLuCCzTjVhAT/sY5e3OKrN4hcO/2
DdspkMVgFuFn6oFlT85M/XgMfsfHP60QJ+8hCtczuG/g8be0iXTYCuizjJBrMrYT1Ia+9j859l18
U9U5vstEr2VmzS/+aAq/6mIACxuQhZlqkCgtNVMPQPiKUkne5MPcS3zyGpHovo7dLonyLD+mcErt
QQWMUhrBcaTyLajhqDekX8LIIUtOG5PuG05rad98nrgTM5/Jtdzrj0ZT9uMQUmL/vsGb7Nvy653A
vk+/AjDyVq2E9mPL0R6PJ8H/VJsCG8Jk+1fJsUkl2+tkNSm4X1XzS0nqKEebSvF0IYw10QxOq+eF
N+TxrAjPuWmXDUjbjlNiALcZm/e+gcYne40DDDK68hIMDtsZWiTMW+aVBUnRpH1u9LpGPFRZWX4g
MJHze4OrT99g4zMMVlBzob03Jj4EfzvXXdHKOAf5+XfAxP+xD0pim8V3CzSu9u6vjJvTWRNCaCP/
ceBZK4EILHJh8TMy9nl/sGh69LtOpxQIb0jgMYcCpEXnXK8unR6libQzr+yEfg81j8DjFGIQrFuv
TUZhLp5KwuCyP0K1cJSr3ZqUxG03ziX51hEy4HvDH+DaC8h4lAztQR9ArgPGtNrdC9HB+B0e7+gN
wRqHNQrs7ZwPAjpcb9ewyfvBvLaI/qQgck4cAyOSikDYBrVVL+SzpN0uDAz1t8965f6ScZQkTK+L
8TqfxpaV4604OV6nYRl3yHq+x+wzISatJBTzoci5wEPAhx2AZf7l4TPyHSyyJ9mRPw0yy6eSJz0Q
dG9l0XqYZdzXux4DlpWO8PZLdE7NExNHoXS3aAa5QjbR/5jH2G5ht3cZTxHghtsRTmR9Ry3VWbsh
iOCKqGL9XfzMUDIuUHFenNBa3GbDBNKqzxx9eb19bCxCbyr0h3UdC2PgCrlCg7sGs4oMwYKao62M
CDzLEEELAGpyPFco1b5h/jpmgJEZgIKZzGJXnQeQoZHhmjAApNrVVPHIc/KfUznSFkQw3Hj6960W
rctj9kagSKKBffvTYBNflmnaZknwFvBz9ajGoZO1q8M6M3THYybEN3yigKnADVK4GDwXZCDMzgDW
qJwsaWdmvXYPlfTqnyl2HP0if6axy4870kAlEOhkVO20cocrCuat5Tp53B2n36KQQiwGnfEcBznH
ULw/iwUyEWpLRzbo638fZoyrxIiPnbKqUsXqMom0ukH0XUjieNJEkCJi2Emrdx01IXUzwwNyg8qK
5ZhMzLcsfKaAlbG4IBKmoEcL3t2ECoVQZIUt0WHiT4ZKzawt/C6B0TcsGcjYA0bu8P5LsYosIoVr
m+i2MbDU5B2rYEhZDOuXTupofp9U/sjLscywCEFSv9ySO7En7j/WVi2nhCx2Qepj+I6qYzpUx4gD
2hatv3evJdhE8WzPcWDUTBhWczY9U9OuSKYzj3HwZHml8GSxmnYCJg6N5bnqtjM9CtjouQIbmfqD
o1jU9C3vlqNlAYRmOvWhsQ0mg/7EqH7MIwfdI4okyVH5s4JLtYjwLw3yixaBmKNiIIUqL3c9HMRf
fWFOYLZw1k8cjljx/5DBB65HdgReh3hYdBXI2Y735n2lNZ8CVcDeqJFmv3nnBIoaLuV7SabP5rFT
TBf3K7PpOrJs0UEslBXoyP4Gh8eYborjOLTjWn/9d/w7jV/QX3zQnvjjYyr0UIiLYEzOzteLzPye
MGPuLk36mJerwOZO0e3PGHDltA1wr1Jnbxxb2QUU6ac0p4vnSuTT3luzF95c84OpnOV/xSA/m0YN
9aZMH160FFQdVv/Oex8aa7XskhNeGS9UYYlKxLZXuMTM7t5u1dfU3eZpDMMRpUdFUiwfJrhP0ogL
3GLLHESdkhH69KtVxBhASz9sTS97z5r72tn9eS4pmlXi7wvx5dy05k2r6iSlnyUcPL/rYAtJ3s7g
iCgYmkgcW60O1yrT557mozg4/m2IWlHNb0+VsIBuhB6NJx+6Phl3Uae3T1E8YEnNTt2MkhEXrke/
mb6qGS/RrxI/X8Tvk+IClNu6X1cJhP0L+y5qTUDErnWGUb+GFpvgUiRS+1TVvgFzrO0DP9SmZyLq
N9E2ohmRNMj5QkxVBeks2gZeyTzDIn8nSJPwD3DDvKI7iwiAcwZtpeWyMkz+6vObG3cHyIxGm/7K
iuHxzVrjI7ZFVMA9IGwGkUwYVTzvhJlaxI4R8EZVGniwcDg3fHUsoREaxmQCJ8ek4ErTB5PvMXek
yTFMCPJ6NqWToRJyilC8imhqD4FEStRleeb9RaO3gmaj9t9Q/WDLDXp3WVW90i87+HS20xL6LN6h
sK1CaicrpZl0XTTPWVmq688VXyYOZdVXVaZH2k3rlSiQHHq8XTmZcVVc54PAarfAfErylvM8JN/+
cUxmnVl2eUqfViZfNmIllgU4WG5CwwDN0CAHxykNTG7/b4SIfcl96gCwAcugCR5+oofb0nPf0Ax9
+V4J0jICQ1uNTyDr4GkmiDAVz6Z4hGhYqHL7ThxH201bNPP2rejGVEMJk0tLHRWFdLAoqOgPQ4ZJ
I+fsgptGagp7YmKUnabaDRTMBr93bq3smH+BF4C/Dp8bfqVDHlAzgfISeykoO3bOL4SVxWJS0WuH
53boM0g6iM+vXe0Y3fbG+37oXXoOFhAGnpESzxfEVZte5WJKlmQpl0j0xIDaP9xKy+aGmGpEz6Q/
6YtNpzvu07CMS/I3yvU6rUJxsVYi4kcauPdy0qGomCYiJfPEuIvAEzNyJvfby+l94YIhMhLq+GJE
k2WdI7ukiFgTRusO05tHUg2nwW9/Sv/jRuHDjg5fvXX8+CRasJ5MTj40cOdf7OQhhnk8c/y8bJ4F
lXnKOeWyc6Bs02n349WKSr8UxLbu6tBnArA8Wh/sgLrxt1nI6uSv/VWWMvtplS8+clsg+o05dqgB
PZdnrlBnEwK7E2eyukIRF93Jkyflc+DZSfW2uqAI2qnf18+oRHRavdydw9SgmOEzQvqpk4xgg0L2
mT8yTUhErgNGKrk247XVHEhUCIqZvmLnxXLJa8gPU8LUA3N/cn+OHC3cQnpC+8SDicYURwo73+oh
p9/HhsF2kZFPE6rsNYneNaPmZF4CqT3kBtHHyjlhdRqfOzTDZ4sbnFSItgGIcZtYmRs3ZaNjKaZe
Z9Tk1/hnxcMIPBaiR2bu/XP5LiEJH/ovHBr28nKDlb9dX9TilP4NZMEoxUnBoFCNiFIi2PwjoFrU
1eBsImy71YDVllcUdrEgxgY1uuoIz4BKUR1+OKk1lC1QF9z4DAYfBZ84WTb82giynn0hYoZKzaWg
4BX1+7WiYIm7w4cZtSkNgZ0eYEkW4ZVeh2P9xdzM8RV5l8bsaiU4nZ1U36iZgZuVhN1pSe848zcJ
KFqzBLvEST2bM00v3pSdAxl1noekBQTTzdIYDjHTIqxp90FPnc871QsmK7axIGnzhJAEO8cmNsHy
BZZtQr1buZZszt+mx2RMvT+DbztQYfa5yEg0wxoINFdNvybq8a5Gg5fXB/m4oknt6WM7DFXxYKVv
i+iCYfuYCT/e58tPHaYmxYWWhV4GNMwWF4yV0o+oJF9rNorcxhs5xZYU1viYl4sOb0PNKcA9f3Hr
IKfbDb/wiBuu+CxrqGDb1gDsMdECeZGkb7IRM2ijEAX6LaIGNpI7sNSk7UB67qeEiv4LiE/lkoFh
40MY8dP7sgiHikeM4nmki3wmxWrXMaoAtZiCdEia5khuH1GqxWEYYueu1A82f6bbVYi8ySi+z4DS
qSPUiNd7Pqhgr8bhtzPtyLNPlP1GwUYaVWhu0jTuvPotKj+lXmxSNsduB0VomsQp7Eq1pYgO5fbs
mRDTtn8SnyejKAFqvDmwuVd1Vg9r1Sld0rx0DMROeJHGKXfTvOcXqv3Lhb2eo2fM1JGwk6dHTCyv
WeX2WiYwduEXYIAsa8DfAqmZYJ5vryS3Twq+9FhI4iCyttoqtqgmjNDEMVA2/ugANPHFnu6oRwff
0LiaVS04x4tRgIJEAz4XzhJOefWsZuQU0rYmX/OtW3gAv5XHr0Zb79R4S57tH35xUVXwwfBPVwsH
SXQbqxrcBsdCAbjcsfU1yisRKegedRRWJV1cMHAei5CJx77I6lBQcQqo/jQpX3ba+Dn7qv+txy2y
64vubu+HQctaHURsuC0E9/AvCr+Ky+RD+QHMHOt80NH47eG4HRuPeQkcxa/tH43UZCaEc+s+ZXji
1saqGgOSswaAPiRztBneZL6337yIbzg6VPvsDmjaXZUH+YRsYxKuoC61g/tFbDyPrYzvPmd4PhBW
i3k+pFbl/NjIuHbfGlYFitNf6EHMb2J1HmImeXZdqvAgtdp2G+TzkD8Uk7OHKeSDd5451LLEeDrV
YMAOhymjv10Vs+Ima7tNQkPEZUao6FK8cqRhIzgwarqTeU4GnhYUZHRYf2fvQQaT7Ms4G9gj6qhR
u61PlG2H7+YxJExPxnFucqRwCzcCVLAHACMATfqJFgwDN5rPPU1LS3kK1rrmWEtlio4Rgb2aex1z
jriOkH2BYGTlGJxnQ/hYjYMmjbiGhcCngN790hysGkiUysZKmA1CplNlwOjCjc/b90PEN9mFZxV9
82g46Gdezkokgn+hoENbTXvwjLajOr0eWNwIkf48j45FPMiJRShISoXYbtH2sYo7fP6cIETYC8g7
XxJoSpQQH6+o/YiAYBRE521NmKt1dtHdN3bArmPd6CCPOYk30/LtlLl9wGbIxglKLygkEE2p8tFh
chPL3DysvGebMexqeVgiWkj8+Sc0AZKedPOfAdXzeOeDuqNmh06zi7NDsgcYZNDMS7UnBM8VAu6/
DiQQuzEPT/Bj64wJz9nBhEPOJvXEMAUyZ1DXrra6oJqzPW8focJkJdeV+tDQEXU/e2NABFGdxWzU
Gdam7RHV8JzaLQGefsdkZVAcJyq1M5fJ03mO4+GPfxWsFOZyAnbwsdmc6M+U3wOkiHBZxqIy5w3j
H3aYD5FAZiIMg0vjX7i4284thhCnF2mmXsvQUu7kOsrQNyvWj5MCKyJMBN6C8te/cP6BJiTHyxSV
228O514NFD6RcllXvtRcVhgEDRYQY+R9QOkKUyvZxOjca004VY0+wJc2PmZKk/YuD0Y3QmAtLr/9
O5DTmSk3+SU4hlQwLezbzLyyJxKUwNkxFMWIiVZD1lvVpKcaWv/nsRQFw75t7UKGm/02Cfvh+r0y
nE9O9jGxwpLePdkUAplwfV6uXeYURDLqOuUOFcpqjS1E44xjJncGReLSVF5tZUUr+ObnlsxFVY+D
yOc/fjakhiUJaUMZLwxePLh8DF/wx0Rcos3F4/T8TBQVOc9kkQ7W+VYDRt3IB00H9vV3okZ7NFpD
veJM9PROm+tg1u0uc5cCqiBOZfSfb2XrNOMc9BAK7VdyWzApHsXK6I112E6WkvLfyhU5CQWkQhl4
jnDE3HwzO41T883khpPT3li2QtKYvu30yBQeEzpvjZfBLRK8omcK9nXzNSguMz9JJM5oFykouI0a
QYuf7LiZeKwMR3D3QdxwR8l+ynA83XnDS47gd7R+AH4UkgQ84IxcX5hQUJEi+gqG7fY9OwZxeklZ
VAoMEOzcld6Lvrn4siECHmCTtQ/2c3DWEuPOsl0dV3t9Vr4kw1NFZPIJtr+7jkm2AEvlbhOpRAbb
0Fhp1lIQDJNyILEb3mYe4T9b6SvdCUc7bmnJoFRQTS30QYNCu55qWwNR58YqTitmp7+AiT+8bI2F
Xzk6oL05VsCcf/ZoyDb/cSja68CtLGoT8xxnPwtq++MfDsDNsbR6rwJUHCbfFzxVHoubyepiHxhg
gQsFtw6PGopMmWzWluehPI/HoGzu4PFfBEqraulJagjqzhA4zesIgkweikitgyjRVXf+9/cGsXrq
B4H7rjls2VvxHsqUN+l54P18DzfabZu6h2o+Os9ltNly8E4zHvnnTEpKepDiQcwUl9yEv1t/Lwy3
V7VUZz6OYSox8S240OWBtdlmEHePr7DKhDgJfVeFyGb97JcNnfMmktsz/49iogxwttfi5WX8Kf9N
zXzi2vC42/MEI8QzBjNAcmqSoTH7m67pTSsMTaVPcHUcNFIuYbsQI1gL56pKmxaYQ3LBSElSrYXE
gXMKhuWhFPfhNJsJpAN1i2WQi/ot8zm9OhF8cn8taTpb1dsUg8t12FucdbNvkVVdoXhuuqs7TIhd
nIn1i2eY6iPMuMhf49c6K4DEG6L+NEDLpK+YvTbz847JaaXC9zlC2SeC5R2NnKSCWr1w1BXtcrzE
2dzkKP708Wtro0kqf2+5lQ8kAUyL4VOJCIHWdZXlHUbvzL0PWY94TaSJYPYEJSDoIEenAmYNgyz5
j7hNxW2Cm8f5unvTyYaTwaID+e405rIShoIiNVJ4wYGMkVMZgKANhZY5s4BxcI2TJSOPZTiflRCM
oepnRPvvesqmG1axx6gjejEAbP483OjUZ/+wkqrGeo01zxRiEk5LGWPEzVHVfmJxeVXD6Tk4JDN7
PujoqQu68QzqCIP2lTd77U8moRuRISL03dbXgPgD0qrptwpvqO+wVIGuN8cl32RH05gb0GuQXDFR
38Y71tTGjHtmuSV7nDQgnyM8hghMzuhaIGMThQA0HUy5HkBtEk99at3wC/NKRqhO+nXCRgjJEalt
PETmXDYKR0DowKo33aEUEa6O12jh1f3GJUiSivF4jIRyerndv2HBRH6TZZRqxbhjG70iKwhJz5YQ
CnBKq+BCl9HsWv9pso4scMm9kOvUAlTXEAOwy7KCdh0chuTCdzZu+FqULLppZfzjXAqxhzf5AeX3
6iYY2p8Uo/PB1ttllZMhkatw3tbPENyzmDe6A603iOZ2EQHrMf3uaQ0pf+Sp9uRc1IPJPkash+YH
2YKHvwur0BKcRRzZ1vsErxq1WwLs/KD1nMx3vXWa78u14q/kdztHEekx8F57lnVTPku1kwVLqpz/
9h4nnVeq3HwAY3aUm5qxBkH3CH+ri1vGWOM4WoVZfxb7FxGo/aN8lmDHsdtFxOMJnjGbdMJngY0F
Td644+rn6OMYUpYQaIpUkd+yHOd4LhzQLUfN/ZlnWcjIlI05Eoc9EXYTmGrliLNcBKmCHDurGjvB
E00LLoXJcAil8v7/FVfV3Ub2r3H6ckEbyatPo9P9vAaDp1AmhiKf/FedQSazvQf5hV4MsVCCQ5qR
BGlvm/0/4F9VUQTkMk4HCXtLpcOxspYGGWVAH+PwVMB3FjoyRiTCLfuJGwlXSPYH/seTNNjlU88I
szbE0BILSior+2JBbP6ZwPmmcqkNLuAT9u8j7vfmSYwDNpfJAgcWXIb+k08HsiiIE7W0t3oNqBQ3
oVOyPkwYlqJ5Ds9KanE6oD6jUInwrJtoSb57WCFQ2eWsJcQYmcsGo0zgiMBVK/jm2ZnHBRMKO8I2
VpDutvEkUkCZlPiagT4fC2+XbPKlyWbSisyxDWg0BjKPK1DDmp90Pspb9bS6fRuzxtkOWRHq4eNQ
oxJagSf6GUSm6AjdEQf5jQc1JheVRjf5SRez6rB9j3xm5tmFeh7nMgdq5Bm9z6z5Y7WspHTJ+Qe8
d5Um3DY9kqICVXLPOdBah291PDJluLQWVpf8T3Mmn/01Cky9KLTQc8WHrljVXUXq5NlYQhgCHuAi
MBnUhtlQ/nP/fAnLgySU6l/YI0vVpvt+nfAyo+Npbb63RJTArZpeBLTQ/MRWOulsSd0Sgb93PVRw
9QFhOUnYOfADYXjXEj8trY0l0IOMqBm6rig7Z3Wg8Ev3svZL4Pf+Ttb1AoJmvlISOVsALJynpRFe
XYgo/wOsQmw9TjFBfEAdSWPh3r8IgkbwgEQqghlBdt8q+MtXyHpbFF++3CFLiQvpby1b/cIfY8qA
9LUrXEhKHPMVSMqmQbF7yeWfegZKN7Lh6o3EsTYY5X9ye4T3sXK4yguuJ8eCo4ljyTkV80Az3LWr
mWOr3e3gDet5ptdaj0rrXTfkSlhxipvqg2aSf51Vg+1eb+gjR8fgR9OmMzp5wRkb96gGhCetCl9u
eIA3Sf93UtEUEyCsVpWtyrcVrMGw1/FHnelWMLQgu/YVZApFfaFywTxR8Jc3KamBNh0Ekg0nEYeB
EEGNmEJxLER0TbhH8XSOToH4nU20X2uGDWIvv3jI8Kzxq0iSVO+KZ4HYSjqscQ7wf5prqvALDFTX
9Af27sF7R1E2M/c0wBrGu0NRTm5fDTW7sCYnMPtL+qFA/sws/sd+0kVouRp+yIn8aidTejCoDCmf
lVzTJuJY1b+aIBhIznPwxHFfwALCz5T3uKIp33HsAyFR0ri5/FTk6lKGljxgnHMXhoqMH3N0eenj
PbpFhl71CsZB/DURaBXBiYA2N+bHVgkWMFHP57jRYGlLNNWFfqZiHIJ6Lo47i2YrkmFwRNYpUxLJ
IXd/0Xgdjv/WZYKEouvJBS7kDwoLpu3rpNp/7x/4vUMf1r9gQz7K3p57f5CKRyZI47BvPYOdKDcD
uiKTXt6+kIwn7X0nnX6rKOxBjBknw1DafQzeKItHpuUjkEufy1R8useImmwuilfZ8jRPGUs9Ifaf
3NoYqPeMHmU8sxA0Nhz3QqrJBkCIgmVKJ82GqDdyFKoJSSUFfhBEHPdZnpc6D7tPPcLqwdx3BUfI
WbEQMtfnxdnK0xQ+RUcRfUaXLySWVVw3ikR2qj1E7sh2mW0KXiDV8x6wC/8GdPNA3viFpYSZ0S3+
vW2m5XaJDf+d0L0UuOt9uzBCeSL8CRYBJkoi4X07p6BxAkCE6o9WbFisT+XuZRrk12wGrsn1VSKR
1pgpJjdZbQ1atG69h35oLdNctjUY4Ka9Ii2OZc/707Sgsu8u3YcEMJ75WO0yZU14cDhaDJV4OU9T
Ju/OYsEZ4NB8v6UJ+ij7dYd4hZ6bOUB8fAbAC6keOW5hggn9RsboHOHUqxrIgVa720VGeWZTESOS
rLG2CuByjoaWI9sDs/QHOkFfz5tAt0dQQrSTsamDFts7Mphjr3EqX/c+mkXJ02/wm9BfQOYEpMvh
MBtjw0RrISSPjtCAypTHkcevQqd15Xq0Wi8Dm/0M8oBI0b61eCOx2J+fvs7mn9j6tPcQBfcBV7R8
Po3Kx5fYpWZ6HBO25fBkKOmFgl9JQP0O+OKO9PzHSeiW4dbsqTPgtNZkeDXk89nPURlT+607KL30
YOm67h/ZjI5+kicArMaNxr7dJeaY/6+Y2JxpLJ0mEU7x83L6n4YoGbabsfoVm2ruUtr3adOn9aqR
QdIlZW3eHBtvR/2HIIJgRcVO/1VO55TDw1HJV5u1HAMBtWoR8HbV4KUY3lq6vab+LSaO/HNO6yC4
6qgS6SHOZ+yi2tydP0DiqCgLgEGGtBVAcBmsvWfiKeHPyXo9ZnVbURJY9dLAmFjrO9UWBjwETaF6
Y2v7SixxK0qPBhwfBzDqyNqICbIS9IQ5Bo3NlTYSmVMWI5iQkILNrXdW5HaU9N/+Z4Iekw1aBeGw
vnpjjBYfX37tcrYiYV5Ghj3C7DbfhhiG8SVkRKs1sk3R9dH+hNLvF4UR1VJjSx6j1t8sEPUTkt5P
AjyescaYBKc1ISpBGaPMatzQelkL6XHFD0u6sWbVVEdBHTafbmtdUNi6SYzUHmCKNt7YwKCmTDHr
c9y+4XnkP3/vddfR9zQaQO3UHeJpKjoqk2l5Z423UpHBiJ5Rt5aGhcGR0SkEIskJAm71PzOpjZnf
U14KU+vnOnm91j04gHpu+2iVICmpLib0ucDh4D8kTlzoGqJN0GBE7qCyQn0O+7Jcw5lOEsV7MF9B
3zN3AL/IsDOoJVc7daMUAfYNY8kBbS5V3+loGNtfhdPMP9VFHYN5+0ruKI+iNv51FP2+faxnZymX
qh+xQWnlZU5tprwboUrmy2t4ln1LlKlt9CxAGnooaMSwSbOTltMYZqcFpatZ/7DwocWJe9KZV+kJ
3+bwwJEpoeziY/LseR9hjIeuObT9V80oK9bJBJcGWIv3+KvMARdDP9HewPYwBUTAoWWDH+dsGWw2
eL5qEmrotb74FnHc6wf8JM/O4SVwNpR9MFR9dd8wuca5EVgTzkugwFMUE9Rq7ElICsXPo381oHFh
MrLreMbsyhb9WhBGGz3pr+ZGooTAhPLug+6J+IiDhBQ3F+wBEtmu6sHwfbEdOvVF/DldUsPmzG49
NC8fCIHG/iD6eBOznuU6ypIwLY2JjnwQafK+4nnYaJFN0DnMgvgZZLrbdanGltu3PMaisUw1k4bz
/qJLgHFp3zFSxbAeIgh7IjpFi0oeO8+HFca4ZFLbz8eTifoo6P8Ctw6bpJd5CQDE/3WdNMcgD6+g
YDq1lkFY3f9YME9osVeA+9wvpH0CVWPBluhwLl08TAe6EU94KwqLh4t5pultSE3aqo512dZhYvcr
rUeAHZKYlwClu7La3VFsJkNm2EauthHAsc2zYH0IyzThWtsXmhgF5m1DIaDGnOdBSHUgiHSLKHtN
ZcUPBeAsGogGLOesOEjDGwG2rw4x2eDsdYTopXmFEJJ02r4/Y9tkE55ijXfSSyR2Tk4FR4lRo4x/
owQLwKGhjM2ukcawXWnjySg6eHMYuzTnWY5HlZQ3pAg0bhRFwx7I8haVoCSepa3K6xL9fP84BhBt
nSyfe4/j5BiuC29cfzAtGBonlLfhvrIYxTrDoRvUcRC5jFtyQf29bos5fj08KUIHwLF1nL0Bk5UU
80R51wXCvDiFKv+l7ctW/G1YtGxLeVT3cokNRM7rOCOlayuksyiGXqUVi/VFuQWp/BAm7rXPq34U
ePEQTsB9tV4+Fp6FdKsGrywQHzhC2ILjJ2RsKQ8REyYRcH1mPW2E/O1WjdA6h+g9VfMQDTUxsZkm
5P2WQ8h14HS6bU0Fn53cE2GgPR0FIfab5btwNHilDVDyhUz+bUQn9JCrO3tIkQi8hXlvRK6upYDL
ss5jnRel4WQxNfq3HrheyBFB2nJETY5KQFdYcdFFchuOK2PQkWMKFRSMpLAw6rHZdD1bn8+masXp
FzmXf9In0DEWW/IgKbSIsIVhMhAZct0whnCMuVNvUcsIENf32wHI0+kLrv/00vW4Sdi6o7/KqRIK
Cx8ns5NHxt42E6eiMEvZIh+L7xiMHVSQLP2Zs/nsBrkczm5GjqrPVIRTWcIHRXQvTEAv37KHl9HN
xDNnd/B6DY7izlHBqFsnCrgxzvTAH/ef23bldvAwyGS6iybWYBVFtfurjmmmoRIG+3iT6c6lVyzm
FwyYqjmH9TmHXwgj7OcAFL+XCTzVOOjY0BkecXUe+mtcWf25/MDiTu4VUsSOJCRVvzdqiZ+eXeaj
72SiNiyUVTDjreOdn9ppUi7bhXJvRjcvpL4Z0Bp3TbqxXWOUjD1vV8yyIzevKG5CemZ+dp/sutly
NOmF6iAXAw6bXxHkb3viud/sf7eBYC9ZVo2g8vBggZVGijWmumS8ahU2kbL7nL/RtJoYr5MOQh7i
3cG0YUHojp/Nhlpda9t/I+S8yt6ly9VupZL7MqhuJ4hl70iUOzMAP2oueP/pnuopnb6K3eHA/W3G
8xlGbg7n8OhFtmHodM6YPOVrq/H5j3DrLMLmHSyZj5EhdIJWg2+qRf1UUlgp/3y64BuNO+QZvVJB
MY8TqdGZ52ptsa5t+qvl1hI/3uVNCnb64JGsT71xMgM883ewn/8L9uKk5y7jxo50UY6N/I+cg2cw
y/dJUEyiaKH10ZMND/x6+sDCUh4goatNQnskJlv/s+So0cRQ9TgJWosWFpkU6FHbkRmPg8deDjFJ
geK6kE8uInk4dgmeh9kxeKn7MV80yzpi4fI2HgjQV+ztUHMyX91PcBwIZBiqu6OcqGWv/mFhqcON
jmSsdfFEXe6PGfP+6XBtN4+KAjQ5zFIEHojBg6JfhVaulNHOWaviv+zy4vgrA/J9AA0jwbx00/Mg
XDxi+PAAulyerv+ekE+p+3FzP7XrzqnijXHWCuV2As2+w7EVz1lGJsU54ySFZaror4QZDDg406c4
fLzx+n1k+fHZjYQ6XwW8OgEmjVjXCdhqiSzwVHhMVRWL/lIQ02sCxg9S3EB54X37TkJ804Waai8v
ShLNr1eoMxN5T+hxISJ02KwCm7wj7gLhJJRZynMwyAbQNddJu0VGsWhLkB5fNu1u0C8ItvF2QXId
SNTgprR/rnxyFqA5BB1znMqv59v3lngbHEGlq5eMKLAnKExFGAQe3N9Zvv+0h91OstIYF46sSyAD
/ANLZVLhu/qc6yMa5fZFoiNqRBcuk15zaakLPD6WNjOUQIhZ2RBbDzt4bud1EiZuXBkpkF5fVxJp
pTiH+xvfenqGYzY1jPheDKJlm55C40qWncPP5Xo1W6Gf3klwhJxdocFouR+VVFQrgGH+W1MECuYL
BzV1tBkjXb9sZnOYfVO31lmmg5ghpB3ieZssMqESufpQ8Q6W84Pg3atDAlPHU+YoApDvHHmjPzoB
nUO51g8rFiNuohkmJMWoVrE3ZuVdNJ5TLV6XE4MlqA5MHM8o4BrxsjegW2/B3btUaUTBzyvv7L14
/8zdjt8NmnYuvTu1PG3UiMvwgeaBz5CtLa1GwmDCDz8WR89Vn1DIo0exuA6iUwqNlDRPTCDxNpbj
iew498mJ13bP2SmQzdZHIR/YOLNQoroYXfVo3pyGtlf6czE9ZRidxld0L4tuoFui/at5GvqZoTfS
G6rh6654FQdcgVMqg6vBgaZPxHKemEm3kQmoZIkIxzCSL+f3b/hChvHqynG4v1ZQgzes0X6NeAHl
6qZQIEC9ID2hTgN+Eju48MJ8mR1FM56wreZtpRjO4YKfgivghR8hZkoHz5EmlXamZ3QLJmoTW9Qx
66ukuuyYzqYh+7snnDJ8s7dm/mmgepkV/X2EFPb/QzPjylgdYNgHIWkAVsB6XmayM2wtV7tiwp19
MYyPo+R4NY+LlBIi9yYjwwzzOY2dyBRrndDENmYwb5M/AfK72/gkIqDZXbHEpVFx61+hkWgiwwUW
EJ38ekz/mIbjCBS1kHhWYspRKrhIf20VoQe5GRh1zjPa3J/0GKXyD8nX4aqWV9fI/VbbjvhnDn1W
Pw+PrmeA9jrNslYHw4uJ2Z4QXh1EgVH5oTe3f8aPMQEM6hQ7tJ+6b9+wur3h1l060hQlbVBO+4HV
KTxoVCzypTNabtYrTQ9Zx71GcUA/SVbi1yYeH/sJvk6YCRHOzgXYDI87rA0fhlTw079JHKseWG88
rN+sjM6ejaryfgqCPYsBpdDeVBWiIkEgn5u26gibl2+1Clo/eV3KXe8eOTd7AVxOJR8V4xMu9M5l
hTAcFTkd/BaktyP/w959C/KMe3A+UAa7pqT74vQNe1tmyE7ul2WYowUT3n4XO4V+xaBKyny7ThzF
fxAYc1anpZvu/6YTBW/RtCLHza55E5Wax2XMkEiaCWKPUUMVq0yFCN0WwBV2PoKS8esBu9bn1Nfe
FM1U+yhOHbPyO89B4juJR7Olys+EffdGBBtP8hg3xqClMvV/axxqdQiDt1aWMA2R+4H3WmCoPyFm
i35NTTQu2rH6rIzaR2/vGvIZh3QrP3aLzvIbQlQPLoBZJyap5EKpWZ5F+BP+AUCeGmKzfX18WNBk
9WEtK8wf4wzSqbe76TUxox+x3Qf0ejpP7ZY9CN0oK7v1L0OTCig2UUL+y/bxIyNSsfbiMuIsYVko
mQ37/wksLNNN2cyqxw7jIwcyLpdoxQrNJCCeHfLmHXxkiyWR+V45QT31swqhgRW9HGtXNlBxnPcS
ASoP9ZyMG+B3Sybj+HGYTki1THwLjJwXC0YYgy0LPPSilLJolal08sINnWPZeQG9hzSkHgyBAmIf
fbpp4bNJD0j1NEL0eFd7ZaW7XgZJ8K5tV/kvpXMVzxiMNcYxgtT7VmdKeHLQAhH4Kyn+u/a1ynTe
6veF40gLpFlVc8D96LzGJeC+H2CgZupz5t1D4qgAVMQfjAfoB3Cm8R7/+EFH6ihPkSEBLfoa/ChU
ugkJazuyg7dIAAk8vvtKdyUzf60O53tybsz7hzT9NPWMrmimiW/qKLhGizqixoUxOQv45TK5xkY8
ss/+FTf8qnM3Thd8qqf/T+fugwxIlMhvtGN/ujj96nj6ozaW3JrElmKYOKcJmgH7m0EnVCJNXiN7
unAwPVE5qMu52sz6DRt9ThojrLFjfJiwXN2pCHTTR5AgHjaI95xHnl9pMPRTNUqoTkJ1dFSU12jq
o0f+URvHV01i0D10IcT+CNHogSrSeBySa0Ks3c0Nb3ok+H2u1dGepUZOWot89U1ggvYNq8K+HM27
K5ZF43sJUm4zfoxidJWw77Xq4PutbeGLh8zYoWU69YQLxiVEpahrb6s7RAQ+qCqme033yL7s1jnY
38nQjjBE4P07Uoe0mrRC8m/kaRtzhG7hPPrh+0fBx/XCKQgaEKK8MfSvd6fOmWsLWdqyL6eIH52b
vBC6HCxgr5KTVV+dxpfrT7Nl9hYVxcxmmjGWgftOgO3qK9PUin+Ha8MOayY8jx8fPMWYO3f4zlar
vaUGffu0FDAfqqHcXadjOM6oVesQZJZWub9I6BdKfceY5WRQJJAodaf8AJWgKgW8IKosX7/Hbmlu
fXrcVrPz+ciSSU59o+qrOW1yiUX+GXw+JCPz0ROYGK4AONOR59nC3Mc2noiKX7jJFTHykObpAgFS
tNGmIrM9QLjaQoq2XqW/Rf9mXU7RmzqpFbr+m3j/zlgjkHfoA6hdjcsOM+5SiFMbUqMu2TN7NvCY
Eds0mv5s1+7xGEP+CQl/5ef6wcI7PBidEJouHQuyE/9qLstUJqNW7NJ2qgRwz43hGB96JNDDTs0A
LKiYAWBA7hDtCF83NSTPImo07m5LVk7syWOaUdN5S7hhqRAUALyW6ZCz0FFKKwPU1Qf7UvYqAVZE
Ag3iTsLZlXPOlFOz9yEtng8db9vlwnGePxCJJE54ISJ6Lj9JdcBB6At9hzDGzL/JkMlRIQk/Q6aY
dQEP+WZxdU+84a5ooQopF2H6q87vPbqEP8q/b1kVRrju+BxaJ4fLk33+WnbRl7OrnKFYFdFk7oHn
G4ZOCxvLz12tvoioheAVL4xyl4OHjS9y0W34LeWhh1lSfgUnhCK1ttwx5fc6+rdp59BaVsrZmWGk
safztEtd54GKikEw0ezevdMYNxH5cOE+t371KpaNj2HxtYeNspfT0VLpf6OzxMP2qbNRAgllXggZ
nbaRHAeWvrsK49+oNdRoDu/dDMqlB3nca7usSFJQLvbcjX3CuLOFbx0QP8e2fvBGtH0kN/giMDuH
MN8sLYedxWvZtIwOrWXHi8fTW2b3ONHLhtKZxxLkCeHJBTaMGG1RsE08R+freD0no6HyLy2eBf68
JOAqSbKyenK8LwWMunstvnApeb/0ZMhroeAHIU4NppHMg62l63YoNzRpE07r6AmNyhsehXVF4g6h
MDBQ6boUBxPmqgkv6N1IILuJcBAWG/gpLdimcdH0LyAIr+lPMkfEL94FvUQfENpAFBT/ewJnbGSW
LiYv4tfrlWi2efahX4rn9n9kooIiyYcHqod/LUzj1VfWPVL+sSvZb3bmRSDE3DQ7xzjbhTpksDYN
Zg2I55ynz6PRb4PEJtOAic3mRwSgVNXjyTteVwiVamOeyyxQRQXmd8HrOk93n3ewiQgt7ndO+lTX
/SXgprzMFwkNjvLbYVJa2EE6zIXAu24lPNZjOyqCvKQ4HueZPpRXlLZ6EKqfXTggdubr+srPtS2m
mZqYphQa38MV2ekwZJ721gqnW61Tk0Qk4e+vWZTYNQg8JSxHpPrLVNqC+QZroEdRIIgHCl3QneRf
0nGIhR+Hs6PjOuAXlD4sW+FOc/u643lms0dTkEo+UaxnpgW5VEMtmvGuo3ab+iP6SYEsXVrplc1l
pUuAgeEh1LR3yTlsVF5LJSmeDHm32oeklCRoJnpRQRO1GYX2f+MLhutOIqKFtbujXzWZrZ9dfWhu
96U1vfrqmZHOryscB9suT2C/u+VXR8xP3+xVUBrGv8rbsVt0Sc7ueuMhu7XtL/ljV0w+WAQyhWV9
FrGN7CkaXKteArFRvfLmE5zPG8k4Z8APOAGz977yUCrzzxNXxPMu1RPIyCcv9ZCyo5475YgA2/mc
ythjPPpFU/+LyKLVIKxV8F8DHLc7w05OipZOxlxCUZ8NQGY4Df/CwC4FdUoxx5Jw64SAB31mRb6U
DBmzw7BlQPMGcK8kH76xkYwOuumcy9WGuUQcJ5823KCgeRL4NQTKD1XPb1fFYFpMYETfPbIq8Lpp
7NQ8fLDSGAGpd8QsE4BbrPXMBN+aqkLpdPUddPX3WzAlA0vVTTFZGcPabFnDBSv4ghTmAn7h63/L
tBZOnbDwH6oJIY9IPGLA+jnmJa0jgNbgox470JYtg8WgSWxprmhFjNhSAjVG8LUVylbotj0Or3MI
hKbJHlH4Sr2TgPX0lfhx+eBxd20ERywrTPPQ79G+Nc99Vstrg3+V3gL7dzoBbT3g1BD/G30HggNU
lZaW6RwYptqODo/OSu0OaCG8PeaUfG+iDdLVN8nmwaRVLbi1Y8CNADKqsgbI5Od33xXkHQ51TcQq
fJMP83+vgia1v+TN2xCBtMGZj/Zt9l+XTUVCKdwjevOoqa7eqAt0yxlL0+iYzWN9X+1XV13gv0p/
jPWb05Uza7eYGSfl1M/VcjQqFPlzVnEWpFJaHmZo3GpkXxx5p1H+qU2ajJpzK177ShwHR3LgB8Xy
gmc5zHFrDcbLSxjP1skvIpyP0NcLQp149pZmyNsqPribL94oEKUCeRAs+YvhVaw97d6nnMsxr9Ns
OCjKRq81LV8FymB0mhsX+BMf6qPrUzgBXkChtfIjFNV1POJ6wn8tIgcyjLRnMTI3hmGRrfRpj2XM
pQVKmYwLbc7Vqx5OkP1KyWWhuvbOF2l5nm/7YVqFlMozI4WS6vx07/zUJnjcgOvVtYYH3ReVIl04
voZ6c+ZdgTNv9McGL8Q2fVKdeZC76Sl6eV+r22D471wELbAz3LEn2buXkIpV6NZQfDAQCxNc1FDs
Bzpbev255I0pNabna7YDLNQyQ8tvpImNFNf+Xa7XwG33oJAKylMCreNJwzirVh3CRchvbEoB9eY1
miKQmKOcxjG9Qi1B7EeESlC14aHr2WAxjkzWv3a1kbAxE0X2iymK4Dsl3sUXEB+LGdk1inW6y3eL
ScwrADnjMebFTWnELa6pHFafJ0e3azB5xSbt84gPT46qB77wM/M14RlMYWMFuhJQdzO0vt2g/iqL
PB83NhEZGFzPDonAsqrOXa5vET+9P7QjaEDpB5Ihfjil4HKNeLKzaflLAH5GgXaU72U/bynZaVUw
9z66aj/k+3vUnl8xsNxAM4zPFBXdFP1OIyH4DEanwd6exnzBJW77J1cCBRC7WaKy0fGMnaH1DtAm
1+x5iEcQiYVleMcNrz4uKuLxfuN3y7oQubqp9Hug9AZ6WFFf4z6cXePUZeRjhZPoCGMEOdtjxYvm
IFGaFso4ufeBzYeuWk/xODP/DUhGRSg8i+lOrELMNuhvXzsOArBWvO/WD9S1A6tB02cP/a7xcHAw
9vg6q1k+rlybFk9+wY5IbmJ5jC3RdQ7a2t9W5m+8vk8kbM5+UeAKPCJzXa98+SVMKeaPShBeZhuv
imz7mdRVQ0aCFGhK7KK4M3qv3k5Hmth8CDNn3/774ZJg5xwDySLaYHmxNYTFeOZ0Vi0sEfhJwaro
F0QTlVnZhWiJsbBVLBdpe9iPkkCQXiEh/3mNiplccdzmR6elC+ZS5yR2/TK/SSyDzLr49Vlnl0yU
6JErtD0HhsB+LRDHZ1njr++6hZ9dDw0jSnYB63a5fXFObaThgEtrsAi7awcbF0FGW9yOCLlZuETw
OEofHN4muofBnawPrCv9l7MHdcLJWUuZ4xEfZPFehN/RBeeHgZBNWtow0ngfTvalzJ+PP9N8kODY
r22o3rtyVYxwsPLfeBmj/nX+bLT/uikR+FRfIUWSwzcQ/627Z6MRxuf/o0cWToNOgC8qaEiGwDIo
mav3Gj1q7t0a4a+3Qz9Dd1TZ5D60rgBnWSH5XmPcU+PTBh4aDf+HhkqpIO0sFfouS3fYZ2S8NrCb
D0om7O7kJNV49lulw1TNjOJVKhgZfQNfAiI3HivoxsfIhH5uGGr1UYg1kvf3iMyGu8PFlTbntpe3
cRnCTbTZmouG8MTDi0dxEE3jbczs09fZ2xa2HPoCis05LRzZ3hXid3bF4LpxQuqm/WbxO1NT8DIW
ORZ+40y90I2o89tgR7loMtaChdQ8WQOX2X6KQ8AD1CWtO/hShLzalWm0nNwPE/47hQV3CCI8Nzjo
VnQQDigAa1EMUiLyOZbGo48WbT9HcF9/a+wdeyJ6KzdYNUviKXH3LtJTXciNkIQx9AyiaAdUUh1m
VUUM1SNB3zVRU2oyABI/OlF2ZI7MRVratu7XF8MEB2aX0LC+tplqo8h0ab5DImgsm99Y69gvQgQp
aAMIkuNpylCkLjhgdIjK9lrI1mYrSnyTeVqTMjhrV6kfOdI6JpoaWf8sTfwSnsJYdsp5B0HIlfCm
QuJmmADEEG6tltTD+s2KPTZbVvLgnjU3YGhUqGX1CPy3dxpxjmc/ydGrC20y9R2/1aMAfSzKXH2p
u87sPNp3NaNNPzR2z2hVkIzE/8vqbLqu0TSbs8nJ/MFeTv7QI+i0iBtZGc5rPPh6cpUbRih1SAFz
A6DULVOEgVeLyNONk4ChLCosTnP74mYIIP6BdC0+EYa7g9XR/ohhYkElgQWABC6VOzGd1Kcm1e3L
Ko9oicy9VSAugUWHYCgjA+eeBE2oXhl3V2BTVYWpE4XnvYJ27GSU8iwtJwJ5hsgVVSzh/ES/Jz+V
qgeRDVUdD9s5LEh5j0MRaR+nAykUPKOs8LoeVaQKe2Kvr7mT5+PIayhbJhnoZ/QZ3RHJUa+tqCQB
pCqh0Yk/FTyUh5R79BCIHOok/3/CZGnHwy2Ps88V7sQ0Ev+0lWzJ3/GVDV74Q1JaxTQT59Q6GxkE
UgV/b9ZUMg5BbIUq1rxbN44lRSMQMDoIZ83lXXYaZi/qHu+SJKyoQeELw80d09gKoqMYEJEDNKTz
OJlqD3kylUWw3+FSgjsZhdktV2DlzUAp5eeMAtOHRvas2jFXDRSGMmaEwNgELFLXtASPmpJX2A33
Y5/5MvM0X4gzs+F+LRc2wRzlNfO7X4VARgP0z0snRwt5KXUOX0vqfULn7ywQP3S0zIbp3dNVEZpT
yuG78hFoAsZ4wcvl3kwXmwWehIzb/FDVQChATQ3FOzWVwlqc5NISTfLgPumQDpol1zCLahUWRjjl
daWp0OCI3jQxycmk1a0IL0u8+xzCFrkHr0tzuq5+Ac3u38e9Vrpp8In+hdE6z2z8hZOuev4IZbt0
CO+f1zHbcno6Y2KriskrZZXYWij3SUaQBH0WtTwVdWJr22jp2GqLmJ8UZr8Jxjwc76ISK/C7C5aJ
DwW1r2l/YW+yOLIqPz0qLBU7X7hzRXsxyLNa8qpEOkPgbVHKNqtdsIXQktb2JUQ1qJoERDpcqVWZ
g9/yMcnLqc55TqWqt8lgwLheSTi3ULaVqitRMyPyxj9o2Rtiz+/I2pbiOUr1Yy4m3Xg/wq0SHqT3
7NPYXeB+nJiR4KKnmxDHco7n0naikJ3sTAurNoiTkR2fcJ5/7800AplwcNatvMANT8DcmCOFolqX
7AQs3yGy798r5qN7vH/EWkisFgrFY54eaGLfySusWv1tyyR0Biye6C/ftuuUS/v4wC1EoOUXMH87
ZPFhO6nXppw/T4psY3xGPsAROIgPbVry2yfxWQ+qpUkn4t7/NZkJX6f4DacZhmmi61m+6qDV5L5P
31nYcA4g8040kTx9qjkfRMtPiLH7Lsq1SJjJWDG6N3BamuHkt/N6NkoP8X6b0JuyQpSir1u5Opse
NZWfSd7eGMEjatvaIUTD27Me/l6mhfg+ci5RF6EuYrJg0fWgHkaVGjV7iJyJgBKpy/AEjS7qRo1l
A98TJATZXJQl9qQ/TT9bVHKGzR703DkiaKJl07yoY7FdXo8OjTflOJBYTpiMSUwKgAmTRq8TXUXa
fNNLF5xx0uw000lSqrLStAUmJYqhvNyh6AGikYrIQhdQvr7JflGhy3aV2QDDZc/W1Mx+75e7cWX8
LF+o7F/M0lpwMzoFdjc3zWZi07kwoZHdM7QZ9YIA7wb8L6p6e2pXICejYbwiBZveacPxNfzbOjj/
3ZcTdS+jspbDDTEaovSXaXq8398gOSdY8be3TSBeGrAjdASd1hW/LuCNYmu88Tuudn8HHqi7m6QK
9Qqe7tqeaovIGt8XoYWDf/gdclhb8GM6AsKEZqQe/4MgTRRD93m5Pu/en6g3XFP2dkJ1fwUyxLXb
0yxq2aaBy6/tFhvqzeRIHCHzANaPLN5PbLkozJKBZNwLDaGDT9m6fE+A91wLpbmll8ehEs+IBVks
uKVMPAgvPHi8MbQjJCEyp231UyKekTuyzng20fWhGFnDJ2Ntu8DoUUBEaXcrgIuiyF6UDNhcvMTs
GUN+ql13eZ+SgkAKks63Rj010/uhI3fAOYw8J8oMMXC7fGTg9NVlonvlYqHCHP8UYKqqBEuddhEP
1Lpa5zLSXuXjukhIirFRjG2x2n6h+PcSJb4R5wmkNialCl8j6Dz677UcGiVktwgHFEw8b4Kr+wJB
6Bivad9Kp5QheIt/EbZ4pgtMdLzsBysZzNhQtYweLIeb82B420z5WYtmW6WKy+o0UtAVipLBA5QX
QHysddGaKz1XbkOx5O/O/1lo5elN2RM2MZx90pIHFCUYBhFTcntRBv3R75kFMxyz8r3/PjBYKhGp
IdWc5BH5FsuLGq+PO68JvVd2sRWMDpdOciwXCj2k3EZ+tVzGT0ijcy1BIv6+ir6DuuGj3uuhDfD8
zz+VRDB6k5nh7xeaUVM1ZO+RJS3QjcFzvblmvz3p7QSzqiyhObA+Ghm4QdeM5krRAsVISA1J4C8D
+ND4jo++LltNrjMFbmeEiL+X1ofONIgzBQ5bI6wmthaz6G/BzgP9Vu0UBj5CFNG7kv3sb+wTZkZl
JB4KnOUvsWvTwEpEeqsk0syzZEtFvyNHxGsmR1HGas3T15h21y5EmnpzMUPGxkN9ZnJNDhMFeuF6
HnQdkFGLG38IUlaItXFXj4an2d2FlIzZnqWqbiAY3apRU6hMbvZPOEnQXvoSlX0TtvIoQTIzxFFT
YYD/IP943sMtFKKAXakXSXTZffIuiSG8K40PL+hsnIJn0UgcFC1MoGsfR65qsFr4LD4zMcqHjo2F
91f+/c2H2sb0Yqcpfr3sj5f6iYvCRAyS+5WxqIbrH3010V1S+LjPUS6aD2ShGlc075vlydmumScG
2ykCqteji2bZTUjfLr/Fo0hlwVXWgRCe259fE4HIJa5rioTfutrwym+/0snE+Dn+BtJLXJuNlD6i
K/mgq5pSXaNwK24pu2ZJsdZRQc/Z/2HsOlnWQw4RUmgAeTO9PL/bZGe+esYzSXBQhZ2xXmBJ2pjK
GrJzuCG3+Nv0LxuGWqMKFPvSbNV/LLmEa1nIhxzLws9R06/ylpCLHz0cLUns/DVxVFFoUHUqvZrh
xq1GmPNjIm0sN67O3ubyExT6O8bcAr/FDTsJ5AfGalhLTMZ6IfxLSL3RDGhWBzJ1coCDVoOiK2SC
o9tIwKUK8SxYyND5DWdvaKc1aklCfWB51/5k7PZfyteQ7YzOuQZNB/APe/ifHrUDgVUVqdowyQ5K
mSh8kTWYXpdyCPQtx8xtYd1xGtWRdYm6dRlXj0ObkC1T2aNeIPOwM+ZrwmZCQUDkC+ZSVvA3l1kB
SvdSBNL4sv5Y6SueecLjln44H1jIdT0QjHQVHRFlYI2LpEzYnjHNhEvlHWg6WOvVpXolstk39CjP
4FwrHQuWarmW+9+7vb0QqL4YklLWFXiLc60iVgl6TdKZ7thKRY8Z00iY5KNkmBhc1BkjDbn8zzIs
1Rt9YVQjOqenHZFAifoOfDblG82RHibj9pDuP1pEHglI/x3Ph7T1sySaVwrRtgbGgzhiB7xzkUNd
YsWUh+sEBm3pZl/ACNukhGNI6Eo3RMdQwBh6l1WZF/287SeqVA7t6vuTqPGfhrQWkdMIaskxSoFN
vnxCtu/cdRVU0WuULJzG9ADrHL21UKYxMLZUxZRrMKC2WePN/k1i+XKSksnvP2ebvdkOugOp/QEV
U4jRlMEODzx3R+/UIpYBGvKnDpTip4FCp5iPGVMX01hoPzVQOiosI5JxopNBHHG+CQZC5E/WjsM5
Ac1P3z16cQWU9io5CzwKYVd7Pu9FvydAXzmW1F3Dp2YF/4Y5Ejh+KxWBMGgmMZsB/NrSbSJg6Zmn
B0T35BYQIJ6FsttmhU3dddtr7b2ot90V/FnnCGi6jMIWzxJEqtM+ESRSzp0wUl2+//fj3mRGMM2m
TS+aIhinElkOiVqJ5/Cmo5e9w4UvGFnVpckn4x6EEiHxGHSqfmp5OBQAQJfhToId3E0LlnB5IYNf
GrSHyUv3uJdnq3//uUZoefp39MAqJk8IAwF5uyV1abukeSyNvY6lruPFU0aixUCTusqvF2zUsJfg
LXGftHZcKyOfCZ5i/hIAMSeKuYKhv3a82W0cw/mpsBkEyEm8yZleWjH+uq+0bXMmICxdDEX3zVqw
WvUmcXfR1ooqa2BfFL4HWG7gn5x169Wiwgy76fxve2v3woHFjNuDO31sBldZWoeybxQLUY3xtGSg
aHVXHDtW0biwzIiiphpBLP9EjxkMIRs7qEHAGWeu+91dd1y26ef2XNds59FNjuAMB8cNjHat8mwa
Fyj2nlSjQxPHrBlJczynn4fnsSwpaGC+W9Uma0sx9x8j6iZXz6+3i16wyqpGuldxJ9vmo732Fo3l
6L0DOtoG1goO68HV61trOR85i4WqKEbaBPz9tg1ln4/XAsntFaJLCweTY8Q8TE4CH1iR+N/jdcOa
DRCSagN0ltaVcr+KWJD7jI0fvxm81lpDC6nvcu1BMxw0hDLD1JEJSHEw6zax2FqD/khJsBcWisYT
ILiZ0RuXQEw/1xARVnYQ2s4eJqJS6MU2eLlEwDFYNlt9y8t1titM3jxMJLXcydl/esOccjwAJxyl
aoBz/Ea+Q+Cxti4hiMcWXDKH9ci6KZul0NHz5vKlqz1eSUyJTMZV9fWyC1WKkfmzfnrxNqgJb9HC
Azoj+leoqrzpZ94rLFSifwzsXHsxtUNsa0cn5RkYesee22kMgk2Zwq4voKyAn39WVQsJUyGAYHp8
g5m1w5+LzYvurzyc/X21DejOX2+V/SPJojWqW//wJ0vb9JEzynpgdfOoTJ/pRZPArkGV/MKOweXa
FAv/xtxjSky5SV91fHQLcHjiWVw75c7kB+dtcMa+Xe9S7wqIN6HgBULHq6FsY4YPlIeRFZ4llRfq
JKrC9RvCGYJFZnVOD/OLGSTWL8OQVQYf7wWsyNz5dOSJMXzCCZIecFKrON3ygW5aRhNG8plcAFxq
N0UQ+bwz4TlZYOorPv0O3xdp1c3Xq3eAfK1SEJvZeLefq62CVqv3s9gCvvPzwsE/10vu52zCYvje
/Tttgh8DUSBg3uWKu5Du3q65SVVf+ZFS4RtJppTSoN8IKnunHxc8Edr7G5nQzhodu7H7hvO9N178
DDIzf9juA7VeroP1j5TT/1Te8frs/Ut+ByZ7ysm2YZl9iuuNhVUfRMHqtRiSaOF+0bxVbCnXm7tD
ZVaueN1mQpjbSYiixJDsSjA5oh20V9o6UvLPujyLofLXQvpCfchm/p1IzG5tFBugbacEO2fbDhbP
BMZEhFNuXMzsnF3Vy7HzpnBnFz6v3WSXrnG7UxIhN0aNXDbJqlqwm2PFJVO+xiKxOIrIBH/iirXN
uPg/r8LnR1bQFvuJHSw1e8glTL9LGWxiP8SOLpVjfJLkZ6rczX0mtVgm91wnVruWExTZEWjJGIQK
ic/G/qk/qnLW9R45qHtQUaMgRNTWE1Vec82YmbrJMMqAW9+pa6kUskJl3I2ZbRkLDSwKFNlh45p8
/4XWEAZPtjMRfwNvHUdVEJuDF5OoT8w0oFifEYIF4DjFSbSjlQNYjvlcby1l5iaa2yNjHFyWNSm+
M77WnHggee1/iSV2lmScoCyX7f45zQJtR34rkUnhvULS39wiPaZlHHRL8UkCE4tksMs2pl0jmsHQ
7/3NMYRb9iE05YdnbLjRopjcDbgA834AcCVR+LWyBuIhhgpeevPCW0xS1PQ5S6IdQnqyRNrXvHER
Qv0yTMmaMAa90Dh3bUBB8HKhWp47EAfBEZ0xVLm8Foy7EI/DAf0ggfC8F3w5MTOFTD8FBhrjx4k4
ZVuJE7+2VWzum8Azqg4fK1/2lvUQPNuBefx4joFLwFkS0HW3dspgzy0+5JdxqohdmQ4GsqB8NDdW
GO4DkTJOIz+u4aC6cU8HENcKJ7aMRqD4SeyA+j9S0lSbApOAv7Lz0iILrDJoHQsTvbE/P1Tg7OHn
OJFqq5XVZlAKPor1xRAX7TXYi8RLnpzCa4Jf3ROy3fsn8C/EuRxV/9t9Wu4DScMJ6rU6uCx2dBR9
fmnhaifzI3SU4N0nvRSbFaZpM3XhiT1r08PgDAtiM98SyFUjbNwTb0fZgDlYcel49Ax/jXySoZoO
lggdSJB4Ei3j2p4hgwP0YAhgF1gOKDFyPwze7fICQMFfCF42xgeKmPyNzDTIHglzbUE4IwTWUQLP
hSfzeGv356OTAvu2gzeHzYjOC6rsfniIFrxNVCTwTqIMOEH0Ye/84s6VX7ytF3ZVrBa52gNfCsS1
xGDrAapIyVOwR8D9Hn6LhgSrzjbOEgOztg624+dQzu1TEA6ZUhHW3hhbesrpY+MUtJRVD0mJBqed
tfmgpaz1DiuoWs9l8SpDvvqmblvTTmZjYtPsdfoNTqy5n3E7RaTyYmGTlzmx8+YQO9rRORUQz6nc
P3mdkx0g1UZ4FEvIkL4h0apaFPJK0YfxYfiGhCI08WurpURSvrcRGU4cz+s66AWE9AzM0pg0fnNu
2NjHSIWVtszPPDgftRaFWzVA+7xkM+M7QbKk7YgCZLMDf9jsB0awWgOmGxnjPHlwPfL0fBcaOICK
R4CMtiugLsWTocY02AmZYqjiG2xVjZeP2j8f1L3Zttt66RP4JQ4LPinkhTaznR754++DSzut6L3g
49hoU96ma/KXhD4FY30q6JzBM6hcw/SpJaTd3bV5thVSGHF2O4ujgSNqv/Q9Ww87O7oJfkiaDPX0
/ba9XMmZp7woY/BmSJqzLuEgOzhXdSIw0L173mEq6wP9iNvzni0Q4D1UNp6P6J9D45bHtsHzSx1G
vQZhsvwKAeuvre2UJQkbKLskiSKKBM7EbM2cioWTpkdIAzNiDt5Ls1kBOphKf3Dq7kOAQ7edvC6Z
XSPsQW5ETdM862M43QxOp8PNqq5J85/bjTN/6/7AfUHbm9wbTRoDglGFwMAcrn7v5GsyLQQqUAJn
bCys5QE39e8TIZBoE7bsINEFXgNiB5oTZ9ZSbkmUw1LZTSJ9UkyNhNIhIV0o85tp5CRoFadKa5f5
RLhCr90CtfQ/KDYl+0OwiFi+JGCRGe93cCfTXKG2UknFqyqaRM17dRx5dNQwZo5gofc0tFD67C5Q
MAEctv/ZjAzqEGGfjOlx2aFxBH2wAn5umUcVT4CJ+UUhTbzQoRjhQPXpgmv7qdTylJvo0BnVhLZV
/9daOOppDebizqZDm1PSJy3cjy90AJDyqfM4fPIokXb3kHZsdhgGKMq7AdmFUwmlALkquRUtjUym
45HyxTfuWcrV/dj5G6YHRVm9OxHp41EaVG6fFTJYbUaABaHPBWmuR49wPhSI5f8HUsnqO3coFkLl
Sq/PMKwnMN15QZOC1HdfJfTd/IOfjQxHwggbuTcLEmc3D/chEdfYQv3rBvpPeWaE4Z+RkP/++V1R
wrJo4BE0fGRr+Ehow+9+VfXqEtxP1y0BSKveWCVnu1vjSL07XtBVovOp9nd/6AwmV3qn5A4OVhSW
jHwvwoxPS3pr5NqAcN5SPSKS9MgsJZIlArzCi5Gl1fR1CcXF7tR2C+vEf1oY+W7qfDGt39hYoEYL
utofxLCg9wn1eH7BoQELYSImSRHnzbjvew6BAKyeiFFe+aCmqk8ZbMSPhlTJtCVm948yoNFOgYBM
I+5NMCD1STJoP0WKHhi65sjc8CSqaHbUjhuCXpnclTNsUXPMGxD1SdAab9sAFQyFJZQTHLB9ZbM7
TYCe1nf5DK16j4O7Xj1gxbKahPKCKiLXZoKi4k4yv+XKP2JBUZTau3djxhGl5c26hcFRaqnMUHbs
Qgm8lU0Qa4U1p9wlo/K08OSdJsALX3NaMO6snGc8Wi8nh6tt40iJMAhlUWthShk3GO3ow/4HeA8V
KpNudstt0RZHzY8ebdIU6iapey64o7pXn4j1pc7vaV2prA+y9qMJQaMinUeuhQ0QfX8f8LbLn3EH
KpJeYYyz7juBKPLm5yM9TZO6zZbANvX0XHAu/LQmomlF3uQEJVXl0yodQG0b5QZF27/WX98REJIi
jBwqWNmWabJXiEhmwVF1Ad8TlmUUUmwGkKpjjuIiBj8EKRIB7/OjkbvpgZ89R+vXzNHz46JwWaWF
oLYoQXQoNhwqbj4JK/Ifvwf/tyWCm01njIPhUvr6+NpxUvW4Qp475LEtCjSZ4HG5kt5WRIB4lot8
2GIE5ySn5ck5BYM9cR34W37tO7XRpA7w76GMPMiLUFLoJ1v1TYggxVWv2btEBm4HhdihYcbrVSux
RRFCxKOMKER+J1iNWplM9jVtXlgWE1v57pnmV7cf72xzxyFS8m1j1jMyNW7uN3EOvXTKfVdV0mLP
SlyaMWrsEXUm0ohthKYzw2gET5AXgjRhc1kq5JAGHWheAQemjLK8tlLhskpk4KjTJzCbfmCBUHdR
jaFrktrr9aaEBijANaRFb7OEDhLjoaW8PzChuqfCibExriWk8FAaUzMvfO2ZtSlND1YKcInBVLFj
OHMne6H943XEL0ychgfUIr9k5HlfRYOZJ2q5IPrzNFnVd4xsKpONNt/rm8xzaWQpfyytNPluWx5o
iDYNDhwcvr7HfInc+xgC1oDkbSXwwvYCq+hghvAsu8KSoIN6GwBYubfMlsXzwfL8/Wi6aqQFUyCj
tSX8vCNLLySPs4HBRecvkaz26aSZNB3Z/yHwj2auKZHo398pPUgK3ECQRd8Bnpt8hXIcpcq60In8
aIjuMvt9GQfmnc8vvJ0PKwTjSDoz2HrqvdezggjDXi7UpGtSpWS5xfgUzXIZnZREwnAT0yWLGSa+
0qOJWfYizJM0niTe5F1v5KEt0xMG7YQpO4jpisMJYmc2KzhpYj0HUdx4kkfOvPXS0qBKKS1qsdit
otBLVYqsmwdOgzPlO1qxf+HfjExjqitf/0TC8C+iwHrVcWeupw7lqUO3BfX18arPKho8QqNyrmzj
Mm7DjAPT8Dw1YJD2iee71OJ+UodH7D+hYVB+gHSZF+PUDWkKZzSBPJH+aJyl7eHkOs5N2HXo81iU
l06SVq2GhlZMHL8aFT2AzGZFgI8d8eudR0J4F7YZUuekm5fF7uGdfBVWU+8p99lf0AvwT8g6wCZ1
vAwZ0L7rCqHN4UfQipwZg6LZot/BSFG4oX4CxxRNkjelN9dIzD7Tj8vKrodmy3+o70TWkRHVT12F
468dRgdZY4TOs8OXZWBJoiUiFpvEFmWc3r/SC6uIqJ3MOu70Y/4w/RgT8AOvGXT1tjtBPXqaeiL7
j7ifcJdNxZ8EX3sGDCbE7243l5jfP7uhS9utW7hBNBwIW2PKcANVKqibA7E26ldi7UaRbFW0RXrq
5edKKdbxvnbgwrTo+gXXoIBxnBwaTnZ7ET3UaNZkdeqQkdj4cd05OpwpspehGpvKuNZIrr/teOzl
3t3eGa1X66gX9kqxA0BG/uoyAc3pHjHTOCE+l8rp9G6didtPtDHN/mg+4PkX2hRC3zFdUulCRlgQ
k2fmXYFJGcKGkYnwUwRv4AhDTl2WWasgDCsy6I9p4YR7Y6wcR0NtlZtBtb05hfDDNkl+Rh1WSgHu
TVmCpew0yeEWwRUBnQaZ76oW36O9FjVX+ZF8IerbbQozKlP3HoHvIghCmnnfcN23fRL8qfo9sCBJ
YdAhJ3JHDCvICqgld4Pj4RAYrPH06hL9iaLdeXDVmxE9xRtKqfBqCsI9DcYlSJgFlL8ffrGUgYRg
yMOF2xDKJclIxpjgezgDTt3UDj+WMSuQ/JRkV8AvNTXvs1Q8hM4oymFSb4v7OlrmZ55DzGIsoShA
6xYOEoqThS7ctv8EaiwEPvfusBuKIwiXfSdjq3xCpKZeP2sEZ0KlgkyPr05NqzxPX2zDVL0J9FEi
yul3eEO2gr4YQ55C1OsDs4LFTQPMbTj7de1B1o7rTZcuSYC7+sl8+nlRwh+GlzQHXVe6xKYYbkCz
5dNTp+znFXmQcS6tbKNCsq2LG1Fu1bxMfD64igsInCNx8ilspjPDjDgN4C9sJgDkc0lCPTDbt0o1
QWFLjrpZiDLeB65uLDq+Nz4zj0xKPqo5p6UTRjiPv5EnCLbf2COUt528HsWub7WrmzVfbY6FVlZT
KqVU/hfhCy2dgjG4HHpkgQSWr6vi62F5MyLoTkeLfPH3+y2aZKa7vwV1/jxByd2O5qhAs1D3p177
YirUPATjyZouHbGWuQro9tcz8o+hMErV/EcOhNJKdORgGMSrxHreFGm7betNrs1Pa6fMN7xxIm1o
ey1oHMT2YuV4axkjMp3JsSOE0iPf0vkyZGtntF//lNqZXkFhe2898bmJqeqz08gdIBhaLSOK1dA5
LZ04OwjHLoca1eAPRvNGA8KHUEksa44ymUzDuxFKaGBA9YuBb1dXxCTZpwZXh4WVbMcM2rWCKAf8
sYZuy8SC0rurWibUPxoxcUHh+YhLFnvNQxw+ikOF44oAJitRXrgo/hjulxtQM++TPoVQ+pJVclLK
j6Y21dwuNeGw5/HpPxEHIAKtAi41TWiH6iDIMhdmy76vS3iX10loIPAlZzZRbDJDJlXpvnqjIgXY
t/W7LyYMqgxvd3+hXitS2MJsgFTY1kGlT/T1HHkaXUmuFx966TFEoYVMbe9ScVZ8kh2MRL/AM+r5
neI1WuHTjZqfQ0ag5Ki18yFpxA64WaBXavQqbP0ZglWk3PHZcljVoJ29x6zBnV1SuCrNJcB6qXFi
ZmT6IKtpxavax4HYJB07SctfNquSBMXB8SQY9vIcLW4LqDzBfBgLkMbmqgnYXsdrJeG4Vsu+h0aI
G+N77MMyYvRO2/XiDdatWc/vcUGWzm5ux5UKvYIA1sCykIY+W5s5FSCeutpxC9nZjWC0wfRHgXjz
UyYDFcFa6hpcwsNH7uQCvvI26Oh4bNbGMJpKK8OP5I/y0GEAsbRp61Rdpp7Gw1C1oyeYzws4TFfl
hOgdk6zfzmyyGgKVzj9utge9yKtielW6MqfkqBEGLtvWrDI1NeAbuhTrnZ3DPPk3IyW3dav2bVUd
XeXqV+XztoA+R5GyVx6wxYM2QzStNQRCY5f1CycPw3x0f44zGaw5B51/kHkEJS/kZdTPnaR/erXP
guVbwj6vywlIbTc6RFHQ7Up5Mm0Lw7znfy8AeBMZVYRRqRyRQYu7YM992o+FNTo8LKFcpwuocrRE
cCEWULVbVKoyuzQceHlkhuxXd+kuuIiL504sKlS26l22qF1F0R+BNScQpl9Rn8bgxKuty+lBEYrM
VT9YHRMa8d1hjqG7mpJTbbPHNt4uvdsw2s2+X4nd7GSrHijiQGlCFQwu+EESqZcD5Z7EIr1/sVzI
GwAE4I8r0lNRHSrkp2EA5iC1wv18zUN7Ntx3bpI25CDgljkUUyFHC4XH17VWcYwuyglvz+n3+WvA
KuZmqxa8LE5OTb40Uie1O02oD/V6oGFhvd+ryyiitXXDtGV1W3+wAXXo1YCQYeWxzzCoktEBBc3J
DGk1XT6i9sbc7//IOlvRKsuuo2MXleuRnUciKcBrWPuIUhvuCwqdZBLrL57WyBWHvRHYwwfV5uYs
+7E6CqF2mQlRT4/ms0b+92MbzHVqcGg6SVsPo0EF0hlXgAzjJwwGbc4HMgQDfenDNrd9eT5zpuLg
ytkj4tmxBjSwb63hB1Uwt3Er1C4/Pfe/uuBJ5Rb0AEXN9m7nHaLct7IJwknKLd6zZWPExyRM4zJ+
q0OOSuIOVU2H+DLgKQQqD6m2M10CpV7DqXoQWTSbBZ2ebutixP5LW5pRjksD/VeZzhdrr/YRQIIp
+HuHEmwB5Sq+HHT6PTO3v4IaaSTRKxGijoTWravX24g568XRiWeZAsm/dLyNWT+HkkFsoGMZUyaG
NNfJ+gvgr/I2NydAIFjyc029dOlAWYhJ8hdL8nSet0TLlDnHeenmwX1RXgD/KzjwF+gJjz557g3n
7HXxwkpeyAWLTIkcyi35TaOSEnuFlleD9fDYCqxEDmBwW6nywcpYRu5EHOXWExi+NCoK8JeKrBjL
8fFDOOARC55sUd7tAPhdOSMIZsN0QdAaMHGhMwcEViyrGU5h0XvllzGBhYdoSmnHMz2wzks67jyq
Ay9s8EKnjMjlQozMqSFB4nTVm/16mjkkNxlvpGDx9fzTPqclzwPmXsMvE6egaIqUaanZtb7LGFtu
+yw8+bkwS3l/nAsWXePRA16sfEcL4X64pkK7FRBu2IAFau9gG64rwt3DAqIsAQArA8t2T8i4yx4Z
lzz+GRILOZESk5rCiOmKeSmbuLeWpm08jI4AEUzRgAEZg0PKI+aSv5pfcIP4lK6JtB82iHdLaoKT
YKsMkX9tBL9du8wHeNBO+yGA8V0OeY6KG4NefNItL6gvTn55rsk3qD77hRIjVq2XwsCDEFfIHakO
FQOKVNm6ygraVz89jPXgN0Tg7P1Y/Ih9jtYgkHNByPsZl9O3qEi6ZaRf7e4pgQj2ZS8jBE7u2IP+
yrhGvXrvsC1h1B+uc/6cbxod6n5rFfKkQm48bpFcBzzJ0AdKoAD/wA1T53wl+rQ4egsh2bjAlif9
kz68kg5bw1eCsPXoenMMk39AnrYTsw0unrzUPzT0lXSc8HgqMR2UBzoWAjP/hscdPnM0Wvm1llCu
Ce2fH6ZS1459CrchFHXyGx053GLvzRSGM1QGgwNEBGdRLlFLQvkzLWDgjxnwuJ1SXey6+RW6nxQ0
b5daM2wCCxj6eUQJ89SsLazBkWxLaRJNYmD3mBhW+HlmhEarb5Wn8sg8btDtrWmi/XyaWsW88xyn
//uz6nPWb1HDCQdAWVh4C1LYkckHl9kbUVazoeYWwopnjKMJs1bYwhs4rs43TrWNxjIjvSn9Q7mo
hJvH6PHk58CP+tzukcLVQCuBr3vAZWm7ZAw98stvzsWZv/5OzL0OL0UkR9vSfFRVObyMCVXssVFq
AJa6PS1EajQSl4xlqZSJZbSRh2cr+K/Qac5MEQBAb5VZZSI0IfT00uNml8tnuTYuCdn09XPiGEJa
VFqFihxc4S8IiruguG7T7Hf+NjdyS1a2hoXWx4+rVIqQzP21t5TsGtiRNi6EYHGGG3nsVOwlmolC
djVFnOAn3DT2P6WEdD+bJlkHkSgmEtobwUZf8erVq03tPEJu7iKoZQVWapxJG8gRsPqL/6QXC/bU
+kLSRTJIcgpKZyry8DAgtGvNsq8S4TOYxLndw/u0EJELVSahptv1GE5lgu70zfCqRSqZicKNxaC5
pdc5ndfg1mbjXhGIEhcsUz50HPU2qCbyJDq7OQfVPAege9sKvo3pfsLdwOouSomYUNAKbX/KiXTZ
z4I+QXjYTpAq3OmIN0x0SmeOvaOIbVWnHgggnbMFJMLUFFgF/qC6q8BePt7ASdtMFYO0w2bkP+en
zYVAiUlzg9RCPZe1mmiT+ioA9WdukIWI55z2qFbGILH/dDMFWWm4ZxBeFALhn/90yKEjJj+F/HnX
QTrFSZG7xmFJMdS9UB9atxcNPPnrum4GuHSf3PySjGgjUg56bxC+jDapjmLN3j1TdODYJVp6VJcK
TLTP1muAjytqElERx6zOO9m6XT4+HkHgOserSlGQPfTzsMDXUMZL+yDgD8wp8DsdLZB/jk4/6emt
qqtLvIIfWRuEfU4tiA2NjPHtF+v/jTMH5DSnWePynbceRyrPAyYdWXvd872JITPto+BzK8SS0ilF
tRSYz0BoLk+DJfPncRcofjF4AR6CnshdGo7lSo60AfA3Eus877aN5jDR+l9bpdafgLg/kLkFCZbw
+AWNkQ1GOlP9L2B0867IrQhf+K36O4NlXY7GBINNYaMDRsmiVqU9fifI9vDppM8JX+eXwh0IJC1v
FORJMQ8PB0t+nlDB2iKeYtfBzut3mAOdcHaMyCs3OZih7+0WPSwyNDh9mYrV+PPi6AqDc1xzqHNR
kXn0rD/9F0I+MIBpc+wPf2mh6w5s/oVp+A1i68d2LJdN84Rfhp487YlAjl/WYqRObj0L50OiWISN
eg6s5q1EntIosByZltVnSKgGFB+sCAlUvKa4OqXM0JpLbOYot0h49xyXShPzGBoGSVNMbCAj7ihq
gs6LXYcSlYJgAlwO/7uojnYLn2NcmnEdEOy03xTuKaxYOQXvznk6Oji7RcMfKCK7eOnDM91OXOZ0
6k+0S5Kv3IOMgsoH7tqx6sQZ9GM8OJVGnEm7DwMcbCpd1Apcp/Mq72DHrFHpDYsU5N7M/j0uFaCe
D5ETAd3l13fm0rATbMlvtYFReRJNC9WICIt50NywBYUhEK5ss59CQvDD/30OHpSPvb/RJ/VDa5EQ
RZbJqjg/XUr+xpkk6DI5Jorv7oYgfWP6ybttIHuqS6tD/xBK+tk5/K65uyZA6ZmN+pm4LImOgSWg
o8bJX53JqokK9LdP0KUTunMR9s0cHhdNoGpppfWmf2EIx0U7Nc/FN1A/sxsFIZ+we4fY2id85aSB
fSGeQNtVovUp0A34dhq6dOl/Qns+GxOFVMzhy7i3hSyUqUHgRJlhmzqaV4X/wIQbiPtEEGSrAJag
iHT8HjGDr7HSHxe5Sm+208j0Wr0RvnbkehhwWmDwtNeHBx2bGnby62Yf7YkHqqEzKK5zz2zqxfkJ
pXquS/dqduQsupmhjGWHOnfux+3hrHdtpl66jVWGL9aJGe1uX/eLLzv67FOoWc1VDlAFFgqC8O1M
YIhnZyghzeaQ5GCo0Lf2iPpyTv4YXNCz1Si1tUe+LeoohAH0QauXK9TbRalZGwLkcRUWLEA4kJ2Q
mzahcm8hdW0i4huOYqCXMINGRHEmE35kVbrqXAyfR7nbcPHQITApFLrlsRb2lFz+rCOryUCWWg8I
7LymSVn5o5iwM70eMkdR3d/9jWUeUXqmDf+53/Nj0BgdrjG8S2LHzUX70Wx0W1NRGevyef7mrmrR
czNhwE3LqVDizb8Ty6ufAZgNUJTyEyM8ALnZcr2hjPsfJXYgzeQ8Gc5008vtuxZ8Z4Q2rn/tDLCN
K4mE6s+iwA+otBiMkp90x3qFZOoOKFU+KVE8kqBArrEcS8NR57kmcqxNrNGBNsTFOcZzER4s3vME
/8EMP7uYNwU65mKWyA8IoMbzgG3J+ALsJduTNr+TrbUygIIlspu/+XFCQr1/tuQduQshOzMziPk/
MV61bFXZqxeCtvFD9xM6lLyCwIDU5oVTxZPWOQ2Soxw1FAYYfXJIIabhH/h9CtO5OeQzHch9mpR9
/+iDcosXWT2G85JyCJqFoFsUWMIAZOZmtnlV/vJ7vFidMrJgyZHwk2u5+napAORM66C5AEm/WnpJ
0OpdB8mdrnkk5Q5TNP23lixFiaDz35X1Lj5Lip1+pmeDLrkb9LosIOs1JUi/jMFq58alRb4bMGRI
b+O94NaI+56XhfGPWsyaELM+S8RCIrUmjcE8reWEAOJViPBaBRk+wYK97VdAPR+HbtlahBef8Vmo
WbJ4ntA2MKDRbJrR9J0rmAPZH2kd7oK1NNItn8EkWZuvK7xPI4dsjy2X3CzXIgq4zixqwvw3mlID
eQ7JXj2cID73PvOKsIzAHakzAukShIm40n7c8fhGqHbbHRRAlofCKzodutw7QdvHxzPsSrDqDk4S
2nHk6DX7GQczCqRW6afeDW9BkKo7yke9wjcH4oEQ2KQ9/jhbj/83OgeAeW06bonNwGq9Pug58+rA
9TyFDiYaDAvQeB8ZLczkWhbK2/PB3aYojiI9HSAGD0vt6PXoTEpCLgc/awL5FhDmyH0mciP9SUJc
pGuhKUzVHjk1c+c31rdg0otJP1Db/WGvtQ9J0Cdi0qACSJkepgkOtTSSzPMzp/A5086MI66PCuZp
6aEEfeUhAFqQVXWsyDw2MhdAHMecvbbek9u90w6EAQhdgL0ZgYiSbbR9plTWhonrJ+QgslswuD9C
e8AWybDvCepm6t9lq38Jul7x+18WllW+ibTlsL56/avLgPkV4UapWKZnRBLEbBNgvTgr5EWKkzHZ
4lKEmbDQeUuUGCbtEs54g5/PKAxgCeZexH1A3Vsv6wUFaOHWyY/8yIW8o4InpmjgIdhPEnXf0nKl
Jh194RqQhcSMVYHnSUl41tbDiTPWfn+mNwsVHL8PxGTzGKe7Js2Ul2hEKu6kPuXV45H3Fg6CgDmU
UygneTjWrH4pN8pKrUuwz3RLMXuV2YGX2w2kk1ycEzf/wtCwZW9cWrFVwWGCcfImyadD71FP6MTe
Z1bIienjSZPf+hr4xAjIp3IveumSKAVkwEvcb32iG1VVEpwHl9B0WckL1OTETHrf2wjyxrcHl3kp
vpREWDGEMrBg3TMp7GCpDt7dEkH7Tpm/TjJgNXIlltM644hJyH8oGtDlY/0STJhAXk9Jggut8nl9
Scu77PpiZzREuoZUTXQgdnTEHcWatFmVQVIfAJVEOj7hQHrT4Ve+nqEKO+jdsooTp17AezLFbdB5
0/7J3dRobVaNa2oSqemwdDGzg7pn+6XSqFjspayglNp4z88ncZze97M8BczmwCig9Zqe/iLxu583
g+bVWPsX5s81EmCvyV9nYStHnBoMw4E0bC6HOBaAgHOyNry6wg0vng/RKcIb86DSu9QtyRlz+I8O
6g6KCcD5BBU9vsPfDaC20QPSBHJPFjjDCzRtF/orlsybTtUsTohf9duyNJuDpEhnuWtR+1sZlAY0
rJZIbjwpheSiClO1+thKWt4+UQ1Qw/fSCTUvXhxsGkvKmL7Mwt0j25sIRIPMsyd797dvUTxq7KoF
PQQNAUGzBt5COXl/ibWNVKGdBr+kSIlBo9+j3twh+lusdiJEzokHoM0Yh/A1L8e2Q7hvSX2r6jQl
yKTZr67ft7OXFamoCf9jGnCBs3iGD5EPUBKwfzS3AscjIVxRyzZox67EXkISccCw2FzG7QmpcIKs
T7SkZ4iOlsyiWBOFuCZNhxjuJJTtZQOOHqkxGYR1mxm2a2ImyHTlrMbEVex7Pm3MUx7TW+pvtVhW
1iA6cCDPQ5ro9PK2iC3IpaAeglpbzPgvD4XnT/+mr+awzbjUvW4YbUXendgXgWb/HhQ/iswhFemJ
s75p5adXn2VIEUBTRulX/x4JLkvl0uQkSR0JEepC2piob7pzydoH1kqzEzCEL3oYJwCsM0Kyp5+N
1cNUIkyNmjFET3uNSz563t4gUEu8EMqpl4PZyOT+G0tmZ4ajDEZyKXbTAy8+QtCp+t+S4iwGOP2w
QVqYghxUQ1A9VDliiQYglI8ZT7RsAXeanDYc3P8uJ3gMDGeLA0TkdyiqXqTqJymx3fo2lOErlRgp
UKiZYY0CO5rl7W34PlSyINCdZvnyMhyY1CnStTxLb12hjXcU2vrInZUMLNhz232yGI0CVbYHuf2R
xJvpRAlwm/Gsrfa3fjgee954Dyk1mHlk9DzHKcZK0stbdyxQH8R4O4eKU0pFzw/F6V96c+C/z98d
O2OD3DhPHpctU5AU6CU5b2n+UpaIOJEcjKCfIqNmWZPB1vmvhNk0HsAv3Bk3dbZ8JPNLnWK7ZR68
pkGxa2vJZ31XOeZrq28q3VwVwgkyi1NkfY+mETm8oS5DVIjhqzKKxmnOoN2w116L9ikobY1qjpmB
N1pGqvXiLxL7+n4N81EWTHCzkuTfVmURYL9ePdaJxBpIT5G0F6MyHgBvwVMz8cN35tPgsOt+56me
7shw2SJ/bC2J16ZvDO1foM9KXLAu7FJgm6ynUmseDDvFoai53QS0i5Dx7OJ83C9OEnJq7Yg9hLA0
zcG9kmU7xREXQRKp6c0y9Dl1NhV5CB04ld+SyjZ7NDVuubNTph7vso4Pfy1qZJRX9M7VQxaEvUko
0LWncX+tz1anLUSDx+mqpb/ekd4z1iTPtf5gFVYMZENQKmGJ2dB7sWFZ3G5zzbb31VbbX5rBb+VU
495PkPmT+8h7vmeO7wk5izI4xQ/ultJ4W4muXDgN8wx4nnMWseeKcjK7HJXmmVGn4RMyn8dxfPAR
Y8nGBEQ8K0K7P+yjPxfb7TUx484pvG0XoKcXh/vcgOhO5UROwwKX7q1ilb7TNQYKZlZuCKNKKMoe
PdsFFNcPb+O++Cb3CWYO9uvuAm+jhuvmLWxaNcNdy09PTRlIs2zax6i7UmLNJkjPMXSQaxbhDecG
B3Sn4tQeeWCPpbZERCYCT2WNDe+Nduy2k9Wfou2vdF/4918VHcPTHm9b/GAq5nJ18cZuHsQUFx/n
KeLzg5JHdMpS0BxlykOwjK5O2Qcey0rRVohaKFiYMacpsAlMtkaRBXfAs43Uwx+M5EJJCdwG3MM4
AaNGR5zZkvfSwYHQbHS9RqIoLDXg/YyCH3P3YqwMq4ql/tKOBhVOhEv2LWpQybW5yKWeYR5x9vAi
361XhvHtesCqJhsQJ1UM3fzq3quUXqftrKnfkCSzaoQ/NUTC9jx0zOGgV6HdrEUoBvFnAbyqksuP
oZ9WjlnkmEecNhqngkRQPkpKqW67GPelirtfqiieRWRTPASbrwuQAf8QNJG/rqx20inMPabBDrFb
schlk4Wkyg9vNDFoL2Zc85k05fKi/VSh+Vd3t1dCpswejplpFi7bjGwOGWNQVPFaSC5d/H54Omni
KyP7k4pScB2rOQqn2069nd41crkBAlJ+jkCFIr1LHIjZB083dLs7ryqhPIU8ek9RilKGpZ/ODo13
ffB0gdzDdlXGA5eIy82NItnaRqme2UrULItP8NjK6KsZWlgXHD/g/6KuyeZ5lkDxTi9FbE/6eMJ/
PpeD8ieFTSLiRWqcTL7GIEebMbfsPzC7MnHiHDvUQRGsAFkTU5rjpKZUGIqVLKDHWJCK3HNGr5ZT
p3hUyiqq1IDvLv0/GkIPgOMqTkYeKyaJC0lI8D5iURNAUA5vHNUkTI0Yb8UZs02fATgEWbyk+iX+
zgMYiIg2SivAMXOo1GmFbh687Cdv76NiFRgaRq0nDrpd0qvHwpqbTD3Osov9M49RFzfoaqSR/+ty
4g1X/lSfs2jtNrxeQBBX7T+3gvR2C8T9RTHPa6mbXEvgstv8eRiHxQwImk1Uq6S+DXcxMJieVbj5
qBlL3B0CB12HqJsLt3PsdIYTimxEvokMp7/phvdN5l3A1GXK77kxbx0JO25Q7jPgkVEE6XmJhYOZ
YvqwmVAUtbdHwFaFB68rhh+hn7JGIBe/EwFlEymGbYXMG3oKJZavH1BlLBsoDAiDASTG7+86YFJq
hGT0iqRMKo3HsDIntcc+sD9e/ceNn5pKF6n6v3hM3EzrcmoRbqMJc95CaPIZebMraoL1JxMlZaEq
NnBw673Hwk4tHL2AjHGnA/ahwbkTWX29nip218FTmtcwgPr+UuBWc4PIVswnG8L8uWIIyLUyolWL
TO0TEBM6vF0u6vkjwuiDvshyFttJjn/IqWc4VYfPmfKEvY4W7CN3tg5RgtVFE6vB+fnCS5ux14jF
LffZ+nReVbjMzvGGDGn50OXo+uHBoynhYy6+jlxQX8quIY/377KTZfRfVunSquf9dftLIxBUI82s
b3yG2/afQ3R+FoXb3aooOWIlMx1mms/AlhsVHCLUmc/W2rti4cIT0nLDozgm+eXSrzZMryTEeFc+
KDebYSUBUkbc2kctifcS1I6a/yJY1QfnLb9PlxdijkM9NrFDxL+khsOFS/tQA4EE4Oa096gwQMzK
fhXxQbvJhtpMGpSN/IF7CIrpsHK1ItNKcJWOC8fY40AcHbvlqNvuPVtlVisLrQ/4yfRihKUevtGG
BVhWKIoSRXyONYSLXrLlM/7GGTLraBYTc1wGOXwF1maix+30cYlZdBSxcgpOuPziEbGZdjC8rgwD
QjIkQ8/TeEkxCSqukZ8VSfIVE0iERxkmMQ1eaMBGHLHFwik7hOudmL6+RmWe32uNRo1PdXKvmSF7
3GP6tfpyAJ/GhmhxmYgIqh2TrdS3cF5gWnKiboa5bdAgmYPhZl6whQgKqMMhOmtZHyIr5pAiX1Ae
pVX1qIQfpW8H3csrD52pgKSlUhJd2tAY8X/vGAOM2ChN7JEEdGBMz0XSEBnHpJ6bC765dIvjapoZ
1Cx4QvOAt6e+al7griGVTI+BLcrqavBAD/Z+mDMPKpYkxWXgy4oRVeHE8pKsK08YGRcAsJJuz+qH
fKOBvtmeBDPiWMGdQ0w44qcYeb1B2B/FGYnRwMGC8sQ2GtLzRPXoDYvbW7vEC1BSCt/t/Wvcm153
N3rUSfNriHZGUaiUTpE0AdR5YXPQ50kcLH9XGr/v+KEIOyzH1yByS/AZ/+b/6B8DKhLVq4Y7deyM
SFnTx/VSNh/UR5jkZ+QG9h5J2G7YiH+4EzeH+91xJwaLCi8vloSG+cClsKPzQNUohixBSA7qaCUr
aRq49khz8WpCkWWy1nMn71sD0YT0P7qqMzQgpDP5X22uZekGXOOCHL2sh54gXZrTTaHLO9vOUejK
eQ3ItoSMXffgJNeq/y7jgwOsvWn2uYN1BaTUUS0EPzM/0hCtDuLry1aBz0l3w9jXA0ay1FqrB5OE
AyFDh1o7rYMTYHhyJV0xzTIOX2lQeloWXlmzXoWqiLBdzNF8Oyquqf76jGt1MuBuMv5b1dVi3SkO
Wu5A6chi0g7LR/oiCtVE3XV9SEcDOW01Lbtlcx1pt3mRbL1DlaPpA+V+bhQEUAiCw6NxToPoULba
BgkCBz+uMXfsQ2h2xykqfDWyE9ZSfsmieqxFR5FpgTCrQb96VpZD65SNqqBCmCK0worQTx0iOApz
/OvTQImHaDJWNFHif7SdQPqjAJV/oK2brEXLO/x7j7aL9/JrrorYUQHHZ/7QBl+z3UlOf27hcW5F
8pQ0g8t/6abI0FcioLgi08D5nT+W51rmeQLoqgTM7E+H5Frqi/PnQKHvSPYoli2n5oYZ9lMHeHNF
EoFkaBixhDN4326VDRPAIVjZ+AQkfG5Agjr+MvNrnJQoc33zjp4Q0VoAdsXQJiPCNi4PPseve9r5
GhKRDhQHoKKU6DVTBnVmsp1Etvfd0L18Fx9teTZGtgAaWSp7DEj5LIy1QT0L5oBbjRorHLAUwSFO
8PoMMor80cjWSKIsGXt1Es5C2qs+Xs76wrWZqAF6xJRfjNqsQ5ue+/DoWYmy8Bb4y0Xrppo/+zp/
sdqwcmbLXpMSmHKFxVkK81I6PtQ9koUg3d5QjT49FYAdVvGPJi/MrJqAwOvGQ7ZSpbim6GawFuxz
qcQF92EJf9meW+38R16LpKuEo6voP4dL5jasa/NmoqKs6yQVnqholkK0KnMYdlNU/I361h4MzMLg
IY+JSN4+QRQVd3yvLA7cZ4pdg8Q7kDjOYn91MQ8xyNfC2pBbEcaweNUt7Fxn8Y2YclFvtbzLv2T6
MEoMkaU2pEuJOKDiSH+/i6UenFqRUdFbBR0U7uZm4hnrTWmml3v5gKbdDPR9Z9XBo8RMGVHt1Lye
sk9JzXeDABjMBnZgQ6q+pgFeXM9JVTRcq+2W4UZ56qKQl9S86YBispvgwbRBxftIXqLxnnmZ6YIb
VSMuHG3UAgb1fy7vtVRR+q5HwzpklAMH4cJqwjq7mbFhS+NafIDSP5A72E36dMf1LKvN5B7UazfB
xggN+HQvMhJLOWKMMCDu7my/ouVyKHLug201CeWJsgsPWFuT+W1u6RJSaAYMx1xRjIIGyHgnnWXf
mfiIlc0HWbqPXHU+U59ODhR5CB0jq/K8GykznThP70TmU23NWTGMx7PDAfUskq+pzRtGOLka9V45
T4OEWIKeF6zv3+/0dmX2DPxp3qygXQ2/yHvhLanBk26j8mWMJyDTfFzPb/P1ewKfDheZSMmjdebQ
LhxPgmUSmt9koKgrldcc569d/qvwfkfljdP5nal+1G3dRht+KL4UjKRbvYnu+9xL9APenHDUS28H
TAw0GmiAehorZuYx4+GGKSw9ggCzcH7Yp1DLCGPZ/n7cMp9n7iialrV2nPZePIzz0EwkZBWgmpTb
VQoRD8K8y2hEL1HwuXRyyn2/STSDl6bEDMg9lPRtPWwc7r8eeTB8LXWlhZab0qNE+EcKp5UGcRqR
ZKsnC95tHW958K0US2C0euBVZOs/ZfEg9Ak9VLp0BrjNkvrB19W9tsszIhq7zQds6/LKtmPjQiY1
pkyqHuo1z69cmLw7XluSu59trOpa4OuU9JytH4lot71vCjxq/8ZJICLRAAJOEozp2xmnv/tjZQkw
jRRamv1uP16os7NsBx9YOy8UQJHwnZn1UhLVdVX0KIaXHiRMuNCUJjDe1q1uXUMOGO3Ki715xp21
n6u3fEC5t4UqVzSnWAIEqo/FJLt6H0Z4YcGRDdtHkLdA/bfc0iIowq4eVuh66aQJDsxlPhOIuicz
288tLJ4xFLU2gjRaspw2OHQX91PEYgILP3dwQjk/NtqYHvTJSVQEmLdVor2rj/ihRl5PIGs581lf
nFv4XXRh5UgSkIhh/RAojdpUGuHmuNYYKgLUIK/7Z3XcuA4mswCtLHvyzzGCL1U6JQXLflhYwIUa
dLr5LCrvPxVLOpEGA5ybcktSo6pSrrzS2MIfdMrouxlwEs+bePjBpo1n0sOXUt+Mw87rRgWqw9XX
2SANVLzs3jzBNlF+0QWD2rcn5o4a99a1tZ3xb/ZbqgaK1bKmYxAN8qR2WPDX0OgolcW0rC1yOtu2
QyMJmZGXW8RVgW2s7qUlAG/DcYwxaKep75Z8e0007eCgpOL6v8T/9LHjNfNl7ZFbjaIsVNP8jkP4
g9FBESEwwnZwQdmRu+4Y3FEJhjqsn2f5pr/hXRB5Kv37gonC6tMefXWp/1nINBpRpn4MhwsihHiW
K1FArMDl+zi4QaeP2whWDldFQqdjmh2dgp5dQN3l5p21aZ+ZVm4OdJWB7kH0A4cHrPHNZv7eenjg
ncH5OVRK4AbeREZ43cRh/ExQC/fj13aT/nuoVD5ZClo9a/ERow1OY6rxbq2SA6b+oAaGuNhJ8tZb
W8BXYWAk11PB2UwGUQ6uzvBWgCenh8U4RiXnK28bRO9gOAlG6SOoiMnuYuVg8BfRPJ1Znl9btDQ5
hHgRWbjx+HAkE6CCMYIqZL6pTTnduJd9gqNj3QXWY3MTh4ofdsl725jibliHTz+U2u7ErXyazJVA
NdqljI7tvDDqeUh44qPESEZEbprJBqdCxYL77WWJ3mMcjO/Ry1ucOHWUm870gPSEp7Nozwr9DC+/
iLW8BBOwhGdepyl8OrYiEg3nIFGWCf45wxIkv3uo4IDzj4st+JXnrzBXKA9TdFZRoLIn9SXOMZe6
p6YpAiuev/hOjy4LZ+F2+P+frHWaF6aTqSd+zooMDNLb92ZHuv/2AONwwQUnJ4asHQCLZU/+kgNx
CX6ROd8jkVFQqVgG2cYOtSAtlCqa55R6KnelM7on3YeFMf9x6BNBijHS/fd9S1mPaZyPW5jYcsi6
DA0KbfOA6nvspLW2U/oYr0pnQUknOKDlwuyqqBzaQUH1IKIfiI/TwICFzNCzkuE2Umad/7b83sao
EI3oOgGb7Q/SBUuh4j8bf2vP41X+JFeO5NiGef92slVfno5HNeGOk8OqsNRKpHDs0h/IJHYt26wv
jJbc203TpFZ7pzgh1xqlbWHVdmWFeQycg4YZpcSI0yFpIpKiE6lp+CglznqDrnpa2wYxgo/2unKp
FcXj+huiswWQuX9Ok2tiqBCXrZ/82l3V6BgCJ6ID65pP5Uq9eZytb9EtElOqusk8iPDeO0WzdHjB
XDlm2B3cmGFyamMR3U30VFtPeH5/s2rpsgb12LJWfNsOgjp7UulaiIwXQdl6mdbE5Zbj1aXPs/z0
qpxLAxInL+/1KDZSneJWURFLI7+9RK24Hyy41KJpqB0l2QEXHbZaF/9hACiwYpr30V1Uglr9Y+Wc
mGKpXtahxYO/P0HLpU2FilgzrnQHXFk8zgeHpXEcYcDExKbwkbcBrFj645MKwQhfpUuTHbqznLGM
yfP6BB4nEHwPRqywiXSJyoRykjzUHB6YbznGnkKV+/yMjwMBSjnJ7GIkLMWKbRqdNLfESw7RAxJJ
g61MvsRdbLCki0CBnglSi2UL2lMf+OcxGz6Gm5Qg9YfCiyV6n0mSSi1IsjifPl7WmzHMzVjvLUHP
5pS9Wvbhuq7Jm6L1FLGLSSkHdvFeFgvCO4OxL7J5hbUTnRftbdrysmFMsdm+gbSQvK5Rui0ldc9V
Hr7Q+UFcraK//q8bD0tan6bdChav8cuLVpHSkVa5GAuo2lbDkyWENn6rrvDEjcRbW0jZLtQ4ch5Y
wd03moAKptIrSwpYt8chIS/y4m02fdzLSKO2KtBttbegLX5d1H272XNV9zeUyhrR8PHzPCOpRKqV
FcafrnNdjNFzELWIbZiP1B59wFgnyFMrC5kYx/zYeGa3JZbFJFB9aIXwd1LdRTmTmnpNdjRLMTxg
BKZrsK0aWgNKE4jOlSGXh0VmVWs5NkuWD1VHazCM9fVdOC4z3tt/mRqyXVJquOhQICnNvaRPDpl8
JuRVJfnf1xMOSaejVXKtgtyA0Yb9Js8kajsL/JhHWUigTUSp156vc9E6WYPj6UJ9ECd4cCFgEfQV
OhUYOGVK5EESIva29/66IDn8dTWlVlc/CO7SN3XDh3WqNHPYfE6K05oqpck/K5FxCbOR98nu/2Bi
uh/rINslf8cszGbEu89sys6IxlQ919hS/m9Ylh1ViyDB3dj22mI7Bd99wcu2AeUBvtrvyD4F6lrZ
f4CF7gphzW1GOAhfJ1x+inxSFfaPtLQ5l50UTiKt+MU+BsbHs3wTDUdLIXiPIQxOZjQv/Js9O7sI
tKbiqdKuQjpxMwkJSD8mu9W5QEsjJykevCn3ajNXZba5JCqQOiuYj945YoSZbnpuBgLftVON2ySf
FkKZIg/GqwpCm9yQr9vmt2MKr9upECyQ22NEfStj1xGkjxTSVeCB6rT93p2uir3DPwtyRPof0WxE
YeFksdfH58oU38L8yhzUVBIyS0X/7Lbw5X3l+mKDQ/KGlc9r+rCUckhUovfV39QhQKHcKlHVsWFT
aUYnKkrmG1jb/rBv8YPx12dLH5mCaTBf28WER09Ls2lGGteJgxZrAHmjBI7JOJbFcdFTmBFr3q3i
gh0AvcSC+3Wl4a1bw7Vrta4B/CvfpGkmoNtRu1zEnAodGmDVL9nim5PqaKzB/wu4z69DIRf+cJTP
rxqQ1HT+OV1eMwb8YR8XpqzDMcai0egHrhuUVfoRQcA8n1Gkh/5NWRUpy5mw13JVXporcWgt/dq/
anNglWgQPsL+Gp8fiO9HeVDvHV9BZUqJ3XTJsvXKIgLoj9r8zqAmeF7fs3POzdvmWKNgXTr81tUK
N1pTgkVENAE5Tcwtfthc5m5pwXglbv0/gyL69l/7QJ0Y5BV/GNMuH1eC7LwIvW4elVVhSMwdAqwW
jbXnOir6BKQ3Qy06D/pdexVN2JDaL/e+/sGy3cWbksJH+YLxVijB8hz1MP+8sHFn6QHXzPe++7+i
A33fwZ5HAVfR66vNroluvMRXSIc0FOlGd2nNIYSRICdebgz/gLzAT4Vbt0BZ9Ct55x3LaExnO4O/
F7pkG/BHToJDJQjU8ae6d+V5OHcJJZHARwxVpGcLsWoJtsSSvOVQFCUpJsi9/+WVG2SXEwW2Zf0M
4835kifmlG4UPCYmfhldhKMUdQS+iZP/8sx/CTAmoKoX5G/pWOpNXH9/7YrXNHsHLgrmzxOsf6dg
Apg9G7pf0DnB4B2jzD6M1tiU6q5eh5zEeBQ5yFqJoT/xxcSb00yRa3NjgkK4rLlJhCOwodaogERJ
wc89ItsPsFVAYwknqwTA3vtjic5QGsGeR/7vOrbaEyJ4PAp27NDJGThctBL1UVlUNaGJGwU1C4JO
TUyL1U8rfivhvpG3kN4+mJIwMJfw9Fr9bkpBIpa/U1D68jN1uVE8QDXOa0E7y2zUDoIkE7Aj6hYt
L3yXJhcwqUc3DkQXgpxmz942qLVi3WqluFRDfkKYGY4WsD3OJRJJ7v8JQd+32hvI4JzeC1yAg1XI
+G3seEgZhuBdUcYpuNiGnCWbzvzLrd0Im2hR1xnA5AyOQtGBcWGSuik4/NT4B8Ff5gmDzcdozbAI
y94TzN1aCTgUe8zOL/rgB8g+eL8jHWU0g4VUvHXfFBItB+PFFrafgzbMxGp9Vs7CG3GdHuLsBcU1
qNHhOF7Xd8qRgqZ0i6WR/mKPlrrN5+42LmQXBQOuC7lv5IN7JW24OvmBIRIQ5F9WU+/QUwPCVaAO
sGw/9cllC6CJd8uISyAwrEDXMN8XGdJAccd6LpIJZ5OvAA52ghmxVfn1qsFXzx9yz9d3MHuq+Hai
XezR3NtT374QNhYJ2TeHHFAdzise0qKEqftiKGPuVXHHRQJ2U92LO5nha6rxwi6ii3H7FidQ0cCG
X6v8ht5sVtYB++D6vCbySdTIbllP4/67mWAZD8I7hIh8kBZKNMg/SMAQZEfIf4TGNOE7R2O9FKOD
b+fM4aHXhnGn/ALI0Pb4x+LmtJe7H01KBT5uD1Hu+POib5aiSHDoaAlTY4jG1p9uea0hcZNA6MKc
kIL90pdtX8efGdqD6GcZ20VgkSvfWTqW+SC8rCz90i2k936Jzr+wk7OAoALZlMp49vujR8y0Rfpl
2IHvzZy/tKzA0VqFBbi/zVn0kPA26WAeXcXB8+NoEzpSv4F6o9SDSNO2KQ+nlgO/s8/cqgBVmmsK
IjIzWFX5+QY/igOL+bIOaOZvPzHzbq0e4IpXk3Ih6cc0nD5CxF5AN3pCfVqzVYGO+JKtfUTAFyzm
hxjsptayc7v6RJmt2mSR1pWH5bMphOd1E6d18+1DgxAHP2MswT2f/BhZtiUOBr6R0B5sev6ijo2s
VcI5/+hAuzDjyX90d2EtU6IL4Zb14QD2VEL0uWOTjJlpDKoQnaai9RlX2GmHbJAdEgSaXuZq0mYI
HQq+HZCYxd+U32W0DihDOnduqR/lGFSRmTQ8msmOuxBoGk4nsFoT+pXrblB5OlgOjCwvA+MkfS/K
/wPpul5PJc5jG7bSrvfkrPX0sHaoYsRYxYPCWbhtcS+nChfz8Q9tuNSIbYHlglyOX1Hsx0h2HM8N
r80vd3rdHfPltUcyXdw1hQTiY5N0yrU47XWoylge7zV3hqakPoL+Kp+ZVUzP094JwRZQFqp/GFvI
SiLE+CmTNmtveh4CSsMB0rnqZ+nERXRbwSsjMGsZCe0MH3oK3kXBaSZKlyE48fuYqT/B0VPbquNJ
CsqkCa6IGDydWabLzg9EggJ+ut+LfR82GgW+LPL7Ae48i1y5A3OuU3J5cDjWaYUnH23h/bAjtshv
fKV4UCrfLCWtRGNT/WPZBK07ql6VEQzgu5MXW4FV03dRd96hIpeUbUJ98DhgX6jddQsJDzxiKsFw
LBlzaMdaWQ8XK/h8W+oV0i/ll2g/twtPI14v5HlUYj/MgqDtnKEK2nj7MxIeKh8Jqlp3qCP9RoF4
Vu3wtGfAWDnT9cBjgjDAUVJTA6i0j+jt0ileMsNL0DsNuTjZxhfM2EPQTG44eqF+2IDfj0FRt6sn
qs6uxONaV2X5lfdCldodcNjfygtC8Qz4gcnJZ3Z6TREwwsE2R83hhcMCy7tSq+GUIL76EiuAHBlp
LUeMPX8eAoKzPRFW7IaTvN/YC5TC4IfrpLZJq4y7XhCAbzzzNk0oT4bxHoF0A6iuCcoyRXD0X8YC
YbT1ZW5Bvmde7jOFhMhoFNoEJlUi6j/LtXNxk7Sy0JPZmCwKVicOjgnNTxUPhud+pBULmRXohuEV
dMqY/xiHChcWNVauup9YCorGDnEblO6eeletba0EgTl+Yx7PSsMv+yYpcNhmxDVVb1ftFj524VE1
hNDPKTPmTcm2Ioje6/+MkC2L7FstO5Lr74YlAGDfvwxxaEd2JPW3oatzq690zkpnArvdrIM0k2KM
jyOd1sgsOxRp31AMZ6JDSdDDVH2EPS0Bib4QRBWvzHFeHvlE/ViJkyrCEykiaJ0BFNcxLGbyPYVT
lco72rbLoeUU1CHUIhiehvgrkunxLyQuWwN4C/ccMc31uK5UHc9ppzgkUM6enSazmtypgQJmGz5Z
nE4kHWNTALV5g5Dc6lKZiC3LI2HayIuwn3jStpFcSueExtuB0qq6PdtxnzcFAKUTJ067oV1yktIN
D/s6LH4X9CqKgqtI/6aLLEpEMFEvqTsM7b0+77Mdda8J1tcaswMZnKj8EDaWCqdeSMNyP6ol7KGI
Z1EjrYkrtT60KzZ52ZDD5mtMF7juy6rpyWDYdAHylytTnJ1+Ibm2b8gUouNIbaB6GTofS/iakr+h
9ltemwPhy+Qz23LbmQIsjMj0WvS/0YJU0zHA1EBQG8GgK1jLvbzSVyVdUlL8E6Hegnt1iQN+2h3b
YGJ8KZSIXmkpl18/FAnXXL6yv3yZo8rXiBP6xitT3SIkFTkf4o9S7CIrJMj5CzHfV9OXNFmHk+Vw
CZyA8XaYIFdQH7fC8QW7p1sFeAK9Td/pcRp9gdj8t8IKo2skUquiVZM7b6eMjdHATKPYlE8zvNsh
M3Hp3qx0t3PGPC+dQ85cRQgY4+1qJmhfxj4f5YfPJvUlrsx9g/FX8d39b4vpYKdjRKmV28gmx+fe
ofv8T6WX5xSZJuJDaLZ/P6JJsWuXbygAE3LTyGtow3kDfJ8hOTk91hWXW7dqcJ4aay0QK94NBikY
TFobd3zPkh39d4Mgp5zKrV3WmnljZPwQf7sey4ZCISh/WkGQTDzpxnM0s+5H5iDv4QAe5YO6fCz/
RxXx6g3UPwe6l6gKlogWJklvD3g5rOoMb+TzLAgv2h9d3a0BTzKggoJ8VF19+a5B/+IcZUe4TPqL
oL+dalUapTVCb9oplWXGo3EzhGBC5Zjcru50TlggWHIWzQTDqQneK1ZGJ22LLFol4KXZh6cH0jhE
nw0F9XdwMTj4NOXFNJPFTLJHkdUbnFTAY825srM7VFEQsBMisrvIDYCNmTYzFxI715keObSVwQuk
irNCO01eVL9wldKty+Xw4U/YNKWIZ1QyPaXyX35XMR3BDehCF+UJpBDm5yMH9RlWt/cqms+v4xaJ
kmfRaHDfvcL0PC705FKorbjPu32En0w1K5AbA1lMhgAthB9o+I6+H/fnT98tKdYsKVNrsJXewHZH
Dq9ROd+xAtOqlnIgkkXjpzwGWcyODRyAi2DhrZHzRvh+Mlq3P++SEH1RtzXtpT/7rMTP7mslCQGi
/pl2CuuHE4f7tN0guMm3PwgrHiQoQn6Dbs82ti+4HrY8ciTG1fp1IN6IrigvK8CV+Z50NOke2FPo
KvqYY632+zNqmwiVa3vzIfIT97EP/RPt57BtMfFBmm0zyawSqkSpeB5Suxz578hApfMv3USdIZ4+
jyzBKvIcUXSm278sdV+GQD29NFsgpm+nd6OLyXwoBP66tZohxChx8nGAioLP4jjpuIrbrJDbEJb5
1aqNMav3D22/xFrPwMB76SCRZnja3Nn0W2gHLvMOQwKg4VzCiZSqVwNUXcYr4wD8DOkBL5+RH9cb
DjB4IaJOTq1CAvND/2RMnY8FhgX/ZSbf4r4+FVt2/0lb/GSpSwGnXGeGroSL0TrFi+CszWoP82OW
Oa6BNGaD3C7XzN8fvPhiob8VMl90X+olMl/iONZO/evw6eID/EK4+NqWHMY1DoF6AW1nqfimEnFk
wy/rQLo4L4FPdd37Y7k3xWEdlW3TEkYoEw6wDP7bu+JfkBFQfCJma59ch3bX3cNr8hHEbjL5glG7
QLTPUifbqGhhR4cxUraw7yUsWt+q5YjV2kCd2Ql6CdWaNXBo4Cqe2iXpAqIGI9ziqnZAv0tbVyAz
QzazjJmnd+OGt4uPufdcEK8CLeXFo1srJulmJPekU8O4Je1hYhGTRn8aA6JBolDx6IKhQdkmiq1z
I3YiwDfQXCtMw6med4OTsAXfVKmHwXYPRhGrbXqrFO4S1GsOVO1axzNsE7GjO4R90h8Jvyh1O6sy
lmj7jLv4paG5nhujikms+GUaw3PCKxPo3uQkEKxylgV0DMf9AQJtA39Tm/3TfB+axuHR8JFcnNfB
3pCOp6jmJbkDfgLMY/QuP7f8o35I6xH7hg75CnV61u2sJVJtivhcw4BVkX1Ub3HweOBgBn6M9g1k
6pgNeuo9AM7FFBffBBQFKtGSO/EYB0jH6HcZDIvDrYARREjJLeMndwBX+eNsBKTpxwhQjEos1K8X
Xo7vaqQQu/GIxIn2YEMhlf4ONPtizfFSMQhILGcsd9w8CX9WUC1wAgMml+OXaC+seeQSFw26Dm+O
d6CQ6Q0J2Khf343eAd4+bX/VleMf6oAp0tu2bNOwC3pS9SfQmCuJAfrCm1RPDDQQtBJGqsJX+wgQ
iVUp9zLcdQcQVFfrOuz15Jg6zea4UTqzaZQ32PTpJVW2dH+ZCtf01gNBSr/HZHMgRo5x51aoS3EB
fRBo+SXLrjX//+KaYBo9SUqU59BKbnWF9rH773fibqn3jFyNPlhk1Sc/mWASQ2bHOBn1hoFfSUS+
vJXOaiJRmqxejRFRK+qrSvnE9lCPYd8L0tpNUBHvOTvdL64nSsa3xWhBOxqB7fkpyzBlEtoMYng6
EXdT4VGQxC5gv17C6qHr+oBF6nhSBcR275j0i/b7Y7iJjMKjYo4qoeRRDy0xz5Mu3vZJVZ8JBlUC
hyO7YZefqyC3O0AddDiwrniRlCyC0U3uK+h6bYkJRGs57piqV7nx6blhOazt/LnWngX1Jbm3SQvD
ABbKI8qYZdXwNNqZyq5uQa1NMRpxaiUTkD6edmTWeq6VlzIgk54Q+KWkwNNWrfZkTPmlViUH7n5S
g3+eytybfgtMtbStVg5G8y28mFhR48jVIWKy6E4F1agMdxLwhyijZwb/q+3BRVgLkJb9iqUj5d9w
Iljbladwj0QRZlotJsPp33frmSnHnKVphDalZeqLVFPKuSsrV+3p5v4WpnWIKJ46Rnjp3va7j79I
3m4G7xFtB2sxZWCp1gwvZ6+VRzA9JURLwTXacTYSnY3MLnqmYPlbbI8ViZYhteFDlU4m2VJ8V3Hh
0JDkHqKkxvveYzJtzvRVZ2y8ZC0o11zuW1k1XQj5SwOpMSD5ajusQyZO9iANGTmY7mUHFaFI3g2n
aTHK+vujqiMCkWyIikbkfey+wW1xlJHZ4bVgisEMJzpfjVF0iQB/DG6adUQxEgWmoOORu3IS1Cil
pUZn4ccUs6qaHv8lc0xO6uhWhXOCKFtBgLyRPeD8jvcmA8u6tKokHICS1HH/mB4hKv3CQBWAG0W0
m1Oql3Kp5zPr7zEY/Z/BhhsUAciwqm8ut1sbQY4bhCuUwNlG37+SEX19PleYJsw4QJY/s67MFCKY
zBM5IGz90Td6sVJZJwM1McMVZYggZw+Ka9NJ2uJ75AJMauYUmycv5Y4woLNv0VDk1hGMGJzzoCi3
dwTPmMFDvK9ig7vOtJ6S9tUUAtHsriMfTKjMCTNYkgUrsj+v30YhNgx75zEpZwC7ylK6oXtXbYZY
ee8xif1hHWyeZYW0+Zu3AjCI5OfFH5y+e7f9w9FQZvfO/Z9uvMA/IVYv6nFKw+os/87xhc+MEFZB
kylU1F66+nwNW1pVxQHz1jk5Mz5EDn87R7xY61ROt4CVSmiiywFjZmvw7T9bdB+umF1E6b/mm8NV
kfHcOKHdG2Ur8/hO5JDKZixLx3QJKWpCLSfjLRlLLBm8Ls+QfG9DGj+VqNiA5ajlGtApkd5m6QIc
sGcLnH88HhEjW69BlqyU4vn+ZBfHM+FhffU4diXSGPPfjh2GaOWcFK0a+2J7TsAvABHR96r7DhVp
3TEzmUQcfgYQQja1btzSs5U9qyxznOj+EcGRGg66E7pP/sqMLJKgb2O1QGWKxx4zM5CJtYnxpohk
qVO/E+S4zr89dmXOpgrlgnebsFD3CWu9bMdiTbny64CGgud6V+zJfLs50H0LcJ1D49yIwF4Ud+to
9C3A4Wv/5u031o7eHJtNr+lU7wmQezWdEgWb5i1sGGhHgSpoC8UHDhKKLnh8LTOS8Y9Wh2NeodjK
mre4xB2aTPHO/DzDTGY/h1lzu9H74ilKQRjnF8CphZ+RfHSy0S6DIskpuSZtqQWRDFOT4sGYv7EW
dkXZj6Fs+Gy1YxE2np58Q3aKysAgYV2TjjiCAQIyaBRo1xqPZEhKJLaAlxlp/cVQTImLO7OK0ymR
Il1CwTrTey+9g3HKMkm15va0FZ78s9ZGs12gF8foWYkSbV2o9QSTIgoA1aTasXLOz9WUDHGr/VzW
6OsF1Ky1B4TdYkzQvKWLJnrADNrT8galnglO7IqoFmwMnRhRzyVy51IH8Dxy9jT1jzPDTjjCeUeZ
zl7Vo3PBEF2I5hHo+LEQNHHxijGF6g8l2Y2mxsOleQbvefsQ1M0ATG9uAaZet3vSRO91xtuCMTk+
ARy4/k3ra5GxaJ2m2r6QHEOsL8kw8pMsToAVR1uZv9qZwPBKmiwxocvu68ojgvh9vmKs2186qa2m
3dFwzyr/98bUSsui0+BYegyxac1Ymaew751LTzBTajfR9b5Gp8B9TPZVaiBM5s4IgpsN0BC4AzDB
OKnMXIkeLXGYpMtiGjh0obnr6aGc2d6nCf55/3AvY0vx9KJ/Up8TgPt8ysn7Wt3ARMn83tcthj+I
j0qTs4EM2dIoY8z9A5DAUUTuelpFhoel8Wl8vGH0irihRz7hYZ+NekXUIeSWGiaEhuOC8DlikSPm
YGJbENCOwrFcL+/zBZ4K3JW5brJa30zJo+HAMUcGajosR7u6K1c3I8zIAj9zyC7l5ozO3uWV66fA
vU+PswMP5Hs+4c7HULDmmKJ+eLPBYS9gKZemOfs3suFlh7tBh1kuYCzGyPS/zWc4b3Qg9LahDoE+
dQIEBJmK9SZl/9mrXYaLfuoVBhoCXRUiu9n4tku6SzlHrImYHGG6HksZKaPc/wvZvRbsOUVPEyII
MGhZV3AHDcPD6WGxSZCYYNucds8afVPaeK5a5Ss1VYNm9rYf3ODz8xpSKlwUD4v6pBfjeLby6vu+
V7y9tvgpXot61ve/3rhkVUtbAZ4DwlT7XkYswEp9f3PhYAxKvhJD6aCOYIDCs3okZ/p+hWFFM0Nv
HmLKptUx8QNQMkop/2zzVZlAVR7pK7/svraofz64QwmlVh4TR65JRpCLUhhHOCYXzH7sCTAp4g0T
tdknEvnPWiMe8os5+LAImneUrsKEnkmqCrKT1tFrYFGw5dJcAeROkel9EmhRSeOm0JyjAp24NyQu
NNjAfXIjttibTa0Ir8KRY+Vk8ZOd1MCxo6Ejqn/AngSw2HYlmw6JtGk0Gysf3HZrBAidMntHyMPI
qIHQgVkET3Ll5AZ9OGdB/sWb59DnokFjNIkD3wcKjSYQkl87d//2sMvUwK7rhJ2ZVHuPfud6VA83
k5661Vkxx4JwgBvn2QxcCQwo47sCZVu0Fb8xTh1EDqRB5MnQhOKfleQVV82ktsBYX1HmofX5ZxUm
ZDcrmsfbbcCUccOGSRIFJ7pCNK2mKa/cQOHac8U2yiPLjSy59t+Mh4cc/YlBDCoC5dKktcmbXXxj
3OnS4qdf7zunxjP2i3iRRBt5vOOYVSlQIVJBg4xJqlRzYFHp7ZcmvU8aUHx1d3AswLxSKQygsjHA
KNdgdOSfgtTfBpVXVj+/yvCPpxv+EJC+xxvP9L6riEqoL1COVgtKtAytmNMbsR4t4CCrLKc2CG99
qkZ+c1TqG4h/8u0MRoUt7/UfT2YyLexvyM+qbNwXOxEW5QcGjJSOEnDL/Q4gwB4XYpxBHcuYg7V+
Eq2BjQNTMgBZ3FSdLAdrA4ddn5MRNthw3KITCjgpUY3Zz0e6bqy0k0tbbPApRzr5QU6+YG1NH7Og
R3TXEWVTrLZlZMv92uXTpulQpiY5Zt3r6xw8MRrUZau/Lm4EZH4rHQzYfF41+RsSnIIZfeGg6/Pg
vmeiWr3A9Wh6SN4+aKac4srrj9t9xQlldY3UTNfwb66HOGSRx3AseN+xbQcXnYs2AsKH22xfOxng
GRGsSWsHq+ceIY53cvugqxe0kL8I1/5XdpUsawb8L4NSqknOjjlB/ojVZ8o9T+J4g2gDhGaNzSPV
hDNupbVP3HowZGhSBHFM8qJ/SwCmlR7yPOH8GVyr2ygC6deJYbSZoD+mr5vMFvOnswDX1ZRBDkLM
5mSXecehMSHcIwOu9ulq2XVzBBxAPIsus58XKuanGJ6RC/H8C1tJtBUstUUvvOiEdNMicOcYVrFr
XKlrn1stJF3YgnUBMpyNVGjDvB6bcSyio48p1kIIUmNjMeJQpQBy20lzh81IQqwUsRiYPCbqhOh7
nHEg+SUWSl4dveRqDVNXpFnysXpxwcJiKFtsH8BZE76q2/oMoO5MN0h+sjtRfkWiL0hExDPHony2
4SXPQmonRjE9ZSvqkZMei1YMP8f3tbcGAX12U02DCaxWZlo/ol3KwNzHmHNDGoAPwZ+13hnxudpQ
KQftdZyQM2fUTu5wYj+ahRX01CtyO7+6age/S6HzED+pvUox+OQK+QMVuNyMqbAQ+/lyFQKiv2q8
gqUVpQmMvdSAj5FlRXvAew8hKGSXIC+W0coYjEO4RccVypPfgMFFrWYfJ5ahawAcnWjBYr0zVTRc
rn+rLY0V6elRtMOsYTVPO7xx8/Zzu4HSoj+YD7Jasz7e58SW9iyF2UZrwI2WvGWLvsgKyTBi76XB
jz8YRGdhCMPjJD42nKUjWXmsqESyFQSRQzmty9H85fgU9Jz587NOGt3+XxDWcom9Cn1Hcc+hPcgb
j/gvyhx7AiRdjdVj3lCVEw6t/OM5kA9FCQQN4bdnmJPJ/vJzTxLtjEHLxT5XIRPPAQOCGHPASsM5
0HbZbZEcUy/uXUMDZfwCZKO26pu7noYvuFnvXYlwzSuESAMstPX01o0iLmGQKM/oHHscVEszNeoJ
9FvtiuSuqh0K8E6FTCww4v45V65Mtppq+ya8BDa/VtJeYe0YezPzkiC6v3AhI9B7yFoiqA8ChkRW
ueIKjOOZUsnP/JpKiLAoAwmL7D1bBBJvBPYOeVcCqVI60WVLjncaiFdDjP9X8eqnD8OPdjfTVboJ
G6+L0y21gVQlYEKZXEDaqhK2vD8W4H+oKf4X2GfJFUo93nLZoRPVtyaIwPXpAr7g/fsc/MH3F+EL
n8Bqs4pT3m8Cw0HlGkTuRMqtTgcg39YT2WW4BszsGEpOgo8UnS58hzkPDRtYtpou4pidEmGljQMB
96oh96IlbdLWFeKpNf01cBMchwDNN1NJbr8YMF/8TgVbiPM1vgAEbcrdt8N7Hv9HJX5dHiwMt/wK
qw1arE5GzgpqG0ykMBkAF3CXS7XaiufkAf5CCMKOWsJnVfMOIP79sfXl0PcFrbUsvuY7wM4dGZB0
IUbx0xGpzGdX4+nrW/lxtaheu96uTu53PJBdIVjxQqAQbUt17WAWgVzXnvUYKjjlkqIgSJRr+Atj
or+mA+w1X4ApOMTm0pHnkD4FGYdIMw80/kuKtkMEcgQKqeioUiZOAl8ABUxm7saH7LG/tBZXxrJt
D1uxL5qKzWhaJ9JNTiD6320ckPB611+z52jHLBu9lU4mmd227aEEmLicFSf03hhbBcUsti1bbsKE
9tf4+1lPc1PFwHmEX+KQ7auPYUKPse2ZgpomgmzTumDWavZZaM86asm+N2FTkHG90CimL3WVsRo7
MB8oRZh9CJecmJSEuvYIYuv6ew1oF9Wx3+utXCVgcQGzXFKPARd2JbQUeFeFrFemiU89JfNBS2YN
dhkWJcz0SouL3oUQVKEYhcVZrHkiLs97ZrqHO5Ao7Nr9AU/t1uvBXaIhdC1/bB+MvwLvh2/gHHxm
rUDhMkiij8u3OIlP99zzlSX/x40bLFyQqpSUiNVknoagMKnvZXqlvH5oe+xAEpbi6aEeFdkKcIhk
DxVyFyO4ybGCg+OMRG+QsO/QOS4axxNyaNCuLcdjrC9TDgn3k3JyQmNfCBOwwWlJmxYe/NpQfdh5
3zAfdgcOJXJ8KjW4k0ffdAMxVm3wn2CrtjcLDMbcoI0lHZflOehkHNg9Ui5KsADqizmDLEgu/Zjr
4KmXHL2XGl/M9AcMHf6NetDXQAdFYmb50peueRebYPI+lU8Aa+NnYu96GqNMXk9Jl0vU7UcdJy4v
3OxgfE1iOu6P3+GQtAPFkJ95aJuv3dj3c3PGtdDeBBuRw+kCXwSnTFi3z9ubFWhEYb3+CPuU/K7M
5OGn7VE60W03G5rP5m3MFYMYEOBtZMY7qNlFEa6fgColVNrWPEZEhWa7MEj0g8hWJlEDm4/df7y0
QEizgX8Qm0riUm44HUxs5FWGMi/g9xqlF6dl3RiG1ZoT7Gow6R1lL8fsfjQs5outp0vTXLN4+4/k
pnjxHfZ6M5tcQgRqgpX+MnjqGw2fpVxjAAshY4Zk1ZcJr74P+DiKdOcWPu8uJvMF9uB/M5OqwqdO
ayB+QeRRLNWfVfGtNkRItN2n64nGF+UjA4VVkLXTOhqyCT5nWPZ02KmYHYi2S+TYWJO8rSReNQhC
dwBzHiqQC57WxK7kA8GhNfVh2+ROisDUjrAZcfn1uWctXlvcc92ovpd2+aaXvoJaKE4dl6+qc4rN
ozSsD2V5W5UNr0zYftLKvqEIMt61V+uvcNMWDMUZ41d/G/ZL6fnB4j4Qd10tIr+Ud+F86Q4E4TAK
/Qn14UlXnhW2izMniibfHtoJpPkmsSqanIPr0ymn6/hbxaKV4Z890ifkvuvfXk82Uhn05Ighx5k0
8SalE/SB3AcdqbnTiVofHARaCTdUBXO6971VA8Jw5E1ZmzqnfG2NtYonmsIgN52SnXC2fkHW3IR/
WDpBI0JLZ65xcD6s0VJzEULgEcvOJiadLUSNvFujnsvXl7tNJX3LZwaxd8FxF3WlxN1OGyILzHZO
Q0UdtxAnWR8OARhLWYlHp2ize/gTGUcNuNQGh6Lgz00B/ONLpLo6DE7t6ezGRrXbUFSAc+iO4Xd8
6K4pKb90xepv/QCImbvabgIWmQeqd5YA063r0Lwckmd2qJyyXPZatv6Dbnk93nc7y5ch4dj3Z6L9
IHy4rWyHzaIru4dA2IZA/vzkDRNJax0kEhuBysj/+oiiIJncGdqPFKgd9YdAXKxHsdCEgLIN7HQE
qLM2SFkroM/Qf195FDU5p5UZyKf4nqCTm0tt4oDSN8dzcxw55+suYI35Kklt7thnBie2z02ymSNK
m9gViVcX+MO8/1JCLUGr/lQFBETOAQg841TtLjkLrBhN7hMF3orjD71QI2A39WuPv3LylS1y61J4
2FvGX2MVXK8E8x08NiTM9ik3rs5y7YtDMGlITcQKX4MlRUhXfyeqYSuewWjZPSha8qfNSJhUvbSP
NpG5gaG+5nGZdbfI/eN8ZlkMHIdmjrGvpRBtbk/fR5tWy0RYUXZVYvjnXWiUIPGf9j3zcblS6k32
K6Rr1fVZqr8vhJVfwsvMylkHs1AjXNgw26dab3C1mIljhVPURZK8h+aufO48H3//y0SkL6vT5a6a
TX2NXkl67J0LlWvHVX4uPD3Q2WMWImdOZPLbGo44aCYHAYarwZpsM+m4XOPa+9ndTs7j9iKO0Two
MF6pp1FS20R5NpqLCNig3tmPFQYkKr9wzMTcpfMrA9Y2IvcgV4eh6qVLcMGIybofOD0FVO2s6NYB
yH2s+/1xTZwdqK1VLMNIy0TZax944qNvOYFSdB34ImMbsKEiN8I1BZbdoKyKOsS2ie3MOPXIfZf/
GUR9EzJfIKnVYtzYYbN9/A03hhIaH9z2qZDKBro1OMdKA0rvhvrIObwG7JbcTYsqLQafEzs1O/XZ
+UV9I8Cyf1AuNbfaqAuqEpD0FCYK8LwbykZDFI2iezYcgR2dxIQX7kVXN8hREFSL0ttK0RuivU/q
WjBAm2ASWcX+ai5wLL7GqGIPP/dZnodlhPvdZVUW8pkiBvyvC6Rk2CZkHITzoZmTRKrXFFl2Bloz
zyzkjNzdIORZOe3EEVWncDvmxGEoMtD+z9BsUq0a/vAbB1Kt8OWXdBs4W5MDd9y0XUtIsRQvVqrr
VGed+LKWMilPqut5mM0apoN2JJLPRvROSvfyxk6CuM2SK0gGjPqPTkYPVAr2u5Iqx/mNb/iyHjOC
lB/nklDgRjIJXiGUUVzPo2+KXpblNUKeTjnSE4eDR1cf6hukPDwmf9EIbBlS0PgtYHqYE6Ub7PSK
ceTa3B5binQ9bfwbSjHM/GTqV75SgkQJpEM09Gzq+ujvhd0dUL5ue9IAd7Y5ETZn5D3SeLegl10r
eNm01cYQ4hTjrWzJ2ZMEONxEdfc5Msw01SXT6GzTPNLj3t4s7f1qlfcRWldfeFsWNX57AII+1B4y
GcqYdTxfMUTLwcEwNIk3wkFe3p5yMx4XuyVippyEMH5TdvcYPG973PVGeHei9KdkA/EklnOdseTw
TIvC5vtCg+mcitH139cPJPus+d8tj47Gw5okilo2njc6HajOYwo7n31VghEoMLqHXvESkEQ7ErRk
QFGSU2QvSYaA3Aat7B2iEArc9h6UMXfdeUKvZcwYvSPjS6qOc6H2/eqMntkn5YqL+BnkFqkS8UBj
rxVeGlynZm1RNSqqkIsEtfXMZSFHuUyryu7L/x12wQPkept5wCHPCjc8nsm9NoBvptMYJ3HpalQT
wbvpPzxsFspNv6BUXzJWYb32+DkQdo8zzSlkFcXmypiweyuLNylVzryOVPpD+ns3zjU5jGwDNepJ
nRRQFw3PCwKNhg6xmjCq3K9m2fQNz4Q/9bUds0ZJ/frmoG76I8dOXe/RfMwQ8/eS7irtc+PtQTzg
SJiq4rd5L43k2TmhZ2r4piMe9+IHXI5yTnQTHCtGCD5aykpiCS2OjmdgdAvFbK+8TBxkgY9Qwd8a
S9Y4rU64biBEENAy4ekpiuXkCcX8ZwLhtwPI7h5vM+dOA6L0oblH+CKXvUugSijQYsx/eE7aiHwK
TF6lZ5km2cSDRBpAZTKYgcvKJfcmCTAqeVN1USZkLxdugV9N3ka5YrEMt9SGpiJ2f3tnvWb7tVyN
KtODD/PQwBbeZ4Xhn3rUrBfVs0vbQbaIKdNgN/8dtZvL6+zFIZhisRrFmKmUSm/tPUSj6Ut+BnQu
c92+OcbIsWzIFYwHI6naG/Oe1YDGfSti0Yp1AFEiGOYbZq9mDTpjbk6F/AVNC3/zrJTbz2zoxS+H
RpZZGIC0k/br9pfkCDmFeFtzIuVhOXKAlUuiplXweuyUd834B0jwF96nzVT4mx1x84+60YCly5cX
e4CC5xb77o0+3JphiSQ8jur1G1+f16RA4dsonrKVrgulE7sZVwKDaIaIXMcTILn0zEhwzxA6sXJA
fxAAcEgLbMG97IsUp/L20PQVQ9AeiK3q2lFgRmquJoMt5krXaAUOW/94lRWmGANB6RNfuuJGVDR9
BRNmXNyjTu+rh8zdBB9xZg0P4PjdVqz7yv0tBRE/QMSNGw2/BQSPiRzCFdKuyK3WaimHlmHhykFg
pJ6ajwaYfela9SGf2hu3xVWIQnsFVMa/0vSNQoOEWK5gBQ/zSMaFXYWOla0TSW7El2jbR+I2D/5b
gP3HzvPhhP4XWlx3AxA0kczJQaJU3hqoyBX6zY7Qo/pf2sQBnVB6pfbWlDVc8mirS7z0gIIbYAun
W/mwbb+LIYNvXA7qsvQuLV8Z03EQ/G5zdjZMnIEqJBtTQFmzkx8mvPrJjec81kiJ4/stwYAxK+Xk
e+BSz5qG5HEV/j+5/JV4gFw0mNdeqBU3urD/eGsDufzSayytyJkcXxQ5UO9jtsvIS7YJE3Ki2V9b
ap4O2rENS5qcmWjlAHYx4GiY9Q87IM/uX7tnysvdmEhtFyP76NH7p8A1/ozg+4kwbHtJ0B7j9YZK
sKQrI/OKK8JVRap14LBJQVmL/MP+eRyF5csGB+0fVZoEhtlrEYKKBfv1awsCL1pT4tiFJ/ebA3H5
niQ4g4QtTuoJzXQzQHKFofuvlOW4AgG3uw6L1kmPDR/YVHYy6PWtTUm/EVm4ZSpcJyipXglAgKNg
OL3D26AFfAkFJxDZYHO+xplfZyrCk8Sh+ntZRRC835ahjRFGjES1tJs0HT6IaDFXxE7ou8ae9CTR
/kFJJO1SD4evCOjXia9uwYrXKvYJWqfzSB2HC2FIHII3civWkiOHRlR7zW+eIPlePRlRgLesh/Br
c95OYSaTJ0vDXCheOr1Ae8SJ+BFFPG0Cn03eCll0d/hO8RxHSlPOLM+JbrG2wFlWSIWU501fS2Vc
kK5Mb6ObjPplbZxIo1OXyPvAhgvbTlWxCAsf5/e3adavtzLCL7w2TcnjDtpuXhb4gUbiLsQLDE/h
A1y2mOUYJxdJNCjpzv9mwfB/rEuLjMYSIN89x0os7sDwhc2PLGaUC8xJAielp89OMji7QX4csQsq
Poh/xjVBnv/lYgk+D7IQ78xUKVcv/GHUA6rRzTFtS9aOwy/55kM7JU77OTqWlGQ3OpN/uNVLWUbt
jXUAwIWp+EaeiaevsD+tvy59SFU4JVkPtnHTUK9O/rPyAjKV7SFbXfvSqqAEEUBK+jBt1eJ8wNfd
9vIWzLf4JZTGygQ3wk6+slifY/Wbkr9cNcH8Zbo4rSOg86WJWwrhVNuTaeRyCDShlTfPyz3fB0Z3
7fJOxZp38PIA+ulrjnpJh9RoAYTG90rE4ozWcyMOeHnoQjaPpjgJcs9Jgvi2Y9pnIvVG7Z5+zFR5
KIHHDe1p5u+I69H9e0Fd0noNIdcnZnJ1AcP/OL9XTLi1MpN0f24ylkcXZwbZvjuFBd0SywFzmifb
ZUnI4dFy5jNaxJolHeVwFQjjdOG772Ja+GE8RTgh/BMOFNPdZoGXpLyUka7uq8Em9HBdYqAKerfL
lems9+Hh0tNF4fd9LuY4UnAC0n4C7tqgWheTZX5ZJNYqtW3rZhN3FSSKiAaLjE1+XXUwkRRw+dfM
/82o2TvzAKCgcGyjcTU53xHKpOHGngL+/xxI4p4BTsZQPmpgnfRBb+n9vBTtdgzF83HNdc6/34T9
XjILG0GDQX2iMkNXIvOu/JIuF76S3+KTbz21S+fR40j4FIxFTLmmJKtkCEYPxyVcJAeaoECnumfd
mcZMlhbtqqQu0gs2q04ZxdjqYgcfrFRguCJwNyrhgLV4TtNxoI7URPfTcNyq1pEL7bUkPQOD/1fY
ZWtESqt2ho7M4atz5f9Toi0RoYgWWy5r/8Y32LKQqiV/AyS8WP2EOJ7RPqOXBEGA/jWJmVgHN0WJ
Gmou+zMHgQCKhFTCxguRMZcKbLjw0w1defC9o2CXPXH1W31bEw0eZ3Kg8kNh9iy3xsLYZZVtHZEQ
zFdqYeKZGALqdiD3NvdakstezbvSlCwptM0WmPeAFDFEQXtXoOKfa6WHVnC4pR2ZUZjg4qApxna9
DGuUKrvhXTQNqcsitCR1Fxc+dQH50/FJOZI7Ex7rEeGzMMC/I7CitK1ul8Hi5wtBoRfyCYhg6SpQ
JZhR8lhB6G4r49mqSJbzYC0xaXN/4NZ1cmrzTQ57bNlcAuEkoAXP9uWZoNAnPmkJAVTywqzH/V0W
FUppsg0okNNBrW1wykDe9CkAreQcRPxYS1qzNf9KkWK/1+eii1jfnMACgKPxBL/Ku6tTt7DmapaM
KvRDQg8IJfMAbwlN4HPyj16S5tQcl4jV1km3zBGGf6pwM+hew0IkzWYTevWpXHXqmyW/15oaSF3A
cqg28d3q9Uv7XOIB/in/Gx0L0CYXHwPXob+Gikr5TnuI+PSv9805ho8CeEPM0IMrNwv12F4+zIRM
W9cQP7Tyz4aNOBAd5QpWjkRgzcS6Z4w+9Qbbn2odShs1VF+LYczZRqr0h+/2q1PrI2onO3YlVpb/
iEErb68NIZMMPtciSVgmNwFmPim9rEk41xO/2JC4REaNSzCAyXNQ+aF6aVq7ZklVVm1OTyiXUR1o
faUWG5zahT7r9lLCqgGTxH5fWacQ0nL5wclor5fpYOjgMnMuIz46g80UlsGLEGxsh8AIFQOYtRCq
FTjvfj7ckQoalrKYwLBEwM1TR5vha5Lzq0qEEVCNgZ690R/6TkenxxOOz7Z6TZuRUtfRK87EA6q+
KpxHVLhAoGlWXK2xHl4EfmnLLNN+FZO63w9SoQ5JjSuxksedWQP/uFK1N/QPtCw9WTp7HSQVWTeY
NkBMm5PZahooTSsN7FWsWVpI9vd7t98E0IIQ5VsaI5027neUi1dDcxV0Eqyv/64r7aF01vO9Pymt
Nxq0jbASkRq+EtTEslCr5PVklHEekXV/PshfMoy2vm7w6LqPvjZr0e8NdvDB9fGDA6LqwTTepL/x
dnYSKr/sdOE10aVFlocIPO9MzZFcWJNpu9fC0vPGpfa42wGkOWbhSdmGYS0ke3JvFAaQvEuF73I7
xK0brc6gXB7X7nV6Md2KGO9S7/LKWJUbxl+XnZrEyN5JJuNJqb7H4EuFNhxnElNN5Ly3HLOxrhg8
hvz4w+dhO+kSa8ZcFKxu454qR6gw3GFW4OVM4QfmkohXWOXmhyLJBjjBcujbkKkBMTXUNy/4MCb6
GGm0GhI+ATOFUWy114JeaWo0Fllc/DqqeKTg/7NX4CU4MSmxyERxW91TuLkyz1eRmAtn510ZO5+u
UHHURfrX3YdUyV2imZAhWUP4Vb0fH0JbFx3bSbzLqHlH+v8oKsIyzEyJAhFev4Vgjx9wXpC4FdQm
9JAFPewn+eKOkelKrjHnewUQOUXZvXEjbGXhBpgJptElQ3oaksXa5NfH5BhqkePdRexCyee9vmrN
Xva1URvUZHuqjCXPZe7dJ7A+NP8MRp3lM1/lSveRrBsameDzgnVo9NdW+fi7lNZ9C4+GsmO7G+Nt
+9JEJpXwv+LQKx+rTmLwFD3R10UbndjyahrYn+MD0aN4vB7kVahzSr2+WreYbhj7mISkTWrOsdZ5
mkzQnyQz0C1ljIR/7S5LVQ4oQkq0W3QiX44yGEUYUThXrpwT7B5MfqlEPbjNEJJk6YbnJuYDC7LF
VAAleN7Ad0DpmE3MK1z133/CjBp8nF9e132I83Fe+NW1F8ytD3wkjNlZ47/mpKOg31riIhTW1hnM
oHc/ozhm/jFcX5+jfgkZKj98QIdGp/4z4Ged5BuezGcu2FatFHOldd3WYnQmUBGbbdKOXK4Wr8eI
i/o8j/zU3reQBs+ndefjg6/vlco0zZ+oWMru15X3tOZab9aIFRByrvq78vhR6Id/xQ5ULTBWnDJ/
3fr6f6jkbTn/74krQnyustt1wmOglljBpaXWt1tq+ko6tTX9/9veyLH0f/J/WWmtjHc1eyLP/I8j
CjeScJxLKP2bv21Ycsv3MHxwqqvGzgVjSUZgv5ljlOwTKMSfHyY3kzIS7WuNNT5HklO2x637FpdU
e0lhPMPgZFn5MIypXVIUIev6QlkFvCynaGJOSNq77StqRIYEA5WonUwmhbRGgXd+rvcxc3yhIm8s
up3+ZyEIysafSuDDdE9/nx2WX4Ttw5HDPhkR7oosPvG3vYuaNMN4ShYb0qMhm7JX2RAs32LWjaOv
p3HuqvpMWA6udo0zU+CgxJKeDPv7NChX9xWGG3Ax6jvh6WpIJAQMMvKmMXvKSqDD/c4DTwPdNMkc
QKLN+Ke6qbFERZ3IGLbzxl0D/y4qwE0ys6BvrUJXheFDvYw1YF8BlRVLsrnUwx6lywoygNq5P+Hk
uXL7CktK2uvB4cCfj+u0LtCdZ8zN2apO8hZ8HVB85TIi+YC8THExZ8IMLB8t08YHLZoXZ8jit6hb
IKjwxbqFvdaHVsrI+CtR9OD7KaXxp38NGETdWkPPqkhsxMDU9xzpuswNWkhmBeRBMpNFwytxatCF
3a9bQ0hxsXjdLOUN3AbVpUOcNhDPvheBzBtpE7uXs9beMcBqD1zybjt4A/wbQCtUJbLAmnWzJUyq
poNdp7lFQf0BRX7tI3bg/N713HudL6ca6uUHyWvd07A9K3wfYUbN1x4taI2CS0M+GLASWAx/o4ol
nym0gawGvkQoKgSldtqcH+B6jPPrtBd6vaGTMIMGvMrO9A/ESMJUPvJyky6TzZMhX6uXa7xLOIeF
BFR5PY/mh5kWH6h+DtLPFI0Y+l3T8sLUgv/nkYxy/zwSwXQuFkzwY4+EO+S1mdaDDPelFbbTwM90
M7PtXjTgkCJY74iiZgv5ERd7QWHY6ES3/oxKUHT0x2TnTl89ZPO9ySndM+NOzIWN4ngQFdBaBQR/
BixExbUz04FAYCMcPbnsZPFFXYgmK8Qi++rVICR9W7odJfmp2Ut66A8k93Dpra4zkmiNNF44lEwT
uME9B0rIZn2UuvF+mNd8Kr68c2y0qdscyI9edOS1egjOHdDqEhPDJwceWfT3a3XGBFBBJMm4cKDv
SW9JolOs2l73Za++MAUcNlWpwmZuzU4j++AWPgLvOPQ18kTxrUe6LJzF2AziWhq67b7UdL0y2tSN
nGxuehDWIaRPfLnvppkmqWWx2lVu4mL+TU7tBNYWrO6daL3c16NIpJp89LyRRe1BlnuLCUuGcNoT
HA1Dsw34wnHnmghiPMZCKHVt1ZlxqSCH70sLnYya5EqC3/dfGc5B187eKljZfIGlSaOX70vOWGQt
AriHw/cn1EV0CjrHvlt3ttvS4drvpkkPD5IfXlT3+zxBXj5VtBBWHNG6lfHcB/CDsoG48AvoLwd4
CpHhznRTtT87prjQ6em+7EvTvpvllRLSVHxg/8pB4w9okbO4Vb+Kfgf15GTJgPUADgT80aA1rDWs
qcv7DxaKRQroJ6cjWdFh0nTh1UtS5LOwgudkmka2RbhEHMu0nCvg2zvpezZxL/SZ1jmos5CMOBnF
wVbkm0M5rxyQewcvQDyFPF5LdmfwJ9q8TzKNXBrQOvM2y47daq1SJkyR2eAsnEmV+ZIKPhWKFe9i
XPNa3XioONGl50V1fiQ+mlutmd2sqMmOhyD1gmXGDat0+jDxJUSHhrXpnM1mbyf2W2KHiocYwoUm
NJ3XhkDb3Q65D+8Zxm/BuyXAV9FlIlVx4sFxmD75Cs/56N5gppWQ4prQUX53t9i1fQG3gFbtjymX
G8CA86LIXBOVDthnqr7zJAiK2gWfFfCTxRKvipYnOv4f1MGt1cLAkMHtjfVMCH4AbY/jA9kfRZfJ
Ou9JGxF3/Hu3edm7PO0sspoV2W3tu5H2tHGVS/MKPBNKBwFTlsc9O+da7R6utX8Y7evMHIGLGewz
RdrKpfhtPtiqEeTot8UZ9kVH055E0O5BIJT2osPNl8IbkWu+X3VvDdEx0Qkg0PHCIZQ8nPxXzFeH
977gpfZkknMK6N4Ojvi/k819ags7bQqLbW2oF/HNS99ow1o7ZNLruPX8Pp3vOPB1zLSk+0BikHdq
DdOYGiVx34YUaRUnQUMfvWMoQ7XrMAK5Fdv7bPMJfNT/Hl/aKqBxrr3wUrOyXqM0dDFp88+GFJ+N
kefnpC8gu9O+PfHzWMkfcU6t66Ws/TG5pHbjc7sidYHMhqT2NiZOajey3sV6otpQy0kXx/OZCNss
tQ7REDbTuhJyJr8v1FxmUcdp1YYbnHhCpXdDiywcB81Fc7E2jYMAJPYi2vMGnaz1b/DbmCc35z3f
9G2U+sCScEcSWryJ0FBGJLZFPiQOu8UmRIT5YM1Awe6q9W2Ktl6JIm8QdCgJoy5o0JCN40oTW7mv
UC1+A4w4sJVxs3INMObHx7/pMJU/R9tdjwDbo5Co73/ZK0x85oktl0fr8yhj4UNwR4E5YVBqE9zd
YLXcFPab5w3Spsi+9PCsuVxk1bn8eNYlz7QAGRi/aS5v9ftLccAMtchP/gHyjsOy0XrGGSF9nSIq
Qh2j98aC9yh1JSyTxZJhWcSlyD2qeXPaklJAUFfNwxR0cPgyFq7/2m9f0UDEvPRPEyBojLbla1Hk
C+Chd4PBHOHsK5hrY5RN9ygXn5WxN5sNqV3sJdEgZ+0NacMDvw2Xdq35MzmkLOfFo6LxhYRTmakh
eTYQlX1uClgG1X9PMTKJg6dYaOgMcmumEiZmU2WV5AGWv9yc9m2PHNRYfveLMDdxnazp2TZ4Itjp
HGoAeXyesPv1LtJQxK392j7Cvy047fn1cOgxNXKqStWz+MHTm0YV/5LcrPUZugLLE5zQXxJ3T8fj
kb1BPzOWVRSx0y3QDLF9e7G3c7gKRhUv8QUNA9zzlLugFR2rUThWUW+YYwltbwgFEVHeFoOvRpoy
0Wn6ZfTkuWh+Kqk8xPJxHbioh0zRaiOCquTEzNWSR+Za7BLLIIssjxHrvzUOP8/LSJ9TU+SwT07j
CBHeMD56h/9Le9nB6F1zd2mQywoyhzyv9uh56ZF4OegVZJ7IlYTj8UFYR3udWY/2uPewR8010oB6
A979ZAd1SL4GIc/cjicrrXrvd6bVkgrbeoBlFbBoUS9fbJxU6mJYZHbfQpQPoo4z9AHW7Rp1TDGY
/kvGcDulIBEOMj+/5gjY664MXziTEBN6pf5VklLMxl7KO0OwEsItK8HwqMHGdWaE5/vtIYyCwsAg
YSihoNFuHdjfAmDaI/M8HRge0ZtljByWB6Z+IdS7ST5WLU9+RC2wW+vCfl7FH5YjWE41yNSaJChz
1+JELzKp/F8NirGux/gRSrwf8gKb5J0+unny6DusbKOoqGoq2i1gNiyvADJztoyXOR/u9Onp7Tl1
URwi7gWLiIg7wXC+G46HjcNdVVZ1TKDgpSgy1qItyqTPWtjV/aIW4hQ0ju4a8F9mwZgbu+8qqYZp
eMi4g5ZI4ffaCyfRh01rWvT4MNmxjv1ko+ZPC9iuqpw6Ngq5boEo7k4lkfj2XjaS3Ld+YG+X8+6Y
IWkakq38Ad9RzHbeqlR39IO7owZVWTQK9U3Rx5QlXj51it3joWieCSBmRqOIyqPpsVM1FGz1VQTO
Jy6A5rTFk+mJrtFnzbWhM9FozDiYGgmUV3RhiH87/+tK9nl82zJ6P1WDH35br74bMDlWRT1Q570U
DhTWregEt1VduS+2S/um3TTDuY66zXfc9+4bdepbHiIbAykbqW1Mt5Gj4mITXfI4v656KNPb2zVO
iq1iktSx1AiepE4wJut2KqeqsrzYovDmhFVQy2Y3pZd8ZswUDP4d1ZUUwq1gOuL+UGekb5FFAdTN
ftnXzZHVE+hmIkq1PVRQWgfyRTSvdfBuj8hROEIhthoQHMM5gB816DjQq7yjzsh8JlKvrdAPuxDF
iT/TIzbuEw0uCIgUDSeX9wvYpAXXQkwjSvbgWH7L5yaR751cTnzq9JbJ6mqQEeioFxjoTawvnjJz
cKi7Dgdumiz6uU1/tkFYddZldGs4thXUMw+TNDtgXCjSHBc8yrNgYp4d1MiuL3p49Jf7frFJ7Yk9
VGegfCzFvHvC++nSCIGvbECNEGJ/kP+dtngHFBkKYubv/A7BlyBnhuvtYyAKenSt2MwCGW4k/yDW
qUnYdXNIwnkC+iYCt5YT1OcMNP5gzsJrERhAX9XfDk9GMeu6GXtzMLqKcagi30f6W9nk+azN3WRf
N22NU6FLwsq8uECGY93XptIPqeN2BNYlZO208cXfIpOXynPdsKhVTldbbUOqNPQ15BSSGgkdMHl7
VhBAGXGyRa7Gkdb/kBtcFWr8Ou/cyRfYR5or3UcHf5YLtHtx7bpdw8Lqk8D3jDpHRPkVCgek0N3n
8ydKLFrO/wLOtfFjsvhvJVj0vfpFLL+SJ4qgBligAXG5er9mIVx+VGRcxfltAzniezlKESqS68wD
+N6qEl2+8icb2ETCteVOW6p3TW6vhiX5rlxJyeCNUwKlu0NJr2q4MovO0HByXC+JkyZveygb2cZM
Y02iR5Py+YqZCFICXpkBuZmyi8uMEhwZ153x9+dQgT988AOhBwlySLAE66ad2incgKbYx7lMPiI8
gfieiRkROT+faPxkRPNWxlwigcawQl88LSgA3XXqj5VGLuXkg2EYuKlWrfKZ2N9Jmi+Tn0neMeWq
+YtO5XToaj685GvU3yOMiQ6K7T/HARcC33vdHejdxcA9K9pIxceaKX9+EGPmo8oolpKX189MkMNq
PffJBvZuIu0xSj+mtuoSknlSTo/2EFvzseWfNmV6X0s7u/uRoXFSz0kCbCWWnwJ+emYf+B4XqByj
5bjYAkXykD/P6vl3KofUA3Nl9Zz1zqURFgvPbymrpbAcIxGh26QS2Z0xKZxgHY38iGUE0QaEskID
vRfg/bWvsRwdzzienwk+dcZa0AUXM9RHKcV3Da6A9dlKH9Dm2Abwmk8ZvdS7hsd5F6D/pWMd2Fw0
LzpVY8yj6L3LUUiaQvw7hEO78SwH9d9SlyshlYn/FCmF4V8xZfBkKPN3uVBCCmn7bVLYUz4oykAt
/G+hzv/At/R5t89l/MxdVzwvRiaj5v9lr34jLvUJz9tp5TIC6G71vVbUMPMGPaaFiEwAHqkUQRmS
ui6h1EjTx+Y5wgr+LbwBgWtin8Lqp3IPSJzF+DmVWNGnOJ6qpZCvuwwQLcGDVCXxJ+auwtSd/Xwj
S+GlQwZttIh+zBsUu4g/w8Xk1uNJbBNunoiuyZkpOon0rNe7zXE2nOMT9pfQzmGHiIILJ69zkIYg
cXPMCTtg1r9F9yKLIYNBncNGh0je+ZJQREobf9OUpolZunHgm/7Kn9SqR3+bV0zNkoXdwknXIyOb
br5paYTjL1ruxkK6yOIMzqgztxaiJMGInW5abf857765llP+kLHxZ2o3yEXzlVaweWomS9Z8CKM2
jra/Mzt+JhV6iXDV5nrBR9tg7r0zYBr9bRihNiqVWMA3113oTJdVQs2EGw0VVfNEdV0znvB9aWnV
XKhXI6HTwDARkUiuCM2cPKPDp8VSi5Qld44kdwwoqY9SWcpPu2NR6uSTh52KuztYQ54yVZzYCBUg
1CA5ZlP/S7otqK1kro8yOb31V84JWjjNyJ5LjEY3dsWjW8XKaKeKbWj/HHT/XcTyQs0vN13NUIFO
py//dqwTYTYF1iLp2SZNzfrhAFjrBc68M+p6e0+zNLRQnEI/mPFJKkCGO7F0A90I2bTN+6cGEaak
ie/Za1iC7GS6V6wdbTuUxDuU4jgCUaH3KMexu0LbHLZLttnho32dCpUMNcJ8lhGBy9nLqCyh4/ft
QL+rbfxAdL63OZu/s2PUyiwhE5avIfB+n02CECFIG/f4//F8IVD5qSC8MqoXmfq0xmYhTASdCUFl
ImDymuFg7/CIjkRsrRu7a21RnD41pALs7pHBvibAN8c1DosurondPN6A4V635iRYbCCa49fu8FDR
PnLMCwXLWlLzDXiahx2+TlrlHJ6+oSUmyTi6slenwtqshS4UCeR91davlYO2rZFxmMsI8LQ2jxX2
2t7oMoxOgoaWnrthgIRk1ICwfnO6M4y2IW1zKz2kb83YiBwKOaq+uUVQm30pxMv66ZQvuPKovvza
yZpyGfo/sXFXx7WchhXLWSooV0vhruy9fUzEXfIqJTkFZbbag2qC8Jk80glxb5hacDTVn6AnCvti
+iGlf9qfM8RLmBoHTQRqhVhu7uKk36uggPIxTrRVY3lyorm7fReAOZ44k/D/O372wS9EMt49aUso
TpzWbEvBLduOV/C7OwGdBPA5lB3S2Y/e8bn0T8ys1Wzw1EupSM4T8n3iwaKii/KgRmXMG5uvzaSU
pnKkxdtO5iKHC4rejuZrtXjIGwDvSNODR5wfwEtQxSmqXE0bbzZgvryxZyy1F00T8LuOOsBKOqH/
tbo6szBL0/pBUEiptb1MP730ZP4/m9LVs3/XqFoGXTZfx176on5HasOoj43byBPUwuUWYWDPpF9S
VGmwZxnbOCx+N1LnPGzbBlKO/plKhLkOsWrpovz2EM1IEy9/GipOo/bWqOYGhWLfEMTh6LDzUR8d
30WClMlKdaDHiXRjgX+3ayo08+lg92lbIUPbU2RkaZdutbmslrgDp5Vtr3wiArIwuNU1foUjEk8C
iuGfzUj27gGYFPJdafrrIzhjjJM8yar44OJ4y8QnG32xd40CGlnJ23+qPYenp4NvN0oeiwIQYe2n
l0uQuNZ8ve12CWepfsOd6wcMU6ceui9k/fMZnd6zJ7zhoHHWEDaF22HdJPqR5sSKg0mnzyuvr+Vq
HhHPfHslvwVYGBRC8tXG4z1TSLBV4s+z8o7/YwZ50P8hKtd6xwj00lDdNziV/TzczgXvoAb3pBjq
s0FSYSRnPt9lWIU0GhIllRdJsLzmb8gmIfU+IIT0I7CH1zttKYR+dkk8Dd1WbXFDnMYtx2g9Qfsh
IYaNjJKk+g4vAWTAXTYOnUTfuYT3y+RWU/KA0NkDdnbGSeN9MBUHOQBSKcmymxcetCdRvBeE0zpw
5DuU84YjJTK5DPOvMA5NSB40C7619+TgrotGd6IZ1pFgI6BWL/hoYtiZY1s3Izbtm2jDYRgLQrqz
LLQvyPT63GcLW4rol3nGMsnsSNtNa1tOiCV+6+e7O0i8cNiIjldwq7ljh8/ALxbvMVpach8RhnCu
m6NTwnSC+HQYkvBw7oGxCzzy2MwILb+lSWr5gthv3tnOiUAm+uSGVnulrceO6OkvN14J/EenC5zH
fYCzldBR/EgN8nhFs0Eojb/xlUJK2+UDvDvOzsShYa26u3mcOlwYAARGPZu0RXdfZoUTpSW8eK7o
EKnMH7vOAnYlR+aotpcnxNc3ubX9FrRzvqKnrpJcMvpAzoTcxRSpdzmTN/gu9R7d2ipmnsjNvJYw
Cl7fEiJrfizI8pfxSrJdfELZe56d6Th53PhqbQ/hCkw/Sv+qpeW1WiDws/7hlOwsxeGH1KMwj9Bo
JY81J2deoh4Ar23X4jk/LhiSB01swTBKXrZ7/EJ9wjT8sE8ceuNMY3q3rGaMrfoKLl4YYqv8Yku8
xd4ro01rWkEwBwbre4hiWp5X68ZZwLXU1lP6TRW7kFCjkALpgHc7uZfIuBZODfYFYuT8mIWiZaS4
72BKWPMvhd7hW1FKzicVwko3ExmAZoqJIvgorO/GKgrXCQ6pAxttzhoXrwthIfzLvYSV6FGj1KHs
owybxm+GKNCxCJxRXLhhDHBal6XtWXIytnQVIPWEFLWaLhMu6oI0lKdFCnI51OS/RDWPZCt0/EYW
fT/ggSPPi8gDmUGQnPBF0j5+Z844ldNp0pzfIoAtiZAFilSEvRa2KPu3a5WB2ION+LnRgFVNluGG
4psi5/26BrJOa8Odcw+xPb+kZltgLJN8TutPBmwVQ/OLl9/bJQorgMZSFwxajdRDzsyOKH1xfHhY
+YaUOAw9en18KnbAAIsTsCxPSmA1tOW0NmBzeklksUqzGRywO+T4QvQzdcw9nCgBGsxLh00s/Ckx
6fUu9vM7RNtiFDCwGbGwy0hmZ9wKDG2zze06UNzkn56FBiYaL3h4tCha5PrVizBLpLLU2dQoCo5J
67wzyv8t5iIOSUTTd4IdYERVfl7PUTfU1QJgbT4Lw+D4ZOXQVKrt7XfDjhSLA+7KyF0UUD1dW6BE
jtA2JWYB05YNVI1w6p0Z9iQOFYCIGP1o4MJXEjxMg/HTZQbuhCT06xYx+0mZiLo79d9KIBQYkNiv
r96THBj/C6LmdpjDzBN3Hb+dvoghmDkotNshH4A1sBlHsYsMKqEPfFF5ULjw6Zks8BJ9YW9qYhlp
Fx6qPNiv3YzhgTRBEjqe69Rj2JelJh8/K60KpKVtGqCrc5Xx1SDGauLP+A1bV1lmNUzKCR7NE9Hf
16qde+cu5rVeSKLHfGbn4B2GXMuvTmN4y/Q8xrEzyiLdjCcXYnuEyRa9EZ19d/isMefJjiHDayqE
NTeru2pykVE75KpjtSRqW3l61Sy+XJuq42oMz/+vgyJcSNWt2AzLj972Is0CXoJUjIF5pTs999Ne
Uy1lCChV1N5scSSEug9muXqxaFtPBGCV3tMKIq/NcxjAPxuWLgkvFzWtRpaHM8zi+J1Ea/ONzyvx
FGZewglDEhoOpNoE3h5gkQNMU3XaKS8QdaeKkCQu9Rx+O/JOehda5oOtDax4YMIybNk0ovqG9qWl
/6AiR+WI1eDnr+Q5C2ncjRWi/4cqOAGotzVwuI1wNA56fmTw4i15MrH9jNf4aBEBkWaIYcUtHQ5n
cJLSeiTiGNFr63I46BFF8d7Nt9wlWvBafoHSSr4Q1xNJAjjdjxWf7NJADPeMJqDLSmHBwtzQUjft
iHZ8IPpIYX/qO1uW6Z2s6HR9YviwzAQ95+oIaWJsaHAYvyGnwhwkR05MfKT0EreXxWfd04BtV0B6
rbcMUTwiqR8G+WBe7gC2Wl1KbJkgHB1CftJibQc4pcgrirfdKknZ3cyNHUZmcNcm6y+SO7FvlelF
u9M3V+LTxwSI3HkA5W2co7U0yQDeO24wzbWwgUmNppexkPuFqzZi60zloIdvYs+BYOJIhX90xIo3
PfCKHfrn+L0E8657RQ9n0MmiCOEqe6UKWgxZKExcv7KMqFeFCOWI6KgznZxJ/l2DcpwTekGV/LXO
adtq9ooiUIMQZXdOPJjWsCKp7pwYVzvFI5bKKy2i4dBWEtbMfnNXy3B0kI2DK/SmedLC3s/tf+1p
rrlbpGztWVQ6Rpvx/M9gZ0E/UyXgGmFr9H1ktrXHkaZ3Tqu0IHbWSGuDyN1AdYaHa1cTvNEkRAP3
eJ0KWh0MIn1VpZOyjXT/qQIFETeeRc84VELenFGPi0pLlPcGfOxhyP1ZMqIcESf9rvMiZXuMtshG
LMk7CtP1WFQny3A2e3H+4PJCsUJpun9hpj/T5xPCYI/6wHw5x4LbmuDZpPeDYlfGoIMxdQs/mxal
+w6cQudqSH+G5tijB+sdjxJbJdRZQw3ZnrWvXYWvzPO1NgRmW/3oz0nd6EhQnA+sLCOVK+RGg3Kb
NhqY5zgODJzxLNw10xXPNY0TnbW1683sJq8hY4So7cXFF1P0BqdXYZ89BCv3WtDFwwB8FfcsOGsA
yKFQQxaXaTpy/nnJP2cR7rSOlm0BlUK/E+T/jPq1weVcw9PwHIZPZuqMuthPzbuuqFAGuhA0Tthz
/NLkMYvZ6sDGYF85pwygAxdsdVUZDOWWgcfeRi40uuouyyN8zt3D3XtPXELyy1VZMoXrLJwl9gEA
/WOcD8ucFPIFByj7gTDB1HhLCZ09k9KOHUFISy7Swd6W9a0NYDkpMzn3Q8WlvbEADrFocg1UOqjs
uHoQ06k1ousPQTZZuDpqojyZwYXsPjdlGlMVnjNPr9cgABq3WHjlQF5vJfygEir7gPBJZefTYDtf
peAomgeijKV9xptdtv6W4C5SXUzxYvY5N5hmiN1X887Tk3WK0ImR5IWx3a6hqBKanT4/C8kCoQbO
s1SEQii8U4+xoNRp+yb4ZAmgkgLej5WipUSCxAtviPlM2YB+62Dwlwi+7CIzs5Z4IT270ywthvQ8
0VYPq5IP3P0BGZc8vxHcP2GzqSEAxt+ZW2jul5HxgiCyvZYEcysqSHzU2wRbu916pVINflTZZ+bC
odU5RxjxjJMy82rAhnN4CmTv09CtO1wT7PjUfi96lcEj2ZipMJpsW7pK6ZHooEKpK4Uvts4XHcrP
MTfimVkvi2O74sTFJzuI2hV/KtOfXxDg5L77q7EzkSeLRUi0R915QeIVZNJbK4GoE6OfsAJ5l88v
unwIZEnRDF4f3GXkCfPlAtc0MrT2Igg5+uvfSBTonttFsB4oCo4KIDhAqY6stT7rroBiJfLAvzqg
ZPHhb+HCI6+vAeUjaGemDcSmtfxGMCEWyG7EL/LihQxc/+yXTyO1jAqK0VPZVv3d70+Y6Fk/MknB
l7FnEZ2j6gAOVrekD1TE8uJ62Nzs0UA7FIUy0W8Ptr8BqjEODJ5QzNBPgLpJYP33LoJhKs15pJgv
jYuwmTdGPaN2nHmqh3SBT+xUzPAPV0xEmnFab99OX1qbNCoJjhAbIsLsIAdpzKGW7UW1T6weeuSt
pmAjn6cRadGtAJZDPYXUgr+nvcQuYybCA4DRx/HP73FzHBNhYc2Cly1nkOeIdaFE2SZvPAaZpdkA
oo5FlkSD4pmMt7l1ISYoHYLdKqYfK9ZmkIPkVPcoHnl0HaDYormpD86YJpSEZrtVYS88bRKz8ZUj
rLnZATxF5j0voTpDP+Gwd51kwVmjSJsJdc85/VLbqAfkSIEtzyF6o1LLk2ETZYVlVIgHtld/PYqA
4iqDmrY9UbIia1DeWeuddjV4OLgTGghUbbzxVAg5TWD3fU0achSdxYvlmy3daBdUeRWC6NdE5AR4
kN9JT2YkGexGfqTbz9z9/tTeqVVQ38H9rmqfFY27Z+38GdmyL5dcKKyS44meeobZKY24Y61mcxBp
t/2WrEzFRw7LHRjZvtaOeKRRe1J0SjpUVmaXsi9Tt3z4JxBicr7ppH8GQAWVokeb5aIDYRznUbDT
R7lO0FZfjMvy3HUwdK5aVPNZHL/GaT/12QM9AwKoUS31YmOHvzJSEKGGaVRgBSHqT2r6I4FJrrwf
p76EBVEv4T4uZz6qhhLkt7hZQ+6RmA0l5LcMB/K2vm7Yc/E/MPYheOwgjQ5YXpeG+jHDA9ovuBl5
WgnPdYNWzZ9kAeDBXIt696VpdyuJwPLeLlS4ODiIprNFwNMGaASZ8pLx1u8YN+1+eVuEPa3wyG4A
CLTxpMQe9YhBvULriEeyjtfAmWBAx7rzLYGJ35aGR+uBzEJN9rpYtilp2dpy+4PGZQYpW/LzDimw
yYQQbP9z/EJG5n0L4jQgtkuMORBjNzlubUE2uQhwNRSrykhia6lQNRljLclBP3POvBfctRkEkr22
DwisQniOYwwJftdx5et6B59TQXBDVddNI0vy4ppa4j/TiUnnoUmMfPEZWUFdWpnf2/n9uNLSzr55
qQtkzYvSmX3muCTFm+L7z5e3oRfImDS92OLyy3VagKHcv0Dq5ChQKtT4iX5lbXCkmWXp/HVIo0fz
8fGflk4g8f8oCyCAbv+ZgyO1JtTxSXEFJQRI2cpSVYrdin/NdzdZ4b8HhuVZhDIYi0a2OEv5H0Jb
vv+W/zquxyKdOwqXHl6QWuEAc6dcRaTq+E8SO6RaBpj4cmUgXB2KrCMW9XjGeQWgcYS/bK0dq7Lp
6kYPvaE5aPSyxUD6XA60cx6N2o01EyHLfEyxL9hiqwzzD7/SO0zsE/eM6Ry/0gH7nmpDKenZxQBb
7rXlRLWjNNRPSM7gQZqFR3sVder9dVBr4YNUfmf8Bpc9ooxzN7VuTE6UuH1vf2S/o9b2sMuDqEZo
9gub+QhLFaNvDu/R+F23jRs5APouKSdmZjxm0EDpb12WOWdaWaacKbiQjZ45RKgw4369Be4cE9dU
B9tlucOdIN+alSg5f39b4ovWn98wWxBX4oc2XXAhZVyAqTZcpkz3VLLqOLeGFNKCzY27mbQ3SPyK
f76817lBVycw2GWjtwc0fv/GLPnZmAR6jFFyUg7VHHDBQUyqlotZoTQyyoml/nP4FF2PIVrxU8/A
N0GcU9sS1HNWZ/u0st7NhoB6sLQC3dLxQlrgi+56b29ufMntz4EOoTVna4GMlAsFfnqC0GlZFRtu
QY0BGorq449jpYthcla4+tR7K9Ab21u55rNxXGvB1ZTu553IBA7vZ7YK+bP5zBYGkShwuGiRw1lZ
8lyQz9HGL00ut1g/UAB7Ve63Dq42dUO7Z6izNFx/88iWdj8f/54NC1VjWStWDEz8wHvfT4zEmLQb
cKIEXiPcqRii9/Li2oRYt5yrMLtLj2y/EwNdOLVQhXuZb0agU9H3R58ZFr17ZypE32tqyS6qpFFP
K4/pWUK7+E4V3O/uflc5C5S0x1t0tXzkRuWkrbeoZxEZzoNMuGJcAsIKVIMLx+p26N+5wqD9E0h6
8EO9S3w8Exwy9qXFWi/sbAbcPdeLRQYR17QsVjFEQ0jBD7DCT6QTFvZZBVzuqi9BOilDQn7O0Jc4
UEb6CXJAS9asc0ys3DIB71BflN3bMzpdyCCEZl0K+2ljbbCiEn/qZE/R1BA+NZLtH+9jltaAIODq
8/N0chL2YSijEVbO78XrhSEUsZDtkYAVByptzDnc1eT9smTuClIFCfOjTEG0Yj5Ug39AmBvA5scm
JAOkdsnzRK+gdZiGuE8t907yRTCmsC9nOwtsU5wvB34I8oYmjTvMT0cRZidqP2UJBVPSjDziOgbp
J7U4OVdZZgeaaEBCf9CxVLFHqwed1XK8LyrbCFJK16aO04s7+vAroCTfJXREB3fU4FCGNRLE/uts
f2NX7EOwN00prhpMA25zBXBpTIBoWHzwRXqe+wXhYDXDCRenVo0RbRt+0MsvJPRhfnvvx4JdAAJl
+pf7W7Jf2CgecqSiQO88X5eQoG+wOQF1d/vx8Zuy9ebEFOjz04T5RDGT6eMf2dqIgzNT9hZQzC+J
0ehEKgkpnMKj+i9Rp52MGtPIqNtEpKd3Q7KuAZYqOtHtywmcQ08p8XEfowKYwA+sZR9B/HjKpGdV
ql7+nX1AFaKX9mXP+WZezHaxiZhTPtCABmwLnPdjdejUczRV8vhSHwaEzErb47621Sx7Uljb+Fjh
hb5ZyNzfsYLVlI8QFfeEJ+SulUTzMBRHobSBx/+Si9J6jlXW9RsxvgzHma7i2fYFBMb9fFwKMIkk
WOJBjxo+0habavpdbcZo5kymO0nG2GhC+Zl4gQwxoDoBrKIegCX/cNGPRRCsJqo0WzBzY9tVZrPC
xAVSbV6lwBDMs9ibzPLw9Mgz/YtUS+DFQbYvs+0wTX7ZmERo7Lx+Vs7yen1Twp1nGJGm4bEt9UsV
Tz/9K/GotAflhy0ph8Je/g1LftTV09AYp/n0jflkNIm1qEb++MeV9NwNft/Z++m3LD+Atr7SsxbP
vc5gG39DM3rqNrtaXjJ7Do7gXLQaqQ76WocN9qLhkyUSYkaZjYdhrNqNFxFntsIk3PvKZoB9OaYV
pgvwkIoORaLh+TLFa6HeiN6sQfC4Dgphyopa+Eqf7xeED40UOuNdKbe8TWZ3ra5qbJLAEsnYJlvY
+5/iOP0pg5c3sINwA82D95fQf2sCFN03OkB2n/absdQqfxXvBRC7PF6tyTVUYdKgQh2yVQLQF9DS
lHLEMpcKQ1AVRpBRIvnZuJvHHR5kYCn7o/ACaHIbhLj3iCO3cmuSZgN7pw4hdupmQQR6RJVIyzGu
+TAXCmiA5C1y8dzhvjn1DznP7O/ISo57xfg0moFOunkvwnvn6dz4MChM4ZdNgdB4G7DskZYgLpEs
liJdIlNW4eUPqLMJyu+B3ZQ6gmg+HKJBxDvlZ6n48DBAakdJvJp2U23D9N4GozyhtYMagzhmI1qe
njdsmvdz5CuzqOLnGhUo49XeNJsOAFlcmmxkZtuSgbXTF6LA610FnjcxSnjaPIZZDoeEZ+sxxYS8
zn/Ucwh5WggFNLPV4rVXGGf0vnEhBGQD77J41nz2x0arA+Ci2AQC6xPRJ7xjrY2CpHZOacDIeBX7
KivflNHoqSKQ8kEknF3WdhI1gdcE9eZoYR5A7pZW6iR5MUx8bjVfAloGH4xdFU/GpyKxQC+rGy0s
2Q4CYd+q715eUxEgDwuzfSnsQG772jB0ELbpAd1Ocs2NLtAGzSfJNtjTakeP0EEOmbwtRlXK7pDi
YOZlnaHmNMJqab0YrdyHK2cJj7KaR9+JAFkN7u6Z/hit5V8OrzOxuQXryavnA5e4jCMCoAFLgBzn
9HYkmoTE1g2H07uDAk/DXDiLDPdU83nQzVLsgMy2rimNlxKSuH4ZWr4xyeiUl4TD9/LeXfg7Rb/1
mxzHniesxjy+DXGO76aWVmJMHDCSUxUjcSbtwUC7OYTVLLnPxm/scc088kPuCpoq8UnlXKu4yQ5M
q7IcsyxtufxpQdUOUzXh3JKT2VlZLErL4ZdJ6Om+sqOdrKim5rS4B3axFyJdOvufWVkk570JxcwG
OW2xy52joF0XWkW6lPLk4i4Jp+C/7oOK86dZbpTS9Cj4Sa70GXEm4UamJZgOCPBoNLKjc2b0qsCh
X//CTJtoNN/8RkHuK0IPUMEF/QSmYS9mAMn4ycx+ZBlO6Z2PZTl3M6+xoA/pa3/XXwCdq+yCS+mc
KY9xnLUnJYmMUA3R+UkFCIqEozLijK5dpPx4zAo9v8L0kBpswfq7pxclCp4LEhETI49w0yfHFtQF
8sYcE/T54aEIus2eMOtd+fny72aJ0Sw4VjOyAegX9L0N3wMoUQueyubXmSVF+NQ1mxTkYjnBL/qo
ixRXeEBlOUIZA3o/N9Ve79LD6wX3k8xbmQOQBs5Qi3D6EWqT25pmT6wfL7kJ71rvQE1se6pRtQZe
YPXIXISUQCWcyHxwgf5hpg1FpSsYEuzFgnqm0Q0QmNmXuCLDbNQKYvRt5JEex4d2NdVW/mloA+pz
kJjRID08LXScjGx49yOHaGvhqXWK3H3MKVt8+JEOo8T5dgXsGa1klFp+RA57c/8qvA5bCT/7vZdN
NhTjonB1cDdbzb+jkiPEI6XcuL+BwYBxuy8Ur10ddfsJAojc48QzrOiBnDppXknIsupwuGuvnkS+
rIJMhzhe1k8aNKf7JWjviUzjhGcFlPPHCj0xv6OzwIAI7AVuQZ4rI+ND3qwVUZeqfkhNjKDsU8t+
b8YS/B/hQM2q5YdMU/CgTH6QwFPEmIGoqMjbQktkY8ny9GKVr0TmUQrDxnCC4hcwYhfM10jAlI+7
9l0A/sQh8BoU0k67rjzH+nFuNwuMpNoZOIQzNxSQYRMs/hEE3NqZGoSfVqTc2LutNVVQfi/SOFa/
4JStegTKCHsNxKbrcOI8RbpnR3ViFj36MvqdGP9GTCA5MU7aSgqC9X3gfGy5wm7oFVIdfygcZrVc
DwifXV79Yob/npmbvxqTKc4zEnCLKUYmFNviulBcQRKT+WMrU50MzlkoIow/tpj7wA+HN3czOzto
BE9txtyi4DLdvA0911QOPKWYXreX328aqEtol3EwVxwmNbeZEltJDqHn+ov4u8Njw+rimXEKZEqP
P8PNiBwH7Mn7qWthbnE9TZeuPTqIK58anFk5HkXSNeL7Hay7qIFBgGLpVGNzVlxBJP1uNsrN54xJ
bdz7+7Br3Jt1bzqxae9oiYLa29XzXsrRekRT51dtawGhxvGiVuM2STL2xOCHDsY9m0LEVay1RwMg
xL9XmK3rklD8qzFG9N7JBu1htyqvrb8n6t/MN5TNEHhfgYqf8/oay3fZDXckFz5josVXJcX1pmbO
pFs3CJWb4yllv4S5eErCRtf/XIHgzi8n/Pu+kpcsD4F3BuWrH06H5/AiSVjGHKHDgbOeyKwWHPN4
Lu5+dt8qZuUTGzn2BqWEt7DMgzH+DJPqSx0k1FCtsMtklUMNcfhHDw0ozIJyUwJ1/DJsFNpx0vGj
9TpTNty0OCwhTP4o6A2gDFEXQWk0iLBNgz39j1gFoyEklBuKgU3vC1xgBiL9MV9QjxWQvxAM/9fF
hZjVei7WRWWQQaOoMVGXz29bMl/M0haX5PhANbmOd2HkXQV6FDW2oOAYrorqbDzLbJZNjrMBb6wc
A6fltbv1XxveJTV1XyG4AhHZqn66PDusQP6nA2HkxWr/Q+nkU6Mnzy/wIhvufQ+auF0demp4WFRj
aL1XN1waIrNRlD76sKGNYp3S4LAKif5l/z0lfTw0kK+Se6nLizhsuYiL8BKYxiGHl8a0FFJIaoay
dA/8g3J3SFHBIo5w8tVUbmWSiO/4Zz1at8SIhQSFA6jI5ug9BDREeOjLRTjDSSWiPLFdP5RzJS1U
4sEOTbWNZQNMiuO1JuvAdEwPLG8l6VXTpFVGERDceHRmO170xTeS+aJsqmmuNl7sIYDVCxbnZpfI
2mZbSczvUVHyFgwNhZTFdcHZ5c76kpMkU5cdCZFrTZLqjp2lrY6slWo6buwD95LnIvsSqVY3d7FD
0m7lHZ/Vobj1S+S1mUPZR1stPcWQFa9D63tDZvIKu3VUmF9dleoxBvqaKlaif6ThKv6ZwDA0K2DY
EAE5jh6vpYQNWiXK1iu2Bsm9ZjwBer5hfgwVljJS+dwjmuGPl7hi0KUrM8DsRtoda+b3t20AGJ2Q
mGFoo/EXQhPhif9b/NllmIw7QPDDHDztBt+U0K1MmcXDEp7DBKSV/hFvGItOVPcNO8vMhlSBDWc8
nWPr0CexMmWj+JSwqIMJ9wVXkMjO4tWBhiGasSpNV/Be4M/k/fLaZeRawvxOg7c5ovziPS7SKTuJ
x9yV4sGXdRPmj3HMdHx4w5n0hFt3lRLoxcj3gwMoEXWOjAORVXDvotO0ZAQ1vSMt+lXqSjZFVDkB
n2dulqGSEvMstwjCLSZiiGX+PIgtp6TIuOWVwCPwJA/dotEAurxbMswt34B6fYXpGMG5R1r60LkV
uJLvmaehVUEqDcxk4yJMmnaA3vTJEAb1VlzjMn+v6dqWC1kAmnQfk8rDu13aRnlGro/paKvHYOpb
Ecnc/o2MnO4KpFcOQMC3hX+XH4eHD4a49YVmxp8gaZ3DuTaRPKZIbsCt6ZUA5KD8fj/3rZddqzgQ
0jSWIqwfzH8LWGlKY8fLrKXX8Hung9kYbyGsA5vCGAR+ZaLLx/QPdXSwrs7Fw05S2rn1R/gKsFyT
f4uJluvH784RFWq7RMDxVE7P09nPamPNnRMZYP5NhtbsiHlUpCOS4iTy4FUJR+O9jhouaOlzL9hT
63yp2DDNTW10YfD3f84pWW33li1DKdKWpOhpYhxhmc2hUz62oE0h0feliAMZ0vOziIzngL+TMP/B
PQylQDItMmIXZM2hN5izClwaf3jPGKSQUFvHvhTQhtrj6NmTm5AsgZtrqCPu5opnK5nGRYk/HU8J
yi5bENLsJ3zGGc/gf+nTuuTVJAxJA4AcLvbyPcuqfCjujxJSYDXqGMQKRexeZuH0ZPU8p5hfkQ4F
xXtV6O6ALgw3eMgt/0dzAgLzubOPbS3Rse0WYxkI9wxWTyQvn8rbqvmTGN7SM4Mg5YpNDuDWL5Nb
yQLkNA5cbl0CNhSgKCiy1XwCxldxtlwB1dQ3Cpqn/uSa8YrMzzott3JQGpqjIvw/MtbY0MaEI8te
KAtQS9GoWrgyCO5V7aU6vNpMqF8wKDWDT5adGFG+66DL7ghFZmAQ0b2DWaXfV660SG3apNSHx9MS
IU7Ak2s7WFCuW2PKhKYf0NhXgL/ZppoJGBnXEUI8RXDeYg43v6HgJ8VZjo77ndZlpu0Bzp5snd0h
1cmfz7wLO/8SgC2fYw/Mf9suenYLje4ur1LGhcEl8nc8x8TJZmWqxHSFtAeZkzjUUFoGM2S2tgDv
C+9qKMu54xAqSo/Q6qs7bTFwKRsB4pFnr+cG3r+X73f/jjRmeXmylT5aCwPlsim1GaE4EQl7Vvim
xTNdeBaltoYuQfsIJucFwOOJOpbptGyE8Ek+PxXa/WEYCjdEabLxjjDx/oCHybh/BTYPLyi2DMnm
aV+wB9Pgxrr8iNogZ1LEU95YntNO3qAQQKnJi7TqEu5gQOADsiUi0DubZkyM5TBy9Oh8tRnTB+g/
6xx4JYB8sHEeiO1s9Wx0ysVJsWz1+nIPzBl8hxmJvV9klR0unCO4mHLMj1aa2eD9rvGcyqvI5kJh
EINS54nCK3mXJI7ENSf5qa7xORgkGZt1Q2/4Ze3eTBTfDP3wTUS4HB2KTdJ0ZdRF10Mj44N0J8ak
ZdMNWM7pbr4Rb+mFY0FP6ygd7BzolubaGe4X2vA2TjxnkIxKz6KVVT1ZiVdEORMRkmnSD1pt02nC
OQfZNM7gooEBMt7YMxrzoMqYif3DXyRFty+Uh2RVP7QDAw28yxtyWcumcy9yMga28SrcYnBf2Xv8
k2rIj08uNW2kmOMKbAld0RTGZADebLkqzNGKEQR5bOD7pLXQ+4jKKkKRTE555WJzW8qkbyj+nk4o
/1Tfhxn2K6VXaILSMxjMIbx6mipwVqAxrv+CHH4ct9yWSIlW8yzyGgd2YsWXP4PzHYkyrA1tZraF
Qp5UiizZZZf3V182Qs14AC0Zz0Kfh5zb6L7nDdeqolVGZskNapGzRP7jf5BXPtDeSV1QNV2TnE3t
oTIQ3gpahMqOuFduoPJDzz1HyfaU4lqYKrGC8qwOoKQ4w5WWcMO7D4TnaNKM0DmfTh9z14sMsBPm
e82BJniQZfTZTvh2JqNjQlshvYvtUdNsTJggF+9IS7e5Fs6fVkfVx/TYYo3C8JuRkQteeyJxcuj8
hwLq+kUJRw/7U38CbGW14oAdFhWa7BcTGnbp8w7ezoZFFwb/G1i8x+iIzcVe6aZmwIAHIuvfW59E
itJ6t/YmX3emnzbr9oDIeRfK++5slGAAi/YrQ4j6sp7Lpe38h4bb7DnbTVbkBD9U2QQJqSSldKk7
DvqCi5oSM6dLG4CBKJiATpyE+Q6qIsjYKVnCCB+0R9pIdW6DooDGIAwQXrVl2N1JOaVHl04AT3Kz
5yJURZUlk7T92CRdOUVRkux17uMA2NckhVBpJWcq9Pp/bWxuoHT1tojHQsrPHzQ38smGDDoGVqwX
/QgPiCqjxWcckyVIJFqGyEqi+EjBBEzdZ1ZQFIJ1JMw3r0+8+knVMB5tJO8TvWQ7LrQHhvrAxtTU
PDqkrcz74lFOifeNohYUhz5o3+Q96VtkI8QFad2cP8hAwD+annxaDKAUR77uUSg142LI7WrRK0ib
ta+Fwmh6alnV/3xB/5B+RvvHewCOkLsZg8DginD7R10VfBbRQAwtjnDbDBSROj5wIIx/ONMA8AXh
zYT9dpEu5cp8X9VChuuWBNqXEv1NU5P82JSFqCtX9C510aZ3s35nDbPj8Rn6pZNT5/nG1IVx+Rvp
UmSUyljmSE6dOAbWVPgqqatmknmZlnHtDs4Rw6Ktfy/gbWWzzRaB7RqdaNHGpmkkK9ga6DqBAQVO
sjkQj0eHFmtic2f+MwlcfXNklZJErM7Rej5s1vRcAszqmVraGsuBHHJRDaTc+/l4bOP3FO+tPeJ2
ki5Tz1xKyCmem6f94jrHWya/XJXdGXY0cVtk18bf/a5jRJbSUWfFnJ1PCzIJ//ixIIfWmQzlUGYl
hUT1Fc5zEk0RCnsRpv2HgyCjXGppFQxWEEEIAZd0QsMm2TrlK1TbSghyyXbduXRqJLQGiQYfI4gS
PEvPx45YYw+RWl/woPzZZwqn6XlTcEmI5I9aBreHzfAVGXkF93pPrsAYM1Dcm6R/c7VvYg9fRgLC
YhjmpluD28zJLOQKhm4VZwGfE9A1b5uZqC36PORHP8FoV1JKlrz3lF8Qy4gVjshTWy8DVWi1+rTs
9vD/n83qot71Py4Yb8AlgYespF/XMn1IFQ3EAezXynmSVsXfamVsT5GB50R4EGZVioRhZyWmC4Xg
rvJ7zVvU3fobCXt4X1DPyiDHykq2+RxEx4sbftC4AYeiklnhulLAix5G7AzRlpkR371Enx+cp9dz
168U9trRHlPyEOfyfmxMHLqbtLQzQh3UT/0MbGtFTlrcaQ/aINKZt359i1W36weLo32F3CHjpMVe
qP0ej+fv3VSn89ebYGBPe4pEYwvX+sY9ubZOlDJr1fyOOy8AGJ7TW4x1zAuO/V1wnKHJ8DuHjMUe
AEWYIhagH4xyPuV7eQhh+2TwkIisjQXn59/il2G4wq+jYA0AM5nu1Me48KT+XKkDzRQ5BKSPpg+a
w31Lk4iZZKkxCPHURlnpUtfu8cddyBohbVf2zMITnzIiw53oFXvlWM4n9qpRJjnK4dCmnaU9Hlfr
1M6m10GE9XqvUjtvAF5l+lVd2/FqCme608wh/gmCMNeVu7cu0AvTcaN4qiZnXmztAGR5vcaN48Dl
HtIAuUyoft5xrWHTKz5n3yhPEL1KEwtQFjQPBMEORrGVfniqiz2ivHVzGHFGXYlCclLILO4+7oBi
KzFTtEO/Ehg/JuX1znS3KUi5P3mj41m+7ovA/mYB5j2WVS4mYf4++haOglyV8c2fhjAaVB5890UQ
mDsxMtzDw8EycjvYbUUHi9My7D44MBoqXI5QDBnFOv+yUlSTP5E2RnxXesXZJgYvwe6JzjLEqKGY
gYPm9gt7NSWNQcb41yMiEtyPmbNOWIfd+R2ez4Docf2vVp4B/UASrrbNwQNju8DNz+8dArofFxCo
BS4FSZKVFYHjasnjzqiY7GqtJz0IB13deG5itKmB8POz5obDxmtUu4d1zu9hnXH+HjB6k/cQEbKP
o04Mfhdb5OxH8YsX6xHxX4gou++4NxOfii4wDEZapCJ/Kx+33ZV8CO8qO6sfNbXBso1Iv9AHgQJQ
f/1V9O4EhHocgOPbfbJNs1hiWDtMOmWXQ0YjMhV+h2RdFSZk9wOIijonxdmMoqMUVzxxmVYGsVZi
Fdie6PAD3ra68NBP5QK58mWFnoi4qDnGVy+XQJxxtO9wKQAfoHT98XnpTaeUdjoWzf3hKgvvJfwy
9OB0zLn9+4GZcJYdlTLb7jq5iPm4ZKfO0tN3gLp5IveN3YpD+60/Jc8NTVGu5DRY/hUyWUlYd0+v
efPGQX8wColY53UYQTfoXnxDLTIZmcdm/aoPT1p9gfenzTuVV6iv28/b7/ksKmbAk6aXo3F9Sh4T
crrnIvlmh28iNwuj3ZLNRaCXPPfOlIfJl3tmSGjLRhcPxib03h3oaFT8kgeGOfD8VobgaNlvDh9+
BZKb5RRuYNgoKe8GGrPxzpww7OBpBKbCRev3NhgE81rjlL9TzU44zKC4zyAqc34u+4rnL0uVKmJr
8S43IfNq1pG9LSqlxNAhIUJJ37zLJ0KK/kfoDHCQLGu+wmIQycka+Hh0WJzGuvBUcilVAk91qifM
/niUBgHh2PLHHQFaD/ZJell/qrlojX6yw9XiefrribnbfzvN+PItU84uyjhMjT8pJ4YuHQWYOJn6
6G2KKeK89pptEsCBR15rRTKRFTcJxio2HG9arUwwNJtx6G8T5bhZaUrhSw+pnjZ4ZJtagiGBGlK3
BsaIJvDH+uDUxW1RR6M9wQq6YpaHWApcH6Yc/dgXRzY/KXI8mk4U1zXCC3ek1Z07vGH6VeNw1/tB
e1ysq/rZqtXKcYKAYQUnH5sCuLrROG3KFit3SplkdaN8b+qjJhTVXPxj1LHk2pMuiQpWriCSeMsQ
7WYRDf9dK6nxce/6QcfffWFfFKBpbeFE1MWLlUTb5JIyPq+ScVn4PufDzU5mfc3I82/rGauut0tQ
80quDf7zbEXIO4fXcUrY9SwIDXBL7RKvWEjVc9q9g6oPreKmUEvIlt275BEv9rlE50q7bNxT3j4Q
RZ56stsGb8ARZh36617TWgWn/ZNES2fIegX/rpGTAXqaGuxSrc+1hG0kPbPlKayuw0pA7ahlQ1Z+
taQbVUomXqGuSNmIn/FVxiA5taJdDBjIRtd4X3x+v7/i5nP3vzD1PSbJbEQ86HLvw1XwQ5nQ1age
rwdpo+LFeZib8RlOuZdWJuzQf8JPjEaSK4Zk4gTxrEay65jnkxijSOPYKQoDL1AgZo1tjg0Y/Rp0
GnHJMqXWTSotdWrQJZLByvO2b9my2DUAKu11vfJmPhJ55t4G1tLkLb6/MStSJ5fr16y6sHg7CiCL
3dJ3SP/2c5LJPEfBlmoiPsAVRxePXs8QPrI1S76hYPN9/6fgMQq1V1YftBbSf2rf3T/HaT0E/VVo
JM7DIBpYCyOuYMAP6xaAQq1i212kTlJKMWKI1Letl3FshFDwYsMNj1ZxdTKsAmJSPH5cOn2dNr0E
E98Z+o1/zX+fFToa4U9/irB8HRpENyBYinrEisAvWDW853LEX1wNPwkrT72S/NGWTCy3sZtC4JHc
2pxFvpH4rTt9waeVaNQ75w3So8ZH5K5bYQOVD1GewRmzhfY4idPfoyz45hMcrOy79lvAXxvkDEJw
Jm8xI41sH96Ma99SZfQSyYc75SD/z46DO/4wPCWl8SBcfN68B7lHciTIT20MGfxYWVRTK72QPIyL
itH/B4atq+J5zMC9/J1YmamYryS69l/N11pj7x10HEhjOnKrP1PVFBKD5TlApesxXGc5NOlcmk6u
E7drdYsw+hK4erLwYa4t/hKf01LEapgmTdjrM3UH3FzLXXLDs3DmKCXNCoaL/RtYG9OVsMUM2PRI
30z4fLA3ZJq7Aq9wv8cxwsh4IEqxTMq8C2yOYVJZ985VrzKvEYWkC8W4NMlJBiJplM+qSBh4krb2
AvSLjTa3bwI9GuGMIXe6ZJrrT2UfeU+VLBslU0ts1VMs1BjtNhzkkoDY3CH/L3/bVnipQmSimPhR
TTufmhIvO6LHya14uVxdfcCybnZAZ4/sKEvC/0OVC2+wXuun3nwtjQuefZcYDT9aOPtpZb15PdgV
LOiSlvOt+lhHe98BUABWTx2gHs/YBXiC0FrtEFkAOcHC37plbhcqaZBrkBo/5UU/3G3mH+hizzhd
yTNhyhkqsx+AMpELlRUyXaUYm0p2skOCIUOxXA+TAYff/v8dXwDeLPWK5ePAqKq1VHDo4aMXKSh0
pUSHzUs5OPueVGuPBl/leP5SCn642zim5KZ+7O55+KK3SB9pr1R0jYJd7fUliV9xWdvtSYiFZTdN
utPZnBZZhvg5UemSK+O8VYmzo4BAZq/+vfNBmhXgiaKzX8pLV/rpYvsu+MavvsmcBfvDF/q8JkH2
X4XunPAOV0nCNSFc6B2wV/RQ7pCHrgiTY7xer76Zw+x0JEMAK9moO34EBU6Ix3Yc8sFJvVWtnuT2
NMgWoAN6QJF28BjelRM4guEtmMGaI3HUPAEk8Acy1lZmrqXEHrfsiVREwjbi98hqk1hdUSieX4Ol
Huj+3fLMO5oLcb85Lv2Tx0PO5ZKkduMSYUlN8IqXLPIErU423riBlbySDEMIv0v168sCNS10zePi
BcdiaRoEv3JVODHaGziplbenDmr6Ff/asD+ZsHCt86yJVY03NtMpRFsJ6EzMSG1qjUZUwN7pE8JZ
t9BFzFi/1PVVqVBKv5NLQaGcys1Lj65PMulfBcbktdfRPnHdzMb+n2czdDkzyEDY880oAFSHH1bn
0p38c2SojuPNwKKYgjhg2MIkmfg0pQhbIykk1LYecaaBmv0RXisJum1Bkf5xZsx5ym/zsJgdkCXM
ohm7soVOKVyBHqXgk46nRmCiwHGONw/1og9CdZiSvGnzd+JSsuTQuwrsjmpXcz1AO7QaG5dW0Pjf
ZyEgpRRaWB+yiPyJcM/bgC5oKuiDM026dA7gM/5lO5LuxTm7njniKBxpaiKIfba/v0/xsCTC64Be
67j15MWcN75OmgExwEENekF3kni8+ySUMatq+hnQQXJhG7dd+sUqyHY0zcAAGx1qfsr+AQegs/7Z
P8wfym5D8GBOL86JhGC76P+Dwrv91s5GpW9GyhycYHjt96/cfoj7iozshKswSZrfpmnr25Z8OZ8S
1Z7JEE3T09PujRYwLGYAiQIrhxoILsSA237ZTJjMm19Ai6/dkUfL7RliWO3Zr4oMHriJ2N1RGzL9
Ugy7CzlUn4WF/nDSi2AXstg23q1hkfUkK6FHh1qRGe9b9oOizuWk5MQ4FLYckFkULMM02DwJrtRX
wVsZJh3swo5llScCh767ym673Lt/oywLuAGcbxkKR/Gnp9me5rVqcrau5/dkykZicbk7HYyVN2a/
m2NJhwzml+wlFEvyPCiHHieaety8r0CnCt5qH8ayH0hTAZeT/SmBM8QBBV/fSyeY0k7PocRDGK+T
CNuQrvp3zvrwkLaj/Q+JVhuv81upiU5UM2mfAVpxiCr/CV0LHfnBUg7bXyaUi+7zm9tUtiZ+ixKj
sNbwRI8pOLAToaHOiVG4Sdm6nIenqFBqnTlTOBPOVXvrulw6T3p4gW8WcbShmQqMsrkgI/mk9iv1
tTdF5glBXLuI1J1AjouRrGioKIit7+rYvs2hV1vlo2dQnuFWWb0sQT8SGjVSA1ffkElXls4wzYSA
QjpvbLqMngDn3lnXxDrAmJ0GZCcY6f66fG+/jnb0wG6Gi0Uj2ogpqMyoJzTvZHmzt+/FeI4GgWUd
wyL+AZsokqSsdzfYpcCOv9eqcrJgHBHQaqVSGSN6BylDQ/MJ1BwTgkk3QJsbg4qD8462RHkiFxAC
tGjkCif3lBYe66O3WR4+8lPc+7SRIiWMexPV43G5uY6SduhX40tUesZHZN6G6ovyYR8XMGXlj34u
0M9e+OQtXMxRRHrxSxpFzG7p2qPnS0xLTp9ZQWJ6A7SzcCY0MDcBVdltuhKUuOExdKQNBYDnMbiI
7TLU2BHhpw7cqVR7ihJBMFHOiy1hCQq3hD7yLBg18QfMrBZEe+x+IAO4bg8Z3e+5yFjwZpb9IWFF
OMX2mQecbv0TegXLrwiSX+HWiq+R5ggmdt2POgpdw0cH8xPlf8PWgKVex3S7rbxI0vZnf3fWMCUC
sBYnszHtJmd/CQcu1PazV/xNQUcc4zR4JlpDxHlzdeflRU/CW2gvAfcYrssUBYCLvYnqXgjfirMb
far2kDFjnxCwrAvEmfhTx6B9xDGuTX65UoXLWdT+YFhqtivN/N/DRbLx2k5joR5qvh7GwYLyCRCl
LpdHF63tCKPApeQtZbDp7jyasqtjZDrX1PGOQW/7SbxS0KKie0Tn+OnvHnbwhh10AHKExowbTb7D
0lvPV1waxZMxCVuSZ13QZWe7rHpbBZFvFgPIEIm2/B8ERoBCdy/0VHDazk5EAtB+7BxVtjqMoFX4
6iogxAXzLP+9+dl6W9SxY1969RBf4kf8EhfAdmxw4jctc0RdUO8gmxi7DDXYTynN+AIiY6e2AATY
/iyphwvbImdXQJK+nyRtcx7a6gDyvse5PpU86BZr+0xnum59qxA094qmkXPpaaZlxnWdl7JxUoRf
kZjE6+OMcyfqSXuaI6mWMqxTraHYvNkSdeNtnWrjOVtGccQZFLNs3RgOFq0IKL800eVX9ge7xRxQ
nkS0nhHBGx9E90gf9drvZRE2kS8UJ7mS9Qy1njYiVQSArS1t0xF7Ddd6qBdxy+5uUoPuUUjjJOoV
wilWCbrSQD7J0EdCn5e3rq4SN/pjezw5vcjjMNKGmOeIVdXBs3RxUSm4YRucK+Z3j+I//8XNSjD7
jrrmh8crWiWJBMk0nHDaJa3sn0J6HBNXBfsJORbs6uu3Uy0KCcYfW7JG4BMsEJMSFyxFAi/oyihF
OpfTb48rh/oqWew9+xWM03jFpdaUEPj6dnAsPTdPRDKm2kOGvxcRI7KfivPZuSIcriaIeSJS4EnM
XeN4ELEimTQBny44RT+RBLZ18mjoKM3NvSsm1X4OnxI1sSOSx8KgR+yifW77VFRHm+K73OXUbN1N
cEQBCF8JcMCs+/UMy56bwOmV0hlbZdIRtcZi6O0ENDjA56n2eUUf7UAtHQ5s+gbRxHCS+9RCTuLl
GAXGCRy/Br9l+b6FFdsxoMWkX5iOiwYW9TajZFC2qwjj5fczMvqyxJ4wRpO9xC3eHqEWcfe5ds1W
BRKrmzbBg4riZB1isANAT0pnCAawjt4qYeK4CN0fVOtDlTSnOWF3FwT/CceZFh1kfKN7Zx/gAhuO
LTN1oBDxSYTjdDoyL1+AXoRtPaZHhKLPnHYpm8tjIPFtJIyicsymxc0FrR+wfnNTAvzANCw/psub
gfC/9pp316eNVjusAC+bk6nZw4Pj/xl8J2JkTAwhA40zu2gfUXb0xalDI4Qlh6r4LiYXvyEsI0v2
fg+s/fQxY+YlTLZW8BoKVZEp+DMnDLCWI0WG+LKAcMsvNEL3xN48Gs1IVDVLUw719zemrDn+boVN
iuk+I3yswo77UxJgfjHohscmKDacwnkwbOHMe8fiR9bDix3mlX4Ec/u8du7oIxZmir8B7Tcc1iVV
wRzFBYlcFMNzdWVsDDlS7IFRdTTK05Vr4CsFMfIkYtf18S4KPaDHGyWG5xy0Q9UmrXOxbvooUJV3
kkl6nflz0Hb0XHsga05y3v//5qwAs467yz5C39HTMW8BJjdO85j3ufXltw+TZMJACvpdiWP3bnMe
4h2fMuMfn38TrcVoMF3WnbG8pKZI2vTlDk4POyAZRkEbb6Z5E2pmHMszCid/zp3dpdMeCHFFWrJV
RQ0sk0hLX0ngCqhLSO+NriUcmOHgs6TcN+e5zI2TDeX+kKK9Z1fL+GJUtrYaLJHd9j8vVCSxZgoA
/KTHGxd/bifjWgJX/CBf9GvI2C/efcAtb+pQ/desiANpD0X9XR8+l+zXUKRSxMwFqGR7bJH34BLf
SG+4XeoceaGvgwKLM3P+XE2lmHEPdyia/ebtb9RobgnhGFc7iecANtuCbmanvsM42AFxMO3mWFz8
3KyqQqKjP/blB2SGJoRwwJgwuDwGxxCHJm+RX3pwHz6ya8wV9JHpDVhjKbuWH+ieFgGQpNMV1Fua
4l9OU7QzuTweC5q1eeGR2NXJrZgs+/uFQODoKRTbOL5oog7jfyxpFuXe2xFv8R79Ctxl/WRuDvax
ETiYJBDtbcRWpJqoVqdCw6r3LvPMWcb8PoTsinjez7tZBX0nlcjwEeOadoe6NvIOja48W0a5ObF5
LANxZrvmbg980iVes8E/i4Nl6rO2BA52FOGsxhpMVHcU6Kk2s1qayWQ6ngs8FtwlAdAXvfq2AiTw
SQ4xNwR0WX9N0Z0lP5aeIUIhTA2etaZJJLtxXdwG2/1K0tFReNdL20j/eknL7HKppRqxy38nk4Fj
AG66hR2LmUoLK4zyYhb5hfCLJ8onUGPHMeRPo/LunOpBiBuqgP33TbZ2TDi1N5CQ0wJsF7HCYNT3
kSULt7rWVmMHdEHVIsQuBCnPkNcP1QJg0nZ1exNRt9V0AdxLQE5uhtouDAawCI1dnkg1DliQm7AB
IKlLqHfciS83sW0wKyz317cTKXEEI1y2eASpM4LDwy4Nrd5Iq+5vG6KrcMGNPy141+CHNuOUbILI
UyDBx+TTuqPx40olOFdgMs8/B2XJSS0hiSKaXtxONjuNUPzHSMHgTjqeVsAIwBZEF7lt369UEoRV
SIazQbwVz/5rsdFmSubP+rNMs8K1wdoYLTAMHTWQjv94/4pWuKsPWylj3KpGnjOx7Mvu1lp4N15b
nM4BT0D6O8gxaTNE7Y4V+THF4TQSsRYR40DksVmmdTPk+NuwlyipU5ChrrVE2Ryixb75xu9scLiM
kXGqSy0vBuuPRKRNJyK3k6SgOW8yd/4DY/b4BB2G7TS+nsXDDtDGBioQAyFHotWP2ncBdRc81qxc
ZdracXtY0S4T2XGDMgHxIRjmPZyV36tf++4A5V/Fm4nNi2g8FeEvJT5jU4g6gVQnySpMuEHPv6Ct
97uQh2IM/SQ/WQ50j71+zi3yhxvbLwhsiZj0pHmYZsM3bh8wD8sFk2TtcRfcxmI2QaCenDJcUNf5
fGUgq8o4ilqtvVGADlFdXQHzTlzo0YE1aOMcQ2jmB51QnJmT/5zc0w80FgVQ7YCFsCbKwFB8BRSe
P/xVbqBzhYnAfkxoQDNSCkU4U2Wiy7b/WHRBmJMk6/xwZQoAIj1upCjVLsbl7ySy6QPJfqEZMiBE
rNoB9y0DZgIhUsGlt7qBycw16zlJrBy68znHEkKF+1rFnPshE74OEVXbGTaHVb0l5Amq6I2s8Ltc
HInInh8/q9y0sN0BbQjRHdHbMZBq7ktJwVTknKOqDUBjaEX6HWbgXutSuzWFgVVckmnH6sEyBw+s
XwMHj409xolJ/u08mQKPjcoi3mBcsUicrnOznE6uX/mPiMAmlznfA0fvK55Ymq6+6SSdOcTU9yYp
S7VnJJ/rDvALWxK0bw2R29Ucf4zjNLT8jv2fZEAv8KwBjsO/3ulGWEwCejx4Em8WNVrxrr5cTjvm
qJe+0boE1hnJDuT9QLQ7iRsAd8X6QxvESY1/rEqbive9nmBXsGfkmQlilD9LAlvvlxkU9TbK3GW4
dQFrKglJOCdkANTg/DEzoIcZ56pxCrp5ox+/EIaE6Ii4M5hmciDbIctkmW9gKsWNkMmvp4SfXaaz
z4uCAxiXlXr+Ex9JC9kCcOfdHRWzmODTPEiXvXsF3x5Qrn0qB68y1qpuv75B4JaKB12z3T2Bu08c
kw+Vd9P6R3VjwgZnn0DtUwrAXTBPO9eDK40vsdK/UX7M+CLNU6/wJPQTrXJMObPNEZChVAwRQye7
q95IJgyXL/QnkxoQMP4gkT8oxkeO3fVuDEIvTlHtPRM7LcHmef2zm8t95zg+RT/tYSwUPVolFpG8
OpOWKjfmeB8xJZ1njkziDIGghlNPuTkN6ltRVycVXJbi9loMd4YJmFNCsjiCm3NAWCrtE4jSAXk3
xWZ6Drtm/8TNvL80YS+IKAeYdclMqa9P5G5+p91R/hXDltmAbD53gm5G8M/WOMNZtAvgEuLi8ERC
l5KYBKiSX6xgBOJEEKKM0N4g+x4WLSgzxtpA2Him54QLEW/ZjBtvwSF8MWY8R9MHQW43i78xqlpW
fjs+Q7BuniF3+SDoCsIe03cGf9xpcClQGAFaaBgVDQe6iG1e8RI3paZ9tl3ykVwtz2F77iPfsBbF
vpkxQtF5kRBfRu5z/YpMO8ZeLOJdhkJQKpUjeLCObSeaCsF0pIGed6q5uWsbG9MkDtc9ShBCs1rI
aLsbU9J9n4EXY9T/chXqQ/RA9BP8sQc97NT/QTSNCDkvvXAH66c0N2s5qDYzpLp56Aeu7GFD+XJb
qrMhH5ArfGe7N2E8M2FRsrtcj1O7/YxzfE/uIx4/RgdncLFM4oqHY87mzuDpas29mNYU+2WlbUhv
pO2stBcntPIe3yDSMDExMjnZ6Z2QdqqTL09dsWEWiugrKszNENu6lW4P4nP1wj0oHTyIiOkF3Sxp
lCi2tHHblIPR9KBdlB4S4zybI0H9ZM4pcw2iOOxbYMbSf1TYHnwEuYtY2gQXaHDDJq4mf/s5MktO
lqIq5WYBekggO8ZgaUcWd0LW5bQSfb4eyO9Ymtv9FiDq5OXBGnFH0fAAKaQuBeEFhWQ/IqK/Onpf
1oJKeS1t/MtZBkqAqG8pmNBUn2qUM2zqTRM2xpd9u+w9vSGpFRXCqui/ptX+2VHV1sMrh2gW1IK5
VE9JXm2SuKOUNkP4eydXThk5H6hHr78h+/7vgPnS7URgceS+g+2eJQKEF1joebhsG/5tvuXKf4qE
kmsvC6jGzfY50oOP8I7P9QA/M72+cCWqVNKtWgcC3ikQAn48XoUJb5p7PpxDfhJhSFwvcouZKDy8
QLnJUUMD8TKHsWrBeTnfVklSRR5OVb6V/YBYCuGmv87R8iF4Fu/ir78dMevLcdXyHXYqAuINwvkA
5/LAecDyzK7IHeUl0+z7Z9epBAZxUMOXTCd4/3/KyiTzOuUpyH/AmIk6g+lkbrXdd30JFIEnumlS
p5ZIOv1yPupdKwpgzJHI+CrXRlo3+ldNnSSDlhhXIzby5JekYUtBc+yE5h8j5PM1J9vDL9gVehW4
I3dXAv/sX7VQMh9UDk7/p1+9m2X/JJRfhGOP9HURUneaN02CqDtV0mG0q9+HASvDe7FeNjM91nBw
H/5JMDxIyzaDqLj9QkDZkG86dstQCLGw23dQic7AALnbw1UWC3kZtVL7vrVh/djPxTFXvwNSBEnN
p41Nj1uqvHXfbINm7NpBBwNbvg/rOXGyEz6xRW8/Won4ZbbMXCqMii2FQDJ2sb/ySaj0CBGdj9cv
yAaS69PW7hdI5Zs1Nvkxgtxtfqc1sxQoUG3QhEdjF0eRCxulOW8hdhdvayrgDmLwTRPPZyYAgSxP
XXoo/pMTIirw89gRGMdzU3Bi13d+tnn7CvNcu+Jfz7r912uviIvmExn/rwfOt7p8YmalP5jxR2nk
BZzTZn5397h356qAzbpX36mSGN2gU2mOZtXE1NwIndsWgVn0S+CopZT+/Ao7/cWRMAfirf89A0Ri
j0MnmU1dROD3pWbMs7MPX/Tl5CdSSCffEFgz6SAZC5wKPuWjzI9L0eBsfSHLF4aeLUccOKW7jBCz
y/6H0Hj/6Ke1iUfDmTkVTD0DDfbqJMejtV9rkN5POgG/qIVa7enMUb5ZjBOcUawKPtd/lEkuNSOt
EfH4Vm7Z+Y12CVemHL/sQ1uji/LjahYoSRHWrFcwm/gNb3PlJY9jYc6Q/b02PCw41T2qg+kJ2/LU
V2tZH2LiMRMmGcSePJniewTqOz+eQ4+Gfict/deS+dJmbTJ6KfYV+MLgn2roKhoSGz3BI8xInA9x
x4UjUJz2Ff6ITd8FuJq3K3ACmBYd5RmPbdKOcKo9S3OoOeKjkTAijllC4s4O7FZRBVbm/oxOrHes
YliOwt94h1WjeJV7Wn+XPuXjL8Ov7e0eyJLaPdzHKfo7i1ncycdwidn/1E1UNcvv5dMrA6k52YR5
2bkxOlV79VeepFaXR0N7NDUNXQXD1KgIa0Wo62ltrCGwo5Vu+gNU7q9C56/W13JwGJBQJjuw0E+z
7Z8mY5f22S4la7m2UZd5zgLLxxkrng8vjoJzwstyWpPRjU8sTYYzoanQ+6VIyItGF3Rp1scXXFwM
U/zyER4HuHlhJwc93I5IA/bMTFGFaWL0hc4kB1WC2S9zebI7UIEgP5UJvF181ax0RmfAsV1P7axS
aGkbGdRrsT1vH8A2n+EB45hzC5NghlIzolgfGqgxmr7hao8slt8BQAC32/iR/EWgUOY+1NeiKqJ9
KvkI1dpV8D4pYn8hzBiTU5HOyF9bUK14kb6GIhEzof52ao4Pr9jyPj+W7OlsWCdj3foUwc1TqvQR
90AHZNaR8vdqrLep/KOj6J2c0vEeuU2wFYcxbG/sE8rKTq+1qfP/2u5ydKi4rqIPt1tvry8e8LBz
jGrKwLpbQMEF6gurcc02mpKOXe3uK4CAAoN9KG07b0VhX2TAR9GFBR1Zsf6jCB8lCz7fqSxMtMnE
m9cKr7QaqAh+kycPOJPQsVatG41GRNRkdOMkVlupkC5Cp3PDLjBZrOxuFesTFq7lRoLGoyKOobDz
Xnhq7q1qAeZ9hRH48s8+RT/zXw6Zdh56cDdtgzBrWEOrvhaIvntik4vmA75BYq0bzH5+tpYiVSIu
lyPaRSoDm0Yrf7Ft2jS8OMTMtuXXtdyc4NH0zLue4VMWBCicNZ19VgUGn4O/j8l0+Pnp3JO8kfku
BLPdMiurxyF82BVcRqL3YA4uHjZVESglW4CU9YxO4CXl+O+3qtWxiwlm5+VXaz8XjrOWZ4xrxtfM
+rtF6TBecrWDsleN4foXX/W2b9fqpMDKK2LSQ+EfPVZ6BgwoQltBBdOvpQnvDe/eXNQDrEQNOEZE
jsuAKbrxjVi0t/bYJwua6H2u1LACljHMiTFEmZ+vcjsYwUs0lTTTzTX8xYWv6eZUJFsU77t+c6JN
f6l6giw+HIvl5mYmIvkDZT9i4SK1j91x2nPHzchgGrCIoE6NCnYTjy70E5aU8liNoqVF0JfD817K
SuFx+YCj3rYf1LeeqVeG6oproVWaci0dM5pj9wpSdP8I6J8IC4RsafzJvxdNb/qtWGjjzhWm9RWu
k9Ag9lfbzNUUc6V+jzgcTPIAJnkPmxwgovEo20Mqi49VAG5DbbqknI1R+lEoL4WEtbpKg7RAbRRS
oJ12UINK6sZSMpBxllG98yAtnfu940qJK7OQHwCHnF/rm0gyV3kbLQplV2WFWEl9Seo/GjgObzhf
I9cuhr5xfehsKQ8N4DLUxAskLq/nbRSLj83itM4lqMeYlHHcp9mDRzDbBi5REpFVamRm5y/pc2Hw
ZehlWMwdwDjFQ3BiwbHK7+yZPUtRihzYB2LcsOAno4Rg0HcrBRTSJ1wh/jriHlodFeeoSu8AN+mY
i/mPNFjc/l+xGwzOVRhvCK2D3QhWoFri7yA7/uQi1ltPvhtZsF2eKNFUHpP16Epjv12KS9PGQ+gW
Vgl4vJTUrpVTMEWklUG7epEVCOPjkpPTZZd68R6pBWavr2q+8ghcVvxd3cKKVK0u7jckDk/7ixgl
E+vsIk9RsIAraK5EPtOcxaBWL+1Gs+sson+CS3Xxvct4MUe/gZniFoZYDzenICpgZWo8xLHL2QM3
mdcZLcF5EV2H5YxUEcEPC9FiRLCj3onOJcP4BRfXnX4uHNJ/TrRrAE9vMVr0wvqaAfTO94RjGW3y
5F0OIdCXsTSp5CZPDU1gYVNF7rBtqGlXZ06CzNroonXfKPCDRemHID5mIlrYCQ7pIFHIgtKDRX/I
NmQiw0xMzSnY828ztYMH8+IKQfA/4sru6pmb0XKj6+Dd60laDk2nB6k8vEIdrUwoSow72GE+fs6Q
9nUhQf+j1d6RgXMZGmu9LqXDJyhHNFH6c76Dedion7nSUCLmgb1bMVPAxT1OkkWZtaywJLh7PlPc
aRV/3C3UTNQF3ISpKrpnYLg2WMYBgIio4sj3PMgYOYHwxDwOZBk/FW3SVVCq/GB1ru6nNXr9nQ9h
OqL0DzTatgfspnPGx744Kq7cjTb2+z6OKdEdVUOx8TSo8+Bs0I/VpQu/CvQBVqoB82BxU3GWOywZ
MTU5c6emgmq7CPS+oyJkiqih5RUsRx34dtjWQvjDL+DUQaU/z8xjJlWSUGfmDxbXhr8lAklsJkBZ
JAKWGvcBoG5yt7B76VGSWC2rohqDlWjHJ8eIBnn3Y1LS8QKXK3KEE0xgxsP8S2pjPSZaMtOF5816
V29MozVC0RS+urihPhLcSyryT/dDEO7tc258EKi0oH9+9HVFd3Xc1bltm1RIQq2ZJAio+TZmg1wr
L83LM0gZDm3/uUb0K6ozw7FNzyIK5ZvaKSdBkxJQR+fhk11QMNgsmnppgSMXUTakNppA6ZqJaC61
xVjjYbOhFOTMJg8JEDRWj44qadH2oCpCqMCVJmaG2fPrv2aUAl54/lGwQfmbmhMryW8xklTV5eIx
lIxe7DSvuhZjR75K3qdnTm2cbnJwDHbGwRK8tbbIA+35nDxwZu2XV8zNUvXDmFRZYU+xdmfHvsKi
R3DpX9GDToxXa8YQDCAV2obkkCg2G6b+HIQ1dGjvI8yl9ExWEL2z/OfPjBcKskkp8QY5SWrLOiQn
qt97OPLBUvePSBG8k3081wtCOlLYA6J9n7aInX2HtyH1MsCKzakTmka/sAxdwoOlAKgFHLU4OC1o
5Jq8cd4/smMsjJqEYtF3b6RfY246qPKcgJlZY/weLynGJZXi182naL+i18Zxfkj5kpGdA9Z7xiJk
bASsZaUHqmBC9j3XpuLeLAxo4MaDKwnlzo4Pd3fol8xgqYNL11F6ffJK78QpTBIPg+2JV+ZZvgCE
GRxaDcHmqC7OY6B0ssVBvcKoWxRPkFEEtzdDB8GJiO9gBoAvDchZa1BmQVx8jltMutWmEOIri1Ww
4Fqf7om0vItiw9DvrBInM+5FWZZ09+hhcDRe2VxSe/EGSBWNmvccIPefYIs9AoawDUrytd2qjni6
oS1zy5rd1ifv3jlmliJHPfz4ILodzcnXw2zDpuSmRaVIteNTn78OHhKBwy7f9694C5muY8If7pJ6
vNtxT/CegQaul5tZ/ILoYw4qm+KG884pU4POlnA1+qHslGhk/71GcrddjzXpspteMmcCftUiEnte
qt67zGSIyLE7TXj5iErEOHfWcYc24lZAdfue2V3orRo5ogwbb/MltrjiKReK3NCeVUwNlJMiEpgT
GdstBJtPwVg2wuyADA2ivsqVq132W0Up1GXshar9w4B9+u6BXc6vM0RCirgwkNdT1neRLP2+qRs9
Y92g/x6Afjea31CSRZBdx+xx68J1+Hj9e18GysodRDEA9pn8iE0WmsgkpwS7Gca31FxqAIVN2R0G
O+kcgRTPocPyTjF17Jqh5OCu6YxVd2BNQJME59+wxcSCTABYAIaNntNTHvgbJcT/60gc3rGtLIB8
dachVv2mhH429xCJdzXLbvwVClEP9Fl8m0qTEt+qdQRUZ4vhl8nlD2GdQYU8eSHH858oFPM0at1p
Dch4wHqQ/GwReqo/0M9D25Cu1Upn5q19JFfTITBI8dPTMOehk3dMzfLdGoPK9EULRp++IfSBmPxj
Fniv01D+5yV8hBZidKnW0g0rIIPp86CbCKptomcr8dVLAb7ar4hU0NbneurW0PpfzTJlB1eX7Fq8
G7R/jVgUG3Mw6OoiM/67sQR3CgufAf5Aqnd/UKAiUtqCTOXqCPHlWVCzQY3WOB/UuMJqDqZpiz/t
mxKF0IOrzMn7ZGtbDbvj9xhCS4dF+XVQm8c067JkZYpgc8QdN+JQmmcIGLOVYeYLWsUBJhsodU5k
TTjCqtH0DSdVoGHdT0Mie3rPP2hN0MrYkYwcZ2T8GtBIta459VkoVlnEawJa2N6W/Vz4eO+hzoIA
e7zNpzb9i6QAp6BRGpfjM6SoFBTi5y8deamEr1F7YDlDQE++tdf1nN/usPR2UTXFfk0IdvDkPsvy
9VBT2BvADN/gkPFl/L++VViasjX17pAP6sXEYUcg2z5k3Asa5UNVpRMRbN5E/Ezb88dy3Z3rPV5k
TjfcceWFMNmOfUeACvAFVslkqu1riz6Hxrc7lfXkPZupnHi+EoiFsqxTQCaqkOvp/vRAjBOZXzei
vgezo0u8lCsJM0nw8+yPCRnvyV1n7HKQsQHNkBWxQ11yhudfZ5tN+YYU6TglHNYly1qlSNDdFRhL
tn1ncFKUMQ84zuBX0JvIeGCGoAIs0iuqiFhloIuHZ2CTesceEvRXURMdMi6pcHOmpWTDA9Z+T6FP
DR5CqvWevF7FOqPeZqd/jHJxXk7viHfPx++RM0aic9ZVfZ/LdWadabVnoVmp5rsXawjpCAIFVIZq
eaECVnUMeW7VcZcFe9P2b7AK6LYy/K/SNPYAb9Rq9x4daUK+6aS5asLRUMcW0oDvqCpDFnAlfTos
3v5w+mQd6L6L/fVlkb7ygwyh7vux+vB1BCbEDNTYtSjJLUij/06HWhVfwdw1fTqT98/ZplE1BlOK
qrIuMgZR5s5BGUeHzggMR5ntkuTxmLSNc0N5A8iycZnHob5c+aoS9biWcPl713jKkfzqtFgyx+wl
n0VnKirW2APjPkzG2OsDqZ4Jxa4kIUVCjnzLdwYj/CWf+J8Qf0bmSw17IXoTUJpiKTpO6/TPRs7s
unNlA2nl5SmcAY/rXQ51y6FzQMvRAlnzBmmKJP2AzBTcVOc8/ynsEJ5bbfmRP0BnKPkgzJ65r9Gr
165u54RBzKeAPsGPBipNFGP/K+d2qEQNHIQ+WeipKVpvEgjWsO2XbqDX3werI5N5riTL4ij6fqNW
pHeop6qkD14TvbQHir7Y2q3vPrh/tJ4Avrf+AmNehnbAJf+ys1v/yGnPa1afXG5E80NSUA7QxF5N
cAuvss6vim92rvaXLp6RugV3kWfBGZeD3qGfp41Q52juxc6i3eLuBPLcO8F2viuPY4Tx4Kw2M/z8
+JX4TlFfS5Af7xF8jJrhvbrM5EMJyXThiSW+zQlfPgCm/NZSCsjNrr8JsKQ+basW15MUm7CHIfBD
/CV2rprl4Y81owRB82y3clyASJbprM3F9sonAeAelTTYGzE0srH19YLwfkOrGTNmSlcwGvQn1Sq2
0RdjAYxspO2308JlHo1ZgyqUvhHu6sFlAoiYvLa1WAJkBfZ/CSC5oSlZqxgFHDL55sdcn0nXsrC5
u1XrKRAX77hqcyHFPmaPNR/GFqgSdpmuRQlJ3CPNNb1zgHL1mJq3n2y+/5TpXCNihcUSPT2zlnAC
gXe/neC0RIMrieTNwx1R94LiyRU+obsN/Ka0fbSZ2JxdA5r9vCwn+U3bWM57DWmJTCg35+Ai5r+x
RlQQXFNUCKp5eD3IIsBT2oZAZymC216CEFZtrBzq7SxAbRk1+Q5GuV1xrOguvfS5xX0SUhKwkIOh
DXObbmqN+W9VTncCFwBIDrvO5YN1Bixa4CWEaXfRaXpXgnY6AY16KqpaXSnJB3+QPVxkIQ4Ue9T4
iHHXcA2KoBICEf0hY0pCddtHlwxQJXBPhXxs65njOQCtiDqwWCMIU5+swMMfMc8cGBRry1kmd9Df
zI6Y1KpAlzqijxOLJX7CXKd7ExdHua/FkYoEdXj7VwHv1HaIA841BKHfSY8lYUSGWCOgU0ETX0Z2
ydyEEI2ViBneIw3Dv9e+Il01MeA0nU+rhEZjITws+s/X7OgN7fIkg6XiH+ofD/jbLFxC9Jpy6k8u
WxzVH/hQfQHWu0Kbdout4rKUNMzUhyRR9582/inNcbD70wlpV3Qo5zkYT7rmL9uFZlgrPr5o3HOZ
KrOkPXvH3AUx14ePuH/umTIDCpIGaU9WRJY1q8F2MnTNoAkOfxTCAqOiHwlaZcVjTKa7ogKWIHXW
9cYsCNHvraPpSlDFsFqipEKiXugsvbT2TXeEhW3ikWMm01MnpLhewfv4KdbjT8oqXKAJs4h0O+/f
w4QRsvd5PZFVt/8SlMXQEuNRHijopi9ky2hkflZR4VM7ci5DN2AHDpPg9e5MDYrbgWs0x+3/cUFc
YA48jksChQ9uCuQafKKq8P8NlyvWZtU26oYxHfyuhpkHefDjLegKzur2iuvHw96dmt63TaA1u0cw
3D3bzrfOvBsmbC+X5GyHwiTLPgLl/cASLPuFmFDMTxDzzyTzDzol5g0fDZf4LYo/h4QVXMI7/Chh
wJBBMICRWDSL7wY5tPdcs9+JOYER0E4sSPfCgnpKOYtk8c+JXpMFO6dQdW4IPmpONEncZZ5JuDTt
qklwmCOzqcVpQMW12IfraqtKS3eB6gBbnVyLYZxwi3yDTrYLj0uSQv4tWWrwRr5QtmN0Kk690CaQ
sZUfa7ROX06LuMKV1Z1A1d9upggFeYj0QnrdMUyx+qpxYrmNBkJyqD6zVxwcNKrVR15pcKQv2x4y
ojGzkqTmjsaJtg/KBmiW0/O/w/jcVOHtYDjyjqiKIIpe+N6q1CQ9BgRlAmjKhiTcjIuAhElW6v5N
Xxe42qAxk/U236G5KgZaxA6wd2VjFoOePsqOLqzij9ubtAjZrB4i/AgeaSaO0UOB0GSQpk9Tde2m
UpU+vyY4Gjr314sAD3i3S7Mu04x5zuo6fhSVuLmnS6dNRC8+mfi4ya0flXqu46loQI4ppRYbs1bJ
fn5XOf8nXyuJkPUT+N0xliewY0trYTkk1jpArqzE2lkNackUhNpFOAEuttpTyy3vyBKg46IADgBk
VNKZn+pfmAgO0aqR4ITnAlCasPfSjbmJipQIFEj0N6P1wBh7ayrryv6TepkAMzLrVjCeLFrGsDM0
aZuuTsLlk0tQMLRgtvE+D3ypg8gnZVl4dFIJw8Dzv4VzdsytvfX2RdTJA7+Hd0nMAvrEFkNk2PJs
yT1kBiwUta87pfxetg4nuNNOBV4y4Z7NaO3xvSZ4pww/dISMT+seyzd3QSmTnsP6i74lKHE3KzXV
8pigStpxU1TtNoPhYKbpbutGj55LjqYq/ZBw2eOQfKyzc7LNX4vmY0gdKE7IFuqX75vorth6P4JN
MQfObdzhD5yZNcl7UtBHQtV/iErDyyQmf+FZkTpSbiTaUG0t9gv9/QmZsh4UyyaluQWcms2bDOyo
9ZUtJrYVb8z+eTwNG6vGL1dc97/Skc06hvFP6/nXhzLKHyEtzh/nuvB9eHmARuGj8OS7nCIH6rkt
70oU2gQfKXtJnnyUAM9194VrVN8tz82q1YZV1xwmWAXTvkyRJE4D7pqd1kaOlq2hVeDDmyVoMQii
qH5CGMgt2ik1vGLQxbrEFwc2JaYU6bhfq4y3vIc9JLruccd3/CnyAywOTGnjL6FX8sTXGoYDnsZh
QLayrLijURwWquLVx9L8yb1ZYvVIebzK7pQAqGNX4eRScr1eD/7wQkAU6zUSmfuyhg5ness9qdiY
w+uavByTzcjNFc0YJSh1QDjLMGP6mIEhaTloiaJCTwf/oj9MWFoUkDw6WEbXroI2zi8Mx04bVFyy
bMFlIiAT4Y9y8S+bbnQGioKBqLILP9lkcrV9E/tFg6Hq1APQOOGBCUC4VmyqHnvvzBrZ5nHBTFeJ
TtdH0PuUbtmudRBAMyfnCtjV1nAlshXPHVzBLjpcf7WDfSHC6i/jmA9+qgOzW0eUQRwsu/BjXw/K
1qWah2VhRjm0edu54wh8HiABoug7ksOEhCWL2vnfSFXB/xd0ODAcf2wlD5uytfEOuv/EsRmA6PtZ
gKY0FXoqldT34hC8HgLJU4aLt7ElnWEFBSqFlMv1j6QDwpZtE3DH8A9l/oP4okaam8tJjA9XhSbr
BNPTN0gQ70nQauTx3xyCFxkOZ7lHyedU/YOc6no44FtsECZ7Ix4cGyhhQvJTIsMh7OW7Tn4+TOcV
sBDMXcLABDe2OkbszxLHKACyZ2x7RZYdYz/X82VXClIFe2K4yMg5oqpJ2yf6gpOlTS/+ikspx2by
h9JXQW05sCbeM4hzPBRKjh2lRV/tVmcWcrmJnZuvkc0cW1m40hyw6b8Ew8VeIwcv5YeXxSR/yZas
APAUVvaEDQ6/wZlA+xCNb2QRRPlP2+oQfa9LfY36KoosG0BE5s2Nl+APJA9aWzR8VgFeN4xtHHTm
fJTY49k8vci3fPykw37kQ+jljHf8iDs5ZmbktQ7MRIUR10j7LN0Kph47dZThNyMfZ5SBcyAFQcuX
11wD2o+bL7Ooc7sLR7UIoWSh2KxN2tfO0Ro6SjVp8m7nK9pm/s25c9IlUz7FvqzkMeRI8TAasu4o
90x8U2N6YRQEQ9jua0Wjf3X4gbAS5Elf3gNiLn5K36rKiUwRQBs3j8dkTUA+ewITkl/1mePnSXzs
e7IK4LekKqZrvV7f85xGQCVPJR85TH9/Dcd/ousqB+JS47bEvh/roYNbxrrtyogu7XHm8A/XbskG
yj2SK+7ogyXD26MZCfshtKEQIgp/dKF4QMabJ0kom6rLSF8W8ch4L61wSs3/K0TGjH3WmPjbtj2D
5gc7raVO4LieE80ZLF5GKXJ09RWsRbXz1WLbRXteqz5Yc/nwcCmUSV41W8B1bSxv6NzVqfHDmGj8
6Hsola5VAeD684n7jCURg0X2oGq4V+CO3RyxuFNjYcEC/6iwKvOG9ENENyiOM+gZ+//TGtwZbQvT
EJmLo1pgSyP59KMReDu3dogckTYL34r8ErgLdufAgNZKDim8pH8WO/Y1uGi5I03hNipitc6H8eV+
E7jgHe9O05+sA2A3MphKYbgS8vJRMYL3xRPLDZrc18NLwiRWyrsGw3uP4eSDIj0KnGrcBlgnNILZ
V0yBuwagOtC/hMJCcUQR3xA/V6DQl+li2VJ2SY2w+/DHWj7rsWaWmfPgaLQSgG+eKxWKbbJCjlS5
EKzXi8fnrLIlKTxkomDT+bmkOl//BsT3QAI+sb1rxGHS7OdqAGyBeUbs9VYP5oEo6emM5hMFvz5N
0jUDhQFxuBcYHcfGdce7ejAlUAtHDxNnCvd/CSrHf9oN4xd0us10tfpFgQMLiSjUMBwblkj9tjAQ
3zTaLMi8/x3NYkDeU1IuG0wbxWY/3Sp30g2VPSpZS5vCxMKSfdBnfrm1g1hUtDwpwBVrWOwk3p3R
Wmt8XiA1ZZ8WzYAXOaTuO7ASLK5P5cb0+BmRuj/3qwTOtDOWXiEbYbxs1bTvlYgsZQT6u09rwdJE
ZInFdUc2UO0FTDR3A+kFyD1CMFbPf1N/gewHiDckXNTgcEIMqeWRZeiWi2++/wRO9FtWDnvB1H4g
UNtuJmMPkHDN0fH6dl4CCgGA3NbDusIel5hJGsg2LzmZCAqmyeS8VuJjmzLyIrHH+jab+/+TF3bB
DYrRzhWHbGnkHWky2uIldpP0ox8Ivu5kwKyxwKGbAJCTZMvIpcFDTHKjM+l5Sbq7ZkNcq1+pe2do
zQQnuV/4z9V+0Ynvc1x89DwWqpacv0XLTnj7hANNCD5r9eOzr0oPNtCa+CeLWb3pDWapHAaex5eh
re2VDCyy1xhqVkKLvfo2x4vHPTQyUcL8VXwJ7J2x6bjq68tz2Z4P2LgI8i6bW9QER/vC742RtaCs
lDlT+GY8IbAWJ+CUrMlTpT0Bh2fBzvztrAD/gjImFGKtqHcCuBO8q2diVdOvPmgDdjQRMyyIF8Gm
hvGR5OWnQyLO2ResuKxb9/utpKlHD5fsqcLvVLepSTzne8bYuFPCashkRN5QSh/v6+CnqqZaCFEN
LYow9aGSRL1vYulGKbxMio9ExCyIvcPYmo+f7AFZK/1Wuxk+u4pSTrbcHrqrCB7igQlvbVxTl4aS
/wZhWUEve2i1LujfnDQmy+O1vOJox+ZtSpZmTeEi9gscKgx5icoOAhWMOIoEBwe8XTzPrmWyfUUj
exPl+N34VQ4M6b7PTW8qhRATeKqf9oGZjERCiAf9kS2zxjewB6ZHpRI+Ekwa7NrrGeMQoh9Ty837
v4oPgdUsYxDMmHi7lH/1Se9a3AvmzX1rWTiHjfjL55XKQAUkSHb3PQoj7+XXsvEoJ85Bpc4Zn//Z
RRTFbD5yS341RQ7jX4WK6GnnTdX7m3587Ebs9VCutfFTrEEfs240ErEbebHsKTehvu+sPp9YHZZ/
6+u6egv3Ksm+Cn7xN+x/cGJvGh62Epenrdg8B/M9gq7iyZhITfH1ra6ikL6v4A0FPxhyx5enCL3b
wwpXxnY2TZ8t8vc8IKIYQ9hAcbS3L3StZ1We6xApbs3b8jThOq4C0apb1Ztz3lwG3RwFFmqnLpwr
HjvWLYnEws4XUht6A0Z9QVTcEJg45n/f1UX+eP8So1Fi0p9n/pMB7pi3ngC9bcDqH7LMmPFxbmhI
BDsdaW0wsxoS5Pv57ZNPB1gYdEZxlx3SMk1PwR77feLW6uEvOA5NOK6amJp0Hi7egG+nb3tY7TU/
9kDZjS9zN6lxlpOMz5FVrImU1gM8v4jaY40Yyeci2omxTqJw+HZWLG1YUTFtj8Hiq/5Yqc2OpIk/
sQmfmBtVRZJRyoc7PjzT8JKFQVhGm0BTr9FBEY5jdTbNmwMN5tmv4L20nhDgQybRGOFwP72JGW70
lUay2Ayp8fQhAP7wRTWxi2eSIHoXk2PD4sRcyXI8OIyCNl2kDl+MSMiNXzehbvr1yc9KWbWUhBqB
2VACpYYVGOxsOgJ2kFOFHivzs6kPfZQRI2aCyhLPdawA6/zxsh1he+krAJ+NI+szIR7zmbm3iHf+
IRlLxMyZ/x65Uop1aaVhW/RejgnsQpmQhjqkLz0Eflb5DiBcmo05ZhWATB0G5HYap5zVNpsUnjcs
O9csNR02WkuiwX09WaAq7gWuNnqYBkMlKbpA+QOnRFfiOc4eznjG6RCAddVod/ncOkJJQRglYGvU
9BKkxEuGxHIbhHS3vZznXKWwjhQdTS5Es1CATkwhGFLLn7kcZKFHHVRGueZJEZ015cuKNKWjAsua
ney8kCF811NmwD2NynN+pgwzvWY04r16G56H3dfh1rapFj0kEY+dzbNgERh+Xlli+GWcLVZEyDaz
ICGKNwHqOz4Y7Pn6Fabn6DbxAbQBD3ahXl2tvnW/SArGZZFsHYduzV1qMuT2Ad+NhmF9CzyQo3ow
EjCFNF4NqqMQjIhnaDhjyromcu3V5A2bJ/K7DBPMNWCvFDNKwGAkQmjgHw2vVG5aJID9W12cOjnO
JCylGQDbNtzYCexsYlyp44doD5n4ARFSpJt0dMEosNlTnSYur0cIm6SGUaPrkffEhq7nW+lLLK6Q
T9kL0iCpaKalqUvcN1mDNthB+yZWOmrWzcV/GjEPf8qQ7JKRJS58azWSLDRZhbPh4cmNz95pCybk
SaR5F7xPnsLUiQs+Eu4UyG/42aZA8yMPEwiC0tl4oS4l8RDBRhPhqkEfKw5nnFV/hdI4OtF7kEm5
Vzp/82/qKHUSJu2cT9QAl97qYNAsQ5+p8hy3CtXJYdMcDagYWijPvsf6OK0+dQR+/FgtPNysn2vm
GxWDMPywVULiBmkGf/hIKTbvrPtnUooObEWHoWqHDTTo8dfs1TrV92L+VUKI2ow6qp6i74WQZ1jz
EazchfynwhB+nCbAW8S4K8TjZ6AAaGfigPR9mI5QBa2e6KmDX0V1kSPUDG0ojSFcNFtK13t4EBZY
4phhD/18klFM0PwhnX8QKZ5CGB8VY2jOzeR9QMy/lnxFpZUpsujyS2cgJcE6mndYzuizoSHY0Smq
DI4yb4mkhTxScU2nE1qhej5LlaVB1mYjn0eKfksiv5PBA+98PBCH9K9uZJ4YsurKpIzD868FvF1X
SLINeK0FCvDgNxqa0PU0TrwJlFve6HcZ42ZPYivLWsLRBEa63F9ODMxgwcwOgKitMsGZN4YNOgzJ
48YLvgdvenIEtoKjz5/N3HO5AK+TQTeqsHXsMBp6AYhG+Wj26z+ufdlJ+JLuf0CUoKGeLMPKo4L+
Rm9nLlI13DhiFWNADPNo6zH8lV5aDcxGCaBA+bwVi7ZLe7E/lTb1jgwxYpLirrEQ5lJ30qEPOwaq
ymh3wup9eT2P0wDVYas6g74TFoccwJFzD4HQ2FoMCWEaQD416O5DNGMok+D2D7FJ5xJxfglsX+rJ
Ibi2+kVlZoHbdOIiqLBlCaj45x4RKlwvRrh6Wh8ihMPNYfK9CnzEwsOcnQEalHvHvpmZURaQrh75
VTeTnk7XsrhbF6H2lLIjcZ51uBdxqlNSswIsjfj8JRLtlG44QwQDslN19Rms5G5UE8faf9ktLaJ7
/Ec4nIOmje1kqd8OkhJi1z8cMevMH+7X5CjIBJaDWpkkNp8Jbyv+I0hfsdedbeTKUcV84DbWMEJW
WG1HJfUnp+eHQep6ncdVR5uqKCNFVLCrIWWKB1TiDYWPWvbwveF3WwENIzJqj9gIbERUmX7bCIlv
VjwyNOmvVBVpsQqDvYGvSLoFjhjx4jyO1ViJUAF9TAEwmawwObHY9tdU+dzXDDT1JvF7VstD/7yX
bNo9W5D7dcwOW6VQkP42iC+FMDAhrePBa7qd5wpD/Ny2jZDVtXUfxbgTmN9bQhr2ps3Go2rdnZtr
5PdlmDcYvuP3di313cg63F9bxuCo033CES5vEi5GnVWdRAqZVxGlCP9aB49P/JsYHaW3nOis1Ua4
tUNKHmc0cn5+tuRUddt/AxjjJ0GEkJjadnr+TGosgfX0D2L/NZ2uQj1hqExzRR+zhyT3Jr5NlMcd
Mu61v8RLkFOv6CO+Az/j1cFEGnmYewYhCsNae29fNwamwy9PP5FPOolXMkVJfe0KobdoqS+mcHHB
6lxmckfqwd8wUWwueFCjKX+zuUmoM5QWEti3p7NlS4S/QEiJgdtUkk3ksJ/xrmKXNZzOyUnXP68I
F93qLQ+foprYA9xpYBGdeXWS3rQBWIC2iyxRDdrXA0WaazEc4eu5CKE7RRsvFSz/L1j38RaOC4M0
DtWrUpuGSrsbDiRpfPNxvhK1IMJPSf58Tu/Y3pZumCwOSVVeEpCz+/n1A4RqMZ55pOlMrPGNuPfn
kOziJ7Rn7IT/FXypIV+NepFrplX5lJKnOU2SpPHAe6TAtj627RTOwm30a7Xi5RnXOeuiwq9pfxN8
MXZl/NujDMAlLXAVpUMZUwXhwAssreF+VfkZya+T0HBco1cWBToSf0IEbkg3eqU/q/rSH8/+sIFF
7uJDKZAEiaPZCGgFSKeRwAg1/Xvy/vLwRfrRPOECOm0YinClpQQPkROq3Woc4BGp/EvLjFq3KPy+
R889jrxSOboYqsPPfSnNPeWbXxcvqomyaftpU7EdHp2llCqQVWwzR4wnE0Za4NCiovrstUblTUqP
nIpuW6+wiG/UW2TOcS5LAm6A6JzAqlC6Ufx0YsPA+CpA4zsetS5eAq6eTl9Skb9ZBv87sA7tLFBf
iA07CppdpA9ptmBKaJumz88QjwZOBRI507PRUIIzd40DZQMeFiMGxY4LE5RvAEvMq9YqNLmn3P0v
xDWarnSX8JGlUN4e7S/wCDPKnLuxfDacVCcJrTNWReixqvaIEHgzkpzF4KgLbYYLSAAgJ4lKPngR
+Ik1w5LgDUqJt1fsEwSvdEvKlortYFdqnJtpZ1hQ+/A5yW89MUibD8nZEitcWKJIAmjMlXrDu3dd
h2o+ifS37TexrZQZaNuBhwQ50s3inpmoCesN5UnkNwsAXhmQ75fM+fFd9nz9AWKQzBreFn4lVGbu
7muoD8rq6AZHYSSnZBfGv+13t5DbtO89jlws7FogHOc5eOIZYAWWN9g9V/Q/aiw/bRdc93LzjAOG
Vm3pnrabbxjqbiIXaomfy2rc+3JEiZlvy1G9v3ztLLroiaKWMUbRJh4IdTRM4MMyU/SLstEwwsIO
mgM9KtMRgi/ngF6rmpVXn5TnE52IAWu579hmK7CInie4K38TiPOyAFnM2luuOUWBwhGcEXhNRgnn
1x+s/ECXxt2AVAftFGWgMHiNJD5nQIzbsAhsG78aI+cBpSnpoS+R2zAKW9MOs/9xTvmPu93KZ6yg
nJaVDViw9nmREplWPfEPx9ikz2Kmye0AhQ9+RbtYj4y6AxZhsmD1NwKKasHkAOpceo+QQnl0k/WC
IqcUrciP3qrfNcfQPFfkuRGJtJOZun7LaC83voU0emkjVMfTYh3kGfI6iIJyp1+9r+v9+9J3+y0x
ZwdeenQWxNCoqMNw3PaDJOfu9j6HZwU8kgzisoiYrjlfPXqKNEeK9Jou2YehaRM7m58NsxcOPwMB
CIGGU7e59Uefb0J2dqUZxYlnfL4oLsIxn8C4GAEBiHW1rUnMvFCbcwDQnYVVodlXijX8zm+M4Rc4
TFwcvN1hSrVj1uAc2WZDPSYJGRefkjd8GV4+q3OlpGAmrJu1nQaK2It7mK3ySEPDKvfDaTRPWZL/
6wtBynmmq6kLRNuO76poUTMd/1Rp7/ClclgwU8IGEARCcYkp/zPbBV5Y6kRxWw8sbWkrN1Y3xfJa
PD4vDjhRPXkO3aNfM6UVGplcHZbN3mUD+FRKt+rOjtsUpQJpCTqJKGRPAVywb7eZJ2NOLDMYmKUx
HFldRPqIYT+ohh9v97EBHAvrMNAkYk5NzEZFUbeqL3miC0kNOx9gQ5IJkdqAjLpe3AVMBdrVp1tr
WgMe7u+wIsMcsnZEtTDk7jd3LJVum4IkZKKK5KubQSR3CY27pDJAJ2IJwqMHfoNICjZqhFdiR2uc
BjODFi2IBysgxmMsl/zKdQblAx5OaEpg6EHsCZF/Oy4IkvIZlb4QQdAj2br0uob3N0lek9zWsFd3
I5XL2mQkVSp1aoHWhWTLV6jr4T6VlAJFQsPsNnn9gFH3M46rvH+OXNRcIgtB8Z9iMkUTxyPx+J1g
nxVI0OGaCwraKkW0lC1TBTgHDZYycmLJEFBUVdsDEuVQagx1KSBdKW0pxc7Gs4iP7v7dxmHQfs42
v5lDFrQieo6tG8Z2okR1B4Sft9O3H3a/PgZ5j5pwLt2entv0TATwE/7pu4PNpj2dgq/vUcWNPAXR
bpmwzUBJRQrPMaatMsmbAhenc3sUKEH3/LwBiNEblT3JxYAalWdjXWU6avwvvFp4DhYM5XQ4UpG0
wh0C4J0sZXFTKq34Scy7miCX9auYXA3d400k2Xu6dv35CrZ+7MV1zoc1ht0gZgg8NuNFeKhPJSs3
U8pq7+cYyeV3FSQ4sq9Or19Zxaw2YKsmqyQUUgQng21GhN+TScClkg+1ol89DEEmhamcKiZRFOt4
UOeq2apWYGdBIyL49UkyPXNUqGiA/bCmKrhixFSVTTi50nDTT4Sxx8/vswX7UIyhQ3Wdt0307s1v
j2vj3pJqfc/VvfyY8CvA1UV/lHAq+WGNUf8UTUuTL/f8xMQozmMtCC2VRCII0GR3a3P2BYaO+wX7
1r5qtsGTHfWbnDhcmrARqWGJ0xeubzPfu6y/oJkw00juEz2US3zxaTNVL3nqIJDzbaLvJJoSkcUv
yR4zvfelAS+jWriVNHWHP+yllUmQznmGGp9lUsZVmPco6cDR5hzy13GJVyGl9ItWQ+F3+svIPOwv
TZUSFygWRZX5j3w2Nj+8KGk2iclBfYlnIquaGLtrIgZ3gkQZYQZ4R0j/mGKjTQvhQy4diETR4rru
1i7vVjoXS31CO5PY5hLeRXMNEoh1we6cA3PO0KO1RPRGpGhD+kKguzd1Ig5s47asaMzI7Z4OtNNs
lODdn4oCWxmRiA4aSIQpKuxJM8xIUc0WIc0WDoepOgoxx6BW6mdnXPd4iCl9aCyUcV+u2C7Z+tG+
nnFZ03g1UG3UHosWMMxCZE5SKjs8sJfx1DIUjCh+2b/Te+ReKbyIRPDKOD+bugsteE9O67OStWzb
evnGSlwnaK7LDW2nUv4x76rDahSGhaUiWbr5OC65kEQNpFZF52qmoE02lE4ruzgTx/FXgAFtAVJV
4bNBScKlZWmtPEOBjWKmYnq6DgVjug6v7ezHlhL+OHI2FHsGwOk8bjUUydBE5tIQNgm3EHf5mh0v
NF1hZMU7atzbfN6E7XEKMmdc4OzhTq7iRIk3CMIMo/TiCBnlWCTgjTIs4jW48WefI2G0ttX+pTIS
x396WWRZEm055nXAKp/NlbbuWPi6Qxyb44vTGDKld03BTJZl9lOdqrifscEj2a/8cEig+Yvp4lqI
7uP4pWdGM7iF2JV5OkOt8uaPR3u8CB2f5Gz+P05EU6vnzDWNFvKVeIbaC+YVPbA3/NLDwBYWxl9f
IB2Buzlav5pwdjATq/apaZPrqUAmo2lOWRrPuVpdFBD0wYNUxKtCDwYGaaPjbq/Ah5V2qhFZaOF3
TDT9wXNuko9xSEr5pYfIXKCdMlNWvYkDaeJhu24+RONsWPSTNq6I1yjya8kQiu/UYghLbpuOeR3A
VnK5/z7juBiqtXDiJ93a4oftY7U8SeMR/vf8Mn/kemLnN5OeQXS2ps4l5FQnSbJgdW8BipazRlwf
eepMXsPOR5/KnvqFidLEILvHuCPCE7wY4YFj4X2C1df6hcgJrc7HXsxtVHgPKPzwOCCMJ1+NLO3Y
K80cD0uKTrJtKcUDOe2E/9TzZ1APopOBj+hpBQZ7pH6xo3AYBnCNi2zrll54XPJ5lfJFM4z4QAc/
pRqkhlx/m20gHMXycuyb369khOh4YzIgnYbIojyVYdk7iETQXw46f90Cb30RAi0EByTG/eup/D1i
3ab1VdIkjdLZplHCgJoP/k9G7FeDcsZ+IwwMZHGs6WtIgpBMVxfQ6pjKTEJ/u2CH7yg8NirMVe1D
GqcMZrlMGDK3vXKmgn/MlU+cRCzo3vfVFD+Bg9UwgGG2RZoTaLi0thFoNpFfTVhoAz4SAm1TmY6u
Zr3r5m1tukBvSQshmN0Mt+605qEW/qhs30l53N/lTPjAfcz6j2/PT+bDTclALzZTk3C44Ad2rGf2
V/faCoVBNY6X7FSxjulw+23grKUquvWAeI6gtrYwoqjHZurtwWwu1uURIUDJSYGpXlVr3BjiZvSs
ZXitG2br3nprm4HRbHWcRyStPjzW2thiwPrQNeRVgikDTeiMw9eCcis/6x78JMCiItBrgmhjhi1Z
teuQLi2A1wY2/16BQIul5wcRqcxVXg8+iW9W8J0QDDF8RyPimL5e2SBhESIRCpdI89TeU7HOkMZT
H5E0YlYJ3XMB2Rkon8HznThmJiP9qQIzgxIjemKIy8AfHXSI+0LM3TjDi+cw48LgVTidHAwqQ6um
iJMpEPMqD9fKLe5lnL5YlADt8aD6KPjGaqBLzvFDPKCd6j5/gXlQ/P6TOpuYmHKOdx3O8CQujTsj
vlmOOY0EmW8I+lM590osdlpF+EfTM7KyLOB7+RNjkVIJ3uWxhqwzwFKt0JQ0j2CypoHEeaohKs+c
HtRoYcPRe800SpCER7fXTQPQvRpg7TxKu18Wen8C9gNUKDIbnivJ1COUQxCHpvq90Db1OZ4Oeubt
ZsQhNV3zd7yHk3kckII48jXUA10adI7W7krsuWMyNH0cQfJZGk4YLCao5s7FgnEOdF/G2tJ+zhtW
p2J/0yq4NfkVRdg+PcKniLMB58GbeFaVpkZluUUBkxCADmm4YlNpNzARgqYXubPyRIPxpW5ifCcD
PXXW5l3cpKWKAs7PUOdy1vJDLiwIcg/qWYxv+rbX9pbgDXMF2oXeofT63tnR6NwFB4mIMjBnZf8B
SR2z1p4WVoSaaak3JqEMdYOb7oSVFkN/5oMtMkZ5Et6HB+8XXThd8kRSvDZsqBTPHcbMRNPD2IgI
vT/1tC6s+NdTQ7Z872wC9fD/xSDEG6lDbGVSjP6CL/fuPVJiXrrMVpYcYrM3N0LqKZCpMB2C6o2O
WwDXt2CQe+oJJN7dZVXF0hFOy2wh2CUP6yMQSFF19zZg2U/bByJ8uO1ic4YXJ/OJzaZh2Zk0HCGV
DadS6eaC765b6JPx7UBfFkHdCPZH477xhG7Y2JIlGA41QYm3GNYn/8KCO1lHkuMNQvGUX4OpQ0KI
8UzI/4A1oy8jXMyFh/07Sd3hOJTi0wZlX1wjGl7Yr/Zd3VAwGHjtBN430CAtSxa1MQyDH5DI+wpH
k6LzbmYDIJf4a0QHMguVqXUpVPck7p1tnDtajHWc0MxADp3sRa04002FNITVB6iDnkP5WDz/pssw
28aqHIGzURI0wulAoztXRV7j+Kusng06b8odNNYxyF7ToqtFZM/o0M9BxvWscIlCS2ZAw71O6Jtd
WvhJI+o429+nkOeNSbdnCuAPNC2uXLvwEF35b1Yc1kwljaeednX/BoGOK5P5kD7kIoo1+lbF2/8x
ZDz0UEnxQMSr4o90VDVoK6UW27jKcIHoZ0rEDPledyYZe7vLhldikodCJscBLujFNduTzT7h0vAK
1rgtBXV/4W5RaC/04znsZYplPI5BUSL6C4DQApVZyKovIuT82oQAqHeSvg7MKHhT5ne3DMEqV8CC
+OOjOmNiitp8wtUim5MVp+X1OKM5zRGffkfE/pkXZnBiazcY8eZjnz57imK+wuFqAriNCEvvRoef
SeNE2aOwQEuiz0ig2WJ21ECuu7yfYFPhT6rLCount4bZsChgCW24LXIABFth1AtHKMo1h0kMUdDW
9hGd+wYso0NhYlcx8BjY/ydJK/GBHYF9E6smloLMeczPaFok6OktUPR86zf3F17IiNOGmEo11PNJ
YG5p8CSehmZgmUGcSLOnMup3f0ntzkiG+J2M1xi3tJdU5VMix+NfuoQCq2qo0QIyVy5yn1W3Rl5D
+/UWP/OpRrRK3e6wakHIKli9gZznV/3l2WIkSYb4epAeHNJmtYe5xqnJNhvvFEsDj5IhdMEGFjel
bY+mjyPvUca9MUrdHuzYT4GYp4KJXSlhIUOzN3TP+0VCI/LreNZVhWBW1kXb7ZSJZoOLaXs1DYbg
MY7dvZ9njRdekuF1bs3bb9jxQ5ZIEuv0NkY1a3aVJe9WgMtRiFhasnyCiJHEcsf0lpzgzxs8CiN5
vmLTKUPAYY+jIXvw+KCV8ELHaRVYSVqesIlsT/27ar9hApej7pXwlddXx2LEeFxwgcqcTYJU/0sR
diqju6SqgHJcfDCtmd5giyPMr51rQSSwFPQRF8krO8foszVunuPYnSxRYzYyHqlmAT01ghzVqK78
JbsQMErWwoMlsmSZQAqYrAEknSppKOqB0M7Qe0naLc4GSekmbb6CEdhfb/LfIn706z9R0svvHihP
ug3uziL3Ot5NQaVDUtmlcgY+jHIfU1Q+n8dQhnsRLlVjPaPTeP4pds0xxPEOGC2nqyzBpRzaoOAv
HYrfIiYbGqgKK32E0yJTJFQIgX8dphdWWH665JuNiVI3+T3wo45GzO1q9j6St9f3BQFNGm0H5Al8
ZIFM/1EILH1t5JiSPBWu6N+7yIp2IkYbb4agke1oJTGAqZUTYdA9YjGLwhOdFeuI7uVsRxPcnbBd
m02U4pR1Kg6cs0J9NC3LRBu6s4g0602rtqH2donqEkBKE2L1lqkSKfS8d/4XtXrhsJNgqqcJ1akS
rGMd7+sbEzyxNwlRI+iMxORsrYCKyv0V3xGv/CdzFcG05tiWUbaMk73wniNslnJlkE+M9iv5aD+c
cZXO+NgEdR9zxMU2W6dpujDIX4EtmrO/N1snI1nf3FpWZGrd5jq7tVwjU8Eyg5VO35VQXCmqtOg+
NPuM6Iban8mgOnVWNn2hEJOh7uayjEb6znEi3wUjpYnPbmAJDQWGpnb21MmGLIg66FkppaikjiOP
8Ix9SyHW1gxlUnhHDD9pOe+0W3WvlTDBUZLl3qENqqJat3qvAO0v4Jhy0ejdL2EblHHJFzr2Su0v
8wiStOmRr6Vy2R4gR4aKVgXR868E+y+VBlx/TrZiwxugcSehogbHHMCVLhNu0zP9kEfjXv0N7JVT
mSpgtA22nB/liTtnVFuZ1iyT8i0rEUK8+QEm+8kT8E4tPzn5D4eniD4al1ra0X7VS3Y1Rig/cyr6
7cNDNXrGXSrD1vZ7hYU0k+O8GgXAM85hz31KlG4VgpProOWoTqTZj4VCXMuv8RucE+mAfqEkcppc
2EtJzj4FevcoM4rrxEI95tKj48V+5dJiL7J4gIlF1SPV+vvB7IbuMke5RHXvKVcWm4F/lQ+0cANm
rXxKRf4dIQKeGBK9XhiOn51/MTYKyqf4tkpyNG6LTG7UymUW96myQg7OWl2/lMTHnAp9Hw+S6CXW
ZXLLBKZpWTtuO0aH5PfhppMKlWKnV/bqO4N/uDKmw5yV0LWfg7LAvjGMv9aWrVtQvCjUTPJzCiIW
QBGGv83Kr4L4XsHW7F1MeEGZoRLahE8o4JiG9+aEKml9Sp8ttX5txFLD4zkYY85uu5+yxDDsCP/6
H88jg/6bsxlocwq1z9jq/jJ7TKf6wvnrm1sbzTk0MUuXjomJg6j6TamIchPZLsF5i/NdkLuC0zuC
Ur4LoIGn86FJw5GnGgFVQMukVDsmLEgppItJPkMyZevQSbaNzs6CfKmetneSRb72K7DWmNFSE3c4
nmxCjLDWDf2WNUkwXY1h+7nd6RR4znCUT1YWaDgvtfJGdsrb0EnFKtdtpcE62nzq8+RuhY6QmgHn
NsIY61YqQ6aZaaL/YWMNVU3CnBKtB2bSFN5BdNopmlRhsJxXH/OdBF212+brJUeNHhEISkyn+R7T
+1AYzfVPPgAyI9wO4V5Gw3LZkYGWKGpBr3OPK9Nu+GnTVaYJIEdgW1AXJgTHMpdnQ9PX9K8Zk6Zb
TNH6ZIlGJ4eM/IRvQAps6Um45VFmEl4cVNvmr0tmPbFlqOHeFyrRGDAvffThP0nwCdWRbicZOKPV
na+jfDZ+qmsMchn8LTV1xWtqYHKt7+TKElcVNt+Hf8Ej3MKBjEdENvrACk8BAdPBJ9saDUBKqgTw
ws9mngsRWYRxziFrJIQPmV7vbpOtF222n2wLO2L1ZLzqXjBIOUD/FX3xMX+qKH5F8RiX9w1f/8jO
VZq7DiAOt8y4uPCcbbm7WKEivO9z0OOfripIMC+MSREAHHPirCoK2QbS3s2Gd+Kazy/CJl+8NrE7
5xy5D6x8gabbe1RK6J/MxS1HPf0e8Azv/QLimqxLemDzzpvd/32RuEYN2qsZgKuAbrSRUO8kh8dI
8NEb7C0ND/BGPwBI1nDkMVVJAu3hfceEjxmDdhmN9hcnE5QkAqhG70LcK78Z1BI0yd2sk33fqNpc
+EnXKoEr/1ymMpTxjnIgEWcuKGpkUK+MQ0nNYgDYJwQweAxcVLlXsCz+5qx+dKBksfuoMSFReG2c
IsBEfj96T9eU0rheGq/swTCfZhr2j7D08cvWCVcNbmdUkY8tNojrBgDNbUCAwVrStLshPSkJIc1L
6ziw6tktXqCNXhULFFiVHE6DWQIe3S3WzH8Cmck+GLMoRVwFY/+bqvZJH7/4dl6xqyxY8l8SN8hn
196YsaCqqB+Z7TafwqcRC+oAlD/dOfmqH64Q57cQmDEu3PVJtwXLYzWZzrSmC4MZhBGBDRj19+Vf
Xa1FiheyXnjRWQvxKZaa5HmCrKoqFYsuUMff88MVxSOBqhKKA+FQsy7c87WwxXc/3SoAk4cVz2Sg
psrDJf86m4q/TKxf5Rcqe/mC1DgU4MyljGJhMX3HEeb3BT7KPnBYLOaEraKzNopl870Jd/3Gr9yU
9lhe2lPYRpr5QRrpVXKBw+iDtIkCuBsy/463KIY1Pz8wdI68yR+HxDAB+n7kIGeoJIaHmvmb3Kqt
pnyW2PKoMeZIen8wQfEdiniqDuUcLlSZMqEREO2rEPgTU+G4iNxQ70BSPy7wvLvl/MiFr9FQy9zJ
FN71YX/LKPnPvijNp4W9d86SEMf3qfZPdjExxrg4aCWaLUfnCDRCOBd5pNN0cYOhjP0g4DCf0PM0
qJkPH4j4n+iSRW8h4p/NUoHUvQiwI6Rqyc2MfvUh0Qn9SpkVhMnvKre0ZKLZLMcguHDk3rj15oTo
1prDeFbRg6g4+8bsjrdA8rvwFS0foNaUFfCtC7yEeD6A2CBI98/68kIY/ttEzhf5q8rChHl5+ozi
vrucZDHnddmWNGp9GMFbA7PJZHaUY8fCxsXjjqBPbGekbREz3N3Nz5xhzzzuZxJnAx3SQ5kwYOqf
Nx6wFfxU71zc8OurEkJmPdueP2AhyPZgN2veO9If7EM7OIwpav9D39zYYPm4Cc8qN/+ZRJXsgP9I
5BS/BM0XRmzYAD5k1Jtq8A+LQjiAfDpQnnKZSRS1tq4+LEHXg/2KnlNlJ9tsVjMA4hQ+mXpFgrvn
Q2mXA0b5vBh4RDQz33iIkZ+hW0l7wrFD2jAr70gFzQq8POOQBXWFWKaVaAK8bETYPaOZE0Uq/yOb
t0Y8IDIDJzpEPY+sNv1wfQ8vnM7xURVIfQvhSMDutRsN0azBwM3pvYbrx/ZqvCJyES4oGi1/1bPe
qOSFsdDODo+FSjstjOB3dcQhcE0sCyG0IapD0s+JDTvXdbdoij3WEI3/xATdM//8k3Bk5KVBTQgr
OfVmLnvNu2zbEKNLIN+uJG3LUhBIIXbiuBd1kUtKjUra9UQrYEu9ur2XNgjqOc4i4ziqeZyUy0jg
JRJLAby9aChQWL91DxcUVv6GAihiY6Fx1ykigNztl3HmEXSWEVnF45kFDCAgmgUm4Xkti+RdLvSk
JdPZoygcPf7TWmLLgiQnQ4OTRfBkFxYchc/hDzLuNnBoQPvGGC/Jol/pwIzPXeGWEuxet2TKD3b1
eh9INwC+lX1x/wWIt+ED5aaFRl0VF+s3n/RHgdfG+Eaw0jv035kDSAQfmA4vKp3lpiWkrUcdXYs3
oTnbt87ucxCUyJLPARfkRaGOs13LzSt7zHrCVHSyJbZEwAYNcu7YpxzyJ5dCRucnDof/IQSm04iF
ry8ykW6wxDA0FGc34ePQXwx8gNaaXjtWyst+VU0uCVmUOacT6TbJGMCTZR3Y23r1GqIoozxUa555
78Yu5vY+RY7GYKS/TNDiPh9p7NSUZNjhUFbF4w0s1ziCdbb6Iad4CtZT2RzfaX8mh235FUwu3km0
ECwH3jOLHrWoGtAUCej3hAalksqAah86/tyQPLe/t/fmh8DR5FlSA7FK8HSlXwpO+dDG2AyzFloZ
AtM6isSYMOnchJdDh66l9P4PcobkaxcH0A/8jgh9hRBczQ80MvM7aSpjrvaKU5dxaGOrrOj/dhkL
EUgsgcLnbHqHxvykV+/yT0ejs7K36ep8TGSFnByFSYpZL4O3SWymWlhheMmcy9PnD22j8IiiWPiQ
ixtBQhSHXW6ecbqCYWnf62WhekHDwQeujyjniPITLEo4P8b2lPTwl7bAasfimH1IPei3JXJLGS3w
WY8v7cTTiRb7SwzW6MGuAM9SSXEE/wWFLflWrctD2yQHy1N3fStK09pigSefpmYzcjE9ipUU0+hZ
65IvE1YZu5Ir2zAXZxhBgQhJ/m4FTo3MpZBoBQ6UaCt3nnoBaVUIXTMqfxLdajSRpbE7RRaPiMZ4
c8tMkldqfwVRaeLzOiiVk97YdqiHm2tRlx1+4EcctWvuRDRwhcXp270A0VLEsMwJYCMsX2QwhzMD
/KG2AP4fkP+soqVJnaZnf6aRxQfAVKfJjPXekGQpILHECuiBbMU9TXqhl8mm+ENBlfchmj7bpAfB
Gj9j6uFDf4V/7kXycMH4LSyGXSvymwIb8BKVUebOdPyz1MrJLbf8dIxEJ/o8Jc1WVC3E1NyC1K1w
ghrf5UCjO7w6kyX+r7L4QSzP0jgKJ7dkpSqOmU4UNuCP0B4um2Ng8x2JVrz+4e64Ye5HtjPBQsZk
nc5HmksiXfTa0F3Bp3CzCPGU1yev6KLNwYHQk20MhbFs9CmTbOXEAE2Z0mzvcDRvPHn69VYExKQT
4Iy7FS8aa1Dfab4zemDZiGO/Efbm/I0dukBSshFbyjTh2V7JN9ftE+QPvXVo2K2nAPjnYOPlr8SD
WV3cNMj61ao7uaJllfMSON3MJyuuK/MdRKHjjnW1bV1egBf4tHSlcNI2L0SGURIDwkoTylP9SErE
n2gxrLVBJWgletf9Q5RWAzJV1J33oWssa1uIvIQDTBYgxpard+4VBsgAetpEclhtC7AC3hXpMMBr
kgwulNwq9Sg8/28MpH+egPpTLBlYkHcPFxsnkKyQ3KDMOmyQnDWX55xe0017eFCZIwRfBde1aGAI
VoOXVYcFWzLRvgCxdzCuU6amqUC52BgckkLdmfGQ1262EAaz+5Gmx854agOKra4qmWPrBTsk3Cxd
Evo6XLUpCCn4pEYa0Ng65AbCetNGluYx7kwMBhiDuGG85tVPU5REAkLRVETV4yFrBTRKqwrUk1xk
jtliV8HELBW8zBEsa6rvoyQI1rfEcsoinfL6VCpQSxUObxjgOCbDGN32cA7y3Tewxy9HuYXrYkdf
VWsHN73hdPEzCILpJ+VpiUUCOGCe1Ri30ISL33+oqN+vLzXBzEfIwa3Z2034RAlV4v9RZBddWBqm
ET9NVuIvfQYeH401Fa0CYYJtkyB3sLr2RQzQp/by7g2AuXffcUNwysyvqnaoxbGdXZtRxsJMQWLe
7zUk694tWu5BXS/a/dXS0uZG90HpRCriT7Cqq0c6Bd26MAv1IEyfnV5zkjUjlyH/0ByG018ktJ5f
GxAU56MinSMTpP9zTwJc4ZAu1RCC/BYcPr1WYRB90y2XbhipbVBTVBNv7VRxvHah5TuSnWdv3xs6
QL7wkbTkx7Bz5YDXs/flhENN1639WAKNr3tD8talKoUaYJiStO/Xodaz5g79/r6xqXeqbANO/edZ
4J7BczUSqjx/ckF6oRMLqLh2p9JpyE6ql0/JsGsxu36Vct+rKPyT6mSc2kmqHwXRm1Nc5EgiYu/R
Zn5qzo7fZy6KBn3v7QsuJQ6YzSJyl8TMwhClPCxDk1peKEEHmXzXze60pLpussO8vg2oITw2hx7X
mnzTnXGSJgUDKVb6Yw/UQU8KiMldvz44bpDzhSmyLLDrL6qRIbDpS34eGYkUtDiuMh9TCVE65DZe
UU3H+j+Ae87YxVzStLoBtrIs0S8Vi+tPzC8LeqRoH+JR6jT7hUOIi8jh8fqYAXNuy1AjChPx3nkK
eCERuOnBvV6Q9lKrg5GEFD6hzftc7SgEWpsZ5PIyLdGKjDbim95nY7azHZMQKDtlCMi3+ojQ/mIq
pJ1s5FVTMgfl+k46x0NdgzLQ6MVVrkGM7wthM/4L+GjJhZbspB2TcH+nQZXA3XdyVxsmCF/JG5gl
UYDedMQ6RqVwbzePYMpNRQpDP0E5u7tlANrFXnbklfLREpSnQgkqFAPjdYrM44OvYA2qEONGo945
lTivyDbzOIca2HnVULIqbDMnV2XvJhz78RDmIi9z0kJwrtE7A0HcfWVLrf62ue6/jlS88DaUoiAI
GH4UPObVmFJ4BS2dx9izKCzl8khuMpLWHpKsC2LQCK/sFvMI6rnUaQUwXrv42KaHpcpVUee7RFbH
5ob5IEb2Xlh17genr00myS+0pIjQ7HUHIvRnoZ4GIreFp/hGRqerjTShMoMJsWFfV1Ixjl0vmUXb
dNMbLTg3wUULX0zI16ZYqDA7MdJgG8a5KlBCGd8hMV0MQaAUmkCVpVsDjRd2kcT3lbcfkUg+nNQl
mrpz+JYwb4T6CjBv0Ns3nQcqSx+vrwySMQlH1Y/lpQoYL7PsbrM1m5w+z7pOCZbXpfb0y9qS1tQ4
IVl0sR1KN8BC9TgnV3Ye/Z5AsqnQXXSRI8Yue9lbMkCcVHrmOO8X6lP/7kRAlqYRMeHHHGYg367Y
N0m1mrMSG0KpCNXZQYMtwLs7vr9HbakpWylz04QaICOn6gUtSi4M8td75D2EJe6e5aB0cZpa+bq2
2Fnl0fifZLjt4VHcVA3OhNC/iKUjGUA9hwEtRztiVqOqeIxBVBA2RucaXtPuAsilXt+FtRcXu5vN
qRsPSc7unUTjPH/r0nLCMpmrhsRRVn+1Pd/UiAEfCbTJ2iOdNkgXjxGzRxZ8wKnn9Bl4Xwp0yD/N
yPw89zdwfd/66vRIkCAtsWMh+frjlj4ep/FbSzyHe8NGirCLb2vKyzVjrWbl52YfvoQvCPgz+0ic
OLQR14w0Iud6GecNwgS8x/oYOppaiOGM8vORsqr3qHdcAX5XWHwPjOCVQ89aLYsY1vKjxZj828Ew
DRpkTPsB6Td5ULL7n+OKnL7iaqGZtRKULX/O2RlybJUa1BxUcoh0gAQNq+1Gp3gg+rGHeG8Pfpu0
oNmDEnQKZ0VQCxnTO8/EN7WNWv4KhwXgmUxyD3qJW3EZWjMl0cj82baOeAHruuM1Qm6i+k/SYZCc
55Nrkqwz2vcwl7LCWJbIVsh/RJFCDP8FRcaGny/GAdxWnHK5qo4w90VzYzt8y/auV5Dpp50TdZsc
qYQQuNK9qjr4QxzWNN4G/Ie334nextzRMlMsxy9o+jBZ26kcXzyp3RqGkP44FBgw4sUtFLNxOP42
2gemUoDUt9ozBKSOy1w+uJPnjWCRRLBbLx9iJPRo62d724S7+JX4c/HBVnncQ2G6bgk5KYngeHXG
O8tLhupCONTtf7w9MQS+REBmx1WZvtxYM1kCT72ucTEq8XTZe0fMz8VoKveOhuatgTm4h2VQkyvo
6nazQTay7UX7rkJlXEfg6S+zR9wyspaRds124VCli85M+j1DhWYPvOalRSwJC0MkyPjeHiXBeAu/
Mg+y1GTJGMLtTHZhISSFtYxc/1OjZFNTMWTUPrEpYApdwzVjt63/Lr5CxIzjkxxWlYdkdVUv/csK
zRhK8RyrsLOGMtoSclKdDmOrPlctBzyKR6HYzaPlXX6wmYJsq/j+hE9G1Ly6S8PJKc8xVQ8qdK5A
y8mfRKqUfJMQi7ROuuE1EV4w4ggNXtR/67Ca0CJ9Xw8+nj5dPHmYEgOVpAwACvcEwGHInpZEQK4Q
X2b9asYI68csuuCBI+MpUGHMWgTV5lB5Xm1NoRoNhhWolYyobq2oi5KER192NA4NogCutWQu77uF
bqyrtrt+OA01yafZ3buqqa34AWP5XW0R/Y9Hst7RouJonf7r8hyj9IJV/tCTMtBA9jvXegoqZRr6
a7uKnmgjV3jccROL6AVH2DO5DHHd5QgSimHEq5L1aDgzSy7ziTv2gAymEHw0yP/D6Wrh/pazBtuf
NiWgnxDdjpn/XefYLhrDxv7tEDbrpxNVM2ljzWV+E3yscr1bsSvPN/eF4Q2+khW4YFSiDpjcBuCS
NUOufFrMOfUeoNjcA19/rPe0j6WhlRfTRh+zvRFoi8Bn1AJBogHX6GwsXjtGlTOPKnWWnFdD/iUu
5DkaVnnTpWVC23ZroCtPuy9niC/RhP/cfSYmj6y3CeD7QspdpyKGOx/dxxXYZWjXUogNJ4ih8nyr
aLmXdi3xhcM3WTaT/j4I87rpjgMJmitYQzXrBspYcZ2HR8BJzWcuC499X+JRmkqJbwG8QEhMc4wH
BEC2vZhCCLoCCulRti+TTbX+/8PmsqHAZAPlt4m0f+vP/sGq1k+O7ekhDDvfS0/8DKTXR3LSt4qi
36KNWzL+PujgZKhhNptMLv9+NkkWap/MNS0O94oylZaxco9q0yphd/7xPZyZee0DwyaKxtCG2ejB
Kv/+DSsp7fjN+4iXi1m7W+p2fq0rVm7yiJLKvyCuItnXdB4GvXbQ0x3c8w65X0LdYk/8swBJFeR/
4pi1zEEO6ojX69ZDIe6qdYvzIwzvIs2dTfM4QIpZsNaI5dlKArH968B6LfWlSvVvPzdzoqIQ9i3n
fFahxcriO2u1qXATtMY3aH0VVv5akM7Kg5voF09091/3BlXkeEH5+jGeEeNWQMDXyDU84QWoxTH4
4IEezyUR/uPd2iS2EkB2Zf2KIpqc01duM18fVBpG7HJ0IUXN+7LtLORGrn4u6Xo6r/tEY5n1R1HS
mV5UJGM3RowpH7CCnuxlQg4dVAOUg1rURCpWCQPIPcrmUzpBtO9Y37N2uLXpwr9GuxKxl/03umEd
oogvQQWs9z6SxDrMOzZ9cJlS+HbTe0z6R2+655PPUp9NnbIup0B0O9O+J4fdx4WjQhoU9yeenmND
eSx9xj7QPAtFynRi1HcXTuoqybQo77Doh8OeAoQu/uUBkvGtzvf+DcI/mHbPyE5ed7nMTHpgws56
2HShyJoZtF0EmgCCeA0rMdMXP9bDqd8Na6K0zq7UnuVCWPrWwt8XfkiVlwNnqXwVvfABK8gZDKfa
c1LcTe3yPfO0DYvcGzQOGbwV/PgtaDgThnQb+sAn5km3AuuJJe6a2h3amtA1JyuxL0h6MAY7JGq4
IeYK/cxlROtIX9Uf4KFLxSisU/C86zo/N7uPdQAFTiuyjbn9/cF1emOuatFPG44MgvFPvHb074IW
h0mcVJ7xlWV3G9qDPn9/nTGM9oUi/5PNwDfS2NhS8aTXHNsW32R/zLzykxfGA1IOQOHr0SYH2oiQ
Fg0BLv2jfndUG95pasHKE+p8F4cC4nm3hRbXygazIHLmtWF3J9WbElaFRW/c7OWN1Lft2TZ15Y2h
D+fwISMYHUl5M+UPH4i7Wp/mHrxcmFGP4N90OkmSHXUrKqtOWcZPQ09cWSdCplB7qt0xnLNZYzJK
IJsc7WKi/A7dEdl6BnS6ngVjyvtaWnrrLd1xnR3FnvrFEmWPWvBsSGl9ybsMnHO4q8mgKlBroYWT
At1QxCbmYV/Jb3boZZtaRcR/P6u5MP6IQfjwDm41XT9eZRoWbYTiDE90CqQ+gF2VT8lE0OTsk7hC
RDk41ysCqAmrNPZDhDtCO1WbFyKCXqO/0euOTVUTixBO8lvSx+gl5R3hwkYOxcn4zpLOhyz6kzEt
9qadqzvNDPAOrR1w29G3E75yEj/NKkhYFXIIyFGz5OpNs7kRDAVEBpaM+YLaJCKcU839JmLHfQbD
ZLjnj7FViffBXmd8UJGfrq3lUNc9zlpafQUHwxLWhfWCgdRXF64+dxeOIp1J1Qn44cNppU7oDgxS
+Syn+tm9vNGJOugvWn/GFtZIz30wXXeBM6Vdw1x6XZZ4SKmJk/dDYNCXPUhoa+KnwKtfoHYf5ca8
toUBZDtIE4qKoEnh/TKOoVyjnyQ9/xMIWoGnWgei694EISY0Lzg1wuE+kCOJWMt8PZp02x3hwDCU
MsRj0ci1sDNlMSuHDDH1qT6nlEK0HzjIO7qSDKx2XuwvMuXS4dw6vwpQCitl0Crv+SyAfGDk4GOM
db+A4w5Al+6GDkUPHeusbRsLFwEsYnPxJ61/XkTbTKxcmshKxFttvyT6UH9ABeJRRgrEOHn50k6Q
d5j2iRwtcuFSKO7l2DJOGzDbUio0+g4qDbPvbbrb/kXbenp+3X3MIc0iVlFMSi4rdHawr6cQzzWU
Jed86kYi0HJICRp2Tx/xB24ZwyYGsF3wQaTl1pV7o1JXbeRNOr2ng5THS2rrwyT5WEGKShzQXZda
CFwWOpAAvYHAwrbFNE3NQH0NoDLO+BDdQxuca3R2iZi7FjhGTBGJkvbMgukvQLn6T2aUOy8Xg+i8
FE7SBMTEiS3qj/irTd2GV7F8FJpQbG1DzCJiDtNHakQKkYdbq/wbtRgZY4RTSGmEJZerCXj4JNG7
l0h2aUL7CGQo8acbvwRda57oOc4ZaHE6vLoOZJ4CUdK/2Ffbxg7UUoAEaVF9HM5ZyuCR9eD2Wpe0
17hqYURXzkUQ/O4SWXU6YDfiJyRUfr7JL3zGwzFtNpY37v44rpe8DJVUH6WBPEnzflB2vWghpdwO
u6UxrGJ39M/W88yyLsunBd7jqh8dxZad6yOOxjM7HpTPDHuH8p0d4fqjwF1GNrXryM9wlWhqVEzk
XnjfVRrCIhODKlIkXIHXclwALUM2prAt2gPtJIR+liaYPXjuBiWu+ql+McpRD/9pOqrIBjfymJm2
tlZb/X9TVpPeiBQ1vV+1Ew4c0KH63KDMwQk53Te2Z6gi7Y7y5j7fjMEEEsrr0/qoNWO29GBykXCJ
G5C7AhGezZGzK32bFkqKyQz4ySvx0qYtDiIF22NoaiA/Dan1GqVH4bQ5UW/q+GZZtjd0aGlQUNcZ
6IWBYpM+TtR2oN2j/3AIUuh2Ah+Mvq3x4l0ez8/At7/1bEDOx+mExxfouvDccEBrHCl9DGIISm3W
lEibDHaouuK42qYFxNFm4N20M3vRNg6LtsPh/yapZPT4KN/ciXAkdlpoTj1GIgN8zzPBvZeqz3wq
GFjqpe/KexoWmn/g4Uwvqhrwg2bLBSt5OsNFXTaQrITOE2FzbEzkawhtZ4uZ/BHN7Ly2Ep8YRp91
s2Bhuf+5ortrD+B3+k6RbqsfI2mud+VXxjNj/1JYNaPql779H2lgTOCj1d0u0KdVetNwc+FJeAwW
+9xr5Ea0EVH2tWn850TtnUaVaGtuZ0lkr4ZY6lCNHWuiyht16sf7BiBhy6sufBBbXqFGArpFuN8k
2l4KP9xoF64AGtIqzScAQXym5y/i3FHryt4DVhjVgIgTFMAfwdJ0vTCQKFP6BVMncowgw7Avrzut
4IJ8xf/AyHoWFitlYtFTTxNhu963xWp8zyXbCyu0qnc2GCKSoUuHuIKktMAD+kfFvzw/FusjNafc
fbKCMu9DJD6LDyG30ZzQPVRz7qB8DWbajBEXUAGRYoCKdpIhk+XzosXsP8KfXA97QZUMUT9talVc
VCUfeAQvYRElPkeBWlMo5bLvIHytm6vMLTQRJDykTcrmtzeU6rlGSblN+eazIQ6GVEks4yKdMoz4
yvFiMa6OiLRRtel5UH2CCXB34TptxWwPZv0BUCy5dIpA2UM0uJk+DBQlowflnz8Wnxxqf3KJkMej
501d+V+pa8e/g2Qpw70e6S38U7AfR9l12JS0LroaCwNRFgJlordShHkeVGtepPbxZUqva6w+C1KM
/R2uptO3O2pUdtS6+mMyZ7hR9MRDkVVJ060uj4SVp+l8r4t5fNKeL66QMW0L9znSssXNZMTVQWiX
T+Xh5moaWIe8TPnuXggaKliye/wZ+74di08EqlNAIyu+tI/h5+C4lU5EFXkvR4atY7F0w9T4MmmH
hoFsMbRMGdH49NfmKeL6x5n1IrXUHmzDDabRGN3YxrTykExTDCxv05ygrEx6sG+YMBtheJc7T7le
waOzS3NowHP8GKb/0yhHFoyQJ5u76Dt+Kyqyb4MMEzCgHHgBQBNNuHrVQ4SeuUQJpXlMmtaqlFzY
+gS0u9Hd7mK7GfsSfgjbxkyEMoTFWclBsTGghwcMErVSRfb9kRxwbC2j56IaP/jN/9RHeWIVXvSS
MUj8Zp1zwYugDBY87akDM2EJj3qN4zgmJ18+AwPqseb/oBQWiJk7isZRZnmk4PyLoWO//IyK1WG/
5t9BaZcokZXPreUKLo2JEeurt0K9FVRbOWuCDP17l+B1Df/5DDfsn7dET0MKjlB6SSYsXrDmwzlc
hTJqyzjK2YFzMe0gR9sRiXdqUEgaoBOwefCzwNvr2ZVwNk723vbX+48u1PnNoQZZUiyOcYRLgKK1
O89ZHUOlbwcZRx3pobU9L4KK2da5RCGjlAXKZ2tNG+a8ZSBR8G9SzzfPhYwhlAGq3zk1zJsVPdf1
baCVlJ0Wz5YjY+qCNSezXuPzBixmsWWbMS010OxDQk+GhURIGyXM/NqBOYyz8julNHt7yXame5Be
YzUJUbGc7VxhDPLjeDtKZMkQzWaJZ9k7C6NWQQwyGrf/pU8KpuolSmxLUt/FSCa9frUOoj0s0+U+
QbpLozWAgBZ23SSzCrEPEOpA7A9HnqRi4+/RHOcJqmX+pyngZ8bOH3ip2iwing7ys0E5rRp5FLdq
wsCtmiSlnha9PomQujHhla0JgShHzaNtIx8+4+Z6L+hSo+niI+HTTuhn62vIH3mU8lqlDxwwU/J0
unvBcBT2fzcF702IKxQhLBJokrpktSagY8XNsYUFJYj9TbHasdf/TAb2ferNBZ/dis3Ces4MX59Z
iiG0xM3Kl6CfhnXQRcxrMEwcSaMj1khKC9iPVKtcApEEurq3Eikc3iAPiz2gWex4+ArHN8mnFqcU
xlLEOCvrOcU39qf8FErf2esRhIqUjhFPvc7yZVj+w/xI2wqAWvPJ890VGAzBQG1w0eh1B+IfuctJ
60wDg/cbDZM0L+Rsrcczp7uowlHF1hhQ40yctmN+6LpZlJrQ1s8XnwfEFtHtyBEBV4olvrf2nmnX
0QPdcarRqpFj3dTDULpK+jWfb05sf5MZOZLjpCIlNjGjXFkam0kWbx9gzQAVkpFX1R5HpgIqcT3Q
Spwqqi1FC9Dr8w++F2oLF1zGIZw1Wrneh18G/HWnUt69YTakP+fvwBfJoxR0pTekxoubDI5EYoRC
LYxIZIUsFeejWCLOSs5mItEGZWnFRvitSympq07tS6CFAN9IjjZkZG/XkFsa9jp/+/459V/Zu8HB
Ov3OzKtGTnoZ7Mf8NyCcqVTV1v7IZKm+lvot/Lkcz0E96XCQvmnmaFGcqCJagazUO3m385nytHy3
VuXVfOc9OLJOU5kfdbez2WAKtemTiklDQClbnewwhpn7rz16qTfVeT8GnuTACFDMEiZit5crNtvo
NFCnyBg5wd5kU484gOui+tYmQAXQRErfkASVOz1JSvUd3jTClPwgEWV1rfFBGruLOa4k9Zg/7R98
MfZ7oLm/LjvgzRNGxReo7ULmskJer303FNJiHg0Wa+fuK4yberYOZamUKYjGxwWJRxXnI6MQPTJw
xShwKBqb6G4kgQY6buRb8L7ivtd9h0R0e8U/gKSsm6cljscaGuQHpMovg6gNsxp9VQDpsqRbQ732
+a4SKJDK+3jjGEom+0ZnVt4dmtJXFceAwYGKIudBfW91eCfAWZJHBsnn2CAzEGqYmftg82iPbmeO
T/YEryymniBfE38/pmZ2i6I1lowb82/+998PybVxD5Vg4qfaVjifP0LGQeC5l66jtKE3lf0HMUX6
jc90Kuzf8eku40CuJ0ouMVzfz/fK9mPXLtMD1U+v/3I7kvsK07Weeh3hvE0pJhp9YT2J6Qb0ewG7
QzWMiIvQbCygPRDP974vA1xs0kxji+hAardiUyS2YP/OHbI7Euu1oCeYtDUVVBopd+Q0otra1+B2
bdADfOq0PeT+OFI5MEv0qI1oasauWddq2hChXUgD0MNs0E2XYzTVVZwdDu1+fjNP5lRqV+CqQgQH
8TvQKGQJbFpkmyzlmdcWBlEASOzxPrsoCuHnlJ2My7k/kkO0jcwkxmdjA0BYbHanXGkaqZDZ/jt6
zt1zVzu5r/h8gBfIsVd2K9D+hd2j43mFqY/ODQBbfN76DAXIF9cJvoBZpHIxn3fJgzM0vyt47NJe
OacYx9/IJIKAANcyNtRz+9+DLE8cNrAVX94i5TL2y2WflcmlDuD6hjyq/h16BsTvn3zJADsh8Bct
b3oXz4gYEdojoHlxpq07545cNuE1kZV+zrglXSLKvUCXYBtV8kVqTmzdNfeg6X5wAGHEZLvl33w4
DM6sau7SP2/yuJOPx7jYocF4B5Bt11mVQ1PyYh3vz9/DGCFAahFTUsG/N8J1vqmN388PEgDUVYs2
GtMIZ8gc2ozHVLNRG3HDT2J6V6Aj0j0zs6o8K3X02vn9dAYS4uudkmxQSkoBuKOxZPqgdGLF1UTc
zYcKSu0XBjfs68BOLk27Bf7qKT0I6ZP93RA2qzGImmDd0AVFtviU2depoLZuaKhw9i+SyKZFlZ1G
NQbe5t4sQFg/Nt1R91diNcI93tryybtlPL2LrHzvNR2WfK7b26aP2bmfvH0Vr3DTLQfD5cyxTuLO
rWyKotnBw9CeK7XJTwyLPSrCLjNuXM3KqEb+R5evJkbFpEw+fTIBhdg1MMJ7xDj+CdHVfXFPtKEt
nHhaczH7duftBrmIlBr8Sabb/nXJRj1FJshzZyXrQDPrJrgKHP0ZN4SEamEp743kTFI2i+RLNazx
EvHIQes8pXUkrV1n3kaLwKmc+rNoR7JPJxVgJhbyNzuX2j7Vo0FEHm7i3CExmKvldPcS2IoMLijo
dyUI5xGwhn7TUGL6MYtbTpNopGegJCUz2B9wZ3RPZskIQkHdzC5vSj89yvgM8nuN0lFhepxxxaPd
zg4U0u44oPWtznmx7bsrDyLZ9kIJF9Mq8LBCAU86hCONZeF9WQH3u5rWSotqAxHAjyttrYd3fA/8
bSD1fPLP/lK1vt0gAeCYIpxgkxVffPpEf72KCnoUiZzu2BGo6bDizKwm32GqrQ1WuASYHkDLH++y
B9f3U0ZfYb4CUCw2lWarLGLukQpQx9ytWx4PLJdiOnY4bVFkjJQFCCYc0oP3Gj8HfBrYpb19JdO+
Wm0KdTYD4Ah3wbf/QJP0vRQvf97DLGdeyQ6OHQSq2DVwJfiY0mzNuYJcGQ2aoL/2Vk0CaWHpnSeJ
BvY4k2Zev/QzcqD4IeKIBJtBQ/88R1ItZryIu6Xw6R5F0jkWxWKxZAPOFr+E04Q3H4eo0m3jU+GX
SnRI6PeuMnVqZAPsIx48oUdRADT3+YC98S6cekUOCQ1k2NO0sJlwhhKceCqKNIUlYRhan2s3N+m7
Ic86MAoK9L2XisIz8Y8Q/hDadkKmJz1dEFir3zA/lH2h9CHFaOLRZ4bIvBT3tH03yyir+NBRG/fV
Li20lHkF26PuWDJasxdDGbPFb88Z9+P1ovjip9KT7zJPv0td8o1w6rFAFpev2QF2V/bs+lrExuw9
DblSkzjSPEmFVphChWl0i+SPPjnDfTiNMS/vV74L6pTcR9d2XrA6tS/XMBir5UZpVyQ0ff0LXg7Y
Kg0Qp/bwrYPYdlM8kzKjKNu/I4BH0smpZLBGb/uUOz7HaWAA6dcc9nlM1++m9syS1Zy8YxT68X6n
SXPAi23DMaGxW8j0q9AdKBYYgKGd8+/fkEf4xL1AP8HYr16yfeW7Etmw19QXE5o58q1sLNRs9yaT
DjET4qjvm+cd3i1PWC9jMg1n3K0GVgfmQOSxQIIdpNgc/FNmjjsrRkmZfwpcqnd60Ieidbm71FDD
0zQsXlvNG360JP0VQgSo5lK5NaTu6M+/9UiJukpg8OX+ke7MDPHHc20DR/dNamKwrMbL/iUNW1SH
NGPGwjIqbLi962msJGzADTOpw1vhSWDPRDq2TCnuUhIbYPZ7KoQL+3Zc97DQCJaf3U++4iMvsb/p
3yir/YqAXRPcHMatGupXmvu/D/isyuXHTQ1vzHHzRv7xH/xL1BobRqiPo7AQu21ETwuHGQgtrDVD
LRK6t5/TqFvye2go1eUlJ3NdZM4/WN5DBoAkmbX+QrSsAz4mComQ8FPizvz1PkzbwYewka/tJ9/m
1rNLat3br9HMKmtALx8sNFHIU3khyfYyAEsOXn3yTSHhwla90FmmUiIjIf1c6SAehGCt54bJtDt6
mUWqB39Sn0rT6N3BkxfCr0T0M9o+9SEKxQj9NLuYtgc27YoN2eCo7G67IDDv+RaUfmbWGW7UDi0E
PZX3VfTPNw6ZuxS86FUsw7hW4makLZbZ9Pe/IFGVRFkW/YrpacpgfqMyyAPZNevkmHIDqn9uIH79
cVb9K04XCBanVVMwDVk9R7i+cKQWUqiI4isejjluWM+QxO4FwdIKaFHnO0CnEcEgOKfRyDtf7a9x
BQNLwHFoFJyKUpPTEb/V4WClq5xhq+UZ0k+5Z//ajq7yx68z5vYHqJxKxVT1jm9Lo06SVf3ZlUGO
cjG9ElojJt4Jo6DjFAI/jSFMIxIveWQ+bN5eqiudQlVllPfqMTT/u8odwqk9cdY6H6BBEsJEVWs8
Q5JZvX6KAliSBd0Ar5uL/8G0fS+VbaejM1eKobgRsoKNXUYNBv6CMpoAI4sqtOb1uq0Fvyfd9WNg
ZHEqFQd52cGX0HzS67ORYxNaqsA/hxvVW9yzkzMOED7wD61kzpUhZZgrc8uTyNH2KMAgxRWOatZP
pC9JvNtTy4uG4crLve2zl+XXPWfU3dhZAAFVY6xqX3HoZdbkTskQyQZESFGotucq8rMkY15VbaeB
Iypi/32SFpghSaFBzxLwrjvf/70VTElxZfQWi76e9EGOXGiUXND2nf7JC9lZDngobp2U1gw2kGrs
29Hldjty2usM+FajRYSErPOkmCJBMxa2i3wf/FvR70aVReAKJZ7BAABHO55bZ0NOV+rpBcHo5ird
rh7ek2bdC53NXEH58PjM1fD7V2HnHR5aodiq85rn5C3SRBRudmD79r/52Jbj+WhS975zi7TXdOMF
jmXqzhWWBJiidV5cS4AnnXiOsG3gZ877HchmzMJnErYP5A6Lv2nI2M+L3ypebvNH0JEsUqymD9/k
axpFSpylPSX1pUULdq/PzwBUW1wsrJyxYLsiCri41HAtng2b6RdpHmhiJ0b0I8k7qduPN82BqHCP
jUOgXK7ehqHgikL/ejhXiSYk+ZL2orOfFL5lkmOyNrOdObMYfv0J7jQGh1pHvc99846c2KezrY7A
Pvvn4kqcjZPD7cX2tI2WGJg0hBkh+xgvYA8C+jHkzTyMiCgZjvH9I00j/xzaHsxBF5Esrhmziz2B
3lhPV8+IMyuPw1/mUI5lU8nFMgnvr6VtvSPljRKK269MJqpE8d0YLtC2teSMy7cKXDtVJw4f21MU
oN/yMUiuR+eBI1UjJF6g4vmxWgPbWeDg3bIDG6whLT6KrDHsQU0aP3dYXEj0ng4n4pGa2/16zaUf
IMWQkdrvzGNZIe1rPWPhN9Xsb24u6RUYiWcymBQZHnCG2e3zIL6cYqWwJkq6uA0z60EabL+fDBhZ
rcdHeiqGBwd0euy6tJekgfPC/2rz3ep0BMhLYaN6YOb83eCsQDOm11KGN0h1F5JK8EdoF4ZYXTs6
OoJOnozwBe8p0MKtiMMR4rrKngw/VqXIyzRmu9yQJAcs70C1WJPhFh69SvPaTHirrY7n37HSTDfR
dTO02gyzG0VW1/3+KcUx0EaXUDOWhR+Za+U0U0gwWNFw+BGozl0Oi4Os2ubKigY/+yZOxTV22jLv
UjPWt6BS1Q79eujPz/de4hR5mzLFlAu9yF8C1vijcG9B/ayjaRSCt+HSbbM2UOIOhM40ywxqhFkN
mbcJyWIKwNjsuY8nbjBfbpJTFtPkx9y0cOQza5sNUI8rSL0uW2Qt4c9EzKUoqpQNZtfLz4x/N8p6
pNkmIWRy4o0yEtglCVdNyGxwyT70z5p7mjhn9JV4GycTH4OXJeVuURxSczypCln+qxgyLlMMNoKf
VzRfg++QeE5e4bAkKOTrapRRGm3pAcBHNU2iIDx3owuHRZfbU9Y/KlMI6TuOyCvEO3bYbT3pl7bt
3oR2cZwq8+mySFNZupqIiIlrUMOnJtOG9/2fcjVDV3Uic3v9bk6ZOXqBwsueIfRzrXZZwPR+gErf
shb272bVyQ9PjCC/L9taBRDPb966KBsZa6JbPqLJ4lRpNIqudC38n5AnppXQewLmlxNYdYBcRlwb
y0s+FbMmZp6XblDZYQws1HZa61Rcc1O206gkEwIhViz/FXXMVQtalwbMBijJ5+aOoRv3iG0joIpl
EAXYedlEpxzA+h0F8QC23evzXigTZrdKrXCPVOTJB32nZJvx/Z/16jQ4xnS3vcXlTSCEef1sAHMx
lkLniGSAF1wL5yhkGqaGjqrkCJggLL24uGevbUYilMIkCspJESWHkIj0Cq1pgE8f0XeojW1OtP9L
ncqMLF0TL04OuSXkuNEgn6robC68XlQz940hpT3ha1kAK0esV0eVv7+nbHO47vaNyJd68K5TBNK2
ZGRcIQb5x4FpZR/Sgjbt1ykuVcmT+iwW2wpRWDJabHIt5LRqIO5maTMzwt+BGgVopOHJ7W8KnQbB
UNXviU07/oIoR6S1AC/VaSNFSwylBhooBoxLcpnIveJkHLBHGggljbIgpTi3qPe0/VkzMZuYmxPX
Frv+L8eDmpwqc0Ey15IboYbXYfL7r0rzTUQqYB2LzRQtqumLOZUq7fRsmezrQDLLlZZ+gWMt4oqV
WwAGSWJQD/B6sU/hSlwhTg/6uJhedUc8CQsefKRo2PnEGGt6mV9vOV1dEFyiywUskUu20JKj6L0k
tLpWF1S72+Y7AxzWhdwkpTto+nVxz40SA+CyZAlIpExZc+htfjGwwm1Fw5yjcRoDI5Z4ffRj8i+5
ynwXv9tQ3CQsN7SdRh1LRnCJK51RfVwPR7DJV289HUXqCRSBAW0hC0JSokDmOpYpe5Uks1eWi+9s
OHFQHoKB6yi6oUHTy5q+Jfko2qUxDePg4XaT+g4xMwBR0kylSJyWF1S/bw83hHBgOMzDLfoqSlso
YpjyY6TczbGXokQ3xvWcwyPNYf8WA3XVZBXz0OuA9ciVLzBf/CFGSGPHRwng2KI2zNCOdQh1NHeI
PgWFnirCRx9FgKonMohCDg9HK4wGgp6zPKk0Jknczf9vr+YwiENqWoDEI7ZUDs61TJhm1Gr8N/q7
wra8vUQk9KRbrl1nl9KquiF/LQhlBf+1pqjlk/VRFoSM29ojBuHAbTNvBrDAiZYrPLg9ZIhUkJ61
2gsOaG5PsW/ZplOZOs1hxDlfDjS+kC19gw5iQSngIuJTem7cy7bkmDH7cpcKxvd0+Ki8OqHYGDKs
KFIL5xmEKLkuS0pSs2V+pqg6UytN82WggveN1ENl/AzISVzfzvEm99z2/a5OpsTjDD6iDP0kXOXC
XbZzc0oY2yl14JgYea5igZbsTgWnoRCuf1tAfkCkZS08/Awx7kU8vjftu7EFO5coh5qUUQnm2Fcr
/7H9jEYsr0+dpKegW9rEI2M47iT/h80oudRyW7dkIk2tEYXI48ekGxBfERLQ3tXcITsHgWjRxB/b
kFVp4qvba/saY6+K6QD4HQ1kJtEGtKn2PvvB9C2BZgffysAq/cZo/VH///gheeZDg3OO91cbKCFR
3apIO+gbhdO1Az1B1ebPSUWXh7WBKHesItxZ9nISsA/rEa+wuUH/wJhlqwhX35BWvqiHiFv0N7EC
OtVKA6ehbUVfufIviBJFVNOOLL+NLWNBInQTP+5n6JJt+1cEFs8HEo0pm3n8zaRHWWq4Ax90V1LL
H8H+fO/heo7kd66DzUXU9POjjOTvD7j08CdGhfYAlt8q8StJs6iXFRu3UDlNoa5OdBJVA4t3NGLv
aZLq+Y7F2rSeVWWrm9uNZ/2Wzj/EpX5GlQ0ZKeTcHQHGR0viyCINiWxF+VcgJwbD4JJZO6dZGA1K
GP9+6/Gl24DKmbcCyfsJL3XdZ2KJVVBfER+WvkSxkKggoyIrdU3ywIsf32T9JZdXvdgJ0JVjFW80
p3o3QOMdjp2ZTEiqRaosAbxys4y84pMlHSMDqoL9w0FwS0b3bS6/0Ox5zovZNCOEr6/mCU3zk/rz
IkT9Ghbfa++CIxG6M8O3uhoTiSIRt+ryUh/+7M0PbRcb2HIC5DbedX0SgwETQpPsnFAlXTzh+EL5
ERZ6dL7XfPMjD9tpxRf9XMPoMb/GuU876RgqOG7WiJ48US+K/10++p5HWh5CAQTIXefvl+j2i1em
7on+j/9FkyftOlyS0Ej84IjNlN/v5qxoX44CrIJ+AWi8O5HeTLqy0ROBqG/U3N5QNhjnglNlO9na
Keb7Me+YvZ4tUOZd10NllIjutdAFmwNFKcMtz0eflIzKoB9E6c6LiKvoqACXD5aKCZtI4+KZQnqF
XcpuGP6iVrlV5yN/beKeZhGjRy6BJwdGolc3NunTeR1lLRry8hju4v058aaeyD+19jW5MQVOI7nC
Ky2n7Dxmh8nBYvFlsi5aa5PDrJEvAweloXDdS16d6tCj5Y9rAI+g+cVGQjc4lP0UFXklvfeV4Mgp
r5c6+hQYfomo41wQl42yXZZ4FLKahjeRnTR/hjykbc3Hx80iDchwQV5Wb31uDC2HzLn2Q/HKH+7z
orUJWIoP3yIYhTpvoCkEt87d7cvZ/JwCo8jIFcRTQC3LJYMPfeeajxk/qWtmImmUf8FAmTzbh5Sz
FdreesGmnyH1D7ZiFXcqOPqZF997q2pW/I0rjz2+cJCegGFdsAcwobkegMu/gDEHdLxUYLl7RVGK
RPjgwbKBTSvB2jqvpAg9FvD0PHxsx74l/hqot0NgU7AD25h5ZkVGpRCoSmvcPc5D2Hxg5SgbRlot
wyXm6mhBr8q5tscEsqlHU24JenMOmDcM3x1ceHECLJensutY/tVP/pZCP3Z7C40B7ImkSovMGmP0
j8gQng2ti3G/MR0RscQXjsuZwyUTfgWivjbQsA7o8nvImnK8vzExW+ql3vFYBo1oUnzonWiHibZC
f8DVryveFle/58wWqs5rm8y0z13n5/4ycbFe8Eho52UDoD0o8flSag78+7Jr10SEcbUXRrgFXy8m
1KsWT6gNOnLzYa/1NuC3BNxGLvZ+I8CR2TzbHyG0SkNzgp/J8l/CX5OB5inn3CXn/9W7eaPwMZHr
4wqWkQ6Vz5B1/t5Oj58qo4c+RJFb0nnFj7AB/drcn2Q7TPPTA4/gs57nav2TMa8cnDfu1iwLPjvA
jf6EQjo7H9zNxxEm1OxsmaB1B2YPGMdvtiOSkvqT6Xd8e+XcrMj2oBS61fKikfMFzPk2sgEZ+rBm
cSme/JzrEFe6nBLxT/iV4cUlBTZoqwTieDHTqbcP4vxdR2GPmNKbntTqdwogUFDfw7GiFlMSqkWS
cWGUTKJwJAUBlz38zePNCF40Z7EtH4DwUbU8oNKjejCAH3rycCFimjh+DyS7HPh/dUpLEfOXuffj
ad8wmVO93sOvyHMyF2MxFcxV/2TVrlsSiTMTTFODsVAREBwE8TylUXpfz2n0zj+I7Qm9u2KgH3sC
Yz0/ZGWRJt460UVPNk8fvz/1VZhnYYAyr9eM8LdV3DLfjlk4x2IInQW7Ho2sN66W4tdympbQxFia
ZVR2j7qTveOgKwjQ2lu9HKqpmTEuBhEtnq73IXsvr7A52RV0y2Qg0onjkOlvDcXF5jRlIUuvRJD7
GQa0bvQIJW6O70lOmcomojaHF7CwHkwZvOxVE8xbVTAo//04ytqZyC8oZKyV2t/TgGAOUtgHyoAp
jld6PbxxxFkcEJnR9VCKNUcHwRbJOTb5YvoSuBwnSz5HPOCL/MbQROqXK/MXlo4lDaVAjuGB2RJA
ITCfJKMM37Qs/eodyJI58d947yfe02WfvzV5KpVJmvGXtzWRaNat+1HmZ6KnxB9CUzonXpx1dd2B
9dOqxd6bkr14celQ1pffT2otdC7hgkuXh83o/+6OFn5vyLLBTsxkrwHkl9NIrqCPa2fh3/HGnFab
4r045XQA4W8efCI3Tho3phuefiUXeR7DVx/OuZVqElTdii+CgCxA3P+7kTcoinppI7vA538yHsqj
wDqyP/yFAD5BViZLZz1Ek1gIhbzPLg/8lJkWhCxl2cdDIEHs7Dwc7DSkeUn3407eNFhoLe0Z/z+/
lU/HRpsSDuJXJJmAa352jDgdqUlF3cnkABQthIFZOvzAe32KJUKDwq2ksUc9mp50Eldu1fe0/wfj
8JVGj/yEgaROhbqvkk2Pt6rFq4dUTLYpRCCqCFdDh5igURmE7jAeaWDoOZXfAVIMIeGt/aWCTL9t
yzInOScyyjY3T+X69etsCNNcxUk8aNwOrSrnGQae0MYvinn3pxi75+6iD8QvH4iO0oYvGt90Ybb1
9i1FJ5umiy8ZvuB5e9Zl0OTn3aQgDO0aEga0vKIA2qNmeHCCHVEarPITg/F01NzghZzmf1s/kNHE
T32vBxGqHVRoMK+dALzdYIGZWK0/HKNSrarZil6BWGDRp8DUBrdDp25V6kvbNWFXfecxvMUS00tW
tEkjqJzvg8rTpyIOOcIBFrnnSdcuf5VM1g8qtQErrOAKrelRLcH84/2DTmaHLDlSYlU5rDR5qxDK
moVAsCbH+V1ax/p7RXrKV1XPXj3gauoHd+U7LV2zWXO827U27R2j/TlDMn21BXl443alSk5cgJS4
mGKs9nPYEzE/y+Iz8Ny9s1JiPFHB9oFSJG4InVwfvMAs/dbTOr64QHEPxHhyEc/9mtQj+FFXd+//
x978xrYteafPIsCOi93uPfi2KyaC9fUK1IsftG2LdPcwCHmLMaSbw9wffKSjggPFTgRxLqLptv0D
4Zmme+UbY3LskWPBHP1ST41H7eHB7jp6Plxd2xdaXG1DD5RSvxF49QYeqamaVqgJebUykIbHc4Tj
wg0/cZhW6vFJLdxZulht0LLlMUMgj61F0y3ibUNvZDLcLGtLQKy64r3eJ8MtCT3SJWDkPiwdduE6
7J0mBu3297UrUga6kFMmKWxB/D3FEFjkjFC3z+YX5hPwV9vm9kWdgxFUlZJBmJKxGOKTY95w4rGs
52JBtD9s6Pm2Wdy4XMVfzz+H7FSNOBC4iCw+t/92UoW/Ut3IuhRzsvHSSaS3JYPuryrJLyT8Zny7
xK0AonmFpHc/NM6QMCNwmq1Z56ErczM8KvkvD2hitFV6vNxTPpx5164K+SvuboOx7oG1yi0YD1fZ
VTr1gH2Bicnbi7vKQKUWVrjIj6awfKytjlvhMJuYg+cA+ooDCz6HTNCdRGFYy8peLKNfCYNbIxZT
XbydNCbwjihLLlZ6EJtEms8KRwUw1g4WMiNBxwwTV68FujDtBJQYMrIkmXwSPTnPc4yYFkJL1wcX
1CwtO5TNZJDdKPqYixLRxSKlzb24aRPlkG+8B+g8s5aXfZ98b++8PaOOor2wIsSKlmZvotLq61mo
GBDibsZZhZJ0x5icU3uktaMfbtgp4PXH4g6WbWJGRwCQ2yZNnnPOR5eANh9a3mRUCei5tOYclud2
K0bmDlIlGVEVkb5RxiQm2g3ee8UDWRPDMEEjsxeWE0gdUgC3Y5fP0FHuDokstbIb+pvFGUNHVps+
nf8wL9xHpM31JXLfIIroPhrhDXo8OJL5ONpIg2tvkCDj4a+0w8OuU5AyXuG6afzOQ2fKimu8cJ0H
AjJvvIORd8J42OpfDMz+n6gliD5q9QpTspGJN/vq37QLi86TevhcPS3W9Ct4hBQew+DRfM2YFvh3
syQ4s9OejRZnO0SecLNftfYzHfLOz/9adGYE8FM50/QyqyjF7k146TugQf5OuCaAw92rwuxI0T+n
BkloO8fQCK/b6GCsJDZB6S5iz+59C+/oFDBLS1ufruaEeH+S9S1jeucSObRMrjXSS9fzs7ohV3Nh
waUGjZpA1MMg/wlrmAt6UjHCJtUVc1NXMwP9lWev0n8H1SRl3XhrGRNO19Pu9ayAVSLvI4gQxF54
ox8mpNiDDXfBO3wuqNKug4juuqpWhMhms3sCbG+guB4AwBojM5/ShcFxgmR0PqThMNmwmthOdFdl
8rldtylQdCnlzvVK3DLf/hufz/HIAwBEMbaZkPnHjq8BlUfmn+ppxs4RMwetOIeKuWNAHKaNusDU
oqqA0m2s0FEQm4f94P0kkDzZvc0NDz4DKBOZK9CQldcrCRb98Nf98Tv3zCDjWu6TaWtpe494KFhb
xzXeDqbPXZB/pdhhhqkXNtoyoK+UpJhUSYb1p9Qd+B/u8XYhjXmtEUM68eC938MLurrv1/MA1A3+
BftS5dGWpTSDodgFDKgu9b6wVLGcgfVmGiGfKnzubJfccG+GcPorxhU9psWEsOQF4/kQ2FUafXPj
/2tAIz8Ni4FvxtQsTQnrIRpMLbnp3PZavVVG8dbvYjy6pC4Rcxk/kPTgyVXZ3HmD5MohkilYxq8q
0oKw0I9RN70YgJhkL6Tf0MyKwZP0OJxJPWGxJ1F7LxFMPaM70xH39Oqtf8Dv/7iylMoSLSbg4waz
fx0o1FN6d/vS66cZhpbt/SW4XxoQwOcIF84lZa/qrz+0yv9lqvbstV8ueQsXHZ7FrdsehiTG75dQ
3TSdxJ7AOU9jfRAqDfnVod7pBuWfRFfwwWUyyBgPPZh4kp5tH9rkLwXgM8rsQsfWk96GTfgjyg/o
FSJBuQ3nF71ERPFGnb2e0Il0A7CyEnMrod6A4Dd7SZkf84vqe9NB4wzPVTabcsXIom+kdhZ89WHw
e74sUp2pN0i7CtTI4RqVX1XKDYAYA0KDauWhmp5hkuNdXnd7eKvvamIQ2Mvpm47TBbRMyx5P5RLw
lePt68ro/qG2yHzse449Jb2By/rBOk8ZQ0YAf6twxCF98h5EVKuhqf+eXanexk/TtGDrZrfN/MM2
hYpXTTnH+As7JA+Py8Ig8AJV3sD7tZosYCtVPyMabd+qK8R4KQjRXS/Dxetqt/iSruJTF2dvJPUl
ydCMyCCuZhsjNKpYDArwfE2w065bLQtdpazV1PmERXDTAwwoa1kYwy9DZcasoI9TP0VikwI2ld+1
a4jkrdnDY/0tyEXD/RlqSpwQNnrRBHDC9abB6NSCx4viCeRbWj+MnS40EZU5phZHnXugu92wai9S
5vSTpxhpJW6C854pymPzqhbxpJIw93U6usTCOCY+rIYJO4cCRtd9IdcTBKhY79W174/6A/QiVa02
rYL6BTU1md2u5njC93nbIu+Nvn7xZ3QYH3FSEW1GcJ67rT5tVxv1zv+f0NrWR1RTZ3VOYmZIMfPX
p9jQ3fP50ypVczluXjMFb8cXecmSdukSghV9orktNLtmP65SDMoNTI04nYH1Lr9aVb5dIORdmFak
CM8S5po690tv8u+o+eS6BPdFE7u5kET3OmH0+keOR07TEICRIJ0SkAqKLBcVZatD6L2G+TkhtJQ6
xZgmGK71dNoRC98796EC9uFg2DD6+Sn90Jt143yackK2AFQY6ZSOXryHYa/WavDFjvXUh0MTwYsV
L1j4xo2c0K3xoJmH0EYONbeigelkcBRTUuOab9yUjk/Jm4Vd16gMXONu8qmfAoHe39ZfaKpZ+lvp
PHQi6yl0U6uyLRV74N/BZVPbJPMzNAMekGu9P8xh5+7CwGnrW8qlpMHh58iwvWdNqrcYZcSHFa+j
4prxsvGAa9nkIfX8zN4/otdRUYAsFYh4Z9DFCbtje2+A38Uiqy01ZPDBHRyZ1t2qX4asas7SfhXi
vTe7wVx9xAARZCajA/Nbax68HKBvol3OvasaRodop2zrSziNTMg5dXtdX245xylww9xDetkMs/gc
GfXdO9z4eaGV8FJilrYWx1GrNV9lWjP8e2FB2+B2x1mcaLumrRwYx3uJGZ8b9uApEq20f1sFTM1F
OcMN6q+uEOy7oH4UDXMIDdg6Vx4PHRYoI4TrwpO8qWKPXEmOUsq5O1+NgFhPxegJt7r/et3nfL24
1Ofp3rm92/pJ4jrgsWFbOMqdfWPrNVRQMNoeB6JVDHDvN7K8u1O35Zo1RiBlhc5MiHQfLY0h3t5W
A+8PsI7IN8PM0cvyO1nhMjkoxmQ32anxPc/U581iij8kk6+b6HNFkm1dV1ta7vcdbtWe9IQsTRM7
TLx5R5b4GA4uZGGYHhanr+/kv/0hUvp2KLFyfLc/KQEFFEjXU8vmF8tsTNTqdEIeKB7VegSTnPYO
cfpfX6V2eQCdnqYOpTCm1igKO5f/KJBGN/TkNDExmHBA0MLUtfmuqxBIgJA57LwjTqj069ZI7/st
xdfO3W9BxkAbonR0y9PKOwlDLubeIBSSZ2ouVGXoqxzCTsvu7dcOvQcBd2zAZrEGRZWA+GIJtGdB
D4T9LDTG9DnlQDl0y7wceL6tMkk7zrtIW+Fw/tYij9bUfzt/zpUDMdUlqjGlex3x6Ne5lBvGnK3A
PszPVGF+5Zf1lr9wcJoyakrjDlcyf3lUt23SHmNvLVwLgF03SEvOQK3gHky8+6TlhEXC99ni1Brz
gvym+nmPWp96B3EEjB1BORJ6/KnyVnN6L6KHLYOfZncD5N7QtwrnXHmW3ote206ezR1kAQIz3zMD
XFsVy99DsWI/rmYCuopuVXYQxhF8lAmWX9jpKNP5I/c8ZaJvVgLxrK6IT+UBJRybi+D8q834zRQv
gBkwF1VFhqqrT/D2ZR027IdZpV4GYKKKlc8sZ61kzF3w+LrmVl80+zk57j7P4cr9iq3WMVbIGt+X
DERmEVM6B8jbJMWXSg0UtUSUGUH4ottcP/1PVRUnCpVSND+GolwT7GiBnpDNm8hB6HtuPGroQIA2
QqEo/6Ou1eaL59ToOJttSIcITd/SuZdWZatBV2LoY3505awDYaucYggenp27wr0iqsH1/kJS16+i
WUoocRUg4uhu9Nq6FFQB7Zej6wCwzGVlwiHx6uZ4+DZkz2aHO1I+idTI9Cz/ka/NliCGZV2VihnL
fH2R6t20OB+OCll1D4BhPhwhl1rSFEtWxxFpFZARn0TSAEFB6JvzcCp/7fpTog1Ieyzr/UkkWF1+
CXsSD1OpuiMzaGJQxZ650rY2K2vJBpgQ03ObuTDLjA7ZvYytMYcLwbYd/v5X+meALhhsM7uOLWZr
LDwiLv0xftlTxAlvMqu4/MEolB2d8P8Q+bwK/KVz1fEBGuKKe4dKGcWMsJt9M5dPVKIvC4R66s1y
9fyOdn3iTIQ4qBdAqan6tukKiw/Zxud4gMDaRZuSDT8HyZ4e+8UdhRQLc2lkgwnNmqI15+HYtwid
1Zncnft3jAUGm0A9zTB4F/eYNJzGvCyinoiUY7qo366cVXJsUVP1eRPHqesKXyqYMNfPiF0UnQUy
T6/o0vjFA0+OeXRQS/3HyFjZjfucsPwR0U3IFtzc+HWhGmDM/eGXuyK6EcFkmtTEYJTe1i8XPSJ4
uanIIVpujfAaA1q7nNDbcv+w1CsZZQu87FI8lVimPG3CZP2KAplrpryJldYyRiNMIfMjDMM+gs52
QdyG15D+VKiXHNcAaZLrwTAjb1p7oam1Aw5PfcOlW7o1ZfCajVzewY6pnaZ3FMK7BfeC13WRW4ne
os/yrFqbSTMoDdVWTa0qrIMNtukK3oijJSX+jPJCatdYU97WYawb4iG1YqV//X10AAC8ofD2SLWV
4XxReunm/xACjRfKpsQaNQUSK6M3aZS+GeU7V0NCJC2DWT4xx4WKezeqo3fawaz8bWoE2kqrHDVp
YZAcF2F9/3JFjKP8OIrn17peqp+JETsk/YJUeHTWk3Jz8bTEnDe5dvdUA8zVIkegiaQUL2que0gh
e70rRAD3aOsR7GdScG6o3oLp5qPrpktvm0EVrMVqLaLzQyrpcocBJ4BCJpE+dC8sg06Ejy3dD9wD
XwS0R1R8REXu6jrss+Pk1vJkLHmcaY3i2/jcnPGAam97vyU5VWWNM52a0yKvfQHz/EXf/WE5bflh
X0mUHu3cIUaSCURSjKRDeyp96adWEJZ4bXITbSyJj0oZ8vo9gIcvMofgm4dM63jXfVy2xT4EcHsd
aj4yP15Y7vVX5uu22R0hmRvIpKNYI53ti6V4RyNZW2EFboDYXE4lk6h73sSFQ9BX/gRkPdgBijJn
kKtfehmX6ue/uDSK8IiJrgCNUPt4phfGCbTi55f6TeMB8Z0nHP5uXUtM/p6gzwnla7tlfg8clWTd
7Ionk7UHrM5N8nmhKeC573m0NnCE5ApgjnfzBjmkPUinDbXFh/p6imtxgam4QnYErjHV9Rxko4xW
IR/jBlzNQiXb2Hozob99vXmEJIPf4rmoE9I98jxh94j7CBbxg9tBVyaHNnDYjzt1erQFW0YpLJcp
0+3jfYvcsSPFrGYYajLNeA3UdssqwRwT1VtdoxRx7KNXs2IW7NfUjO7tLzqF9bjPotUnWl9yQ03R
3osPY8gEZxmiGmsN5bX+03Kf1sIZGYRM2yFxUDQWOyXbEDcpd4WdCofYIdwuZCtHIBStqvsi+85k
zPLNkoKtRr8fAxZ7NA6BfO/HDusK6ZPdbPDvpXtBp0vPavPfXm1DE5WwwEuK+Sl2PF/Iuhb7/xI7
FuZSUZh7+I2aIM/5VvyX72i8Yb3qIVgTeYlLVBYC4QEk+Za+YjfvX7C429M90/fop/5gRFdeWEJA
rCoCYUAGtVECYz3NpQ4MPJnAv1Ubo/vfxnihTyfVU45rBHZaj4SkUG3ENvmnHcdJwJHok1RFODvj
MOANEY7kbIlc7phnDZXzenEWJmmran6gM+sXs669pb3c83EzIMfOIN2VtC2Cf8QtJEhsyZA2oJ2u
R4zF3rxp76aCS3zHgq/sefCZ2w/uLyXRMJCOhsv1qDOQNFxeu6KWVCbFzHfXKont6QZAmksAth2j
Zzi74ToGZm3+brMJb8gVwMh+DjP0rK07RD5Jzv8rY9ZJHyqmMsY+tr85kaxZQDb7CKPZ9Zn8GA9b
9vcweMdaImsEP+fhyK85yiOA1eDao+DTmjszj+Jk5M4wnQ7UFx/HSI+iF0zSAe0M3NajWJelA4ql
PaLPTX+VdqTuLxCsOsZp+0ECQ3+wb44L57K3YaHkg7qOmPDoK2eZIbQzy2ixkw01rpTANFQROFWD
KX72c8xTj8wlQLbFJ9j30sH5kMHi+c2N1WfQK5NZH3PJgxdn7Hsak1C5Rf8s3OjNd1oDcf4zf0bX
xbh2vu5dUVxDOh4WW8uiMErmnMndK3Xg6iI9MnLsIJp81H99h8QxA+WwqIMi/3z8NLCdbWzI/K8O
AHvD0B1tv6qJONbvR8MUCYuhwK+DxVMWM1zgdsjALW3WyCcd+HjgDfROe53rPuEEv49hUDq8sTAt
cjUJgmkDX1ODgO+1VWM5N0lmsCSrqUBxm3aDlRmTE6HGJPqzr6W4ULRAhaeupMcmD3hO5bfLyzU0
eThnT0pjcd+UroYX1BJl8Svate0xlWEptTY53dLCYSlCG+US9K+x6keERUbozBIV2GvamAgJc0uz
MNwUdczx3k59fEwLMajvaTNZ5vxN5zTGmV7L7zHgMClWin4XWA2PvHrhC76dlFrCekyYWao1DWf7
4dL9CLNg4INmw2H6YWb6NkjcF4PE50b20Bgt42AEjf7d3zg+CoPkNdIMsiWr0XWaSijVw+MoGAz3
mBdJr1SIvDSn+zkyiBXdGYPx6nMrsVb6Gn4ZFmxHcsMad43vfMXXXOeLUm2JkfBsNuFZoljRyC5x
SQwyjefGBqqctQGj/fV+m9nhpvj1/cg56Ql0LazCMm5Vt7G3wuWKYTcwiMUVmYFObXCTe4GpwXTV
NaCG/M0jmAZH3T08OAU064NShNXXD9ymKbFMHnOU7lucoBy4oqt0e5GuOQT3XKzT3G2CMcG+RC5S
CTboKkXomgbxiJNIpEmRvk0LcDI/45+F7c4GNIt4FKsKqNRqZYxARNFXUZQs2XDW2Bb/+rA+FCb1
q2j92pr5a/xlQ+3gkT5ZZ2/eJqduXZWE6SBvlO00+FZSpmPP5j2RmiTE9rzkKhwrTl6bNr22CpGX
Sdgxnd36C3eTkN0HlOyVLEDdEHP6soehR1AsJVb7+lNW1a8HICDhUOhU3vUFe2S3UXF2NJ8dNbtz
KQlbjrXGxw+iq8BzX8aTKVe8egTtyH2ZgfTygtyNyZwUJbo8NmKXsaKaW+x5UfIMdYrJKfgf+Ara
CBKA9Ok/TwenCpQ/P45FjxXOVirJIYyiM4SGDZp7LrRFb1c0pm+zrhgIWQmcXnBWbB7HHvMUbHOz
sa9HOHIdIXZw1zXwocXApODjq1jUpZLgybapZ+CoCOyVRYyAXrHsIWyyC1Ze0eRSzGV8X2/LEYGd
nsmb8McIC4dywPPpVSb1efpKdRk35fQ/8LAHddjHAkVH2jfMkUIo5gzngqb8QJqbld4yUGd8US7N
lxozoE37M0geA9GaFDDMvVCNpkNjkyVfa4NY6eY7MnP7QV1XY4V0X5XUOL9r8gBKexN0RnM5ypav
lmj8fcm3s1dJIwixW7a2WOdLtsC5uz9bwurdTvj5iXfMFCEWyDNewTVz0P3QePm8qIv40nuHFWsY
z+EfAK3q/8TUq2nXdBIs1al6oeHmnpZpbLdwT06+eWRRx+YXIhYoDgK0jyB6rq5TXS02ohn1Uyhj
GW3b8xbelQq7RRfY7VGls9m8sBRi8P+ihyrDnG6az0h9DERRjzq+BvxJdacXK0W/Y6Bisl12PAi6
Gb0p9nPiHbxZCJwYtnCHTxrKuGRbKsh0KCEvJfF81N9QgWLOhCA2i5DsgsGA2kFhMa1kVizBD79Y
fcH+6Mwdto4NVIl9krFYL/xRHfoFuclwZV90kWriG3j6YK48hCnY11Br2lfpJ1gtkeBRFKxL86x5
oktxv+sQJ4DVjCs7NvcAO5/pjev8Oo3XaKhOai0GVB1jXBVAdtoXhNH+NvhpZ9/GnEiKy/5N39se
U5RVzgS+uoOs7L1QPTD6SH0VCVe7EQwm4ADuadZyvlo4NFD/bcDz0fo3OzkT+8t1FOSeJRkr0XZa
c7mtwWZ+PNs5lvbWyNyQwvs0sVNYqt7/woSMvkdsPua4GtM1iQx7ir+m4IA3SjVg5s/BERShl5gm
fdOrI+L9vHsIeFt2Gm7Gd/c1L2O1uR9rFaZ3aq/EvkjEOXRmAd9NgUstHpDjnUGULW7Z+f1nxwM2
jDe6CvPEYNw5+sngxvX1H3/gum7Sr/4THzjY0UTUDiR0dc3nYoDKMDFO4X0A9WUU8/4RKqAeXEDY
MHeKLzkaVjSyIFicVWzilZawyhklwIE/E+6c3KPTMS6vqb4WKDwTrc1UHHGjwF57GDrdZFRA6QbU
ACV/a2SJizOpZsBtU+ipR/cxUjLrdMT0e/d8RKRHYvBXXl0nz37GRfyVACDvtqZGAvEi6+C3B9Jp
xQ+Qf/iQIo8lwhNHEf5n8fLlQA8Bh5wC+WRpxUj38p+2VZk9j90Mjug83CAnSh3AfWV41a3MThun
b8V9wu6GrEdcyjENv52xwfgNmgDQein8ywA30PIg0xXCfhWcN74V/6U0sRbdw33F1lFg5kjNSrKi
+lioOIhJj323XUgB1IquEjvV/BKhYBqGaoaF30N3QnTtIM8uCRWKF55/syBzt5bHCJEHDhxgWEfL
93LGQfvJ/G8wrcrmCIfyNr67/mdSrd8XIVI0BnEOvj2w+zTmxPlBL3/Eqpz21MHeSGCg7DePzTNc
cNwfJn5Lzr2ntpdRCSK/935P63IivsuTN98qZOcb2vEbOb95CD3PhEloL+WOTnZ1J4HGeMTBA+eY
iPngvRm1jSqpoxxWOP8aCBnJ3IiSdOgpRoLoFpwtO1M/4WMqkkDHjcxgwVSj48qPZsUI7yBNRYeS
ZBE/brwEWMpfvBA53K75K0Sa9/CrWWfd/TRoe01TFgB1ysruNbPhLzZef8yH5roEPwxiGjvH4HbQ
1fcPvbyPTaU+P//y6pwtMi/cN/GLqT3jo9Am6wICNnWuhln333wDmxNE2n9fH3k+AlRB4Qh8qYp5
/NW5bohDTqaQUTYLhajJe+i8+NYpkFTaJY97UBEAgBsExiZj3J/OxJF9N1AhcULY9Vkmug81nPLx
PuWfM7XUUDe4kR1usbon0PGP55ny5GuJcKk+2FPP6P7N7m/Zv0e0SaVqvs0O6rBfCdRTNz3epPEJ
RSsCe6ghNfxSDzEqn6k3o1pQxctJhn72wziojRDB74aD95xc5Rx8D29KfQckDycsoYZDbknYiLKU
oFmZ2HTciXdJ7s06J5z34NiZ1yz1RI383rU8JXpml0DNQ5Rzem43d8nFs7ooz3xKQ9+d2HW49Ipj
/By+Di93MCtq4kyZ9Bj+Tg3IEJwK/5LNIZWOjDVmqD5uFuo1f6oAs2LDtf0ehfr3xOPvjZlgvh22
woIYkqsOMlEO6sclit+usjyObsnWnyid/FdHS/i8/9WQx+m9QXMAbhG8QAm8G8aL7SQsgYe5CE5Q
tdIMhpIYj0rZiguBzgCrdapVO7szzTaKnWWeFvfCuE4c/Y1wocE0YH5ap4RKlhPdAyqlyx0P9zOm
ZxTsObvClkXGo3EL2djVIv+sAtlcOXXckaqIESiFRo+vYU2umUf9zLv5b8Obwimc3EDYWN8Ts/NW
46sGbJ1JPgYw/qs2DkmGcIj4QrZHlZbrcwC6rAWNQCopW5+6B/gjJkzGs06RGa8UTwM9Akbgg1jB
hfIyNwzIiclt9owPuUaoeY8nA08i8Hq5eFNkTYl9A98gMQcPjHccJyQIhJ1X3NsaDq2hjZp89qzC
bAGB+kQQ9B/1OJiKl2zEj4xK8RtaYlaGdaWYDOwKKutYqFYgR7T7UH8P4Xwr9X/42XXi7m5dyxWo
5C3PEjuZgZuvNM93J+UmKacdfE5dY3CgB3QkRov3Kb1FhAn1aSsitAkdCIhLdFukGPpUdEfZrTAQ
AIrGxwIXlmq7PyGwkXzPX373MVYN4wISBP9hus9IcXcRDSaIOAy2cwQB8FDdrYSunI4pZ59xtoRB
Q9JtWXcM7lnmuFNm6s+YSROd4bulMH+jxmaCbef/ICcQmDx01IbydbpKxXXOVLDAUph9Bs+YNSB+
qbx4gwNQ2/c1+aYCZFMUkWgXfPYzxMVt9CZOWodyYurnjFZeaeQ8WoJGysPTajsGamWdma6mcsw9
chHdb71WNvsdYR6e1lE6YLiz1+DLN4HDgARKH4wlJhrMO9wcULPl7w+5gFEJwiKrdydUQjiNqO4k
L5xDfij7ObEDnobzFR3jn6RhvhbfVgKy/fGU5BBBbJAZnMVOUia4vR6WCkHyCIsNtvo0SVzy7QB2
LfpGKrqVnqmIU/k77ejFoBS6CbtuM9JYp4alvwC74yDQL13J7HtbyApm4b8BXv1+cQu5jYbnIAJa
czKgzECD3nTPWujTiAhIMTgPa6kpHMsfBSw7YnQbzr6v5JM9jrbiJ7YqX9NbTAxOflzmhorDFCB1
uaPRn8YQsbehCnfi8PQWo6c/jpgjfbvZMtv26O/syd1CSvzog/l3P7BKwM5LHtUY0U3m3SLCM7eh
KyyhEDPiPr8kYjeylQm0AlCgHxw6VXD0WICMBgmjW1utWWvO1ShM9g7XEkVV83reGApwIrNJCqXY
AaninUQhpHlOTTsfGr2142b0Y303GXhBy50xyCFv8s6lMwtNigboobyZpej3EgjFWS8qX3qHbpai
BXUjkSrv0SmA/OyhNFm/Q4P9KU4yYUmzeEXzPhGh6dwo9Nq5sRbTKFV9ObxkhqcKHxZVMTzc1J9q
t40JZ498tabigt3yGaRgMS5l9baHIWMmQt5W2+N/JwdI4GER2gFA//NIi+muPoLY5MB1HwluWAuP
mkKobgPQn+LVHPXTlqV0PRft01TD/cKxGckJupb+WVCw0nODe9eqKmEnfIqf9AYtedT0vTQpAA3k
m4jl9C1WgisgImSUEpqiiqSlxe4lNEaHtnR2PvHWHv19HJ4abz8JNIA9Cqvl3e+1tctYgtlgpW/R
WuAJ1MVu09HJZWrVGv1Uh+mddIkDYU/Nkqe1+92OEjleMClwmokQuM5IYY8Ho/9fD6exTivNxTaz
utsvayQmZvXy0bomQ/fyXrVBDN04VjAH2SiTiwO1cc6EHsLGRPjRPosAGo92OOMj8aQDA6VBqsjq
2BrvSTQT3eMWS9AK2Pe3Ua2Ob59wHn6BHGSNCFWqYxpgsnhHhvcXo9Td7D9ps18lnuT1jeJazofk
gSSDjgJ/iYgSAsSYqGfZV0s5wuojoTnxXKmbdYmYvBsdb3yzfxbUzfwoRpGNOnZ4vg01074zForI
1T4nMvDFWdR7+u7cAxU2Ys2SCUIdckNHno77R6iHqy6f9UQbAQOPGGdrVcAAgbUx7IvKG5pgLQUK
FM92R5sslylsSXitWzYu82KHy7fF08+y8D8qra4mMpOHGZsrTYPdm9Nf435eW90o3+DPLZEHmXBa
HIOy/UGNZq3yxnFcbXJHNbaA/6/IgXldnj9WtuOhSxFv4i6WYA8LFvQSDAP62hwk3beKwucekK0T
2ZyVLnI6mFBS+NWf8EZx90c+rgy8686xA8GVMVUQD9UaD3M1pueTFP6q+Kj5k99IbyZl6szmu6vu
9Dw+jQ02r6v56SHdhDFJlUik1rJpSN9msiQ/+j0+7GbZ4N6zhTk82kTYYLTPrkTy9rQmoFMjLxfD
9tKnMyQvDuwzGSWFcSsh7s/K5KZ5sPGfieFXkJOANLJFX+cdVaspWPy04s6DPKjEQ8UHfli3ilet
+xVbt75Ka0KoCKGo3iH3ZpBi0DVYSQghQD3vYat3O8tMmjLJzT+3Ccl7v7qVaNV3kLfIWcj285A+
uBZ9lrJUUp3nB3qizUOZwphfvA9xBtChKLofgmyG1q3XlzA2+H9hIPxgA5WjNd3LCRZD/quI6+I9
IkHibhSSuMvCNrVFySxhVVsFfvj9zWbBgrFSL0guUSpKZxL8BnvKICDcmn0ruzVrGMFrMaToZxUh
2g8u5aAIlrlgsbHLA+3k/uwUe5iCq+LDqQ38FVkgiHDx62HBCalfUSDkbxfZgmEfJFdslfbMOzEu
DM+BZp5QA8Jvf9fyBuATf4JCJjceXO5bS8wNTnMqoYgCC7QPDYuuo3ekh8jN4xAFHwLOJcF3fBdC
nFX3Jp/yR5aBH7AtAtyMGXYRTOGR+REQo6JxuqfE4atlAKeKR2epWtWeb/6x5JwdaGdf4swYY4NB
fvZ3wL6APKH6xRoSStqDbK7hCr4/NF05TIdV8lpjYop10n6FLcMrb8F4JYA7XPJm1mxKtRxrkjom
99b4pOKgzC8Kgq+y/08POIc6/7BpRxFuHMBrLOGWRarWOWXQR9iyCnLGuIx8kWdYYdW3awFu47U/
wP5j2/a45+1Gu9suY0MI3NvtZOt298CFhnSSXaIwdzpEgEQmjVwnBo9Db1ONc7Q+oPY0/Afyr2DU
/s0RPLyYklSvNBw6IWPcFowJF+WOKk7botJWWX+dEP0yWLxLYIX/98Zg+uPgJye2ZqVFVlmE+YBv
2IZmANLG90uyC32rSYobbrLPEe+LdOUaTcb48coSqBkqhZ6aVv7+k5v4GvjRl0iSxpNcCjY/KkZ7
BtZ97NQsjFPv6a5J9Nr2dFdTVWOpmW9EdLd4WQ3ZGHAmO+J9aEiUBhvNnW5qpNG8h2ZfXFgyqvKC
MUL1BoKeKUor+taD4/x6Z8yM+r1OOFDr2/8UcZqD71d0WYGfsomIDLqwGfafaq33ifN7Hmgu/Epf
GmS+6Tyw4HLnwGbeyhK3vKRyexHpSr766h5pqBhjegnKHadWZpBxIduNAkltm81wSbKv1O6Vb4yi
r96csYFaCGDuVKNT07hbdkyPFjfnmwcx4amqYZ2ZODKAG8qoMw3QnSotPD3BlObGhztjHKJev5jl
wku4CG0XoGxLvngdtAt2SJAnPdhzRMau/hLVAJF5+pHj4iS4fEvEEmIPIjWu6W5BMSoozJMb2b3c
B3JwdoVhAxW1o3mMJuUM35X7YJhyi1J2ihl6ZCfrh2PTE8OThDV+fQXF+qdcZb71FxBR+QX9YDuo
+v2I8FDC+1SX6J+wk+yZCru1PJlv6+ZUCvLWgohkcO3dEwSkgEcST5ofJSBMscl7w6m+OgWSK8jV
aZXKPDlWsIc+NokWgZVi9tl0i2dJsign00XWIgj6RvDUM+dj/yFejrw5clgWEy+RegdUJNvbBepe
V2/llYMRKiKMDtdrnxxXIoaqleLOQ5noLc8QTiZQvQMEb/k7usuYcG+0AhjRH7i0cS+0YwE6kxIC
UAwlEXyXHLahG0OoZNdfJfDhfgVvdXFOuOLopHAjjVp2OVLHvAetA7BcMjTkUi7qmzRQpPvLvX6P
bhAqoSkKDJo3ziPmtJ/J2qxEIUwwfGdkzs8hqcOLt2MKww81w2VKs5JrS0F8bIMLWY+dhGhtVZuW
kEuRLMbu2oK8nPweSgePl2WnQNMK++xeSs/jpu1Fb2monWvLBrhZFz+LCrb+hW5dYDsxLvBOOY9K
16ibOc3a14KkbuiVi4Z/Tank2w8qKD8hEE6ieizjNNZBHW25TSYgTh3ZFMwnH81W1C4jte0OtFrU
8m0OFkAJhnxYoYrFAxxrOyCLFrDTkHfJvjHUn+0lqypARzuEcxGJmfItMxG6EaKnZyrTF+FYCCOo
sQAb6yrXmj5DhgxluUuMstv5rTLy9H5PIXr1dAEJKjKichn/+yFQtmhAFzuTMaRIpJB7KIrFDsyO
DHO6b9lEh1/7B63xRqIWI9vDopAXHWrxbsIK5MnPO0lI2IcAt01P6u+kLF9lnS9x5sWI7HyxEdK7
Sa787xaS+DmD2vqIDJbjXvOxP1Kden8FHwOopHiQ2jVvDPqtxZ938q4pHpFE/LVVxJxcUNTf0Rwv
lPXiMdN3cxL7cFEe9vJXvY/R+u+SkefkIqjpWXGzNn1HMLZHyV+DFcQsnyP7Ta2g21/UkR52Umug
mYghyGWXsMKT6tCJVrX1j9ariBFyMbq18/ULgTOX9m3C36X5jQzFZXUT+PNF4U/7SBkDA3N9gQK8
FpMrh7Q7yrKUIxvuX53Ivaq+gT9OVmdUEIpH19IdXmpyBeNPQf98tLX1Ytq+DrhCw+dGokhgqgN9
CO+EKM0+gl/5UsN4SoDJlN3/pyEbtZzo6pIghJOoW5DLdwPePukQ3hcG/gPr8ZJ+FcEpSdDRvuOt
Obg2cSIoIItaIMJ1Tc/3pVA5u2LCT5Lr2TYep+VcQ5G1IBkEujIL1q1tvdGrfQfekiEcikCRHPdd
GwzmeMGhdxtSRPm/xatCOPU4gWhXhUROqBEC7+0ybPCSbf3MZx6sRjpg4v0EEvWCaSM0ItvVDYGv
x3musI/tuW+EYw1/4Rk5GrN+9nXQ7iLfMKB0p0r7dcBAHXnBWRpOAMv6Cxm/uL4Vdojx4peW9sWm
QRe6RVBcrg3K1NsoF/n/JV91K8wpQ+fPtJd3raTDWZ/eepqaQK6H1gymG/5ExJTziFutvTVWN+pR
KmBj8flhMR+hFTPrwY8bzkkFwgWBug1tIGrsy1VoKvRxH/bVEK+cbxWp6sIkTKMHTbgF45Rh7QHe
qMZijntso9m5/xsm5dRw2RWeY+T8g3RM0ab5dHtgIi5letp8CtlcuQqxeDbgYUxY1jriKegzmEjs
KKnrCo8gP+V6pSdtW08xjryADZp4k3GsSo2+/wqDPbuA5X98zc1UAoZPm4OO1ktxZrrVEVwUvbLg
a5VJmnA4SkYchd/CBkg6DEK5ZYjWQh7QUyok8fnlucorQ6Abut/z16X0zbnyZGhAuESIpdd4Fr+K
9LZmRPR3UjGqJYIUxAf0ljRP/NfSUdZObQL6MseScB94v5jJzo+8rzokZ6ZYzrligeZmItBia2sH
blm7nEB30HJWj7v8XY+RAKrUeIGj9nuZXv3HnSMwts0BRMDkagwITWU7L/7TVONMvq4eDpVVjrcm
jUQb2EKYkQ85xVyC4qy7ZYAlw3Pwr9nXUjtuw/q2fu7kQ38IvwbfQfORGvxAIh0a+Sg9vbsKbp3+
nE+kW5vU0G99o3qm0uzG0F3Kbp1YqpG6+qlY0laYHxSTNzT3DNAhv9cZTL99KXquBEq/5fy3sADQ
+PIEaRArfJch52FjLPvl8abR0bFxcOR1WKUstDN8F/XcdExI68pBlBbZENZLB+fTMINRVMeXoX0z
UXBwQSaNeO82cDTb/Zekcx37gWeCk0xTk/KHmOHNRRJJ24Q6baQ1O72Hxi6qs2fMFagAFPHtCywm
7Qzpycl/sfR2YwmH5CI5ZOH3LVTKT5SMBhjo/0iiwCF4e3qnVp++wVh2tFygRUv0mZRifrmpH8bi
t+bUjqBbC5I4n7bL3UltUwGhThoIFr5GwrtyhNeolFVBPQ2kXUI3Xe6sOxcHfhQ5W0xHh4KHWIfE
pLoFeSDoxS8mjoe/fmWFipZZfhqdfa3omsEOBMBhbrVKATIIPD+dNsw5hVipnJclN8mRvYiwd9rF
Wwv1O+zIvZTvSVCYrNdU0ZzRdATsTDVhWTLOw3NB3bOOjOWO0aigaYupxBiXQ0k5S/eJMibJYK1z
e3rNEiXJf/lhDM9jx01Q84n450FV3sDLJwOzAOFudTh0CGZQGfbenFkOwfEG73OJZrXX865P0OC0
Gfwy00wH2fdrDJoPtY6pPHfKx8xayCc//WxnnSQRNnrpRcidQ/Cm77lmhtKmUDxVDgbw15l1V+jn
otehyYxGFSfG8e5+S5LJQlKIoIOuyEW5RDPRUMfvDaR7k/oHKaqGvo33+8bKhIR50O405mU3cMQt
jpkbfQ73kAByKIRfFRXynE3coKn4AnhQOmtaLDOq5RcdJz7mHfAtfAbWoooqvAznq8O6X+5r6SjI
qx43YKZ/kW43auDLYkvT5VYdAujD+0p2iYpuc2xM8Z82oxAb6hvAa+TM0RElpuubHex2mlKSkgI7
ziH+ZShn660Ne+Q/bJ4tv5xtGoNx1fvBraMVxgKC9I2cQNYc7Gad3FVrI30xTETbV1TEZ4iiTyrw
IHbiIyk1SgFr89SJpezzqtjtDSycxw9wfSFe7xTBqMbKEEqOX+FW3NsIkRi2c9NtqvZJpOOoHGhj
PVjX1hAfIHLrxGvWPXr976Q4HgkAIGiB0BhNeiCxLtD22dzudFPLaweGY+jU/rx7w2wE8U8R9XL7
LNyEigq5JlE4q6YeRgD7Jz7k0AMxaw5Q4MxQDlaXw6WdtGgaNupI4sRR6XtJb11GgCJOCOMKluVC
653287KOPbdB8WdnUkizFG41wxzfSoavcaqaFM1tiFUucU9qdjJw/zjs21VyYp3yz+JAc6l2KnDu
Ax5aYdHnF42V5Fh5HOrFiEI4n/VfMN2Q8USkHu+nyU3ujmpI/K/XufyOjCjLm28FIfZQh3usJTAJ
6RYwzVJLCuDhu1kW1ngy4p2xlHIMHkH6Kvlb6J55OECdPrq8NhbSOzwhtNoQaII8txOat48f6kYb
0Jz77RG6IpXlhYwFl3xp061hFeM/rwG+C6CZehE/trIDkNKLI758IbShLpt6e3kKeNMJJWKMPyzv
GmjXtjIVRdeyxtg6lWsJXJn2Ag6d1XV8kT6njI+iIbWFPSaCtGjb6xVffVX1r+VkbMhKCJXVoU2s
9H8Yi6XvDSe8GFEjigvDS7aDOPoQXiQhj8J/LPzzAyuM+D2YLxrS2iQYRcstPDOPVYnr0lex1tlj
ZYDAdkuj4pdskr+fRQcW0yKsPxAUHGUTVAbJWMfUl/QIYbK+IGKVowH3My6+4voqC2h0uH6x0cNf
HsOIcB5aJWJ63ey1uxnGV/TyCI7DCuAZHzizSFUlzaDHEvZenS6cozAMyEsUJzk9JxQjCRc8zRmX
TN0kyEWlgEh0cpbu6U//h3eAhgEWrUzsSoqvusmg+nP/J1/jn8ZG5pCBVF+Sa5eTz9wfn5JSEjkK
5tKJtFXq/fvSUahZ1Oobrxkf+vd21yRS68lbdWIuPB7amMjdypOCqwr8F0Wi1Rgb+GII1dpLW6II
Rm+m6alepUEMcUVWxUwMujRWFQ1VDwHl4frhC0j7XfL6OmH67LlHmF+Blkt7mL9Tpjs7WQYoXoRT
94KUCkCefFyimJDWeJs89fiPm0cZkaTP//AB4niUZOPxuPqkgiGEb5jOlJre2lqJQB3DJCEyXk8b
s4xLWKRX5Qi1GWvUUvksV3+nGoMo6qsCR3FaGQuPAJYtrj7RiE1BoOlaKZZWItg8vpxPefOu7CFW
uJ7VxWNQa3tvqLNyyElLJvnECpUnsXBvUdKGASSQSz+/mS9DjIkgjCr77YAQjUIhfhO9JvFO9Y80
Myp+2q3RjfO34DpwWggSeuOPrR0Ufb7J/YufpS4Oji7iY3NcZ1aiNh+AiNAwHng+vn5m1OLJwUF1
IM5VqUo8G/SNUnf+0pl8yunx187nUOo2Wg0XxA+aq3n3EXhdzyGwsDZYdWPnO5vLdNQcTZ3ftGKA
aCxaSYgVtiKdi9y56aJbLIkmRUpTLveD9REZJJLKJoT1s79VjYFSSVIUvKwO4YKNDdDUuALXIcxc
pQbrNK4AqA5y7a9J3/TcfoVbqPt8lyMM23Ccwqao8C7yzgX6qnvQESOdGWX59z++U/HmSI8UovSG
Vj05Q3VbT+JwyHEjoWc2bDJafa7dRDkCfwC1H8GhYoFsS+rVX9cLzYK1QCtYqGyJwAMfo2LSNcjb
8sQDHVeozi7bC2dLI3oErnMFMPYwRmazcbmYRll1Qnzstl5Ox/F2nE/IdIAteuijovb07Fs6u+jZ
f45pyUJeA8rkiRWMJX63WjL4ZJedk3gMpM+FVYd96zsWUIzFxJI3uwiP8l4iOJmjWiUPqCUVgLMU
pNJRfvkU56/4pe+JTD6vY7ele4rPpyECRbOWOHnusg5kqNy13rL0XmfL073x1gLsnmxZZB1BUX87
fS0vAv14oMia6F/ckQKlSKx//lccZH6ZNHUpk/t8+gSY+ZosYf8GVAsdn0xI5dfilcShbxUNun6i
VHfcPu7X13henyEfpsn/j/xwm+ARNGX+/hefP8ub67gjMQnTbGVYrkQ2+Ard0TYQmG2Vfrzxc0QO
8RZ2ZzLUgqcCCePaSHm0UgLyCFj9h/BMuX8Rze2EI825s4YHqKNHAtSrsHlbGcEC1bu56zP3/GVh
WaiCocCJVMdqBOi6QZFKesfqF7EKU60FNtv65GSz5PnO5da1lxi7KxHCFx5/klrB+/t7fmFG5gUZ
t3eI4YxtekAAajBcfHcwjhJCbdCgw2RNpOClKWX2gvmbVXNwICHdPNDKI3gspBBmhPKNfouJ5DrD
+BAmjX8lkUuvvF3TNrt3YCxK1bfTKvmhG29r8OOC6mV9eUfjuSX8XSDzf3QLhywTViMxSmAxT0iu
yEPy+2EFQ+rhBXpNcX0Er0njhnzQRjiHC1TeGsb1JsJSs6rr6/jpzy74EfI6bfkObShO28VoSAU+
d+sdD/UBnAPQgvXrA3bW7D0tFsi6f1TNn4ATqZi60yhamwe/nkft0pyaKsIcZW7kOKqnZDPB2ixP
PKlPs3NiN1tEx5BlzcqVETqS1WNqcKkyuJbQPRtg3kEFPbPFjTjDZzIfYekcboFgiknlY3BUd6G0
HXFEiykQs+8I92FL3kYDjcb9waKdiEfcSxHtTMBWZwp+WMaqTUIq94fOUfxHCpi69dm6p4zVCBlU
Dp25MSRUN9FOPwOk/vsxsXRyCztyKYIWqsxGoFRc0CGh1KEdg1GXgrmY4cVwswKDW3QMjGaN44L6
Eq9rTsFjPLazL3xYLXfIIzFxQL00DEhiOMTzzKTZxqQDgRg4T+Xmip9q1vkBE2jPU3bNjZezouOf
QZUmV3zA+GqLzK/v8sVSo3bKhLcWnRdef4CsQCVkfw87+WI4A269j71ZkckJ71gM1E+2XToVGBM/
TaH40KEGvdAKKk9lRi84BAE5VDTBnoM4KAJa4rA6zX+T7Wk6fwHuEIN98z5QUL/tbOA783UgpNTw
Txzp+yGN+CxEP59UxraIDmU+LEcSBz+clNhZhfAVBYluFfcaxqupYzkBQIF++4J9IKGmHVxyd+8U
+TZX1hcLfeHVM4NDrB45ls7KfNda+WsQn9Lk8u6h3WsyHQ41zep7OVtafoRtK5E0GivKJPO438rJ
8Uy90Vky7pVPxLMNZhWmOVznCNxUz//5Ya1IctXiZCqRYsJJecyCstR7RXT5ftk1zXp54P4ZX1Ez
iMxxUuKaa9JoGQmBKJwF8az6GdOQx9vNbNAcRODl8YOFtjSFCV53Fz8BGMPwATc86TK9ict/iYIx
qHnk24kRfG0Hw7oZq8kBx9UdjQhQyM7/A38i/UXViDvXy0HczEcWQ7uYaAMe1zeY5XZSsKRXSFYl
N/tre1evhAgldsfPhUcW2D1q6tUejPnUtuIkziIcxPOgkVKew7wdaGjp5FGIWKqUbN6K7PWQq8fx
cbywFhFMyp8p93Xb+XsyGHkZf9PxZkdCz2ZjIM19DzGI4ltQfdAY8Fq0UaZCpOjaJiNK3VfIjF9L
llgR1pFjBNn+0Iafj1Yi/nB6xWB1hJujMHH8pilHlzyw8IaWaaRlWpmKRl1VrYQ9pbbdlHaWrzk4
KF2QOeuYYbXk+ql31liMmko4VghMwIvRRqvJZMR2eUVkJB/NFTKvLtdbb8IiiwhrNH6YQLJod4YG
2wyK5q3QJnNJSf/bIjZY3LMfM2toAe3W1EuoxuPwZ26NFWSZJoKmlXN9gDoz1zUmaD6onWd82K7s
PnoVkN2UZMleqI81xJxOCVeqfKSSyM+M7UGAfU8TMDTzLie+3JtwVOcAJ13btDwOAWnSFfYGTkru
uUkV12lJvZaRJL7bg2lkkIoZCUyWVNBCa3yFIvxbBUhM+uGDqsbog8sAYIHlqmP6jx5rSpFmZANf
fcOy66QxNlW3SR6fHRiezgyKwN0hFe/vGKNgQ/JHWcHaOqY6O/J8kjiTOW2PUHRnPNoPIkRP7Zj+
oUAnsS4RLpLs3TOjcA3xm+siKeKRbVBGiysUxc9xCCO2S5KqumCY3wPOdbikKDYUbP0yiKPnbu7/
1j6tXoBEvwaKe0c/ERtOtC/2PQTJKqzh9+xEHOtHAcycPtZCTRHUVaSpUC0bwnCKyO+v3uMa/uIS
4Kw9dqpKrWDdaQK/vkZMLyneqJh/ultKcmEP8GQ6aoTn8XIsrYwWE7BE7xKKFkuoaZOHIsKpw3Q+
LhrZfQi+xgpd5t+faxZmUa1BjS1rGBJviVe6otG1joCol069adtHVwsCVGpuawhxp64tUd4BXmz8
pJGgMOHOEHTexrsRwME59sKq73rr++kb90B2XBLs42xfkbV4OxP9XjD1hRCc4sj+avkmC4GoHyjA
7/l7Bzzv4jVVsDxqHICDKhgByV6SuNA0ogqt4CcCscn3p5PEjpcCuv+0n0OpdX9u9nv9KM3fvd1g
II7WPnBJW9+Ayo+EWj1x6e0E3bfnw483KaqgviypkP8UsshaVSlG5YuQyRgAtPiJcbJ9f/azvSNS
XZ5JXP7QzdBckTSl6QGT70155uDJEoppv7ZBuMEZiIPfvSKgRzlZNV7uKVaZ98SyopRKzRhd3KH3
jbUe6Wtib8WJYxnsaZYoPuTfGCg63ey6ocY5o8yQvPR2CSougW/2K+l08a2d6qP6BU3BpeA0MR1b
6vYehIN0NhzHk80uoNjEcTr8r+YaNhFJi8iCZHLbIbykwFzbRbylc4OE/k9savqybWAh07L0w4CS
Dn5p0JxnN5mB5qCdVwsGMr2DDNj5mnh012838UGcodV/M/yT3QL7Ig6JMn06JBA4tVH+/nz0goHe
1qFnLfmnoUYdFH19oAZxuEscxr4yBTk59oHWYHdd5eS6rV3kUfRQ1gp875rc8gyr5kSGXLuMnP+f
yK1XSHycUjjkU40q6KUsY7XGxjftWvSXj0bAvayQlOjmXoPUi571AJGIHydXLVHoGWgqgTm2vIGE
HlvXk3v8M/9et4qrQPn94Ke+PGkCoSpL2iihOFsZqlG9ClIFl6tBKDoy1/zzbYS10NlvL7f1SWM7
kg2cw1TDv0/go9IxtSDDLbSq8RA6WTBsqq0a7EENygNcL4ntGUGDNc30DVKivGQhedc3SOkssDP7
99ezGElJhGpTx4JYZazjpdPJwym7Rs1Cers1PZCMmS3EpezWK2zYdPuP9b3DVqkcPreWebx7Q5t4
2QnR4rvNlPOh5+NJbZ2XyvRDyA3DqJpdmjTFsp/jpv70PL0rmD0ivl36HwI29YBaN4GT03vq3V4B
3Lk+EAr57QtFIY3IVoZIafC33gccV2kyW7qMjxdn0i3itFLk3HY3yHmazWTM6HakIm+DORxfowtq
UVOcBJWRgY/ymjuxUekCTqXUGQHbsNc3tx7qCW1NSg5BYIe3+1xjJyPGwOrt0HJxXs19yQ+bUWYY
YGjZn1yvzJEO+fWl3S1wEYJCxGtRjY8ok1rjhP343KCggtltdzB9p/9p34hhL6bCDsxd7sq2gzWQ
h0Os4EeU+YGd3nM096MJPK2ZhFZoXaj2fet7rL75xsC5v5ArpxaZSNHDJp86prnVjgmitAjJ+B/+
X5T42SqT9CZT50WnP4t0Lw+XdP9U/g1W/hXz+vRrzrjHNwOzYz2xe8GyGlL/HLJt/P/gNZgITR3/
YGuyf4XRvCvX476Yis6aeYM9GHb1ZPgiqEdiDASBIH7Lyx+V9U7lK5ukL51mHbjxgtlgOYreltIP
2F/1X+5hB4vy2ShVK9NttfYaXZ+2uNgIXNUm92nrNFnsD8Bdidhit+5oxAETfHc50lvmQ5XyZj7/
utenXr3DEbBbssKe9MQEDWT4UqzZvgqYol2vAK7ZcG9tNGThp5peMPTgtGaegMK7TbvzxaTQOnSE
BvLAidpcgSMstOHtumA6s4UMNBWkfeDaupZvfH9yVLEYAIHx85xGZqa72xv+H7sEOAYz7u/FRHDQ
WAvC7cmlXrWAKUIsqmIboEnyqivi+gtm+0Y+6xXTdugkTBaXjuaXU5SoFTY0dfQo6nWsOFT0Q1d+
acsWzElj9GNufYHwxZ+dvoMKo/o7RW+i0QR8mCyN8kTg39yHyO2/uvPMjdtFvA0AcOfg37PB3tJl
X4iLM962FxMl1pUUUa4ixM4z7ASoaFB0VMPt4lIzlMyuGbGr43tEuOCGFEqhEEhqjlF7wzG1A5UH
f/Sag5/bRKOdv2JFp0ZjrdPtqXbOytZum8bChMKExjRDiDwLiusYnbAihaaRzYtX15mJxvyJMd9I
OY35J4sV5Ns4IQ4kWbhI4ozH17ne5AXQN6UUpZvRWK7x50YpiuV8LUIPbL7EG5Q7oBHw51iCr3Dc
oZ9RxF2KXy2FSKZ7H9Lpf4UF+jI0xtjrpThqGSEToavM4cUdNsLMLdsmJMbIsXs2uy7mEaWdK9HR
zqurOOfybm6OYMZSH0wk5BOFS9X+Cyg4iIwjK0nOoDzOb85sBjoCZvYTAALxA3CSjxbk+FmptgrD
/CxJvXIIh4Y9lbzPghsVe6xDQxpyRfc14/xmxEc5JmbAj13T5TjUY6pQNSNzEC152+jV66wYXaGT
wovVoRjJwr00cm7MeCmkn5tlre5+BUfiX1OalPzX+G6RoYakzNERCVDx5lu0dqRrO+VGcSswGBvF
nT6p7xQu4hhtppoxZIgAZBkR19HLClkrFdJecD/nLjO4QOd5vZW/Nuu8WEka/4Aeo11TRYvyIFCd
IQOrBJ7IfKx7mx6SIjb8zUUToy0hjLNk6zahwcrYqKqhIetmSpwPK89UK4XGqPohK1W4161Uspse
8wJvHxAm0pgqtUPU2NuzIW10HKeubhIuoXwz8IzjqgRRpmaFtsQn9rzvN31S9jWqOlY3QX6uupSo
9v8SjKeEnFAAyHOkwphEYWbgDd67JJkkAXs0Pvm5mPW1YYiZ7bjf9Sz3Rzl2I+UrclNmJKlxW23Y
Asg1myoj7jOszZyV+VZFwhbr1tO/cpHZqZYpOPNDUXdE5bdfRYuaA7UbPoFtXnEjIjGqzlQRRLfy
GaQ0FKi5boBBGP1H0hG3OaM97iCCjP92bY/NQaMZwqHzQo4Kf5st5L1yXprywZMZhw3HS4hhb0Tt
C2GgGzzYH5rKANBhu25XjVjYwbL43+SfSFSI81fqk1v0IBtkjGfiWe/rvo37q7FDfI2RGKd+pzMP
Js+towIM+ewKp5ejwljBlx1rH2eC3ow2frb3EZ/jhas9XYic2p965ctDWS7bWYMb++lusIp2OJOM
Qlz8onJ4Vx1Kf3KgHlcYo4i3ZO2U8IZN9ju/LRuFywHWqlEXV3wJirYxtCPwS0ihTKHk3HmG8klN
ADdzzSD89aFLteLzr0QOND2uPMFcR3MYOPLXsfE5FeJaw6CHAMGMqJ1h6ZWVsvKR6dhO7DwmSVl6
bNauUuFxgUQ/TSbJNMmElRg5ML+RoF85nxO1AVYmb/MyYEjcs4WKOqRXk2VMYDd6OJyvfzmtidO3
fWwixAWm2pMXrp0IaM2lQa4FcuJwaOiORc8kHNOzzqA/g+S06D/ILujNqHgpQYobO2E2P8F6NShd
abld/zz+tHUfxC1Q1TSdK/McaFiR4x8RZOXLeHjTcimt3vXWKTi2XDaRfry1No9YL28wKu3nDzQl
7mm43KC59mi8IbJY5JhzeDKZ7h1K3ywiPiYm+n44mzl/7tXsnMj3fOylz/EbLn9VUYlEcOmsykuk
nF5H4Z69rd1hroUQhgHWiIVfifqULURuEb4O2t7Ir98sjEmFmnofRHBbs6RwT/3FWhR08o3ZWJSy
E/EpxUb0CnbhfJkDjGhAeEu1NcHBactr4Uh3QGxQsbPBlPVNsAUup5/ejUjsOkD+VJxwXE+mGr33
rp4Z2VdOTF3fQ+w5V+ANwlb/48vFjIfsLmlblUSUM5b5Q52u+euXbWjpWdrAYOhKjUP3eM7VlY1w
FiPEHEepJvq7CagYWVqcILRSP27XrXrxPbIYaJVh9UvIBuQndhDWUXnqw3b76Uw3yRFBe99zHE+E
zHv5x77w3c+1Tp6o4Jw75Tt3RMgvtF8ImaZf1sXIo6yLP/H6r3FQEjd7l8s38pUZUjuIn5blGONP
+5eRfkaRWSVXyOYye81dTn/lOgO2gjNrnwoVB8n2DXSPLEy2hWX9CeWmQMM0DyIVtZcPq2NOD4TD
++PJeoxjR7Eb80sMsl29BooWIoztNJUDuWi8udsFKKWO4IYpOLdjXY9HCoRsGVDEuUnv41a0QaQb
+HBhmbYiREDA7QnCjoV7Jm+UB3OJ8Bgn7trVDUrdrIHF7Mc0zeTyQeaD05h+1IeZ94PDENJTj82k
8fK94Dr2krROQVWpOJ1a2MfY9MiHg9YfICg7u26TK3DQkIyPMXa765kAqUfwkeD962dKH9Nu+6t2
/vxEo3F3TYmIKRBFahnEUJ+OhsdKXw38fvZEubNtEfMqu3JKK7YF+GqIfp/gkhVFKS7vm3CWhcVT
deCt4uuC4Xcl4F1FQoh76OdgUK4EvxXCUzBbe+XfB11PCi+f67NypaaX8Q1nlfD5yS6PGzZGWvPG
bah+01NcnijrpbB5v+W3/sGp91XKDqU0GxiDWqMzri1/5S5/JeAQWfixeT/k78N8nCSBw1ZfY17B
XrPyxsgoiD4Wg7fzp0vDRVN1NxJ4NMU0w09NPfgp2jfSiZefaf8kYZYNhO1KkKoRDgZHpwHZVMtW
dkkBee7Q1boL8pAKlOfXm33VFMpumCwbO1BtNkvPSlkwOTi6tjiyGght+qWzAtVuhlnPU60Ch7Vs
FvsrujAojFNfsiqcShvE2q/hp44fynHXY+9uVudTz8wDaR/TE7m/85RSR4ngXhB8omLQFrAYt4wQ
H6P+tVH1y9brIR96UYuFJB1ksYa/2qg9qdYGWTHDUSQDs0kRVKKbtWrVXwL1AC/ZzaU2j0wkKgs9
tsz+MmFjVblls9jq0WJxL/DWrSsUDeA2ph3CsP1QS3MNGApIfXc7HwWSEo8MfO99V2gIJXl89/pF
oxsqZFSA41f26ABA+ZLIUrLq8sJ31pHDvuxwAyzqZyaA2udOhl9HrPmFmohVZMi2mev37uOKojW9
n+r0bWyOuurNbcX1rDc4N4Lx+Nz+0ygaWbTdHNad8Y8oLRRgI//bcXLMJNuOBDXt7moAefkYTelf
3WXpq/EXRzWTW5Js3CVJMCyujojqFVB+d13FL9q+Wg5baTdTHSFMSfOX+ZxOJ24Sp13D7Xf4zBWH
Ma5P8GVFgrbrZ3DwjDl2E2p7fo8v4hOgMb+MDHAdFInbJCnOdxluTYDPtC3/iroiPTazIFZ+fZ6Y
3pY5NsmhbwD6oU4K4lKzkGAnUvyIqIvQAtxScuCxVEY7FQObtxAPcJB21pbg+gab1yvGccb1AwAo
Eynm0VyvuPWk998IXTouSTz7aATH2TOBVZEPiZ+BPObIrdJ48O+whPJEL/V+0uAXQWMNT0rFNl7n
tbC2o0LnUEZGGozhhLSW1Y26JGs42bmA9+jZM6lFoaWu7g6cnwXLj9OWPQ8Ep5zvET+r+BhAJAux
SuE/7T1YEkOgnXy+BYYpU0Pbtm5A1czSemLa3BpN6KNvqfBevAU8p3ap13IwHJU4jiZdKLXOeXK3
ShI2orulBlkdHuIcjXY/jSaSNdKEHSM8XT64NGSdKLpQ3Is3a8Eo7gZoBh8a2HeW1TM717ITymqL
uNbaxSE6EP0qA+yC6EuXV5akM64pciLzkZTwf6RFv0pEakS1bSb0xM9dHKAt3rn+Q77LveldT16j
fEZ1tiEPMWoseVsZqh5uwDqNxj7tlo9xijN+IXrxd4JW6V/cBVxSo+5uaRsjFi0Gp3ShywhnCDvT
oUK8AJYXRinF8QWnqln0zCIgCozG96XfoLVZh3WYDPcjPT3csGN4h0db4idFHRk1C83Q1lZJ3ukK
7VCG9W5N3xnyFTVljPFUFczro/iYPP5lNxjxl2pOSquU5QNkGSfufVbFhpho0wlcLscFqd8FZx6A
/rggFkjMGJgO1IGCGzeyp1AJFR6n6fpjFb3uXKg+0Yb/BYsJ6ADv1CyIpk3E3lJKtdUT2LhiqDsp
YlJvL3laCXHlV+BVagBAIO5f1MPSos5ul6VXaPERoAQyDV8cTl0aU2WfaKmm8S2JiJsiGR0Y5F4u
HtRrrL72HiY1cYDIM2QbQwsUo9VTfV8Pb+BRc0X0G3yS/SfB8HxW1xav+5iHGf1COlOUctvIiUVu
cvzECMq4BKYoszWr8BS8XnxbUyRnaeVu6hm895Ks+XA1DIDwQA2953V6R+8V++EnU9CUKxncqv8x
Oab07hlntyTEygkH9m/7nfv5q4F1QLUo2OHNXd9QInj5JVUFlNHgQ/JFhWJAA7dt0UEPaKUtXK4q
fpzBmSOrc5C8+bsTz0SWMFaUnpsKZp9TS9IU76q7S6LBisFZC6otmLnpcuBLnZuP4AvLXUH15Ggn
u75HK0qBhXsfoOzrxgxw/GP817rJ07lJjxP3uUFnNrbUZ7Y61JnOzObXEfaEvVeWsnbPtkXgRcju
VHrBA+nWgUXQarAbQjiBVtVlEN0BW/WlXGvBCizQTr42XpJStaS9Zlb67qJzOBjea9OZ1+/FTk54
p7LAwgpp23N79LlSbYB054+zhahxLyOzPDRM8lgInn+ffv5I6KoP12C97m7mLutgg8BsurCMUUq8
7ROHnIn1yU0geuPNfOD5SI2Wk2IMy/o0Z43qfHIIbcz0PTFE4tgNQrcBA7u7l0PbXntbUCqYpE4S
G4DGVO6LEAQb63knABeGIZ3N7MsITjr0Mm5PUipgh9IVw4MaYCymFAVkAwwRr04fKR/YJc/wUx0G
3aY2ar73u1mMIIL2d4+1d+lfj1MgWWtj0EfVoOYb9pw1kSgesufDt9zROso4zvgjDaSOpn0KD0l7
7QdIpnOahzSf1fuG8++XM6OjFQOeRXzZfnedhiMxgpDuwcVTtCIXCa9rq0lOrrtHwUBZ1v5WOjXa
CTUbtmbzktu2eLfTafCJOP48hBFwGAlw8OkZYWdcjjnuJdxIiiTfFv553DkDCU3IwzO0XUke0E74
fU+g0Nu6E0vn+PHc8Cov3R2RcjIjKLbmt6JpIZUJBcjPzjdW9upwxp54Cvvu7ciXwOBK2j4jaIoI
KU8bgImopPgcJC8YpRT+oLVmhkNrpq/Xcl/2wMfW2pBh1AeHw6LJOo0QJSxdYtl/uKPgHfiRlj5w
F9O8RMF2nhJGe7zv7Q7K1DoNoKhOPAvm4th5XJYSUMK+4hK+KUtP9IzY4/Rq7/d6ibjvejgGc3gz
CDNf/aA/Bjrbmq0fSQOvkQFBKnwss8aTSm4pHw5xa+ozYZf9cBvRA/q3F/tSf76MDhEAtMVkkuez
88oOwSCDNKZtlWL2q9+3gEQOscQNWTI+JLvUWPO9I6ZoxJWy2xrlW8b1ERRRBmT4x/OSnVC3Vu8i
Yt/SQgF3QOasc4bDVkAunvzT4HFtO9MNbDJPob4hvCp5kngicJ5MlxV9/GLQ9ofcwB3LMFg3pjc3
wkNSWbf64J5fxDzdCS7fkquEU3ytuKXh3+4WUdtow8MmFp58h/DWB1dDpeZ5b7OwtliS6j+HkCux
vB1VK5+evWl7UwdNbCrZrwbYJ03jjLAuM1rQd57+uAmgRP/HiTXseMHHCmVnTGmxNhhUc8clfAy0
CGk2uXeJXeD7fstMuHh/dmI4M8W78lY0PH85PUneFMmnqR8rONJPLH26sOi1AlNQyKHZGivO8VoD
pir/5ZaIHcFd/MVFk73wQL28nWWeQlSBrNcstdj3OQCTyDcjcgX13K622jkMDCbiAKsa5DuncfVh
EwYpUBystCCud/4bgJPEmyqVAJ/OWSvacLggqJ7ILz0UyDEH8+KlfbnVpKbJqlqf0fX1b8+cQN2x
GclEbefz23M7wsXi+wuJWLs8mV/Wnjgvh//wqAmyF7LnGe3WHSSKjqjpfmTLRso5ID+bxu0zAOKi
KZmX5j3QKU9jSHpYksWcPMx/6pjcY3YjiJ/yb5zA0PBoOliG13+QEqyJDw49bMRPxptubmT9Ag/J
RS4lE4GdoFBgCDFfvbfgrBCZa0IBZNvshqehfp1O/3CN4nWeLbWnKd2he5xQp5I6tGgjqGHrO+oy
S73cP5qYnF5Ntn+89a3rN05B8+XtYlKFNz1HTPcPWDvkheZMnt1xeWOrAxswe9LYxHcL9w9x8xpS
FH9fFHCxljTX3hNYh9jAWgDXH4XSryUZLaHFWfI/OBigyTeIU2cqURP3zb9qMh1igz4l4cTtKqGV
hLfKh+StxlmZW1nBRmAcauwk5TVxgJOtB3wq9XwSXjdwfs1jvhc/Clyhzsfg0aWukAeVsJF8hcB7
pCFLUOgqGcsAtBiAGPEfObASqJ6FpEZ6keRtqKp04nr6WcwVbQAlRR3tl6D5g6agS0tPzYnda64V
jx2jeiLRjd4ooxEIpRbQSc+NMWoGlaIGBTGXheywdWsF6RrKFt22EcskDdkFfOOEqwfiY6iDT9Kw
L58kEtQJdso/7EgJNf6ZG6mdByAzyRhY0x3x2RVLW21B2eegrEdRB6zFoGjKm2ih44tw67uRqVPH
3AtyOQdnp43IRQdXq6dMjwjyKcR2WGTpn2+Y0GBREUr8RUbKX5Zqal2lNX/tpYMCKjYpi/+djWbl
K8Zh5pe6QQeib95rzMa9/4Sj/nuiABwLKMjHoTIqO9vJLQCzz74jnwIc8Ue3PJS8tMmqfpiGlRhf
v/up62+PKbLVxuursixY9gr1o1r3QLVNIjkwW+Fbfjr2iuVxTx2eyM32Q421J9pzw/C5eTGVf+tX
z++yWDDN6sdDq6hQnYcVwinKtcI0ggBkwc8JVYSLrnhDM5DnQlY4k2deD1MOhCLmHBNfOCAdjVxZ
D3mdk1AFY6gFmm719VXO/qU+FwUIfIQc2W6pebrixWqnk5aBxZnTLz87CSPw7rFiFlZANOeLTmRF
H5aV6TZon3gaNIDMyfIaj5STMAAF5cZXlR7d72gHTFh2FrLPR6rB+X2a+gS+SY/9HhcQP/K8lGyp
dQhUN8cYhjc/pPhYl6cHW1q1mKdIiq4olT23cwYMxEI03V6AYvIfKBNaZzi+jJyFEicI6N5qQYOS
b9VotmbR1JLgq6LVFt0QfS6mWIo1iECIQXLhOEsl8t78uqsmSVn8JVmilMkOmQFzc8r/Oag9gowc
lI8X0suRnqS1SMkDBTFcPxCRAT45XJlCn5JrfU7LtAO4uoDMpsVvcLJ4nkaRwlN4JvMkg3OWYPZb
PEQZPay/1KPBTdudi6pGlGUpbRe4mzbbOT1YHJOi7/1fzlKzL7qL9GvSEm6jzgcypxAdUn8JscWb
6rC01729LR9cx519nvQIsAp9nG/xVc0Tardn6GAyl6eMsMhHoz2Z4hERg/p9x7q+GkbOvm6ad4Dd
I1eE8mq4HaC37YIZIAOooSHsYOzCGWkJKn23IAYipJ+2W6E2EavMgLmH6shsPEPUX2NHMpHxa7Ns
FUkGYtxIDXyHUfJ4KyJLN07zQgqSd7dxibCfc1XoR5HH40mHxB8yg287Yeo4Gdntgr8SJ/eywSjw
az3AQHDl1j1nm46VNB/6SPpDy/csnnOVtfI1o331ihR1mHUDh6vZHuSUqdiOMMPLaHqj1HvMOWQe
mclXc8oBgvo027qdbY0Lu8wdaPN7DD/eSVG570lEymdH6E59acq2NBfk7cY/nTvCYmH6Iv+nwfnJ
fQn9AfIwGwpM6BDarO/K3+g0Fl084NsP6MVEPQJtgE2/Hfco2i/NNoUAaTsKj6vMaP08KoURmaan
F50QiAPEopKig7Xe/mydhMVwxjzFKcyhowHGyN79zwd6pJRkpd3gyKhffMBBG04Ukj82c6TZeE25
YIhlI5KbB3accPy2bhNDo/+zAL3B/2IwcoAiKI/UckJDYr/ZGb3TMI7p972paxp4P11SSA+m6yTk
79aYq3U1NzSD0Lv4QEPpBnmPlpzcdolTZ2obq2ZW4Dr/IEKGQdP7aGlamfF+8SA6wzMTH/Peri+O
PPlCRiX2bZYgNSclua8j9uF5MuKlPBfBM25/KEk3LcNJAPpWEK8AAuhYKEjv4f5QajgbEOEEqNU4
qfxh9qAhdn1LWNkVgDtTifBn9lDJd1CmGIeO/+Y4YkJXruegxGImVegEiemDvLcqYVGeyEKMWRFp
5qzFsC2dXY1p64HWJtINbsh8kwiCZXRXfgsTT6a/W/yYMR6gzox1/8Sk7HF9qIu/tDYAqZ1vZUuz
VlWRYz32eL4YGp5oUjtEUlPFVndljDGkX37FGYdUe1KIt0m2oj3l4x6OEH4kSvgxx7okb9TOkJue
gwVyfrC+CM3G/gYTJdNaDo8CrzIUiqTcDAMKJ2sgqha13xUUugAzUK+Qz7h8NZHGvmXEpTeR3LFF
2PCpyWNKJ9Ccg6pMP/fI9UG7rmhamPaUUcNEsqLrPRVFy7dpNhh2B2TC8r9kAckFEyqq9JBNoE+Q
wv4l0nN/w0RHq5yc0CmQsNdI1iMcQdXBUwOx2lRIro88aC9mnlcNMllPkcQ1WeVpAv3J1s1Gsf7J
IdBWMIUYgz5wkkgQWthR3gr4AYrngvqY0DA1SadyeysAdZV1TwosCwSUbxIRC6bcfQ2K6r+huWx3
CBU8x3cV2KOVtbIOoAAuiGSK1t6f+wCkihTuUBgfgmZMPawTPekHCPawec7tMFQrS8pGq1LL0NYx
SRi5xKeRyaRsOTdZl0j4aYHOvgetnxlYH6RAU+nKAJxp2eQqIiGjyvXrs1N6K5hRzA+3mqrcw9rD
MH867sWBlm5E5VrGoHWtyPGXN9nzCvVpi+vRfJRwLOXNmNGG75QhvudpKYQb9cT9uWjRMBYtuVNO
fUFRxdxUB8qOb3z7EX0O//LxkJU4jnzABDeSvZNmJYa5EzVQdgO5EZ0xuI1FF+eGC8VukRrequcD
GZAOfLzj5wMKlN4gtMIbRuJFevQzOITKIWvLa/+gimSzdAPcDuQhCcFhlYav0sMBTYAMW19EYNHH
il6GFz5nfFRgivbG+vzl04edi9sw2t/8Gx1n0J6Igilpf9GYM1kEhbG9A0uU4MccmCeIftQCIF7l
cm/nuEyn6tWqqwGN3qUMWLqxwYVQyDaJqV9ul9ucW0nvP8nfgcTzJgycFCOX/p2t6GWRlabWez3g
5qiFbJ7gH4JI/C7erwmZ7FPy2ZeLiot5jv6nD4CSqkmOVAPNyu5jix4JguE9vtNHK0hGFcTJG22z
ZWikigN4LJFFkce+YVzifeYGJ8Y4vH4KY8SCZvM+NyrZd7wW1ZN4MO8Z9OVsjLJGLdnkivRdrdDY
zx2/TzxEt6IQ9Ejsu/N83gIBVJV+kUlf++yp8o2PZx5aU7DFa7RirZYINRJK8pUNw18+qZ6wu0V7
iHMfSYsC4rpVgJiYjbUqrolRGveru8BJhWiA2mH3gPuPalqO940yPzRAN3+JvnqhCcy3HgQnbavb
pjM4V50dNMC7lAR6QpJnT7cWV3RcIhJfE/yjeKV2FiLGsG+ThLdU3QD8wpr30xmaxH2/wt18ORKR
GAIXuuta9kgEZeIDy2G9PTVM78zknc3pXIIuqTPMRxf7Uw+uYlbbT8c1lDddS3naJSjIM/CoFoIl
EDdqupp16xLU6crDRIEmJ5YZISjGzlLsAiFmdgzYdT6dg7L41UsHyH03MLouAkvQQrkCkbgcw8Et
tQc2Uvy0U5VbehVVDjY77ZWL6fK8+GE64ZZoDVTTdcqVGo9ztTt0qDFpyluYOefuOyY69tbdq2IS
aCjZUPbd02wy12yA0cUenurGkS3M2FDQ19AFnNsSfA/OAD4kA5iAuA/fd2NFLc/UYqkcBES6r7Yi
RCdWhBQchBeBNMVTsTXctEijRJ0Koqp+9TanYQN5V14eKVW3awT+8CH0kDznQPiSmOdMPVUKyIYe
BxYSmPsVQTQD1wyyRtQlp5jnLxwkq+TuBODm8zgcxPwKuI2IV9xIEA8Q34Crajm5F7TJw+YmnRVp
lgva/luWSoYOwB44bQsGXk8jA6UEOHQZtzjaqLeaBtJbulipkm47GsW54/Oa9JrPdMc91cNhUN03
97Y7CfHuwKoLudQdL456EypqjKZPWXwG8VlvR6mF+l9JEv6+eGKpcwCnjmgiuDsd55OPw+8TkG8a
vBTgdGFiQMtpLLvxLK2LfrgFmlgnX6YiNeWNXOuwZ2LjPHXKN60Jrf0WHHKjwEtyDCtBkOAjQfhQ
W2+Ch0px23sQpxoZMPng0kp+7wJSprST1/bwKKxRckeVYbh6bM+ohZPxtSImRTFDcAxQCrMSQQaB
YTu1RriqCZiHGlRgIkmpV0AMb2qSxgafzapEK46hyhqqQrAEZPVYyQ0iWoqrAceLsy1Ea1aH4rFn
kbAgIg/CRewuSvCFm+Q2AewM1hH5jKApJfA4Wfx5jXrZVBgshu6FUM1mOJYfIDiCjclCAyyFtmty
tLwU6MT092o8/6ena3w+mlxnZIAfM4nvOy9MXwVbd3aGuzmHDFhFFxyFMMZtSQoJOsX22YUbiX3Q
5deaN7xd7+iq0eDTbt1nTGoNagAKybebBNb/A6XpOE24GcUuMBsKuhI8qUdJ72EdxjxN8LKHAqZB
F3lM9rXZXQKOR3X8Qi3bRDUXUVlaJy9yVfMyHJ88wWTlfmaXQNRnWMK/hPMD+4bkm3CjnncdCMFM
U0LaooujA28Q16QQ4Y/PHpedIrbom4S9fXp60n/uK6ZebN8l6lIKETlVV+v8oqeIfVQ2tjJrMiFQ
3bcBda/9x21szMYOHncoDTWk11Ipr83Q2Mu+zswRMMFZ1+CXuhZA6dkwPXzowzQqoxkSB5EjDD3b
tfDg+VCLUrP6KUinz4Emsw+7oOH7+H2HLPFR4mdqOXczdznQfUwpKGOmKFxLOC50zY+jkz72cp7Z
g3m3y4GCFLO1D/sy13JN5wrS5zSRDRUkbpUt0Gn+cHSj/NGVvIRdZgZqCJpXum7ot70N2U3ns8TG
UwlpjRAXliq809UDv6M3bD7o0DRbUcSGES21KtcV4vXVzM9bnvCVhFN+8+lO/0qH7FV8HIweLdqn
rxnIVK97tvhaYEPb4rmx2ljUMjeobMCP5TFx4xoFPzpC6zoJ0tMrNAklQGv9L2W6RIlEGSGWg9B4
723wfrqvy8sPKxudt7Z2EEQ9vV4P4vdZUrz29sCBycv/qLJO0/PSgfeK9wuZcH7PDJSZ4i13lF1N
vFwh+TOJrFNduT/T01a6ysNc29Id393/ciONpa+BLB6fXLRe31SC89pm3ecwJukKuZsKGWSv/pjh
wqjIN5yMH8F1ecpMq4iTHi77Vh844fKsrAWHvCGtw1wAXvUfXcoW6HeDdyW6Ahe0sRUD9hVN308m
+HjtgeraU6I7B1RCSVQTZ4yYdTJF8ZFOlKFhRMxjuKyBsY81cbGk9Bx3+m0wc8nZe0zDu6IbIefa
uXseVHUSHu0q9dSlHygkqVBnr/stTcbZHSpQGwYjRZwGr/5n2PUXuCKuYllwC6iL4lra2KZQbHKG
A5BZoPh72TBghl3JVtJLZczCzkMRVViOcI4u9ofeymN6iIwA9qLzvgwKFdLy8UUnG5aBIPBeWSKf
lmMv+yV2nDN4udmzFfmtgDkje4YFmn64r+DsakDlwxqDugU6lvxjHS2cPHclr6IGUKQd0W8NpVDX
U02qyR6n8671ZESzoHWMOQqKxiZCQcGGZOn3ylHQTKxC8b6mmSK9YjerjMvyxt0B4g+StUF60kF+
0lylVes2wsQfTgwIprHcyNfa3uSDdjFQ2o/Bap8j4wvl+ESAJivKSdCie1jPUA5gV/9xU95kJaUt
0t/zt0FIbDvDOtuY6VJ5IATwEv8HONVdG6tIlM7UJTLh0d/pzv1Mos9cgMbNcgc0n2T4ACo2q4uy
V1Vs2woPnpfiEpYIXgHTrN5T3O2l/+ggl1cJ4GYxSegz/8n5iy+Id7NWY+AjDNh3FpekE8twBCOS
+fJPH3WL9WkJsB4pHP7HC/QuipvHy9H4xF95/zpQNNgKfyoZX4lx7480o5XJRpAridehTrpHM0lB
ChvCyUp00cigV9CVx3N6zX4vg8nEd67YQiDg6fAS0qMZyh5vToFLp+c2WyBg7NxWA20YNiM0VXOE
rZtm3fkJbTu3EPK7OKJ4akVhoYSiMheJLfDOrcJLjl5WLRbcjHT0lMhKJKAvtBRTps0r1gELgyJt
ApDdYnkvrZmZbAdUWN3LmrsKptUhO2iYgH2FrSMTQprqsxFCswOm3sEgOxWaHk5/Z6/oOQk3Pfpn
LqCCwmTe4+un4swfTkk+JiZ6Xgdkx4sdRc2k8echavprb1NjmHSrk2QC1Njkcq6rzmsXEpVNNtbw
k0oKzYQ5gHq1GHLXWn+OUEL5DfAU3Lu0+4cjjbu9guiIdtV6sYbHXlHI1et6xQJ8RRrhtm+m1/QB
AykKZjQUUmZtWtfhBIXeCUQNr6nFBZYjxqLEMRKKVN5HZWneywUnxX2Esf19B1tH/jjNZU/0+2JF
d6QbI0LT1yMXljtxTz5SdrjxvwaUeivJ7+23cxUEzILtLwO5a/+Dp+y1vPD2sSMNzchcQV/9fuTQ
h2rJcPPNH9rrNBCiXS6K2XBvca03BAqM2sxWjg4MOs/zaIbaXPNUhbjTBc9AEQQTVF57RTA3PGSB
4IlcIvX3ORc7EEN5HzJdSWjq5NIHYhI0Bm6WlrtVuyksqveaARD8welFC8q5p9KnELtzM7E3HwwL
F6nbROnrox5g9XRKXDry9Ot2VlGcLgWni/zfBD5mDfXYzccPdzXyQnKjHWD/uoyCjC6fUkWjAwqv
/Wx8S3oW5I4wupaGrFPB/c4HXnefyZGiGFx348sMOR9V9TKe/GTcAJXQzevI+6uqKzYV3dWEeE5v
IgBpItknavzKARP5lDU9OQzmbdLi3ed30hj2HR8nDhxyKAHivzMNBg/5lZIfzbet0gNyLcbJ5orK
AJqSb4EtSNGErkHa+jp8AdOFCHeiUk5K+X3kGlZA0yKaNGXv3xwlYX3Eu9hgbFqKMrOF+ApKIsur
7aYRyLrnQ/+MYMAu6Wou1urQtiiRAMG4niKMMT5GkQR+9ifwaYPu4dj5dnnmJo9jwCeKWRJh1dwG
vC1Fsf9uvuiToviz/B32WC9iizEJpKnZlVCwFZv7P1iBeEnnplU06iwzYoRuvZli4VsPmr5xeZKg
gwujOwtmq3mGYgFUdRB1H0ZUC2k+Y4VixfEmSKXCeZj+e5MLjVPFAo9GGHqmGYDURAgiE8XAjkc6
McRjB17e1Rq1S3MOvS4lo6FbM9ejs3qGFuzUowGM41k6XOe1FQDJ9ryVKwwD4PGn+Mhav/8ZeSt9
h+XIYrYGiH4gMMRlAAi/Dsu3l0bAtGgKbsUltTvjRBvElR+kY12IBY2A501KY4C5jRIAlvtzR7xt
Mo8qW1eEr3FDTnNp1vDqfRX9CgjB6huF9z8qbSPs84tuocuPSHWhVUZ5DuvaOUOYSU4xYU9Re6lq
IAWuekY3gL9tqUqGz5IkgVmkmq3xTpfsq2ewLtOop8PRAhjbN3cK9gcOHqeeNXdVTJN45G2KVvK6
mgSQF+H7qZNkenmio1m4jN3W3nLdImb2HAjIi5t5AlecgeqdLI2IG+ZuhUCqm/6ukst1/Iflfd0s
wRHEgoLMxtHbKPldr/hCNFCE++5wYhB58iaaLVUmMR1vMKt5AFnwRDSjO9dLwUDgupB8Eh7FS9Id
QlyBNi3Tibnv45KY5r2qIwUFhKo2E/5Tmo/yk0HH+m/+81c+eW7T9HSinmGEP2L91WajXdwVkc/T
22+r5N6sDV1F6EbQ9rG3vt/Ar/DWxGb2Sor7YcQOHj5S+Fuy/7cP5qBD6tORjeU2YvvTFPP7A936
wgEe0E6cnqtaJn1+XCjuyT5vZKq070jNc2UzgR/FIOuUNlX23tNAbW3N4S53nKr2NDIpQFNkVfLr
A3GNcQ4Ss5bekkstd5tgHkZiRcCrea5sxC45q0lj8uE3dL1gNVlyjffnck1YOF55ZRz7TZEqPfec
NDg981a593N/+/UTFBzbUaoF+05L68B9fpaExqq6H1tu6LIg4iH9+9BUnDhyIypbShHCKHmKYFYp
xSMD5j3oG50ydBh4FO7E8OijTmg9g7OsFXo3nskVAf0AYopoO/E/ZcdbkF21YASVDLdEYwM/gyH5
jjbdS/Bx1M0UAzDBsz6CvuWkbyhRx+61GRvt1APHh+ac2HXDXgQy0E+MVzC/vlkbxk+QvkMTGS8k
X0HrIeh6k70iXqZ45yjINYbPFSSJ0s5EzA/c7gQlDIHEGt/yQMZxO+bLi9GLfDNMkfpi/O+VceQP
3DreRKwAetj3qkQtZXgd4+0ByM5jhu/oa+GOasxY/GCbmTe0z481TBRdojFGLVQbcFu5hzRIyFfz
XjU5bnuG+nWcm8x+5jBebQcLbW86341hQOSsea6Dr64urCm/6k2mrL1q6wc7/olAYEiKHNb4Xqke
JTQT5kRPV+5HQtXqn+xq9LmGQQNAOdGEiU0CmfH6cJTzs/boZ1wFAjhS1lq0vOLjFH6W9Pwfj77q
Bz1efyeUuKzx3HNpjKV3YfxzBOE/+FDk2jPIVHWTnv3doJ+s9qBGoV9RYs4k89nXmVTkYTyU24Xz
LmsadyGjBM5AhQkJ3KfGxLJKdSC4PGjkK4Qpo2IchhNAw4oUnC6Jfc4gUo8UTulIqwTbpSP79IeW
nRIhvQJvmb/V+oW2F6NJJSJw3jJNYLm8uGIL07AvWR0ffVdilB0VIKQ/hLD3toqvIg7GQ2SLMaW8
cBNY1K3tcR/2vn/GvFigd5KNWlEIsw61WpJt35KCRE4pFr2HR1b2/pghwoO2BFDCGOPv541zc0cZ
DM1LgGt7F6A7xqOGSFoV2WTKiBQqcqzDsSreqMht5vJc87NePT+Qe/ceP9sFLf6GyG/R6zyov5g1
0d4b7Z314mruhfkh5Z0hqQf0wQUY615cN41hateBfo18L/Kp1+BtgxQ123FP5nYrc9JZw+usqut4
VCyUTbUymyIcuTonH9LYHHJGilP7bGF6zHBvMwMWaGuHTVosRAm6vHnFVd68yLcgdHn31+RHWuoQ
E9WivCW01zmWV+m/wkuaFhWe1QMGjeD/vOYAtH2A3dC9y3Dk1jndiwe5wwguFbmpIK2kC/rEo/4y
/AN+kPH/uv0dmRX9i0eTWrFu3LlxjwXdy3BBc6Qudetl0iFFuegsBrUTSwRy8E45GTLsjNOx7rnQ
xBZpKF7qGrbijLHxRTwOjyp7ziZDafpT9dRboS6gcKusCaRzzshQrP1TAP+sOk4iN2Bby7ATSuaH
K2BzwWpORJGZj6Y+SAhhmQ6OxrAT7BVLsUprqJYnLMgArv3id857P/HAcrX67C06zGohNxwb0a78
azT/ETgCpFzz3XUeEijE2Sqs5lwAOb999hDSlBxKllCrplXQ/ybHgNkSdW+U7UF3a74ZY5vEZFd6
bu7yH/AAmsAD6H+cnBSzlO4BIRYp+sPV/a/FqNq4LW+2G4cKMTbL3nnGxW7JNusvLvo3WBr4vXts
UEN+NbH2qhFoOul//Upca9hCFltNfhmFBmW2MtVFZA3Yj96jHp6fl7jvcVCnj7a0DQq1ifTD/JGX
16ZTNzezt75rqRd2sMSqLo0goph7fDkMJxsAxvbSxs383NofLWorOXAflgqQqCnd1s8rhUC1Fwzd
Y2hhyTdfAZky2Gfzq3cTcjBrot9hMpPqEfGM2/7TKnSOdYXUEmBmA1L8+mbhpTMs+RiA36OkIOki
lPRh1mfL+Q/aSiSe8x54ekDcW5JcjRRYL8R3XBau5j1BzdcDESiLLuMsUhNljUKOJqjas6DAxYeL
rqh8OVzZ1mMUZdH2UTl6pqYdyQiBDRIK4YE85SbwopyUwe0Tjx6qwHv+zgq2NJ2ggKJ5nE2k8RvR
1jYwubNcro44tpyQoonIBTw9CGKIySFKYVBVNW5wb9mebWykK79GRM0ES4ldxjJN3kKDsquAmS9Q
9+I0ONotIvQoxxgxsStBNf0Vo0fhvbNmMgjjTWQCOW5S3OgjAH9MbkkyWl86Dc3qQfYATWCX3O0Y
vFpMKohK/k/ywPAW0CgGZi9b4rxEVhUMdsUOqWqwfzyywjE5NrrI1NXLCMS+tT3e7MMcB74uU1VK
ZHa1mxwT2S+7/s8k+nHKhvPuxiLtB5l7VE25Pyy/QLI08sMYEKgSg2XqT/xsvuQirXzrK0k3uD5B
UfrTq0m2W7pUS0MgyKPREofpQ6N6u5WlDyqZQT98skRmc2J8kEGWud1F3QMiC9IWJx89qdyjqrYx
4o+gzSadc+wOFMJHo3TFVcIGLDiVUZ8Pnvm/BeZGfT8N/GCwETWvbGUKDRzg6TRm5Gd5Gq9aP+7U
tEvreZenI/tKAEFLwyLzSmPQEAQufXIlRsdQgexmZ3aMU61HIxAfejHB3C1ZDva2fEQu4VYG0nrw
9dsIo7FrbhHII7ukC+5E9youiLcakiRkyfwZ9Rd85+v3sQapw3NAL/s5823CXz8j8EUhhK7+0/KP
kg7hILY1e5FTb/J03W/M36eETvabEk2oEVQuMZB5u8KoLz48FdICKlb4nwZ6PogqVrXHaDo72Eea
p/YUxyTeWTJXKTnXv2iZvbvdT61q4TkRHtv8ECUneDtp6Llz2Ek8FVR+y4IVemVLiblKpNyO/CgM
tRdNrWoD34bCLghEi7ibxjSS75hSOM+5wQx3RpMhHRa2LEJEH9c0avSYSQ6ReaExQDW2hVCn/esk
IVMnhK8cvlibbC0QB4Ug7KPV5BApA5TW8gSEJqCXX52ZnJf+MEaGkwooshf5EaiULSNqEowKfUHO
GrbMm/L80UVBcYY45rylLq0qTGDu7Sy1GVAUXKnjgSnQKYGA+/HkmZV4DbxM3Z/+po34JBA10uOt
rh+oCFZQIjyLOsVEjCeUoB19v9xI+RxG7uFbg/g6kbVoA0svNCQBxxQ0QfPc341/1PUTXTHzmhq7
gFYnap/XVZG0cHHTfEzm8PvTwT3kbXpcR2aAgT8hN+7W+TCbHKNoJ1E7cWgoa7WNVOvr0vRhNNyf
IX1m6R6qK+4FoBigvesmdKFlFaVSuUA/M+0QiyO6zrd3r0uF08/93GzFrtduCEkCUwBi+JflR8cK
ynuvfbXcLsYudPdy0bpzXK+CsFTvDrbmopaPY4M9RWWm94D11+sCIghM5UzK5GRmjKCjSX5KEQC2
9KV5LgSbQ9wIqAyVTG+GQw+USOzkFGOuRskJkYHt34wB5fFFDEIilxCq/9NeW5PODnGpKH8Pq68J
EeM7EdUPG4ncHijQyc4k83/CQDuZxQmi8tL/Y4NA8aILXo6ugBF6n8y8nYqaWCNnJoDAPVSjcu8L
NZeuPmeIcaf6W6Shllbk7L352pSu70b2nivYLbLaxHagOI7PS1+TZTkm2XoKJCm/ZPytdFF7rbaq
uKU374o3CAYBuKPw3H6MGR9fonMOXK/3/qslhNBdxgG6I8mQsmW0koWHvNXLjgam3UWbhVISVrCu
9d9QFBoWhQf6QHLTs94DeYzuw8qD3NYKb9Skzn1LMMRhzy7CqAZy5SjnZfNHuMl5IFjMqLbBahOz
0wFmxHCTTM/OE4qm8lqRtpmw8unMh6XkihHSvSOZ+PQW330uuTNdybC9iQlKniTcTJ8F11PFCu0P
Oj+0E9ChZ28SobRXyedMgqejXslphFYsj9ZFh9OO/gOKXlx/DqGv+EWmtAT+arwa84bKgYvqN2pI
z1ZqP79f+KYcx1Z2WGu0+BFceerAxx9j0wxpm5/YZhtdhJLl9eN/CtM+JtBdhN1GnnsIEOLVyQ7p
TaHpcX3v6To8r5keFM4U0TVaPext/3F7t++GPZ+aiSzAM4A2StnGhDW8vHraDG3dxWl5TKuc7Jrz
HrZnC8QTDMfyQYWB0Ehodq51EGYGuoP1WT5mHX5OFdH4rA96lMc+6bOAaM6z7UiWjfQP5rksEv9w
UeTwIvnt2+rdb3X3qF+o68I3r/jFtCg6td8zIao2QjOLn0Szo5/YPv0WLyvtrIh899r83ps/H25+
/ucAVBVEAbrjzquX6YKtU/vZVMxOh53TNYis8M/SRuub/4DddBoSPdDqzm33Ovx2aHdL9vqVVOPg
2hObyn/jwk87608sIgydJbjh4Eg2GDjzXTcWoy2b4iuyEhajuz8wVyBomp81UIMQEh/eWGdZKstX
PGv3Zb26pJZL3BAuhshPZKmIzAvR8eVuDyzO9FZKhxq1seE5zy22EDs7scY3B9Ompoanc/oz2lZm
ygy2+ZSLfRY9HqdfN0R4VTzoEkSHiR9HMFKpxiBbsFhLctHOTdtp8LyMsCeJERFoh/ZcmL+0nTHw
c8Mau2H2c7Z2w3L3YhhpGpkSJ2qezRiScc+8lSvQLLTTOKArCcOBqptODce5MLMhnTQNtrYZT88m
aGV/aVNkh7KuYXInYqgoDGRrvQinB6bGyQ6Lp8+i9A4280RPThupSNkEZ3bu7badsKvEehPmodjN
a8/y6UnEQChB2KSdSeeQh3ctQfUGNscWEDlMnVa2ZYWQwih8ahfcQw6LU6tTge6E8XXdK1Ha0vkM
0QndO2iTM6a/m8EE69CPZ5B1V1Ld56EIaN2Uh9GYMfIzqSnWmrGNcLV2Cl14vbgUq0mnvaDzQOkB
FUT0bCf1Ts2NIhuWMn9Y8RROdS49kFk5BBLJ40RgSfT/P/T4477AOkkK7K7rPKIaC9s22Z+dznoN
H8/goBiH4vE5KG69W61CC8/2YUo1TUUWqCP+q+Rxw17+blzuB3sZU4ntDroE5lAZRHqDs8BbyPXm
//rDO5w9t9y2zTXYzCNAnbAyxotFj9ATjr2hgIjI3qh26ekLqYy0Ljg4BE2hwH3sGqJOvham4RQ0
x4eDZqmEuUWwJnrg6DAv7riwEVBG8e9DwDsL6yIdRmm3ItUyVk6tMI/Rvz16tAcvrn03DK5jk9fk
zE8O08CqBlLsMmGe10vk3xxrDhyBjojmzSCEuAEnuPXbxcynehrczgdqH8UWYAIXf0UVKlDaUkWg
AM2i0J/3/dMCzMD+kh+DMeNiEPmmw4S3JPRoii4MWHuDED6inck0zK+4LYT7MltlZq/h515FyX/y
5eCejgCBU2fhT3232jtOigHzdUPvY+1gvmu6SjQkmHYeIsPT0Z08mm/2Z1PH9ciWzA3snphSe8Yd
FAyx9Myx80LVWWyHAybDrQgNKDxSBTJsAVhMMCVv1JbzNyKNPJ+ryugruosxPTD2M1kk1hnIQUUT
m2SHSKEqVqYBF/7D3KAfTs/znGh6MIFI17Antj4ej9+nJriWXn38z/x4ZTkrc0vsnyR0/dqclAgD
GmGzqwhxcGzi+vYyHvWkprxlRkK0W2rKZA0vmGxj4zcyiUQZ9bBAPvwsbCV3+2GNj9r+a4SmsvY5
Tep6/PzU1Sbv9unevqQCDly8K26x8yWizmGMTK8T9ViUyo2o/jcxd2UhbYXgShMPXgvAMrbsiuOe
gWTwn1i9NsBkqaI4yOi8jKBQKyow5+vHb1tV/yXUfwtFLKU49bdTtZIGpueYuCTlVims05fBxKjg
LMCP3ffgKrTKoALl2jZ7tNuX/1qebrs3gNYplsTwJ9wd+lRu6pyRhKVMGMQA1DM+bb+Kd/kd2h4r
zHscX7l9nkLPquBmIMXPeI7fGpJruDz0JU2j/BHbIaLlEWoOLWaTPJYFC4m4tf+TzuRsHUS2OTO1
57iefHzT2C+LWp0+jxhcS/KCNw+mLK0XK2DSGRBJLun/OfSfsp7WFylzidzRe1KacuyMpzEM2vaN
3a/wNlEuVxHG+6yg92uDD1J4BrljxDUlZANhJFs0t/DjJv4T6PYy9EiuGAnMnpUZ8gRHlaVzGNKf
YMt1QHqYMJsQ/CexEahAOBh31rXpR+Dx1iYP1UYijgyAuxllp18CvmU0APJAT2KmaeznYwEgUjEy
+58zAgHRp0lTo57pwH5Er49YyuH8HtzKF0PUkF4N3uIeed6/VR85WfNjATnMJg5SOzcUMNh81BRc
DejruxOiJtYdsDk79uttFSg96SzwEMmRTARPsKMHxUP8kKnKM/uIegNHzbWyeU1eqhkyGng54Zjp
PV+bYt6tldnaqVvX7jzP2qSZ+N3TPvV44kebuWpZn69W51mptSemApBIMIEqdchaS7UT8d/H2Nyb
Aatn6032UcFW2+FjVc/QTDpeV7UpVXss47Lsd9mI0NaVmljzxawSturJqyc7sYYfqxupqRecp/+k
glviQgQvZTUb9jrzRqiXwdLz2xxKuPES/YQDlyshO/pH+YhHUcwlxPD6eIT4zsWcVrLkfvX+6rT9
LpHUU7AR0HzQmN1W/CixgVc7v1qMouxF1r89sGk2eCgMmUnfpreURZlQ51SNT6m5b6d+v860gWck
YFWPJWyaAOQsUVnNcdW6kVTGVUx155wE6eGsN/3wb+XR6Emll87DcnfQi//ZtCsO4+NlkOdS2ksL
8Fme8hrVtrBxgMnXX+UDUC1+Ykx5eDKG7zhkvY8ufPUlpyiU5A4s8XubpAeqvkDO1kf63KyKjIRa
Dn6XRB64a5GOBZ5RlUTcLi1V4rbpIENJiQIiXjU9W3/FWrgHXVKLnFYvn2tKLk1BoKwmm7UhVyrL
NWQq9Go86Rp2F1fK6nIfFQ4opnXmrfliPkSIPCmLQ/zjxIJAxkbUV6xJSBfVz7NHKvLvfqnNihzV
Tig25BoAogqcE0SIhVpCC/8h7Uyflik23WEmyx1SHG0csRqULZlnMbDcSbKS5LY6FvMdrphmL75E
QzxsH9gg/fy6lXtvQhaImY/QYdzBUugRvh1la+LbLreYV1A2b+zeZ/zn2/s4Wyn1P1re08JqNtHL
3qbIza7XbPHtR4gd54KsREW426azIECBpDCRNncOQYOgfwMl7Z7ihTxkU5kgy9ibPw1J7OeSOp4V
BImiRUs3V3Ebczl/U0rMe4buk/0An1q0oGM22EgBcE2tk61KW610jvOS3+lPOoZUmZfva2JavHtV
tJkTMnwm4PmXXKPjbpe0daTM8XMq4V6D/n4HfjiGLWkMtt/35IWs7MPWm5K0ykXaK5CGdMJ6NqgH
GaYQBVwle9zXCGFyCVYMnHhaOhxdsCEq0SXt+Jiao1aC9wIqXEC0hU/9Na9YhEgYV07hfv0vUY2h
GWx/OwxCJzvTULnGLMMARKu3S/ErfC4zWsicX6aykQcJHSySq3VMKBxtmnlcqwPW2pOSVIB1FLb7
oRcbdU3cSzdwqcxS/zpyg+hd4PxDxZbJnwGbCjZQbdkPin2mE4gKTlDywX6UtoIrj8V2RYdhZFOH
G4RK+W9OYSErqPNJb8YEf5DpZpHgjNU4rAO37hpUVGhlLQr4GwXe7u6pKCBWI7X8xDPtg2JR48Zx
VPMd9VT/8NWPZIG70rpEdIx5J3D335SqiDaWOoHcT49py7L25bZ7xPa47u1XKStMGZ4Z7OvIlhU2
W8ztES9Vsvdza3MoNCSf4J6sIvcPSL1AvvF6+YwvHp1sZ+xdjmsDFzAvZOvB2StSztDyUkFA5vy0
fRjMmE8GgATza7z2ykntwlwjx5nNqlfGtE2A5FNWUwI70Qp9d6fIBqhtP8iKTYttfcgNd9iu82Iz
w+tPYS5e8vRBLCGcoSx69XgQz+11/IOh+n4slEsOjSTQBn/Is8Xk9b6TMVLIZLrxrkw7U+wAVMZQ
G5pdx1Ol7LAazSTfEVXxtHn0o5UCXitXEFcnwPgWWIvHjGBYLEx7COGicD6Mi3T6EPMvJfnu8w7b
P6J4ndCrCMtBFi4wSZ6i0M9SpY6sX/OVxkZmoFlMFbZK5jHNs+P7eWHzOzs+H1fnmCtMSoIZ5R+E
4MSrqTSaIao4ZZZhNRoRAWS4vJbxrMlgT330Fv+XQOuD6SWp2NLJmoTSxV0ivEPkJBBCWhuGkJ05
prS1JwcdrhAfdkIFsgbXNoyRD42ELphBVjR5ztl2lQmi7QGTxqtrRiIbycP6+7kmojtl8/YPmWQY
iPuNneewX7kPE+5EJ2AFv+eHhJG/ksi1e0pi9Xv45B4i+cVMQUSQgvS1EAFX7meux3za5NTLt3RT
W/EDitRthYayorRrCTTX3TR9PLbgKhhhx6uIhLRjk/2iWEHMIrRqVrq67sf+Ni128TAp5Oj1pj0b
zuOl2Lsio2GJ9N++0g27/+7LPCpkQph/LHeccoVTzGkvL67w0MCeenmQHnjnRrZP2f1NDfjwVnZ4
iwmztmpu93wLJ0CU7Ij76d1tXcnUo7s5deNvtkP19keK+Vs79IftptSTuwSTOSOwnHaujGzb5iOh
cD3QupBBMI4ZZ7MWGVvpe0U+89ChC2lSFwanheuDcUsuMaZ9RT9gpZWiznFwZejDwe4/SMe8dPB+
DKq6tz3YKWe5WM33p6wNXmvYicNJRwEgh/QE8Na9bp3Z2zBqESQTpgBRMws2pEyt+sM7GKtdHBr1
E9RqK+LQgJBZdsXi3C2tKxreuE5ak6MdkZfWoSWcVtxbxBOxYTg9qVdJ/Y0iu6LocmFiyYWhdnVw
tSQVBXhAHQlVkhklvj+zAqVjMtoDpvWiVuPI421HE0inb1ekJmXiga1knnSvoVdI0NyxrEEFeZwj
fQvRqCTyeMZyrYPazcCLkHw4z4MNl1nHgAuMLMyjZw1NWD/CzxJenWsRcEOmrL0d1FFtYQKcqK6t
SwGV9bpaE6cNQ0Dw6Kum5Xw2a1p0rIiLD4cH1EAeZQxI9vwi7UkLquZLWmJu0YMIgZwhuQ5iMebM
hY0U21heYm2lTmOel1DTvlAtKQObMuSciw8hakKRgx6s/9+t0rzdY8i2Bs68tFsq2FnXCISLWWJs
/258PIBp/ykbMwwUkTNqsSsV47zc9idwCE3Fx1TEhYSdXIKySLEZ/6phpYoW4stFu++dI1VseGPj
pXpGNOSOClFDF/TswzTEBTB3ALE6etegBG0SvZZ2Z60/+Upzat/MftVMay7sw9QHEUQXBJY4IY8C
xuRdu+O6LXh4wPLjyoDd+Z1Q5pBtVWBsZydM/mh6X0e5Wa87qczM0FbfKLvmYV7YdeHzTaoOFQV8
JLxbt22GaG5ItH6ui/jyDr4pwXL/k/aSFLdBZNc09RK++a13ECzgCYLzZK79XkaUX+JtHMJHHt3Q
czvzLf5vfv7qbQPaiNPMxdZxdIgPk4kf4HZfl4fOXUPvKb/6Gr/TW3JGNvs1qSpPhFQtk3i8+tSB
zywCyG60LADbjMqOft716ttiXk+5u5oRSTgQN6zBRVvyEhTLbv+SeJ3tDHWt7mf9nB1j7pQ9YENR
+1vLJILzH+LBksg6YnA0TqqOI7z5T2W0fk2L3MMVhyLy7cnbOL7BrPkQuDMSMF7M/0L3cw4/6wWb
F8fovCR0GDjt7ZsHJpK210UCJZSe7y1hWOnjpm3uMVI+SEq5JP24URnqG7i/RPOUuzRbgQdo9Z8v
eNUv/4qaU6okPiHiiDAlcuFb/P/UdCXBpOQNYD8YMqD7S9cop+d19jKLK/9vkXQpkBTqpPQRTpGy
nRu2Aa2Kt4ggQuGKXFBPzMqgt7GCzmgHT34rUASxo192sTdtqgNtAsIlvJNWdquKA5iwtknYG/+0
NmFTpbudI4ZEOarOYpaeOJTz5U0RzjRpLT+dMUFx+ljuNbH7ZW2lSto9ZUa4Xc6owXjUJ2qTnKwN
NdxsqqMdUk0kDbA3LtkbteK3RwWLq4nSh6yOZS0zY+VD6BuWRBPDRZx7FPvhaKa/2lZnJi/aTHig
fyQ21yxxjnjhPS/rcAPr8VwMU81EZlL/RqV1aisziYxZcEv+Yp1yS0ymjbaPJ0j3iOKoEGHYiDOc
Nhp8Yg1SXtudvX4icCBvizaVFQYc7sLYGZeJn/WIHJEgIoF281ETDQr0UarNf1MRA+9HPpAYfGjv
5oJmuqbNANMbS7cVhS3JZ+3n4NDdhXU2GS5iK/vdRcBWHq0AfIDCxkxvbUEDvt3eQ9awRzPaTmQV
mgLpvQhlT8pqv43ePDzrKHbJZeeJr4Dgf7P42qZfLc9CsDSPwOn2vDc9f9kvROYuoegkxZbarIzN
XoUPLqwluQIHydsjE/kS9gdm34/hMdbILo4vFhtnmQfvkuKXR/gMIIROjCgEh4lj/BIEo8FZ4eta
3p2g9rodpLrRZVllixMFq/zYAf4/GGBWzETK1ZUcMX7jx4nxvbbpDD+tqfaMecQA7Xi6SxX2L41N
r+f/7ObSV6QC/wQY5uQrU5o9FM+1OsUeYAGZ984cnTxzu+SWIqqFmVR6qKIvSMnZle8Q9jXiUGq1
JdpG6o7dfSMTpLCvAkmTrFng7naVJo26p9tqGhx0Z9ynXDYwVUUa4flpI2xSuFQyj/wLApYWcnO5
aJ+OpxZIgS8tPVeqjTvSj2/BLUnHqyOdRRL0/pR2hIoPQYvpT8rWylu1nmdRjdnZtogx2SzJgINM
/okPe23gSYx0g5X88N+pQzThYHITeM5Cg5uZywTOJComJubpI1C33h8kJO5DBm3Qq1FQSKzh48D9
itg115mOUcZzFfej5m9XhwC8AvU4+ZquMb7Z3t6YTGajXvExOrcSBsR6DcIP46iyB0ZzSM/Uq5ks
BnkEmXyPlcENocDRbgBt0dYJhj8V4OwNqBmry7Iz8KnCFGRa1PI1U/jz6NjOHpBBG4nQ3v6dE0Lz
QPvdsCQVemCodikOD8C448UeMV8yZlEYxkzl3mr1+S/SlbH9y/7ikt5UahG3acZ8LPG9a9QlGz2N
8YmJejC9obgB0VADqbC+Pr3cL7Up+52IgsfJby6AISCaZUius/cBUQSFMutkFzdkry/hRQeZPAFq
+K4IWL0LNBhME1S6HRiXeTPjqFNYNrcW3aFvBmsre5OhhxP57ETXRvfhNXBdKAcmUxWO5Nftzij9
s0szUMUseeZn9SqwRmklMMhj90y3ADhhi7993PDh9Vk4b7XmGbVst+s//zhvE51qxEuvt0Wlppw7
u/ybVK+4d2RrBNHO64xgA0JzZu6q6qEeL5TRiBxwSzH4rcPB3xYCvCzxjlOIXVX/4KG3pDu31CGz
YWSMi4pH3nsaxzhki2YKYnAOzse6R0jeQV4PNIuXyTx/BE1AL72ucrt4DBzMZ2HZZayGOQrDuCxF
K+t9Q5/302BJaCCSGOTpWidv03xLZqtVOrQKjIL1Ya8onmMmPlRPB/Tvkpg/fLncV3f40JdL4Zzk
CavThd1cryauDZmDgii7l5H9PxBwgizW3kJhrMvWimzTUOGAUi3bXb7KqeQIGrWP6achyFg2evsm
rtuZRjaTyi83k8+sxXT3PgRqLZZi7G2X96a9ok9e7WOxbFn/43CGXhzJrjyeJa5HjS5xjUl42Kmn
Y+QjFwZWyaXdbf8dCT8tWg+XFSJ/QIBUOQXVJpwR6HfW1ctJuqnrhBuJZ+0iENwL3RXUQxOWDrGG
B+ekQrpqcRpJfwGsFUd7SDzmNh4r8goTO8tb5FHG3hqoWnChQLxzcHf3y0BcdRNPy+nNKh30DWud
ftu4nTXdrFqwcRYHLB9LavJTvuVXYFY5Fcdg+4+flAaPMl5oO9g3BZ1cTpbbiptIvSFMgA9Lpd7J
x628NxHdIWBNXxLQHN1Q9n5MuhScqpKBQrUQSGiqiDAbo2sE43dcBNRdftjrz7OO+HeXsiL426Di
ya1OhHNkUqr2yN3vbGz4L0glmtQMb5eHeni+jkmEOO+0IeTs3X0191C0z5ZuUuc+y7jWWRU5HQrD
WGt7y89e7YQRT7ReF73On3EtWHzzB/egOsLcbPmrqIsZfWY3Ng2EC+/NX4aUyikiBLpnkT7hW2t5
FfIbIdwkLDlq6O2OZys6BIzhGTdF+xxvG7/xR9AAjy2eNc8p5iY+9/LiAJEnLNGZptL/+9nE7ncP
5ADVwJ4JaOjZNGjhofVQcOqldVstpMcUfUMPuv8ZpJXWrV7BpX4orWTY1qei7mO0O18mmp6pHuqw
bnNIGSszci+cvV+nIT9RKtz0ZpxS8zF1pSCeluWYUTNy5urwlqM9rKD5BZaTX2mpL+oVWli/Ko2U
ixAqPldgVPaiMlfXIQ4Td1IW7QuuGu5INv9uRv0U4tjm2EIGkfH6Sp1GUymAhHUQw24NLWp0oFr0
DFEUvbxBql8H9CiByLGEHQa65PY9inN003uIoEeqd1G3tFDVB+2jkob8AJtiehoD9PmhFAuyzDL0
QvzHc8JBWX0ACnNY0eI/hoUf3sOJfqDh8i7MfyAh9U8LPDBAkhtY9yWkT+89yyk8wGW1aa4LtQQl
sKzsnDwJTzhfFATBszkKs0RDEWBLf/gv/4+fXP+cWpEoD9cLHc5e7dEydMqPF7YbQo3Ur9MXv9Fu
TI7Egk9DaxQeBIKfKCJVa2DjhG0Aar5GahXXYQe4dehtbWethlNtPw2Gu5WjwR+Fhl2HXXUCcb4R
bpq1iH3tK9ZLIc/rgFSI5ZA4My0X0azAZLqPVn6Vc5nx+r1SGA7vQaSdRV8vrFRvgMe2ky6Y6r7S
Z72nD3yXEkbc70mWXwJ13p6KMEzdFeB+ngIrcOwlQCuVelvjBH/BwgoFiZuDeb0zLkHpAsGJCF9Z
nNXAYUb+eEKXxYF8wkkB0K2Thq7NnhqeEtC6S0C1euYZtiw9rF6b+HyKtdjAYQ/FMwcWK8j3d/k0
udwWAaPZbW80EAtLMnAjfxe088iFU41YwEH0sWazeDnMIjr+33rCGHXr9jP1tpayAOqccg6sY4C5
HOIYgeapBb+ICF3hJSELfGnrgW77eTPTJ8eqFVqiLIIvV86s3a8SJNbgJv8QLY7tDyjgL4k5udpB
Elo8fIPlJoFjGrU+TWaxQNL0Vk+AbaZZedHZHpywZAJ6Qc2AXRovn3sDUuT4676UG46KCWVdVkEe
1VBaugVmZ19x1qbZtzXysk67RmD5/RyDrVLgO2B5nUeCi+EVfbI6EW7sBXD0Z1VtQtxQqODShGJ+
WvN0gXH3ZIYPSKrfbkpC7J1Tu4uwbCO5jV/54xTaU1f01Ti71lbeBABrAr0zSl/iUzx05KhPyVRc
G/QNbq8tFzaAiAm6OaEdYQildqk7AYRn6gVEJ8YqXUEptBsxAX4GrI7kTJwbnL7jrho2kaGcRe+x
Lia0BsP4J1UyQyWXWt90ii6woJESWddhRFKxHuA69+ni/6Yg8eBwIlOkT+dS5oxwsoulafTNknkc
Qx0FpBbbHn+ieBPkU9CALQeFGQTZROjlohq1+5HHapzH5SKQl8M+gIc+iAp07Jj0zgwSVSteuVDu
v5G9wm9+RzerPqO4IeQahfN54tVDSTiiXwlXo6rPR5PUFDJYh4trE6i72w1iiJetonVLHPMbVzRY
9b5qoiBWHpU6Wq4IrCJOo4tUzm2NoJnmECwnYFR19knA7y3hI418dN/L/fnnwVYIpb5v6PJhrlrq
ICNxPlGJGfPyH6PbwnJG4QxyFr36/i7Itr/CMGx4TS2FPoGF4chguHR+6sEXUQSG6pRP1TGladb1
RYeAJ3Xk6m2qH2wfuaeASsxeYpNvR+sNMKNKid7PwGhCOz8qAPJ3bVVlqFI4qRUsyoYWkyznV4++
W085O6JMSjlCdBhXONCYNz3kaWvRuPJ9Xw8HqyzgI8mObizD171T+7Dx8QZKiZ2ram4xCS13Vwi8
mi0av7BbsV5LGgdlF5bTBx479H5NsuWvpUlsflPqrErWdTK9H84onY/soeDou/9/Ap80BeJcLbtp
RaucbhLjJGDxU2Oe/4K3T2y+7oFBFnRbEjXtUz7l158c1vGwmQ1U65rzIYpBGOm6+CXd+LAGivi+
FXRY7aAr/PVMB2ECv+dUJElTNIw6zYbn0uNmPUSgZQrxI4oToamlgc0Kric9DUEEC7dfsueiUgHO
FbnZFLcgvRWxcgPubfv/aLemkLuv/qOnwieLJsax/IloqCm4nxiozPSut/ylxwloKInyJYAtpY64
r4A+wNbzhAQloOGTj461ovCchGZRT48WTXC+leOg7nx0uIx5cQs7MKI9q+iLXeltAFzupA32909G
SvxdYA3s3QdYR/g8MLA4pNdvYobkyOYzii4D0L1L6VvYM/MWm6gaOBxXoUIkghLwllexIfZOHIGt
lEScVrTA3tLyVVJheJiH1azW3FFeqXg2WHKwiK6bUT/EdcAm0d22sgB11U8mJCCYLhTm1zUZGgeH
UGy8zhCH1qmE/C3z652pErrGW/bBt0kIMJcgWgZjbtKRb1a/DX0vgC5YYFHKseRunjEmv/aphpDM
wwaLeBHk2rz4e9amE2aRWYQAZCp5vH/KksZjzpOMMHTn9VJLvoVS4VaFQhD6IoIxdiLP2NTvaO8m
HAlNvhH/250JzDWxIHRb7fIawHlTKSgWyoRsGTWZDq00CAZfhfaAhNle/qvVbl/fOxyGVvX7gl93
7W5yRZlFf7Js1KP9WpVpkf0q+7ZLIlc3aSdna+aJ3Dd1V3hdX3yAMeA77XD4F/pBejPMjR6uAoS6
rq/ECGO1ChdmEbx5Rb2toaHvUJw2g3TKtDHpxQWOWQsZyXe8idizRqIekF5DERW+eIldaG3T16Ib
R45GKOYeaA20XEmmm5SGoFfxDdabD5WbUlSCaQmDPRkt8xusLZCW35E3F151TVIa7erO+VtDulml
a7uxLkA5y1MTWSSmW00KFosLrCA9ShZHAgCefx1ezquwRXykdfxiZdVBAbQ+0sM8hcmkMPB0iM3i
SIdwf4BxcJGWiTi6QVJGy4721GeAMoVJ4XOfyfg+CrD8g6IaI7KXGtvGYgERbdU76w0bneOLYbZR
QhEIwg/2Eu12F51uLP7LPLTW0Uhids/oqEMnmwv6z3KriPJIC9deKywqTf8L39YytWv6cvynsLlq
pYGqsAHxqWxGk7t7kLtRTiGkw5mhybjnvO/zk1Y+iPSKBLDEvFmvQ2M78g/KeFtii1i6QI4z3ARu
5nbAPO0v2jg/68KbaJMTaG+SP1Dv+M/yqcyy56tGfimix1Zm619EREMqrRxyjcdAKCL5sRpcgm1h
m9O1B/MvQz8fFVzRwmf4HkUI7UPu+NDgJ7QBqAfUmXx6uErsXEK5tb/pRSr+pIezOuu6CBn8qTq4
cKpOD9GzX7ySwgZLDIvroGg7WIgSF8T2CDn6WsTxPFPsueUvOGvfAv3WU0dRFieKwT0SGa4+8DMp
bSgG0svr+BMX397K2fgxjCfgED2CG5uCPAu5t/8vgOl9DjZ+ZmY6uz4QWGbkrhhEBvh7yajeSi3e
+TupWa7Nit4RjYElp74DYqoKrFi2hfyhTMWLF6n91fHj0yZO/u+8osvcaNBMESvDjnYCOJrR/B3K
TioQDhOesQJQNQxg3YSDEwujqVFcAa5EAQs7o0Un1XdWIahE8tWVTrwz2zTeg3N4Xcqw6ZwiEc9P
/QCcT3tV0xnJ09rMzw3f49YT/CR+UoyRXbzZwEqdo0rc70ZfQ5vWpbAasUsMxQa6gLo5adstELfG
puOc4sLr0jsoK6w96mAFvAQYQDG6YECYOpMqKO7LydOmTsPXfq3zRNSt8bn1ce+Pn1ACs8KkPUI9
rpiFNIPdnSej+uuPn4hMHaW0oUd/AZiMInwb6u3CheWVnyMGj8Lp8g2/X/qJqCxm3okF1Mr64iws
Pc8JDNqV41hYUocAl2OpOLlDus1JtDkEQ4E/DwsH4fRAIAd6h5cQoYRfaMMrcBZkcUAAyLdcSOhz
lmcPVVTDQPlXxyUf2uuj1eUN/8ESA9w97kYk9onSGDkvxou4hV4/Hzd4EYKp2k6Lb5a2y3N5FGOO
4DO7LtLoGTwGTXjKbHK0nVLNJ+soc82kXfd2Roor7nOPv2ph/BZOO1HDu/784o3dhh9/fT29cuOb
N39UGw9JXWUTApc//A19ZHWpL6pkacsOgUTD+CKna1rMR8lyMMalnOgmlsghIPAipjbF+O4v4y0b
wl403dVWKSU9UslRD1DFevmc9JpdfwbSBEpNIzj8tRQKZhgMrF41qQiRb6wot8J/645+vXAHeolB
wpG26xp7r23wHA9drXj4WVpuJh2N0ZhNpQvf1RUUFep4PjtPvQsQNX1I3kpYEdYvgPovy8IqG35J
6oYb730M5GWacvozOD4JJPv0P7VvxXNRcWXpb8Oa/M8jrr1gM0FbTlNompRQYNdNp6UmGUOFCUAg
okcDY1t/Tacc9/moapp9IvL0ogVmbZNO3X5K131+iQ6Ao4H1a6rDD7A6PsXssglq/+RSsCuf6UfZ
3shc/lf671aEX4CGS1CqV6heDNaFFI8ii8cO6He+QojiQyhgQDbJsnnosWOzIJ7gTrTf7NPPucyS
L6cDg2vfqz5smxIiiwKX7zJKDue0kmBtidOTpG7i9ywEVEGJoeQo3jwhMW0fjoyqq5qeOwd0KqNg
TYbciv2Eh6yvIGWpjCGO1ZK/X8opGMkZMCRN693zwDNmbj5jLj8JoRsd5nSflFUg/p6+l2sS7qmt
p+pqcFknRpBzGxnRjXvf5iIb2cVo4Jk2Cqhv/wekYbAkzpOmkoA0eT5PTKZssXDMyXKskVUZLBB8
V2hzvdKHg+p7vG5962vs6nAplK8MMqmbF77CpXLIOVLPlm/z86EZDdRBLbXpzCsXZjDRvmvvmm8R
O1FehqvQ1D+HORgBhnn07yGLc+E9c1XeroZO4nGkV7YFR9JKtuTIFxiV4l30rLPJou0U6TBc/1fr
8GKJAuDSA1LtObIXXPt+aSkyPoRAQwHl6yjtVFN53MuSm6YlVenYJNubClImj/t0e4+k/XJOSPWw
FzhWq//bNtS/dEhITRRRptwP02ZLupPk57hUq1+uBQvNnZkTP9f2F1ILbnDyww4Wbw+HvGzLUPJb
KzxqTB48PhzyBB9r65UTjA5Q4dfZ1Or8hYoKzo9NzQTqJz52X7RVhNaecIyyJjEyPF1GsOXwiD7C
xI0VR1EBIt1vZTid0bW3Pgr4ZtK5enC/lFsGwpNVi5tU2SiC2OrbgU8lXfivn0O/CtN3xAd9PV2l
yENXNr6yrfMzBvmkjr81hudUvYGLbCqwD18LSTdrZjgxuD92zJpqY0RmRCawp7b4BIlBy5w8047y
e3Sp6dbb+IejqAV+y3FtH9aiCdTl6WW3XCJ80QE2JQGRxwkZiUDiR0WShr+NYLF8Zney49ElaHVB
fDarl7emXDJBJUKL64Imo3kGV1AUDfIz0GOCxMiTOQoBm3CeoIZjk9RLfEW2fRxkxo2mlT3pb6fY
m2x+KlAT+ElmfA8VcN9dnz9kflFgo/5JfAVRvsthKELgCtmMr2fTEBf9lyRDErmCH0ORF6uv+O7L
Do1PdS6Oy0gmoPJ7nuixGLGAx4f7FkWFCvgz7KFkDDQP2BgatytFMN9rhBUJQ96p/QG5i8Y8AfCx
HiSv/ouUfjxlWcqurGbmp9cbO9o+wHydsAMmC68mlI21bvOBQbOGgFHwVuDjJcOyU8GIKveV3aU6
diwVhOdb3PLtXKNYSWlbjWKin56hr1FXsmbe0WJJ6GapjVewQSpqyDBWijStgSgoS+BWg3bRjV2q
gUnvrD9d1EImkd0sTciG9krrSvpGCbXg/MTw/leenOOCtOKUC+0Cyvd5Vzcw/huuXpGBoBLfiGBN
fiarDQlbUEh2DkDYzN74fSW5R+QF8lIUBN61AxRreIL5Yp4TWE7JmccBdBc3F2IHVt0yLwPteLMO
/+Ma9DOtLGBtGDn9WKCgqqCDTjl4yCtsHNUykrRzu/C9ia09Eu95JpS+BOldAxatLox6WWEspSW+
35H4Yc5PA4yofFxw5KMhdOd8FzZlopIJ+5l8Sct43D2H2A0vvK6qjQeW42FbDW16pOI3TQVMCYfU
ICCVacFButyk1koRjFtEuGpBwZUMY5yHHNyZ1gRoBci9Ijoa5IyWkUK+vs51u81sVpEiyYLFvH2h
8qvyKr92SB+qg4P0YqayphKG5322Q7xA0UYi7rwT33u0+/XZVe58mpK/WkJzfe9MnPsK8pTXzt3c
6acW1+dvz5AlPxH2ePz9sH5W4CBfr4Jm/nTBkRAzh12GRVDscgQJbUQ5o+Q0VdvzlGpNBo5/rVxw
8Pnad7lcbc7CEcwg8+mb/HHzQGJ2Ja7+MWMNDje/AvjGzPYLk1zqTl3pwvj2+46L/5lHpkd1X0Kq
mtUIf5l0rg2K2qxhqgWQ0rP9FVos/h+xfz0BGVMUlJtRpiijzMDAwlEeJpLFtP/ZN1jCLlYoznyB
fidDoCyKKX2bUSBJBNlJQM3A8N/XN9AuqiwW5BvsVTyy8Zwc0R3TLOEIkbPa8sM9XMTvW4u7g87b
BnKZcEjsfOutHqceY85qPy7c/T1OPE+VNbe9git3LH3mlnsKanJNKd51BNyTxundSjpfcAzzV8oN
bTmgLBB/6FZ2ccsacZVsegxsiLCdXcovNbbH3oNS8SImz2dDEwLZ7BQXQJNwF/1dr+r5JyjqCWzH
APCZcqPykM2Izmx9uKbieNewggG2OwxB/cf4E5mvtBri14KhLSzUdCG98lHt85F2Y10ezZ7Nsu+o
2aNCE0tdgMS6U1Y2BKSUBmwd4Tg1QpWhpC93tC+aXT22eplaAlb0p9FtmtUX3BAoC47ZYawsFZd/
eUkeEK/MZJzEs11iWpqBq3mUhN0hBst5mFlWbV7VYt4hNzaRTFdQwhKJ2oimK4VhDtKGfVL56pLl
ZCYz3+n9Tzhx+p88teSIjwPjDceFYEPowSBIRbKa5EozvQa4fhiP3NKBGqD9Lr2Lm6HJ8wtW1kwJ
H0Ob5O8jrRuipLy0C4R2e0dhAsWKGxXJAIFDR+3LscwKV3Si1XK0E+DWCHXbEc3OraBoLa2u+5fR
VilN+PlsfwoyYNvD9RG3ZuqHlDY3E/TFuKjpyYOkg7D4kc1xFKncFUboUBisn1PS3kgT+lWznWly
1h6B1Ny3UOMnEYmFU3kagEewJyV2sTuUoWvuMQ7rJzyAYKhigGmtijNSfPjnv8U7nsr2+Mu02LuE
3qSc71bAYCHCz0+qBzPwuCTd79I/SMIq/stHkj1kVSvU1IaaZhoRaPY33HrfIylk5LcipawvLoh2
pZ3pMAMBXyqdzoNHEQpVOpy0fCnS5pB2CEwephiz4TGI4lqXTYz8HdbJMtJ7dI75Si9BCSYvu867
odQd8jQ2cY4tHjrslCAGJKXMO3Bdxy3TOt/UUmgJByAcKm2Ti7x4O2eqoXvBD3hCqMu/AQ8FTY8m
3hYTdh7PR8agQseR9McYk2NsKbWtMQD542Qd3fimNXYdG5TsR7dBM9QKHC9heN1naoNPAnGA5KFF
h+RT5pOFL4FaXhcXf5Qfj3y4WAsq2aI4bea2PjJLLWienQNVMuKzAyoTaRkM6VRniCmaUichbjlX
TuZ677DsJ4bknL1065dsco1ZKwMzS9Mo73rJqQw+6Nyoj4/bZJfWJKdzXBi3Hu4hwHaJ3fKuWYFn
O7iB1OA+TrCXfFjFBAYWojT+3N4mNGGnF5JydyDOqudZcwolp5M8bqiqcBKKcX+JbH/CXNrTWTeL
Mg0m86vgj/MfeG+heAFZgLlR74zC3X32GqklhDQrgUBT9BNgNt47APWhlMvoCSR3aDHTSlR40iyk
gaNAX3Xcu9L0iH73o5Fod6ztC+UUWrdBgQhhyDGTAVyEXdMpFTwYvOEnfQ4zBwVm/9zIM6FNStVD
5tSO1tzB45AMi2o30O5UCnKzd3jWr37NkKQyRtcWNnuXhQ/LmPUsBFaYwVhi+9OlII5NY9R85tEs
XqC5h21g0NQCeC7iMmyWoMrks3at/GMN4Sdv7EAh+Kd+UNfo6N4jCNKrA60yze1q7enJ79/HxEYD
L9dfjPTipoo/5GzrFZFNdXDawDS9SMzR+U+ewDyDBlRrSUn7wIr9rnqfXHOoCeOGqSttl99c4wot
6YmgfFnMiB7djCPPaRMAK9GZBFHtwEWy8BGfr+2G9q5mkP6YYoO4kE3TVD7ENTA5DE7+sfPpTecS
hR+HTqbHbPDHAQIW5N/UXcXRubYtUlZ6mQHpTvkSYFQZNAEAADwcEtNicYeBqMRHmVba7D+PA6Wn
aauh/fwRhUvcSTNMx/HWeYjg8a0FY2m3b0S6uceuhs/qdLSclVnNCo9qmq3sqmSkoc3fyWYxc+FL
SWEz4A18Tu4nQx3lKLY6bwcb1wXBWP4UzkkXI/ZYTeeCPFtTPBVh5YWtNgDgJTx+GutXV72Pzqaj
BwvKoVjyIwrIF1regtKHymIADXRiLen6Ai9OrPFpiYvc/CO1C/gQFPXYquBXMKvK92zOslq2lcx2
4u5qIbfareOMbzrWOj7GTxkD9wweQwb8YjGoVXzerJ18BF8Tsl1Nd+4NhdTBg2savki2n3O46lXx
/Kw3MX5D9LE5yK/DEjlbgDbAn7LKt13isFVdOWlCZwjh30oKr/VBtr2SWel8WxJ3U8TZ83pj5RmJ
by68YKsaW1JS2QoCZ/0bBdY9FnH3J9Alms1/aN3ljm0OYbgLEyMTgoseMNW0XrF4X+UKLjILT+9n
QaWtRBxwoRL9sSgjmAIQN5sJbVYYv2d4kBjQhhLEAQZ7EmyclUDwbHUjd7tJWL1aQXrt9tiB5bdE
7u7nUCUhI4+/qdRjjOJU6HO9Wimlh7S6uF0XR9WhsTmlowHsx9E8D3Dmvnnm1tBXhmoLQr04lCbz
+tE17Y3d2HPTY6sb+LGqdocUXC3XvTJrS6g3i/W9zfIAR7minCZcs/2hdNDap5jNZsi+MbfluIPY
Cxoz/LX/XV4PgYCoDknu8Fw/trbqRG7hagzZ6isYL5N0g6V6y+G8OiGj41JK8HVznHLUWbsvYmuz
0WPsR+z363MmSguYma1Sc3Itt/ZKTwUunoKO4Y8TYofT+NqBFdnvyrI6CCs8bU/1t3M+ExfYGNRo
OVREN/ZSkfx0KT6Z+mycKNMVtRht6ymrbfHbyKfr/BcVTxs5iYaJSDyyAz7KEibAGf4TwvSdBdNN
WcAmIFuWq548Nww1OyGEmpoEvNS8vbpHAiZKFrU2ExC3lLQJ3p7n5LeCUtN10ihBneG3VfBPd8p2
g2LaiDsf8qJstPBZIMHaycorx6Zy8ELhWeEYgEdLkSzplaDkd6ngPtsg0l9kb4UZDjVVjfqu5Bj7
hxt7wBG0GrMnk72U/tbpmRaX++ehqPfcnzJ6hdzLRA+89KqsQ/x17qqRZf2us3YqVv/CdxTIZNdA
KEBf3FZW2stoEy9tKQHrTWCXYqiaZMWiOrka2YhjpzJc9ZxDKseD+5T3rVzsJdwCaNhtCU62+JS9
tZR9rbHgNZlL28iidoGu6ypzlmDYGjoFzGqgmMku5woFhx94pvTMQjZMeFxLwgCajeJmkIsF40/U
WP93adg0j6SxwO5r/+7w+brlMPwestOqBp0oC4DIbMALEJ5sGoBofdHlX9hKRLiFRPJUediKq+Ra
rrIhKjfZ/8cvIwfKfWConnBVQe+78Qey5GBQfLDCHGAdDC+E1jmkg5E0HjFwWKjLGCgQdclT3rmq
6m2lxq3qe6fNPNfXkbnPWjPc8QBRyAOxIkXHNxhm+oaumDeCogCea4fe8AYAA+zcS0WEWPRuO4uQ
LdAt0OmirdGWBOAlTh5koRWrJsqLCSYX3C35isnLUjiRPrM2lQZZNLXyzEt2LrQ8FwLfxIE8bW3r
DPmDYdGXSfpwQs1OOIaERvl/Dhx/uIT7t+MsCqr741sVQSbdY4X+r9O7tnVIjcDehaxwo7ASqkPl
BQbrrt3yQb5tdlO1aVrlqay3OOYyXI4rPoQZaBuGYH+DuEKFpdk0BYZ3PGIwq8Jv9+gTpvXr6Q+A
8VyApyux7I9QwaRXBzXXJmjq8b4RBz8YoKFr/cPG678W7W9lvwRl4DLW5CjZgmtsUdyZQswbE1F6
hqORhxjHP/cyVqNLxnXYi+JRN/q/PYYLfQzBywWAx7q9SjKvXQrTfp4cKCfmOZmEEipZrNR9O25p
6J5HeIX8Id1iSVB5E4erJzBZI271VFC4rdojyGHlwoXzko9MmnKZ9aHwCuZdJZ+PlWdWYsn+jWpk
cK6kID4HOA1/5UxTv+2K9NzNCj+JPTF/ehRY3lweNI4q5SmDSfOlF9KQIdaqOeVkMcR+sSu9nu00
v8gMYRmYOb/cl5HdJzpoF66iQw+HuZqY+cg8C/OJYu2zbRR3LrszgnthmKXcDUVqDc95nvSxLB8Y
PXUtxcvMjzEVbQQWtTZOvQ28yp6SInMhP9NbA12R+1qK3tYjH1lAVzQ6r0vb1510//Cey/YEQxNy
dU0gGoiDV1CrWX8ToXnJEQ+CyJWGeulveUGNGAQVj9qCNFbevHxX7ogsPmyDuDyDyDsCwcG7TQ59
bT3xFegacg/dqdA0fABYNt/TGDIQqHl5NHljlwH73bjZLpbvJJGrZDodCFXKyakcCQwuDM+HePOk
BEW74YWrDb+VSp3nVOwXYIvyXphKal/40Mvi3/2nFgYrs7lEu8GthfSNHue6W4bOT33EVU/YGU/8
v+p7Dz7BmkdwabofZn5I+0mBmJJPdw4m5fiqnrV4o2EZgPVQbLkbetG1iYctbXUKwQdCwz9gGrXb
0S4txFNL1y+5ADyN+yL0kd2sxHHRgZTGWSNZrODIRFzblu4bKaElXyFmq3GkliFM8G5UcAGBAeZy
ES+fiIuBJJCZhFV+7r4T3g52LX3Jloq41pFosCTToFXCjloPh0q3oDeMeSZSj2637z1Pdq95ecuZ
UmFAUGuv49DOodceZHNtKNyF+XqDCmpFz9IC9Y8sVJbOc7wX/5bASQTZwe4hI2Z2lpkXnZ1j+g02
4qMyQwFfbrPiQedDB9LccRxbegIdC63v04yKrF7Rg6D+v089RRW6g0bkaKOU0IPlryBKfbvYp1N5
rWP6opYc8a4REQ01AX0jEoFNsQAjFYhZERbDknHOP0/aCpu1XklAR8R2Hd9F5atnqePX6kzI5m8s
u0X+UiMYxfuCFQSfNROIV7FU1AqsSJRfcIfn4KhePSziXiJK3YtyAbax07BFappZTyg4BA9kAwJz
52Vdl2oFiwc5XATUSgj5Qht3cG8IoIldwqXLCOmq/MYFfX/8fSw3BEoJyDX9S6yt8dD6GGrj2liz
vePOlmOJLLJxgUjZsurPJWxBNoQ882t3NvT2OfEYLVAWs/KayPeG1/oAfW2U6jNPB/wJ0lztB3Si
YrGXpUUkuzHjsQP+t/e9VtF+P61ovBbnZwWiy8dV2mTzHRzqvYYKP9aonXlEc32gY6jO43uEMhV8
8LZmJRjSseMLdlQZjAyBSP9pIxYtHR4LdEpWV++tL8Dq4+oIWjsP81a6qs97NpiiIjhSjOdm6UI8
yCLse3pmZ4LnuXg3xKmJbGpNyAbkFNeyWkIBe3wqNgWPWlqf9Kh7u4sxUJBVaLGYQdRTn0INIXGl
4lK89SPJP2IH6sxIN9MUnBU39qC2s6RXYbtEWwlw6c5+hePLf6jKr+W05kxL/V6TYwOBw315+Dsv
X2rrfznM32qKKpDg/QrRjRyToL3O91nT15L5ytH6ImzIc691R1aWmgm9KfW+GtBU4waqPRTSEPm9
LrE04p76JEYu50/U2wr8c7DoEhv8yG7FXTF1T/7QOc27D43T2LbcefYUeEEs7nmnrJTGj2sL8r6+
hc3Y+MPKXFAnkgZ4ZFsf/lAJFr3m23njAVKXT+AnwU2qqGutQc9NF8gNdr1UrnmpbxV7iP4fYOLD
4U/GhJpUhMKiNRQPhUsmMQNmuomcRiaEWzmKZy4nbHkVqMll+UtgsGbaBhrQH4ucThPyHoeDPHoJ
ABWSoi7p7tqO31F3TEzEZSgmRVZdf2+aKx424hGFWlQSq26Cf7w3A+JV7CtY6mlXGZ6rCLefXKXf
Nnf5u/7NXuLk+Wpf1j5NyPjCkJpH4/M8+//2twZ2XnvaiAl3xsLZPljE6Zt0i8LolBDaj+aZel5B
ifIKWWTdoEYSKnBOi9lrCgK/dR3j+022a037f7ZiKoBBgwrBnYXa1eC8q7FdZOLiQ4yYVSDQEp3+
zu35+mgeNIpxNJeozqeL5tRvAvf1zQyIjHHWGBSTlJPu1IQwiha4PtN+6M2Dl8LqEDEnhqX+SkRo
i6jsZ3X2tSt1lNG/wbfYH5JOsv+y5KJyk1ngPn960RDvHEhGhQ1ldRnzKVfYyq4WhRHgkiYD62cE
T1bU362vqzZXy/t82mRW61OE+CLOc1YffO557xpe2FFRVWHHG1vKwh98Rns2HNugF2fA+YU+efBN
QlpUxByXTb9I/G0gkVZEb+8JhnP6tDptoJdZuJnmDOAbDeQ46MNrVD1SAsGywGesVnrFKSYdI5/+
MFu+ENID4DAbw1PXkQea5XfT6356ihCz+Q72CJUirtI6gvZCKxC/Iqbrj8qcgAmmK/B/s4/p4R/w
4FtMBmJPpVls0IcEb571Eo9FeBcc8P54L699tLyT3YzgfYNG4DPbJ+07el9PurPrIALcqAZ0SYAr
y2o20SBQe6Ot9zPX7J7lQa8c5JL5rWypVSZa6NrPXtWUvUwWqj7Pg1EOpmEhqIVUu23Nxg5lRxLT
TtY2R7nxp00nhOzXOREf49PifJQKkSrfrFBn5kJc/x3tCXWQUBdGD8Y4Jr0g2vxNjvJp6JYJ+8XI
c18GJ0Ih+hrxC3IoVfjPG3VUnmGNw4tp6DHKcz8z8s/9ffXJRGtdx/0XDMFUR4KNM9L0U09vZpqF
MmbVYxD6Gk3+DUpXu67/I7wSZ1yUuyUvkGkKAQVKnwHUWhgReVryKRW8Lyy3sUfPlX06oChKM+TO
yjMljKt0ukhQ3JAlUVPHjnITmZntlj5uaMcjushqMRzT28tzvIWockFA18qn+gafcenD+ed3h/Ql
xIpNOLCCtev+HFj856ZS88k5O8N78xVEF88gz1I4+Sjxn5QrKsJxu/dt1rd4xLhMTGe3Zb6MVTAA
vxqV1gNdKjabCskreuZfj9STEqv8SeixGSnaGUY75nYPGuZQPyHBVpoHf0wDuc3lQlcucNjVE8Mg
nXBzw9rH7Dbj62WC8BzOBONjoivF/4RAQvbqycXW6OrbbWxDQNTIAtg2FF6t9K8u5Lg/zGxJUVpL
td32KfD9scasFC9IqLVjWhq5kgl4jq1YKZt9ywFnTBVOM71svkME9xpcXSNITxL9UPBGrSdkElBy
2gT6sbbiM/EUwdo7CxsG7Z/P5QPB/wTwQ6POe030KIuDtuui/rxCrAON37hDz4R0Zf9eorvBCvgH
kdnw4CD64m6xjkKNl0YUva14swfSAaubnZqv4+XrqVJ9oTX+U5gcDML/7OnwuTuPQiWb0Xj8+Lq9
6NSd2ZVdxl64LQuVkOBkkC8Nd+wEO26G7U93LMFPbZw00CzWVY4rRVl8//T+vp7nRJhBPRuo59mj
zMjrudHc6Kx+EEhuzqYj6Wl5A6R0up0TE1m10UaQxvtDB1/OT3CYC+nMTtBEUlScNnwATRnR/dB5
8zssvkqxPb5KHN/StI6jeU0mx+tTj1N2d3akCNTGvVBtP8/fijGuCbu8rNMt8tZx5ITOdqrtpC8f
5TK/C2FWACqx1z0As0FrPT71xV8bug8hevmWkm2hIDatVv13iwI9uh7OnnvdM+TIgJyTABBi6NO2
ndWcgwa7bZJiJMOgd/tR1WcwqCQi6Rfr/zhrrhx35HxIs7IC/y0bfSCVXOr6ld8dhPFUi+eHudLS
HGm1v3pz5gfUORt2tDrC5s8S4XcVbb6ABRP+yFlev/fPiOs6P036m73NoKii1NCjuYuZ7kSADXuK
ndGrrVbCJzaqRoPI9Ojvlhn2NbnZDfIqxhaK7etnXaV9ys8WLvB11lA9FABXnxB8ZGU22r50EPra
SDjslPC7jltSZxp3IYui+p5P2QWMP0mQOAaWcS9i6pKOJhTSxx0qrJVuVwlCjH6nGwMq4vnRq6yy
bidrRTSO5UVGB6YDnBTKcyWmY26M4Y3C5gsDFUOZ0I+OEHqtjEXWJAyKT0Xf1jzq4rR1EiE9BTzI
LDpl/Pzb4Y7uSGaHx90FogUeiZHZM+AXrfXYunuYzrhigEpl1T/3ih3mBT0eoNTwtVFkp2ngH0my
0I5uO6d3Eijh6x5HgVXI1uZzfu0XvTLC3+/zRTKW5ohTq7LnuCYS7XMVT2Vvhp375XOfR6hGER5/
Sniy+8oFlRTqV6oyiBxGrwTjh/nvsOo/dDxqaHnifSwz5DpGZrRNsDoy24Cp5Ix88px0/L6qnWk1
K3gWbMb8dPjIM1kYeIzYoJJyVj9OtD0vaI8SiHVU8gbnHqAR8P1bJmaXXVohZN28E4Mn/g7jy0Ud
cyaoXoDVlu0R4ea0Sp8DyuEnvtN+UPfMp6EOYCPo/sOyK2c7mKjTRFomQrxV1FsWtOsn6IN0Em7C
UPTIPeZtIh6ygSwj2zT7oGc6tDQeL+11hx23Guz49DG6QKve77dAPXjIRkax3lrj/lzpLKtB34FZ
qbnRA29zbHVGl74l00Lwa830xLnJfhsmj8qwYOeMLvhe8Sj/suO1myLxHcbiV6o0p7khLhZC7KGI
dnl7cZBu1CJl0vPvFDmRZPD2yBqiUO2HbbLlgRSx3loEm+47EXX3rfioxHsxiNcuuWHYrZ4WfQGg
IX1dc/XQZfPh7qK78bZa2sH3C1kIpAHfcEyDeWwhPR1IohRp2LzIQ/g9zLnXWHvDGgU1GjzRbpK5
k5gH7slm1XYT4H8rwJetMVZmyMXKdUWazaKXcJz1+1SuQRESb2tRmMb6ihG3rfzuD9ZX4MtiC/rj
kCUEpyT2OuqnzaUspHWhzjqPQ+uHxeuVuYY2J2/83fx58IyiBLOwJcJR/XTbf5VztSjGyy2ht/Mv
IvtnBBX0wWwv+APwybjw1II8F1AljdtJQiEnqddR2EoELGnV0ZrKXY+FNaPI42egiQsCpzn5CFp5
5CNTYZqaOgFt+8UoHFgF0CUsad6HswKhP4Q+hamVxmrBe2PoobxQbl8rp5bjDSEaWAJqQYqKydbP
aoubOKPPzEF5NeKZ71KUmQ/HDraG3tra+TcoP8uCMxwfsJKakTuJ9ad0zizCtIg6DZERPs1sno7K
akmnL/vyQ3j2Rodtx66nNW/BaKsKW/QMBiIgbLwc45DFOH+9z4QO84vTZzv63TnS7dgNQ4tkQcrm
wLfY/DBTXkOTxnyJQiatZFJqpoPX6EerWiKuQFyKFfwUwOkrQ5/P4VxRsNA7U/zyfUvXM0a4ZVRt
UDP6E92+iv/rdMjTuLugooebGp2kg6pEXA2dSU6AN5nztwL7KG/NZZzWyx2CWFXLkwzjXMDLnwRo
nPU1ky4B1kgWU6+4kZMBBkCZZSlZ5iKao4lL7cy3OUh3U8VX3w+LLk4fXEpi06uo3xl2kcYRUgNq
tUiqulu9Dg/rM+ySeuyLShkhd4Y4aaXJIvo2g5qspHZzsDa5Pphx5kBC8lcIKXFl3a8303Ho01vp
+xlnyZZKQlTbE4SCQRaJZHxvYwqUGuYkR/Aarnxb4/9ENyLDP5cuLYjRwsrqlMhOI7c6vdheAceh
lQrUt8i7nJJ256jqvf7vJ377Cy33MEYibZcA7SMzSS3kZOaAVu/+RR96DWNJD9OROjkLh5U89dvk
EBk4Ne9JQhVxiCisG6UYEDVxyTUq8AgUGJA8Ozzv0MH02I9gsiIgyyjj5RkojzDOMW2t+ZsdfzfJ
bx0KBtPKM96rOud7nX7AtKZMX4OcrcNFKW7OJV3N5xZ4sUzq2i4EvGv07QSerDz4Kv5msNBiu/mK
x96JwSIgyQWTM2txwSW70doVKMksqhvjLUC0BCP1Y50RCCiAfdv/XJ50iwGSbA5DzIXDoHXS2d04
EwZoTMQtzOayW+Qr+VpjVaVmM0J739UnX4Jq4c0kZsljAnnDuCRIuCSzxgCgNwM/nhQbVO6LcVZg
U6wUArCkhDVupsvca1L4/tY+3bN88ctJHih1TBs/KdHSxKpMxZTzuGwDzSAwevN6Q0V5IphsJT0J
KR6+KEUIWabrPfZy+a0+ps3C7uTLlefs9haC4crRFQjEfe9QYonkyYecG+qUEn+cilFAPCJ4MTAL
YgDFFNWxAUe2dW7unxLYwZfT1qjtciI0HjgSbx8zEVU1YeU6tpCrzOEDQbxBWcchhX8DOqP7FRos
BmX9Rfz/ooWaDYDwiKXVxVGoJloKkRIdX7arHRf/h6c2JKbkDVtn8fL8gCuoCpVFrYScK1o/NRWw
Wp8h0gI/Ngc8ti4s03npA9Ar2w/9AcdLS5QGV9ZU/O38bl0MfdODq3ayvxpRpUsdhTCMJO7johw5
CGsQ7qnfqAI2HkkETTabpJ89MIH14VjvJqT+4DmfvUqRVF0mSHSiCn7gvfDQbdctb+x+Lvp5gK14
vRUb1td2EOir1/Q7fgC9GgdZuNiPR25rgAogfqbJNCCtKVAktaHWCXII0jX8/0RJzt6G96VHD8rf
mB/xpJx4OtG2tJzT0HpASXYFcPqJNVH3iksPFJkTSB7YvtpqnvFbOVOkPf4jIVjNCO3vyPI0G/SC
JcqsUJvQZCY/ZXPsuITOpxarjB6pwKiRayf7YPU20z+zB2CqDgGQksyh3sm2QLJbvZw4WhMm8UNl
rTPYU75qyuA2mjc9eHKoJZNwYH3WRGEuVBYP9fnRixazGhf0CGVoVcNp+U0zI+cYllYyBfhM+xSX
t7Fjn/OdL8LAquE5nwhnF+MJPHziimsa7zvuZW+rScYG914jTcO9vj3urplIL4RwGaQMsU11rxCV
MYvuvuJch6i3cY3DHnjM87uTL3NNUpi2mniHpdeSG46TQtfl54TTtIeg4ZnrY7eXxsr4o7WzlId6
NlL5eTCRYLJ6oV2VOvdk1HMFhGYrbPVD4KZF2y3+xvHaIEXEEqGhx20m857xhE8R7bF2CwYHOZ3+
iwwoTHcfncwJbVpyzj5+YP5YFxFNHJNnkR6K9FVYboiDgGP6M3RXdwpnMjV1j/9P+ds+y4us98Hf
LaB7uxYuppELDjclI/gcsocqHq0CYoOqMYpcRYpoij3a3yH4X5F00zzKqlfoXErkvCluoixPuCfb
qUg5ef/6+aY5h85v8RIW38pjURR3a5csF6voI+HftukCbRX6pQQFRjpmWBOf0QDQRE+JLR6zZ5qW
Mf735Ap4abm+ssTq01rcfBUXp9HhKA+FZRa6ldj9B1TIxXDchCXfHfdA2l4E43aEzaL0mqaxuklz
S71H/dpswFylGRIi08S4VfnooYgyuhykNjpCnfaohREpM+Tia9a4jbKjsLqIc7R4Xq4MREw5YuVw
oKCocDKTfknvC9RlKRNiN1hrMA9L5auUbrB4v3JEc3TlSsyozY08FF5v8VSwUKCAIcS5Cs8HdUZJ
Rfn2mj7+pz7OfxFOFxCgs0J0WVcYJmPf2GygeXUeUq5XayURD4J8wWP4RRozjTyiS0c+PVJXwH7u
cn6i8vBe6BfKzwHjKkUVu9Wb5G1eUN+w/byLiL+x8XCyJOB3InlJeq6sseYPawVt7BHroi4NJBRO
3JZoEBclUJDc5sibX67Y+VZfAxaAf418KnO7DBXa0PaJQSiKRqG/4Y1GFV/yZaSyF93OCvxFppT+
OZ3OOeHUBBkHQ0pysqI3+Mqe3fVIO8MO1q2xKi0WCN8SoOIaQgwM/kIr1y3BuI9F/ys7M7rkeuzV
npvfepeFfgCiE6Z3f4QYWhomPSJd9M7UTZN9FEkDRtzRxTpJfHa8xSqVjQ/0TKLnTzqr20RWcOKp
jnAJlPBuVhw+9ptKexuskf9l4U75lP5YvUeTtBWqIFGm5HNOwfIW4ZkHmzAzNAmQisuccT4bF1CJ
L43wwG7jIoYPHUkY8EQG1yiMtwk9zeDhWJsiweLHz2haSzPr4YgfYRRPSjHov3q30CW9v3FQDjbv
g8Ps/2Nq32J68dDB3isJr2bgWeOS9KBwTyJjkvwnoguF8ppcFCxUqaFVa+X/ocADoujQpoqEPviI
AE8fwYcAtFDK7mp6A0LgNSkSZdnTu/nWhrDh2Vy5go+ehhtT4ba/i0mQphQYDD6pPKchNDwYGsFm
k/yHC10W4A/+7oJDHY6RWc4FjbZ+TRH/apW+b5rCOYJu5gSl+wN0ZXGNSgXD5ZXEA6+Z8LVjtLHW
TqPlj61lu4ulU2uJBqQ+/BYdITiqHqtjdOM8RpU4u72Z5VB8eDJwrFseS195qsqJfDThbJeuYa0O
fFOGLfiw4oB0YKlee2+nICxgWsTXVjwoXy5Q5odom1CvpY4ewGK7qaGMLP1DtualZU6hjlABZiLR
Xr7xh15ZQSof8fciTtR9YCWBh2ahx+WPlrxtVwr9896bDBt+6N5S2babaW64qySTLzpDpAox5jZu
nWZxR/bmXrV0wolmFGTT5NRcjRRhrmyYbNNTnxE5aAY/9i54Jk9AbmXZ2ECc4knvTUP6ii8VOk/u
sQM1vY/Br+8nVthVfxqGPUoumV6HQqwyJByRkyeSs9QJ397mJbovWZu7paivTrSlcxyJeR/FooYw
QT2ajH3oe3qytzdUnw27++dAnpht11Go+c+dbqUukZQ/EtEjwAa3EXm3FS1l3pWhiWUyQrL1cckG
JHT+61c1flasCFpDXIrSERrbV0ssf5klNgVuFPugFPwl5KjX081vqcUuU0r9r5V1z/NqAlFS8zyb
H2QNYGeF+4x3OMXs9/cO91WJfYE6XFEn8lZi1mLNuXGlN7YAFrnBQfkDQ+ZM0d+uVIYXFGWI8yXa
vfT2vtW3ecIfrQOTrUz7ay6Zzwqd5BoJ5rQnR65E4b8eCFFH7SJJE+j1cQZBtZ9aVwXzEHdCcwW7
scfkh0ce7CxXkq9tapUa9Y0gg3yGFAB2d16PkZiXnR69I/4RUaIohrnNRANMamRqPJWPQ1GRv8jv
sZ79oNbV50pDbLWDPhNWpIrxUqv1IE0G8twT9ECxSkSFKl5xGuWBCEVYKwFEQ+jbwJld0W9hKBWE
1SKMGnIeJ/j38kinEs2jpAXuorQwSCqVB7RuXUHW09fEhdSSjBaLTE495NttgahaZBTQx/rsqZ+/
lSmHv89Cx/e1a5WQqw6PGu7jFjDS58Yy8NCjrw3tpAPRFW0nRJSv6tvRR5R29YSz2Ip+bOwyfWbS
L5Na+YlXmw8PQSu2FKk92Q0FeMLBfMABGwYwpDlkVg8X/hfqFOuJlVE2N/KUTmQx55IRhW6x7PZI
0ORBt5bb1cuWCrINJ/r1TzhWoopl/JIYGNpL58tgOiY/16xNGPic1aH1FI1Bpmbv+IYqOS70nNBm
hQUP8Q+9LwWT5+JDlofhyg5ZS0BNtGJ7sgqpeWKZosSyr0lefE4yew4rbM5k93xDWPbS+P+NRd+n
CHLBsi31fSqo5IkFLltQ06jyPt6Wn2sonZ8XXuYmSRZ63LK96iJTynI5AWIbS1EmfzcVDtlqt0P6
Rzq2WQGYmLHNMs36tD5Boym8xkzShG7miPwEH/gIh/07CENv/Dl0nXPcImRTpZ+V3+i9efAP1aPj
Rx8ylBSa8dWa5w+fOtAitZ5s1Ou1k1HsB3X8CIBNNsSR1B9GaPU++9ciA2rGT/ml0zFpwsSWISYt
M0rOjt9mktpI2QzXj9CD50qv31yx9JDzjwNMuRRF3BGpnO3puEXyZHYFjcIwlR0zFmRnPGJ24wkq
1q+rr+KpQ3DbWJy4Spxtmqk9tnCO5WBMd2fqf3jdo4xnM5t8T//pENRgLgwkOI9n9b7HKKrb0/eq
VF98VpPIsw7n8bqhxq1MUVEWIA3VlNobohZEOfbV+l6SLq9qRt24xGllEPRTrXwwVuCPwU6U36KQ
Xxe3rWaNerajrsNlqv2CVdY4PdWwZz5RZ5xKToHPoDDmrbZGrZvLg4UW0fnvSJrmF0nSFzA3pyzO
bSRCXSTiJL8B2w4yMW1Vh6cO8U3SMKonqHZQBUSoHGGmoSjjdv0WpyC2UgV9DTBAGZONuR5t4KJG
5KyDKvrGfcPrkWf3kKx6fVxp+QJT19uPU6hJz4YgR3T4Wvmp06Gm5FBI/BUDOvlBZer6GMRVq1Lv
Eh1/si+RMMetUELF0j6tmbeFHrhZM6i5F8RUX+1jxP1TIAAOSZRxV0zSUrCJycQW1Minervdgkbf
p2ue33MBiiyuV4GFPLtgf1l9MwZ4LjoyISuy7t6FqG6nG5b1V93oNRi6Ue0o5yOZqNZb9+61gOpD
/xwwc6DZJ5VK9tTWSRSzx+BIUJB1jkYJ/v+rIvUmnykPE06PGnr7SxglujzD0iQVnnD3mmlQTyoW
Xq4DtpEOJ0+0yoY/vVz0VvXRfcj8Toj3bqXofQa0KHY9klz6RdqjCRYR30qYHHedYnDyoYjBolGj
xc4a2SUXAnlTTvkmXJuRht7VOBOejau8W4+qtvIpBJYwHsujsUCEDva1IUoqJDAOi3Y6otoOJT24
442fcD8Wme1fLKiVJLQjKcHS/CfeUVfVZVEDmncR9NRvHZz/GOnBdBQ3aErzqwsaR2VMTiRM5Snh
sPWJCGz4YmLzr5UpM4Ukus6w6F4ZXQV4ky+QSuU9X8lxyrLfNQbyAqvAmW/s3b5+QKo91JlILI2s
biH33zvHxfOiXlr/2JPQLVMh/MnE/yRqGu49LmGKNgplbBXQ18OXLh6js2caz105569Uoztdv6Li
oq8j3Bn6LES6rPMIer+2/lJTquMz5NzK3M9bAUjEKMnrV7LWr7Qw1By89GWqUGHIPv7YhR+13ObW
QufmPiDfUhfweIV0n006NCvZsuuty4l6P6PwUmd4QuYtLP3ZkzlB93IVlSWbFOIlch4XyB7dMTek
BTbEL6bz59BRBheoW+vac3sXUCYYwzbfxZEs1mNfw+VghD/IPFerd03lF0VDbkmGE8i14+vOA5jO
WcmaoUb9I+TYnGbu25UCCS8IopTPo4asgjsxD2UDZ9c0tuLFtKFCqq1uNymNnt6Yq3Jj/PsBdLss
DZACYGxfv4BZT98rJ/jAEMDpQZqv+/MQ+zpf8Q5EfRuei9br+BroVvbUTtUYVwsGzR76O+Sd04yx
NV3As6iVqSPmxa17CCPR/vCNpwlD1yIRgya1xfG8rXmdl98cl6B5vuNXFl1pT3BZ4Nk4eRkmFlZ9
BhWmJSFtmQhUkYqun6nwpoQJwEHfYmN1cCG2MV4bPmPnFRGBla5vGP6pPffGypacYOiV05j+MXn5
OVnpUf5Mugb5XjnmkANgyCTZ6KnMxfTZb/KbJ1KQ15KkWngYxt6zSN0yppJ7zVLGQcVpLWKoyl2H
TFCiPVwsqWUSD9FEXkG/ZRuzUCXOVxF0Ux/RDVdW6FYULFcP8SH+7OrtBZZpw8DN7KpcXXj83TaD
Rudn91FhscSZP6w8yeHWa3cx8OcXW56D/y0yHx2JV/pCerZPIHmclWDsMn9fZT9ugzH7BkcT7tiE
IP8Haitct1Jc3UCWx3WFVMFN8Md/HYWWt5BFeFapu9js4SIbEsIImVfJYn3Zhw7ZzYrdmbIiz60q
uruG1z/ohAqvQJ9SgF+viHeRJX7f6AwLPjXyNJpY5ynZuX5p2b9i+vI3oOuILuYyH7hvOeLMUvB1
0I0y8/1OnAQuYZnhrg3Typ+sBF5fu2Ad2em4Azms+uAEVGVNKsNYex2JxMVsiF5EFU0zCxEBDh+M
HGDZuACYFR7h2VZuPZak956c7sSfjBj4f8psI2VWEXF8CmhCrm+vZcB9hCaSmhnvq1gUSp3e9/rM
VbW2MvCNHortW+hAIenSvNitp+wDFpCIktHOtLm0HeuLBQkcmWBnB2k9leLUr/4euGAwjifTpIt9
qGH8S77Ar/NvvmDgfzsVrW1Nd3IfJTAFwAkk9qnmQbrrj0p8XsHo8epIa5JINr4Q9KNWGx4OPWQ/
7Q7r2Oj7STa6qqDLPvm+abKiFXD8kiY09yU75MpoEXp/969f4YXIBUVPUDbeu87z+rN0bl7PtVEd
G0vcHH4USsc3/iFPDVkQAF8ED/0OMSSTOMvKXL8MwUayxNU/1wWTjs5j29Pymf9kRmY0SgJmHVSy
0jJRzo4J6aYiI6hzbjKA9z9IJRWXSkk4cwh+6xGhJhI5dWViSgiMMUIEd5BIVb5N8Px/szTQcHDP
79G+snhwo4rQvseUXMmgei1rmOhwnbkUNI/3ZLkPL+GJgPOvc7MI1X1qcBuDX7LorzIioOX4v1LX
PYby+UrujwTkz92tlEfOSmrlAYRbocb1OEWryTo2PRyhdOaatMsvrvNuJ/TvuLGQoIWPRI1xNEFS
G5W7W9hpAKLFEOjpLzZJe3Tt0MxNaUxdJaqaKGW3+xRVFVPY3agkVTIeEQStl3FKidGQzxH3tuLT
8bvXDU9jPcpMIFjUu4MI03t6t2xqCfCDGUPO0fqQzuvd6P+dw1RthYi860enttN4Ti8BAyG3QUL2
S6SyDNTmt3pVzdtQQ/+KQIPmKTxVjtATmWTEJ9PITptMqISiewjepyGLu54hSpiJNmXm8xEfg+BW
q+BNb1v26hNwWWUa6aXhkiy+qVhAfIm/uyOOXu38BRLy5kIzOyULJ8hvWi42j/R3wVoQvfkHksnN
us5tvHtRT7OPtooqSzkslK/dixReY0jvuiNUT3gKJOugdkWZ0ODju3HsS+RcZB4wrhwtPCISSOQX
N1W7d0xYbCREdObG7IfnXoppttZ/LbEASoHnvqxxa104ROMOUXU8e/Zl1AF/vLOkdSBlcOUuSKAX
NEqQ7TBOr290EmndgpI0ElAJGI1ExqjCj0KHyr9Nzj2UIlOeKw971M2I0O5Hu66HxsN2aLC6SSyW
B5pivY8NonzbDgKF9/6BPAUgYDf8B80L6FhkZLUdETFWHjcBik/+gCjVFwxg8QlRxXGfWneufYHS
Ne/7GiTQM1s2cmqk8b1cCwTUX9G7zWBTmJPk0dzm+qaaePv3Cd9T/GohkdZ1QvoncrxNu8jXdbZ5
NdiA33/XcqxNFfrgDaH+M3UfhEzRvKvm+21y401d7xPSQRlhE9rY30B2/dWEnWEhWP9ex8UHq0bz
yc6QsQZsfMCRAOPcwzBDEcgsisjpOfBbR2u7AXq01dhfYLvbn2Ts0dUxKBCpIgDBi+sPsveBWbZN
CNzEOTF6e0Nk7G4MZJHx9iyiF00HNrxgJXtm/JJZvWKhzmZnS5EIeJHoKNGRirMISQ3cRjEGjfU/
L0n9Y19XC6CFEEWlsF2ixqKPWuIHHsead1lDvi/weNbsmB6Q7tyaIRFqLEJM5RaCrmBDFrHDPV/Q
Wl2hurG1V+UK8+LnPxnEpCBi2gm3QCGwQbhF69KlmxHLktm0VcwSRwR9xjVjKKM98uXzgMQ/Fre3
3nPXmu+Tv0n1HiEj+f9cSu/vGejUXrjLI/SWoZKliGmLPxGvwFO+97/oToarWUyZYDQGqeWxfvkm
T0nDMF8djFKTjCF7uAyfi2lkiN7o++My5DrqObVGQeGiv3EEQxE+96gygEGAw+sf139i+RzuB3T3
EHpg5KoAwKexpQmYCtVtsAY5+JxAfFjOr+lWQ5UgqC9WQvW0wg8wvLWV/4D0PqKeZkR8+o0vYLV9
ir6oWJ7LSWrwX7VaJ0wvRULGJHGPJe1F4Hhm/zxEaKoeRg7PS6F7XI93NnEY7AQXdX8yvbHuVLr2
7BuyQD0rsfvU43+qGeZen2is3zwQofAKloypM7oU1iIdDUH6a0Xb79Q54nS+KPY1SUGmzHgRWu2n
B51c46zH4zAzJ9lHbQgTM9R8yfVM8t+sjSSm53Vgu8Z4UO3il/KmYt9Q4ynq51VJ484KC9ECTG5s
ZjjVjOnFXwakoz7jVFxvGTWS2kHO5GRHCWwjw/nv+IHoTLL3IAB5/JsYGT+xvdXdPxnU3BjLizr9
GV4nOC+uI6ZMuz4cTZPRQ/DtfP8zqANPXHW3mWLMB1yt+wZe8miRsT3DfJpsuwHeu8mLg6AUofQJ
gIRBDZzwIutx/HK6kzklotvD3taCskXXCso/h88BcJBd4W0+gbZJFyzgmMFrsqehEokKpKuucztI
67oPSeCDmV9GOZuXqHkEmXb/44hXomDStMQjnxwS1xp7Jo0//iIcFhn67lTYj7F21NcXba/pXhDO
xpkuDz3c6810NNtEniM930/hb+ah1Rn9gQL1DPeuODE2wAD1Bts8I+K1ZQQPql8I2c8xHeTAKWLY
e3ddTswfnMltBtbXOJPlPaI56SOpUJXmxP7ETG/xrL0SQY6B5ENsndOofIvWg2A5h1ERfk+Gc0mJ
sb3pbzsgVZAbbKQ3z4cfBw0AkkTqHGfEFfK95dIVJOXvZDLC3F3Tvj+rROKlCi3XNOVjq5YNMnTS
+AkIPVOYw3pVNeNBibyB6R3l1tmC7r8pA7/hczgyDB80kgiP6m52Dsei9i6o/Mmh5A27qI11FjKO
+MeUTbLijCqmYrT3iPAlENoLUvvbxM9DEUQggHg4JzSWVT8NywzIktBt2ML8MQZmHSMXQI4k0gr+
zsmtO74Y/czWjlm0WKRgCPbAX+RPd9yC42qf2JG4SMq8ycVKdz40rsWyE6tT1J004UjzO6ZYJXSu
cnlJV2Z6nc/T/FBbGxHQxhOhB30f5KYqHKUmfQZW8d3609xlWfQqW0QjYFNpjYKvRAq/G8UYl1Ib
V6mP3bkL5jpJS5qQ04Falz+kgB4UsCyoOFCWMgvrPiuEK86GMAApRA/yOQ8qARX/R8ukCyvnTe9p
3689dGgcW2q1WYzA3zkH6H8X2OxGrzuofh+1G+jyMkL8oe9LhqyPJKBS2ue2QVW02ug7CAR3eEYl
Ug2bYmSk+Shc3b5WMgoZ/2wj4KbZ1FTtVANe5y4Bz+fMlkcYXGMJDHytUabYsfFcYEo4TXi5kgiQ
CpTQ8rLWKyX4XGRgTaDJG5ufnX/mcCdjSNT44gMPzPhyRvsAA2Te0aeSk/384y19NFCZXyUu9kD8
J5/Gi5Uc2aIxRxVgjIDCsWP7EFloEceHLk80wqnRyHheq5k+agkM2EWGDzcpAqBFZdPHr0P9bULR
pmr6ZYELeL9UaOtfh1CQVvVMShIUNBCXg9i/+vuEMPb7PKeNDAnEqiz1Ln4DZk0HVzjKl2HI1jFy
O+xvP7PZ/SdWYkVLZYdOqle8+bCwzHQec3C9qL2nAnUkkAOOLX+OaV1vQ42PnZrU2EB1u8iWi1xp
p8vR9JIhUDD8XNk7MTWNC1PD4BLL+razHM/T+ONQQ0Yx7DuWKsUUefYZGt5nqQxwdZ9Lad8iEXZ/
UVezUDV04laV2vPyDW/g7oPo7P6qDcmwRKR+kKzcsNBi16hmBZHM1IxK/jiQ79tsOcAlDdDuucZ6
b+m7WZmD3I3h1QzBds9QgqfzEKwFUkD9+qAWOpgJFwOsu5FmClmi4ZV5M+hz5BitpbD9EJcC/kGi
bleUr3cmDlZAhVfCVTgwo5e1+SPUCg5AP16PHpPLvbvcqmEKiHibEQvOtfQjAduwwk9BG6TWdn6r
xEjyVYfskwY1k8syo29rzl/CDH6ivKBUymiyH2YAjAy723Ysvs97NXr3FKug7ndzvIM2xhGag5JD
cBsSnovv4w71P4wZZGawlTdvFjxLJZ4HS6CPFMKqKQuvh5ungjTu7utDPLHGAOxN2+yiBLblMmqH
T9rIMEiIcT6d5ltCJuNLrnk+w4d0ivI2MrJxETilM5xfoyajxlpwnp7h3weDTjufNeodHqxhcYvW
R8KpH4kMYbwVi089Wn838LXKBr/CUFwgo1whmWGN0sYtx9GhUn8jMeC5aYduBDGeGMdga7iPeQ+b
8rYzZZ8TRGHTYQpnvrIUkmkPQrGmKrGmQc4EDokiGjcXSh1NWTXJG1q2ZPLfjfBZs47UDNYt1sZb
pJEy5QmZnK7Y7xIzivLdwUlvm1HOIb3VVCC8G+veszX9+8sB/cTAb6QucybWB9BJfaqw0xUowDTW
lSMGOB6hFRx7u6sGt95wrPGsZIDvYCNBiTtQ7SvQm7Yb1qdrMNxkhbcg9GC8p5IdJa5zxal22A0U
6WRO9Ow/SVOhwy9w1zJuY+LsLxM9KKExVmh25X10YPo+Lz2/MD2lOooJvJkOIWSeeyUHPQ9YE0iK
2nsUkDGEUbVkYfvebToez1jfDqXsEKxYnYDluLuWsdosnXxZ6OKVPOBFipIyz5miGGFCzKT0tZM+
GNmLP3FSB1d7lNBu70s+1ClY52rxMHoovYk9PoQMj5fWaF5sKEfAP42K90MH6NZu4zXd2ZuTwo2y
q/8Ly5E1g1wMK3qqonbokS+pp/PoMKP2bnsVvKh42OUBP4v7TBGUU5u7KzmArvZvUBCp2CtUEsQr
Kkd8CFJKv/mti7zO1p9awHmyaRRjMPelVzNe3bBPrvtDZ6huDrXMwI0s0m/J3iVGNOdm1GOUuXPX
wBNNr3lfjR+1YVPOPuo9HTG8kUaX1xyqDw7sqGrpLkeI3tUm9+C/IiIz8Tq1CI0EwObyGFMBEVWT
SPkClmRKu+kEwt+c2m2iCf1NCXSE4sVkPeoh+R+KSRqMwJHLdk7+u9ORiJ4MBrJGnpxG7NQwHnPv
O8nu2Ju/i2NjZp5Iod0rsiRN3ah1ouphNd59mE0odWFeMYZ454O2t+DCxQbd/7oFHT01UrwNuHR8
fLDtRAcXlG6oD6UEdBlvYXcerPyHQbXMioXzQrLT4aDuYro6YXIXlj5VeHZI8dtVccRV48KunWWd
RtEx0op6RArcMNZyGVRnrdyiwFdy0DfNGBLx8LRKPSV0ATEoPkseOBZcSj5/0CZsoV0og5p3nPUi
cliqOvdnGdqSh10ZUVXRP7pf/K9KNCwdCZxirrsE5pzdxEBgZeWnLmW2n7FRHYmKMNEOJZRmpkXS
F687b2fEInZwVO2EIK6JQpKNa2JT0fJsbm1e65YWCc1xj3iRpR8e00Le4iKkNJjp/nXqMMlIA2P5
EECEGV2veImJwTuV5CgE3us3anRdK0H0SdcwmfJR9Ak0IVN8jWGxcePJ0QYXvJmylcmp70KNgzc3
8nLav2SEX16xg2uSxv0mw2qSVPJJHCGHT0LeqWSCYOAdhmys6hCIGvq8wJDgnCDivBXrrmAVCq+B
ylPWTAIkIQP43r0DudpEDdBcqaw9tmHAgrZszyJWF/gC1HM+OmZBwGYXj6yXSpRlJSEEu+MRNbim
fxFD/wQBIoMqxwkhYgh8nIqOGeX1F+sTNIOjXzgrl6I9V621WXKyAVoDWP99oF9Wu3CEUToyTjhs
M6MFQSoHhPh/Ru87+tQKAeyHrNezma6brMUM7J+XdXA2tND4iQ+JJrYthW/z0SUdh3hynsSNk/HQ
XRXkEmzVy3Z1c/XqqI/SbBsbau2+I3Awaaj1UT8J+fEd2wsAIoW5RxEEqVOAQuePgK6Ixafdt8zw
yGjUT9EpbDyknXecO/Bt+7kHpIBBy3D89oOvWVLH68Acvpssu8DAzZJZLfrAkkQsbYNExOgA6vOS
cTMsudob04Ch7aEluhld9sgLhzn1NwR11E1CwiAWe5NdJTsqVvVvI/Fs5aG6f4HbAJS0ldxIxDzv
E1CW+9mDYc5xL8FyBvLGqLQdpsVag7/CA/qNYn9fiFNxwPvPquc3bajdqQttZq4P0jugaq3n0Kyw
sL7qAaIDTNrAA1hiaVr6T8EjzTC8yjIw2e/rXqzEwP8h/8a5rNibt6Q4JYC90CafGDzkUh33lJk0
Msse2cec9FahnWM+E6Kcwgtf/q7HUqGUO5CA0qlf8QNeVlHSNShWMq2K7MQxbgsuUoAZ6vW4s1Cm
C3PsCAve8dCYaYP7TzDnmPd/7+jk2e7i9CQQx6OejLC0P+GpyDlfIDJmhJiAktMRHeo6Xxkjh+Wg
jnJtScGm7LIDCiRk1tweAifB/x8iCLm2OQ7DvpRuRrgg5vVaOLbTqsItHxqK5plTEDphJIf/t79I
3NVtDRrqnpT6UbI8OM0GW4AhDTVI0hGnTlx429OoW8Upa76rIv4s4fbxzmNxCQyL7EyPH70kN/Dc
F0EJe5UKurm0OnOtfM0nuJJfUgdSKjFvWhOlrq1URULE33lGv5TjLE1rrIkJCRjDBbgG1UgctVlP
dX2bGzKEDyvhwyEh1sC4act5phT6Cz6UPqP07hM8MSxK23Z2TUWVcqIRuTfGT2CC1RSBkz0/2WMz
Dl4D9Re26/1E1Xv7odnWBxGnDRyC55ewCJz8p9KrGlrZUNpyX+fejcp7t5dua0XVYmgBHuY23tEJ
zjQNzh4lQWtMm2aYv3W4cpJFZdmtHRGqGUIG34B3PQHN/O0GKQF91fNLA36DRaIZtUs6r8rnzH4P
Bcsj473mQSS8hldx5qrBY4MnAfruJBdF9g+fxp3IpcnQqum5OFjz6Qf/J+YLn7EmpvETjbOc1N0u
OgDpQTpI1ddFyoV5uTVa7SbrCBWtRo8ZEAxJc8Rb4eR9bYK3Vpb1TDJ+3Mc6Tm0oVgAIaAtKUR7e
LMakgKi7mob2VjSJny+KSy50gEp1Y0QVqKHqToSDKspABEwVptzsEmLVw5gvCEF4Rc2e7Et7Srkr
w0/CsgI2nY4uBkqDJYYE098tKPw2S0X4GffkiFSTlwlX1fAxuqZRKC61LqYpEs9XTLiy+/6yD7Q/
kzJRN+fR0vZntsJQeAD1+/fUhkZe6AXFJuyfqXdN+nimJyrZnVMQKNUiYf1dWGgm5X4TywPvt4Ms
IsBk9RwegIs5uwD6k1QqGCxwfh5txWGJqt7bbwNTs4m+BSscikJXC818tONSKSsb0SCldESsFga1
2QanlNDJCabRPHaSVgX+4/D9C7LyjC3oN62+24ELwNjIaxCZB9Hm96GvUqWxMs1y27GWqG1sP36B
UQT71Y6IpWbyQv8ldXSW/br847e1QqQeI5WmF+5rg5O+EW0Pn5sOveW7MPq9gHSuUBRSWz4jU9zk
ZU1SeU5JctBY0TSYbvLJ9wz2CApvvT4vvNp+stQ00C1IvPCo53ybmu8Pw6NoAYwweYSNBy4+fu4g
3Xgmr1poUNIllVeM8XCIvnsX9ycLyI5e3jjHN3JubKblPXp42nWSgVSQXKUEjnv2P6VpAO1qHz9W
cDS8NIN1w2edkmtW1tsK3lZKC2UJfaVExQLg6c+S7T1Jqq/s4M1CdoGDSGjBe7pBBjJSuz/BG0Pv
mAKC3BnylUG1P1dGAmYSM12KDdBoM4pwUOBqDJ+UPrd62ImTggYP26Is1dWQEi8jLGpMnvimaSNA
nw3r+spUOGSbYKLeeuO9NBO4fzkHS4TnBasL58gpW1mIA+KjlvevQOC13vcTNLhhxE3ca0mOewMV
IXOP80jI5v3OGE3F3vSSIdHffJrMTH/3L9ohrjsZAFajiP2x3qIzF/vBWd6vKWw4wjVotxq+R1ih
qyc83Nzp31vrWpL++HrmF76IIC4o+oVXkuC4n2aAzwAH26JX/xc6WM/krYk3bSB51xxsjVlr0NJf
BDOzzR5HFQKuLwnka7LXZ3CxWuUbKN/9zW3HQIqPlyM0dyTaoDoTexihcWkxEg/mYlyAwYVdQ4PD
UjZAahVQVBnERf7k7i9gOBuqHyt3vGFwr++2YLXgqpIdH0dS9S68c0umD4Jyve6/T0js044ah0gH
qFQUm/jTt6z6e47VAH9bc/2MOmUaBnHckMWuOVN6/BiV0ivVZ1Vh4MbTkz0CsgyCK2j7oEPHqyqV
aVxX+QJSDfk8193b6qposjKtXEQ3RImqDPuuqSrW0cZhdOktLr0pchd64WvQbw2x+3xad7dux9Fq
idqCTxQ2/FfM2nkCEw4QhrdqMKKEjlULJQ2CsRQi/A7p3T93PdGBYAv3uw9qoATVBhlQTTsZu8KC
6n1PnQEPc5I5szVXdRoBexNKVCYyL6SMOR491lz31zYEsW6F+7qmmaUsPAXN/EXsmeiccA440UqP
H3ZPARREqNE4LcCb3OfSDBo+IqquyLC5PPsQBdbdNgoJ1kAbizad8a6YeEBVgIlwuQOyAkuy1gVJ
Umv8o1jkBdNHa0APep05CFT8kj06bj8FDx9uhwtF49ceLshUHiKj/b5I3UAovTDqKQXefAxjblOk
CGIEMqww34qdNsWk3WDVNcLlsAlJ9sjH7XFZ3mykpo4Kt50z1SIxDvCEiL3YmxpiRx7V/y280SB+
cKhZao5TFXhAbp58I9xfSSmRFJYjo08gPGgF9vdLufn1G+Q+EpVdA01oa1qbXKs7OLfy5/whudUn
IvMpaHFTuSXukjX/dRUOR2a6rvQhDE7kxT/mAeppTo11xBulW2yZqUWwnlQUOEkyIS5Z55bMNqF9
tSI+drMrfBp07nw0OfMddu6bgnzsPA/om9iBqenRYnasgR2Njl7HhDtpFwRkLOv0a6sRBFOE/p6M
wq4Js167K3PppgqjN5dnNSq0IAHVG9C0uEgNVbtMLe96GIm++xeWJGsavzW5w3U1cjl6/q59NvQC
4NOJjKkZwMyzjYacNd4F2EFlxaCFmEkB8FGS4ZM5TZg5qSKatUbsriP8Pj9+r8Oo7uVnfHJGYK4o
3/lcctvj2fcwWj0K0+BfiRGERKhWtoTz4k3Su+x7Xh/IZ+hXeQddbVop6yYuXdKnYYmiB+rYhlar
AtLriXlTLs09KQ7/YbKcyyoato3nldIUD7ln2avghCs4BbwInFXCgRyTXC7zPR+tRr/CSXaXa4wQ
9eeq2fuU4DAyvZRh0Otr+QhOMHKsZ2o63f4n3s3XPF2JApFFd8W+SBTjrfdJ9tNpJgbMloG0zG8S
EJj7+/KmD5QcpinvxvZC4fApseXIzX6E8I/aWPaO5eU24URX1GNwPLD3T196lruHeoayj/Z367X2
WSnWJf6bDTFMAprQ0UH5bPy7DBM5zaQJ/lvNt4HKx9ObTKg9rISO4Z0Z0WjCccx1/19fol/+wGN2
buPmQ/4Ff7MRPCCiHa/u6AEVpjJKmYy9PQqd9Y8UjYk0G2MWIDfzYmST2jVs+EhGlQgZuZZW3/pY
mWRmlJvzdwFFwN/6/wzypVuin0Hyna8wojy6j4u4dlB7Zf2nGYF3ogpTf/ZG0bNbreh3cnrL+WvZ
pkdj8m9EZnufpE5Nk0csxHjff5EsL1fNE/PcSBoMsDBCdpfCaeZv8iMjyh/WHyyoycQJY5gapvNV
1aFEoeoeM/XfBYRzC/wUT9J2+dunb6BNaHIA96D/fRbGlCaMBOv6dxAUF2GbuACMnOrSaazFYBMU
Fl87n/OzzoI1yiQra+NNbXpFmrwWYcZKXqAb4J0Pey/bWGEX7rPIW1RS1tiJLXXJeh19TChf1Mny
qhHqCjM2slVktze7MBQf/peQUxUJXGsrasYHIwfCGD1bosKFcAzAUyOOc+oZLfOxEHj0NbFCaNVA
gI+rnT5tSM0WtINo6Iy+AqABPefRUCyAInXB45BU3z1Pjg6Z/7MsQFBxzExCCecdkiE7np1VQ7E3
iFoMsXmxzgoGm4AFQ2y3+QfCMpQiKJUPYepqU62xVLgJkE000oB+AEpGv54LWDVaENBP1fhtFCKB
D12BO98OF49Hw39ZNd0vAEU6D5GYcv7e71Oq0AaokzNSZSD9YnVSWoXZDtJ/rtCrYbCAptSw3TyC
Or+BUiBNbWwJeBYaWTxLBaGzyeqVLCH5Ot27wA1j9XWsOmmGV6JsR7FsvmD3E4HdEtDrUrD0MqLJ
gtMo2/aTZewYBszWZO5v1qoeLWgn0nF7h9fV8ODD6auzUirFnAX3bk7vra7gJJKBOLW6J1zFN8XD
i/W+Ikig56bTbJu1an71ql5NyPVuXHiDebZRATjMcB4IfXJRtU081UWlbUi1Q0gWt7rPeVCbsyZS
Tu9eoTftlmN3yj29gDlLLl04PzZFzzwefTT4L87Mf8kvKrjm+Bvd2drkGBtryOjsqW2c9sKGAvys
OcvsJKRhcC9Z7gGE9pQmMeGQ3O8A/5iDT1XmuDBNQELCGzcPxkdDN/fQdfX1rUE/jciZsmZjYiNr
YWdvaSgYplU8+I6UUXxs7p5cmvv8TsyTD67+fVsGiNh7tr3FTE90yjYF2/MLYrCH9RdGvhHBRAbm
Al7v0+04l0BEbua//0U1x1hkktqcDn+3Qr36FVQsREIajqKA8X4buVshQkxAPbDrZbufnquvZCBp
O/+0XeMV/Kqi5vXziJ230nrfKG6OhdK5/ry/u2w/+qD8w0rw+OOOvDy+QR4Yl6jhWgbJQxpxY8B8
ERikihNgRmNNzZuAYkpuGghg8Kao1QxsHIzhxN0nmsRAM7CQ560GTGU5SEA4wEUaaep45uIEF+zc
ZJrYSMJTAZ7Tdt4+q702ioGFU7wrmNe3FwDgRkiegKvdAn/18ZJTB5bQhoPVafGQGA7DeQWDW+fG
k4/Sm4EvpLxfbhMbDg3E61f6yI10rYdkfIKdYgdbEQMMsIm4IwZ+g9PYGxMw/y0w/PHo8epjGJke
g9Ls4OJEs0Sn9SeWkzKVodcePzJzqi+EUmP4VftQP1WHTXmuxOY5iuimi17lnJFr5CAJRs8vmz3w
QpMjrA+X8H9X4lPXdzWHwk/0eyBgFwgKcGLyC1ZkvvNnZvej6GslrOHBYjXPnEcx/Bh3J4XP8WWe
78ciuJaY1ehlva46XNq5ZtIMBbU78TfyYpHe9hh0zZZaYxyJW8gcHVoejk/AIFUt4KCg4V4aKR0t
gv523TBDp20+3EWtb9Q0wmcKikRRx18G5vqe025DDjF6qdnDXMx7FkUAcsQirYhLR5jrTL5pe373
T+0jAxemRNEpBkcKogM5+edAZ8n6fUgO9e7HdqFGIagA9dFgiNH5Bszn/BgYW0DZkLLgPJnMGm1a
LgCr6UL4qg0VYGtpoW0z/19OdJ1b8+pBSOCDDVcnvAMtD8O3S2b4DoQ5e+MLmDrODIb7YnxGQ6SD
Tw5E9b44xqWsmCQwyF1TcaXDcPvx5nxczmWCu77zR3Iyo7G6eOA4HEeWVrGgfDi9DxDauszIjmbV
pXKpw+tANzHRLj1khm3gjwtyJOrU2yO9cEHp6z7lSDAufKzBZJE7UxLG+wnACbfZBwVc0gaQ1xNY
AImTDUWLVIXN2xaETq9DWwuXgJfdKILSh625l9iKM4xT0ULohZX08UOtmWpOy7xfQl/sC6yP652Q
TcKLyxyHrNzaTyGSU3KWlHbpBm5Nn0KuXGDOHsXE5n0vmz5y+cMkhPEFVfgfyGtA9sqhnZrwA/m9
DRl3CD5WxicX3HdZ0An0yEc0lbpGWKNtKgWhoNmZzgihPzzdAPHB8m2v3iqO/OCbyr5+qoRLYDbp
sZkoeAivG4Z5kqllqQqDHko+BIsWfkUa4DSjjo91TuBFi4apnC4pojKvJpG8VG2ca/gek46FzwjL
sI8ip83P6Bmjm+myXuD53pea17QaEVCvJyZq13yffzS1YgHWgRy06LJ0GoUqYp48TSjfgOH7fD4y
7Wb7+HnIhc/tu0Ly/TRgErMfPwXTM89V4Y4iFrxXcuKVZHqO+PMzPehslA1oLkhW8YlPZNNkMGhB
V6WpHzZnpLCf3iliUybOqgz9uw7JgHBUMJmETOQ34Z3x9PEGKy9I7DcC6la19M30tjsPBvAFtcPe
AoetGe5CqouQRH7Cifk6Dkd3NfmhXuf2+KElY10BxZoHK5zuEJF24N3laqYGCNZaYxEGoTM/eWMj
7atcf1kCvgYuLdxGGiMPy2VZ5wqH0mJ2C/s6lrc3zfZHk0FV333TO6yj4AaLmxBv4+8of91JeX/S
AMSfdc97AN+U33w/jh0NAuggmMUyQh+NHdSuLDwH+1XwDMrOs90g6k2Rsr4pGrFxyDA/bg/OlmE/
omMd7Boe1ygIXR5SqynMu2e0lDs6L/yynczyvqRS+nhxLAPUfvYXijOahqsQUeh/zw3nY8Mk7OI1
UDNPtRRGRq2OrytlNE9ZuOUDlLaDjCBB39WraK7xeAxmyd+dVT9ig400IzAB/LFZ9CIAI5n403xl
yFqJkjmymI+edHpBEdKa9fRsd0aFHS0A8HreMMol/Bjam+U7FPkoMPO4pTq63UbEMmTdu+IZYZBP
TpS+irKTnjik8jBJ6ki09k1pdDID3XlJyxJNfi+WhmAD7TzD2xV0j44QcJ3mcijd/ZK2dmZ+H6kq
zGMpsPznZHjIa7oV0vgyYPchxtd5WC8ANfc/+xavrTqPC16zxarkJGlOcfwzEjxDkUl3dcTEETCb
QAEHFECEDLZxRcs/WvLtCFapQZ0A+Tp83xjoR1+SveJsHYl0jPNBnm6JYY2Z0fzj713zJjP0MqmF
h4L7fK9dSeIC+3a7K0haE7y7uvlxV3GFT/Tj2QEZWfZx9YSlojjRNCXIQl5yoP5c5P6XRM2fOf0u
me2Mu+0Mq+5a+4IKCBtSd4dHUggfpb4LhhFRUjXsDnz99BxLEYIAXWHeDMYUepaIjRswWM6BE8Dk
SleV7TV88w1+kyZKJidrDdosgc8eReUPS2DnAwAe62jcmneoNDyQCQ24gosW+1XoF+wqMaM9/pIs
NcwQxCeAnQjuIlnGS8N2BXBPrPGetOxb3oyY71z6rcvEollCbM1UBsw/wIAHH0z4mnIhQE6+06do
AyrTpWUms/I377PFUMFjgeeSz6N0+40rbsIJ7q2I9id3CLDhNv8Ha4B7fGSdAKP2FOTvm2jt22GL
QDjcYLZc3L80kHFT8pINVv2PDEiKRuTnrDPLwVJm/JOI4/2gJ3YM475S9OG4R+gTVjJnEawJNX2U
CNXs672bKRMDemEH+ESfha5Qe1vMZj84WUjRRd/C/0hUv54G+qtThtXjC9zzzMEx1dRVXgA/dmSg
c1pAAEauspXcDavAUTR+IWYM2cA+5uttJzCDMqsxY0qQNfG3s8xeYR4twL5vPT3wUtDxnkTrqqCw
iMcGhPnae+PKzt/IwaSb5wfScEm4OwbWI9xIPPSiEHB/n7N5z4KYrVBbPiSL6fCc07oeeTzAhNaP
e4HtTYKq5+4+BCPB75qIO1szi0cpjazteF9X02dtXJSg+ZeykqRvEQQjlCbqtsMcAyWIrN4XnUQz
wPt0hinSFfzE8rxlsDEHTx1T6g4QhgmM38lWmTRMK/nwZgNXn98F4wNhiY+93I237OHMd7xH9wb6
Q4VhG2E9JDmybJYQvmv452QQelP+DvHTlSQIyzN9BgbhQEnuDFtQtAG+Dwyu1L+ExTqAXJ57dStb
sZuNR8HSPiqdC9vyDnI+8QWrOZWcQ303tjWIqpA2lLIgpnQD5xuWTuXBYII+v0xrCLHzE/jjs32Q
VKKw3z41ifzMZBrjpVpnp8NfU/OM88OAfM6AmmHVlmroQoXEI+/WS7cveZA/k0U36rQEzf0IJuy8
3IUihAKC34DFy0g8Yl5q6cyndrdhN/Oc01c3n5Kjm97/njOL48GozygEaI3squkdqGiKS71at/oB
/jboXk+XvRSIefufKbB1fhtdJCztz1kPC7ISmhnNXuy9pYR4xYmSnIkvzf30AgU5NnqY9NR+LQgr
bU8axtdFHiueO3gGAP7GtqDBVTlSpDnucKWQ83HEeqPpx9fx40/po+sFEcUiIgP4f89bSb+xpf21
uxkq90VdqUGIZiSacE0XjLW486D0OARsuwSHQgjWMVMsAM8CdBpUxxKdaDYxpQ0vznK3EJakkrFR
hpH0T+yF6AX7WwMe22/USG9EourqCd+q7/hMMR91+X8wjY8SPlKbV1nhRkrjmKks5fXFAqlRWP3s
ZYwk1O3WgXcI1J/sCrX1Pf7euQffW3nuUpK0z0lo79tRUPfNSmafX+fN/g/sNjNE6Uc4bmUNlSvj
YiJ11AIBAUzZfaN8FxQ/uBS0TXs6NowmVdvNOLby5DOZuWPj8KcyZVaoh7/ZUjTfNc/M9kren2Gj
mvQ7cyYR5/jD3hD6sD3HVLrchd9cse0MwT81fiZykmvHp40P5K8WHUQGAMJTIjG1GzMg5GSE/fQW
uhIAB7jOpXRKXcDqU8sfD6fSILZtoG8IueTkWf02F172Gxb5xLiTYRxwlxqJMSQ5gpAsmolcssNK
3K/iaA/ym7xGrGrLE4WxEiAeyCHRdYDo+qkQneO3lrq8LOIjWqA3UzgflvM6vPMJp0arRn3qGz1o
L5Qbm7S5prec8WC+ueDDm1sVIOfPnPtM2Hp1llXZEkNnJSoDuWOxCTqz4MYIR+hNVoThRBEDRqOs
HAXu0Xd17yzLUEID4/8WhWAkfm5vMbgCmkACvmOmZTIxwlUqdmal0AMohT+NALQDRK9rGm79yEym
xfGh8UFi3D1GiKeGW3w7rVQ1ZWxpcYlDBekAqGoeh1WqoMktS3he/tCx8GoDEW3D9rjAbGaEaqls
zazO7IOIrGKLjkwAndhcRYJ6N9kU/U7gM4PmsXlh4ACcqf+zhTUX8PiJEu4hpTRpcuqXsB7QO2A6
kOTFxzdmOVarR/2QfqHIviMNKarNuDZBZa6VAPN1NYLHm/+Qbd5tbYubiZT7+FGRR92+gbiHMLQC
k3jEJ5/DLvPcvYwQxD/PZ4t40dGrxe6cCVkS1h27z41Rq4H6JEg/PqKrxUUSLAvx8DTIzP7jgT5L
EHT8jb8ETR+wVolQqqZ/mupKGVRTw3hwwX7qS/Ygr1og4o5JeHd93ndtKuFsXKxijPV8cKL59qPZ
p/r3fcr5WpTltTIhe/lSHSDp260K71UAlis3ggLA5oe/djcOz6pz1HdddY6rd9MIRLQaqHOcAHf4
JY+wmdQPuDq2BVvtPoR2sefvoli87UfHkyLiijcqUniYFFP+VwGrlVa59+4p/ui22VRA+6MV5qGd
u1/Nz9glwNU96g4U0d2ncZ+wPZZ4CjiHpOwAl/ndPaQXMdb7brw9mJy1t4hefN4DwneiqlLuyQH/
qAIqqSppa5B0AqYS8SfSLomgmDCB4gLcInlSp4ZiJ9A7mZmDCAjhqkYkJ/FNOCcqW2mmNto/wWkW
gl9gc/j2W2hr4EWKIvy4TgcipILhP+CHdg6CWhKVREQs/W6CO65k98s6SQ1d9hGlHh1GzkUccoTL
KxTUaQLcFVW90jnoqIWAGOJN9CZCFqCo5vx90LM8PjsSV368iVsiiMNPCXaZ3/5R+gUrBy9rL/Px
2+10iPkA0mTlj//SM575x5eNjjW36yDpu23pXw8Bd61p4Xt/ulEtoH3QoMqcc08VDXkjw++XPVBV
+FkuZyenLH4hPW30n+cTLzRpjpwTL5enhU4QmgC8G0LDWniRsAimIh9wZ8qoRd38QY3E7eMAKbkT
AySJ8ZgtJFLhaug9wgZlZ2xSEkKJz76cX8VMvPyfbvkBzrlNnW3eb1JdCqjr/sJbYxpUiZgoWTGK
AyCaTz8bzcpkC9BpzMb6eZMG+3DGE9qCsUWkhMDmVE7273tNZoiU6LopyQPP7elaY04mL5txFymb
pQUeo5sn5wQlOHSOqxFUCdBaGVb4kvpsZOa1pNRQar0Key6U/UYi9KgepgVUBeqnDHKgRuygT9pQ
mCOJQ7otTS3JwqfOivFUmI9gxqjqEJ4ZslfSZtVyKMWM4wPVAYClZ9MiCi3HIVA31Y8Ct1MEv1XB
w1k2eRn95FRZm4puFnv4Hx82bxc9rmnAlRi80EdN3aJikHX8EL60+nTYc4xV9eOuxo19AdeG+Gz8
M8ThTl8z/hf/3kd/UQIOjWniIw+vq1+t2zQs6xZRCRLwOWyiAlyh8/pkUxCcsIBncTI0lanCqQ5O
qJix+3oJg4Nygl+iU8YdQKE8HBb0H+/oIU4e28NJ24N4zPLfZjFPKBxEorWgaOgLiNXno6vSYt25
yYaBu5bDUl7OihZJsyr+WAjyjAF3MgTPx4ZK8XxkUzeHIhZuMJe7yYPaRCMkfcTfxVilvlDCRDAX
k9HN9CV5byk4vPptKZ83XnzkS2GTEFks8pixpG3nIH31C1v694DqblYaPITI77FktmSxCcz96vV7
SV2Du8mirR5qZc2olYjf7Xfa///+++78roMbZXtAwXmrmzRi0Akh49p57yovccFpCoO+xl8WxLzL
S+7uOQXsXBQDTlqlMvlkz4QWIUykIfJVuw0nG3S1U26rgSxonL/NdrssxVhEk0cAjNbkUqaBywSP
P+YvU/+z/AVJCjqhkA40FJ4K1x8A18/87Dsf+DAZiwYAp6dCPbi5TCD3J2ImD1wSPPcrVlHeLVvx
Ss2ZYu59rJ6r8k1FMTV484Mit1+6N7HsXbAboeNIOFTTVtHrSu9QTs6qgxTD3RIymHi+Ghzjjz1U
zZ2UoPnmh/XvsZ5r+ZFPnpSLtM/aW0aGoSRdNaBPAcQMP/SUNYqbr4ITNoXSfjn6QegielK2RDxD
VNc/OZ6Vg5lZQkzVi7Zg9q/QiVr2YinNYixlX3KYSlAxz648TXdgVLsfKPP05s0OntUAiOlm5fdr
GdH4K61rpuzM8uqRcEXbQ6GjWMfKr+UL3gH8TkZT2isETjnHrHZkf1Qv5++nFEZHWWGeb2PV2pOE
eMoypWGNP0tC5M463aXTgf/wiH3oqOV54Jpj6gcjm4XTN2TY6Rll2lLhLo6q+4j25nLrVmSWNOK8
lOfHBEq7un3uIg+l1Gl9LlrK41MjGNvnT8+5yX24dlJzh1i1ZVJrk/v2s7sEYt8m4DKexwb1pCgL
xmaLcC578DAHd5zkLZlTDzjT9nnnwv6n47fDhw4Jfbql01Oxm2LM1ZUyJ65O4deA8lirCJ6rDLVk
GSkIAALwzY9mJYSH4oagldq2SymfmLr85GME2XHsNM8afTz6KbBIYchlNaqzC7y6H17vwnKawnAC
SUzh6ztI7c838kn2tMdiPfP20in2zrLTrp/LpxXRPQO/UOvoDAFpZnfml8aszSDy7GRQg8pijukL
pnxPmq00aPnujJkJZSvcZCFMadgLkwFgkEQEERWfY5wMOwc+De/bp/C1EEOUpsf3xpTjjMe/YE8D
1J+O2LpGbCY6LC8Y2oq6dl2kJjMxgpuc9EKhzyoZSfh7xgKQst8KF/fsuV/642/QBFIinsCUcOsn
Sj2kAR16jNzs5rh3xh+/vEM3BW3NIvw1M4H1z6p1V/+bkikIviC0ZBVKcLwJ3O9lEpMaqDU/qIcj
0+6x1rAidGsWZPLQF62u702hWXGbNlF9Cv87Glct1cu5yf5KgAqHFB9vC/gigjk0eYRpSCvvKCKF
41uqsyjINi+mgpdaS13FiY324K8JfleOxpZfpmzYNZNWPkcZkD8MfBJBE0V2qdveAE80CThZCvF9
iQ1sfaE7OvCLoylf1RcQILEWs9d7ny2ioE9PPcC+lGYli0Kr5EBc6djXEu11y1DjMd1uKyKLp3lv
V0U+Lr4wi76bTlqyaxnA5GE31vyX6+9RXV2/iZsP8ZMGNXfDGlr3kxzmZypQJvPaQgerrpAEpvd/
WzsRweZbyLc/+iQLxr11IaIls09RCnKI/x7opmSz1vUC7di7p7svHwEERrIATvsEZYGArS8Y5O8h
bTo9B7bmVT1fg538O2jOwsJ6EzFbjO8xdK3dR1ksS9p0ApksWzns3Q8XLIDoCmjK+i2r+afg8O5b
ZkDPi7cEjRp4h6WNxyk3P4ua48ZWL8vtuPJ5Qumsyf0FLh4GwwPWmNOJnPUstyEvmAhbxT61wC25
gKYqF0ZcgjEN/6hVKGu++tRPvRcH7g8YTpu5P5++qiRpq3+Otf/c4x7P9Qv97Y1UgNMKnpwxFk2T
xUFC0BD9d8sVN5TZf1lQgXkQ/FP8wUx1yYDWhyHWvrl9QnkgsGzXPzXDm64jW8d3LdTmEOJyyN4K
rImLTTx0ZM6CltGpwwEi5JYutZKQZD0ZESjjnIfs+4Qx41J82Nn8i/3A0GDUjFHcBKaUKzXUmwuN
iciB/72DEgF96y0ymsM1Nq8Miwoi020hNngqkffwPFIrpjiTcJpaEcuoGuQWpWdRB2HfxKmvUJPj
9H3bhJ968rfHbpm9YxRIUKndTUCR6DQUjIyLkqpPv1P2dTEIJeHU41u52C0KxvtGCUKBOzFkEHQn
pSjsxzIC5r61Ize21MzTmPUvZloIrO9BBwgtJEoIAtsAWy1AWO+IrLM5V5N5NBYwZ6ky/k7LZHc1
Y5sceAxf6tem+uFrHLzYZfF951LqeVutlE8zXqUNi2VbHgodxTNy+lsq0AZdrejhau/hhKR9rUyy
yDRUUnd7K230KhOwhuQKoDkuIO0Bniae0NJdfPyYtl4JiFd4kHCfVn3qM/r3ArqhLTcmUpVnbkRN
7Jl1QY0wQtECcXIeYjZ4v3/6nhED0X9HAuqXwR0n81IcXbDU5XX7vbOsRt135hga2o10Y7Rf8iP4
dm9GfJ6TWpf8StWgcY84XugQdc7Umla77y2yOOSdLPyjkI/b7syy/8sNxauBpWa3UDnhJ/wzmVHW
ppynO65YTK90yv+pVnkx4UZWmvxHal8w2n2XW2J0GPYAGcf86HjJcnCerHO8tM3Rz8QNo9dk2j0i
/XYIl01bOv8uBchxm9dv5P4TGDuYHJJwHroMzzuFLfFPQmumrmuZOcX5xa8VBV/9d6mh4TMRzSx5
hS1t7qpsWWoiaItRwHtnKvxTGRYu4HxzZNb6sB5wSVatZAAlp7nJVQ6OGPFdJ1RqUWT4+fq/Kq78
ZhbsragiPaBn9ifpuac7hIgKeb5KWqyDbNJ1ppXLvqgqWjmDM4ufdrYR0bTuhjDASabvbMlXArza
3XMp3t/Db9OE/FlBp5zt4hNsVy0VNs3yfgK0UVCwdnR72YVDQ5H0JovV6IEW2k3DVZxAbSHeoz8u
Pf7K4y7dwU//U+JihkPpe7Z/m2ot6uDzaXluFIOKa0Zp2c3ROEVU4A9Zvm97i5d0h49AVQc0nLB2
3i+sjldD7JbeBhIIoqXJNiLgT1XE0/a70NxwsJN2zNSDLaFstSZEAKmPr5SMwxbtpXRNRgJra6Lp
MH/7oCuzKq1ieJjjN5nwGCbPWUpuhZVgl9OO53rS34MXLvabLMF2OO7zkaoORTUZdOkVlrCqG7to
rJR6h6PQKMBIsrpPMiepGbYksirMcE8/xIBWObFT5kFx9TGn0OUO5UiN7MZ93QKk87i3nUsb5PMF
LlGIx4NUEqsQoPqn79JXv70+YNMDkuDR+Tf5/qY4CzXjn59h0GBzaY3qMcHEAbZGKy1dyeo1dxRl
mhYS7O8Z6Bvu6jFF45vvPDsyZrB7Vhk3tNZ1Qi5eZdWn82HmJQ2OKJ5V5k1ymFPg23WiqpNspE+z
U12ZzbTugnWQdW0q35BFclt4N4G0bqO/bX0395CoZ+e7w3p34Bk7KbWtiBaFN+RV2WinO8Yl6yxO
dMh6ajgvFioW2auDENeHz1TBoqEZLVsA6XL9d7rbt0d7JlY8paiJhrbxUvCltJne6ceDbWjag4d4
Df2KhMu7KoZqGcqoK8Qx173b8mj8/qrq+qApyh4+RqeC7rYFwMZgzCt/dvfhp+cVUtX0yJeUKUJy
0bx3beHVxgTVXAW9ui4ui5bbKsfOk0w9p/64ovFtUIjKG1L2SKU1LcbU/YQ/Fizxl/Hl0aUJgT3q
liqBnlcnorAoonL4d4I4kjDBExS5UwDdW0rfaQ3pzi5h8WPccb7AIctJ2d33wgP/0VtRXMTf1ksi
gPOzq31wzT6MZbuGqCKAkcoix4x1XAAphFEszN6oivbIYcPxX72a/nSR56SAMvUzHnt+Jb+eajPQ
VgZCcSEAaQLEWzdJxrEjrvjl6HZHKelPS/6i1GRgWFyCqPCUvNnSCXoHAYpapQFXAX5Qrqku5I7p
GNWbdMHIJy6Y7RZ1mAeIyW/eLgBm5fjDhlxkiI6/m6FdIx/gqgWlBu/ktjiq94wccIpoHa+9lt8U
VRgWm7rO/tipeCqOUyYaZ35bd9zp+/toIpstJPiHaXCkGkTO+uk9ROO2wDB55XNSTCNpYd8iYmiZ
repnFKxwC5jNmYODfwEg+3qTqw+MEVYeo+qpV183moG7rR6nPU8iuBpQEGtuX8462BttQaa4jwz9
wzp5PWVZTIG+SQjmdtASr3MI7nJ1hB2Y0FRSDXXdKgd2QBT7XLWYFxO+DM9nmwQXA5tl1wByi0RM
Be7Ur1GGFXTijRW0WYw4S9lUpeLYoRj2KZ82GDSTxbmV62DTzWihOxYP3OwGjP2H1dB2k5TSa4wg
28sV5dcN+DOk/KZP+h7AKRMCEW2g6P0JsjJEIMLpctcNR5KUqF8oLtd4c6JonQR57Tyvvj3s4R5x
AvTwb4AjlbpiR92tTKkBCEKnivz4qgo7W8uFbCEKCPPinVHMdzBN29SjIaAo1w240KRu9hGhuDb9
qbkTs6wKXgGC08yNoU6yi0Iv7E6TAy/aP1VZCYedzB4OWuanNb5LXFKwHDwaOn8QJDqWRiZGBrjB
aqe92wm0MNwEMAfOLwzxwyj2W0nm+wKlYD0tfxOp6TeQ8qt2M8yBy1Bo+fH2yYxJW++vSnSZVIhM
KvUVkEhb+RaQPt6+sUfDo2tkhwGq3cv5nSceIuB0R3Y6C3P9Ca93Sr/RE1bXDRiyFdAHhEKFGJ2y
YuEZxjEwgq1PnUE95d0OkEnLbex91dLd2P1rBSiGF7WKwcEBl4DUUblnaDPnXerlYZX45zYznn/R
rjH8VMVc+ydDVQ27el7VsGKFTJyHi/1v+ZG5i1f9uEiEpuhX8kM00gjtQ4Lue3KzjhyOuw1ujOPx
t4T6kwhUFZIkNyHGis4phJqMY0rYIOOHgUZjdPwJgSp2XcumbEJerRP6weADlyNVs3MTwHvtOV24
UzTkGrYIz6H1/aao8/wH2LqFc+mW5yoJUww9OCVT41s0oU68+qTluycJlK2KIpQB9Hh/LTWzqLZs
oeWkXeFQBBqmTCCtoEL1GhxFUYJp5ugZo/fBcJjX0fl0cKllagNlHo3RFFualO2w0AGj1ltsK3Vg
TAhmptb7SlODRY3tbnf5UnxxshmoHm0QvlSNWCRxflUd0sBVexcLDJXeydALXhJLkixShD3TE0Mx
kkQX9IFKv90+S4aPTgRVWsPw1W5ZJJK/A/atIQdTvUL32lFqHc3iGOj5ATbdteT8kDqKShHraZqI
PlEqbpPECbR4RMYyY0mifhL078iEcmalTSWfg0JcEHLURc5AGMnQW8HYC4plT+we4XLm3PVudff4
j3l9AOjHa0AWZSYZ9I2XMlZhln5487J0r/jiuB1gjaFk59wxRfNsaC03drb7Ss8vtCQbHyZ9nSF7
DOUm0OrhJFC76GtMBkjUNagaq8TiGvTyxsPkxtV53ScI03mU1DqeBJdAvnttGuONjyS7F/qkW0Ty
6WxTCHYLvqKyRwEq9MPBN46KO6dZV7CKtJHcdDXNnyKUd9Bt2N0CKKhSuF4yyAr7Vj8/AzqCKKmI
ydpcmBQFBUV3LQ/G2JmFyqyeUs7wumCPg/W7px/RcnZM0JYpdDBfRaGuIeBxBcdw/gL1WHzL/PJ/
nfXo3qRFV7XGPFitO1soVk9r9nQcq8uapscGW/3MKkNX/40ejK1u5qlTXOMvemTiJyWhkU8ceQ/n
ZViu1e1uQALxd+RS0LXznEDohIu0sNwecZvrmgk9iI/Z3t+H4djsPjb2CzUmHBhzu0QCPtFnmABN
n0O8MS9zARd++vexyExVx3o9FY9dyLNQ9l+LTJ72rk1UY3BLoxFAFWl1k0QdQ5qooFkY4I6+cNJO
T9NX8XunZGOH431+Wt0qU8nMOcg9QbKSRNvA4F/4bVfxvuusXiMI+1lwjLEoahXoxPkCBvOe5UoZ
JVI52lEPzX2nkf0dyDoUQUNUqR3digOBQcl9ndEf5i4nt90SsifSJpZfVRaiD5OVgJjcckxSSruW
d6cBWqomUEaEYZS3jxA7sC4ttZySnlDzpE8b1Wo8L9TXeGt9wDBu+C0KMd+zRMfg+P9G/FPn8ghM
j3IZ7kp9+awTzZ+Q3HBlHujklNL7K8o8ZmaT1I17ixqrTo3RbL6h67qjiOh0XOTW4nMobyOCSA+j
VO/VueUz1PbZcKZagWfDfknZCJ36wya2gHf4iuqiNydMLS/bnD78N7byojLfP4c++nl+M9kOJaW/
ADuF8e8bmm9ceszwsJNhd2GkXVOubPmIKEa7FxhuJTMqHkwjdUWLXdvwNGy/qHJQDq7qKz2EYVqz
XMN4CCgsaE5FbK5m4FsLL7L4soX9G/sIyBuLG6Fue4VuDs+mJ5h7W+sM9EcTD+8bcVHP5Vp6nKf/
Dp3LDizxw1D2Y1KMZXkzVdBK+psJyP+ipG1zP5bzcpDdYDgHHHV149LiSeGCMz5CJAdV5qOaNmeg
pKK8HpHmChv5Dy/KXCd/FUVG2yoqH8MbGQGBtOa5uPU6TDMOleV83YeKvj5LFx80xDf0HNgq58rF
1ANEXos+s/q+Afwww3v1M7IMeKAEyLvh1fCWoe7WFtXqwAYNl3+BriRO8ARAhSHX5ZuIFaAdfJUz
Ox1/hCYiPy1pbbE7fFQtVX4Nx5/f8wieQyTNH8z+qvTfkJUjv4vMmq9jgUucC/xXmHhx7sRUsExs
acOiKEirbhuQPwE/XjjkSN0z+bpPRIbw8xgEuq9C1NO5oVYxnC7ZrXI2ywy/1W6NH8CM7Ud40ebs
kkPS+kwEt3Vyr+nGM6nHLu6XUKPMwpyLMKELRsvmktt+xcVYMhYGDlQwG4MJxPhEXPmZQgub72LJ
oWivBMPBc9KT9+Ay9s+OGZuKg8zFEukCXNnaYIBYnu3jtNsD5TKBW6Mmi3XS33ofvVMC8k246I6T
CwOCXj+oSzl9ZNVGjZaeq3UQkrkp1ThrIVEUPxB2WPwnVUSK0rcxn08qIhchqcSyNxvoIswp+t3J
pPBGtIYQGSorcx3gUmIVFpF6GO21sfZzz8btVJqK2bsdWj89znOGXMp0nxQNMmU72rwilS0SRgSh
i//aMsmEb4vK7etnBP5mjm6Ui3SgXx0H6OHzbM7FwIAru0Iks/yqTDSYgl1ewvSa/l8IjCnOliBK
Svm0tiMlAY+3W6j3ODH7vMIGjkzJV7xk8uUd01FRF5096u5TqeUE900cNseFCWHX1mf1K18ZQcCx
1lyGZc4Rnf1NpiZsdfH8P6e0nYep/bErCKj2y4Azc7+77v3GNERkDuv2or3p0FWYAlEpAEvaP9om
ttkn4kqrsSxvaQ5Qc9FKxRZDaloRnZWQJY4vpw52XTCYlEU7+CHfwWDGMDvVgTbuMnAwcWhQEurz
xe4I3zOJ2PG69eYBlFHupOChGLDZBoKbWCvgSSxSGFZO3E44Cafc5c5/AIwNZAf36EslepKi3UzL
HRGwufWuR4QfyUiWBzN7APLZDl/GEZbTBMDImxzZr/iNx19PrLxN0ZQvkmJOhRX+wFN7j/8Rvs1Q
KeIDi6srVdvesH5HYpoQ4rWgrD+asJjPM7uMw1oSAa7+vMGHmjjP/dWEQCJAc6yet0SNEF982wu+
HA+44OX1dMdtOOOr1fBiSSyBbz9iklbtgzC1L0FBet8xXOd3ZKKJIqSbXMZOgNTfgGF8grV1ffPa
eSc9wgCvPVm9/CPOOLGDoES+6T2e5ggNpskHoy4dP1z2zMs5LxV1Ddn6uO8QP2+bf6t/ziTn62it
5FpGDN3WxfECEh55P7xur5PPK5JMz4WFfWge5WBHP66Ro8zck4u0YL/rdYum7P+Tgf9G2FkjoTtQ
2NYEcEjwXF21lPcVuz/hbNqKToB3sMlKm9nw2v9imPOqJgTrwqj/AfGy7f+dRmlMoOgWUzIOM9I9
jZgiNmZgPGs4C+di6J67DKKu8NQnSM2NQXrHLgf5Mz8TBnv52GyZPTl3iEZ+CDW7MaHKX4sR1MXx
vy4Fi4QKCoZq7Beh+TlkcVQ1Lbsfc/NzoAf58XSYGxVIPmCy4JYO+kCu3JcnQEFZBuCiUIgiOhHQ
e0wdwH9giPZMsR+jsqIAYmPdG5+uPMH73rTcW5MY1sGYNAWnBdzdA2kmzTUT2cPWK+9D3UrHNQA0
Gt/y59jfB5PQt6kCd5jvftHbbVcKsPvVkID34C6bHzlgYE63NlqeGSEM1sklSeFIjtyWoKnmgpEG
5eEuw0c8/t9wQTF7KWKIcedHgoWNtAHiKfe8BZT/c+GkhNlwH0FncZkAcqOyPQa2AYdbCN8e4KKa
kswbYK6q5UxAuaxe2ytgSkyW3kKa2CNIthqbWI4eTrPwfWKQMeNyoRNHcjG62FcDV/QRDOZ14pKv
U413Y6/BUj3FITh8qgyolQcNBPmNLsl93UUh6Rr+WrxWlzE+XmxwhgghiL/EzLmuO61wWFPJSjdU
ldJwxuWqnrXD5BgJdZxrVrULjk3Lo/g31EoTeYshv9wGCkoq4picKknlo4mi2/ZOr6QAWrWqCxpI
AKMsnoUX/80+Gsg36Z5cIUcXdHxfHOqFe80Sl+JBs5XsF/WIx/OQpfiNnaemxkjfcVIqJIsu7js+
oYOQAtk3O8iEt7QuA314wGizuUoLKaNAVrj/dfYRGs7UbUiMXtG1JkbBrBMzzXB3qOeaiCa9SBih
LZ/BGEAicfczxJS4xy79csi7DgRbDyeNehxwIMWLLwVdv+SzM5WgQna9IJomEyCEgifDsOA421z7
jGtofBSGRem/nkWd5wmPRVYEkmvCmOMYcrYseZJEVgSqK/qDxQOEMKr9B4JgiruS5aYFyuChpvtq
tvKL76R8Jw+YLC4Pfl8jGc/ijPZeM25r6Dyzt2o8zTd2g7wksqAYfqWyDJbgR5D8E8hXQmUElJFV
zF0XIXUDDzBv5ERaEW3sLtZPmaydyK4aDC50kBy78R+K4D7Q6OQt4mRJp0r/UwdRqD0PQCfPCaIe
B5DR90uAp4/OAGdwbxE7dcgM0rVAnR/LZw7IvJYL4Q0gwLxhVnjVo289gbAC5fpeR+bOft0IZHA9
3EwcHYypT4uJm1SZnSlyi0llOdRzcxrkGQQeOBQZp4bCbFSVKkOrRu2DNbjX/n+9+gijxsrSPsYW
QYYwZ2GQhVfBSGlfg6nSwNrZp1/+BgefUMvrXnaigXwX1AJa8FpHlP5lg71BhKGiQbmG2cpAJn2a
2Hm/0Neu1dMeO02mPt/29DWlj/IQo7BBbRDnLyUYgxufnBvzJRw/cMnmXtDXZ1PODUICIyj6XJtH
zslijURAJ2rZDG1AY3tXfWRigVTHHIo9hBbc0K4S3/BiK1R7lEeQKVVTd9+LBwfpH+DHdqPU5SjE
Av2iDit3jbLIBvGfawYsaLej6EcoQgOgaBfm2MPDfRX7QM9dwc+FyVGHIWzWAvNhNu4QRGBgwEDy
IQheTB631JMVruPROGxDzcOFGYMYJUvMPAEnQp2sPj66GLAzfsyh54AMZzPZcG/5I9uSAsZqtmYE
nISDPy27MfkA04zax1nIIIURtBohoFDZQvvhF6psIiSCdK4tMtpkIF/ulwldW1MW2JAZouXs0CIF
mE/1y7V3WsfrKP1mSVeZ7L/NIV4VSoroN0wCekfB9sTnMs9mten97kJL6UchCDl7M+0oM153yZI7
uv4C3bMidnPeTktMHDnqPrHQwjZkOMNqcCd4SXFca5qeBN2mTX4F6zwydxXwm3DwTXtM40eEa5xm
Hu7GdViAGSP4UUVyUJ1WORc44WlSR8cayuR5xzmsFa/D8U94uBuPit9hRaljHA+WRAGS+YWtRGYw
iMZ/B6fQ/t2JktxpXVqOHLHUonjc+vqy1rzuAeubhHUjw5SD0QeVrMm/lJXDvaBbJNL4R3TFqOVo
yagRyBMZg2SgglotjosA8QBiSbXDUvx6i63H2Mrc318N19Mw3c7Rlajf9umy5D1C+//bdwAOBIIM
FuKZNuB4B6TJfBWMn5fsBwXLrhFY8yblxIMYEaXcEpC5rwyXKDH/V9w0orRGD/q4ZRo66DznI9fg
XhQiIqmbPgL21+mUtE43dvlkcsGyUZUXrGX8PqIwO9ejYP/VddXLnGOWAh3JCeLP+nzhXIhizhGY
FllxYuDCop7tnhsxCGc/vmnvi3w5xs+wgAXcuNwDgKTe/eC6TjsuClqyzD5q1BLSJqEN+uiLeLl5
LxOElNdTfqzjG+c/lb3Qk4kkZtdH/9DYnm9dU+jxRuzxZpm5WrqtAymEAoiyjyF/if0/hKSeIzbP
gWJdZIQL3Opz2mhp4ksR0zpPBoQ59N42bGyz7k+f+4ImDP2fHkFrZ3cPnjoVwftTmDJoKY2KF9cy
4SKQwcsFBZvJFhIGu7VNsAZfQfXXCRHfELNNL2A0wco2z8pD/nmPeUGum4kMhH7/DUcEiQ/TQNeH
/kT1AtTivF5ALl7pZp3d+VFDpSt6WqJkWJ0kQeBMdv+5oqkppz2jyU2H/OVuHDUtkL5alGbj05Aa
/5Nv+iam+U1jga4Eh+HMVoAj58h+8apcuD34OdZT21MWcy9vY3fJbsGTyqA+EbdnhYM2OsoA2IHw
yLUlfHYghbAJdTsK+K22Jdjh8lqW/Z/UytnXun1T6IP2Tl7Yx6vhxCPY4bJoccf+uj1EUkrr2ePl
zqJrIqUR7JvEEGP2DbIa5D9unLHoCX9TvOKDOEiuOtWnlhZcTnw4nE1TiP687JXYvgwi43NHfBDF
gnqdnk4FOMep6KA8AbhQReEFyi0b7hSpwJpoDkM6NWg7yG5NcB7tkaCrQpwU2dBsF+HNsa4Jb+B3
qBNksoL3Lt7SodGrEIy1eM6eYu8/LDRVOy8zx92HfNo9Lpk4Woam6CFah1st5xAprPBDgPblE+ks
VTvB1EMS8Rc+EVfRyT+m2ePiGgmA12UjameuZRwr55xfB8g5KG6hsZrwUfRMlVuuKjG+3hcFADtI
DJPqhTFXeT+lG1a0//d9zwizH4C8RfVbHDnxwC3vbIPGmzMozcnTOgcFeRP9HTfc1Hep34+reLDK
SNvrRz/RJ9SgSyLVQro9QXHpS4XT2oJRn6lheCAeeBz0t74qlTrLHt3I/gsTL0Ng/XuiRKNb7wAm
PULuFWLH77knCnNhgyOLUs/U6GKxV6ykmSprwnOJ3p54SC3qyThz6RsCQJpPdz10/Pi0nXIOlhM2
D+etYIKFdZSnDQ4ZrMNNXvnvUCuacZ97jc9AeiO1RzRxbXZBzfuqGh5b6O0jWSeh1RLYgctZ7WL0
jJAvJHGmCoNnXXJJ2mVvcnz8xsLTzHN1Vd3de3tDbfdZNjlDVUy2pFFD5KtO7F3mBAEm0tqmVoVi
WhbU6nsPPCdQLw0S/HRrGtM6UlaTjhSIWdJzwJzQMX5Q/NNpWs9I+5IZBGc0g9+/o/zr1fVNLmLA
f+l2EtxjBoMKUojo47+9AOblBw7K44ZT9+dcm2N/tkK8JyXS5ctKGNjJvOjew3kGlHBj9vdxzuEs
9gq6e3sMbvKUOif8MbXIt8zjgO33WnbNHvVqNo0+v94mxRh8xfzln0xVbn564NxFpTxcYXwB7DpS
UaNiRjWEh8woeBjS/OQyZjdgya+C7heSC4lNv90ErRjeLgcPm6aGOQKDWKz+k1b/3czidzXt3lRv
ztXQOhH3i/EPLvHPiZyAM8BaFLcHpgFuXfYafgT0ZZBeOAzetI4VkI8m67dpKWENLWIRp9jxwzB/
nNu/PReQOri+y/muY9+6WaEVGpVPAYH0KWPY69pdRzEt+OzIkPK3tUIcDwCs9MKn1EaS1HGSD2S9
llxdrcfsvjjeXmlB7KZ1zk+T1kCruVYbujbGxV+VNz5yLTx5KXMCvtHiQkQ5AZDlczxRzzfhCS2Y
qWJPkqwUFg3HOMpEsUDLxvQc+dKwXJwSPLtTWdaD75+vw5SV9wiKyCeu9W0y4qWeFM5yn3ALinoc
FfBqaiEAgZjDwoyr+E2Tra1QuZNXdbAmAbh35gNRI4TJAebplS8zYbK8wOENt3Xj8cIMBDWFrMYy
y3Nn96bDS9LZcVNuK62OzEazXQ2mZasFdVLt2MthFjA0cRqPN82JNGaD1dYiXpYdOeJWqxobWshc
URNfkcmKCR34yTfiXoXh7OzKVv1S0YQ5YrKPct1ML70gUw5qwwMfigIFzcSBByaZz0exXjLUsQhr
2OKJ+EqiSQEqcdM6ATGET8Lsy7ewTEbTqklDwKtr+KHNeJXAQ2uBDp1rMZn31jCQQXujD4Tn3S8d
x/ihDzDeTywlsubnG3PdSURF/MKrDQ9YnrDZ88H+P/rgJRACaPXrlsFGzgE3OQX00L95+bwMaE8O
zrJm2Vx7WRKiIfRJ/aZTT2kp+5k/V/K0z6RT9zk6xPSx3c72DWMM3QAQGuNDx/xYnS1Phw8IRPRp
hgN+YSYYJ76H/U4jZUnrcjR5LLK/eHScVt/1VWRwhzyraD2+q13R6xebKzfg6nURUUV5jYRuD6Fa
G5c5L9Cw/gmHYxcevMhFftZcwdm6QFhPibAgSCak2mRNGWtXtZvV6LVDQG7MKle+TOEIvHTEG15q
cgzGidiFiWTijT3NErNtjsn7bxFJwsSv/uH3B1Op2jeygFWH1iHSab7dgoaM86US7i0i+cQj3jML
fg/DWqZuUdbgf1idHTm6z6qvO0KoDYt0cjpuk55dsHvZOWprh/SQA4xUKnngxh5sLMsP3opCEp7D
UnBnLnPN66Vwjo5gX0gHtY5g3Wd1BdxaYpOegT8pC0JsZy6BsJie7kALURwGg6wxguxkU/hvxoqz
MtvI0xnbSOKkp9LZWintWp+pr2VGtteMTSV2O9tdZl8c0AaiyndEdw5MkSVw6iYuYVE1ib58jObV
ZZtSXpcKbwYZ5xwNfCxwCqtYIuh1ifOm6AY54EkPOot+ttWtQA47FqB6m3lszxGP1+sKHwyvJtxf
T8A6FFg6gBto1iFf3T8w/SycW9DpGm+2KAiSk76oCR9yrBBU/14vCcVBZsyJOB3v8r4nb2dnuJ0S
RRngToGRMv65gqXJP4vqNVj5fsr0oVaHgxJB0K0lsxj1uI9lRMz6dM3r2sLhAr8PTKz7V27zstd9
Cy7rntZu6CVDK6a9vAO/02WU0R4Wx9GJ9XAbtdHUBXKSbxJtSSDvlyuu2LLzUsa1anIXdkXsXljV
bYx37lUqoUGrssDVtZxzQihQSgcGbhboG1lHVSh9OIAErUfz6vqYSQybLet6nbLQ+m8u/odr7HDQ
3o5dS7WPAYfRm8wMItOgIC5KFYFSRK5uEcoaVbXey3FWqVn0CaxrE4pXbGBmDr5oExuA9cN+tNKy
UgK7FrP7bOgGLSfkFF/y7hHKDuV3CBJv/wPgIfasb6B2bONTbUc9YEOhpe7bv8ZeuJFP3+wSXWFk
nCKaDRpHNHsDA7Ku7yoLGlF8c1A9fIDZykgA5utCeuivT/GlCGDO8XWRjqV/p8AzzZveYdSO9p+N
oIjT/bbdB1lhklBKQm1Cx2xhOwGj1WJzYRlk2HDTZpb8BULKDbPvm7V9vh8Sjmyryn9WYdg+KNsq
aTRN2t229BCbcyItLmeewj81R5igk2Qg7dnN2Q1iiexkmQDU491JECNYeevV0bHDwX2p97rzxexn
cXm/W586krRHqqmDapA+PLQdF2AcWCGj9fNnxtN9uEiAJOmzGaeK9kEX992aBL5ZYadPtosG2+8u
86sSVJ9eVPI18WDFuVRG87cXri+1j7BmlG+B7HxEJ6RNouCsIPAK5kUba1CgAiVAl3R1JO40zaK+
4sBuG97tQ8AFhbOQn4tucobX32ickD3ssBtcaF7rjHRnB/Hdm+8PdycroTauIHEH1z0B4HqzCJSO
clDgWDv939U6NWuFptP9IFEOjpIa0l/r5LdCgF68IxE51mv6xTxV3YRme91lBx+ZlTMHCZzRdnk7
LmonD423Qe8LFbrglPXHoqcOfVGAKevCevBLPC4XeCrnNmWSS6Jz8HHO0E1Hu2qP/ggDV5hIHan0
H0KsR/JTG9MyeB3KFnYnboZItV+UbCUl8hiraPjK5TjMHAKM/6+q6jcNOz5ihSr/o/x8h9SbokMK
F/QCy3boETHRQoTzmuXpWcaa4k1dZBgK4HdTyGRv7xESo003yxTdszeuway9BwRiIY6KhpL+3tKN
b8wubyVfWpaMnFxRDNYkNqYc88n+gd3UqSfl1q9YRVecpKz8B4nhBO1UmbhGEVtiMjKtKSePDH5A
7idvJhv+5Nia/Pwwo0ugQR6mAlOu92q0jmLoLoTzAg9f2UBGxvoi270v68P3wcjbqbIo2QJib0Jl
8cLNV1zsh1VK91nJ8vYNbEaFGufK/hTWYISUTM7nclg/R7Aktr2J2NldNZ3COZbcSvcU/qgxDDDL
iW2NjZuo3pFiqubLkGNTCALW3IrTGdy7BIptQntz14ioHe9Cu4LjiItqrUQSrCgJSoB0WtgJEj3l
y3dDi5B2Iqcsq/rr0YW5n9ooEkMG9aIe2Sl6WgAC1TUdZ0iwCg9PTAJZ+n9htWTkRyQypenP24gy
bim9mK5oPgiSczrxdgulz0NhUFPKxREYo/rzRE6alMBzDJtGco80J4X0+xoJsvd5Vunl+md4DjxE
Vu7C0gSqRUCYk8jMihXQn29/htcBlPqx8I4GE1oE0l4g73GhsdgU07n9KVH1mTS8vYTCApKwKvcn
JpXr6C2emDQuQPEnnDOXEGT8RaKVB0qaGtOneSoWOjcFBY2SSfIua2zC68eIUUemEgh8P682+2O+
Uiv4aBGVrXiPqsLw72cNjhJKWHvmeUZuyVf7c+hH2u4I9LReBz+5wVBf3YunjQxdUApH1w/kw5xm
AV+r2CknhgNhZ2ynCGxRrbcU6XEfVok1e00SodCekYyLmFttxEiewdjwkNLjS8at7EdLhlD7O6Ce
lNGUR/fLfCcTG1IUn/j5y/+v/bmSnD0+AnnLGcqG5T5wPppjjEaA4cbk8VS5Puttl8qcpLk/WijE
Xb/5pfVngvyT00d50GANdSloeLQny3KeITZFHkeszC1fCKvP9vwZqazcvfK7qmlEyCrL3dIZrnzw
vjjOQSxd4PnqElAD4SVUA77KvfAuIJo0DOtyMQjFNfGsdGWmh8mqgwGwxup5P3QywE6seNVUoHI3
qvJVZ5k3y2E/zu/dXG0p3FFyHmwISk4sPJ1esohakEOoNh/5SyIWIrpZKoF85tgaJTsjiHoehnBy
8tjUF3qVXUMMF94QaguP3MU+nR3wvEJvga8wScYpyLur4gyzSmUg7kAOmXnNf+K3oCbafd0Ae9eT
V4jKIlyQRLsNE8rHHb1fHy1k9Kxjt7ENkx2U3/9CS6PlJvD1+1+A1vtZfXFoLz9Pzwu1yCHDlHan
k2r1CbEm7QXDMy16kno97wnDdAxEBWB0mf6lxfB4hq7iP3XIkoTgKL0VKcZEomh/+lfkciGusKBe
RhKQkkR8CjAopr016BerPcA+GAPfzGEQL3fNagBcZeIDoaiptJOOqJHcs4GtObkALCNH59a82Fg9
yMJ4EbaDzcBEi+5IcxdSxgsvCHBIz4/+bcs3Z71CFM7ANcWaVJGMw2Sr3gZMtDa1EK2zdANt2hqT
gPMs/zh6oAQGEgWWKESAdU80piRJqdA5f9azPFs6uxW4mlMjO1p1vhud/tfOAXRqTvtrwolGwnnc
Xqc0d8ILk97l9t4I5V5xEy5hWhQ6U2fafiVnCqzeZFmTSiP/6OIenGa/mQKKu+Jh70+7UJ5FP1w9
oiHtqAZYTZw4TV1NPJDDVyRrXztT7jNpQJ36Ualmwmw1fZ5Q144su3AxTs0c2ebPoX2HUu/PNhWF
+h+zhJ2F42h5PM2kpD7iB6pU751rTxWMGuqcyQgFc5/+A98xzgXFv1ZMBIQmdd2lfP5y+QWY1Trk
4vLjnyQBZhD+AvmfBrV4RYbXS6BwweoPmRF8EDpYcSMmzPuqzKk6nWDutVzkIVqkQ4r+V8orRBFK
T5w8tYa/SASa5ZBCpYCxP8MCNyiBH/AukJMp5p0d3dVFsEpHI0KOoayJNRT0zIA3h5Q9RKwEwshY
moHivN3zxjrvO83jtxr/wpcCpCYAMbEdDFbIDC8aVHxxb+8GTEayzbB0nP+mSaE6yNRWKvCRj+oD
r1ebRRMe4AFYK8kIWZTYw6l2AGXld/d+v/1LjPzELQJIIEg/BDGGlpUbW6fxlOV9kA47lFH8sqdD
D5MKXab6JjwIhM4rnlHAHfrR9sBo/86wFmwQvYm5Jog41Vg9gjmeFdY5IRI3XrnNSaj3Bs7bTDtC
7xb/roGPyY60HKdFvBpY+QRw24qD7l9vLHsPnuyu/G2LT0bdDMUc4mUzYv9YbHtixGiAu40YfppO
7rIo90r++sWTcAI6C5jl0LCSLMRQzDV8GEMjV2m9oNonLif9/uButJT4F5YMTqtaIqGUIckU5QpW
adthrFVizOCcgdu+qREKTCtnSXg8kpLhlxjQAuEXH2Vpnf+z88Ck7NUhAbgoCvLgqdWYrAYfJYs0
Pgud/TeZG0GMDOjSOmKs1EaagP3KBuL6tDyL5ZJNonoLBNmHC2kYt16X3p0Md6xEhXFGeyjHtgIm
mn/YHJGEe6/3BFdetLZYTgVijQkP6GkItCJzFUYSohVCEgOMOL3cU6WRArn9f+9qRUKG5UAO0KRq
PtZ6MTGzBjXjh3JiIil0Hc7+YssSWJLZ1ZWn5kkt0ewMbGO4PWMJLt+8k5fKlYO6tbBUYvMcSwbV
KWgkLXeiu8wYNJxOXHfTiXYCqiECqpzU/3UoVbNpl3e2uXe5tlLMet48mL3Qgc9yMLSUxfyIdnfl
fTrSOnh0LuNe7VA+OZa1WtO0PCkuha3j9klCEMIacODTrO4JBf6ty+3Txvq8nl5sf8poqJPRvSoa
1SMlwd2otn6a1BOjq8BGjA+sIeSnvNiMgTJC0S60IuoVj5x9JgaFoWAZzSGBygqA/vhvlVPGWg3D
5QktjMR6iVoSeDHRoch9PrcYyA2tTUSB78LyJUO/VcetXFIk/PKm6Cz5RPWVGfhsUdDETM6BHaR0
2GDm9grO6g+UoeEf8a+9KPEXkq19lR4X11ZBrBt0keklrScD5AjYB+Tj5GwjXPW9fzEYOq1FOq8j
Aia7fMx8lRY1vanCZZe7ooNj677OGCuYCDM/WGcnR5GSXgXJbhKI2AtcTwS/qwABi544MXRnrnWf
4lpuVf0rkY0qmLApyp4UcoQbZ3mhlo2FbGaR2fzrSAclNNVbQe4HcBLwU4aiPILVyIRjzeiLrO87
qJkeC7Z1OuH8QbbazIcrY235iRV/qM6EF9xJr+WBteqgPTiUAEc01otDqO3ArBboxy3BDAcIv7cD
htZ7L9PBvlkagdimznbz8ntFd6UzEscfFLja5HGckLtMEvPBiRDhupUJ6LXGMtxCLyLkstOGLiKO
HN26nl8a7txMJKOPg5I3vKh3MM6pe9e5LYJ8YhW8uGi0KYx7g5ZYSMhcFEl6hMDG4NQbexF+S2k0
5M5iBVC5VEagAh7kXAvwza0vw1wAlKxbmeKMfrjPu/MnSklmXUvw9E+x+CIgfBFJiopwhZfvoJDT
Dggl8b0xS0dj3WsVP4onDDHBCkGre0xsJP8i7bh7ERiuNTaPN4qSEBrysC1ssXjhcfBDfaLN60V6
V5i1GgIz2UgrcKYOMYdjW4giyUBYODRH97DCZVQAE6fxA23MgRCvHDzbGGPcV487h5/PWCNFb34v
Hg6Xe1bv2ke96sqscNE37WV5ZXPOtNv2lXnItkZP7T2NgYxGb3RrTDY7+PkWeXjeYWAxlwfhDlC3
UD795XCpppwySc51rhQyjsb2pDhfW6bgsZ74PpKb/FCHTVmJer70uC/0B9f1f7y1GNbdjvyULECc
fB9RfQWTm2IG09v3NGMU0yejQlQJNNa1GJ3nX1ZW0UohSrJbJ/YCtUMhJMsJ6tlfMAppKh53/e6P
IllcMXUVy3/RlzYwatnHd2FTY05tUfzBupH0Kpmr58tTjA+gJxhS9k3eCHWzr8tBnPhdexEuLKq9
3EyqRoL+ye0lLcuAn3etkg1Pgeel7ZkHbzUCwgZtUz6MnhdDKNpwcpez/KwGERxFoWzOJBR4EQrx
bn+TjIsnheolk0u1Z1/+szwPDrdzW9BZXTS9glY+Zh7ZiChktVoJmheHB8kmdvJjk06DdO2Uh+U5
lKMmQySFFvG4dKNA0rMTtcLE3nWeNFw1U1953FTPzRbBkN5VcykFNY1YWeP0KCOTNlOA6p+3HRVH
w9CupfeSxHfhcmNdeeIXp0anSzkadfjfWmoxKbUx4/+DdNlOgud1MmwGzuDsKnYZKW4judKYltzK
SQ7priZA6TItvzORoKoAiaRXvCEj22zFuFux1K+i13XbIXfNhJ9byorp1Yv7hQyfFdUeO9+/mCz5
hJhujkReqfGb8Rja3sgXsHUavVWzhfbYMzT/1z8AIPSk6pdT/m3mdlSkztptMQnDLpKnVLfSx3he
Jyh33a91O80Z8ubk07/eIHTR0MZP0fZW71JJRIIUufilXdMdlg8riLL1/6WXtxVxHk5SqEsX0jJh
p41pcl6XIIC5Ho12n5N5m3WDQfhywW0M0XiORKUD+5felbys3Mq5Dj/no4Ayg0y62lem84voWCAk
VGq84zK7hJwUJSabnzmLCF/ZFjLa37UgKlcBWHnNRVADNcfctYDwTdJiaLUmSrOIvC+Ns/OYnoqr
SuAiF5VYElailnrnwOqEVjWn+j6fbnE83IeuyQdFevrJVoLRlFcClBjsciaIP+KWIst6e85k7MLg
Xhf0fPi5GApPAk89lNosHkoydPWWdLs0c39irkc4dxCkJkw9U3WZdSYrTbwEOe+EAkselOjeV5Gy
0ukrowj4Jk9zuTiH0dBp099wpSaMbk2y2sTivFAuf2yiwKhndHLHV7vDqulniexZod7zFznuwXGq
F49H6PWqtATTcY7JrVWDEAqRNGsP2uR7WcfnxWRaup+W7ATH6AY8RT2+iCasMhszeGZ6IkXASh0O
NYnX0LSzOg17NA2+sJYvU5J15krxj9iG1bSdJRN5PBRiJvPBWEu3zAOP6X6nv3udHl508SFYrfsl
tRwoB+xYPBCp5T8ccbTw27KqYwuAfTyTEzlk97Mno3ZzB109Y0r9rduINSLAebekhO4XYIsDokYb
FWEbSHlxRqz+cIsL5Km2JnTrHLE7YQ54BqVgOSlMvKGWpP1omnDghoLqaVPH/UEQZ7WEdm4eLDZq
1Igui5vl8J6acWHxnC9hrQ+kjlu+vGq9M2u9OCpq4ql1U5hAqEVhECroiGKVRUqB5Cnr1taBN3ia
2P+8Ufgeacv7tdZXpLz1WDUvABwEjnwL5dbtaVbjbQPecsRrJ3cvSpS9MLp5eS3t1XKUHfCKhsPJ
DhRwa78oiIBUAeNlvnA37XAe4dzHlpOKMQ3Hp0rFa62V35ctQzV1laG5gmzh79dkIPzc11qz79jP
7bVZuMX6nny1gES2gt31UhTFsWijsY4R7O0tvws9N4sEZXm4Y8/a1CtYwtDClKmqaz8kwxSezGIv
sfRBqhCPN35YakSjk+do11KLfced0YSu/8H2nQJ2og9HcnR50VBtDsCYcz7ja6pfuWQDNtNQOX67
Z9hy3Gt5SWgixS0X153E0evaWtHX4rwhz63mqkTwHR2qCHZioknwJX0xg9YpZV7gkEoqXl05dFt4
jLOLbTfyLINcFKEbpvt85E/c0EdNtTaC0j3SKY+LCEKXpU5AArm6VyVgbouc2AVkj8hZm+QyZOJN
mhxMkvpH6kvyjuHEh2zoAFaAItIkzu+Vim6HYMGv1GkZM0/vJKnXGWUsVmlbbEw/BUE1UM8LhGVj
iapP0H5shZbSuY+YnvpkPwYb3BOuDntvXu77czMM92JM7jynSZdoYAOgFhX56oLef6bSzgPWtU3S
eB09Nx6SsTvrLNW1MIIQnCi3SG3Oz/WifEoCQCkLN3ywBIc8/3ddzx8TYB9kQHDusGYzwW1BROrY
GrC9YQTWCDZY+x2pBgfUFcaZ1CKgckkEYHTJ/87NsMgKt/iETEkSja9p0p6m6kvIMzZiaXvlUuhb
gCCD12rgOMprX/gnuz+oHR3phpmBNLPrgLSzS6AqkRuGWs9kkIbu7Z+l8ThjGCNgNix+YGnjaLXt
RggWmBsm8MmWE7WlpjgZ0s/zDrcz7heghwQHloHlkf8y6YoodM8dSBYrMxreUBAc2uKk8ekemGxp
tXAjlfqxiqB7KgIPM9CuCGHQdtPKrplQ2i/vBulBFwCgE3Z3xQ9MTesuEAnQKlkGCUnSDQlJy7nY
SqYIht6Vexb2J4oyqpstfdXKjZ4ZT3RvymE4jwMbWq/FL33lq8vVAU9lzl1JiCV4VLPvr5iDG70j
RYrHDA2/OuQtl8FBfUgBxqARf+X1FSfydQdsT5rJv5vjy2euFg57zsTvYVBFXm7EZrIdB6PbdiQW
fibHMmydGKyG3I0gY/L1ZC/szFbE1QADaKd9TIyqSla41Eil0wRSvlstFYTGcTOyOzJqta+qdD5T
wbnY3M+vTPojiaYIw2MEFCKlAX0tHKRDQanTrpRWiHe+aAtFCByagi3iHv7CFvlMYMFl8esJC3RL
QDZUmlu/YDNs4pIEb6bOEp9KS2jH5Cs5HbX7UJO2W0/it7D2fGZpP58947WMETgQ365+jBRpk5Nf
8SIp9ujJtyjORcc6fT1x4+nu6sMMAkdG3ZVrhLF5ViQufb5Zzjhkjw/VaB45OA29UR2ET8HAMkrg
cidkei0GjZWJ1/6Ai6bX0nAg0FP7ZcbdzeBPV17Qk2Mg67Wtg/04Ep9WcJj4Nj9PlpVNPvYxfUGi
dsXfRl3kqHtYUzRS2IH7jORLya3ZLGK5TmpJWa+F3pCJQT0druXW/PFcbw1PM9dpwMY4h0xyUu0e
HJ3ReAPJ1+V7ZHzeLOc7LdQHsCCW9TvYk7jPJkaBDSPPer/PNtTQMYf1cXEQjXZ86RLNNbavgEDA
Vm10eA2zSVLqclQhQvrrgi0w6A2elN30aUj27fIueQmRaZTOiiIQHvdgD/ivKc8Wmm47gI6HvHm+
ASf7eCBo7Y1uAGRnpG8qrkIGK05KBIoDgDLJuiPW9adzd8tm46VVJ8lkJIExb/rP4LXHf6bTnfns
IfZGo+c5yTs/Q3+8to59nUI4++cqTWxu/8xMjLTIGxDETKNtwW6Z6FLz1J8d8kgMbNrJUhQ5cUa2
cEFjk3rr5dVgWte+q68TmYK/f8Wi9WqtBWh0pCETrt2NTAw5NfwxyRBKOskEYQf94r9/lTqTbUEE
HHCJ3F0Gb+Sy5qTSAsmrfTQu/Hf9Ou11FkswlH3sadNF2uJfrbs0EI9efsN4hODOSFJiF5SrV5dp
Rtz11qd1l4Oa7O+Wpht9ZMyIQerDtRpjVYloqG5FMWeGvuegFpOJvUu/rfddDPRmEHeH5EyfY97n
huOZguflmJ1MEF3bz3zE9u2qo94t8gLZrzUamJUKFyqFVakNhxrMEqHs9cdG8y+y4E9Y3u0TgX+A
V8tUnNgu8bHTrqWwvKA7yKwleZys7blPvdCxfDQb3EWlFQdzygqt5gWBirdcryLdQRjI6g0XyERZ
hqq8b3gVsQQPgmZ1hPs7pK2yEcJvwrxpHHKdGU/AhLuYWewOWt/XUErur/tXymij594zfuKqw/An
SFpujBUzUqp27vNpxIpymv4FB7JP+9Ks79UNnzuvU6HQuCGqLL6blYVafo/MrKFsZImnvDnu2Jb2
HpnQx7soW0tKLxXr6wgbcjYOxlwM9OgLc3RMa54wvNX88imkiT7Ps/kevuHCRH8UVQ3syX5sXFmR
31AKv2yhSdxwJ5iWO5heqBJxDDh34WFPQjZtSpus7cZUI2szoz3VQlXTCMoNp6wFheTv/A40mofz
xD56lNeCUyzIZ4rpGp49ntK7PpjemmJYuAeCcKJP4UBiadxA/Bs8ynBBCRnv2FXKkTW9LjLJRstg
MH8Yk5KafXbd4PS57R3MoqgUR3xIhNbt2ufhzQ6UxeQU4kiAd4bV9V9YgavHRgQudi78RedekktP
mg7p0QHExVl7ztwOSnI2zVzG+X8Ve0HfaenM5lj0ZnAceMj8AKuWISiKScghXjNriDI2YhyJ8kcL
oFUHKOEhQfGy/A/a2LyL2VZ0rOWT1HjNiZiXSPoAZuXgS07IecQub57OxI0itStnH3vv4tFutKge
fe6rniO2yA5zcQkpx4s8xKl8j8SUkQrt0oa2gRwrXt51wa0mmYc+4mU8dewg7H27Zs3rcPSATOgH
cckXtsCEY9dUBmNR7ra+sjp5c5Gq5hhpoDsVqZAJD/ieOghzS1Zx9sf8xM4GGuF9TAAS7LtncEJg
wgSO6RHrgAvFaDNyEfGm4Sb08NT70xws8bI+L+6QVMu+F3x8U3+GETKP4eVEjvUmkktz8ZIHG7E1
VDv0ElnBdkO7g617c1/EwZ2Ss8nE1OQZXTuEUlKkdrkPFF/63G98cb5tdb//SJd7C7kW1OwYOmlh
fEJLfWdGgLpom2RrZbvfOq/7UVethUuQOLnXPBh9C2LNsKdqqA+/38xYYYomonnwm1jECpk+ww6L
noudDYFNiCdMmrfj2tUwUEMr6/61L9f24SypPo7rxYxA27aOtTHKscs0Cu2kUR5UJfVvIqZmKGUr
cwHzDlI17hQxeNaPpBCojeslZXFwHJZ9BQAjlMQHEkXpQRIURRjBiabnuLFDc3nuL9OdirGkB4yg
1/UFkMtbLjCFJx4Ia51Pb+w86++rT3nHhZ1wVDBdO0ZgAT+y+8PrehtTLx3ayfjAWpAOFjiZN5cq
a6cyBccq2TB39PI/PX5stlIwUv5Gw75E7/LpDVLuB12uq2iEy0RPXnNh87PiUGT9uOtaVDL2+bGt
vSWY+0lOckwFAIRg036FkbiY3wT8hp58ujLqj2HG/VAEpDnVGWIoVefaS7BdqNnl8lue7Vg7mFu3
teCvTuX7eWQdHYsGv03ldZccxu3jYvac/aAAipYWzKJ0hgU/lZjo8IrO2JEKYtNIM2WYxrBl+aC3
KxzztHAfwouyySM+4b2K5fLKblQ4khms0DFY6Kq96xcKRGFPoz89bHHNxKAK1BWip6Ko0jsN3mch
1s+l6ZMRsVFiHYrWRFyece8Ws0/czt0vAoVz4VMXaqML66f2rf/wpO/HvAA5lXzHCKP8xyQi3bau
i6q+cpzYe4sw4dQCqfb9mDERnkQhe2vjoUpcYjj6KUoY09XRZ7/p0G/6RFlXj/DmAnm6Ee09iLLs
F0H/0Si2jnqirNqA9XgcbxY6CooNMpEPD4B4D5rEhQ5tUwbTkgkKm/Cc4FOLjiMd4G7t+wrDdfOF
4lee141vhFxKFcHr0wY60Ld3I2hk0bLR0Z7AlqSiaTVPkYXeZnU/X+LizlKVL6Uox9zqWgrK223c
e+9d7nl4wlnPBEFDt/eD7ExVTzrlcgFTXtqzUdiB9LhR4A4NGFe/cru3ya/PpL4//xVZjo7viVUP
bhX7UIlRlYZ7J2c4YwIVOBh6azIw5Wsvydp1fZpZQ/zn0X2xWPuD976y4BLd6JHeYjnOcvK41weD
Wn3FY4Gj/0epFfVJ9CyO1Q7in0B/p5elMk97lJRa+R01cS/4CKsPmn0AljwlsdvLzgui+dqwEpRn
IR1UCyBupNm5C8TEFM5KG8lk//4I2ndUfRILte4OGuKlHYCk19tByIHdoeUTscI8lUeE+olKExMj
7XsHz/g+Nlr5WfvsPRLeIBRoTDms0oDx/urgMeKbOb1oRu+CPAcuTWJ1ViGnAdxXqvwRX+dpLMd3
epXLp6sNhBUkPqZCNBthGOEOopTr/ffBanSouyJb+K1pqhn6FIi/Pf/HWOESLkt9cGMLD0rABe+U
p1MreTPxh2MVIIh+siIgJZfhaegNlALZ49XfvlUc35aoJy/FDi503ybdXjRlOTBcmjxab6Ib5g3L
WkVjINeX4MWIlcXpibWjYTzFBzqyah/JscngBS/Gsrp1aYkgFHl0x0svwdJ3CHuaA/l5CNFqyfNC
XV6nEaA/ZSXs53ChJNTdiVCnragPK5IO8zerp5KFYSOHcrYLduLNZl5v2m6lX4iTbqG11bC0SlD4
nGrHdyK+j1x+5FC3DTl49lS6b52RZnHsWdx/Te6u5FokqB60rsxCKHpNrTUwpNQBMqHXtIaMcz4T
V+6/+XHnwLaqNFhjB6kMgGHUo4aK7jV7vEkLcjrnJB5SCNgIG9YRCVLKMME2zHEfA5lK9f8kRWD5
yNJkSqVFIC2Jzzx4vwROLVPU4l8wa54ucSynOVcaJF85tO+c97OOk+pAImJAAQadUt+eK4QqVypv
Ma6Q2SVjeIABeO4jo06WdifOds7SEOyd3XEURagxqgfTMNgTY5868xoVwczsq0pMzwhQC3fI0Cab
UW277YqwtqJB3mivrGuiwNaAEOz0hgTm2mDmpVIADdjUIkFx+IOEifbpVgD8GxBtLsI1E61MnVS4
BsCqbk+hST+ONEIH17MoRZFj7PmqVOQgDnnVc6hTmdTqRDI5DgQYEsWPPvedJHWYFGIuITJYHCpg
TVVFYv1iaWZ/P4KBbMpA71MRDUxmvyNPtZYD0uVYZbl4uVXL/n43aNdvF1NntPLxrGsEdn8HphSl
AvHUFLw5gmU0OB3m4XVhLprAdxvRmOKfAVhezWOthYp9V/5KB7BocbkUY0Wh7nZ2+N6uip0iW4Sy
QXbR7ZgWqvo5qGB6MuhiEw9KfwBM1gc/w8aO7W1kXWUfYKXsuouoVMuaVPYM710UR8/L9IiLjdrU
7VYKQVMxup3xwukc6s9o+mAMPDBkkaTpqKIcVer9YknBYG6vGr2P+KmSwXxxStX2X5BNJ94AmYhw
GowhUNXLH9qt2TlQ0AmmcO47HoI+5+TdiPh0OICM34/r7urcPf3KRLbYrk7utdFf2iWnhFbq8n70
f+aZIJyIHgbc24Fmo1NNZvig2RRi2F9V/7IoNw+6vnV1w8I1p4upT+4U63BcI4FroQS4+i4aUZ78
yk69RXuqzL8b4Xjm4ETdBuUve21u3iutSfHNT0HN4q67RNla0b4O7QAhpJ00L/WTFxSy+Z/1bNUg
WE2ux+aQRjDVLZxAGWpedKNoL11wVvcUNBlep5lTI1Aa+5TP2vP4VksDHvFll+3lzvkRohuUZQUQ
zQlsYYls7LLg8yQtUXDXdP+HAO3SsNtAJpNdUVHSk1DpF32/cH3ncSDwYSQfXCHwG4MSZnmLARO0
zrzx9MgOH2K53ckc4tc+oLd623QG8LEpFfQg7F6oQfLQC6LkI6XICRb6gUGp9d4504ixCsxxSVAp
yRg1TJJG0XZj/SZIytgaZcrcBaIVy0qRDHXs/EplboilcJB/Eec6l157iiuj8k19MatMOGcZzPwi
cZdvSnUs8648bDsobV5W7R8hUBOERbOdazePA0XxUwnkRGlcd+1zT1Brmh0VNf4wPLVWwvlosYaG
eKmhmHNAMf5WSE4BTEtY49th3RLYYfzwoMuuiIBRoXYYgmSYaksHFaQZNza8wO/F5BDsJWRAG+c6
BN6KGqOlYDEdM1CWsDVDyYllEZ4GefVjhTfHc+vDDdtHFQDYbVlrHDKUSnt7LS0Co1I4MjbL8Hke
DzGvuCPgDzdrj4kEvNalSLs+1d1NfCjRbQNeK76UOTP4dPiJ/lzGybFot3MyZ1/dZEDSCZ8oguXL
GxjgzPS/+Ft11Kn/OUrXE5GYWi7YFOTtoI+w0mZaOwiR6y4ZxfWIS11Zu65LOCLf7oGhCD90PIR9
QAipuBDED58fVcrRJGPoHnQLSNqfHBP/Xn0DK0M1BwKGftXvflAYo3AWcT40R+77UFiwslpwTrFQ
6tAt6nsXJBykSQ2tWuhdtrDWR5DzFmlgNB+TF4wo+EqWN1RXkKH27UmGbHDbWiTvqbiL6TBu2+xc
3s+WojQRw1csZXo3rLgk7N95ok/wbyU54rVpck+AaH9N/afwCJIQ4mMAlHtK35CQ7S+t2Weo+BgK
v1HL1Uu7RJSc/zGtWo0J1ujyNd73LdPGpkDRehC3n695npMlgU286AcCvXgTlvLZS6laXd7KvjWl
2T/ULg465rMYND+e+LxpraWhXSS0JdAfNoQHTuHm3kLM/FNkMXhOa6EZJuDt5kqmKKqv8oKBVCCe
oi8JxzMqRKh9CO2QcPGP26cQc7T9G/5BWkXruumPQ89x++PDsOasaiyhm/IepGsoOJbw0XbpsGMM
pXsv2hPccQVNmdu+BMh7RteXzGGo2LzfMq2R2bpwpwHGmCIL8RSLVhj2f5H7SHZMmHkV6hoHqAUd
YVlDxJ0ZM08GgqjZPeg2TEk21JFnUGIYmx/X8V9SKHJy5SgEhD6fQHc9EETDtxfyIeMo6D0OgKQp
YyFHA9b5DM67vN2sN/RrsPVQo0WBhFJ/Dsxyjr4B5EkAWXdXXUYKRovixi+OrHorDuLWAYSFZulL
ZwdQ2CeIb3dyLsWjrIzd8zinZvrvHhxtpPUd+Fz0Wwcq5nT6/BJDq9c2dTnJ+e/8BsrsvScFLDqt
uo8mxvLq+ny2b+ailbe7vISZuYQ2xreo06O7OkK0LyKmUnaoQ5kKD8FRAGPTrvtMqKfb4/ZHXaUb
gynFXEZDaxbXdb+3kQYg437PENsvXT2DhxwsNDM/p29zycKDqV82ATyMAtjX/FpWICqzEDFb1boE
zO+2Ft6AleFDMankRBAgsjgxDjXvH9W5j2TcG/AXQUqIfM8Cs1CMdZVX+I3MCtf9rtHH+Z+MkXv4
Jdi5vFkjzGAKFGyyLCoDA1jLxXzulkFsu0RyfeTTZx3SWbrkfusOFCvDQDtL6td6FT06eegn+FQ1
Hri9oB3VWr2Gw2wIuKoRvz6ruzx6HBgBI8A6XQD845GP5YRmX8QWn+I9JWT8Wui7E66YpSbfoNiK
11HnRa5Yt5apdf1RYlgNWFUP6LGGelLJLWh9mqrgEhkWu+5S7FcBWEp6J2tZYbPe0zmn/wU363dl
K/F1RF8i6v/+MMDGvhiN1NdqnbEhlmW9kwi5NcoTDFzZiMnHGFc2mGRg7qErDUG9YBLP8Dgd2jS8
P0iJUjDh2re5JCrl4fZqTde+sq4z0qH8cHMFzPITuD47gcoqzS8EYMuedDXf0LpGg5LWC4A42AF2
kLTzxle9fUDjacMIf9utoFelnLTvKcE++tiHJ30jOsb2ySTMCJ81GKk0Gl7pNN9aGDuJHYIfOLS7
ch87cSEA/ygWaIw0/tIDaNC7zeLWh2FbGlgs4OIVf1N82rV0DaTzvjdoFQRKVGYmUzpfuTUBgejD
3u2fgb1yn23AObywu0bVmJs4/pw/lZIuBUS1vFhifa9qsT7Pu7l5JxYHHhhmFLgZ2V5L8PDPOH0/
jbuqxTomtTGmKN/S2ZWdFt1cFvWVjmCRWaSEGlgvb0ZQtT6xNEq5rN/3re462ipIQGGzPjHk7/Lk
ygp+LsDVX+VD458i2+U5LcI4x2phiincd7iGJy3hLvVh32YiTn4ZWnIEFF/eGdfOnnDsQ0eCNjo7
KACtA9lLMLLxwSYnUP/AweMHY7hX9QwI9mJ9f9Ki2owYKlbesnRS6Tvxpc7F3POK0/GppKhGYQzT
EpQVWwzz8f8PSftpA0W6zv+wApIqpk8YpLOlGZMpKnaFcqGlV20WHuiDxQPdMdstDBEwt9h6R1Ia
MDPmbCgqRoe4UqV5KVCtMFgvkHjthND9I6St4ZJ/fagqEwNt2u/HiGCZMtwHPd6m9xUBuz9VLujz
96Qg72QVKyyu4uSt/LaexDo8v/EutfOQEpXrpvyeFmzJkVmkfXCJq++Jpp/hXFCmo0vTZ1e6ANrQ
JSPoOlKYGxXTVX6cie811030nBp0dOmhY9CmNoCgiGkGS7kyY62O5ilh9tuxH0wQxvm6Y6OE4vEa
KAKe6Y7Ax0WLTowEtrbyPa7pnOPylREUxlWmdoXaoajatifeIKEdT/bFTh9VLA27rbGw5bDB1pox
XkyxcPhXsb2BgC2+d46cXQpn0Xm617vNPHp9cBzhp6jgx9dBTVKSwy96OZF8QoHfwgWIYvZL88j4
p5cD7m9wPWjXE5/X4+UhTRYhKL57HEEXysO/6oJk8bKTeNiaAG1ncQff/pNacA+FBjgJE5IfXVTQ
yklFlYA3PDwTndF2hDwEwqhI/XfKAy/JS2WA0OWdUIr96/+eIRCRVxdRSOzocwBwC0WlF2oLmWHq
o+EICy+bp00OG4dON0ioQfi/kDG2ceSQeyvnxRsZwVw6mHNQEBiorKljJzCDvljMtAtgBmKvD5X1
h7YfQo0l6IXfzVI3N/7l8Diw99+3DW9oqqgW2M8FtUuSUmJ4qTVEN5Yt9Xj68sqnfw6YF8V6piYV
mXZ91OFQIpopArVtxpaMRS3L0sfH1MCE7NMpurZDF8OI8bc5+g9gOgARRy4c/v6YfyP7MoPo5l4L
dJDaZo2CAsVhLYfIkIk4cR857bFXh8SMGgXGqLx0NpuVa7yVpryZxF7matxxXa0+cEHFJtBQZOJG
bcelCPYruLomg1upMfDjdL06uPv3pcrjJkYBdKQ5T6c6QLY0UIytlHfEUL234VRqd6OC/ZAMkCMw
TjAUNbBLtSA/IP13h0MmgDMcY6SADXO2kOd9Bf5XKoQBhtJ4tGuewKJS0yVwm5Wdy33aLtPwOHuo
GaIyJCrjHGriw4qTK8maLTlxoKiHRnFewzpUSJemsaXx3doUZJ1tbED7YZT2vRh7x2ak2w22SY1D
ecgHd8RAorvb8D4xio5Cv4IfSG457ADBGUouV70zJGyaGV2hjd+HgCmlK9bA8SGDgK7MsIxoA3CD
dijl3rWIceqT0Csv5Bo4gl/Wfn7xTinegsKf2neCcuH3bxFZBNxOHolrApwzMRkWPjoRRkO9Hw+m
ec6NtL9PbYgRy0v6/aDO6XJWfc8SudI6oRyZH9JMFV6GGwdV7Pr7bBEr0yZ/oD1pWtYk5YhXjWlE
xh1JzaGdYRuqqBBxDutgziHQeve0Kh9A06i5XinsT0zhOTVJxicYdORdLqD/yLtNO05iBPkT9jAq
e/WgNbJVEguGZ8I+7VlMZHxhkm7CTlFXfoPZ/cXLXrMCdVx2QMNjZAuxPSzZPy/VOa9Yd9sIJWk+
WoSxmkuUkxViCHQ8oam4H4Z3camYQUtYpiAUvf5XJNEiF82zLcR/RvBTQTjTLkmTP+hp0Qkbp6Nm
O8YaHWL5pRUoRkcjLAdsYGtP6b6WbwrvJ85ukquVpMsxYR6IBgQURWPxtbz1dLItTZ0ns8y6POM3
rnYGfBuNbA2lBmIo/AngzMEcA3Dl7blWV9Qa4eZ4S92G7iUcjbG8xR7iF0EazxcJbd6z3N0KeuQ8
USiaUib2BjM7UfmZNz5K4gWgJjCchI9vCQhl2o2ATiG0rE2DvQ6WIL8ef2C4zzOrmyggIlKz9GsA
A78m75DELeY0+6/ySumGTuA4OoQHi3/b1+pOHn8Chmg2YWmHesmfTvRmAEGzw84NaYaG0eB0TYP2
ZOq6xDlQrCK2QTnJFtmAujyS/vdVGNl5/swdoXxTBCo8X594WKg4E1/Am9JBgLkYWbSdPNESpUBj
Df7amJXRnZYXuXGKcMBI9GwT4OqkjbxZW20P0XLH27NmlXCs+o7QsOCEYnQHWAf/P4vMM2fg/kTj
ZaXQoLP5TzQ0QVZv7D/YV017FCBc2/EsJ5Y9XJwNUKBzV2DRO8HGvResMmiwE55XV1IP6XZMYby8
EATbAma5xNhWZbPQo5IwlVQxJyzNAWLe4kZuegkHKbVaYcvbcoxdxf1Cc3EPcSuGsPx2PsZNFCUi
m5uBntgaHHk3RDpo+pMNY5cisYsrEASgDBC47a6Al5k1elWHOy2x5DWNFrO5aCWy/frgvjkkMlar
pxizW+AyX8LLcLtVlyxUf4UkiRaAqMosaPbPbwLQIdF/qdp8OMPDHIcaIAJqg6GLk3vLKMid9D2N
NcGa8i/tOp2F6vixAOGQcuATD6hjUrKzvHNeOTaAq6a95uj9eAtyOoUpmhtfWFHcgrpdmBjdcBAQ
T8UlS/i+zXutgXu4zmQkj0H9NsKoZF08rZ1UPP993LOuLdRTFO7zFIHcKi3SPYzTl5ZuQ/tsclgd
hLRJzJRTyEENOw8S31YiVVYSE3Lc2gHTTvCwvL8Fv3Y7pDFvJKmBnwU4NDipFXSQNQepLWMw8Ayx
JVpl+ScB3lFSPHY15KmGD/Pg7ovOkJ96Nw9pQx+lAucA0i3E5Wqdnu1lgp8bAVWP5cdz6ubTBTbB
LsizEbGBFgBA1thNAu7yNdsAQSTIPODPrFLvsz8e344T5p81WBcdnvEXx2wTqjeGrFOkJiaxyf7A
vXnqDs8B4PHWC4abH/AQUJuSbSGDzOb7LHcu/097s6MtG88gzubSQoLsEkVsjSK9VCviDi2mm/jd
rc7z12L7UeWEwPVMlIMBgk+RCR1DRih9p/JZNoU0nqiMNNyBrYU8kk4fdzrWUwsMIwLoHgU51c+U
PK6m/yup890GuZPf15lP1k/3Ptu0YLJIRUMRrNFjc83hYNoYY2jlB6FwkRS3YZmDL2NL0GjwlvW5
lGs+/2Bae0FgdL20jenkN0zi1zFqCozSKTjUSRAxEuqgWydNCkn3sjbrM/4ZIYnFEjS50kJVelJq
ygaQGo4CUYQoLkHcmXsWbXn0QN/jWYoUHP4xdbp631D1bBY80x02yEneLJb56borLpiGqiO/4lDa
Vsu4TFW2oxOA2ti401xyqNpme93yjuS8IconTq/6Fz+MC9s0RHTb+JyHF40oPkkH9tcVVyrXAQ/m
XT2ajEGi3SF3Yr3MSdu7GnpJrpThF0t/zuxKWKX7dcK327z1FafQP6lQW3aBuSMV9VxsoALxRmjQ
x3wVRGyNTDLMfupFLrOzGK28GEbBQezXuLbwUH38wZCHybPHadV48jBj1Yp/823S06OGr2JluhK2
mdSukdwf4DJDdkhwh8xh0NkZii8uijOUBLNBZX0mfLiLFbucZLQpY3a4dbj9Gds3wjZBgrKhH17D
JxOufZB0Gyp6CFR9pQ9GNQGPVl+qqpcW1+js2LXOZZQEWyB58GXPTZBu8JfWO4pEMwEkOF5vEaVz
sb5+TpqahJvZkWfSCqHwjXDJIseQ5tJtlvQ6NjFEkByI4uIBnlTeysKPn3Y8Qty4p+S5sOEiWgST
3Bl6Of+n3SA0lWG8kpp3Emaa3oo3Ir0q8IZMYKPM4KTkMSnOLwhzxh0VILIOyaRB/EviSZ4zVVt/
KCj6kHAqUjsQceTZDPuqj4jpRBA2DDwcdB4js5rzQJx+WH0OJ9zS98yWT0w7B1dP1qdNmguJbY6u
zGA8EsP80eOuJTQNc+UFSgVd6pomYEhFeCsaiFODXM8hm2CnJ92qCv5qpfm0et5ZkR0XiddwsjLh
CjUYzoUqsD9RvL7DAEXyiCxr2fuYsSL/XkndHEjsWYqubQnfntDnpSnEVT9H9ZL/EWjbECbkfelZ
yM6vfZevoxpNP62qoCBNRpS9ddc0rYnCBGZ7Fh1jtcd5rme4GfvHzRf4UyobKcMhLZZQHOOzkVap
7kEGJ8pqiPAf+qpl1xDw1kJtt3nEF6gQVaCM3pwrIave4IxQbNpre2/g5QjtcpCveqShdyIBP2aY
fFdRC/IeB/M2ii8I6HFwEtYmd4bqCTKwLAZCJrUmtuJqtYvC/P5XThHcPta6EKB0WEGscsgxUr9T
jHLGdwdL1HejMcBapowJKLW6aVCksa0KitBsXhlLDyINiK0UdToXCsBlltKKcMXqudQyNZ1lzTk5
IXUsdh5xjaxgyo4QgnDLGrw17wKP3qTVzLMCLyvAvMDBx3R0Rn+hQsR4GHMp973ACa+8SSzdEaKP
wsOjbdHmycbZ8R0qdBHLxtrGlFpjVF98jpJak/pQVOZuDSx57zPLL0a0R6/6Tx/Stjkd95p8OVgl
JuirzUBUrHQ9+GMmfYzN2ozqO4/MbzhhjQRcJCK3A/uyw7cF5tm1cEPmEOjjAmMf1BsrVPpt0ON0
+YSQ0TOpZUhYYAfWFdXeHIDoZhfquporW/o2AiutBiPybvSFUXXemo8U51mN9BCObc06IKNVlY0G
++/ux6bacuyIDsWI1C5Opm2SRKil2YcMa+ScGsenhPd6mlEKO9LpIqJc1wk+N+3n3JCmT5XVmekL
tPqz3P8KpbCwzvvWEj3MDMPsjAeVBeaJn0CAnexjeNYvH1kUemKvMq5aUi2Fuyl1UomegfMyW/oZ
bKqrzn4LMYk7/mwD1WUr2VP9WX55d1XWd4gHL+btmhlFP3qx856pAykaReHZUBbaFKlQ6qPParII
R0noo3EGp9TMBx45UOdVJUSGtAbXVYVw3MtpJpdKvzWAHuKw+ULbHaBUIGAJG4eWtpsKirnA+cwL
pwg++3H3XVKUd4z3WmYHXfxO5MXyOuigbFdTyWBnOHa9c/B5szrbEYZqtvyfcafJQna/C+8Ct4eV
6KiwtEaxHooOiTWZq8S/AZ/86NdMqcyOz4hgK/qtMiUtJtkjHTnx7Ujyol1Sw5xqEbrAyEZqqIgw
+ateLVlPo+Le8KbGqlL/IEBmXd31guD+riUep5zGl82osD4hSvnz0CSZTDiKnvKshl3MgXBLXYvK
pBdgOOlmuKmJjTvIa45Hd27L6A6mOIEYl6LM3bPJxT2DYrbZ/TZzlXx4a830WL735t9Bw5gqj8rg
HLCxxLL/99JxuJtLtAh5xOdOOAAWJrUapDEt6YYED8EyRwuB19lI/E1VuIj8ECyN0IH/qOpCtzr3
QUio8SWA0MknzznoCH71Wf4zh37SIcyu7hJ60+B1+WL1PvZPTak4nmDZQ+ytk1tkZ8naHVT9WpFN
o64YzugwRmfVrC1f1+5SD6kkzlArJKXANzgCdQ5aihf7pqAgnM/aFYongcrFSO0zR0+YKWuz3JsD
LNqMwOrjZRRBslDyRVGJk4aaqLXXKJMaj28zdJ0qy50FPbqUo35bzNL9eaRvCJkWOStnBN4XM8fb
+WL4B5/27WfGEuxU1i5ThT74n5E80H1TYsnYpZcuuGAJGiWC3uXmGdW5StSrIim6q3lXB4LuY/97
c4aujffPo+RbDEwF6Xmwk6E3f0PO4bMr5nxWOhgcaz3jFyELZEGDE0i2j0IG6KJ5+1Z5m0irETlN
g6E109yxeLX5JgWiF6idEK5F3KMJq7WXnWHQQAsBENgtzEmrN8IZsVmopWGHBn0b4yF6LhzjtMdI
xsRH0VdX8NBwHFgl8ohkCOKnC0BqvRuzckcupsxCcpgOcuU5KygWFG/ABOsHX1s3gLHETRULwD6L
flTFpOlDfwOHIwxaEV0Wb5aWOvz/7flkYueUX8mTP/MeJPH7Bu+CMen4vuenZ2yOAchA10a0kdFt
6PcNCjgc3UNv1XN2OCrgl9ldfmHLlNzmme+zEVdYhJorM4JhQev4FT5iugt1rYSzEoUJLtG2tdpB
UwxPc5072H5JDKZBpzuWvDZMYSQzkjfqeL4LNdVsG6o3FEDFdjUvgVQOAHSXboeD7CXd+7KmQLoh
Rw9uredrp7JD2R6bikfqKVsYIMS+Xd+GMJYTomjHzUyeUnEedlNM30u+gl7NitP0SFM6wZAefNai
5jt/xWmrcgCnxxtRr0Qo5g2XqCVgbYPUiRt1lcq5peD8nH2qIfgWbaLSndvNMXFa+9o+ReA7tM2u
M+BwRRJe9QNnekykiqaSBZOmBqCPU8TFUHRekoGwR++nmw82V5YJJtJ/NLJcFbEZzGb2InhBhiQV
7yKySc43OL+9bCe89wmCaFw4b2v3fiVDD5/JWrWbO27WvimlR2j9mkNMmG/yVw9FHTla6WO4hsl8
csg746xTHHJYXZv3ZrAyBUjoW5mDSFYqDBVKd+B+dKn3v/da7ZlOFSUXLlJB6XMh8Nyx8JUOTduq
blCEgaJBoNxIEHRhOu7C4OmpbJ9PqrjYb0DQR6JJVPEQp4SSw0mS4ujRlMFPt6HGTyxsHOUzSvk4
jVi5J6qBLGL3dFBk10SHjRzZF7dsUU1OFQo+VefmN6hXsh3QmQRAmvz73c//fbSlCCywP/+v87KY
gUeQarLCI/sCfDYKVqOIQKR+DidhMtdiLTYh4bDhki+2G+f98rlTKoAIzI0T2QNlWuj0IA0twE6L
0LW0ob4OwOJtCzA/eRSK8AeiGDqXqUFs0tBwBul2JngyJMWlo5p3vSbhsIhmcO5BjHFUNKNp8/Gl
S3BE+gWE7MKe44BJa8lAKq4ocO88Pq2BNsalc8kbRYSW9DcKjHgzb3mmo58Mc9gm3gvSNbtpAzbO
m0XuFN3czlxQ9D/noYahEZOWLe1QJBSVxcGsNAdYDfYHRljuEyiv2ERcgpUPDXvnzRMMthMNlkFq
5kOMJFIqW+iloVABTwF6Ql377uIor//iZgvhnaEBjMS+h+4sifJjlLI3d+OddmaMz6UV4FVzPzAB
8g4L/St9yzzkhC8T1YIP6iH1IVBHbXSi5mr0r2PAcququDlopiTAPiIYicUQMkJgLGo7Jgk92MXC
G1QJv5GVmZeg6SbuG3adZ8mN74cPUACOqTCPZpecj0elsyFC/ZZ4oHOgm5/PU9P78yzVMKF81W+b
E8U2IgS3bgXmGMI4a/Za+Ub7oZyrgBLuWXb0aiY4yOSAoydhTcgnsLSKdoPREmRaK3SSVuJiEWgV
EM8pDgB8gvyDSeRybrge2dhcQmXUv76XzJNP8zxm2kHE9M8vvZLMLS0Aaadv8ZzWPYNDyp9C/W96
U17GAYAxhPs75uCr4c7+3YYuveW1jXJkv8YnG67fx/XTY03iTqQMWVSUECtUK4P0PHIpfp500y30
HAq0druglpegLT4bU1gLl1jyvO7sT1Apo6tjyLbtDqx+f2LVGhVJtOP7l0bWa/DIqICPlmppPUUe
wW5d8rOE5obL1EcB8fpmZlioRbF0Jho1wYBZ7h+gp2yirCAYOC5vqPz9N+W61GxFUufDaR1l0LX3
hxPGl809bzVZQ9YtBAHxE5Sw8hXoP1E6D9UWjI8BMbvDEKGtu56M7/t7ULR5QOgBX6c7f/6RUYbw
QyNOT7aCVfXxN1GNilLAo/N+aSWiWlx5Dc9ZMIQcsQmi6SVX37hTdx+XceLDNLCTvnUkLR2ZJjBR
Xg5nurSQXkTYzlVGDKk06ctSsnoBD1K7hwpHmcMrgb6BVPbGZUGTjG+hriMjbsF4rjUgEWv8RjXX
A3/XP927iiYlO50/abkghtXYAychBOM+8GeHMJJXI1B9yV1w/t9jgf+mBuFEUhRIE/TKxVopK0+v
/lFWNDm5Kv0jE0j0rOk22LCGo4re7CxiMmbfCP2mIVQW7P8R8j6ct3wtJxVavhMIWuie2eFUJg8t
VrnBuxm9ZO3OFfDH/RgwZM3mOAAK23yySZFFvwdDqPgwF8tSac3rl/4y8CP5L3S9by0jzDjEf2ls
OKjBBkYPGRsokdWG/clFq4/7zUZxF6DJFwTrdWWkIa0LLkAGH9/0V1u/aa/YP0BYFa3gGLh0762Y
vLE60jgMr18WcXBu2HagoJL6TKJxGvD7tomKsp//srkVukfiyAcsT6P9UEnrqTx/rDSAGwVQnvf7
BhQKP85ljlVUR217J75eHhwl+quD5vmj0ipp1xkOIcg3paoCngY683T56ca3SHK8iB5CCwRBaBU+
j8l/TyxQ5Hsev/L+bRX0WnDrax1Q3AUjONWyI7c3NHfSs2Gf2yysMsmoFthlWwmPsYcvsfqicC1R
CGrLhQL43AqGmZsCAOy2T+hlZwZeSOecZlRBNErbd6nFMJROYMRGBSNdD9qmy+Iaic2YweWvtf5i
EA/15GDmJmBC3r8kW5J3nWJ0Kiqm60MQAX02vm6/a4jnReblt5NXxJmjk/r/9dZUKgQpVz4GgkTX
ziWM7+CZ5su+RFMs+t9Y1kjffzmv0EZ7F84D9cAaGk7PVFg75RTKh0lQs1GsE6turs7XR9Pt55j/
WeYE4lVYpVIg74+lkz/gtyk0sKRMgR147M1EfXyeGikz5ARTdSgqlb+4wKRFjCgbXyknT2sHIceU
tA8nqMnMb6r7p9nra+W5OUT+Qp3Do6tg98USjrsrAq2+WGUoxMjcuEWXZ3zsWNfs52I9M1FCPgpg
cAoZKiR+bRj0FJDNnf/x708fwbzXVOldffrbcZq+WBjyVCQOtDhH7eyASfqWHNa3+s98FBK2X+88
N9yDMTXZELMmy+jwFA0ndm/UmS3AebyBLXFaJbNPLuVIf4EFht9VUdlvWFoNMxdRyfGTWR5+JKAI
FP+7CyH/iaIEb0TNn6z3WTuW+wIroA+uheooMIq2yScPUAMAUVJNsgM8JG+3SGUi5yOKzSIdawFA
xULjEJAkeZJeL7qoVBsaPT+TPmsl7DJrOpZFTNKGCvjtRWRyE+6UsEPriBT7dJ8p0cBb6I37V90g
6z8J5WldVUY+oMQ0EBB2JZady3Uerhuv/snU3GDwGrUpzvmw6lvJsRzdNY448dm33+BUFMLiEqA8
/skRmJHsLCxJQZgRDrnbXD1cUZg6v8eiIDqV4mvFWsBAtXLnI9TOa59fRG+glStZ9VGzxoL0v3sR
ks8q+/q4b7GxAT+EXverFjp/IjiWC9aWZharVuwKSam0SWrzQ9LA8xHziQ0OxlV3GU9q6m6hZjR/
Tx9NkoJq7efDomFu96JEIoqzj80LKqgIbXF/mXMbpUYxxyWMIu74e1fnmlshtpzqzolVZ8CzFEG/
X7mYzm/0WuY5dnwzlDsCiUjr4D4yAVMCePZ9zMXPQIa5/brEnfxnnm0mZASh827pwrMpgFzLCrKB
KrfZuQ+bbe4p9oifrEpN+H+u1uN3MkXeh3SEJBVo0RGychVWCHSeSRGuW5Wc71CTUX1aIt9KJOK/
TapfBuKAuhYxT61TNojgAfW5w/46GtmzNezTjyAH6Va8leFpTFO+RHHJg8ot52xRcGPie1HW0GPd
05XIdtlrN8klVZEMDYb9GkSdZ553taVDgFAziZOU9T2QlO41QWBwuTO5Jnsv64ZgZ0SE/zX0B8qn
g4JwyP4ck0L6THrn1kSkE+uzJAZZp7E78JiZdSxdf9xgqJcQjgTYU2cu0d4uSUTdfanVtvkc9s8+
f2gr8UIuig9eumXOPLf4vDFJX+Cb8RClBl6OLuSmm5KB4FkUATVOeoOBaCovPxgyMnM7G73qK3EL
T1pcsfRc7b1d4pGt4yFUEhRnRq/LBurXoTo+3R4uKinWAX5kSlJktZiXgk0rm+rJEypmHujYKhGi
hW/69dHJ3YbDPo+Z8fQRSXCKpt0t0/QWgwECqDbF0ao3GZZ+TnSl723oeeM9vP43FDpZpQoTCJ/k
fFLFZILR6nB+Mkbd2B+fhOvtLrDpYkHtLoB0HSabIB9vQjQxRjP5HD4J/lg+EY1YatMB+v/690Lj
Tn5vR+jNUPdlyLzUaNdzBF4/Rh+Ed3bd16b/Oiy2tmPjFmgZS8YpG2IeRyb9zTFSa4PG6iDvQ56A
ooULRO6aXN95/lelfhoF/5xAJ2dLQuYoESekaYjVivsoPxuSQCl7mJwRn8+zO6RxND8z/ZmgKjo/
6cgtggS9enOXVpuHmdAvNz1+vTXOm9+JpvAw9qyeoQ8iILxHyGeyxLgFknWQDU/UZmCMofy90uzS
EAHCBwb+Z4BWxqeSgb6LWck7zjhZRpeYllHO6/HpT46Arq8p3odk28Jf60N/SO/6WQ+zgPmMVPii
gj5ts7ULBbK3hdGMjZp4tKEuCXACIoMQK7cftBDaqwJejZ5XRwZ4rux8H75pPIiYLW7JUmkrjkq0
oq/FSBsAWehx88ezkGyqhzrpKWe1Raj+wtU+oZc5Vx9eNaLixhg3l9N7xtMCK0kzUzEXm/i8kDOS
2+DWXcColHsChD6BCQDMQsJLrnLCRB+86/FiKVzHTh2CakadDZ3IGjdFEtQQynCvyXTH3xCjOAjc
xSGAZliGZdrK3nIpYDY/30fH0qvkCiKBPovzd6r18a0BJdJ0Zp+zLdH2j4kb7PddTyX41iQ1lVyI
oCo1BSe0fWUj6xWATzwy3Y+FmIvYeEY8Gqukh3OM8wOME4HrAnZyrDFq4Rc7YK/QEfmXTd4U/WHg
tgc/AQ1U6F3np4SqFnbWtcgBbf7oUQHJ2kXaZlSPVw1nLirL0htFVW6NDFg+GuyY4+8+4EZFwo59
7GkWybDVYFcYP2gYhh7mwi5u70EX1OEY5jTi1XwZp6GG1Vx0glxNGvHOBtmkkWyn6dHwBdqCI3Gz
Rzmeyl90zq0X2ziyNDlChG1vG7RVKVnI3fxBCEhFywEyIlhdbeWQ0pvIFiYt3qxwDXArPsZ1EVvL
2jz4+ERg3j3NSu+a5aPasM6pSaCQoFgiXAhyjXYP0RK6H7vjm5mNASGoG41VsRzguekoHUCL1KWQ
5Ngx3relB67vIKbmtNt/G21IUKbb0/8UfjDyQTaRCbRw5UXz3u2ni58g/ciGPOFK9z9L7/gOXWxS
gVoOyhuApOUBqc/w3e5H3gzf0ZOYwVudZPxcrRW1CSlAIm+SJgQMFU1R94eEZDf7y7NM5aklEqmZ
R0xt7vEyakwf4upTaT24eLfRWT39J8m3gcpdfvw3U9Z/HFYz6uK0y9vyayvUGzdOBM5fsvfU6e4P
tk2HqmYoaMEJUQhlROUOjmdpilxRcj3R82VINa9lFtloTBg/hT9caX4yReRyvozNOVcTez6XE0aI
ZqyOBd0nmNxLot4gtIz9pb4G6667eGW4asq30w5oBYrM52/U/Z2pU3VrL4o6aVrI0N5smRIZMIuA
CVvlAJZkokruSR054dBGU6l+ooH3wP5Xhzbdj5hpFr/9+NF3ikp344CrXwniNH0p4i4Jtr1KzAI9
7RQklABBjNrct2AGniDM6V1ZkDRg7tRa8+3TxIqZ7ZH0Nu21oU3KE0KmfbZ0LBY/QKtpFdSLhVfj
DBLyiUNZtOewjxxbPUg3FJJOhCFLvbOPCebVN4XwCdCYl8RuCmMsnXSEZaNa4srlxdAYEA1Owgnn
8KqvxCYb9Pgrk/tjvV5x4FvWpfPS+DN2gjcfQFJY4RrjH/mrTR6D8gHC+23aSTc9BTMZdS1fnelS
WNyIV3fNAeh3o64futgXVs6FgLhTrEWCRGM9f2wW/zpQ5+Bjh7WWErCc5mtWpDkBzEXzs8GxyaCl
mpGh1Bg03qTHDMR53duTDFeFKAnlULw8/qo8HqBuL/A3bo+Yn5lh98U9jkl73YFbgAJqrAh8eRm5
XJLQMwY9/RZVUI8X32FYINpMnPC3/3dDaCRX4t95PHIlnJXO3bHK2IArfb1b9XE8wHs7lK2QykI5
An7vdx0hBuWZ4gj6mxpAUF+SWfF+1l0rG8yFIn2b18mnNTHDN3qJrZQuUgjD/j3tgmbMaCuMwQmc
FfoXW1NvpCvQZx2iVU7bFr00H5toc2VmS4BXfRzQvTR4Y0e38bTEJbeZECZoN10sF0Zo6WqafL/x
Zw2l3EMZPzntLJ2XpXWLStHcgoRAYTWv4jIJJ2cv+bP10O6Lr9aHFtoIMXRfRtG5N2wHvSk6K2CF
OAufEZcWZ7TgcCczkPBi4OoiORWsre3Ixyzdi430Z3+ZlQUfvW3LKW4lsRqvW8GAa0lIIGNALSpB
lFGD+oGYAQ1OIL8Xc9L3RsSOj5CpjbD5XqBFzguFB7GvBEB8tLioxlk9+wdNpPAAQxWH8+VWaQE3
Fl6xMdh0nscuHDY7ie57hpa8HZv0WpGW/H3r3S9lAIwRuUY9PydJZKadqtstwd0rFmgZz1wr3G8n
s89374maZQ/0dOIvm5zWrzKBMlQ8sjtpj9e2qEHeZ2zGXh+maoCOp/vgyoH9U4ieICURPLIm+l6k
y7qHiDcFZGGDB1CRyFglRL2GFsFYhPdHJI2Cm2Yf2pTmvFPO2ljJPp/hxLFEP7zFtw+MuHHUuMdn
nBbGmZxemVCgBtSMj8qQz9R96COjOamuT83iw0Awj+91nzJ2VbGjOD6zztumpJFcu4ltPJtXv2Vi
2tQnDzvXV6EanJ2f1OIfYORMoXNxgGTpfQ4NmuikJ952AaZpfDhO3rX10fr7TPL08IG4FLcVQU9o
JmUmbOihxKP3qBaoblUiTXex9oipzscalLjDTpUGWf62l6TDQ3oSVXLnZk8xZqJIiFw7Kya0ariG
dRK4bGbpT5ygUK77kyJi77n6Gz5Pafg6wEapwnoc61o0REFVGk8nXXz7Ka0/cEcWF70ZzPINInqK
vPyNrVMY4QR4ylbEDyeJuViGBJAkrZ95qvFcqOwrmLb5Qi3+B0AoulPOyzEaOD55kjs/WYESjVx4
9V4K6uRSQwsfr2w4PyvW84VSDTEy9t3oSJInlkPaWzkn4jzz6Lr6DAJkj1VpgOwsyoZHoJq8xFU8
VHFtW7qtATCqEk8VMWKj+pz66rXBAZGUZP8Yl7dkwfGXtunQqPvPSKn/dCHiMjkq1CC8POIsOXH5
yANKoCyPRdgjaZKTS3acpDdBhoCZ08/Vrg09a1OC9Bo456WLhko9D5u3JJ7ZmCWj/c5fE+29vWm2
yi3gAxySpDsOfsTzGLLCKLu9Oo45WAZN7T88+DsdNjZy6YGIepUiZUVGJ3lM4MRpF4+o/zzFOLNb
fNEB2yHDCYTlcpvj10iU7pLEQEI/lCyr2VZrQRwxHyYZKZ2Kir15gIhHp4DI2dHwSvrc7jYOapuK
MCwn0VRAWnry0BI057+F9ti35OGeM3+RI4EkD+QCWwEIzyyzGwPq/nGA+x4HnhYnt1JdWuZsI7Sz
OamIM45ARUQ14PYaiFY4A6FjUWuLvH+X2AOSmuLbgtal44PowgaeA1j5uVwrlZjz+4LpISNH8lVC
3Y8I1G8favgCCNHYsWPK4YN/7FlfkM9KSwKY9ggW/zxxtSzMVSUUuhyIjT1HYFHPbh5Tm5GC2Yh3
By8D06Iq76kfUN774tzWUCdyRvad2iaQ7Zcn/LuN31QTWudJppny2FcwbUXbAszlUl7zUKhVtq5y
Zs+TQ9l7enLZhz86yRTKcGd3An8bgisAyMry1eJd6xdUaj3//1tblOch4OhkseYfocUulex8w1mJ
17xpYsP8lDs7168Wy0nduzdtCMvFTmdbOhxQj4Dsv1oJCVShetp0A1BzGsEvPHZQDm6N7x4Fk62+
5A1YoRfEpfK5jHNGqm4Y+DHfuIBsIf93u2uTLF6BFbU77hUvx5JVSjdVBDuLcwrTBL2arGT9eE73
6IoHH35MeroIxzQpUL/1cMxW/SU3ihN+qXIwEccOvTrd1V3QallPNdZyG4ADbMBlYIfRLCiOK/IB
NlF77tNhk+yGzOnynE9t3/fVcG3Wn/HcnXp+izYbd3r9TWYWCAY1VapPLad0aihf3OIC+q9Jnln+
Dt4opbJWobRUP7THVRWduGfG87gDCW2AakvxgbkAkiKF8OTRHiv6iHjDvtKs3wDlIDNKuUzE8g4D
nAKagMP7n2IJCzqheFyNMT77mlGmXyyp9rrdq4gzdhqP5XM+1KwEKFGM64tbtuGxV9ZmwBQ6HYxI
cpr0j+USvwXoA1D8B7H9CT4FED+gV4Ji5RuzmQY4OiBorRKoLuOqebG38DP/d1t0NCdemU88QbO6
cvoeBa48pEn6uQMhr71gF7bzmP0MpMTAOQt6Y1uxxDpVkxZvtvpBMRWwjYXPNun12gMldEqONqeK
fFQO59UXHo3sT1Oc2GtfRtk6BWpwZcGeAT/8qbCH4U6Po2ktA2uyTpdMgP0o9LNAg/gd5GwA/aBl
CVwH+/adWZCfpVIwuDOa59t5j1DbOWH0GmwROcLnbSgTNGNr0nUz3f44pQGBQtctA2Xp5flrmidd
NTBMpeZon/LVSiXfEQhxnmBGjRLKl9qtGTXgJk4+pDXovxSMsOPYCcYAO4FoVISPxvUVYcjxPJ38
biv1VNarpZv3RBre+x13wHtl9/Ikorf/39og1Puy18T2MLe2dH1NvXSLqf5TUSFmP9EZkuE3pfvO
7fADRw6xah6fkrz5vfSSDvTcszzJ8N04PBYVFExxbqz90BWnRS7w4jYQzGsIERuzUrVLbT2/kO6b
47kf1s36ne4LHXpoQOF3sSsD5XI3yKKhANzCGN3WRC5S2Laic3SR9ChTwHXKtfAspE9FZBnnuXrq
QcRHjDpo8+6RwjztIS7LtdYqVCGHABS6n6GOa6uEWpLqiw1gG4DSYHdxsxi46n0Y5sCYfTRMBdz0
BO9ZvwQKWtSp5tqMZm04wGq7xP6dzQUEzrS6tb6wXWB6rDSBrOB9FkRRpwWK137ZKkMN2uwTHkn5
hCEt6r0v2f1QeH+mTyaT1XhN4oN/kyD3HUqOm2MJVHbo5eDpglxAHnGkPWonW7Xt9sZDVsbDIs/J
Q1RpXSAInPbz6r214weIKOx+Xsrlf4yaKVQenJQznevM4dP4SN9L0K4+G12J9nja2Wa1/Ur3Nm8b
qBj1TYGp9F4EnzNx3GlUCZ1hBf08/pn4Y1OSUPOf1zpFa98iSg0XE69Hez4zN6DtHZMooOV18T97
Fm+DF2oAB5ZMiZV8VM8VIeAaF06Vj3bZE2vRiALOcwHRwWypex35y15K4X5HP5KNxEfV/U7lbBvb
ewL5Mmpk3OAip3xgt8XZ3HeMndljazakX/6OGB8ct0qjFZ70IFTr6bNzCIk6mi19KVsvTkQeVEZC
j9wU1OKRkTFD5j6nAy8+Fbi+icidRvwJfCFGC7ohRNGYodTDXsK2wRmCf7yXWe9Y/yxYvoZvu5VD
apeJfFLxvrBmFpICog0f6NGoYcdrk4WlKSzoIjFrdEelCl9PL6ogVeMe+seHAt8y1a/BznLlwjla
R7TN6a5rPAMMeKhmjuNlxj0RAvnBlVmxlhV3foNUhtiNcSGHDUxzl+ZWmUSzidYlGH2SwF9ZcyoO
jpeC7z3g9Nos5M+rbTM2xbi9MrsmO/BFPXZOODq5VG+JvfNJgrvT3RduzNdz1ipY9ID62uOqbwBU
yZqNcEZVWTUH0UWBEKu8/TjltPlPamJqNEjqjRtqrKiPS+Dd6bmtNfKMHykEefxOcKzo2ivNl9cy
4BmQukZ1WXSQq1MToPppc8+rVvB19n6paE2tdx/BygE2aHkhACZpfqVGR1izqTQFqxwHWH6XYOMt
pyJfvZWQExNMxF5voxLEWWdnMG54mtAR/iORgP4vE8ifcWFiaeCFiIIryy2I8UCYqils/4YliVKS
puPawp+l2mdK2hngJGgIkoLTy+QJVNuOOq/WeDELDRtARQ3nIkUDj63S5Qn38NpbJGTA7zuHkHqC
0+fZLeeeFTdouJmVGCHqKpBX+A8Iq+IJztWvGo54j4HlAIkputTUk0EqP3P0XxOI18ZN3lyxhNPp
LPhdpHp4iiEuFSPP8qbVM6g4sdG4p/GGJ8Zzv2FE/kp3/lwb7p2c61cY9Z/9x6XRQpj67749/Ie7
5hGFztORA8ctYF8eGwJzHzdh5Fc5DUzSonlUIh393pqAlXW2N0XDis+HrHWqkgpC/54tLna1RVsN
JOkmuSwMw9TnJbIXkZYz/TNMdSV4WQU1uWq7SBrqMpqsWZCyaiwoSHeU8nsAzYuS2lPjpq3pSzBj
dGBv1dIAe+k0NyoSGtm3NLc4x3/ZWFUHDw/2o+XqsNPUA+3wlPvHGM//8cOYydonzyLfql1xGRRZ
fsYllfWaxKjEuVWq9Moyq8D4zP9xuS8Wu0bvcE6hEDz4ZIRcu+wO29GnXj6o/z+/6ook2U8+pvDf
dqvulQbXL6BI+5Mf7P2CqRqyaNhI0fmKyW0n0bjye3iYYNyUJ3CtQMRCbgoevWSeZIXdLbkXNkF9
7lp50qtG1A5aiQ5MeEzrfptjmFMvEx2Unpxzfgwu9+uUO1hXhXUKAT/48brhZ0KO9L8SPlI0QnTo
iZXnaQYztWchsLqED9ZDq1oHrCExaQooAiKO2kQ9jc4r+0o+m1XVlPXpNUBotKkMSofBmm5TrJ5t
fGKT2ukqdAUPcJl2Lp00Wmx9YLfe8Nvb+LXtUjxDLfKUcDr0212negJNHiSZqEY1citW7cSpzpND
0W9Bp8X45amaM0WmwElUgv/Gs93p2TdUH3HuLqAxpraxzUEr2PiVGXlfkqQlGTZC7vxzr+M9Gn6b
1YLAYUCyHtXx+eLEO6Ylbo/29JzpoveG2yW4r0WBPPlMrOSJM1uUEzKvPeSGOWvFtheWCNrRmgHI
vpFwOyUEoqyhxOokplWXueol2z2kMZN96Uj9HqGJzc6/XJchws9CXiIaavwa7c7yJiy+ujDKVZ1R
MBMvYFmTQEzrXjH2JBDsEJo6d5Tt035Zs5S0otit1Jbav2WKUNMxU+8KSHIGsM/oMSW5XlY6z+pc
IlRC793qLcCNriO+q8DHCPBNr/FOVW5fjbSi632DCODdnAtiB0EK6+E2f1NOjtnxVVE0Jy5I1Mlm
RQiFg4osjFUF8Bxs23nOtDQ+dqnrNSIzZF/p/T5ifCLaKt72X9l+m+rlaFxvQjmAIyv6TmB1guRL
1k+FA9BJcbCXUbf+7eKSCdGOOJuOpkOgPsqxF6/fj1QMPOH8ftoEyGeUh6y+Y3+/4MzBBQSpK3vF
F4Paz4PCBaOJV6Pz+JH6qStnOMb3c4ZB/F7RNMk/okFF4RPR6reka6G24urtdT1EaWPhSU1+pGNP
z14KdEtzwh0KFJuEeIZAZIl9NSRDspBM1EpeeFX+HJxjzWQNazH2dZS1l+6mTkdYdb+2qk3RWupy
EBJFPYAkGUCHHIaGZhv7cS5x3ixwd1rfGPP78AkhJkcxjDRpVkQD1Pk7ggqmzmisk9N3pWrKwXGA
cFUsPRJvfnbHSNJFhG9HbbhMwB5NPC2/4ug49gQ8339nguOe43MIpXK9Pr0S2xQqtiUciGHGfKLD
8UgrsuXa2P/zfQi841h2xE8kku34kgpEmZLblFmvhmDl4jotax9gPOPWEcrU+PE3xJt7S8qCj4aM
eUeKGicD39HITfVaLOzV0UdkgCpBug50LS41DB3I8BNEIKlCxRCU1KYFQ3XANttw4Bqo6wl62bqw
FwJj/9KaZeXgxitYhryuvdneTVpfLvWIIA7QHFzvFQVY4C4vawUYBYL9pttgmP6+7nbJGHO2rUAt
ZcvzRvZatJZ137CPdrnsiaFb7p5NM/2FkMCqQKsdPvLkK5hMKdOU4SjSomfNDhIBMhkDaJSl+l7t
J6Kvkr6tQsE4whO2GSB2Y8B5m23kTJn8M6msbAlUfysf3gYLZPqkYSFsBy9obb07HxHj4opquLYZ
TwMVR0fO3kMf0dYJz/qj5dIFFSH3ph32fOk4hEqjlx6SvCCc5T57tMYAhCDLqQ0/DaZ3kGw+iu+i
1GBxf7lJkEDA5KKq9q6YOp8KNNs6jMmn02E+4hlJvEe/vpxuFufDWHkU3cm+i3jezjE4m85nxq2x
Oapu9LO1/5w6toneF7SWv04KiY5cehHBGUOuNI02HQnPPh06ZVdAlzuV0NyhU4WT5BdUgBaXLB0B
WENmFGtPeWZixeHCkG5qRZ/JrFalSvYWHgCuJJ1TMC7U6E3dYYG34qXoVwyxsHPduvIrYNqBWmmX
U3MpMIrLuJyxvN/LZkgOVlORMuawB98nwdYIMSn92f4+Opks/lkTlZw0XYMxUY0dQQrQQLAo64GF
UzORxxWEDHg0nIRaYFzBlDyv0UAV/qU8QAKd1CoRGmEqG8qMVkh2lRNWBFjXf5lPdDlKRmPVWaqs
kk3CvDOFKf6ZisPFtKJOtAY211d4P4jEuFpLTiQCe13AxnYJs2oSMZcOEL+ne47NhNNhMG2FMG3E
dHaFBO4pDv3lKyF1n8hlEGpxolZDgCTEDDfcN/MaMMlvu0vCn0i/karDqfPP2cZU9o6PbqOvJh5Z
OBdQN+a6UpbUegfgD1RKpqW6D8+5EhNoIbhmDrTtKc0d5rRWntsZJqN0HBZmO34/kgibaa4wa7AA
i8Tg6E8Iqp9xmJbHcHBBYHM5mwC0gbe1tZ0ubBffKiQHOvA7eHXeeMNYesKsIU2+hQi/Unp0+0Z+
Mb1pXseJMDyy0miNiV/HXPjgO4s+aTFbEEjZD8qyoKdKFyBTz3Y79zio1LdePFjpo7MU1rt64Ie5
0Hes9wcqtbJ0I80BSHhyYR+J9RspcorGNSzsuw8m8d4ktO+vqdOnxRsQ3eA8ZAcwjxbeBumdbZ9s
AuXTS8qeismb5RMtXEgoel/qB2v1g/JDcp7Vnel0P0mCCegHyAF3oXfihLEeCUH+nuNWdawjvTh+
uN6jyPM4U3KEXkz8iChF18QKiA/FqFpIPc79GzOeuliq6/V8+RUZqhdVPE7UnWYUeoNcMKdE+W9/
QAzF9K1Bxikw+qVgKsx17TzMoFE58OThUICAvNHh1LshfMjWk0sQzOB90SXUUW62iax9MiiqsG15
UYk2MZOyJRhznfHkL9VD9lkcpKlB7objsI8u4BKIr3owrKRqNIP314Mt1EpqG3/SaGTE9QYFKGg5
V9s4svjrljOvQkDLY3cFNbp/StEsdBD5bRbhyf7E7PoTznz04dTUScyx2cWMA9KyEbcHnEuAfkEX
0/f0tzYnzwq9IRWVRJL/q5gPTawPxzFwuaISYWv6Z0Rpdk0U/Kjd2qWM4BAi6dDtQvqyeFA1Zvp9
nVbMLEugW6AyfGkT+eqDoqwdEb9H8N11Pyv4igjCd1IUEGZdQLZfAoIVdR8bXmDehJEO+Sgr7rP3
pKDe4FdtyM6Eo6m54gr5V0zEw4yiglQMzh6ZI97wxof5haJ0wW9FW+fYUFpN2TNslqsqEOLF2xwt
TKGEe6mgwnkEMLj2CcbKCDdcmlnugazldHNNLIIy4NIi46WV0h0r+JxovphdteXW41AyKG6/LCiZ
6PnRDv54rqP8uuE3aI9m4kFTHGmZcAdeHpYrkzcaR7dE53bDV5m5DKrUq1cw4k/WjhKjSn+kgufc
BBJpYQKepd5IuAO5vbcNsn6IvIFztDEqh4/cAqKHR0VktVuFHzDg64lSCYWd/hETFQuNq3MjWeEy
tG4MP9g7kJ9p2e4pPF46tFwN70zf7pQEpRZ29QA6VtjKnTMuefbbQ+oFKnGLn/JqK4mczlqdfzje
+wb8C+vwXc9bwQvHRI4a/EZhTlIJR3xXMlptJscEr+UHb6yEoer75+jb70WVg5UqiuJhcikqfACU
x/ti8OEyA1k8mU+rsVguhQN4KzGdWrckF3IRh2PT8D3NbU3GuUXPABj3WQvCYzcb0ABUT5cddMpJ
oY5FBvK0o+dfDUfk8o7eS0Ki70Cy7OewuCeW62obPSAa7ED1/+iTbdeEZE48cICwBF/a4BB3cR92
1t9Kdk/0DO4kkH5U9vxiOHEvy9YaeojWXaljp3dqFADLYkXkmsNh/F4fQ214FSV2zB1mVFEP5ETZ
NActDPN55u5qwtuyhiIGSZ2E8T7cEnHo3OQxmdMgfRktykAu7mFcCeV5C7JDxd9Wiaw0cMpGQNb+
FpkAZS3fSo/1KCSWQEfsroaPeXYZxBAauGmFCDJr69YYrpbJPWQfq4W9uaUeZryqAGgzQ6a0jbGi
njGSd/1k9SeCqPsNCB+Sz/aCyhpAiyMCfRT0hQ/FdjFj5hNbY2polN5Iwc7L2duk4CUIqhOg8PRk
U45xGndWKt20fmErW95Vm5Poqy94H2hwi7CkpZ33e8MlbZcviZ53HM9AU17BCyAz+bq1TFzR92xs
A5n7sIuMmiJ2Zfevj3G7RZI/XFp+ay9QHIAnIzDaFx+11GvNchIHi6br9uQil43WVWYnDaAqNWoG
BSDLA4icsFXwOL9Rj5PVCY0EdU4yJMLCtwVCM5XhFnMRYvbqnmpNLPqAG92mb26kE+0uImQUln3B
oOmnF23GqkOkW6J3Bza/BC8RrF3P+puKyJjtYHJceTQkO3ACeRAsP5kYuQiH+nLgUizoOfWRAY6F
GjFgfuFkGF6esKu7RextJHDPSSJeGLwGC+1DC8zivZhKzRG83Og8fB+re1K/5vdmVn+IZxnmYh12
f49QA46RjnaDYAR8zGtAWrbv+AiyFQw+gr+reBMevfzvf/gnYzCBCQ3ugsb1Mh/J15K9qpNBP4Zm
4UzsAst3VYbi9gGAx6AjZhW05TAsstRy2+TRJbfl06TuDCkfRj91jE+U21Ix9k6WBWp+fQAXnErL
o3cOYsrk6x4bdT1ZoNDW/Y+oJX5DR6LiUnWhvyM/onqL4u0EsmQOhg6wQEygTUcqikKFY36FLOEf
dujIh9BrgyHF11cMyYIR/GRHNjd3Gs7XVhk0T7j7PF0okH5rYAFf9cfdW+K2Wj5WQdENQ8alehLx
rcNZzDZ6iPf1IkXRs6NsGBmgTDB16ZD1wOSomPRm/n+BlUFExwrhdlh5Zqa/1AQajQld5NDRrkhE
1CTx7FMGfmocme3yWiFX4i57dlG04fSqObWKDwtGAKmdGVAtxkmJ4fthNjRnshxQWxVHxn8kfZK4
Rpqac3xVo0kBqkTeM8PPGUirdlNgA/OLOK+zoN3UPzj0+OfZ3yUOY4lCzXT33gGnpmhLU3nH1MCt
WCGt0aFYLMDe3BGfKOK2K3Wu+fARJozjFvtC1bmwUst2YYiWLozIiRvcczKY77jYtrE4Ouevdoc1
mWwb60ykUsDIILYhh4/jYlLg23CRqUMt3G1IcwRwvyWxuHxsEjz7Tx5irR4Z0w3hm9S9sgppuSLz
opWVksJq37TxVEisLYAlxO6gscp2Sy07cXlSIZIWTMb8G6V62MDoVO4njqjFK0S7BdHGpoEAIBVf
Isu22mQEayUH31Civcr0S/DXIUP8U6eUFOdX2lVP+Pd6GKH/M6WVVQNn1Htp7CvqOYrcCMZQANIH
AvZLlaSQrXJ18cCaJ8aLh+ZjyYxnIhxcL0Mc6y43rSjWiBleT0jUYpF/81sZ6Y0sL5ujxNfCc4Oo
/R+RMfJqHzZIv3g4Jfn02weFzaUlan1v6+Bsf4ySipJIyrKhbKvxN+PKpHwK6+G1r47d6WXfM0w0
XT94VnbVT6LKaCWHR+A+HIPFsbjCcOV0kWYMaPXx+d19GJHFXc0v9ggQCTfT7T21KAY05NzJ6sgt
88bpT1aqXQzvXZBj87+b9ysKVuvOAV/CUQaaCYr0Srrd7Era+OrzJNnN+13aAhONhhjPPRQ7Ai/d
Rltfi3cWXufsMOuYMqaWLUGnjN1s2bzQ/yk3I38nuRXpV30t3T4FpFAyibqXAyxosHJ2HsiO0s1s
EnotuqzSUkVTiUNl95VILvB0X9/QOnl37u9W5qvjsJ5xdLoemOABKjeoayPZweBUscLwb4n8HOz+
WKYwBnc1TZh+vPbflRt/6fUGKMS0/UtgmuF+9oRLawfsCddQ1XsPFsavS40A9y0gRBYrAAQVU+UK
RvA9unCdydpgmoDSzt7THsdQ2XCY2CGMa2J+H+jKzAxpc/fG/mFT/Q1J9ZVI+tJUk3JfStCm0bVF
qZqUHoPu/27RTqlKAMGQmhsIEVHo2EHFyB5YUaZdIU3n1bvHaOcsGmkJaFUB94gnJrk6+a/XitAb
2VgDDX/i/6yvJkIPKpKRkYedy5GkzRVsgCTspVAZ1imAwvPM+7iKj8oSvAMjic98rlC6AU/FZWr2
bzAG7FMRdNlp6AGrujQC8dY46sX4ZKabBgZTuvEt/a2MLBo/DEaWgY1S0t19WC5dZsMmBbvl/xUC
izjeJkJMnV2BGlYa+yQvjoiq9rD9ZKLR3j2kk2tXNv0odKO//5wr6ZFt8HGWNNykQiUSj60zilxU
eKRp+gCGU1BwtWuLjb2xYwVvC9C+QmOk0kbyLpzpiCKiwzRczLhOcvBruh6dGo3B0Y9n9+CN9vgE
AlHmb/2fDD0csBIH4zAGdKqsfR/0eAhcd4JQGaV5l3QBy3Vt30ka2/Hp1WEx11miUZHlLk1NaHYR
l7CU5943A1X+QiJ59xfBRcdNSlVgMnniAbTwgSpOM4RILmLq9LJrAvpTAcFq4WA40HFxvJu9It3J
jgc4rd2P+pfTjiOdyiWd3U/9K6EJ7Am/Buk7+vQjgSwFcYjP8sc5TJbZdnVaH9i2gVBZi36WvUQz
ZvbVQkI9xshfeULGZiCCieJOPvDWGo5DMbatCMSIMpFXvLeOVlDvlhlgw6e076xHW/WLtH2wess9
9thzbhhq0E27JGtZajpoeXFw7EU84GMysLnfE2HHel3zOxS6CFXDd1hgRG3OxpK/SHLNqGmXmZOZ
HOp928fIO2s70tvoWgYxdFmqEwMvNMfJAX9TJrIVoX6kBDlXk11xUdQdH1wa+kCQgpXQgpW3/x/o
R9WBbqzIdqSH66Pyth2aC2ly+6DZl0GtG32ZGleVB9ptY+Mt0eEcC/Og+/pY3y1Iggj4sjC9xleU
HEe2qfWJ73fpGd4jLzdR6RqOKjUxdasiWc79kGil/+XFib6rygnIfRzLvJSLmjzje9IIQnoBMlho
T+oIPlz6b44h42+Krg6bjc4R7i5Ez2Wlv7d9D8lj8na3U08TuFi8w1nuH6MY82+KLz8BHLGDxuJj
3FjRmYd8GPVyc/H34SPeL8bM6aeDMHeKFn0hxbJLgVRTsow7dY5kJ/C2o2SCB9T8NeBqzcOL8CsF
6XEZLc4fAjnG3UvVcIIAZAZ/ACXIADeqMr9p/C0s/cQsU2q9myH8eSjQheLs0ibFLX3Ju/VQ/vBz
gjrc0bJttNB0/q2b1WaX6NY6ayk7046bNjMn2S7A55+Xl/B1I8nrRpYv7XPys6eyij7qUa85C1xw
gDm4igEh5EyhEPhxMgBz63HVrAjVPr4n99SLn6ywMAu635qyGqMDQUYmTqufrqJqbRusVY3+8gEl
yeg9IPSkHepNN5MPEKoS6rsWbMZcLI+CyEZ0ahBTgFEqUnOdBmL2MUECJA2wHeRPVvV7LS2T0iWX
G5C2SXMoveLZPFKYunU9iHkcbM60i7Dz50o8dYNGX5mc2xr2ISm1DAjaB4dr+nNz35jMea2516nc
OSJMl8Jt6kKj7dZFy6fR+ASMHjMSh9Sf5GajE/2OTvSlBZdSPyybN2HQEPJb/HeSERIG/9zVjBSa
KUXxNz7t/D6MrKRoT/T57OAFcDwQyVjptNGcF+wOoBb1jNZirrvE2des++RwymnoxVY8T818sGrh
rh2bysgIzRHHTaUjgmXTVQuPX3mVSjqZsonsBBqpEO9W/N5OBqG+Uvw5K+mTXLvlLbCgvjPfKIWv
xNGCXu1FIaSrT7sMPMnjQ2PxwTw1+owuiGcKjwvXHP8HHLzyF92Ep2G/iAZ+Ey1bFZ//P2hYhzJn
0gOMWYtnQwK7garcHDd03d3TqLCxgQS0Z9hTJK2NeTZGIOwgCtM7HSz66VJEa7TKCBTCXwk+cXt9
+GVSEJxaZBWzLUKG9S+80d2CUep1BIyTuPMB42oz1eppYggY9iZTbLYDEo2cThyXoOW5t5ethPEV
odlHJWLclJHSqkWirYrdoISrzXBLCweieKZUog4c7/TWIcsJlEQUAIU7tBP1TlPzBLfL2f88T1H+
9c4uUSbAujHEaYGxlI1gfu7xStdJHelHKldQB8FsvoJmTnOpylK+bxEE816Cr5VNXMCwbLf8PfQw
teD9r/CHQ6/prUNrhW69epNrJu0fIV0WHKwbi+GimAIYzn+zZtHOglXmAoia3FRt5WbsOAFPjAAM
QDw/urvOaDKe5g8OsAmOWlqDpl7uJtYvV+mRaPbvEGSR2fAvDHUoe/m2dA5ehWT55xkBTTO7qdt0
OQzWnotwiHXhsDC4Q/EI3iZK7/laDnNTg1cq/5DwVRkxSEj//HsFYO6dtWp6hYhymM3NcM0S6p+G
SFFPwTyWm/O4FmOHDhLSzW1RMpYf4Z4O8NVPpiLd5s2SkYIgP9av1T5NzAOFa09LB2OKtvGYrmru
tNwh1DLXx8VTJIzYFjHrP6LTTVWvkAl1APMnyxZ+U5r3+MyY7MH1miwWmEgm04ckGh4lbpjiW3NR
PPdV/RF/3zaNUPDOzyVie0ISrkijiojlo22nKIKecxAqtddZ3Nilfp6jHSlo8i3OgEoOXvHPJ2hV
rcWNINeUrHOomE5oE9vVKbWRWH5sOhLQmH7MTbKjNvs6fGigQNtkvMihvv/1Zo1LPpJcLSCxyO++
wOU0XsOgZOPjk7sKG4iAN6kU9/7MjiC2WCjB93cgF/bLAcBaVTr1XuovEbvRSi8pWU5RhMHn6tFU
PIaZ738JTnr0e9YMdpgSRayzXY85uYR72TW35xlDd0g6w0Nbs3gweKof/oCLWLkmoO1Pfj0bbLpV
LtRJpKKbVa9VoKIj7OmkS8L3Z7akrk8m1kViQUiXwzjSRoL9se2libfvAmIeVsN9es6yGGDvIgX+
+sPsjvUPd6XyM+v/Me2XsSZdQ1iUqe+/Y1/n9eFkJTYXoFWEbECP8eAE7w+Mli3lQ+9lU6PEx1sj
Stt3Q7/hUpIxHYRuUYITJrX8BBwXWx9dluJoISbwqlIGgI94Ih8m68GE9oYLrITlOB4YiVlwSD7H
/GhaXb+nAO51ZWHKm2Fn3QkUZ+R1hgnBnNBcq7KBtcEY+1pcYaiPXaWtWbBfbUr97aV8xhXNu8yW
NaIddwoBuOKofuYpPY2ZvLlUL0C+wQJHoPOpSx5H/+DKRcKBZ+1zbOJX3LcrTrLvm8a6kb48A2yO
29dDtUNyHTSlfsKkUJbmMI66BqqWJO24HggEPlGhbvPu7zmyB+Vu8AOmJWe4JVFgNqJXnlDKpMJQ
2zcNWslZ2xv/T3l7Rka5xT7jt7G+qcpTJ9DXwbjVchMjuTk6OWXp6FJt6TeFdDbRvYfkLXM4odw+
58eIYpgojJZhLP52gE6B9Pr++b+wXbyHuAJBDso3sDseZlBQHLS6daRZTI2SjyZ2qAog6uQbL1gW
evj/Z8o565m1dgrd+2FO7YWDxqYse+VRJMBOluVVp3T+YCrkFupSqYuEV7ualgElS5IyCCt92L26
C8aDnTlRUAGu9eQp6vDWfkkZOC3002rPBc5G/pyjAdi53yOBfJwPS9ACGksDcejnAtJ1ixQsmjd2
ZDDlqFIGa2AJ5O2j4MmOtTrG68mGzuVKaXfkhn2n+oBJuWp+vQAhzQjYZxkqL1QVs/tmFNyuyT9R
F8BDMFYPnGHWzuA8/lcAlE6drMVIV61RIktNDR2ksLnY93U0CJfEGx2CMbM75FmuwPkMYkJpr0+k
ANdWPpBOv4DzLXbYVMy+Tdpk/KLLv5XU6LRpIflxifn8K1BXs8p5eyqZY46bM9A6aiCth5+ELFnY
QR85jtjB5d7u2Se3tSxAj/8/ffvMC1YwqGHOE9YiSZTGZDXVqJixaahhVuvd11tGyNnAf5a5NTbV
UrEPZbsaQmlpk+wq7+b2xTNAlzzBfpdzQaw5o+L2m7/1jnF2pg5hXna4dzNlJrn/FNxWbQ9sr1Xd
kRuD3fJmgYwENvAwXIUOurIag0WdwqfZjI9zZLfFHq5v7aEVok/TAdKLq1z6Y+xa3TwksXw5cUuu
A7W2InK2RtJDxQN03NDkxCEm2tF+NOjpCDBgrzDUoabgjE+Z408upww6oljQb/hwMi8S5qKKl8we
yTPhe5vzzun0eXUsHmwn6rmRMVRpt3u8c4yVPiKmjxQZRRWfFdbNu+j6KwENPzl/wpOd/rxd1rLd
h02Lr+4FpYrO4Iy+GNcfgpRaxTZZkdVtpvB3U0IWzgxx/cQ5keowgoYmVb5LbEAhFvyxKHiVMZs/
MXLOPTVk49/3/6CPXHgOmZMGcpd7vpaeJhWk0nee37+IyzgJWbojRDZ9k93piQxhe1s8kFLMALdQ
BEWHfe0LqG8jn+ojIoWhfLTfat0ALQROYZKEfpaANddzFyK6hn1iuTOabw6KSpV5HjE65Dsy/CmG
pcjUjD/V0e3K9biP4msWKY3JOCcGgwI9OzLIAfgXyPUjHKfAOm4TXyc+SjJAj9VPSGrUrRtziQE2
D0ss/YxXlfjfMjqwfa0lA1grl4BdMrbVwuadh7VhqCcSEfP1MbwYaZGznDYvwKpGLKPPWyttreEq
u5Y/OgYBGmdL7JYqPrr1KzJlAGN07cklZTzu6e+zRfDLcvtIgpo7ZkSk9/l7tBLNgysk/oAAyVqX
ozqhvXrDyJ2UgLn5A3/ErJCitRlytyCeWNUC18K7ShD65trtSlSDX01eNVi6nZiDTJcNkubwcJrI
eRMFivtfKg73gaZkMaeyxdr84R/uwJ7no4gOOcPQwmdu2GijmahZT4XF+doKxM9EHSlC9uPemaRo
Me8pLERDwO5f/Bxr657iQfGb4hi4bB7GpEaIAzWe5gKbO+3blcVh/4v7rwBtMVWuBj/ZBpQuthD/
Xwu0FGnPzVE6esYKbA43vsXodeV2d+Wf4MBqvPGBoAZUHnMtzZeXYyPEFPoGWuFCBMqQLZOaxXYO
IJWLlVFChfcfu3T/0izcPDFH+l9r+6LecClga716zhgoFEynpSF91fFmwK++hyXF0DD7njWVcy7m
kUenbnqHat9/n0wSk9NBS1UBtjK2Txcnyp3TGo/At8t5j2SskR10pjy48JHLulNtI9gobimAYLxT
FO9lSihF25OQvM+vhyPGO++RP1vX3khWJc2G2r/BmKjoRjImg4iCZNXE78q7WgzSbxVHa+22Iv9w
rZN9TnU2rJhujbfoJtci9k/G9Apx6ECsl0vwaYgY/uQ3TvVGdo8lYbXjSPfeB+jLI1cGl6Xy9YTW
jbJFbH88HzxY/bk2OtqHH3Ap0W5/pasJeeDHUzA8LjSnFjk+somVS9PBygsmNvjEcBktbzMCS+0c
WItNipqZ9/BKAY3isIL+2dz/yKuaojSFw4SlKWCewpFyNDnj6aQN8pA/IDDIIUmWmtANi4s4hHSM
ehYXoh/qLcw1TITYZNHZdfbmdiHVPBSil6rnQqtgcLGd+Rgk6V5UKA5tc/KLOQo8QxKUVtb9BlYN
FcShrj8Q5OxqeeGCjPNe94MjEBRz5IusaYmxbI/9L1dttbzbPM6WJWJ4nZG9pb45sQZ0ei0zi/be
C3M/DuA+AFpNi3IpXVOzWiQoUxinbkMT0mvm88ix0bPDRRI+8ZZpKR2h/pwpK3UQT64MR/Q+lidQ
A6Oghj5wnaLg20Me6EDdJy5FYIxtkIwLye7lVUmGlDSH9Bh2EXNpZp8eyThu/Ssn+Uqw0MYWKR8H
nusOIWRHlZmQ7008BNzTsxw9jHQeVAiAe9Jxrk90YJTa+IgvXxHDTY50nUFBeUdqw9I8uebM0jVg
Cj7P3mjvbPMS3otJGhtXcH2VP2LDKrtBseK9ph+SbybOExfnT9nX61n927A1DxJN1P+bAlkNfJk5
FOI7NyWIPayiVnoEMnvdf7S5vCspoQMmVc6ZAOMcnQHe4y8K93/k7t6o+Lyi6Uco1Qg1em3titjR
VJ5d1zCe3+T4C6IlwUa4gCmnTL6HGJLa7pAJTUiud3iv49A1Lk6KaA0C+0RJXHTOHvGp8F42sU2y
eQCKlrtExIiSKQojxQP2Ejri39IqlwEgBGVi7+hFYSwyVn0ADYy5foHoUVjzJoIWIQsVz3x29alK
3Qm9NDjD0Fk0G4mb5GOraa0ZXfKadm2mGUt5/qmlFzk7j7k5Gkqw/378KU03wnq50xQ/NCzC54EC
m6nxw5S/kuXhfXPJhP+QpBb7aUxmq+pITyyd2s3zWX1gtabiBcaWgHClLnbE2Jg0blYdZwwFanUQ
nljCQyrDRVNJM3eUy9zcjTNVGf7z25mYfOmcE624fIFvE0FmSEEML5q21GfoABCV/uzBUG9lZlun
SW+m50v9mT3X4onqlnSfYdMwco2GE5yKSYnJN9fbRfpxaIPtfLaXS6CGaRYMaGDyg+iG+ubRcBcN
zNuMjIYuf3I7zHu8aNSgLCO3/SYbJfohX0Dq4b/KWXMcI1ZtdNrIURVqlyRieMnlszR++ebSmzru
lZeudGV7cvsxgdEA0xibteaIxQRLDtmGOyqdqXVWWOylG/9F1Vxym+2JRg3eALxNDIXuWkFLYA4l
MrbmgdGofJlxXD/d9rtFwiM4QFsk9JnOEu90/TlJ8L8A8R+G98k8J3DYXXv0OIP3RI4wb2ec4OlT
0YEOmmQ/ezK0wuDEH51e6ywW0yh6zHsOsB67X3p+82nK5CIMVX2cJ6a1Liec1PvMWwa33N1NSDnx
tWibNTCazS88XJqT3NhyE4vfq9dJ4Hv4vb4+xretI7BDFfPLVNW9hjUj+BR7IsGAha+a78kMHxoa
LeYWBzigmQa1I/koHyu8NDYnjkqnpLPxa6724PWKpXKQbln14dtXMlU7nhDhX+DNktOGXZGjpvsn
M8b8A5MRfC6EzqXowAHi36CR+gc1/knUtFZU74q2KDnIFjuwTzFCx6Dxa45cPi4qwPINK76UOgFF
OuPHb0PXvfIfvnFdqtsOXte0dQjh4zTEcFOE8ot0Zmjao94/vkYMkNCNrjJKET12fy/i6KIwiw5q
IqOMPyyo6CnADbWqvMHootxs5b6gK3zzjpIzijYg08cciAdZa7PhjhCZrclM0p8vd1acx1YsILyh
asOp8VLLPG3jLEBy/D9qHKxb7vsv5gWgxScJJCh/gBeBts0T/J52iIDJYVbs0yq4l3g0lgmcRr01
2bpnvn2Y4qQN4gn+Y0opk3U05gY+0urtM38G+CdXVn41TzNFboP7o5Um3BDuNbiWx+rVU9rNPzdE
4SXexcE7NkAF/JLVXaHEyyjFWCUAkksG+Syk4mmun+Q9660bVhbYXOD0WAuXZNAfuy6+XmhrJuAa
aAoU9/gKrsIUt7ZDl0hJqQ8X1XuzpL9qx5WIp8efa15wZ1KnddIsjeN+c7Nzw+zLK13YtDpPcP2Y
XWUdEGeXiNlVRsJ9Yi7A5nyy2g5kYBUD50l9ysQ8yvLq/iNtd56jTqyJVAX38dqcbCPLEfDfo4lM
TsAPHaH+JM982Cq74IoG4zsjd7VH1VSHoW9BrpGQbQ572VSp3whAExoaB1iLSY+1vkmjNJyjh0Ve
JP8mvEt/Ucn5It6UN5MEvodqpZI4MDlF1vzR3UW04N4r7JmDiOlPc/A5pFWzpO7Nd/6JCyqpcbRX
UvTdjMInibGy3zD6ATRkaGDN+2E+kPmeFXfhgGCas6u4icygcZp/5VMOEpy27nhJlvJDOjXzApPp
dMrKrBCzxfTPI/e4oACSqSGFw0Kl8Q/EzYwRwA0mpUwI1i/xP7nXwJwSLzSoQ58ihZ9B4+ErFBvZ
Bo+R2Zh4OtUN67v9PCAt0epXWxvcyznmvr6vsX/KgJ3AgfCa9eOZuTiXDRhswWlTIeVqPqeIi4rY
KT4Nzibp3OB8NhDdkEopBUT9meSuFEsOdAugiiO+L9s24cO2jHtORqV7/faMU4UwFDHMJmVQy+DB
CbAmXZ+ckvylDI8+jjurXHoAxqOJd87oVyeCN998ghfDipjs6a2TWcE9E+NdJnQxsnoZWt1gSzEO
SmZbc/FwRITQkD6iU2Qjvi1HzELBZR8ectD/T1COOFoDV/iEwEmhsMcBLAn8wPzMOXtRX6O2WPFJ
sX7JyibRYV02PD2iHDVUCPiSCJ6l9D6N5ie36TS9wb9ppqInqhLdlWFBU5LhRCXQNc6dxR/frT/b
HbPCzEglnUQY1CaVbCZBPfa2gsSxkI8e11gNNroa1XNJRhlknKL5EhIH/4nvTAo5wlkAHqqpiD2o
vPi3QAF1hQ6QJgVJBt5/+BbWf41n0pC7s9clwd5k5tCyRv3g1dTf4uYl0TonQ7Jz58WiD5YA+N+e
ot8RNS5grGEtnIQtMrsI4+G264aWkzFdWnl29Jt2Bv6laRjCDzHredc+MSnu2RS1nX1JTFmUPJay
1wMUTu0regW8kWRL88MPazrljtvqTgbY6mrdl+NXvPznR9s4ryCCJJD4LRPorQrUCAjRx8NAas+K
eBS8jGvDs9SMQYMudGX9kLQ8eGqDrkSnYv3PVh29Ve512XkRCLYkvsV12RBvse9rMv7y1NL4abR7
JTwxwanP+42ZvGx0+Kiqr/4t+FzoCtycI93DltWA4A1ScrwW/gBx4JZAwXrb844AzSCsBythQs2r
sboVyw6jSPWgohHpk6X43pLUmE6TPmQEbTIcb25wqGY7M3IsompwxPtDv3XT7rTLz35mxvZEJ1ji
R1JIsu3cMQWvyVryKlkdVDnmxhkRbCigWNyCcisPxvaAYCAPCdrv2U0KB9ALIezkW//UgNc7dqng
4c3pPO6EnywA3zU0GxTM9cDF7HrCeDG8WnID3wnnSdLIdanEjYZCGZqDeiumoGeHQ6DbE6LFIDr8
BLJ26OzYgJfvi+InZwB6M5LeVqgNSejHSaD5zv1JTYfG0ZrIuU7z0lUCg+DMh0oMsYHftc3Jqiya
/vu7PHkZMocb3quTl7tCNX0sUmw9IpLDhPUElk9VL3JTf/o8/YeTJkTBV9ezNcS8B83r/GjbqZe0
TW0W3rNpNV4glmxFjFgObiInhCGF8pSrtGpStOgQVEnePPTB32m/frpAKBnk/No06S4f7FiqeWp7
29MaO3GKjYPaXiub+YqY8i6pSvOXdmKG61qNZyw9ICDTUJVDb6iopMXcfzA2VExoJdboMc3pP9AC
bYx3OBGqRSIb4rLwVjT/AL+TWKrgSnRBWHltC4UxhFTnCDTrpeltzUMQQFyvuSMKzJSLZvyH3xi9
ifrgiSkiGN3TbKD+cyEwyJpEH9FvpGSx9iUP9MnGynWjkohrxPHVptO3ZoczMHG+Y1gVaPMXYKN1
JKckIZZxki2yL5m4Cr/RfxZoJx1bAcIXgTrBFu3QkUFh833kzGCwbYfUKT13P/GpRf69PPFRDn36
FPDPoh+hSnP0lUyjMiDd8Ea+XpFQnnbsIKBQflYEAWcCu3CkH0hpnUUzHQSIzbvc5muVQtDx3wTu
YJ9pte0wMa7AKJqKYv1V+XPrN/4BkQ+AUk8CeFGJTry2FxGsUvqhF8VN3dM8uLwekLFlmS/4FPXV
Qs7Vc3qZIDt4H3d39Euf+YkZdpK1SLUrpKOO1GICowvS2mqQ7x9rJm/OQLSXMcioNZDQguzvIBQF
L4dMYUZfpJbSxVxRNcGSfMXT6OK2QfjyIVz93YKr4D5Jn8OlSdF//25VM8B7/7KmNSRRgjpTYfv2
UISj8l8H734KsfgNLZGHGMndyhHajabA5OCMaIVzSwsR+3aZm02dkasZqunQqJ9Qk+dMZO0jI9Qm
CvEE8Gyo1e2CXYfTYYk9jTrvsyfk3F7pGCGUPcyLihpSf4P2svYn9BgbUxR9L5FwptSW81XIs60R
Ep6Xr8DNql+JYWIy84sgVHgmqj/fKnqwZIZ4MtE4IQG77msV3uV8gPHDITLYTtiRNtWSp1H7u5V5
ZYdfF6zCQAsmpHdMMvptuEF0ssMIo9knO9GKFdOCBRpQ91wbw1s2shCNPTf8ce6txAVoEoRyfp+q
Og6sQ4eCvWodoSNlhijOpSogrwUZpKK1pvaeU1h08wA+0v7zaQSqsrTva3+kHPvb76dGEmLaAXyL
15KBXpyJADgbk2mKyT3hPTnynPf0daDQb99LwzKgQ3bHcRpvQRthMA11c3CjaZFwxswvorA7lQMY
ZIXpK2/Wcl/Bso+qzWR6n1VUPFmZ+3jESqj0xxc6iEMCP84pyYVOQbbHOkhNe4JKQ9MVUKZcYj+W
WlQaVfcV9RnrFyCEFf/GzG8Y0pH+cmHUxbb45oaHcF3ThaDVXupAnizPn59jlxYLpTvxhv3uwjmv
UO6iuqKIi+BV5zHekuwpkLD9qtMMSjmrUdh5RahNYVaHQcKai0HHFjMVY+w0Yab4Qy/Gy9q3+JdS
x1SJLN0tgFWU7qpzF2hvjShKGAfusgREGIqUsFW9jSuZX3EqmtiJtFe6TzZAZHRJdkbSkhDL7b1i
60sF8b9n5lwRumTRVsHTfmO4EXkLtv/AuDCTeVi96Wwob03IDh0f9Qscjqk1i2QTKRNmOSseT9O5
ypXjSfaOg8VzTuoEMpHIJuMqvAxQ5FEITXSg8YIYsUg8uRbCpVVaZUWn7Ynl0iHgTHhbEIhEIE2b
a2HIp9V8KC8MHpSliZxQzKhnwjSfHP3l52mt2gMywje4e/uaGXtOSxSz4Jg9Q7gi/4Q28aWWDg4l
4DGp7M373raE/AIwQ0/726kKfBdjCnsaOIDM4ne++QU83E8h7uXdfPIk7V5LA7rr2Fr3jQI/EfR0
ARrazH7GjvprkN6PvE7E894o6wysvgWGXpUkdY3BkTWnBV9q/RsPrlGnmaNDYyG0nf385brXE9tt
3FnVh0xsoOFKUCxq1HQ5ekmo8h09Rj5AsV3ka5vIowLEU/QpbXzXVSzXx9GKZ8BU+qA5/KVPQIcG
xxHz3NuVH/3v2vtTynFliAgI02SNNpt5PFIXlJ2uDBYQ1RSi49Qf+eicDFQ3zgh5OzPtVj3y9qZO
nen12KxDr12v+dEXMeoudQGVK7Zp2ppyCp9lcdhbUMqUDMUH8DO3FAcUCBpAL+4Grfpya+OOGFFa
dcYUDkaMTZJ/Qn/siA+Ytmx/lkNrUs1xZ1hKbRnX/+XQPwkVvyvFdiNg1RFuvdcJF8jHsHPbRo+T
ZEXJly90gsc5X3ZM8J2BSU1k4nEXvWKtKVnnOVnGZ8HfPgPskKl3vUzx9t1oopE47o/auBUKz68x
+Y5KCkzEaLQHyCyWiazUExEf9dzWYZynYunRF33CaYkDvqYGLu2IsMgFXluiSrDSZncmGwI1dj7/
eBqCsVos5vLh5P6gVJ2nUKk3IO14n7XbFIwTgLoC7Y8TKPWF7wZ4+3aT9khn6SZgcPPQ3DjTpwrP
At9GDmdzwtLEK/5bdJS0TLI0lBVQe8NKyrg9mUn5f3rDReWA5YZujXZsi7J3AR4UWNe9OscmJkwo
Nvl3T3dfEWiym6wFfx1wl5wPK8eU4GU7p5jQ0V+PKoTi0iaee+9djjc3YTPUNHdJ5w+i6ZfCQ5v9
yQP10pKzwnCE5QBAfQMq5o5ii02KVmGPTeA4IReNSo1moDDbU52iB+wwl+Jv9TjxQhsiiyQgfQv8
WGCatul2Y/hPnRCcOM71VDfPi9hDZ3eRXBWUUqLwkVsDrRYtqg2zH4YYuDsSCHnAVeme655+XA9x
WX6DNe6ypdTd2QhTVmBneSO70jMwgj0JTE1kRhxmrp3nt2YF9+0RRcul3y6RLzC24wkTfhgUTGNz
47ErH+INt0qPgGw/ktjBpNYV9JC1igTYIzXzVUZQP1tXyakonudlRybKJdTvY+TGDn1+4T832SBK
7R6BB4AAwgPK/yu6E4791dhLd0g7IUKS2xNgUy0SRHV6ELq6oitCaWECNn3yo3h9WU+ozuw4yqjm
d6lTvgyc1wTapycVrFlpc4rkTpxHAkjDf6Kxdm1COA7uNeqBKN51xt4cJ7xgDp+MgcRIvaIdvI3e
VNP+o0D1pk2hCmLRcBlDGgVwPy7kURsr8HiJPesWgB8vQz2TmjDEX8RLBCuUwNh/e0oUy0L72UfP
x5buZBu7kZV9YkHk9O0GJQkL2wgPtU2QzzvFXX5VcOF7/s7WSBgukFlv2rbMDnCkg6BZ+sG0rR5x
qpg12fW0LBJKnJPdyC5jWs84XR53yH5u9wAjS6lNojI0D6iLaX++DMhLI4suIvpOgnllNZ8geGuL
xdEYz+DZf7jYCQe2k2uJFcPZh5JrKlAhjIqLHF1A6UV6zVLcUbtEjhzVBtuhrjtI0pok8DD1SSWB
JTIAMe+DKdLY2G+CgkvQw7mKyaskQS9P2VJOGwYgagoge4AyIjAc+fREnAhWctCtX1TPck19t0by
FDwb8F0PQ/EMAVwZFX98TyEkTSHv964g6+1KYvB8Xysxsip4INMg1k/Kg3SqavYTEZFpW626gtm9
JTcMUMqcun++jVcykbayFzET+madWGl8tey3GqGQJZ+ex19kLJe9c8qXHcOxmLZw1YoIIgkaHN9N
ZRic0vnr8oIApfOd55Axq+tx2wkoYaoNlGI9y1R5JuZpLWM1bAHqlEsssRB0jA6YDlDH93unYpnD
hbAKwjiGXHqCK0K5UvZUZ8OlsCG8jCS0B+WZevViYX6uvfL5tQVAJb2nLgQnAL3+HSNw39VdfwIQ
8yjU/bsIu+kMybXaA5O23OeUz3dljaycAp5ysQtjVzKcvaGe+qm7MrhS/H5F01GJfFMwlXp5RP52
5W2o8VOfAK7fi3OBI/OG/pAyV/7yuz3Qu2mSINfq93IVoGSDQbpINGSISKUL6QteNMAlyBFj1l8j
FFo4V1iysw6m/H9LNBRFNlNdd4oB8vz/Xa8/pPW6YDpbT0QhjEHNHNbHiVOhg0IONokC0ap4z0Wd
EssxRgnoUW7Cxxuot5v6J+i3mK8PwovxZDsBV+YF8MtEntyFS4buV8Uryaef36ttOq70v+6mkcOw
A4HV5TRZJ3f5/D6/eQvXx1BBIxkdrvb4VjEFb6ZolOB8wTuQwWrKEZNzLFAm73T2CJX2tNZymTL1
7e//GZmSDL2vdwkNLeQzCmXZe6OydC0s9SpViWVxBBkhf2ttNFfDc/qfIx2lcL/KQr1rG4q/d5Jn
0zjjjOtoK5I9hNdBx+bn5AIIZ2kEcVVILx8pGKOxm5+dm+motajeFwphHg/8TKjDvBMT6Tk/5Kdt
GjCguSLanP3gYfPFN+TdndFf38njWd5yFC2+GE9hCuhdpZwMrJ19OXr7KGqh1UM8Ea+nYr5mND6Z
+q2bU7hgfVCZoXtetqW+WWdIFqTddzi/ib7KVdXoBjhCAN8tCqbj59vjmjWLfoXGxqi6fd1sIvbX
kxY86cH8bCGO6d220cXS2Ki1Y1r5CxBoqqvulv+dCqzwzw7XY+M0HLDbpqdqEDumWyPuftUBb/K8
Gl6oyjROFx8vL4O6+Qn34DxTMSgnjkeZun0zbUvhMhBP2ToUITJIyJl/dNp3UntbZXd2Rh4dQBRs
XV2eKSen4/GmVVRtOV6VctzuYrH3KyUn3xWcppeEG6RwJEH2GQPnglFs9eeAj9PfbEqwoMxPhvHk
nlwQdRDpaiJKo+rXTyRpfx7Rc7PsGUR9mr58z65gDERJUbtu+WAMEcBFxlBa/kXuuTPkgV0ANocR
jfk9NzfssBkdcqRwv93qDE/dzkBwZ9O0Wh2kIRvIC9D+/97ZRPMaElPp5cl8v/s/c9+MJbQ8caGr
cObzxFTXzM7+W+lWF4jN22ufim+BEzRb8/7BC53vwKaeaqdFGdYNDdJs1as91LChDF8WR8TJpeAz
3fUbIArRjxXxWPxk15OkCBlJO7IVgoRp9qSrS1sAP1+QlqB9HnahWn5w7+vs1KxuM0u5ikO9v6lH
3YiFP5I3JxSjGqD7ZSwsyK0HXmT7YWn/U3vrp8bzR8d2ZnOnxFBywTWhk1fT7hhz0diDcxsC5PS1
5OF7za928EzPwhalRYohlihaHIfTNoVadu2avXkNmpNSPbU94VPXA9p9EsDZnskQFqS1fkStI9y7
vtvw9SH5VO3124+bYJZe7vPMXk0hTT74QCnhzjj5+Ur+o56VzOclQGWmN63gxkWsrLRSE46BJJJv
AlRtDez6Zy3IPNBzusCZRz6Mp+ZPjk5aCWmgZPLLalRv5QCEj860HMMIql0Y9eVa4aXAfiXChkMJ
UwiZokTJYD4Arciu67t0oBlkUa6HD6+A8pj7jrHxvQm7Pgd7cdRiqfmvEKuM6MS9sYOLbKNDSMpa
o9+F4gp0lY2oeVZcPoSyvYyu1FXSTo80ZIfdE5q4rhnoH0h4OrmDVfWV5Lh9fHnrcdsUGhxm9Zwp
MN7Aabrawo2ffI8zAaT/DEywjisv+c3oL6QM5Si6aKJt17wTLqruoTVvsyCIR5dYhBR803Sfg/LC
tng1tOXAuy/WT3/3kaZARDKzuFMIpm/ThS1eIzod80fXQHnIrSSSW1wMjLquXVnk0RA4OrCwihUc
uMK4Q5q3RrQNamCXx1igUxDzkZzj9ZWviQS7y0xvrB7+m0yViayYCoNF5oFoACyxViCfdguEHsUR
+xB72F7DzmivMCpYLPV4Yx35msO6CAnKiW2WUhP7jnJ55o7/FEk+8F3OoPlmOakCZhAS3r1vutrE
S2RbjjGZyzGaWZMuljIZkmZ4wHYUMV/PzlGSXlYASOwBt6QI0bCUzGyJqWjO/43/4Yza/4ef3nP4
rFRk6c8FKwUpGsGZumtcMPQSy+EQhej31MI5iMzrXX92cFd8Dr2AQG8I+tJzObXrvbO/CoyAnJ6B
fRiiWQ8WK4pFgYPYWfr+ogUw/yDDLTsc3sP3ootM6T0fcSj/z2kBsIXUMPvyefYA9bWnXu1yjxkv
sIjdsFC/isPKBFwDFdfSFynk1Rp6NvOKyIpGjvBFmQn5UM9aWJDcSaeoXrRlnRfODAnvL70g/vjN
O6sMVRVNAPWDWa2xonfsAXNW3cJxJhu98RsDSiuL44k5pACBZQMpFTkO8spmQaoxhS6DKqMmqY1c
nBrPrVk+Y9ULHM1ctq3SU3k4mnX2u039Dtz0NYTGL0j2gq44zBBKQHyEuJLxfI/wN8BHjTaFRRz6
El24MhgzG68mLaxHgVKxV6xyhoWQN96P06LIgC4dBqS67bVu9iXlZT2dALsp2dVKqib3hNRY0gak
bpdMtHsGapR5SMN2bwFnhG8/kzFIfQKp7oJRQVUDBmTFlHBBn+OtwCajALWl8QKOc7E4AmvmaDoV
tiV7DMQGIzaZCU0OlIIHMbC9H8jDMawIUFgzgHDr7SJorFQl69SVrr+5ttnTa0b2tZU1V2oED/jQ
8I2rr7XWiqUBLOC+wV9tbgiX6rIDrcg5I7GF++/wiugws91U4ysozXEQ3VR8MgzAyN/0XcdVWfkA
gd4fRay8ZyCBDvt875mhYUha5fFgx5Vj0VX7DbfhjqDCAcALhkQbhu2H7s/2JWaeU97WvVHG34ab
AGYDV2B/MBJaWgcjeQMKGvrDchIeVRtH78cSd7FCyou0i7PIlLy1IBKAQdN1q2YiyWfKIZcBicq4
pZgZgH6Q+nuKexmY6Hif/f8jJkPJH1P5zdUngD9H9WFhZFJJIwhzK9RG/ebcKt4CRzwddJyodL39
a4kSOoh8vc4ONKe/tx0mmbrmEU+e7P930JeChw8KPUdWqvcP1oZwqtP5WEwFNp/o9Qnb1+s7UQYX
Q4pYjYNXASp0mpIx14KDdUXlMy+edseg8xD3WXKae3wrZ5AWBD1qylniCIMT3XilWDtToJhwQGH3
yyb6mxq38AXUqNDOekocBaRK/XmA0Tgt/HIFGFQCZm0kNBIChoRK3N4Qjvdvs8r27hO5USBJHLew
5dYxdbu41OXNdGp1tzYRfqwAdmZTTOsIL6KcB9jV+C1OfpvPqS2M/A7V8e+xDnsiv4U38ih0wgN5
rByJalkacWlEBZQRv2A477bTnXMaLIvXwAHaR0pUkdNzo2DkuuXYyxTznufGjCw0VWWOLP+DHQTA
4a1J0QtXTbcMrV5RVwEZz59jm8L0VWc3AzG+q9hquwRhvHV5PO2pMlaoMMZymOdszOXAOI+h+WVm
Kx2BeGx3/O9v4awGzhbEZwJUiG4AWXlEuqqS7/UvRlCq5RzV5ea4fbzYRQvH68naiBo7twUom0Vg
1rr5vVTnYkERGXXypjHJV0Vco0tpInE7GoZDWpkcZf+qHwTg1pSjFofr3VbKbHhJN2tvMv7Em6oH
h6FOdtrhIQXNCQ7RO3uIcZr/P/3cf2ALN6Zm2k8uamCEkzJTnkQwpJZRgYOrYnBnonc39dkmWLUo
Sn6Bhs9FyS/VNI8FsVifVhSWOzy+14D1pL2+4v7HQPpI8bX2dEAOrZe0+AHl4uCBOelWIj9FPAUX
7Ehw6X2585dPW41rsHfLP50evkRRgjccuLt4LTIwFsivzFocSGw5bVxDGV+SYd0jOgSi3SkjoLYJ
5ZV4pHuMMBDTj1/cWB4wWc1a9tH1vU/BrAiY6IAHBu0fzJ00C+ofB/1riNmCeVTHtO/MF6TzR+io
OIDQdhbX59SAEhhuqFK4CpWXVXVHAWd1RrC+LCVr/lt4zR9CpmtB4Z9sBVuVRskNi9WZbCmuUwVn
xNIwzLRa2qomBvXVppb6neJdquzqez5/IYsBZmiAcYCpGRx4obluBNMvX3gGA5U7QxsUgopTzC6o
hSjlnCsTIYA5/fTeEIB3j6s6X1yjSRfeOeu8E+43ngTuT4gbUYDl9UwgROyB7LFGyUT3HL2sprHE
NAtRkkLyCXQQd6i6uaRFfkkPXfuw2eySO+35XTiXWRe1aEw8Hz122rq7tADMdK/9uzJsZv2O/au4
DAqMMJBr7EgGJDvaQoYdbqBNiXDkiEcYQ+HMaKE1cebytV16UHQBORLek8FVDoa7hvXXNxkLoNpT
5CUpnreR8HWuHPouzuK2fwRJ+Y4nnU5WpLDqtbQQyrmKjRnENi5n+Ck9TESdMN86OEL0U2TacXbD
Br9tdtkc/Wf2h9dOcQk3g5rs4PiJQk8EbsBquU0dJIO2cu2mNJsAc9gTbD9WRJeAtbmqGdqF3Vy4
r0UNRF7cBI87+hfHTHvQK4GOo2YBUJ6YDOtiPP/fOAbiQVmDxT5s0GDlNU2eHBLxs5L1wWs5x1Zb
DE0nWcmQxkIhDzwt7dfDlDnXAJaXgAx4A4HYIpOglQ89bfRJ+drwDrMYK3fLMIJZ60xK5PNWADLp
wBffEkfLQl/vCfWbzvl4rrZHIR3NmFgE3CcO87zwB3PYxyiPoSHsuWxTYc/w2u5MeiDwDx4bBgkg
3QHrJ5X3d21MP8j83axFvhycmEF6dBRf4D/kkvrGA/ha4sBWjZtXytjggfbRnr84hSeUVVeaSVRY
7wpI8KY6jRaV/AGlAeghhzqIMyD5Bw6MmEoA/lPgJoOJ+itei7Xc3JXgKbR1clCWL69LPEhF+xP/
xk+NasujOxcbUbeLeYp5JvMZqVHtKMV12PtEbrz0pCG+X4jKB7q2K6nGSU3ctPGNSyOzkARl9jSi
c4h7rBgEkBpjj/f1mZq531VxiRIFRM+Gk1rogza+zIMhkbi9VuF0HZEoiBFsVUhWLm/fDuQTcR3l
dT8nx2tI12uRe+gQt0lVd+iblB8N2xk1LeEvaRFagoiJ+E2yVsWclbx2dJF0mFP05mhm60ybbd2i
psrL3VsTzvf4/XONZZI6+fXhyJg+2tO2O+EaIvjLg2Q9twXJyKLjkwAqu6xCjEluFkTfarwJnd0C
JP1s3ZYUCwQgCbWclYG1gGzGfvR0RFB/DSGMgvsvOujfk/it166HIQrhfc8tpXkgcJxGb0xgO5Kv
qFqyQS2VKHDUpmn/GEhoeZnGvTQIa9z7X4M+E2iZDXVQ79sv6fMVDAVygLPokmIJ6F9DrOmtWOcv
PCtUwKWv0QIgFOD1JfVEZ3dByUV2v4PeYiSDrAsvartGUZM9+OVvjHJW5lbYAClLiwhC0jE56nic
5Gy/JEgweEzb0quX1THyi/4UkqxHlCaxYnmsZEEv6scMr/gmGhpKAP6H5lMQPDb4SGvCHlBGgCmo
3ki6m0ouxUfkPGM7apCPxdBuMXJDGQ4EQdkhHauNhrpY+MptW8grOMJyr/r5Hugxzza2iKSQ2jEu
sPi2ZdYU19BXLTf9fP8PBLLUADozza6U1+omv7fW4WlBwCej5KYPukJysBDb3qEYaW9s5mrro0+W
1CqO3E0CPWBaBB8EoHtPSjKvGI2TB6lJna86YSGTwcIveUvrsQy+fKYKxTE+925rz4uHst/INRUB
QO8klaMdePSA+qGYpVIB/xWTGnm2o6/1lJIsyrH+GYv49U8FgxNA+i/VfdtSeFYwdNDHU1wFN3MV
BN0BwC6fXfqviIVdsU3EMsDdvRBnhTimD1w+56iy+VEvacYkcYq2fCWX3ib91Z/8lpWwQ07XIM9m
OEyXEyg/rjoEhPSr4EZlUN80w/gmxK8zeFjL/A0DYsBCTaSmIQBxfZ6Ze99oHb0F1SKCg+bptLCx
2T4Uru9VlI112p+JV2EbWxotuGLqw4AHsxW/mPpitdP8QmHO2ExTa0+1UvzHP/IEIu4phxd1kMkZ
xnmxn9gcTZDimjDy7b/vtROzqSB3Anoegwsgv9xggX0rlUhkzEbN3zcpa0c+2FpLboOcP9/G1jwh
x/K1x/lHCNDANmquNez0qdPqt6wue3IgdGEDPXVH7CGiKLFW2mxn6vQkQGQIAswE3HBuAHhWLR1r
/Ew/RqdeePiAQzJgXIJwWvEkpHZedOKv5S6++BEl6di3Y4RRVzhaZjlaIg608FMV3HW2AHPmdWeS
EHmmmYBEvV0BUHEie+lrSwCr83BbphSGgxoJYUgZxK+Hf7wIyDKgfUhnoAiwTD0q93DIusn3kZTC
v0PV/vFTIhvcSoablXkwwjP82fBlc4s+Rz9Vhd1twWSjzxgMg8Tq1K4GLlJtvOKdOIQk6AikMP7q
1MGgoMSefn5IbyG0qVXDUvpY3aIovCncDY1dRtbCsBI8g6mzYPd6YmRiKzOLJiZ5bnniTBcYPHTT
U+MF2RPpocFXF2GbV6BG4PsribsedKUaqw8FHDjHHH2FqzqyVieltxRrbhnvJgeOGW/OZtnsRCA7
9oS+k64KKVYgy8VYHU8NSYmalnY62x64z793awXdNKa49Kh5W7SMvM6My+CEItBJqa/pXARQk7Cc
7Rw7SYKZF57GLWb7AjfIZd8VCHO3w2ICihiQ4hsa72D7N2DcHEd7CQUjIR46YKtrtbihxqlTIprr
yokQpiA3VC+XjuaJdVBhcKyJE/s3ulf4EmgbZTI2ysZtxdMmlUpydojC20W3Z5t9+NJRb+iKu28x
wzyKr3zawBMMk1Sh+ykyiSD5qPgQLrAOX65P/YE6OVUVf86GA9vOrADuO2az1zXqNH+hp3U0Yyd6
L7WJOeWjqh3WnHT9Qx6KQPNmoM/nQxVUnEZtI4joELLPpr2dqEDMbrMGj42CoMasnZdwowtJ0eGU
pN69BBD06k9DXyQ8gVenxoJ9htCTMPWQgG5yDtwqzTDW5DsmcyMRWt6MyRYxw4dGJPRyx2G+Fyiu
X5jPJY0jvtH1BES8qKKn3RAEodtcQMRsP/x69hKC/JSPuKdrjv395iJoXT7oVAHLI32J1iidsoo9
Zelgm4kEsqhA87UxzuwTqX048lieaA7YSyvV9p5ulM34heSn0Bc1kFgfxDIt9RaHRZJaQ5PCcUxL
1uM8wIjX8UfLcwdzS7u8E9IMdggXnOHEK337uuJCoqFKU3GZ7VVWIg2IdmTrY3HONphsByfa3Dim
WR8C/bF4AxYzmejX2G5qIt9Wpou0ezG0WdtRrHko+LnY14BcFdmYpnizanUh/hGEJyEhywz2P8Z0
q0J9RWj8lhp8W6GkEqnNRErOtTK1nDAFi/RFJWBZi7/H2TNPyUpj8FYxyL//4i5h2eVvZrowAk6p
GGX6xVLvnobjk9+NohCBk9khlSmFLWvEI5rP8v2q4WiS9fEJZvw0kfEVCQOjJGKWx3sFE0CUjPQm
tB9fr0wJRT7WB6nD735z2rbjxdBU+Wfk13uiPiWF+DAJ8DW+vmiSkGEY+1b+UDZ9fP4S/Zo1+rFL
tPmY0HMKC896b290YvOQVPb27ft9ZrgmdZEXXwrWe//fpVlF+AOu6GOrgcBy3f9cCCPTPeAoj7j1
bQFMuFnKilAAmd6RX9ZMXQWOo8pX1+3zSuR8rKQu9PdhOsZyIlK0NNqzv8MTk0nSuNkgBiOkOVgC
7z4o+a8dw30p2TTIiTLXkegXThJzsCDWUKtVwEFFZyUNeVM9aDFy9qHib1Zdc+Do95xGwuzAXO8s
AMdHsHOjau2L97LdRIeG+m9WqAgU4BupExk+bK1vupMy8lhShjmuxz9xY3Co5Rr2a9im2zDDfey1
coG3Klhfmp+ZLTD9FoUwM4O8R25FC++hJWyYcAdXfsV60AMgHBK/7iHRmr3i0F5JoMc2A5vYa2mr
udbMMusjGNd79/jPcTlnWW2TejwJ4ENUSZBS0A/kvMFsG70iQPl2iku2+vxDUKtngzPbdN5+YDY4
DH+yaWdSLnVB2/UJxUMQ1KrmHwv9xeUimnsO9ne+IlNaXVy/VdbzosMPUtviPcuGEflXcik5MObH
10lKCDzUHfH6il0u/+3GYlwHk8A+6fyXf4ip0406lihDAyRO6Y+0QU8bHw2E6nWhoSCcbJsurSYk
L69OtzHgvnyY71eFANUyfAgczFMnKk0YD31zacJ8uugrr2IOCo1EYpRmwDRM7engmMnTg4UPubgq
oQi2ASzDAN2AI2l85D4FaEJMdNIQwNbbfsZsKUZ3yAItc+/VU92GuSvGHrMVjrBvXUXbqiV/Jb6B
MrY2T6Jc+Hf5zwOokWqBpu+ONRcl0eJyxNJ9viD2CGd81bSGse9R0nIF/tP6zgeKmYbrHaPyjO7X
/1rnZmrONUfCmKS/wFgs8UEHQRa1y/yE5q2BV4P9enQbmvyMUhdY05TqDGqxaz3oUk3ENmkxfFfc
+hJBBe3Br6NFTZ/ls/O4N9qP7kHDe/2xsnwcAGYS6nZlxroBmwoSWfXaCk6O+OD9ucIsdoqOiEIe
nyrMJUuhfXQ0jqND4HmRc4AADY62TQ1WiZzdPWsRUhLbXkFtG9ngvYgMymww07RJ4zJc3GJ+INlX
tMbCXW7jLkaeg6DQlP7GKhVxcEuvpdlh86xHlJckmBC3XPArsoI+vKJI1j7yZNg1dKLhityojh/I
xggtK1hsx1U+DpgU31pxyomQEW6uv1FhNY8WKLuhSoNhHpt+rs3RWBIxlCM+TJTBdva2JxRMXlOL
xF+O7HA5jzj/nYd2zCw4Mn0nfaiKahAYjDeDIxQbChXeyKZZD65jPq2r+xYwDTvGWNDKmCh/kik5
ck++dZ3HUP9K8kCITvPV/5Z9+G/S4mewykMLEVxOzL71CXvjXWmubDCN6bwOV35GuaMTh5SndN5n
gHBtICwvBjAyoONiYlsSvn2eeYyKgFOlUsaxOHVzuyxkXloEzGycnS1YXflVMegjqfYGyjl2bMHc
ZZoO5lKz9zDkQ93Gr385fFKsR1PVuZRFLDCHjwWYeRubQ0USkfSp5G5/NKHxfcRY76G/AlqpWHS3
0rnywbYZYSXjXLcBbqGlZ/DTfpNjem+7CNqrgxTWNR8ILNwnjRKBnsL/swClDQeLQqyhGsaC8MDT
0YuZYQ5iqpdcmWxq19DrBWrrgP3jVaidDzDewOUvGpHHeogOELGyHAQ9Eix+3wieHVw4TBM6eJDd
9v88zhEpHVoZeq42imy6bDCTUWX9nLMxVQkq5abzVR/6x/Bg5MGLsQ3b6z7H2VF99S+xp3oAn3vV
TRjJ/MqDCjHPwaRbutI4thQmH9YXRsNMLT76PEzBdvJL/9qUURW9D0LRx50lTwk7jg8EhU9fYVYH
9uiqVnzypIWkWTmG35p4ffOB2MBevhCLnpiXtHY8s4jO2RibJtiEngwtngqp9En03YgRq1R81og9
b62oCS/bTSOcl9jt3W4h7ph8ZeSz8qXrI92fq1ZBXbK/PoE3XlEzr6XkxL2RMBTICQZzSKh74bBp
4e+tK2mUiSjLkhoO16JzMHwSxODGzNW9IjWYhYWnNAvDjKRRlg1phtZXpIKxpjny0b6GaC7+++WB
/G2mZMLUiZ+pOpkt9UBGtlskw8Bu2l1ZwwXyLwqDylOV0UQwdK2V3l/VewCXdtf3bqGnn+UGCmKa
kOO2VZM0sD6YYu9rPNYjIPRsAVJdemxFX9YN9IjjzbNqPaJwayKsbLJbUvpL7exi2tLx32uqnmxo
EbM5MjI0YFNzvKFnZ/S8BVHNExSYotaWm1s8DO5nDS+dXpt0UPIrMT3MQ50mUqplcN/wzQ02K8xo
I9EBTca6rug0N3w9nbJLjo8zQo5vq/HhAKQuMwMfyq1TmanAl2qQnNfqK3s+gKw7ezk0iXFAOdM+
YP1VCdFV+m5gYTqXjjnyz0o/Kw/STMwpx5hgpDaWiNFAsGtpyO98VisMMK6LXylpCU1WElwG4N3+
/BspMrZ+t7qDVN7VzHLF69u7/g2Dvnx+07mQO+tX5AT6ZZRtVOc7K3DE+/DK8YBOq0ZK/aEiyJyy
y6dkuaFd2J9y33PeKiaVzIUjUrIFTl/SBb02Lc7ScLysLYUfykXThccEMspWn8xmNbuZlQxhZU8g
kAMXv7U+yMZLHrWvef8+db3l4psT560Yt8vRTtjdX4XAe5Lky4qO3WhQm+OdzdOa7Jz6CJ+JEm7Z
ek0pB9V53hYGogR5/nKkB+pBSABrY+D3LHxvmgxVrPG48TeDKvGG2IYRlmoobDl5wL7Niw2BtC41
pyg/biMWHxuFwPOIWi51O4xUd3rgJaX77Sj8Z2LVIduMcIfxAsUUxDaafZTmrqL3E/AcvbvdwGrh
xPXcNMk76vIkt6iUjzGyipZIn8NjVSSXyqrxAtVPQ1i6AwAA5gGfQzZk89+NG/1tBDAbGNmMJZFx
8hOG+Rg0gAb38M3q3nYiqDLt9YXOwTMeWaVAAJJRwtScvKBSYdtp3xFd4lle71nggN7lY+pJdDWc
53lVr4JCbiiD0gWg4PNY8UK7CfXW62DFZWFOpmjqi0x9CfpaZQ9kQ0rflgDUy4Cpgggs/tOuOFbB
cYahrzgrDmSjGL8dgFJyr7HtQFCW1VOi9JHMAnr7I+56gensRaosBngayk+6x/VPiLMF4EJ/r7Zn
nmiQogDje7dd1cPU7ZSr7CSUcuhtmSLlKJWc7Kle36bd5V7quAy82mWe+MeXvLuQHwO6bVUCk02s
7ZfJfF346NDfzpIoJSao/1jxxeUYNiwnlVJ1q/d10li7a1dy3KxjJsQb6t+4mL1yAANwTuBSPZ0c
C3Hi++iVhvbRcSgpNwz8/XZuZ+TaC14qU520ezOsrRQCMspsO/ZF7xtDsooEYodQodXsT/gkfesQ
EbBhqJ7pTpm7uB+seAHCeNgtngrmi3WeCySYvs7PucHS/Jlr19j9NL2FXeSYVSdvU2cfJEMHoZhT
8bzbPMprkyYV6SyBuEziDeurkPGR6FWrCaMz+epPlnF9PzGvcgqjnTWe37MgvvIKvoTTOlL4t9jO
1WcTusmStDzMbEr1PcDwqIctzkiThCk15AGwZus7EOptwcxBSfbiqrbwqP+4cgsua0aYDiUgc6Pv
8bGfD1ClFLoN09ORkZYrntJlgYmLNpuCPrsapfEc7njHSNPo9gJanG93Z0evMjjhn0xqc29ollXf
Gau9ti2fAY9duh8fbuZMCyYcPrg8LrIfj9eht/c5Hi6WEUWpzfK0ahpYTQL6nfWNI2UOhd4HghTT
Q8dfHe+Cdrad5oGip9l7bCiHBTbHVP2KQiUvngb4SPf1DJc+WtXkhYhjiJYTUlXEajeUd9RLCCh/
Oflvg000zUjGxpKyjeesKXQWhUR3tir4qzWhwJfwnNkyHojbajePj05180Q9dONSV/t0OGNOhoE4
4FI8aO4CD+2Y2Cu7QoxOgI09lRmGotz95fJbnffMHL8UnU4cdCtd4dR6dvMDaW7N5YLhPtH6ajwY
kLFC/uL0xXP23ls73krDNbU8UzctX+t5/9dCZx1d1WfapadiI4oMNXGcAdKaoZ7uil3t4FIC1py0
iI6ltrLovotd2vsD0tv+/9JBeHdwXjaY6QRb7v2cpK6EHWgoOSEzFd/3YLa0Itm1iDjls9Mamtd8
J8VmrohWtyaaRZmjWis0sxg8I8SUPGNKGWn2rDZ4Q6htfL1lVl/qGSMbuVcpRX32Q1rcbXCh9Ub5
bwf/mvMS2L9UaGji/Ez27e5HJY8C7hUxkF/wfdZ5hb3O2VFs4gXJxVBa7rB6vk474NAcXRtRoX26
9naxzx33ND+U0Fdb5RyrmlkXiDcBz9Okm9c8gsUUb4biaANfLkTAsQWHu0J6QqEGGPb/y1aoAK6f
eapgfyuf3B6SeuPsIzywfO1YWcAzEVsZeo0rl/mZpZrAfKOdsCD8NxzfhAFArqgFok2UFyIp4/Lf
DnaAQYlZ8XN7tsiDAl7NACpqD4VcADJ+FEznxtDPgjcVN8eE1+zGWZYMaX9kh16lFt94nWOU1/ZD
IGpbHlP0ql+2SvZ1yVm6agv/MOGMEW9nEWZgv18H7W7dUPtyA7Xkud60okKRqPEzrXdVMMEz+6AB
29UjLkm1OfN9WLYx2SVYg7+DXp36Tg2rngAtZsbn79za/6uNCJQeSXFzXiCc0n7tIjVVzm/QVctW
nmYSYA+KCDBNSzuxYPKZ9gZvatYKO7hEqXyIPhUgBW1+8L85aq5dgvwxL2Z83LkV/clobfoAggOK
agKBfsZSzSe0158o+QTg7hEFoy0CU0FpZtCetc5SzvRaCkK/QWJoriMIXWsx86x6Bue1hFDVt/E6
XAWu1U+GIqHcJq/So3pKRJWl0WXzcRPLPZRGNG4W2B/vuU06ko4Zl5MZ4NqTHK5FWtZZycKu7E/+
CMqLtMr9858gKBwT4cCqNi9GKX1Rpdy2LG5TmeDDHQZFc55ZdPAQfXNyJSALTozb3hG0P+iFM+/X
CU4t+/MsvEvthp0XXo/AzAh1oLpiHggoOjbKpuyE/dV6T6vnM4vjH9m1CvL74kdHZQywkTqntE3l
Gi1Oom9vlVNj+hygk9N8Aj0R3feyFKcDNTlss6qNzmOTd40m78XAism5ttDBaKj5+hbGU79D4DL0
xj/VNUtt3UQSlRtLCo6r03nrozrGU3RBL9JFR80uJCGGxIZL+wYbcGLQXMpRnTMsMI1IkQlD9P8S
yC7ws3e2myHxZgSYX7Infp3v8a/aGQxz4kRtVCsRxKhh6HxLXl9OdY0FUgkjrQ7R69uh8xTnOGsj
iDwouCtZ4x0rleDx9zbcT+03hsiD0XMCXrOwJtyTfEZLhPLaFJ9uvjuIR6XTcNe7OQR+4jOdaSMa
bgr2HZYUZlNsGHviR4vEQyenlXmTRykLirkO+kc1ApLz+O7dRPx3MlQ06UX/BGwvcSoUuslUPSC6
5und3wDor7j1fgpQzoeKtZvQL1N+AYelV6KPEgzBOgB0pgdT0544zSk84Cbc9+nSlbAqayNfJ9mv
w3lIxJKBLMlq7WUTpwH0hk7qyv+KSBOkEM1YEy1tu3+Xg1LhdgwvMHE5ejOZ62m97nNnPaUEg+iW
5rEFM/EW0T1QETfxWQL7LoPOaFEKuYnIC0Qr9n/g7GIY7gvy1EPM0lZo7LDPLWbKMA0IseM/w5Tu
5pzYMm5uNhhk54cnIPsaXcAIiGUu8T6NuZdD1y0ru0JoqV1JhvpXsgkF3CyWwcwBgVALh2BgZLAS
drzHSRU1rtIFaljQA8GtWgXUsqM9pwfrDHCreMIMokH/NEXtubiAuubK32dcvZzaMmw8gsVRbUah
oftb6hJweqOMAkBBPKii5sTrEyMvlxuYlODk/cTflhIOXW1KEHRa1e9BfqeDg2qJfjooaIK7QrY8
GKB3KpZIMOVJwRN2R5LxLwp3gDJOGiDI0Toqg1kejEnVdo17X3SzV34NyRy7HQShKqzUc10GeoSw
+0ATUVd8PGGbgyfiDlldYzEdKWxexE8AboX8uoSMUZ2zeXpkST+OfqH+HXHgGpHiASIWVt4mt1Zy
9sgjU1Byiw8WeoNEo9NDQIrFZSdUK8pFsnkXSNOHgKxndklOzQxHo+8tZK+6yHSE8Ce7csyOogV7
iRCKE24Q7+hDZ1k9wKghMLrnJ+MfhFtrDG5NuqlWkliPMNJM6X5VP8YTWuJesi4r6x0vHFdDhjL/
qy6pc9vtM+dldjQb1Q9/jxJ9mhBR5+LT0RbSuzIU5bUd3M6g7C5f4UWZQAEvjIE6mIkYG1DnsRbh
bn8uXN6j/fHcJu3SKN/B5Y4Yb3AFFK/BN+h8PaR86cgg+YQgDx6EWSk3pGknV3ipRyrkqFHa6jEh
o+KI2oiKnIydEnLuph7kkmIMGJI5n2VkbEKM9d/QSBrwbsN1xAmbdmYiR+WIfLLd9tMtHiCbpJV3
tok3/YxsPv1an/4CC0fMjcrxz0rpls/L5IcQbBEGNOXERi6o5MLVduOoRAz5vK+hyl4r4LJPScBK
5sDSpZdlBrLPouh0hexASGM6TBXWvxGqBLWhOmmCLUkYYfATqw2OBIEtZiLSKu9WWYUbClWMN158
Vg7qxuxACac7i1twoDtGZaDNMC7KtVgVKj+g6UkVId6UX1FPEQvI/hLaKJVLk/LU74ziMIPHWqya
jEYtUkEv3MsirsPHVTH5N5Oqpw3rFhy+6w/O3cMgbRE4SpJz9Ifuuycq4s+s0lcJbTCOJL/NoHLD
VboYfOpJhL/dGaRSE3HVJPPhRLPLkNK3xviOmH/+sNBuKxHCD+6CvCSDN3/lpehPMuDIb3+77Lqp
puJg/DWSNpzrZj1/S2ndAjDPvNNnNKg5VeF++0RvS4MJAz/8TMT37NTV69ig9aZ6rFPb/8hjZa9p
+SjbERIibSdXFY1+sKMzK30U9hEKoTWcoYGJDjGtC9PfuxcycxkxdRObVUXdNhi05yBktD+VsHab
4JEAKF+k3lyrVJAAU/amYoVuDbdOqF4haiuYoED3uHG6QEljHku3Td6cy2UjqhNUIOuTWg3uTyCT
RGHWwcvRX2/XBusyycKweuhoNSjGbWIkoTbAr/isM5pPBfdRijwTkX2bURWJD19+OYWIfKbna+nN
NiEHH/eEvl7QqC6zSq0Wo2Nos3da50RhfQWNxA4/C5LA/lIrqxii9G2LX4XtT6elx2sHvEjoPPGQ
0CGRd9u2iivVoyBdR8ASFrdQtD+M/jQAoduYo3J0LTre6l0uMAGmwbnVIRgsMqaAtOQowfxI2qBc
8vnSH88fzctkqmAollYwlCkq55iVRjTc2y8V8Rzf6dn2iZRBkFE7T/l2v5HL+PXXyQJERpkkQ4BV
wBd3jYeA2JOKroNvX8586PZlwTI2qYMVB8LG2w1780o4dPVm9Ip3FFjL8Sf3F7S8dE4e7P8/oevf
fNPZ0Jc0MUUuyYQ4ANWDmhX6+hYeBlE5eZsh8h6qJWVTtrAgGH8pf2lZ45/tlMHjaQpnJ+tKLMpK
cUMAeKVvRbj/wqmt+++kDrpMD+0Ox1DnxYXixcbNCnR+tZgIlDhNslYZsEvDlpOMjwSTT2902csh
b6MKYaAABVwqj+3+7U31FGaARDA2CEwvsqF2eBbknz+NhInpBYvvVX5bjYWUUAuA0BjRCZCOyFRB
zx0HDSP9w/BGBQTFrzindMtfNKLZx5bqXY0PU+eRZtw+BJacxQZ6JFyjaV7nopTzF6wyDJgdQO1V
xIIdfgbww+A7onW2gAaWng0eXwZSikOXCfktETO8vHFxjf7/ABG45SHdVlJXR9ssz5lt3n/Tbvu8
vbrboAHz8QarIsuI98olMFEdCL7xMv91LRnJGhJHp5D4RjszorCd0LV58L96m/2vJS6BoCTN+fHm
IFtpyHWpLlbdw4ryLraSz7HAvcXzTPPL/vgrfLR601Yk4VPscGLQhnzSC+q24zElQKKd62JnVXOh
UDFl51iXIeICblWrBUFOFA8f+nzvR+1H6po5x5CoA7wSGLmmGsL5xRwFvTv4sb7bAUUWrIh6mpjr
BA1Zu3ybXtgO6kl+e6eNdxYHA4nupjufUbHaDifqcxaHWymJhyEmoaNhl5b1tdFkOB7HR+SH9LyE
ept4kqO32U0J0I1lsAD8HnzdwbBVKwsPPnK1niF89nfCqzdm3raHbq91LI8nq5hRP++/MVWw4sL1
ckdjQQ1m2uPiFI0DfCZHnTVX4MfrtVqGLB0nJjBcpxhFiMxZO3ggtJ9H2+7lh73eFsuvgg8KSN4v
sNKu1U4lX2zer2J2TdYt1NnjVnEkFny9Yna2//cPnIGkNru+XUx2v9cwMyfW2pAVK/BI+udSug8F
rNsEWkj89Yv9EmsnxBkZM2ZboK4ph0lkzAknXgsDGI2VcaNO1vc0k9GzYTq8o+rAJmzwT93E/hGM
zh0uYFPLCTZjeGwACUSsblHrfzOOlTMrupvkji+Z2feUn5ZASNIz27uXhqmrrl8BfVqhW+dxBVZG
73cbwinUDjMSMfxQb8XiHG95HNzphH6gKJLdNeDADtqEKK1fnHLSzjhNi2KXGnRTiuJ89STxrvFD
JP7GAaTgaA+denx1XYIeQ77OVnG325D9T+Rs+Lw2IAp7Gg8x97RFDswa1e9GhwTeUzAs/o6bcPF5
4P0XU4bm03ekhcHkSK0K5lVzKGtqth/94+egLXY18r4g6HEkuQrIw60Wfd2bT8Tbf4Ha5OHU5WWF
4Z5fCpdUwRqjjy/GK9uCsUUTO3mSE1ffyI51RHgwbCKs9mW8uOe4mAmRHluw4I0EYWOuZUdrNFr0
0xAGZscsjefuOx8J2wQmkBbAT5LwVZ33VY2Ph3aVJRScom+6HwpqmU+TdNQZF0YGG9n5ffSgb64Z
tzqVf3B32BsZK+6v9Nkal4PO7e3DxFGzYtec1itNIgLF2aC6x9n2NdvxTrctdd/QLd3FZ/MIHTRL
XZQZrJnwcA7/UuaPbfMIk1HZPdvzIcmhILiFYs5HfHVkAetQhczx4iZBKfb2Eet+6q0mk0bVaAkU
udgoikiHsqzjpCiC8jeWNzZJLuz5JDsF2sQtjMBRxYb0FjhuwDzbKAbU57vgL9vP5w/ik3BxXxwk
pjYTjwe6glxHb/Dzk/G9725jKAXoIO6gsvHwInkSlluNwoFl2FCBGr8G8xo6NpQo87r4ykqLKj9m
Y9W98fxgu/DUyPhgmSV1Y9dtClgqLxMX3jsLDOexRwKg2Dt01txolDc83AQD1zYf9aPm2ERrLS6G
YahdJk1fFL8A2bWvDeL6rW2b9MspkkbfOhUf6sbNpdCX73vgAGXXK5ifAkOkUls/+AUebBjahQx/
3bCnL/zx5IlMbymPv7hvXL/iXPFgCcKawgr4iS6RuIg+QbdSigUzpKWBfNbGiPGR9CaFQWvNMnL3
cyV4bIuSZyC1Dw6aioaJiT+fhPWl1NCmpJZQ7tLxhDg0I1yc+FQMKVVGHSnn7O1NEVcB/UwqjyaL
62mxIXxaQb8EFvqnVeRPMV3xEycWQs604HOCva0VwQ4HaggkHPab5zMuJMOyBmcVQV6bHAY2ZsE3
srJ82vr0lcjO+VwhQD+K7OPPukJ20AU9xkXNy2vjSZ6N/7QLk8OHimQ53mCaLYWCbO/Vu5y0NxtV
2FRuLxtPbqKN0hjF2uXj0MRISZyOOsVo6XtbxvMmkLKZmbOph8Qer4KkCXFb3BSyAfwKs7IE+A3D
3nl9OjME1ZnPe3TBj/HREXfb5GORa7Jy48QoVT+NJovLKsuc/wnoWDgvuSPgyUeR82SZ9+dX2QhI
JZrRWcSJZYCalmCImGp1H60LBPaBfp6DPsyPZxtDSFmZDZtJ1Rr7hvxww6Ux3VfFZHlK90JkTtyN
tX6oQs6yoJscRQS9x5FQoyzH7iiJPL3S/f69d+8gmwWMucfdvuza+4QX96xOM4lkca9rBOSdQfRu
JroTBwRsZX7tSkGc+KvG7GvrXDmFT56TUSiJk8wwiymNF+/hpyto2YVYIknWht0G0BWE+GKgJZ/X
hqdO8s6xUAdmRLSt01vi3dPU2eQvcCVzUBI/fEQEIC6r/NUZsf/HhJR4zYT7UOv2xpASctkTybA6
x2YR7iYHpwY8K/c+gWQrRtO9jxnQzCZOjaWFIE984xZGG6Xnue30ilJfMlButgepdcVEI+Xgs0PA
rO+bZCxwMdT4a7GEXrhs0Te7E3WQOZRxDB9141MwXJCK5p0i3+f67OGDWKcqW3213IGFCdRisWy1
tZBkXpNfynec6jNGS4KiDAF+j+h32eBRVRfJIvhReXqG9bAET26iJZ18sDGzUFE2I0M5hoYRlYVC
LpvNCFHlda9QOsIkNg+yLb/QNqxPHH/rSBgPv8+kvk2G3nKeBy9ulLL00FMPEvvwoF2K5aRvw0BX
jInM+4WcxeoU5//6aQyrRS9hUKutZcPJyJO16kn8uhPa3QQD2QjCNrt8eoaNJyhgqmKWlgFhMv7H
+1bvhtDZBMiLPLIFTg3JaqBqaTYxxpX5zGqXDY/o4ZgAKN6gy+r1fOSWpfVG5r5wCcPBlpoN8655
Kk6x6CEOahTreodk94CsXK2GhJV8N4W6fjzGxxi5wsg0bnLkUfny0GW7/wfHW5Qmm3fcLXdSM0Mk
yhQ05xKOtvbMifNAW3wZB/wUeu7Uhf+5Oo14L+hRPDLbQpjtEAeM8ZfuXIiQ1mD+Lpz/u43a8wBD
1ujNoO87O28f2AYx9ktvbSvrXMXQvkkuUuRLuA1Z4f3LezQVFROn6aXqaBetxY+AJkYv0hWL00S8
c9mVeMVv8m/E9NdUJaAXUtRuJjH9allmkQ1gZJBedC+7fhoG1JoLpmNYrZEHrv/4/m+8SFpZZ/g5
sKVaYDNlj9DJMoSUIZv+L8LB1g2jQFdBqlCCqi2TXDLRqGzFQNhE+UgEfM1/KZZXut+f2He4qxcX
8L1bT7C9l6aA+dNdoApDrrnEv7fmNKgpE8HCkn2iOkgGSL/tlUJO/yPWxgvXjUeskYb5730BVRzI
N5BW72XdzddayUAzjG1/4cZp3lez6oi2FquK5pyVgPhzXCfNOwPylavmfL0kposPXjrcDfXNxcgf
W0E5KXHc0CVd5vZrDPeonAXmSt7eX966QqoIfWFeQQbRoPgNiUGX6wXG5FjXjX+n7H8B1BIrS4O+
9HrM2WVr7R4wKf5uL6pWjQCxFa7QciBKw5ZKk+iPFK6CFXS9O2RBRf46XKbC4xuQuf35SmJDOc7g
wKfA/2N9E6YVx8aX7LirQHGczCEKdFiOKsTK6zQxlcCpRzyLIg4fVOdCvzZWRNC7P4YPVqQdQbxf
ryGlbo85M4ojM9Wvyda2sggD/x38EKtJ6EAk1olveUjtLrAKu7BKPHTaFTLiiyKLHu4WRvNr875N
NhX3LQ5EOfph3ULbToQW0dlG2b2roOJE3mq8HHseDlX922G9lmE5oTc4/LUrZMaIEAqtyt/gEOye
vhkghjEJN/5/gCMj0sRFLLjg27lF5vLtNM5VlEX/bjeFqq4EtTnsBZAyJVb+IhM4R+vd0Zu5TSqn
WehYJCYTHjKdZsTfYqD9dGLFsqg4QOWa9wbRsbMD6c4jksSrcqEZoh+xeODNNt3Tdjc+u3D/t6vP
4VoyyP3G79Qy5hDk5FEE77ZlrwdBklZFti++cESJb7DxwZnYuzIkTsLe1hefSgOd3QKYchYDut0d
COmtTHaKcnZjaNxQ/6iuridOUHAcDfLVYoZWrUDs2XM/6XOTZX3DYNZ+xBEhF76rBu9c+jE2p2kU
0SLF7vasIv75r7tr55QnA/K4YMtastfrZDhV/lAU9k7tity79oONdVBhKa4E+Zl5VyalXi62YZ7T
CY6mJw7tduUl/UYGBKeRwJDLR/qXc//lqupiAvUTVrvxTZJnNbBUXl5Zf9RsDrsJKhX3oXFuiKaB
/QLoxqp68Ac5xVrI4SSsdcVhVOFe3GrJA+tsBJ3Y/u9hbQ2ooRyX9sKw6a570aE21Z82nC4rkezd
VPuV1I2SB5oqjlcg/RuQr2MVIu58BcIgxhSsbAPZi6gqa9XDaoXZCzfCp28JWJrm2l2V3cIYienz
+n45n7VkbFUVcFHujVZqBFIxvGLZe8+Odvtu47pVBzgIYAdfVCauCkNvX8SfToEsfvTnCUvhEXD1
3FJMNseCQyt3pG990wB3mNcPrYUXiXvSw0YLGcIQtImEbEyWA/kBF8LOowTBU+XX7sxAfALImagG
Irrmu1j0gAQH6GCaVdj0BiZDsJMrhIw6Yxdbl6eQ+O/9aHhK9uiR0J7Cc1JqiWOJlYO8D2ACM/6p
UJlQWaPUTofR7/4CG5C6gmb33ehJmINnJDEzyIvAhoswVp3o6dZM1JHyN7wOMeTd2apb/qJkVKtF
sWi5w16bM0Vyzlx2odqnJDyjFsMeBhyPMUFsjvBHEuO774zuGI7R/DvE8xMq39h6tsYLz8rhfH5g
HnSOrwb+YxtTqdpFCenLZBMyvNRcEEdzR3INJAa9VoVv69bfbm+fNtZVlCRrB69CxbVQMz8J1jXd
fxQXGwP1Uo2sIpOCZh9Eh+EWscyxhb2mWEhwhYfXFhWfUs+9hpeFueDOSYzyXQguKRfDV3C+178Z
pKnsLM5oltaMuUhkvkGEGViPOcu7tRPWVeby104dBEpzHeV7fZe5/2Fkj2AFOLQqH2qyxYhTnf5x
V2Hvkbxun39c68tiHKZWVC+yjKy9rc4dPKJIDb8l8d3SYe4WsbJeIJUKY71kTH9rOOb5rEBaYQ+z
IsgZXw4dWdP9WzX9lDYL3Nqb2NxmJfqi7GJUAlOtIyQRE6HFxA6CGksnaUrGQGM35hJ3BlWcweqC
KP8bRJXQUi6BrOj6gTKCghwDjgVHCDoAG8DmlX6aPOA5O6Hnzq749V555WPsbL3JxsnMTNAAZrKk
/PZnQiLKKSGQx4xqijjrsjhLyMGlyG/6QOkf3V3805JUYeiGjub0gKfPw7MUFs7aNKYvDYw0yxso
nNDkNij3J4WIMF0LJ2y0EhSgovkVZnTsGoTAGGDN2Wuxv3jJrVeW8E6xkX+gCw3adVVyRZ722IOR
Z1ZiOCJCvufm4c30pjxx2U+GYRPyusgMg/UGSLa+O6FAvBRmZyL1vZ6UACINJeaEoeZ07iK1CgOj
i2a1VIZB3IT1gUJxH6/b3nXMd2+vE5fEyAcEHt0nCNw3InK41+Puc69XeLJ6TPSnWs4OjLNbdplb
/JTZ0YS2lDsNK2wiY4invb+DzsblBIAYMCz0hYgrq9brOuhiR2/Z2p6T2e1J5krpKQjupMqKWI2O
HcoH7Iu6eN1wZ8hi5x7OAFjbOiRZtqI1iO9gdK5jlexL5MZdEo/G9GoASDGNsuix2fRPEIyY6TnZ
ahGmGIMSo9yL5O9HVhcoVxfevuYPXFKyLI9lytU1ek13zNHsXI5vRxYtPvwEYbcZWjobmoAFUlLt
koC6D4H6x0jFFLCOaESalIyGWs62+k+gdW1N9+d5Kwwu6fXw7qghkSjHqBLQ5oSDUtKFQrN5Irya
VXLwi8+KCNbVqRFg35QkWiKFnXQ/tHKZyRMw09I+vg6gUAg7yCszAWzR4dtQHcMxhUDNbJJYG1Y8
S519bKsXxt28dw5F7jq8n/NUcKPcWWeHlo+c4uzIV+6nCFIDwYfs5lgec9JDxZgrqWwYxmGbaGQJ
wWf0QE2qNeBE+YtNjuCvOl64OqAN1yGigIgVzGRhK9N6JgXy/ta86zHnKMWnhi9kQaKNp3nY7k5U
U+7Z344ZGa06IRcgcRMPVR6DSvafirH2v1sF3cndiOuCZKry8heuugpDqcX3z92T8vshbyctgFPh
z9B9BpMy5PDbx+hOj+GvHUNpZqT0+TEoRtYS0hwGTulSBUxcOTRV8MBDwozO+vQZOgCx5qU/ApnV
KUoXpCmf8Jk2E6HW0NT02NEHoiU4tFgyqeHxh0OVwaBLxl3/T16zpF5sIqE9hvbMMKmg0cXIOojX
LTRSt0vH/v22Ga5Xn/AO0JpLzxSQoAkfxFqcIEsHGM33gyDQWRAbn2BAZxXgc2BwxStmDQWc7vDy
32rc5/7zMr/5WQ2Tg4n34dwMzOzr3SfUl97Dx/dvQMxibskJssqfCurDvrqW8eAim5EBpr5lJ0k1
L5LamQ15KT1x7r7EsQ9898+/P+C8oxqXDWkT955sriImit0bt9uuGmRDamc6+otyZmnioCCknRDq
KzybwaJwwATP4OtzF+3Nx1FS2ztgJESzR4g7qasp39uS+CcT/jxXi87//bYDqlkOOGioky9yhvz0
VMjDyXOGqQpcIpRdh7adbtcbSHB3uC/35JTCi7CWuFSNPXrxzDkM+9N2xf7E2q+//ILbpgKlTm8i
p1+7vt0MQ3tmxFlSqCqEwbeV7GgGm+2UaGZYpfQrP6PFbnZ+jn0p4XqEAjVJFo57FHjSfiNFGqN8
tREY4CD27QH336yboPASjtc3py8X/zm8+5Kbtx/l7/q3SmOxqT/DxBQE/Kk4Ead8PRE70rQ2Z+am
o2ztMyGTjGCQoWYY8C5ldTyl2kezPx9B4ObXcQjjgGYcswtT1MOxkPjwZ89wOnCGn+RB6uROeoNc
bNF3oBBCVvxnNLNWex/mT5LCo563MwN2lafof9G3sdBFCsgpzdH80AG7QKCvOBJgoMUz/rg1WuTL
Cf2uG0uc/SBuSUsUlF2iF3IAd5VWIpBnEcRWiu8DdMnEeNO8BLMwPEpKDAkHOArzjPg9ygQ5X/Ue
7RnlON32qW3tg/vETym1yrXf24QG+J+jPHsRf0ZaDJJGMa8ou6ZASUGpRFTnWitrrw9bvKYWt2OQ
l/C2SpcON/ex+ojMbxgGhUxcemCOs/nwM0ffVAm2S/MRmEalc3pbikomHY33hEe5v117Dw459hDH
zBjvQan/xzeQPgWyvMRS5ZCT3Rq7jnbyAwHGARla1Umzq4hRDnqkWbAsJufTjvHAnRMNH46KemDX
uzoTOX5erPrartsR63yqi7rX9TKVIt1ChE8/1RDNQbPDyLgEEojJlEzXeBY4aa2qXvUkINrMl7ic
Mc3XdrV8xq1NggIT7DueXzYqa2S20/RFxdgKZ6pNAL8LhHe4j41og8BjYHqd0Uo5UtycjkCfPUpn
8cJv16M7KcR6CLPe5X0hURCPRcmtxTNocmkuxEnC+EeZHE+A8JEFj0/ryB6ARWtGRK/JQeHVd7MM
lBy9obSFybRg/BFwpKlP118+U2u8I82sgmGI8Mn8mxDaoVnYivPuDrySkwBNhglVSVqPyQSmvzf6
7LjXmxmpHlhrU4ARuNG0HY1wlbqAGvMpQVy9W1DWbLJbaGNjA0F+lZPzjid0j61ZzOPTbKB2f+Q+
PsYsBy1lr5jtCxX+f7mGWij4pDCUiEI1uJvHKnqUosk5ZlXtFR/pQDS6jaDmhns5k9/fi3hN5nJF
XP8GksUtpygI72q0ppkQPhwqErkDu+CDL1FbenhkCrqPGgC1iee/FqJg5KkIULPxHwnAp47Bs5/2
yuzxRQ+7n+0GbJ38EpvWTpTXJLnq/74Z9dbGNOmoKDkyfca9wxQ79rG3FtIGNIrZlrmeiE5FiWFt
nn0cnqJPSUi2lzSPI3ic6BahnRWcEL8hv3eGyhKLSyTeN/f5VEfWf+l+6B+ohKEKbB8j3ht6WVF0
BCfL5yUbT+cDKFy9Kr4gGYlYo+w5VRqpDTCMAG0aFrQZtHfQbFUPbANmGaIfHnOEdQrgMFt5juMa
My4vExd3y3KN11KvT4RWPn0KoswgJnIpaSafuijP+Ek54KmBGoOwoe5c5LdoE5VtbmA6xzAaOKW4
6cx5emKlC9IAPLNJEC3xAUULUCP2iPMZq1JlIUYj8gaiCc36ua7xrAJSlxW/9sJQ4C7fxHdEyyKh
VWa8j2dVH9hztkOhomFyHAOVUQU4cnx7HEJHhF6biJeHpg5yKqxknN9bKRjJzNZLNLGAUF8jgafF
c96RRQKTLI3jqwZz16Gnn+qGEsjYoMfT9FvKPLPJNW1cbXMNuYjs5VaW7x/M+n9PFu4umO4rvs8y
rfjAVSHWbAWFvz/HkZZ3d9X5EMWqwJ9pBdzxF7a8hTtmKqXh1IpjKJKntKKPr1NU0pee1SMWdBnf
7lWQGVFzb0nTBSJaUoMOO5VhvqM27ZAZwGWeoSsC1taW8Z/msrnIgClwK9RakrgA6+FoE7JsZQ4o
jOqeD7MU0+RYZZ+c26ZroYb2Y6Rjsw8fdQlJF9W+i/hfaJN0QL0IMZyihYjdtXPe+fF60tt1K2k6
ik/srEb9LyntupGjBgc0OwFOTF5N9Iku6aacfUTdueIuhOaPKbf1oZ1lKtMKrwUzFkthQAmgHE1b
m4uyCQ9zfRas0h++xRnvNpdnU+oo5+HCGB/b81sDc7H6fLpB2ZxwVf9c1NHkqPin4JzbmiLCYwwK
f34JmHg8rtSvJDGKSXTDG6cHGUaCAfF7lTtBHMYzysBLa6n4tRvkuQG1xxokeOpgJjZtPLHeLp6i
Xool2c4NhRwU1F+npJObMSRC+fydhHMYLSu3E6T3dY9TY80698Go96uIOexv5hhd5AeaSJL4TwFv
ak0YjGFGMCrpmSaNwKJIzp6axqjy0sINmTaudwoolNTHr8J05V6cGvr2dxUtvC96Z2ABx6fBDmWw
l0JJ3Jx3peDfmKUlHkDOUs2V71zDNpeoWqw9+r2Y9gSLRpeQ5jm3ITkZqaHr6AMWrAnLrRzinsEa
0QV/ppJ8QNww4lkXucXvLt8/Y8tR0RtOA6SaAIkWehPM5jlrQVz3SznNHP9TDLjhyZBZdEma3K6S
fWnPeB7hnte0lUBEDHKTl2jFrux5PjNVCkJ+DOa+Ep/gJkK7tSzc73I6PzWAARZOvGc+u2SJGKB4
fgaJdshlG8hoxSGmNDk/ZeNKYCyVk6CyqZJS0HMeEKjkVuHxV5BJIIZn0dSvYxhre8iMyOLleAn9
do+EdMaoQARTi1wd304hdl2vGW/OHhLDeI7diX13MH+pPAGvz+Sa2Md5NUf+E14i9rq40IvbUn6H
6ubqlfQNqssCxFtzZdjPvdBj2/dIb4qj72XVgRELhixtirtOWsZimJVT2IPQvA3uPXgOFA2jM0gZ
aTB/y9YJj7dNYPSOwjv4+Uj4Ej+BUYSYmAkoGyABs4JUjYSHpHxJAKivkosie698Qb2asEzvGdfY
YnFXGSVAGwOWKPUMiLZ/BsJgx8br+dgONHXe/07Qr4XKOa5YPHeX+AQFPMG29XdYDj6wcFHYq0v1
STpD0ibq0p8PQzxAXPnCV1oAW6bzGO3qkZzhM8PtpmF0WfC80iVsEhzVJxqlOmILgL6uS2CkmkbJ
Sq9ozqQFNhG8ZyFs9PQHPHon0oJ47MA0VSAKhsI2kPZDGi2/VxiyoJIcWC3Pj28kINcUyBpjNNKK
Of/CncFZfYd07uerPOYCAhgYSFuqrDRBJm+wFQAMDsoKmvh+T6urZKj+wk0QGT3x3HJ39mnLsf0T
MSUFSWzl6owR49OKhM1LMqclnXpo/nyiv5CagRhYzOaqJkOifSS0vNrmCD1gW+ABmsOTbAcUqC2q
MjDDhBLMnHuUslfD/DQfcFBdmwRD9srWFsmFrtChmftVeVHy/gOikZr9tW68k17dnRo9NYDXnnrs
dqqnZlc+eiFv8n6r6ZSYDuMb4gcHmj0wxM/3rkHOpqy51uz0llTEgdRobAjJ1R53lkzQvEcFIStl
ZXWhzDfSmeTdzgGdHIBKmbNwCBrRrHcCjjSvrO5/E7oO59vdvDiq5oRGWd/tDv8Vn2Bwj8XPwdmq
0yJXMY9sGb/VYpDBY5myzE0/JPYCNMpiiy0A1ityMnG8VrFyoZfvzKXkoIclybwCq6uy+HzdIx3o
uYD1NcSXNyjgaW61DlqhAARUZce94yA93BnYg7LzK7HaQqnEy1SGc2cxpkhMsLycUf/wvu0C+da+
jKQZfpTirQN4kEHOS/dupSJQctvJNWJKTY05uFfJRgKPQzTtxWW755dfj816+L2UJ7mFsdt/eNgj
asauYCm0hhpgsrm4TsTHi77NRar5I7dD3P9Z1OFHw3T9xsxgzignxZXqLE1I4WfygUnwfJB0J2Ui
ltvKyD7zMA6S/QTM0zW107UXqz5HIRdE4hsz32hTZZip+iCKglc80o2gDXf9JxOcRZMsckZeG0eu
7mHV+u/vu5zycc/9xVBBuVDcJ1lw7cR8nNvEHrIlr009aL9/Bxxdcs6ZRwhqR4bfcK0fDXWr0ohG
G8HHMy9Iu/fPpYUWv2vs+eXL4Ysks+wQYmIE/zwCahqMprEx0IJRbGamSuzciFbwbVIfsOm85NzM
e7UIYI/DrcorZXOZN97e7r3gp6BHC7faP5XeEjLS/w021d9XyyESts9/Zv3agmtbg3fp63l3b+hs
9CXqXyCr2kO4aUgqTRpbqYhKAkyNlV9K/8x7DC1stXJcf+2m2Rrl9pXUY0hzPx3wv0gSnT+GBA4i
cqwe25etlnP6ddaLOCQZ8kH0OAOcbtXmOSVcuOGDberEV3p5TysO5tnwiig5YvtI1P1eDTmwiNE1
oqMMXwIhck8fykzLxdx9vI2PdVXl7pmP2ybM9taqPCUZM5o+aOl4dGTop7lxKqBUZvQUydIV3G4r
59WjE3VY8ALJLaHGOWV2oRpBRCqjZABMVoaIhHFj7RqFmwCPunimUFI/pgN5uGJLGIWk18E4TjZe
pECw/Y3QXfUSZ2gtWfivpRjpz3I+4Ncxm2A1jw/1PJeWlBAislc31oGQFkgaYIQhl4UVIKH7DVA4
jYsGfDcu5sXYUCuWnCR3faE3pF+8lWUt17rqvhY/BSXmNVLabVNMv82/vNXce1NXNmicj9uwmL34
RXQwISOSQVkh2igP9x1GFaa+HdfoB/wkTaXSdDcWn+A3GhBIKfnKTyeP3WTletwNiy/JyMfS9yAf
KsSw6GII/vNgfVi+b2Zyx6vYQEjOXJEGRyVOGg1aZlwctJRsv4VQtjsNm8PanMOfoL4LOrq4O97N
QwqwZpgZfEuQe+80pVVRQdJsaWQdBMR23NsW+gkJh72zgN+m2KxxuvgWkBpG043A2/aRKUR9Layt
/cjQ59S361JlT9L8sJU0F4eLsoxoly1sFHDzQE4XCXRtv0nY5qT3bAE2hAEsClRpjNMi6gcO7dit
GtcYbeMZqlYwNIjsoymUTiT9V4nW4xetmwjp2GaLYOsMimYCOkEKgX/78EOlffnPrXSUXq6ZL7K0
ltZUp9cakSv2FzOI1/CB9G4DGQtxNKKEm+omtDlSSho+kn+5Ug5SgtqYsGdA7oZ/sCmW43/IQXRT
hXLy/RlN+RGinOXbGZTsFL6yZYBeMzqKvgqLUS+lISuL2s7JlykkXxXe75iJauF8Q6Wn+CO6bIyo
m8Pw/5GI1zPYSU5LCqLaHRkQwiGDaT1ImqIqgHNcFjNWbRC7geMT/8TSQVLscX0cqNl+dadSM0bE
gT/uAFTIbNNNk6Anp0oxJy+GOdr5TCYp3NmX1nxTRWOFgZwijlLj8glWjPVno2l8HX3xmDW+vppd
rj4VVLDmJb8OS2dGqshtAjXS3nQ8cPJWadggciMJnljpTiEhA9fEoJkQnIycUon75rfm6NBIWODv
a4cp1PRI2vKA2z5eJcWTxg8n1R0Z7SMUvpMq8YqA++TJP1iquNY82VS1e0ptJazCMQXdVZ9aDa3q
f8RYXp8Gm/it7AElDhQd379M44HTkNoVBEkFaj+RDzZX+8dL8Jk/QI4O1sbuhkhtSRvHjA6Sk61o
XCT/NHWQ7KVSiPk/1+FSVjjanToLKCNLtcMf60V/neDnwWScpQOvRFPJLkHT3bRIfPRXng4r04Bo
g2Me5mFsn7cKtwdGPQf7J9PqmjT+5x6JhjV7bVh5rgcqjf7LNg3YGcKJocuvwInNDkOB7G3hKhoK
5O4VDfbrC/TYcB3UXIpdsWqNFXBttL08i5aNIU3TUmyQObm5mVVNtpVDOaAcUjwyONm/wJPH6AGg
mHclOlsAI/bCc/LGA3oOx+7+CIQwoBE4dhCfwddvmsJFa1bx6RYc+GGKAeGqcXt+HfglbBHoxaD8
w9T7WbJyzmGe9x+C5XrIm1rAjxWlIhMlDw5AI3Zx2cQ00MWhjwit0BKQVTCNWJe6IWPbHjNU4Kff
SHxVKtJHZdeYyUuLQe72d3sL7Z7M/M8zqcYI8ks9lWIINDaU9LoC0/lhJIW/hDAUARSfS2J8Ug80
2FSFDGYS8ts1sPDnAzVxNStea9PRJc1loV2L6gk1AePyPXyrfuMCquJ8AwJ6nZS79hgoGrjI02vZ
jowYU273lXSY31jkWLjA4kS1DCYHLUGswpyegh6bcrjv3nmlm0ZrMk1IF/83ixf9GKHa5pPVhDHR
+5f++bVkvu4QPB0AWy2Fx+GfIeulayrmv6gutbx0YaGZst4l7cloFVc8Chb4ijDI0nOtVQKfVxaP
WgSnM8mALmd+EVeYt5DrhjJilwb40Eq0SIgwVz7oImVqTagLUWgabXKMeF6iRnv/M/yMyImLq+ER
Ymqfq5vtSKV+VkGy5JRQt/loaLHaXMdCC+ctz2EO83drucW15U612SZvM3qXj91YOlhYCbQzgokY
71ZNRWBSaZr5PYVVcGdFUrV9AeFoGikH99cNzkNf4PzXwxypyBEkeQ9hojRrR0dfd3w7be61rxVc
FxSbHqDvD0UJMHvkI/Sq2WCi5GixsFCHKoXjESldDfLIt3iXrtBjPoMaNZm2vLanOifNxnA8HyaI
neZChjbzUpWBxvDfOpWCFcTax16SiFaCNP85FerFdlo0jhFtp652acjsyx74gnKvBlHwRe8VzFZ7
FZnHi+FfqOqPSi5NB50Qk6lf1Ak72Lu6vXqB8qNn2XNSrcwor+MhismSfblnKJcNvnTG2D4YjCOE
U9b9DVs2XV9ELFB3G+KzqKts+2r0GIPdyIl6C4yYsGrtxuySd8pEvpxn54Yt9GTkzHu8Pw8xRPdF
fuVXvOQKHaoucjTjFMTB6li+dnaqyAONdLETxtEr/nrQjS/aHhML7mE2D96uj+WQgaW+XFns491O
D//G/2vJjfLzcs8EYQdN3h46BBiwZo+Ctp50A8KcSmdFiyivCH1MKo1Xg61fSEjH2Qcfv524ELVQ
hFlIw+AGESzIeYB+N1Ut80AKFUeBLbR7hLeIE45dwbnTcMl3egHg0xWv2thXoOTfu3my+BU+imdR
2vASZApv/fO/TOMBkeXgnEU+ERrD70uv1aB+KAI2vO1BdGRXpW1lRQdMl4JfHCtpnBmVi5ktzY4X
iFciQOhn8P8RGL9eqNHcmvTuYQPbxqlyfz4IFA2vEhpCHdJAPeFGN5hY4ZH0Sa5IxhyOC+qItLhV
82u7Uy2HKMHhnusce6OxRdHvr2YDqIxN0GVaSaCuvX96bXec0bnIbQvkg2qdVMQOn7pSJsIWEMjb
xOLVaZK+5HtvULu2JPMt34vZ5JWb4OhTEdnIrWiQnvOCIfvA0oUWmxkJhBEnHK8fTE4ftAgmyH3b
jWTvoyiVEzAYL/C94mA+yshgav2iSUGjHtD4hC8u71zefkZ5nHF1W05qohfXIWbdS3vQ8HsY0k3P
iQ6k4Vrut1nAdoepd+BlzklL/x5bfyGvs8kmRBTHVNGob7gN+2wSf8ys1EaKFUxMCo83vlP7y/GV
9p071jPTppYpvY56QT2brfaSxIuQ/ZRRhlrveXCUGx14+pPdAyi3gxCdWgkBmqyJCWid/dFnjVgG
J41XnzLhJ8vOtNubHA4RE3F2MkhalDOCbTS78vqP9r/hQFhgOCJIrgbU4Y8wooUlnr6sAr+w5rDJ
cn2hgab33UR+kk7Y8GcBihQf5v4j3YnCiKKXiW7C9Y8uDh9I70Q6N67MF114v3++0AzBFT+pzKF2
3Kh8V+cdi+cjjD024gwQ8Zlbgem0vruj3M39KO6LuXrGI7ICdbewHuAh0HIBrjmF3hrljYoiM68D
aedzvP241kWFmC5+NPchzkBXI+yseUHFFN/x44ukYstS7CJfu6JnppxFbcnL6yjDa2E/6a2hLtm+
dTpc5mgB9dStFWVb2suQB6jF2GKRmyYemYs+yTj7f0DJwp2NqYqOOKb0QSZ7zHED+AUNdOXgz5eP
w60e9g4znbkgNAJRTWTylr0O9MwRWfpYUgoZMAeSJbJ5CcGYKPGtHvTFMXTaxc+TCGnd515DHuLs
SxUHB1dSimpsQQxH06z9GPs8ig5jVAg6wRcKCfKjlLjVSJ1KLfGP5xjvuZOHeqli2E4814UjdxkU
849x2tRH9SiW1cvbiTp4fmunE5Kc1YLAlSo9wTEV89gL8vF8UylZHvjCf5jiPXAnOcW8T8XvvEXL
7L2sTANIIF6bWc8bgiNbLqvF7i82dmmnsYiKWkoG3eyGRHxtLr1nnqUv4QH+Tib6gQvVdWLmHhBf
RZpd+j2mh7xgRmIYWddXX1rOZ//udiEWZ5KGCRlukPMCGDxn15Z5/6A3Z/7iXaW+cGHJ7hewMx8h
ZGPoImWQaOFem+9675n3AEdV7XrtzpN6TKgFTQmqAKgXbkx/S7R7t7plyZSYad2GoWCOEbktsweb
Q1T117DapLbO4UOS0FU5DQiu1tN2f6Y+TsHVpEMC0ZfSgw0tujqcSW198J4GzwqUry1c/sk8E6sh
HwAhjT05KPmhHsvj4GFfjMK9gY1uCXpz6nkqiDahfBwDEczW+D6/A0shehHO1MqY+2SJEuWQBz18
fWHjDMjyMFC1lgGoRG/Evclk+QCqS8aqZMSqHoPO7e/fBW4rIGt78ho+gQ8yCnjOLwVUyQjFehel
jO7dfc3hFynMe8cAD0stWSiOSu4NNCPs+MpRXMepTRbkZPKVFjAqUn+pNmj+UnSaVuUnn+p6WHvc
a6dVMIiyVi9Rq7mn0ECKRMsQJDxdCG9hqxiNzGffXFpq6ef2cTaLrExiGDn1wLlWTCDO9kxiOYMg
TdWgrmU2y/v4lA6I7D2342b+50eBORz0VCEAbG+O8DVk/pQK38Ck8AyIGhsu2vjmJjZWIJjINUAd
QFCTL4E4EK2c15X1X5+h7O2+g6zuUqR2X+4hSivshol4ew3CKxKFeQI7PkTJSzENGSg6iCa8CvUz
LoRngZIqhCbq8NojYu25/LSNLSnk2W4EZc9cn5xMK41IKc3pmEufnw3Pa5KWxEqyIMRJMe9gV99D
bjbHRPmuzV8rAqA+GN+9EXugkIQnJVLTJfIAg3+/WDY7eyvcQLGNhfmELXB4ZAohtNMJoTww8u+O
RkDLkSx5VQuomxSthmAybFEUmFP5lKO1AgeWWCFoedtCZC+O9SLHnOY08b/umiQUFo6yE0Z8DZBK
QcxGlVNfF7DDbdtNFXE6BMeETcyQK/PFVkKWqvJL+ZSss8fkA9ch1F92Uq9lvW8f5k2gtRsWaiae
h9wzczyq+yTPqMTDEJwzogyPzhOGl6OWPNe/UsBuQv3rtTDVm/biegdmqqZAta762J+URVzG6zii
h9U0bxT8aJ+37OYsD40KyU9CVQnCzBIE7peBrawT5ouGUYqpA1XefIDP5M7zspeQxf1Kwbt9wjxj
TFxS3xdIKOnCtc5R9zdWGiGA5OvlX/0KV9hfFqd1IPzf+tGd/1qgicNbwwP826+GerKhrpgVd9jz
h1PtBw6Es49XloRnrDocLcSJ6LweuArx5B2Y7YGDXOTc47kKisvR52m3AbFi8/rS0emgcUzJulU7
7zSDmfbp4X8ngJrGunLSBq4gcnet+j7Ll+IkyZAjNj6ykzspQwZzXo22f9xNISkhtx4aEzyYk/Fv
IbPo3YmAmdMtzH02rLacKRkNjqP+O87hB7bHWY7J8sJGBi+Czi0BVwO3LNpMzAnrsxrKdqvPVpWq
x/gUayNbxUKaScw9wlkeTi42z9kmBuvEjIVm52wqJ5lBfk8j5XmVhzcIjACYACYMQ4HMHJNk6CyC
YTPG1avfyHb987YrzaVe9An5AVd/oq42Gz0yjckzWi8CwCtnMMfK6uKgbL/6jAMKaWsP2IPBDwML
zSBKyREwarI/s/lS7vC9UT9t6yOGRn1PNwi/W3GGBXBS2n+U3vAlLTXLWX8W4pgz5KFrpBBZHThp
HmXFM/h3CCug9ZJcIxt+wtlmTrnLuPfuuItIhdGKHvBrGQBjht7UaW1mNEd0Sol5PeFjAGwHSF4m
ECcCb7LrHaCwCOTff5K7FqRxtGe1qzK819+ZlhmDs0pVB9scNBK/jOu6xWF3A7atkBYbLLTV0nzh
GJhbrmO5EFC+kfdDaFXme4DC2N3DcZl0zFMfe+NxShNu4EGxPhDioyQKQkIA6HX7deCVpE+HTC7y
rZPkqJEQWki7QMSSmO6mBMw+I5trp9y4zBVUntkQhYGR0HAUjjt4A61hHCx1+xz2oYw0eGuHolN4
uXIHqVibs6z8wVUeeSO/hiYEoGbtBP0h5VCTXP3BPu92572IoumKu4bFaatDS9Rq7poJ7KP9VkOU
HZGjeHPlqmyR3tAzi5gnowg6Naepel7TC81pUrSuLcJcoT5oPGe5safwoAjJv+Mx+iBCXzqL0aGO
qsRzVoxzd0SH42OQs+eCAjmxe7pRw+my70sL88kBrMge0y6kVGdC1t769chgE5MB/91SKutznCpm
1adWG4ekPsSFiqBsax64Rlc+OJ3/NWxHiBlXwI7D0NBIYmIjJfPEAy3z+3PzWm6A7MWCVtWK1XVe
A9Rj8gqb1Qi0hfsFXV8Ty/jgvGfZFTvPM9tMwUI1VDhSbmjS/oeM2hdGfyBAVDWKX8TYgBdGeaFt
CLjJs93seaaX5vpDJZ+7lvP/f7IMp3ydTYWQsY7AmgsuLVwBNi0PEmjZ4K3392brnCg6eSX2C0ua
+v7Qbk+FUyziGB+cUzDrSDD5Tvp64kID7ynQZxrnO7acsFKNGBh2bjtJtDgFKWAvGeKzoXTF8Xn6
LlXX9iBTIdyFu/S1IQ4x81W+dI233WJlqMb5CPwLDt19q6HND2Ha8RNuXPIJgzNoUd8a59HSFFGd
KuzRkDFdtopPd88OAUIf4tqNL2oQ9n8RTj82iXFECrrGIeJZYvNJ2wur9TndJm0pKG+OVdggac08
25AlfDa/WR+tHNAvF4qkCPVaEVUQhgdeMorgjD6g7hhWj7PsbokVEFzPb9r0CG93vP65oY2x59df
SMoL7b1Yojv/2S7G9FQrc2BJMsGDpY72CKOb2TjsM99OGZevju3Ml6NohAHirFJbjTAc7GJiBrgT
SPAMlHRjpzrgzwEfGZs4xr5Rxmkdr+YXWLGMQGpnJcNtB8rAVge6GTcr7EDFvErOtU4q0f/l0XhG
2HS+adX367j09KF3vAg8rL3kS7l5VACq0C09ppzOXJ1bT5aU/DpFr3TNDH9eBbTRhJLEbjATLETh
eGm51oSdztZ+JH8Z48DURXjFOiq1sw+epobLTtrAiKVtIU6TaudgmVeO+tpmU4N21SEJ1YhYiXAE
oNaDGvWIqdRnLtMoOLMQ9PbDwFZ6ELa0T00++IYCNfLOns4VaV+pH9xDsmkm6ARMF/eCWlGOSKMu
ViDlc55HzcWYf+9D+5z/lYlhOWBHnrW+SBFYAJh5Ml3wvSHGC4hDocjp1qPk9hvsdN+C5uO9qJeP
V6ddmfyPui1/Sl0ilz37Ch1XEA2C695zIKgRmW0iBSBXnatu4QFfk57xF7jLJBYXHJT2Jt4gLaq/
O49ZhLDlcsbX0tx72ERFAQYoFV9Nhy1u+6PBZozaTp+JwKvSlr9b+k55vnMKLWtJ7QYBOtueHk7J
87ycE0ZGLim0VfJdHE+3pfmO1zuIv19ep1axoFHs/J2g55tNmf9SEiJELihmfh2aXBE4MgjU1M/e
u+hoQrJO66k8aSxCY4FPDTf6V5o43jHR2tAyuMCHtuF4ZQwJvpGuVOXRcavJ9BYyUuSIrHax3UuN
Z2t02+BQBwJKOW6iFQbYiVFDYcWaSnOpq8JKpzFLFeeki3T1MRUG3rAoVz0V14Bkj5JujbTsdt48
8yoLUD3Wg82oeTkwDJ/XMEMd5A47j4iauUqz8YZdsuxW6xmc/8RlFhPkvPO6TTE/XDM6NFlcSeSS
XQmAk4c3blnz4ACaTDx8RSU3kaIrEz/6Qb9isj7zH6tGM3rV7iuCbgl+PQtQbXOw4wTF6ZvgM9Ig
EKgokSSMhy19R0IerF16u8EVCpSKxyGBf9M1WqwoaIYpFggkI07uTHefqGXybrnGzrXEvtdaXFsw
oF2N60YWbF3ZaFHaq/7SzZVpqllHFtzTyuSR9M7Jlg12kJfEIlHlKBFH6RwspXUVBbxdwEnqcv93
IPtSGVkj4IfgbfyZLI0ls4zSVVUhdDOn4Se5t2pXcAIa1ENA3OyqS9Q51+q3scK/cRcFTZ+S3nRJ
nfYGfY5oyeim/IVL8bSvyeudSED4jTznllCyhbmfyLO4JG/WD4RwdDFIlmTHIjKKl0eiUyHouC2Z
EbAtoPY1kqRkNimOnzA/a2Rud9+DjpXbhfcYPdAXR+w1zGib1YhE1/dBekWXjDLesHOrYjAM3YQG
wmtOaoRLkynM4ybk57oziEep7E/2tMo5rVY9Jue912VJuI3bU69YYqgXbhY8LWxBQgEvHBfsqUQM
gvc7+Nf3FHawfuqHexa0Ceuu/FLme4hej9jYQaNjDdQAQkOrhnd3gNZsgKVo+Hb/S5/goauGhMGP
fjISnZqQKE4oCunEBBgOB4TSkgeRmYPr38Tr+ebXGfuBp7KwGHRzQ6CCQ1wXyLPP5D2/nNRWO87e
RdRDAr+FEvI5zYHKdtRDVRCbV87VdrYuu2abnYirW7oSY8F3grnVObj69L1LW3de8mKcAPfroF89
1xGBWeBYcOITngbXNDDX3XXnfDP0dCE9vqwmZmQWV+VadLIByuFK6H8aBSzwHo8JvB1LiPIo2+Wj
Nu26Mlbe1Zz1BiMJ8238uTAzsV2DdC9UxAY1OteHCiY4eqdQ6ZSSUXTSCcgWPlJ4vN1lmouQg5lQ
u2yF6nQmUnbEJ8GCRAkX7jHpMT1k5QwJxhhHgBcvi6NVye2dAsCwQUSrsLd89Mtdf0ytdPhl0+AH
9J3aXc1PXPpaS82pzwbkWXlq6ev9gBlGpY2+P1vBfYiA7RNEVZrcUqHJtNW86VibAQaQSk5vjDFx
jcqy1eTHLPgp2sJPOD4ZnMfZeIAnNQXXBFHN8OrbHbI/STFBctLypWVJBu+56SGw/RydlwNyeIqt
jF+bdOMHFwj8JA/eA1Wv6F9LWyduEj/EUzYnGaRAPhf6lVGi3/M9YRy59QhlI/lUi9H3W9dL035T
ArCu2DFdQMnSAJniEj2U18fctBDQAcZMFaMlVifLfqa8ji/KkMPOVIof469OVhI5uz9c36H7WfVC
N6n56zAs01ML7s2yfNxerrZMwLCHZy8iXyAlMjbZIleBgaNGsb4JcUcZz02pbpxU4hz2OtNvNw8T
CBSwuPe2QaKamLV55Y8ZrqV8w/p7h2Qeh/EBqpaCwmV3i4YFeqekNNTLpTu5Xdj2juRO8xJTERs9
Jh7Xwxv2U/pDRTuqPy6iUz7TPXPA3PDZJBgRsAuP9EK1t5FNOxipowYv3gAG8vkxoPidzLyZzQpY
5hnJbHKEZsviqdCWBCpsOv8PpjxtdG7LCoxj6Di22TiNw4gdys8Z/wdGkZFam50vr4+zweBEFloN
NnDq1ZW3z1NVV3Nc9fQOozdw4l3LRRqv6aKeylsJq0oKZWX5WHh9ZKgrmimLBXenR+UodGCs+ShJ
GS1q/FFX9ARvXhLjTtFhI2CzYA1q6XvVpvry5ug53JQLbn5ULGSh/6bG1xSsrM7CHWzjXeUWt1FR
NUqYHGhefcQecynce7+ukv+5SVlgRrgbWV4XhMS6wjrME6idbkrSP4a8KIb5vYHOmSMdzsLCtJXv
9NvBj8dt9AkfDIIuxQurCqt/+ldlXFPUQyh2+3i0GrU7apcYylkfT9WUxqr249aYRdvDo3qk3KqT
025KvAgCwa7BNH5p3M9KowL7FyD0Z9Sk8mKdAMa8xCDSc447LjCMZlqOBymYNsT3UgBUebxRgELQ
JOfLjuPHJyH91TVZHdKdIu2ucdpWwetcn/g+KC0IR30i9V8BXnTc99E2klUsjkzywZ728Hzeo6e9
rjvY6mB4+QQ2ZNtfgRmx/bDtm4EF7A0ydCUJrbjHoZaSnGVaSz44wkpQccCifjFuToTzoGe0lJwy
/nBYKB6fu/LWX2QeO5KPy0k7q57w5fecSueOT1Oh0ytMonS+Q3Pg+z+aUQ4Kjyx2fiN7mOoFA9Mr
30/LmoCkq/QDK2m5S1cbPfnDoSu+13/NK6aM7y4WzZXjHu1mrirpPfwiNh5cEuz4wqiE+9eMW2n0
HcJuGcoTSk/zmfVuhJH/6eRRgf4crvPjObKhyN1TAKJciqi8304lp8h0Iqxl8XD4x+12WmybLOnp
PCJX3NgqQXDzrEzMTnVmftWn+9RbJLJkYfJfpQO43VDsqT9WbRegmyzkbIIlrtGghT6Wcp3Ti7B/
TyykhjIgONGSkFVaosXaD6kcA74pI5j3YTM/rJ+TZt1rygrkglrZnhkDcP3NUrhpSn+6HxMSBVlG
K0dFv+kjnWZbzybdkQVc6a3bY2HRguedgujmHNbdjzXNAJ1optEZSH9RqBDSlUtY14R2Mocurmi8
eEX7BUZyWN8JffWw7hkJVRIanbExjwGVsZUOyvAmtY0EUptGAiLUr4t28VbsbU/gwjAduNOkUFlR
D6R/SbNMXySLXFgi9ni/Qy7YWvZmk3V1NCtfDYSCpHJrpHVqDn2PTlEUb2eWA7FfPuiuRGUPKxWK
hW4/z7HDWygpOwfQcP8GQxTEMVVwR81X5Ao1Nkpi4iba0ctjNzJDY7XSWigUlnZuhA1XSw/Inx7w
E+rJ1gdo307gPV3knUaMhmNZZbYZXouoQKJGVu9ALAYqKzrQgGYfgQ5wCllxGuLF561RL1hB56km
/FfsVvb8Sc6rEfXkI0LwnFM8BHj++HDtKK7v/6sWMHTlCW12Vp4LKCTcNqIry4CLY8OiDj8o5giW
8m6Wds3QDNXRaqqneSWhEP021M+25X/Vetss9IcZ2zIClMEwBSOC38eXUgUDXgYlEmmsU5KesvyA
nvObWG1e+SEnWSMLiQRheRe7F+cfmfkIgKIttDAPi1siI2sD973LiEp76xkkCwCbefXKLzKF5UnD
mDyTEw/5Tmz1oqPc5Yy9fKakllop4zE1uJ413Pf2eUf5RHE3k/o/qSNKlyWS9ih5PB9meUjBorit
5r2mpOoapseS3yunLTAHv8DeQ48FXDVrlkyaYEOhKsm9+C/RN5jHDBsl6qavvqFRco0YR8xWsTUS
6kJPZxS2Xe3cZcQHEB7uOjRrdEkG51BwdozWbIVhofelFFDO02GyuRvFSwXRdJAOZLjNmaAGEMMI
0qTfoRIH/7KPbwhpNsc/fQCQUWHGuJD7vtCi8bwohoz2KMtfoEW5wOT9Jo81+XJiS88xybQON8oh
Zko+Mn22Mgtu94bPVdNDc+9H2+wGmHmGC3L5jYR3vKWrcmZm4pKY+5oBs6GwAL8zEP0amPwbbiWp
pWu33kT80W5KznAvQ9XeFluM1v7qrLXg1khCVq/t2jz5mnv+UJO7PgxMfzMyx0V7A82YTbt6ba8N
2zY2Pj6mBps58Esci5qgekCxVIVVHHHgSk+t5GEbSz9vbd8sw9oFNqQnFG1kbHZriM6m5hW7qTDO
WzUFq/Oc7fd5YQa7frJrVvj0fSjPsTZL4WL9xaR3Danw8hniVPiA0P/U9Xirv6UGl7hvVAngRgqA
nWBLePMIB6tM8pdNT7NFvJEiTp/jEqnuOFfgCva1bfyaQexSf9c4Ov6qDoaaAZpalcid3+Gj4hbn
jDMuBHDnIGm9aYeJF2vuEnct5oy2n3YD4VnekMq/uX0PwvuA76Y7VT6zo0fIxvwgj248rZTm1TdZ
prHfnSQysen+uvUvAEKJQ4qSk3Mw4o3R0jHKQADlRD+xcBxmsfiE9L3q4NpEJit0TqY1eqk/FMcE
tSZPKWeIRwJc1NPagB23Z5DK2W/rlyDeOiaFqIZuDYmYCCRooNvLKSr4mRegqI1FpuEh2Ylq6PUn
BhROHF6lnQ9HXPHkWxO23m/74XxToZ/o0JyZVVfoZVPw4jP/lmGCawFPHeDWLcrRm1f891+89T99
NLmqmoTclL023Jta6+MYx07f9nUH078Rf+HgoTxRc7QFUYjOuKPyKgyyNc0Uc2kSC8Rq5+OS1HK/
Aktp4j72nnXTkS8rNqebosWrj57qvGdHHXWMepzU/9qp7mfpkRoW3AmplsyVtquVNspfXN3Nyvzl
mW3iZR6zcDUVI2p3KXXrtqhLC7on/4GI8HKNOUoQaA9KuRkP73cRDT09VWKvSrTTQOXEcxcWjqGW
HH9SlYkpciFBIcn4tUyABQB0YmYOeBf1Fo8B+cZU3CauBQgWrybrBi5A3Mj/2uPQiiUmdJ5Xl/pl
YHNzQppZLvMF8Gyj5GaFuHx6zIiwow4BymkObWoJaITxJ4hm5jGCebdCZQ7/VmqbKoxyFQ90EGkg
uGgGmbrYJZ8c3Q0YKEPsx91ywKGTpQ1jC74h/KfYTf6HLWEgAA2l+Pfzugc+m6dAlK0nrI9rX+uv
CyCUVpAK/teQNiin9CrFV/7dstagJ7wy88sVP6TxE/f0F5iQ6nH93+5f5KehBUDiZSKIEhiakaBt
DqraHbpIKJNzD/jU3DiNdnasGP1WoKIgEbiD2UGAYOsTz7vrKzaByTdTh9SiR0pnyyVzVekinDKR
QEcbCtlvyU6I8MyUz0FNn7XYh0lAEN4obDNnGvnvkiV3aFUaN4QhCBqi3F4Q6M1jsrsQJY9CIUOh
Htd3CIPEkLeve9uQudlIX5xTCgLFR0j0v11AYKzQxNT6GL2DbL9bDiVVy1mnKBSPJNwW/bbyAqbS
4mHwQo321Vl4PJTBDyuGTCCa1TIdVl5zzuOAJZyildHPRp7c9DobNRDQKe0rLyZDY+VMqN2Ux9CV
ea0gQfJ87QcCY++0jsTmXUfpjfSz7NL+sVkg9VsZ28dphoLk94gCkc4Itxch0ySs8v4NdTMn/S6W
5ruY7dxdNohOBXrDx8mK8JNkfnzeDR87EkGC8VAjBW/mwHR7ZsMcUoJUfpc2OGYsEhg67Sh60Gd5
ukL4Ds7Xjx54tck7SStz8fZTA7GGShnFj78J4mO0u3xXs9+QFkv2toj9twU6+4kjMu6I30xm92u3
4LCl2o5qd5z1ATU8Wa3DLo26y4OvxNdN0Eq+3sEfnHGsle6Xmz8Cw7jlduF9aoQ+hSnr1wgwq3XV
LtLeTz/g0j9dJMt1/4X//T6WvNEsC1YgcrHaGOyzPz4IjdOUFeicMCy8Df0Bhz7U8q2jZA1ZOj3S
hPGciJnrMhdyKIr/jDGjgxxF8Cn317siX/QxYIEWAjWzzyh1TbXnbMgLL7nN9T76jwCsgAthRE2i
uAsVGlgDIzslhwK71eIItqENxnIrcomsdJRiitmvr1aWmlK3ErAS1L4r6vqeeTxB0qX81NDrl4/p
vPM2PpDzRpXsPyKJ5H/JgtnWoypEnAaTM56EekqTe6/IzdPYTOzwDRk4LWd8ivDYMpbI/Wf/SqTU
T7QLhRXMN2gdgP+XP38QfBsXUGPWfL/1FQNu4gghDgrBzTBdAHzIcKfle4sR4jl0urMpJGgXbAI7
fuJGoWJPxqc/Vsk+KFxQhkmykm6sOFQ2TC/vFgeSQgyUEH5OF2uBARCkdznbXG0YsUMtDu+CnEQo
aeeJ/IdDz5xmgQUFwmyGsj1ebYHfz3ehuwb3u/aacKkwbbCNaXp/k+F0AlyExiqaXr026c9odiyZ
135lLc8Cc/Eujube0Sjou4CWzesXFDKXndJwneHLrwBLGMY4Q3mjfcVwlpj1tDIo/H8j/ey/8e3Z
vnNISTNdnWkQavYwpsiHtHMdWDZ2zgW6fMqvDim31Ck5C0VSe08Op4GNFo5wW1HKKqucNvPIVJH3
7xoLUzN2KSoeKS6xhy06T1k/lYgWLfQF/eVZFVnTK/oeFeOzLOgMVZa/Kdpi1Xdq9GCr0oj3BqZL
rYavRVFyCc4FC30z811P2UKzns1i2eR7O+/chxWhoJ4n0qZcFs0bXZzwUpUcNz3jnVdQeMTw2kNW
wtMQ1Hd4umKr2FZXyTBpw538Dp8LhgdYf8uDavs4U05CHlzMgY/o3OkQ6KC33ejoA7EM7Vje5faY
Hv0BVn3O1U5B/GNSnQLI15oy0aIVD22DWlOVTus0ef9tCIfVm5jF9i7TSvKEupYUCgXTtalr8Vcd
XRW9GZz94xz0AL4rTO+08GL03arXW3XgaRD5j/6OZHzgSqRWj6oLyjqQJsVljTJ3Fzhsn9sVEe+G
vaU8wtMsmcrVTUTAtHqCvqTtHYDAB+rCp0dlAwZJlZADulo+iuR/WSu2MNF+sihnEMs58nQXqcAo
UrEmZSAxuHrmak/9Jfi+qUoz/o6dZV+xWGYOdGMXArJvlWfk/6ccIj/qC1AjdgDcq0LF89wZFpvD
zg+K2dJ200UqG1X029z89xQKVuyAshsG1CDGT9P+mbt//dRQT7uYs2umd0QO0/zfa6eR/u3AsMU3
ukiKTNNP+FHJoYeGE6GxQmshjtmgZNwdF6jWw+r/5cod7VKP1H6NS6D9NO9sNmPwXtDeUi133wjq
SVChdruZcX9bMr6U0B2uCZH6OY3fV2BrynSjv77cVkwRY03vraitR7nOSiyf1fHhRpldrjBbmCv6
1Fj6KJEx5xRtexTjzXBiQYVCDfX18EvbIE5HxxwsnJK2HsEslaWDgAsEJ1jP/3rz1xKdcB07k6sr
5cTVBU6xh8o8VNIG9dgmNoLNdUEA8gFRE9emW7rnHCbZvHYVKqrhQaz7Ek8YLKrVp0MzVP76X1CA
XUEML0UUmH/O6L2T0WX9R5gaRz0TG2WwolsIHBlorPbB4qHReS3ndDwgv81xG0Qtqk+ET0LiqhOc
oV9M1M6jwYhj1cpi+77M0gPZDcsxfTDOOsMQ2TSFhx/w2O19pwwNL4wqTl23ccvz814+jsnl1TRn
KcsQIeRaD4gKO4JMbAQjb02EcrQ3mWvwlihl4SkFGsGMsirli2lSr1QiyQ/CltWregWk/sd7YRrQ
dWB56B/Pjo+nOJ6+++YQTyCqVvE6CS02OarHH+Ips/QBuP5GD+bm/F+4evoM+EV9RYDnXgfFzq2E
2JXBW8ZEn2Axuc+I0dNeEh7JxyC5MiNNstllypE85D9KVQJPDIeQG95e3obOTdzji0M0Y7vIbi6M
w9eC+3n5iGKIoJ46hHlk93aC+K0ELjFwXE1RREFPSrrcDJBOzI/hzqiqWva9jVEjDosQ01KsGXTd
EM61I042radcLgT6b+SvQSm1HxyIdjV0E3JBLRsie8R9BUzDyeT3mvobsKdn2zxEDy16O5U/fWsV
FrwBklUajrERDygq29blDgnBNw1K8xoZ62JpjMgc98sRnMs6w1bTl4aJYL6vofgb23DOVm6Fc48B
R2UkG+bSBMYMgE9UAncyOLgIvfP1n/qhPrz5MG5U3FTJYCbMzp6xwDjuObAqRGGD7+t1QUpIpdMY
FnCH5rAdxpfg9DpEz8qLuMAdRb8ACf2HBb+abG20OleMqdxSPRZ/NkvMTPwndqET35q8dBxBgxFI
CSyeqf8RfJ4K6JRSxYXpWMp0JE0vqBrO0A8F0CDDXC0JvtAcTdXBc9liAMC1SYFJVtB/xVcXhsvU
NaHlPjfJf44DZoGGXr5rYrgHiAHmMC7f+tNIui95ZQMVV8QCMVGkWd5Nmzf97G2ASTWQQwZfTacr
5+rE2jE2F0MiM03BkNh+RncQ+bY/N1Grb7UpeVpyS1zngcVKNHF754jzK3wCW6gGwfXzq1dYMlNo
/sGHs8Rv6UZPlcvv2WoN9eV1BzmxYH4Bo9ZVbIfOWnWQ0+R/WmRwv5WEd+EQHWG5n4W14S3zcghu
2ugDQVAsiFxhTTT1xaXf6XXvU6YNjFJd/W+iLqxDdbde+twafk1s/mOMEaa/beXo4rAOPQEWXkeM
ND+Oxa6rf/MP8DkOyW/jOiba5hoAFi+J+roiA/Fx9Ai/gmlQ/fj5NtoASkj7uZsFEXYvwhyr3zRD
eSQnl1bT9P6OG12+qiyMQ1XBa6tVYqESO1KOllQXRUZJ7GpkzGKUz0AXvdwTWMH8oW4mThREf8bs
Upo9mzY3CngaSNtbxGviPgqmA+IG1r3hzer8jQpMEXkz0FCUgd1Fo9qsrmxHNJIWYoog3PZfjgSe
zzwbhLNhn/QtwgG4uCYco+9ZURrWuRdcgS9FFBaadbeZ/UQ8mxfb5k13wyHCQmtc8gaimbrrJRWp
Tyi8NvIKCtkIANXm2crcS2Jch7WRowFF8FMUwYDnLnWjca+ko/ev/8gbVDT8jjmrGIrkCe+R7Kxf
5UCl9BF+7/SEophtLacYwYmL7WRH1Jeah2Ke51/I1wjqUZdGpAXJGiLswylMcEogJqvJLSRQGEJU
oBUa9B2BkwD3DkL75n1OXq9IxGO/eebSUTZ/daQZSSzX9HTDf+TULLRmNVXakWWJjhet0Ru8bP2j
LXwSMpy2TpR4EwCkswsswJFNQrFItGd5CaZaTNpwMbyQmr4eF+ZVbquBBCI6C22r93hcsAgQrd4f
lQV3ij3h3UNKeL9BJj8lzYcJBFTbGREMgodPxlkfvDQhZwrzETaRDPNsov4uwnBZSxQ+ZQhzmOgy
yqXAN8+rhVVSB3HNMxyhR7wzRFlXeK3PsjXqnCJIb2zBlcU5LiKZuZiL/nd/mPAIpfsAsut+X6rp
txc/oMURjH++lcZoViqHOjKQXi59iSLPyy+c2+y3AjX/jvL0ImlLOfJCJu/vLzypx/vCbicYXBCl
YJlyZwQuO8pau+cBmr6QujSlj+vg1rjAJ2YgiImr1M4cZmqFKEsfrcH9stD85pvr7E8jPw6H+MOu
n4yPs4ajslsfIf/ynQpeHt9X2ZNSh+HzzqNJ/M+aIqexqVVFLD93LRBQeVpIarJNNmH/ZhJyjFND
ws8gY7JxZ29HjFGgwUNnzkPhNHCS1DujNOhofyM30OSsIGMGV/KCBeUtoZhi1jgpIQaIJWqKSce3
KsaRDIcJRZ2QDW+GpN++Ye26HN5gssOlT1urQ5ZbzeS6OjaAY2D7olJf+L/Zh+Hz/l7wl5z9L3II
2IsEPAhVqh0ZL2YXsIuwNcG32otMBNNETg8yPgV/GuoJtYyQIkMKkv8vTTV1cpdECoI0ouipxwYq
/UcYLI3wr/y19v1B94YStAedby1A3PAqbnqoBC1xFmA/2V2km3VG5+mkHldI9/vR7vRLzu3IAuj1
a2zo6APHxv7Nk/FmVGNE+n9jwCmBEyywYH17AhB+F/vvFf7XfnagerFWMduT9axM/4mKOxAz6T4u
P7voC2mgNyS/irHngvvaZa/RL4t0Blq9/fdKeznuDjMVun24+kLGqVkKkNEloicbfPxYLTArdJb/
02Z9O5mgxbSghM0xfvQTtOIU/MUTget69I701xvouBrkWFT5kps8hSdB1aHxYKfVFR+Ac+faXZp1
nsTP0VaVJZnjceclGcTnQuKVTgVXIaD/efrfOZ+oG/Tj/vS2qMoBSOccPM6tFPUG042NJNDatvMm
wVzQA/Ilarl//oclkI/Lh611aphozcACi2QwdmA2tinxWKlsMRs+1ehZMumyh0W814jt4jwRv2IL
KQ1U6LPNXcY/H9kp5WFxKyONkTXY/+hkiQSNTqMR7zP6DPeNirVuUm8+0XdM/M8weDi8TiBJaTf+
PKNpFPnkiYwFSQLNJLJKEpA/ub4Ufh3sXfJr8OODarrq+6a6GrOoRwOPTgY+Kyk1WVZcyXcRVCRm
AoUUbc2y75f7P9LJMDOfLNsJPVtkdP+0UXiqH0cUke7GIICjZwAt9/+OxU8a/QT7reQBpiZRx42+
9MfJnJihVFEaK0bu+bp7iER8mJwRfhaNzJuqyX8G7P1klJ0/FfgHyjt9tZwHK2+nG68u9U5mCmfm
1yWEZWR++GcHArKKUEUQDnnJUuPWhUPlXcaF2+iFE+Di+REaN71ncdvmroBg7JJvUBggYQUgrxXs
X+881w8ZFMI2b8b2+OOPM+7TUA9N3+on43jjuVZd/jOl6WvYri4oEbpN9huUv3YYJiFduEys8nCW
lvGzZX4GJ4YSuY8XIbTJLRxgc5ovlh+ni48YV/cGA6QZSSpegRt7S9vfbV7E4CJvHcfZa0yt6Ihz
WFk/xANIN6CbIVI3MNA1LGFjdSbJW1xyETsXN6mhDIiVK5/bzLYnIJHCUrdqPgg3hYMK5Feb0tpI
urTDH3Si/pze/SpIN1ET2+j1smcmSC7ktcWWwLTR0dz5rhVEl2YqGbE1hYin93aOeQGfv1Pb88Wq
QaAgwgZ1dEwVEEJdiu7secYKafVtorKvb1slwyfKN8yMT8YestyfOVYYiXaulBVffkoxjElUJ1sl
cSdLQk/k9ok6SAp63mguNvc7za7mk7L/ncJPvJvmV6oD2MbAvrWNbvOE4WZezC5U7DrpXFrjVVex
Ery+BQGkkzuPAXnlX7JT9Q4t+kUfkNJWfDMKLJdQFwgXWUMOvbjnp6jOZTcCduv17c3084/hyZNg
d28bC59J8RJ5044Bsxwpg2dMhbnaLa9S3i9WeBGJmOwSiYMyKhV25DCwxwc8KoPStsLrk3Um5BQn
arfOB+nyjUk0G4pzgz1Zo2P04nlxOuUIMN9+83IKCIp+ntZYbK9AlKzltHVa4cNfmgbX2bvS1yKs
CXWopg3xQDUyN9B1+oegy6UHdqLJYQIui6isCC/i765ZEivsOam3r0HbBa7PCs0YTKW4Fn6Li6Jw
DHQNNVZhU2zt1nvzIXatS7m9OBq/KQYQK/ur9H2gucRAH4pNZLifYz01tSevpA5TVr55y25flgxx
5aOND4A94FI5E5gR1CYJYEx5P64Ik9Obp3VY6WSwysJg0NxDmtteTQRwd/ozcP/C3RsoF51m2xpc
jHo+zH1ISTCySnvxuUIAkgbfwmHc7fwvAmJzobnElugVxcLLHMbB7HG14Uexaui1aX4lqFqNALrO
tX4MmXK9r5ZLbg4sBnBDj5l7gxS6ddPxLcH9IyBv21jWBczL/+KXqmDAw1Uzs/pEVMfNLLiAEAnd
WBxjZ5YVHR84moK2K/qINoZnQ6IxfP4tEm8CsEEbp63Fc4F7VnXGH1c0LJWyDmkKlEE8iKCBcMNC
ByOR20yVMZK43XxBIcT5KZX9uQL3Za5HAbZJ0zHL//EvJ0pFzOR5BnzGxMkfOKCkW5txLno9bG28
Ll2nbdlwsVTPYnTRhiVbwD8oeCgrigoKdZ8Ue2raisX1iSF8/iZ2IgrR0qi2jWev8ApOg2pVzTjj
Ayz5yeSxtT+o/Ivj8tWTmGC5OSaJ448vkS2k1U3+HB/85SmFDDqBbLXzC/EX9e4l4gSiplYrvVZA
WKtq6JPS4BeTKG35InbrHJsGJv8KR1UxJbnAkBSXO7gICSyCieU+IEJG9UL9JuwsWDCbs+fR5BCL
P9QzAmTnIJqmOt9XRAwqcG5FbbvsyE5BmnvwU2TJ4Wf4vMUbhCXBsr6ziILnCOgrAVOWzcjIn6WK
HGOLaSi7Ur5dl4iXYCfQLy+Arc7Hyzj+zptOlkbxby4OHzF5FrRjwlUL1Lb7ZlWCT0sMLYc3QdGq
pKc+uDsuL1IGf6V3tOatQQjd6sK8r7WJoYEvrcO9kP6C7cgux/5LIWFop6rujwJNi2LnU7QXKwS7
/tb3oaRDHaH4Civ/ix4EG6iNzRhNtsOmk9XvHIVfP6kmgE4oTK6BZ/k3xQkmROzFDFO1zfLjZNSV
YrEnKABHSkIXtzCjZ9bGf6Vh3NxhHDN8clLyLtifT+VJLqRg+nO3QE2JcTv+tgkjhiIOM/a0M37y
pZtubApPhq3g7G4zgI2+LAMpQ9DHPJaPjA4N+QPyGC8qQ6cPPYGUngH26+j1agYs10n7OM1ce8+y
3PBlDoJMzdmMtdbIy5JxJ7AXo9lwMLFCJtXClMUXJrwShuuC51mc37T6qZN/e7DU4oh2wzE+HIQ6
HDNNvAhg6+8QJzdvjT6IUYi0BpWnoDw3Y79UXbQqHR/rJ5VmYBMhzSsjDEAmAm9BfwuTAJqB3/SF
WHu24PA7tZ+J/K1f0lT/fDMzD8Qgi98VC+n6P8tXFgyc7RxM8gESsU67xWuqWqhGQLous/d1xqE7
V+PlRUz1ZBm6fdnkz7Kfs+UQsu2yOxaOndVANaWLrbPpjWXxwqNoLdOqRhV/nyKk7m6DWBL8JDmS
nBG+2fthnDaAXZ0l0U2u67C5OZJwGPH3MC9sdeSAo1Qgr+bRtb+LVoZO8rC1JGVEzf7ZeMfkwUFl
WMuzjkmaX7xBW1koMzr18q/Bjxivy8tqngVW9gM/gzS5M5Cm9OTCmXIMgiaDHZEcfTV7dpcK/EL6
lA6LM3F+8rjGo7z2VzIN6Z6v/EYmx2IwlBwk98CHSFFr/paifZR+yptrAYxAQa2+N56xQVPT/zA/
F1ivxGoYcul818XgTVz/1IMq4++RHUu/swW3JpYVvmFEf4W6YDUtxdAXW9piFhJlg4EZZV0UDMNq
ycCIObkSLHA2+39va8OO7pWLaRKZX2CdOKrKSzXJX95P7YeYjypA03GYHCH5ioOIlpD088piBZm8
+mhK9EeDLbpx2rg9QGYCua+1O+k3aXv7nAEtipGdRY1KbSFNz9y823OiLsGxe54tHIvAtmO1uve9
rdGut4gBIerPWCSx4/1yxGTNn6rE00onLSiFjfF75/fjkvGvZyMWgHhvbJ3Sfugo11R3CjjrILa8
LJcbGiKZMAAK8YXspHbsFn4uITzMOwd+njHupWP7P/a+DXa72wg1V++L+yFVWf/trd8S21k+MvHe
CUqAaZacMzmcIM3ZSIWI5qRsIlMBlFpwAaeYYergdBcCb9LQ9i/gyOMpYauu4kE4nJhYF02vuFsC
IH069LdV/SGCxrH7XweJsaMSdbB9yXdRDNAeDUpKsK6AABkcOnJWnx0ZT/9b2sYMuuhsr3mCjK7X
R0Rk20rtQ07uHx0/qWWve+rAjYELfmDivHB9zc3iFntHiLiJ4WluoYCmY5q2aYJsdmRRVly7OXZL
FVfQw36wGJWAtvVChea1EBoxGeUdo4uVkaqvQ5UmLYW5I54mSK1TyluH2qGMLl4P67PxZKFEROB5
0HGJriRZhkg5SNt3e3Fez5c8EjLiKbyA2jmyUpWfAlLuNEclxdB4dNplbtNtoguoai7qQBKzoHtL
M30HRL84w0CU+PZaMnUVC2t97v42BqASJ/G/FrF+QAqy4gWFm4Ybmoi0ihmxQW7afK15ZYKo0U0L
Xcoe9i742eRL6U0R2xBYNEgwSxqy9THyWNXJPCZfi1pAPGuxlnOur6onKKiyW81vb0VODN21lrJz
ZxutQN7wDskGA4saasyjNwBJ20d9qvSL7vxItsumFkL5b3ybG8LLiFq+CZhj4yT1BWFh/3FnwBzb
nT0/RW+c+F5IQ6fPhdyNULz2UCHKjpb7fLsEF6gPEwjhdqtX+VMv2xPqt+YQ9IRMm9KtSb+AHCVp
Bds5n6m3Rly1oRNimnmBBn62bV3fZKKS6qCy+4NB6HQUZcrbpRA8s3r/XXa5aR19V+fZAH5q94i3
ctBFFdxRSUM9OevP+wEUNlQxMXcCLbuwbuYqLWhKxzxywWvS4zERNH9y2PRQH6+gac8sY0yzLG5l
cRTN6GJOa1KYhAeWgxmRFAmaarFHU1K8yg2qdyPqIiF3+GRHvsJ8w77UwaAwMrmWHkyVS3ClN4it
rVBVoP3mAQ9hNVtHeabBEUMZR5neunbfk7x8/SFmmF/TvoxnpkRPpneEoEDZAdoI79RJmqvQEkEA
Ulhu1bxoDa8t4GpPaYLkbblG6ioAPKOIHzO60mBy34lIVcS33DTn87y6Kczv5iE/YxKkkbFQVrz5
dxRUszKH7Fe2n9OGAkwCZv69GAYqlGO2B8Y6ROkRCmUGlBUAaWJttSWgJ3ysTJJheliWZuhB8RTM
CXW+KLvCmq6NabQrXNCBq0UTMeDYtEo5SW303YsVRslM4ncmL8daqcq3iSgdrwY+KgKee7v9jh15
2BK4cctlFB5GK4askGvZ9f4WTNL5dOuFVNrbm3Xz/7+IsoXAvygNkb6X6yFXWPN8sHgv0HrC3jUv
mRs4JM1CHvp7ZZCg38kLJMEAh+OvirKUabSYPlrTrlFzxd1CxA8xnybjVN4rWdbgxzrIbFlUhI03
APBwWajYagK3tWomFhyb/bnWpozY3fwYL2J4KzdNqQycqlJBNTqQgq7lf3DuMcxA84hhgSBpa7pc
F7+ka6l1O80vM40216KZT6fZ3nf4K/u3wGwbYiVoSbhs+1TyMtcibt4eM/yHao+1bE0rTW52l7Wv
lOR9CWnXzZR+nAGDo89nWFoo4nBF/88grxVyF5SY8e+VSqAsSQBqZmI6sMCPT68PQ9y9hOkGK4UB
rHgTpsYXfHNb2MB0jPRprsqyVOEye78KwfYOab9fZmZKJaNwdbYjYSUV/h/+WRfVqL1uFqWOACOa
BRnh/7z13zB7twJL64elulaA9PKxTNatPppshd/iybN58pEEJp+dKk/XUgoVxpZEQMDaDKkXLkpK
lJppPLiYDD20znYP0xHNCtTZ7ldqSpekGtvErxMcfcRymoJXZ21NyBbfjaLCkF2yDeD5EasmIEb+
Ho3LFA+6GlqF9tjHf29lNWz2nY7sEC1Svb+1AERcLNoWXWxtQyvuazOrbg04HUifmkRPFvgvz2Th
TBkFrpejOR6eHUrNkEOZc/sfT9zH7yr5AKcRNcE6+hk2TJBAs8RUzUSQyKnE3qlGYXbQsF91hmRs
/ycTwAxnzFcRsYT8Y9kbrYHLbcMDnibYIQLZv9AziM40PbsbFT88PrmIPH3W00HDAdsvdKztKSqR
1rTbIjB0Ju46wi6ClW6o/aKPfo8q9oAGFYV+aVf9L5YY2mBPBRtspp1TBb93xg/lZSu7kZVx6d+Q
KEZkFOo/iC6Zsl9bA1hebh2dyXwCMK69UGcsS+Hd47zy0g5kQrnitioHstNdjKAobKfKMIi7i6Zw
93gteEBr4RCW8EWWvEb6wgakeMqdRxyryL4ssg06GBAHtcCk3NIuKitHKXeeagq44C2vFYZrPx4U
/CXyu17zgmUdDS2NeXKwN7jB104hghesRlQA8/zJ8Fl9ZbU7CfBxEGVRYKkX2xkgPqNRaAZ9ZeRL
E3DOFe7/JkLzQIEZ0dmdIM52EWV5bnxe6EbGfI3I/XKD1kqYCVp+7vvdfxwjO3P/P7FDP5zkFly7
GDLQr5dpS0cUqvhStF8CM0eJg3hSRC3eETMJ4S+7X9q9o59mqaYgYWMe1kt9n+2wQ6LTLZmHP3/t
8WFrs6Q8ShSkU8D3EmtqNBPJab7cMF3dAMaEwyeTRsjmZ2UZzVBdVkTY2RAhR1La1KcWX60U4IxE
Mv4yZvIqw+PIDK9rcocURcEYhpUmT5SVyzDbNB/RO2Xs5DKqt4XhnyrCeyRdx1HZrxUtk11A8CYF
ECS4w5t0kN9lXz6UdPF3dNyPlsbovfYLkRQ28bcG9Rkgy9nNxNaP9XqYl9phrPUHvLET46h46eTH
8kph4l9PlbC1aWTJcM9R6VhOErm+R1kxUdiqFcwI1n+iCTzMw0/rtPYEF9LcHP6oYfSgArkDYcWm
6bkYHSGQYrp6PpdaU4bs5axqGpGk2nAbwq+q7sqAV41kVlrcs8LhsYpRnex3k+LrDg0q/KQbnQkK
OZMDIe63QVztn8/iS8+DChjXGUJGcpVKkZIiey42+PfXhBGEm+PE4Ea9RCNcbJ0asJftUh6X32O2
mCGaLTpcxWBWRxmzcn2uOABK/jPABR7PP+4cEEHDe5bOrQxqfAJvxpG7iersBR4QsbKfRDMdw6sC
7pjVjcGaPSPvD3jFT9V+MdthVLQ5ZFDZPSHkco2qVw1q2agvDa3aHb7hLkumMKrn3VrZhbMGHyKp
W8yq27FojK7SIjvHeRw2+l5zS6dvDu/9MJgfefrSR4WRvBdW0wlFcRzUP4/BXwBjGP3M/VY4DDja
2A08CnOfdPmzLsHvO1J2SqvS3hv279EyoogF985j0DdKzyImXijyotOY8HipYlqrXeKWnEN4/iEX
Z5BHgY9t5XIZyIP4FM2a+VVUB9f1Z+vEOLkIFLy3jZE1HCN01LxozUaY07M4KmzU4MYfDhf7mCO3
ec9QqqXV/fGMqovlftbJNdAXYXb2Xxqk1EYVJYCQjO+OLkRcPuC57SnktoqXTuSJFWGY7w9cytKf
GaLSjacAxTKURt9AlNjRT0oBtXi3MqUxaYPt63d5udJMgDVxu2kxRAioHmmSagwvrJ9g3M9otc3S
xNIOB1Z0ic2Hdm1Sapq6w8UU8ohcqfT1Dmad0V0olpD74KClXcFhpdvvAo1UEe8RhHqts6NF6m5S
tWE35/8KtXH83fIXWwPygErjUVtRs8sfuDlKIigv+UkBDFoYfa9XAVLWs5fSYDDwNhpUgX1bAnNE
X6MbXcu4Re+avCLCOaaR8dqLPSzOtLMke6afR9wVyjkmUSCtyBtL8bxKk8J6f0xxRg4LCG1DE9+P
2f+LGMvEwIzm3I6JSe5gYSg07u1GypSg7YVXfk/YnZZw0mbwmZun4r+/WZnkPwDuVIOINZ28ND3E
MY8FhlVhZPwIb5LsmgkaJb6/nNdJuFahEpDKAuLEG4fWAOtMqe4IrIEp8vfW+yPWNPW0sPJ+x6+E
KZARHMTTveJ+Bv6/kS5KsUG+d+M8NcKkaL3ja8bdHtmo7f4dI4lTnNcs/QtnUKQsUAYwWWmiF7Ia
jnIZw1/tUodW20XHcYJZAfk87yXIWTTAdiQHuXjB4cVXxx9ZTBAcYmgrcjtgUDWZ32Sd2X/eAQ94
EFoLlAPs9h7bDoxlln863VYXqbcNkl15WPCQH1N+bQbidCdTk0zsRI/pkDyxWnYxmKWAz5ZiSgoi
K1Xqg/oatxuYNsV80F1ICt0c3ddhrA/896Mo9TLGtdzm7QyOgSstGb7hnCSr3G2S4NaPhZprX0Uy
MmvYZN/Tontn050Lm8s/1yh9H5sF6REbRiJUk9i9pWyFRMpqcijQZrHHZbrQqctNdMRQmABkn1lO
fCcxRvaUjCj0C/PamfRF3ejKxmc1K3EC0RTDDxn4R7GaA3eD0XrnMLIi5WxQ4/s7DgnQfiF+ej43
jP9Zrf0jDFdk630FKfbdUOaIgGNB78olry1/XeQcyhxr59eiiSSYO45QtrSFsP59mej6wxq0oAk0
UEJumNRpVppGWGqux98dJA/gaM3ZJMk4C6x/Gbd1+pRPODsUIRtZhur+x7cDN+DykvUO5UClqK4m
g0Yv6jtG3kbTgPPkPgN8n5+eBHfbPOtjuaLChyvSs1qnX+3si3TxPMN0T5gBEs0/nI43EV15FLhr
jWRZAKOIcfSJP0z6sVkTsRGZGYdfGv1qSY3Ane0Q21mlgZtP8q/gkgL5iQaPouCE43zLmI1XmCzJ
rhXGlw5qdRhX7fhmUsCQPoT7NivF5rdjzepr41PAYGm4dOZ7VH7UoRuaSYYs+/s26JeUJ69EaRRw
5/Ya0anbGoI/+SV45Cwxd/raWyxpa7ulmKL+ONoocfncbM0Y3rhuhhIZSPNv2Bc2N1Q1g2HXq3T9
aXk8v4MjB6V8vRYAdVxhRrvkoa3dMp2SNqArGXna1MIwXYrl3e3iilVfDoocAkmf1I/DUu1de28g
7v9Lb2IfLjA7+aQ8mcq0YM7/d+1auFdc39FxOuEAA+y7TVUWAkbphl2rXyd5J1pTKKBvKFUN8MFh
XPow+7xnhyaDSeF3JSPFJHi44Os2YFilLgjyS0FSmccgMm4F4Z+XYBlZjIjAqkWsR1VqsgXeHnM/
D3Nyn18sO8SbFpn6p6l9RApf8BhwbfvdVLyjuFYD/QAtHIizXje/DERuA+kJ1jz2OEDXZ87p6ehh
X9BrbRGhb9lHIVmq1t2f5bInQhzU6TqF+T+UFJkpUW/+ApGtdePGMV3yD27F0BS/5e6VB1KXg/17
hiYhneukcWaaNuCbOfXykBUpWwxvkgMVz3RjibVuCx66AXmVI467xifq6vY0TWH2A4p4cpk2tqBQ
VkpWiTZuAU46vjIvOEbmUNgvamb24yjq57urnLcGKYdCVztb8zG+AczHcl3vU+PuqSJR85HeNMMG
sBYfcwBWwhOnXdLnAhkDzRHtm7KS9DGaJ955nOOyKKhNk3gEbKOrnaADzTw2splkkx8dNNDcDiqz
tfjxmdH2af52ZGXk/CsstGLWdMpN7PnCw+Me+yoZHZS75m/F0uWFW6Qmdrr+ehBfKQNLFX1ybt8U
+QDgCN3nY/b9zDGsbpDPWVMmUlS+mVf1qz698RP3QropyJAILD0WHQMBNfeVMp8pyVy2Yka8/lPI
imrNCLMrVZVCf+/wvx4aNX0g4bHwzUxOfqTdQVF4Q7xW2DxNSSZLbRkO1/gB4SgfgESBcKbOEQow
w6b0fGeTtDm7KtmjFsW1u0ULlaRlm4oHw1zakmT81SLnnG6KADzZcjMMy3SDrpq0Z40J+EAhgrZq
r3ucaKtbHEagiYBKjr33w1URlfUF+1wCf1tIvcsmi0pPe4ikmZVd4wPn0LNvjhgOKpG8k1vZY8gs
ffajV7yM5WneV3v2cN0J6gKHw39c1gevFXhTbFhhYRKEi/KE82aQqxc/r9Ks4YuY6TkcIty6NSxw
EiQLWhFMScbPTjBzuYtscoQEEESKDWGi+uOItLa+tNiU9B1qtr6CKfqI4ENYf4z17KEY/r7DeSwB
tS5rnOwAL525HNSrcMJODgcS24lzsbuyF4wo0qxL5ZHJPyrdw20woWJByqD6nBnLdQCnc9PX8C1h
IWU3By6zBzTOQie7ltz+bAps6xjR74cMSxVSarWRjHGWd5cift78WtvVweHnArZBS894jtL0xHkM
+FlsYPFO31SDp2OX+6eN/XqpujZ13wjkdcdB8w/+NwDpKHGllm0GKcyYnOSmNZ4Yj0l8J6QBt5ax
Ot2ppEJBiAxUKJDlYGzFZn61vO2YODGtzBB8n4MfuCdy7cqFy/74dE+alWm1a6idAz1e3nj+Pi7O
mfXfK3OO+TWHjMV6kkXhR2roT80JnvDFojn4qSMo9LweSJbhnmXBLV7ObeGNw88YZZRAwMnhCpMc
ZHZJBRdsSpC1OK7ItwzzKTrgw+s0eVh7tacMzdc9hGasAND2Jl3jiEGwXRc1P/uAcLZy0nD6i493
Lki6QaS9HNZvs3ZmeUftlkXQKzhGUpv02wroJ/mb1bGAOEtBoJGuXg78sKCt6vq3qldSSAXuOKhb
UyIiXjz3kUOcyPJJSJCJE4A0GITK0zVZ/yGJQ8zQUIm+CRbD0uGxISHX4oceCEHeJRGn8TpcPnhK
wLLj8H0L4GkdeMGUz8HT0GBKm6RDAScPOKf5hyS2OZZ8v7tpcnZCum+ulkRAFdiQJS+FtJJEdxIZ
CRSPZ1lj7PiQGaFxB/4iQNMJ1BYW1qeNRZjVuN2xRRqTbE4A3VDLu92f4zjn6AuaDIHeMWQCkrqV
exdxFWG1cxuWXCbJlrD8WEU5QakeqeWalsBQRcSe3nmlKuqF7dsxoQbqmpN3zEbZgoQRo6TXXbiw
72k/KsGkwaElulIjD8pFzyF2mDD85q2yFN5OqVqGykPQnlJ06LB7VKRMEahCKTXJRqtxiJPFhRpP
7AQ/JpU24zfhbwQn9FqOppNLA5FB4dOP5uzCSgJ0jh2qHOU1xz2GVFdDqPSlUtWaf9xgdfrnSvN3
R3tUQD8rZv9M80HJAOGM3SAjIQ5VLqFZReoniUZBpekJ2xHNBMKnosz8mVgnomQt/QG4bPNJCb9U
T64Ia2oqGgig/7m44Xuz7dcZIhm9O66R8oXgdkgSNXIGdc7m4a2SrQhTegwTpHzAQE2UK2A+OOzC
qU8MUFLfAN/jUqlTiLPSWyVGBjVoW724wzthxoI3TPFwIEt6KTE1arVG915uPS+o44/CpAocDrZc
UDP7LLu+bEIYydm8KsrTHVC+ipVILCOnteMiDoPFVm9Q/THJEErbg8vUmwQMMU/8jGXAFUnVQq7+
tj0npcjxoU9FdtM0Xuxd21/iE0Lmnh+faY2t4bkXVEi/ybf596hkCaAH04i7kTTCUeQCcw5Intko
xMtEBbvrIqM6EnBnmcPc6Vb+E9vTLreh04GAI3i0HQR530WsmTfi+JExmWWYCttUjXbae6mCY1cW
Qiy12zKxsEwE1k9TSNoCV9L5ygBBlIGhccRU6ipJhw8f+V+Mv2PZAlwav+9aHK5Q19WHYSL/WPcl
gnKE1X69txKc92qzE90Pr5/uuVTsWk7QhhTNuDkOZLfe7+UoklsW4wqxXx/soGEhQx1+7TGOPg2b
LrXNPPxJY4+m2cxZ56eso/+pfhUcEMvNAlMEZnwtha1RaL0TSwAPMWTAHj4lPOdTm90wgqzGP4NU
xJE9683xLrUCGPv13ZfydmcYXfRreQ7RhCled2al6P7WhRjwbEbvGpUROkiauOGbyNgSEhJBbaEN
4Qwt3vUHHo0lg6TxeMbTv3A1qp9pviwCCp9tjK1ZngEY6QmfsSnm7XeSRJKGBPTJV7mS/ZyXCPi2
uSTeWFC89hvpqza8Ciah61ZNBdImUWiQEtWhEN8AivpvUtnuxMWr5RH4lSjzjFvZTsEPsEHAa4z4
r5zOZ5CJ5EI1cZ7YL7iyCOwb1fphnEg/YNpY/5j3ZkJEORVTGGsb4kN0qyvIBok26S17DV5cjiBM
RIVJYUKUyj5bx2IDu3S6449+AddUgFjrUsT0dM1botoXKu63ryJSyBWaJCSm+okrbbKbzDpRIbju
jsen2pk4vPukguMFvYBx43ihFZe+pxvpmvaobv/fhvVssZljXJyG9zISqEUUKAcuOx+B7njTocar
7eWZmhZ9C1dlD32tRB1hEai9tTBTrsgxsVXgJeGkY/dnQ4pQmZN+VD6z45gmacDgLAylusMaFpqw
mLTbVEX4uaREkiEUt70ftqpe4ivBRxYn8Wf84Bp64FbXu7uo4om9EVTTf6DKMzgVfZjf5JAQZ3wn
iJiVN//4TQPvLlWURwMB/RiH8hZ40fJSWTfRljin9bKZ60B9LN1m7OFIt7u/v5Z0h8x0oZJ83jpe
clpqjUe30TYbFXQLWvY13eGV1IP3P+Xr4acKmRXwoYK4JjEN7LORgKOtgTXmxJ1HodyBbZtqGIqy
aKSz+KkvGPi+b05ddZUwTfxOj7PqWzvAxBpeIGzhRJoClRYih18YZPbLDCtneWNhoeHNTxJZi2xI
zwDUAym4k8a9kBCrUTCxMWXxqFL/XsnPYHxWbB9Y7yCjTcAx/BD7iNEReJMSTKEWD+yPBJxCgXrg
1bBALynyWJ0fUXYMtdOtbYW+qcjF2GHgN3QQZ7ZHD7PYYJCkTchx7Y8n4dyLGgLVrha4gzkONwy6
dTkdCZ+YF5sXuW1gCrVEja0yP//Qh/PJGdt7PuippOJnU0pnKN+cMqZXLDQZRVXHqkyBYFG6Lvfp
AwtHBPWrNJS3HJWyPzAtt9SpUW+s/iT2lBbcfX1+iIUJAktqyfzosOBHgiLt6DMvaAj71ogo6Ozl
pEkzLsHChXY+n/JtHxPyMlyaAE8ytkQMMsl2oi1ZJR5WmakL/nHtNpbcN1VKll9+vUte2lHYMT7H
hgvTm/KJZHAjB9E8hG8fvuy3AcepUEe7cLI6G8Zvox4UbzcJbTh5kBjEEWuhWn/v3AkrJ1vSZ+aN
i9oZirLIsqLDM/pxbZrmfLwW+kC2JPbTHYh0LXCFLstkXxDnOH1QjTYHXEfAlfUsB4ssXnqjOTs3
kB9/7vKJcl7kY2lAsbzRI4bqRIy95wt2/HW7bRY3S0/8PAJLeEjUEd1Ve9sO1sReaDv7PM7vukVb
dC9e1ySIbyDxrs7xRtNJ+xR5DA5XpII+uFUnnBX0IE9MLE2miJoY3Btr3WF5QGmildp3KHR1ejWN
jl8oDK1xgZJaDuzItx0gNnsU7QSc/JSbNjz6lyWrOncb+KT/VLIEgXgkVXAThGoLIU2EZNscEdeR
kXqtlr5n668YKTFp5goWFyvnAka5EesdctqDGjnNN2DSwG5GogskLv8vR4Avdv0FoHsOHL/CvdeN
m/KI+QGwg60jLKZcdSHYmQzTBhTl4xGwR8pgvnxvIsFzrMeh8GRxAnO0/ZUKY8nqUs1KTD/eQgJ9
4WzTjODoRw4QPn4MiKgOrPOPTPwM//xwQP7BAiHJBe6nkTO8OGlHrxkNkafiL5Bmcg9OhXI3txP/
ENQfVYrvvvlXpW/nJRSpw9MtRvG0L/PmT9NUYTd7ClZSEVFgFaPs8p656uM37c5gmM2V3hu2CTA8
V0kiKQX/4qLB4zWB35++DF9ot0bUrYusOn8KyCje6DJd1wGVcISYOcLIIMYd8+icMRnLImOuDgKx
dMdS1BkT4tX7QcnC26UtYGbRhV5L1qIU/MWoIJ8RcDBRLBWEIYF9r2cQ93PAHnai7KusRrKx5to0
rJZF/2DDpAIH2mlH+ZuxQm8yzenNwiJjaU/3srNlpYHz3Fym/y6npXa1TfhYO7uAuqARmupUnnVX
lp2ha1b9OCn16EFkCw84FYZy3i6xjC3jqkip0lXCAoOP6HnmB/LqrTRlQJEKNe8NEDmaKQQEfcu7
MkAv5iD9M1lQK68EJBL/o9Y81uorPAtX5DJ6obzXqjky9qg0Xec+iO6urrQbYzes0ZvKJhJKvIsW
TdSp83czue5puNkAmYcx/zfxe+9G0iZCq8DjYUfs4VZ0gb570b9L8q+RGOkp0v0VR2KCI13ViWbG
n/BvlFQiLR8Wo0XlnDs8TSGk5Z/WKzqbUUHkDfmp18rU+/1V2U3iTDjhbIrSNX46VCJ4cL9NcVJA
mLDK5iGxdBrFmVPhUau72HOTed/Hl+77fqPKhLTxdOnUlbRd6KgNTR9ILLUbX2SCCPmRq7TX3YY+
t/1fcaXqhezwJSBzOzukf2JrWJPEjqkIuip4jhRE60jUG+9wtp1u+sC8AcI71ZFp9EFJWu8HEE1U
8CtF1cPu6wtRXxWDsKGoi9YHO+h1i5DYzZuFAk3nxJuYLch3eBviJL0l2JjiARyDWlgRXTi2JT9G
CwGq8h04Zt0a/qwf0zH1628M0tl/mh8tsL5IUneKBPZTyvtSG0rZi4FLjwsTH0/x2WMJhRSGllfx
6TShVaatpT6G5aW1Ha5QwPvxE60o9FIhn9pPJkYJsoqyQxCUhlZOEYKS4GPk/vavAZS6K6hOdf1L
NqUWk9CESCllhZrxIX1nPiBc6tWidbgz2+O4ux93v3YxkY/sKEJgDQUg2U9ik0+XeibDSI/1vP5h
OJTSx2yD0SZRZCAXXj3Kj3P6Sgk5FzZlHXjeoyzkpomzgEabIiahCq7am/TOqPeEc8GO7G8rrTZH
lAlkW2KrvH8CYlvHHd7pRdrxv2SoRBjx5+5pEW9+MI2tKFADs9yA/FFVnnFqYm7moynO/eTqTt9C
kMR46b/bNURLZx79XQTwVpM2Ir3eiq1vdzJhbDOec0l0fdXSAJJcNYR+Zx5mOFVBrCekabU5i5Z8
yTugcWmFlo/HPdT+eNrzY9dA5ccy/+wl3sSMNxSdPrK0dv2kTFiqZo/EPksIJYzFRNWwY0UeYWRp
3N9LVft6u7gZRAb+vgAgKjc1gi4uuj2wSLBD08qX+/S9V/EUjnzskVwT2PzapmKaDmS3K6zoaszp
WoNyRDE7kqAG0/vdPnc+HuC2Dy4BDyFdeJCa/koG65/uLIbX0iYTEiQa5+J4WVnsWWLc099wFLdd
wINVvSHmQS/bbQAWWo4lFQHr9E2sVoLQ5BJUDRJmubm3JsCDN63Nkq9B7goONACL6hGTbd14XEZ7
6/zn4ZMKJh8vDhSRA67B18Lllqc0cFtkGFyGidXr+kRl7GvaknOHBadkKavRrhEBShgsHJXc6aEw
h2G0ad8rtQGdKmp2IAKNybD1kPFed0eO9N5fxagtuzhrqcgIj6c6u6Yp8g6zj2WdTCDPQdBkxTw8
k35aOVvg+93V7ZjyChPaGtBK/oNLto2dzm0HYqNWZcusms3Om1ej9G6TV63219s97sTQmhDVXtnw
be/FoFkDKpEDpyji/HL18hEmglgtgQvf/ss22dz9W3/oi0BHrzC7vwNpDK2Aew+aaZVf+v/9g19p
u11Z3Rz+ZrrI50fhl13c8lgJRnLXyU++7Rx3ZuqNGbVj+VIAn6NendZb5rHY1TnX4E2C2RcR1t0Q
yqemGjsJd7Izv5yUIlArsofEHnryOSbGvkc3lBf8wengaILYu2UMN55SduUNsRLbnDrHbbhxjqYx
9i9mj5G6vwXqYQM10nQTOHF6AgIdmF/Rvb7D5BPW8L/GZJVMnR79OyjY/Qu2sSvWZnBxPu6V5FQk
1KDgybu0LBMvXx/BLo49W+fPrdN6PryukX2pMQF9KwgJB3Q7XVDMIFcAbjeG3Qh3vtVD6Rg57yFP
P/bfa3suqH2IuKCnRSxL/4CtP7u4PqByCG9W9meorfhc+vY2HjNelBVoj3Wy3/vW8L7C/JkHFV4c
XO8W0kP+G5/zU3W999YMm+2ffKjXHeD5ru8YscMosw6AreLJtWjO7da3nFSTs1L+g4O7oPXGv7+/
qX86yqbzrFZb9k+8D+UkjHjGMjwczdTXRo6yOpQAYBB6KnzKwtEqSO5Ehci4W3WWtX1zQlEnzaQk
8Zu5yKUkuJ3PbZ26wSvB1DLE9WOtIs4j1IWTHUwQED5mC2kWE/ZDJ868qR2OUmWweLyF30wElC6m
vZ6bRtXCFGoeYl5cUdu+gNQPPJ00zzkeE6Ikkq8rQXmPIfh7+osZMRFJx85/hIgdHLdHOUQvF+wI
IELWAKOOajarahl2xW6gMwdQpYuE+cL01orIYmDZMybI2+i0j24J6gpHsoiyFG8s2piBHa8C+FkX
x/kLvgE7Wg5jdQIE2XPqBQMaHqPsI2PcPbfzTGBW/lQkVrW8U7UiGNEJAfJPvkzS2cJCJfZpNkEt
RPY1P1mxaTsoqTiRm7AWynfZXWYcz5dW6dwPHX5xcqxO8REwX67rEjGWrhROD1iIVo7gO5QRTnok
/YYzs2miOaUFJTa18zFcamAnAJJ3eLgwFmMUE4Yi7fhQEbH1+J9yJ35XprX90YPBqZ8Uiqis2TWz
YsGGENkbdEbW/65rDkcbvYoPxZETZ46IQkvrETamadUygAA4UXfl3DIMMdoaJg4FZPT+Jt1/kUb4
wwV1Tw4UMXtYvGtYU3PSxnbYBv1gb37ZsM1d15N0QFGjgF/AUqrQXJBo/kKS2LmiYyjhf/Llx/Im
w46WJwhPwEH5iNiDtGUohyq/o97FxnQWBXV9ieqQhwRa0BfycI4XckoUs88+ona72JtwlX7M3M3I
PqpOCaUfTqi0Q14ftD6UlACa1fkZvEEb/L7lZVe0i3dU9Uijy302UBRGkmqM5djvgY+kz2HUmjKM
69Mt+cVCRFZkttlWF4zFAfJWv2xdHE/g3lcRZ2DyJFn1/IySFqNJxPMXx9616PVB5whXnrAP071H
7D9yRmmcZksosyTXugoDGDwrU4YYwIrurBzdBiRqk/4Dl/KdP2NNia8akUdp/lKy8kKhoodWV3bI
9ikRY6oQz7VLf6SyRA7RsY91cBR6rEnu9OIATprnYoajikgqi7OiJm+/KiSjSj8jx/px9TaBj7li
YcPB29x6haFfwTC1wAWdvGXo472dsK6T8hDjKKo6iI5qn/Plj9+FQcwOCJBOAHIMldkXDKCPlaz4
zfnAMVLC98e8kjGJevCKCYuELdkxPLg7D/uatGiHM/GBvRe9mLj7xNClw/UWKERze8nydqa7EpVv
m+a6UxO9kHFmF/4RwqUunXUAl0xalv86KI0cALbmG/nWp7b0khSxrhd7dJE8CEPtoymPrZVne1T9
cooaPO0peSe8gmSCBN0u4DPRPzTiu4rwIpC3g9McPezCi0eegVgGgY4b2h+oveX5q802KpljwkzC
Vqy48+zcYg49h2tKt9Vg6kc4yisXwukN96jMMLpWbuPkNVUO9Se1rRxYNsgZNYa3lrq8tE96qU+w
gaOti1Gi3138+Igf8ywtFt9RKzfOHZZ3445ci9mGHYnXW4P0LDM9bEejrxppT9skoLmaEicUsgdn
fM0glT2EkyKsZpTBCwJYNoI3f8W3dhf+k0aTXNT4gNPsVfUw6622J242Vjp1lHJ6WdMlcjwD4mPN
NgZxXppYboEHFLgoGCej24iz1Jh9NWN8kSKOImA6NV9ZdPJXl8oq6adsIA06f+ZbdbJv9T3gqhNR
hr8NRLg+HwZ+KijtPqrcX1dSN/8oyD/mE5vsK9Dhtg8QibNUUwAg0N4lMDyopSVlWypqhD71h6of
2rRVeIOlYxsE7Ays6Qkesvq9YUx4tL9senq6KoevAwe8CzTMfSPt+/qLu1LoiKs4nW3GNIcTLUze
EHkh5yKNWslv710nLxqQE6b92oWWdRMLsHs47xy/oob0OlXBE6hRtO+klXSyRcnnVdti4u7TIDLL
nMl7jlqbPOn8MOg4I1j0E5b/sY5tYuP62pvTMsU6p9DJlUx2DLGD17kTKtVv9Q3fe9c5p5jPDmcl
J9qhw4+jgzUpk9UIsy4EtLP+CpUzlZ98THtdagAiZASsZHkpc9CgrizDQ+O/9JECULCS60MPMg3h
Y5jdUgTYMCYXzFFYjYDoK5jGuGM5QOnC7aYnw80dqiBHxlZ5rRwA/VVynjnuXP1cydihLDTFoL58
AZUD4RNN8VwADho+Y7RMF/vtwPY7DwgdvR5vEVLJKAWw4v4mzNg6ev9kHUtx5cYLFSE8P4INZ3+M
ckxpLuof0YlMQ4BHHV35Qr5SUXhMvBQZsXfJ3dQN79B3/qQuKquABZL2nYdhtqWMilAs2E45ksGa
gtTWJCnQgI0wy07LPSePkY9bmGJF0ZES/VNEgDRqsP34YTd8ItXPozJZAxR8lDcEPoABXPgdW5So
013kN0J5dc4rjJ9USFkxCJaQ1X2nBNJrnGTurMTlYyyp/OXFPlEk3Wb6uKdJKiQfHQO8EispWDpt
4tYdE792K47s/g46f3x4r3/nVvjHG6s50dFtxdsSXt1sVdzlKIGR1TNVYcxhrqqpMI3dUa6yZTnZ
E8oDPw0nrhLRa7VPOZiA3mMOiuYBrgwfnIvo1Efi3hE5eU0bF+p7fzTxhD1+lNIcRzGRIkz4MU+g
dryKadM2jGGGxCYIZCK2TOmBidgXBH13lQh7B/zbSKEg/rk0JAZ+nmhxynReKOQZqZ7tn7LuOb+0
wKEzgZTud2gqV/Qhz2IFfDUcqgmb8vw8QuDUcklvzWdqRo3vKGp2Aj+iagfNoqDLtz3NL7Wi6Rbu
/jUpq9+UNdnPf/Vh+OBRRAb7AmUGqOM1QsYSPLDRR9R2GIeP+nAuCs1quzDx53R+kS531fjC097+
kaucKEGEPJRlaPTbMIFEIY2nSIPLX0nOkws98ahhHDaIHvyBCX8RO/lxR1oqaZr9OMPosAhudq0P
SAo0TNV32BBzClt4X1IhByb4UGpWfU5VPN2BbD5sPjTKuUMKu25S+StF3j0qGU9Z3T7kSiRjSap9
ZU1z+qwkF8Zj5pu3JhOfrS3WZEq850p4nhm5+MVbjp6ir5XteN1fp/QRUZj+oUYiprBdDGFAu6Hi
r6orDFmt8ZgoLLHojV91ewLR3pFc/bP9TwXTQTLaB3/BNaHx3YMPlrRePgj8xvA75HyGhgFbOuq7
nad35BMZfO5F0nJW422B6f/TIQQUQMMpSXwlNMB6agpnJEw7TnfyIUuGWJRHbANJU+U+OueFJmpK
un/886up9ecLVY7p8CpdFnYSIT+d3E3uvEogUYYj+e0kmUK9r/gqdgWLQD5Zrk9iFE/2lUq/5F/d
98XwtMkw4GtMaUME54Lez/zvGg6aTCeSl3SO8ELevIvi+P4F7Nc4VkSBW37jgI9e55/PPkuTEXAf
wDcecs1Phzgdv+ZDVsTzz2H0Ila6+NjZjuLDsBbAfpbUOAwUiwhdbptRY/nodHT4h7B1lFbjMjjF
uPnw9qkOSTItwlijFsKFsGSEx5CMHG9Eh1FEomFbwKB657MaAmBEh/BqbT6RGiHm8Xlfk2V+TG8G
AQHm2Mv3e2eU4shWG2ZlWXgq0y1NeqmDuzY0scHMoG9JfSnd6O+JKMBEiasYCe/bJcMt7TIVOtxh
aRgvkwQ/baYBnox+poQ1AB8czibojorGlldikaZlMOs/42clU7cQ/xdtB2gNwvWK4+YhehKZ3Qe8
JkwgyES7g3C8daNrtQfSn5ZDYt9sNqabXDr2nWLBJpXxs2vqxaLXhlVU6KMaFoMGaLWke0yUJnrD
43/bmcYZHePR9EP8fMkFEeumFU7DZMzEfZqNlzHc887XaIT9shduGtwnGciT3DLJZs6C8UOeswxr
MsSu1yucTLeiqTXafekBmTAl5qwXA+n/qT49Yws4AmHOI+QC9lFzTuaa4hnAvuabzTpcTIuTmfvG
1U4/ucGBGUuaXKn7Hq1pg8PfJFCDVi5htyAJ47DHDL9HbM4FbAyOffifgzuvJ8gukzDdQ1ihCQTO
7VsuDlHxQgQWr64pXoESFgM3w4xDFIG74MLgIGT5saPUlj5tBvrS5hD2lbxnTy4QVamtg1YYiVY2
+IMFSyHOq3JZYgxsi3eT+2I0FNEq6/aZ8XAPazH4YJoTQ8qjU3EXm65Z1eu9bCJK+qRp8knS3VVB
pV1Qv4MdRZlEhRtC4mx1r98Sw8uOkDkGFmOY+LjfUamujzNsxTv4TBn0WuZ4BjoUSLJf3APuNZGe
2Mp1k7FFIy7kYTZTpttTlnxcseX04s8sctASXFFcefY7lcBjDtM/ruXymAwqpG7sOfjOYMrdxxhY
to+XxEOlkh+tMOwsMm6ML4Bj9x50kgx2t54rF9eAJizOQ/Mqp4WWmVIgTCUxiedrUZQI1iFDcvEh
dLEcBiqZ2bZi8eku6sEmRKssdj8g8reTlkCLYwBLuNZ4of6MDXlFpNogQHsDUY10ZIhz7Hyd0dL8
iLlKmmikUVKyQ+w4wXnyl+zbYMiqcoR9+p2F+FqW83ftZoFSCDaBLO5aIWOpmHeO5InjqUrOwPZN
9z0QyOH4s9LTlE3z3CRpYxFlvnXEBhjU+DhO4jP/t/7iX7snfASUPe89xBO1gsF5GCuhjYkPeMIV
TWmivcCidM1Ixwzr1jSiAw8O/O6jvTUDVB8krUF2vMxE0lu61ME1uFJkGiK8r+J7VrrZpC/d4fn6
6gw2CQDsbH5R73tO7ek39CckGdpwcAW6Jb5f/XFNjvH4gXm1roZ54nnnqqwNwAfBxs3YplD3qtfQ
qZ5G2XclRQ9qk3zKncv42neD/p40xkRwEbUA0uFj45Id+w+YWsiAzJNYoLrjBb+Z13x39khw5X1i
GSViDM97uJvg744rHNqAMzLlV16CvWCpORKAsTaas6wgvC9WpGCWTz7j+ZYOD03fgkXHvOIEtb4n
K3PX6LJwZBd1GHuPP3eYBrAcwvJa2LHgv1eHW5NqVN0Ng1GMOABVBcVFJhK6LUBOUw8u+gM/RHc3
oYJaUwcd4pu1dokOzkxJQ36G1C70jPB1JxSkRqL7wu+v/5OXf9V0zazeN78T+M3fNyHPMSq7YTtM
Pj0oMQtp9r1H4Ax47NmT+tKV4S//rO+hzXJoLjSUtnL89RgyOy0iUBfGPAcXTQ7rrs3d1dvqp8sn
Rlf9j7Xb6hJAD7iE800kPet12mpH+OskethsRggP+4tF58kJaza26SkSxcxAk+KewnjZ87yWh0xh
1nbTTSBOvH2raMOMLyHKG+MFnJQFWpgfLpOWUB02IZyjkpMwpkvpLYlasqnjevd6or6d25uZestf
obW/NLIWbvmLRConXkvdMAKnYvvY8QNDoYo8isE8/qZZ7U3z6ekMPldn2DHQlGh7LdMAhEOolvXs
4k7i+IIv6kelfSrq1/66BMDk1cp/Q9LNKUbTvDiRuYLBOihXrz9gY+PXtGmrtqHf2axpk6D86MT3
TXfb1jnGKPLtsQcpH0S0CKcXf7mzVLnMymNs0w33Jfj0PL2se0Q6srLFQlGsMRl/kk7GDHDtYHKv
5sAGggrer0eTW2GMFj2SNfO9l/itEz1jI/qqJOkdnAiALxKKyf7liAb11m+47KDmdGsm8EH8cS5I
j686OnNeT+zAPzjcUubRjWEpMZ9VqrE0gtDluN8eNFiQwbnWHL3P6QalaOmk/3ahOHG1SP5j/vNJ
wRX7BmcOing0RSpT3iXx8s0y62rPla0eg02R6tHWe/MuNFsbHlb7Ky7lW/rHtjQCn9ou8IyJLwLf
xlfQZmGtIJYR+ZNIgZdmdsGO6rVvNIXgaqDXRjUBqepqSjT9QTU/HHNXqorDHDpdsakaVXngvjmJ
nJkIhVYcqplxBh9Nm9AktWYdO0zpsRDCtL/N0TtF4lb13bxrZ6ikGK9+PIZRsdyesGhNYOj76D0z
UTlRS0Ial6Uiwd9P7u8LxKM6hj51JtTroppoMFeKmyzLToFNtajMtluWgpQnQcmcOn1TzCwcIPVm
8oLKDN9SF/CP6LxZF2UnzRxgGaXfqcZbmjWhBTxOta9bHo+xE0pcl9f2f9gamNFC2jt3QTvxybd+
w/HMEU0Udt43ezOJ/AbuLjtawn89B2h0lGXfKQdD0Tr/Iq/xrn8BV8AU4QC9o9H23OpmfipmnHZK
qTJDYrqVf1vE+3ILgaDw3q64MVdjYPfHXovwSGSOaXn4tB7pNxQwVpuMraPty5HfFRQpygGROrpz
usEyfvzpPpCrgRtFlbXwLYcS+ny53zJ9BV88pqOyg0ZHhAX9z/dGt4nk+DzLVZOra5rmsgMf6670
MgYG/WBccdO5ukThywqvKkeT0EMabBzJQW0vLim5EAFQoHk7nUQ3yp+jWqlRITtx+FZrypSSvkG2
A5OVaEBjFiH5L8M8dxdioccBSPx1aafoSVzX2p0pNttsPJABpgS8mHCLGKcqKrbuMhQb2NIMGMsX
4LxFe9ek30xd8+WEnFwyurTFdeKTfqvEkayqNaCpQ6cfBe3JdyQrLTI8Kb3vexamuIE0qCvtSO41
Hc4jOFzMa/RXde3L7zB+d/IPa6DxyEfoqBUWOFXICx8Nc+ADUhXsfRlni+5nH2j4x5JEA8RnyqQM
8SMMbxuswi4ys2GVWw9IXoxrEYfK42+EieK25pUmJ4SqhUfodXf4mZe8Zj1ohif068VzPO7CuUGY
W5eOkfEcvLEqK0vTOatB1lt7pXbzRbmTxE4M4N3bNQt246kRr3IHZYn/PBfLOWKVIadpDdS0M/Bj
zCT2KgCq+5GpK4UpOA47fI6T0uHxtuqact2yBuY8YBIOoPdUhyKLtw8CnOO/bKLut745T8OlcRiE
a2gG2S4WnZueqAtf+DYlQzh8N4w52grt0lvhvX2mf0MQvRr5hBF8AeFiU4Be1w545w0xTqUwVxAU
y93adxVYVs+aNAaBZNFRbhty4aa22QFe8I3s3RhC2RLWEVfSsZDsP4iVECBCj18wrfiSCMJ6OhKc
no/XXGy3x6o6oOg/yde/7fOcrNKuflv34gXneoiKZHs+lCb/f6cG+ebq8sYIvPFSU01w1R47yXkF
Pf+Cyoz//CqY9tsT3oon4aKhG/XsnKcPX7vNvB1KsGxxZe9bZcArzcBRd4xODJNU7tD/eKhMvZ9I
OdV5rBz9uuReCuEeXwOestp989Jv1cJnBr92kDsZW0xjZco4JILvYdtPnRntvJzh44ES7cfWLBRG
BlulaTInrAjrmAipgTFauEY5aERY8+A+LkOa1L1H1ibDCeuUu8fo7LVNRvHA2JNzK3CNoUxK54gx
7xHeatx5tKh1IHwKh9CZFTp/9sz7pd+MVqpcKaHqx4JXs4rHfCJv3Sef2NlYa0Q8kzPzp0Sjbdf2
bRPfPwqXwsEZOdqa+U7QBdirF1IKIldy1COCZQ8Q8MD3V67uCC1quCowi6ADEgDjEhQdatZYPJ+g
EQP1NYWAK+Z4G0iwO22lLDkmsYBCC2IVFvm+2aQ62jD9qJGfkMVUqgPTNRhpu6ELwRYcnT2kVhEu
8J9D+5I91grP8wZp8R27tkxk3wrwFe4fRwYkD2UqgHtL5unRPeJHfN+/waIasbWTt/mm2ns5HTtn
kM3lwgLMXSCaIkKm/1jatRuQ1NWzHHUvu0YzTW+suytmF0worZJl/Q2ZLzgKK83p5JG5G6xdyfE4
0DvBwb1R32Gb6HBbOfP5N0oV1V2k/EZo7JVfAfqZu89TMWcxLpE2G7KHWDIVrcrV1jwN9DNgJas1
SyMV0FoLZWz4B7pHtu761lWiHQcxM8MPNNUC+GjN5uTO44+vwcrDJkuGu/VyXmZRq6D/dYdNpDqT
0txTNuSpbWgSFg2DI3GRO44BjYcocj4nnFFoUQgEUzVZdB+vIl6YWJ3VN0wk9OBViUE9USwP1hHM
An6ryk74ooilf7m9Qf/nFeX2z1V4isHx2AbNEy4/kGa6OPjfoG4flHt+HAuojXZE+UZeB+FkVqRm
AObc1UjzlDML9+oI6ufCg3YL7ps6pghRocAXOfGAKBdpcKN5xCgOBVOmH9tQeljIg1dlJqjMJeUp
qAVFqSf+OPtAcnrc7YhtGbl+JTSCQtht+vCGkWHcOhJxoPcmKs9FW0AhjU5e0h1Ydw6XG/LqUOW4
ZDg84IMta9gEJ3Po9qKTHQDhp3MoO3nDYHfvrWHw59O9gjtZVsmWKVcLvgKtn4HqnRDf4NEuGOam
U+7JalzdppldsiwoUata9ZqtzdPEKMHjINoXzM5cnuzTlbuGPi9eCGMoTbhG1AUJoGbqHfrcJcTb
xcL16RqAlCQw9IdWOZri+jqjWj11UmML8sGClddpvn45nWeo5ypvkxDhc/WYwV0ImUrJg+DZrSkj
yzs2Kuj0KveS9EFjMbLky5Rw4kbPfpcqFudDUh21IVoaQRqiPSe18AXlxjxsZGw0rDiemdimji7/
J/dtQYc+zdaAkzDx51ju2e1xubxxJKKf+izJWGmeqqzcFl1MS4CzAaXD7kmMGU5OuhTzG8VXyINH
yKAvcbTisyKCd5EYyU1j+aVbotxGN0REzcp2QZCqvbuomiofFtzcHq+fXSo68XaaIJzKEks65H/v
SLhOqXOIy1FH5n2hfWbLgcLBuCpfrO1fcZATHFd2Xp4ri2V10rNW4XOb8e7IrR2eCXfXVAs9FoU8
O/SVNf2Jn+gWb7Q8NHSTT1KW+TJP5Kik9MqXV0a8+owQnDtu0C/zKV+Njn5316lTNO1R2LLyGUU5
zmwMd69pCCujPiG+i6ilZmkHWSUnyBQ2vxq0aa9cGsPQqllMfWC4By6gfQ/todH934Su1QdIhtfF
EF2IUd4Brxb2wB9USZlk+T5PFliiOAnba5q/yU3i+fyKSkBCiE6Iko9Zclu1kJN/L+DbUjcRiEx6
dAJddAzBTE71ocrzPjUwDsNyA8/aXP+EF/mlMJBMBlxjy3kjpcY2y6Elv7GlVR3qXnghoahSJNhu
GE6XA8hq8OM24W/2Fkw84LLDLurLHsH6LGGCeeUq70uo/s73DGFi/41kMjqJnAraPrKmAVbkLxN2
pbeTCftZJTLwcBMZEHEs/ApTIV0AGNpqaalFJ6SsTbC6qyL3U0iG2tOy/Da1QCSS1aODiIQJ++SH
9Oh7LsKmALIcOhTyQqcoEW89NCv1BL0UsUdJjH/MNWZN0eoEQj6BFjvTlL8vo/NSqGN/YXVsYVx1
XzOMOVU8Y7g/O3ypGsr7+fwvm5aZzwzGwMYaeEY/fkBuEdofV67SMhUbyGQMANQAAlRdMANwrTdX
QGcpclvcA4G+a9c7qeJUuRfRebUGb49yWIaH8/FmHBT4QIY9wQ+8THrX12QovIqV3XTtFwwBFIpW
jqSb9tVcHNTuvkM+VBnS5arvvuPqUSH+h8n4pNvf7PJdqJNnEugNPHNX98fNPW29P7qdJ6c1WmQH
XxUSlfE3UML4GDQdS0D36XKc5E3BnTFDPuMsNgTtB6WIlDr68kANzDI+gc0aLSrOk1I8ZV/YmD2c
Q0Cv4P0/ZU3PiF2uRj2nzBSnCnA3lFDQLilVXCJDFf6Qd2xVhbkJrFlBdKOMpgNW0SXZJ+7xxgkf
gLJTcntSkS6PV1Ol2T54iP3E1FXQtvaAkOVsgBSIuf+DgPvEY8lx3YkGTTDD0XGRthf6GG8z5lCC
vYQVNJwEA25LBIy2pTQOXL0JxvI2LvqC7JRAaPw1Y2KbhG9qJ25pxY+RDe4AOlSxOjXvcxxaqdTv
uzazX+XR3zwXa72J63J9vUK+b2FjptRNGVXFnelDU/sl7ccgUcg/xdmpHaNAmGY1TM0Je+hNxwib
ui5pa5Uq7Yvz9AgFsLQGAn3CzBT2ybgYPB5L/jsq18vfWhpMLBYv7b5Vh6j/9cv4WA5pWAtwG83l
eEmZAqMUZ5HN2VLDGyCC3goXKjR9Bbu77TCSrbSdtaVc7ckNSnS4Zma+hfWgwOwb9ZAyOa8pjvDa
kJ4tL3krB9oTyITWf7RLd5bvY9I3njnqIXbl9yTjtOEMssjP/2cp15ySFNdnO8Bzb1GVqDgca/6g
1rymQa2dZ8tOj6OBcGwUiL1BbHrajkwV6M7ZORQKzvlCxT2cw84/V0UnsxqRxD3zJBVzVVrTNNUS
gHDdzVR/8/peZ0armazX7mqNT+a7QPZHt1IQf6Evbx49l6INA4c3iRtCfmq5jjBgC96U2oEQ7Idj
c597Owi1pQgcuf7+oLdVuErlG27kXnkr3+a/ECU9U0J35Yg9tJsJrJEO4Ks2s8jMYBVAqqLrNCz6
kd66fmWih9AV6GUzmYaleaLpZsyh3BlMfDRiX78W8ZI2AyRdTECyakWwNKqnikWA7+tlI1/RBbWx
juAxkEaGo3Ylfv4vskcxV8QwXqCuLh2ye/epZnv6Ge3DO6QylGBpxmLhrPVqrbjnQRmCqf9yxjMT
XzWSlyRtsIzIl3yHQfJlRZXUrPo9zDC5yD0nkdBc4BIZG/x5f4RnMN5wS1EnIWcj+PnYoQ2Sl5q+
Z2NJX5SYr0FO1GCelK5Sf+aUO1Gk4+swfhJ+pu+wGv8mM/KemWLvkl3sw7uaNVlTCWFo2SnFltUZ
pjH0LupdEYFEivMDjJAeZyfmUEAV21ueS2LdHUWsYiec14BgctEAoB+1f4nDdRewQkIyFn9NS5pn
vPMfttQ+kM22ujpb6FDvVWAvorZRcn5Rn2FdTsDQ4+iFSPCSGsBgRr//p6jkrt9pyT9PYZHnK0I+
FEi7vrHVcjXP95aL+nimhUsC4Ys2gmrAt9CZQRkW1cdHmdT0fzDcI4Vx9c8GY1vDmPfQ584cXr2i
DSgAAj1sFwvkAHOM12j04Nbq9PL92882CQerUdhdXU1BjLMlbsr/+DDTb9E+zYDGNPe3zTfDAucI
DHD9fEwnIe3ebjNiHgdiC4qgX+2//gJ6ljSLg5b2iTeEl2VPNtqvAGclr+jmoL9DV0s9k8MHfYYk
3GejEdpn8ml8sJ07P95tzDGiieHUo6DON+8up/FWY+ZOfBwdiSby1ryAVCNbpGAxc5oL1qzes166
zoszXSGQzA+yeleAk1oK0ytN1FXvhexKLV0FNsVFs5YbfjnMskJv+qg3jARNhfL3UQUxDNw2QNJE
mFvaRwyP12OF4T+B0T/Gw/pWInjRW+WmlW3CURH9uZS/viNFuF1jwVFs9PsqJyEBCftsZQcVjOF9
4mu6t3CwYR3RSvt8etDpOf08EUUp/jrFqgis0UDDLf/cCHaaeXgEmRkRJwB2SoCFDR7QadxWMrA7
eIo61u7RtJVyxeiioM0eCZ2xR7JeW4RLypwDs5VIyxkCn8pZ5h+gXfX1bRB2KeTkmpHmqYRggswu
/NDrRvOnVC1it6XIEDWyJo/RCSWJkHisFs+rhDp7u3AfQcJrUp4rxmBzw8MUSOGgPJ7MWQajXcar
UAGLBQNbZ4t7LhvyEKA/RZ4gMeUCvZKiCMRC6+LiK5TyrsFBcQbjLYFrjQ1ZO3mgHHoyi/wWcBuO
Ue5KJTC1DhIuLBcad4OAz50BIWplWk1l29LKybAmtI5oDFMAV8anzp2+2fW+HZkrFO8rIuryQoK9
kl876WaFfGcT9qiEMR/cWF+q/m+F+0BkBae8wSFN4wor8ozpdvrWFECL9aH+ieEgCC2+ObjHjbuC
P55E2Vv/sWo1AjCEbZUh589Micqrf/QXirItqplMrzq3JuEWarlT+5sewW7V5s8QkSZyePh4+QX+
DvrlhOr1ZtmSqUCOy23bB9SY2Q3pvqKor4OsutFmMhu02A9xU7iNqwBZTIO06Ketg4F0WWrido2o
Af5mylw9aseOauD+57rMgDh1/QxiCMi6Fmt/ZYgVQ2nd8ykff67JJ1jrE0NFYQ6tjbpseTwqSqlB
mRMEWuoRZdmT/NxnHja3qOwxuAenmn4JxJMElktBF3fX4iQ2zLDgzfy7Z0D2YDmlOf+C8mGHFWGw
v01vWRwasN7d+ctSsvW1AAZyTJdCtFVAqlRWUnsQW+gV7MNCfBPi5z3NgG3K0qaLk2+QKzO2qEwz
MwUC1IJA63DOqcQeT1H3Kj7AS91vFSU1KgZRIyGEkHLsC0ihUIDAzTN2t+jCr+BCvzIgPMDetyK6
fYujckHiuYTUDfFlhaRyli58KTU4D9uPMft2+Aa0xVc6+ejTqMe0JT0HE/FpPgBAjJUZdSELpP0Q
ruoNjZketRPFGsQbMcWD6R97WYFTtWZE/BAVN7//lJT1+Xu5bD1wDQmJ/7Wu1GmsUtAJohSNPHI7
ksD8YK8Rryeyh0zZuIZ3+z/l6dgnQKOvk6mY4478QGZbYplgTD9tbsTGJitDbaxVXYfnX5IxM2fa
1xEKU52U15PxDFoH5N/VBonJXFhPGZT1ibGqBjvkrA62877OBLxmTGiAAaH5lJgepvVjqtUYCS5E
06XWPc+MwhyKSSyKzY1V5K1pHGxpKQuhgeF4CE1TgAFn7DiiZFH4j72Rs2GxdX1RreDXe5zYK2Ma
DySISabvoXqVCgEUBn62tvTRfM3b+vv+SgrLKTpkbEm2jy3rEerbH1z76XBka/bNlhLufnSrgKiT
aEktNPSv1TJ/Q0KtTmNXkayzIC7uiQJsj0yRWxHUtgBTLo0J9IXNsWqZluLyB18fV6QQ2NS29W5g
1qbntJiQyRW5QyhU0FEdlBUFnx7B0TTidw56QH8AnaFrLSt4mQSYw2CHp6fs6RoKYuLH9IBMfTq3
N1gAfoaYw9BdRv5xOh0+fjRHl7+O5A1Abkw1ObupEjm/v/seF97MyMFDqas1c5xQUEYY/xhiimqJ
MnJsCFEaxlL+4jNxDKutJU4ztxnMbTvb0SMkHI2PMttQ64GZdTX1/gqgi6f2sf+Ptun3//92M/6P
Yl4wjQtX8KLV8sO6Mb26+juXP47i9/vlRsDe62STrwzPsWWwMsRi1KlSjxxpjc+gl+de+e2XZhyy
sCoIaoO2vwNmkFNs3xDimLg/77GYep+1tJVgUqSnXNOZbrlYb6s3fMIHfzrn+Jj7HNYsU8Wk+Y8w
1iqqwwI425eygeivZqXgV4ZI139VT2ChyXmhKhoN0uwDltD+DJTiKvcZitpNXGp7p0XtO//sN9a2
b8dmHXpJRjtVQN95BRYGs+qtGSHvjemOIZpgF71b1fmG4ea+2ThXIkFkk8eSikgKdmacOjbbSp9T
ZZf5azJ1CvhLYmigCs7Ey0Wc2T6Sy+0mvARPkHS0MyaEwEH0bJ8FVRnIVcFg5UNCYCITuSVoewvA
VO3p3AK/9McG/a2kwZYWDauonVr0vJ4Qx37qYEgN4KP7inU3gP8PPrijKux+n2njU2q4Tei39jpJ
XXMisrv+KPZk5WPpjxmEhipel+0z506F07K+9BbiMzyhAEaIid65FF1PGewHjJg5oRzs2sR37EAV
L7z8aF9GdOpWkKAro2mpNpArNhkJVCFtEcDdVvcA5dQ6l8Nlv5EGMqP9+RAx7TslZAK3HIkjcIBh
/nI75B052L7uByzBmsEkbYx1gGORTuRxA40MIh/Dxm5ZrstwulT5gGfRGPGcQDT0vR6V20YXg2UT
k5X7+w1+wi9PGxm/Pqpb9cF/ZOOC7ar3Yzr74tacuiqmMFxakugSdGpCevV6vwr3l2dyRh4YSHa+
K3bl0i4Oe1yfB/45PHcy4Y07Jtj5lqkItUE3bkSiPhtHtoPv0a3cY9xiHhIzxc8LqJe9da+cwjOG
tAL2R8D4ar1uwdgCyscbjFTAMheV7zzZZM3Sio1o/v3ghcrtp8NFeTrklVfQECJdCBP00gy+x+jp
8gTNA96vFG0IdpiOPxpW/7PBPatcOvyC0yE3V0Z+ZS0+AKZ2Zls5QtyLV6p2IxAAZsQ51IYSLiQb
CHniXg/gxmy4UDaj2PhnOy4U8eV/hMl6zVg09Y7JlrHfBCZHY+0TcOvn0OsYoVJtWw7HD/9ojMHS
nTBI5N+6PIVrIUWRKLWy+AtFw2D2SlNLz9gfaMZyuqNu1obsvWZgdmDaBvNstUsKQqwNyG/+Iki8
/YtQ++ZhR0K485+cdq4tAKmoE9PDwYmm4JP0ik4zB4fmHhyQtyL9lBpenW3VHAh2IdHB+ejFvJ4j
GHC3vDdc3eb/qv/bU0uVKezcA++Y14twYm7xUVnigeWdpZnNeNj8v87b9+Oae61tT7RqTJIYpbre
CKwW0a9K/VtEoSwS/GJIb1V1yVc3RWunjuA+uAwa2HrEAlyDseJeh9KI/SoxUX8yyukU/20DfGuO
W7al4MxbAFZSm81V5+FZpXO7uPaEsu8tQO9rBp+FuQMRgdNLxxNAL/IzMjBrkqjFHK0fWx1DQ5o7
R41lOQVGYeTPnGXQEQ5lUUHo1SGOyeeWF266u6QKBCN9idVU7xInTAl59iV3iQwOGqzp87jZQfta
epewBauD6rpQrkeZKBzt7ldTzxHHXD3+ENi5F74esTAHmMn+vDIgyiiujs1PYDusJRbzoPr8DF6Z
iBK+XYymNlSlx6Oljrt5ZboaFCMx7J2DCNUALfTeOxavfwcJ6KsOXb1w2+c3xJMvUWxqmk6QPsdn
w84vEFuhQh4xs6s/zkQsIADL2yb50MRth0a9hlCV87ACLTrelaBczxefTuOngwGsTdLLiV+gZuw0
TJRX3xMC+weWbOiZmwQqUtM4LG0NC0L9BRARwbDTxaKI5wwyxHA3GRTJ2ElQoBsskWnkRk6NcGdX
goQcNtWo8CDCBqkpEg6+ZHJs/jmjFpVendCnG/wFGIlENbUSTn5HnxOqskuQY4Hei4LwXqRjD3BW
XxsebBeLgA3KXqFATlQXikrIQmaZQk3IaA7hlZOfmM2sWsmPY1+itxPNQHUhweuhTF+Q6aMEr6PC
LnwVZKOxCtwEWCajHX49GmbJbGEq1mkE1QeXL1SLY2s+lSW3Y5TpmTCGfE5BYOkVT0XOqd+xZdyz
AORXTq8uWx5f7E8FnG5VJzAcAogzxywzng99c0lhNQhyLrRxSJmfy9LwRNOzlQ6JnFIEfXDX8hgj
T13vwsSsvSLWJR1WtDX05rldGVtUct1eF3uF5dk1LuytHziJNAUXjqFIPVdv3jrj5TFww14uu2pQ
wH8fwx1OeQ4vxMEjn97d3NFm/HNxo+JgUmI5o10WwBQf6QgwzGUMKGCAB9XXgp9q3CAPrVvHaODj
JnFo6LlCCHZIviS23Vzy+eWySycW1iV5Rezyu+dNrSpK3WTIi5fQep/1HZTibOF5j4sYB2COt7sW
W34h3ya2wWA1ezQaIoKoQW59dygEclX4Z1sehpBwJGa4BmcuXYvU3z6tIZBlaYil5OmVY1oEm33m
h/t+ZFfB31yIHhouZJ5EOfcrnpnLmKmmL5bAL22XLsiRQJ2jK8yIE8Bxhpix0ZXGQt2RP2TLWg+c
AgOZbd529oK5MiP6UpFX5ymfq9wk+nXaoYrWJvS11KQKo6B0r4BsdBGqXfCVKBKyzZsKg5B6ucVk
Kp7QX5VqNDpvt58/UTTtigJshuZTtaLSLnQwA6nOOzg0j4XWdAz8q6HtkrOdyFrCMUWfak4v1wll
JnyuQHZjaBUa4TFGsBQedKkj/KZEvAdMy5+46nb/NJrpWvrljHIAhsBtL/LK8bijVDJD9Q8jXy/n
NmAXQumvOSQHX7Iqq7lWm/kTsYapj3QvV7G7FpwlswqrGJ7/fX9Ef8YmDlc0QtlpYXkr4/Hflw6T
dqjPkKDFA1DukmmhXSQ5bc5TF9Vjx2srq8zOUdxUNDiOA+eAr6SbMwbRvykly/N4W7xFpLiLAQ72
Z8h+cAA38a/ALekjLE2ARqsoFUtgcIh8lkONkRfilUxX+M4AxWHbOaQrgG2Oti4ojon3z+UAA6/k
3md09/sBsQIJewHbmTJRpuw7Hwz1j9d6jNM4/FuKPbvAy/wzdrr824pnJzyB6yP/iuSa+084bynd
kzvVLv1y9S+iW/bXp9IBnThfRMUIgNUISjYdjy3/APf7ICs6+96sGWdvkRdsGG/vWHzb9GkpolEy
csxKovFvnXwuA5i/eEedBEof9GO5FKYBnBI6Wk9cqShmn9M6FO1mFOfnD3QSSSbGk6HfkBJC6EZB
ansuVE29/GvMnvqIx4jfjzcJj4IB4KeSiJSBeUK9ULf/fRbEMjdgYOgD7Zj0bk223qV5D3xKvjaN
VoIsQm0mQzRaKG4/PZavQ3NpX3ZLzUt0T6M9way2D3On8u1P2lvNNwxZhvW2ia9WGEUPCGljjT4C
0seZzZdYFiY9cBUruj6pvHkmwZ9fBP+p1MUwDZeDPreTeJjKG1YiYYw+5pxN7GiFiVs0WGdjJP+1
zT+oS4Yl2z8NWkhpcMF32NW9QL/OIqZz38nraPaUvTMWUlrL4AY6JDUU/KIJcImkkiLKJTKDzkxB
acskv6cxtMh5XeTUR+LjhPYj2ns7cIK4XEHkenNb97PxUn4uuHeSzE+KUobzssCf7d4iPU7IsHO+
TbDFVH1m7sP0iPqmM2RHwG23cpdma/jlAhpfmPhUSF1JvAAQcYQQuC0QjfW74/BHPLgkboMSeYfp
n5PTqDk04eAIVsfs4dxSNLHWa1vy+0xaTW+IFujOnKhw+kwEnaDom2YSNgynaAvk41RH0O4y9u/P
JEMMXJ/Skm6R70uWaNdP/oWQEBCkeaz5zPy10uoo5Q1oPK8+UQ4PziumcFf+2VcUCu/Wxzhvrpv+
TWUGrgQzrQz0m83NZ31gSt/3napx2byq4XJURMS0/hXNBlBDC7cRTR4gVTBeEilvQjjclA8Df0AD
Z7VggHdJFhLKAD0ahtQM5IsjKYJPkY4d0fuXE1Fg275MjY1nb+H6cW4zBF2jZt0a+I7TwJyJU0EE
n5i5F+zXfMDRF/n2cDVv3weyhlFKcFrhAyo2ImLvVNmBZi5Tn0VsRNvXH4LZxJnUBUrzUms4xClA
YH4wpAewJdqKBb/INlJ+7C7QHTMvdtYSWoakK10bw6JIK9w5/8mf4lCznsEyNfwgfiX/j65qR4Wh
f8xJSc2b7TAfGvxsFwBwRZ+NeKLggNqDPCPoZzjpI9s+69wZ1us2WLwbfzypN1TnHRdNeR9R5KC/
g27J26W1bYRmliRCv4abKDZkxluz+69AH4lyskMecyLzKf5UGwSyDislSFRhpPPenN7ydSFrmI3Z
TdUZuKzIifnrh3IZMRfRbyiM98QfpI3DpjHigOZHOQ45DWGAw9RsSTQkVoTvH+tVhKKBh9+XSR6P
pPgEbcLZg/A6VsWk7omTZsuEgwoPTZXdu01XRyAT/QbxYWGIM/r8HgbriH+THqki/7jMUYdVEYyB
76Ds1c5/q2Ozm6XPBzN5w+Svq88DqGp/9bQJ9evIkAAVq/IwFAviFkFe1eUj/oP7WGShMPqkZdO1
BSRPFX5G09aDRg1fS/ek4s9G+1H0TqRAhtlr9BrJzvRHgUlaP6PUnzgk3MLMW3ZROakHzuMkVz0L
BxCd9hhzcM1gdvpn72bc+kX1h2nJ2VEUnqJ0pPpZmjS/LyqXJc1e+lyknk0aLEXupmdQ5FdASZ1w
AtTKL0JnNr38CQjop8pwnv6KLRXgfKYDYFmfrZmgYtksppzGKiw2vyQ6XnHCNiauhg/IICfAyrLV
MbylTbOG9x2m2i6vfDxE4/+T0cPwVGje9Dhdn3KA6RY8qjDKVWe7SflUgXk5uyp9nzf3O2yg/JB8
KusocdAe/ASx2vekCE26/X7OTbJvt9soHh4RKtTNyinnoBbyfBQG8O9t9xbGSMMwbLRdEpAJkast
lKj1gUXEvIE8nNeG3HfS2L5gXgGKdNn8zaKZ9WbZh6SGBGiDfvcOKaXbypkjY0T350iwoTzHtWMV
jNmGVtweKIbMtbR06sdaZvrDDfhVtXook6l245D7oqoz9wO3+XL49y5ezNWMln7HIkjFOQ/VI7XK
4WIK3UNFBm9qzrApM9SdoBVLgr0a8vhVoUy0ZG0DsPI8yObMBqOE0mBOTk9w/VB9LaK/ioHzWFW9
6vs+hMLiKq+5B6ukgcd+ZbUqj+jetBmwE4JOPYtgN8o/xI2jlFg21A0v6/2ZdKglzMQ/kNz5sDsP
3DhnxtEYn55HLHkxnLrrs8DVmqmpgrkfJV1oowBijWF7ii7nc7LjhYiKG/sd0FPFHWXEniVBk7Ex
vXeICtfbHocqQCvKcvR7x+j6GPsRsZlyyqF3ERDchQpaF71lCdheRxo74ruOt1VNeGcb6dP31IJ+
xbvqiMBBCEKyYFQLM0Ool8J87qX9OT35ODcDKBJMB0X2oev/vMLEGmeiteVMD11c0Yi+9Rnip3Et
R67fVlcEfkX3VFNkDV1wX7KjcDT95eYMOthH/OiNVIYIY7fHfWYWeC5yZRJYIB4tDgByKOQmzRFq
CFUxI8eDb3WYatMFHoQpW4Acm4fdbHYW/5cVZwKhuGeCFiENd4LU6bI1dy7vj7E3FY27tOB9uYEj
tO+lHeS1PULlZCCcd4tbuemo+H0Pjbb1JqV/i2/fHPG0Kk2M/bq6fH3FgMWYw2rGzc4d0e23Llmo
nelzKzWHX81y6C4PZBH5/S1i3fMimOS+YFKUQjGpiPUjw9HJ5+f9VhUh/6GpAojglRdqwhERvbVk
JZANmGPPS9X8DFqJgSqpTW4BnB4VpwHU5FlHIzbx/YTXlC6VOhodNj5szsaj+xSATQVIN/wpyuqZ
gbC7Fmckgz7EpLLi2PZiu6bYzdRMQm0+si97RbVEBaM1BkWEej6Ma9vOe14LTF29N/YvZ3UKEbHW
xjXxGef1AFtvJ4zGXRGph9uM/FPQN6N+CBGRDxYtPW7T0egLwk/XslSeJ/wolO1DjXD8kWVf+vMj
jrrsauOXbkMva87N7cmqH9M2721NC6VBKM8R6215tLasomz3H6iJlmFxEmlt79bc0MZuOZYH+foL
ASdsxjFTajQG6RgLRRAS0Jyu9mxrPTVmZ3I5BFXT7HvW31ITUhW26yWixeiGAqnp1Q1yxDNSKWrG
HyLDbIPUHxYfSG77madOwQcLbmKTGieCZ06bCVTxGSyLatGhfKD5+B88TR1hYmN+ABC1bwlyY3hB
HKJVIec5A2T9nGC/pI3b8yYLXFktQPp0kvhouFxBCZsooHATk6dQMfMhYkciE4qxTk1vPXVR8fZG
F5a/2gvDh7tGdZxR2AC4n6Au2fAQImvvjXq4DybSmo3Xouo9uOar6rTgYubIXZIlJPuCWosrXzBk
1i/sR+bsVYVSwfLPlfJ+0db6XksfUvk1e4lu4jcQciTcm2XLa0KJJxiOAbRMssDkawuDY/PlWmpG
mAZN+CS+CGDeSgIu2wmzTIigQ+XI0uWPpHbV4cOIDuzEe+cgWjQdeBN8i0IrnrvQyls7sAgo1t9W
lKX5fCCPNhzeTOlekRpa11ReIU2Bypzoa8JtIEET2i0ko95kORi5VGkn6V9pywnmKWuLBxCTnw4+
96NXlrsXZTwG/I02IKh/TTeFq67ElqPrbsABNmY0TnWX5a70BHe4LFXcTfDaF7pRzip6L8CmoVWb
fQ3h43NzSCBja/Qvm9GmwsUyVJdRPKvGx3Es6HG6s0wER6afcNzxBHbmuIGwTH52CZ9t94hKAVEV
gc61YX/9xZyQ+Kq4vq3TUs7zryTP10f5zoH02ccVjPM0bfXSHPrBdo+l0qtXFPLp0DmJVyZLOAqL
VHP55N7mfKvPhNYFEtYHUIBItQmS4ZYuNYbAHEzl7M/0FgyHsYcGjHRLtN6Ov5iZ+JUxyx50rfQY
VMk5MiCdtHm1/q4X9yQSRiv7kAbZwwuYCWGIGECi5SU3BgzBRi4io+CZGBIAynu8Ul4dgYWp+ok9
qVwSNPHjvL8iYUTAGFWFRYxmriIvfQ4mbueSL3wG9q9prj0t3e00i+qxP2z5dBAV06dSkhs57/tX
ao37XTS5F/M8R526ge5BxbuUo6zW0MVl5gSXyBNgE7JkFYEycqRX+puHRyU5LPEogZ7jwXptQfoR
qnGX3UmCv92wshwNT1FO3f9E9SKi4zZxQCH/kEjlxmVlFcXi0/tYT4CvR9BeWAxTtqtaCXxnc5h1
HFVSaKmfdtSKR7BSIHQdagfpxbhKjTxD9VU2Y1aTeTKWpEyqfV8X49UlpdbKPXNYyEwnBxZA1dAX
x2iq2QY4CixpCwgxzFggT3Ife5IYLqgXaUxZBf8KuEYECSFMM37CaLS8hi7D/hHWaSQKi1a5tG0Z
LDxOsNBH8aSZ16Pn8OdKZGlhO67GqIuMDT4VmmEOTjL8UP7w/s+nEftkxZBxnwcMaw29LT/gcpH0
ZBw0toy8I6sgKAPg2234+a+CNB8gXkk05tasCZQA2NSEsKO3CstzzrU9N3vf1a1hUX9LsA/44GMZ
0x4dwVAfxFGGAlh+UJmwsQ+z2UpBcXia1LoNi+ovxNEEuQDP9AgCYIhpQp/nF9oTgk8bNF877/eB
PO/wRz+XJ1dMa49hRUdJPCp/mUhcILleZduXB5OJMS1ieEOR2QDECOrFIwzaixEJMGq2gaq/9s+I
ab7LntFmNGGTD6yAIMas+bv/0IWTbviEuocYSDTUCWU70ZLcHzClWhR4dj78Hbybf9xQaZdZbAD0
Z7u3pM1pSRgqfRNxKQht4iPN/whSC4nbTbYmh0zC7RZI0hdOU1pYYQZxsGVP/1nkB6cSUyxh7kn3
JRri/Yl8UTRukT40nqoHLqqZ7yiD3MmiWf87n0OQlZy06htizXxFB92eeW3MlwhZAbWls2fNGUh7
xMC0yO/P+PjFpFlH0ZubtfOL5idFjzW4/2qJgOerOLRONPPk1axHrRmQ7D6BOhoBs9kB5KUSVsAa
p1dbuP5dE/fgq/fILBKDxyYcsrNUPj7ovhugS6Q+drsQsDHlRTh6fH62XqbFg7902D0X5ZK7zIF1
no7gBIBMgKDaT/1mkfjlsgi/OKAVbyufAKfa5glVY2Yqt8jeApoWNiDbgWn7cZft2NgzesitRuOL
HbtrJ9r/2HWbgJ4hRhnUNlmNP5TU9bg/sn63OnauJHprAc4U4UmnM8LhH+9dz9FCXVTO9pmqeJE3
cUIJtZbV+0cTb8G/T4lHDL9eipjr74zeH80zcA4iIA4vs4cfjnbuIsOpQwrq5w1ALJ6VnIXp2IuY
AmTXllrogs+FbwHaHkeAPUnES/xHTIeEWjYZVoqJffurwAH6wsHN7ypABX4FO9EvjUnj9uLYtPjD
0o7hhe4rzbrdeycyikIDEU5yAL5oAZd6/JJB8uxEETCXboYK0LrGhIqG4rCix/qnbXRaWB0dOBeG
iwxBf8kWOk8ODwwqTa0v8cOL0P4bCdwKSsfMEV1ZxxDRAIkPd+MmcYJBT1wVecBevOHqe6lScTK0
bJKUDExNGf+u4TjHaFzg2pYbD5C/mYWf8AGjYM8/8dcZL7+kj2l8hgqTJPEeAK3Q0L8ZHeirahWu
8tUjsDKSenKys/12XbQ6hfpUnzSz9ABqQGpqXhXSIzlOXvMCFFDJp/h+E0hYKO9V+0tzXRHUVFvo
I5TtpBi/uGZ4Mdjx1E8cdmffyvrmgI7WeC5Cb/Wz2q6va+DArzbhEit5rJbKBh0e4L2eGd216RQg
Y+gW4seoO2mlQ9sF4xaeFL2hpXezvIAobM4EKVTiJBQgITreg6WW26DCu7KdW23r009QULXr/NBJ
at2c2yApBUp467vKS7nuxwi91tWxfDy0L7JyQp+wugCtN0FDuky3Q38O4e8SVZdBXvqAwG+BO1w5
iJ00/80iEAZR+YIdh16lVx/QHqKisK2GPkePYY4wsnDzH9owz0MU9ZZr4GJnq56uDKpXTyoqPKxZ
KYbIIwO8l5u8uZfkogtIrXTZ8IwXGt8gxb/KxhtRDUaFKo01NVAzNeCbFmXcems+WySGaRQ5dLy/
mPouvbLWs1TchPyz1OlExebn+hBxwtutiKRJTCdVgbw7S8i+vzWfO92q82gh+pl+x7MlJmHQQPN4
ltg9QjznPa3XWXou1QT8T109C0LmLzMznIA5+RD8uFdxkhyS0W+a07eDfHC1zx/XLomv2vIipyPf
lTAtMAQdZdiCGGDfy3BEnv9pmmhAVEEfgN6mu1LVKauKLaHocNKr0m3obLTOL2MvV9cq20cykzKc
6h43dP8tVAUE/IfPjq21KdjzIuc3vHlcCjwegGkzh5/b9lOw/0z71OIzCe6LHust30gzQc2tNo3D
cU/DUV4HSiZk271seVZvgt091H321K2kqS69T1yv7ECZD2N3T4gLdUz5Mu25oneZCDOpqs+9+nBL
z1AV4stqUy9iIozcsHIbnsXIo4U/1pLUNRQ0rCQNXMdFS3nJoKyy5nXgPwy/L81xjhwV9fFyvjNG
PWVCzHED50EedEac+aoUtcK3R4fPs0vaJYIASLhfQuPdtfF+StDpizkbmQKA5jhhUOBYwAXjob3m
XuecpK7/RsuOYDCzDETbVLqD1IcxWei68NNgm4r6QJkmtvib87YxFc2scGCG/lIVq/l0MkEs6NRI
vkesDUDaTpugV/t0kxaLe5P63R6iSei80G5Ojf+dTqfEuWWO4Sqcn4Pn0D3KZ31D8JqDG6pzPaV1
tWac28/i9T20Zio2Obf1MnQdtRukcP8NY2inPXLgU3sDfrd0VkLnQiy0MRtTYmfajStzsBMHMCx0
UejcfKCLjI/NgbzOP8ToLBOiMSZDMmyLxGHj071cZ4Boxbp95xcrPa/RdfBIl4AaPuLn2TBrKpmt
BX5kG5qHx86fR/Wk/Aqr3OoTXVqrATVwed9PrIdqYjQHhyyr3/gPcMoiE7caUHrGTfUMmZcHLsfi
HpwC72Vrsi25xLSDD7qEnngdE1C56bESupDDPYim2498N6apCEP3Vo1Y427JQjEFiFkouiqt3xrK
rpcAyHlOpMy7GSfxgXkE3AQP/6IZVjFpt2DVFpMEZ9ZGhEnlobv6NKD7RHHfeqwYiAlVnDvci4qn
n2g9KeDBJjcnR2A6DDCdmHdJnpg3gEScuL8vuInzCs44lvAK0AOZj1J7LbGX+IbuEmh1wbbuazB1
djAozYZbEDPkp9B1tNvXZ4VzBjDlOCuSz8RT5DeuFJoaMZeMY03hKRvTLeQZFb9kT1NoAgvKVoU+
wZtztB52OOXvbfcwzYDuekEdhO+6qxcMA0I8J1VX9JY0Ryz4BK9TcoesS5VEiCKmJO1PNNxgYi05
omwirt5dFgRqAXiS2RDTYu0BGSYjeeEF5tBOwl3A3Q7a0p+MxRiDNedl25fgN9xwVasWzG+QOBuK
RYEFnbzRHXlYNIdaXyWYKY1SID0kiT2NtLvN65QbM4VKw0F1x+9cMCwiGeycD1fkokBBKGDGWIeK
S+H5eYtzNUklagtmOcqeupevzSeQQUdksg9cKa1/mKUrTJrD1y5VW2hD3YWLk4OouolH7RyevmKY
e+FzVjPb3KrrcO+hTn9O+FIgyK+UD3betUUPI+efgEIKxJPd44w+sfENbiNQOyiCXrIvuM0pP7za
Xv/cBe17/RLeuC2IX33iGcSPX/SCbHkeqN81l4D2PnY4aYbhdXbX7Cf3BDvULuiFkCqQG/DFXsl7
r6yCb03Y/Lb1VQK9eWHRBJBWKQ3kltxEQIfaUSrcvV41UOrhvmO9X1R2cudVcW/Jo9ehHHp8eT5S
KXvG7aTcY/NzXQNUIQoNzEOzUD2biMEgc4ay5Yr7ZxBBYuejdgVRcsy2O5Ld7EiA9u8xMr5Fg0yX
eYyeX22av+c0PFyzPHVA20a2Kw/FDbZb3Nzw4XDB9eUflh+bWI/57UZcZ6wjx1yxY/LCfFqFTGt0
QF76l+wd2pbaEF6XjTd3V0ILqJN6+AewX8PqJ9xt+X073bwHcgYRbekA0P9+Try8fuxwMEPL7kNC
6epenTvBY8jq8NskF8QA0SDMO/d38JuJc3hENVOtpV/AJ/rC5JwHqsNTOUEweQU7f3MOB0Zd43H0
oWsOSwwUCBAYnPYDmAqGOLk010RTpLyxUI6DiM7HsAOpiM+BBc76Pp43SSbvUX7BMHWpq660Mp7W
A94hiEC9n0wKf9c6K0XSm3t1+FGiHykF8t0CQnxN1/mHIwTdNN1K2OO4HOs8fDmAKT3288X4ZT9R
kBCz8+npCQPcreX2SuT+DE7TdsJIzqM5XSNBkWbm34zui2Gv8Fp7Q/ubhknMnCeDz4hb5QhodVrQ
Tpn6ub+txqJ7w6x6Zx9OMs7pS06P+Li7R0boyqtlouimtbSJlKpFK4ZU/CTRNYRoeG0j6+lb9VWo
qBDsDmwFfTsHgoop+RShUVvKdxIet6wOE7klgTB3gqqOnzauwdu8dp1SlQ8Eoy//N5tklsGzKiUq
Anws0iQwEb/mMpor+34hCl7EaU554fB+Au+qbGQYc8qETwMeCAEv+rXwlDsIFTjkbfwzOd0eo55u
9X3kFo6IVNGBsFVCd8KutiRED8AKWQVFZS65U28wGt96/kg95+bM9v6KmmgJUd/BEbohEOdGcMZ1
vsUuXdbeNRua56vP9HJarsf4JkTHECw4Vv6sJdZmWHMawkGgZUvgzP6YnRHzA0MoVK+bXjjYUfDZ
LasAhLPTClTfNKR07cTRW23AJZAWLQmXVThtegrs0WjGh8Z9Itf38vOvJ8O0dWpbsNHlKtxC9tRY
NnIi+0+sQT2mZqKjiKGa66sdgl216/eKCIwdlUAeF1S06ctEjmT7Naw1XopuTDbK2d4QuMjbCy1G
wI0L0M7iA6jO9Mtf8ttEx+PctLzxyekvWS04MpXG4LE4Q0b27r++SDw2f0vhxbiuBJyd8RYbWVhf
xxgaRlv25O7eb1VpaHt6bEvlIdcXlk3W3D2dY7trroj1QOLgOphDyGhSPdb9fapMudZA3JxyC996
VURn79168elPXf+21vs1nPcY8iawKsVIeEcT45/aqMBPEu8ONBaY0B2iCj0z9dBXIsZmxXKMDK+S
jl7XnD68/WI06QBHoUGh5m1EnKKdwn2y8D1Bo7pVEMHaDheA9gdHkg1yMun3SFcgUhAXr1K6oPi2
OwsVkt0Vdmtbu0pK2/DgQeNU0xyvdRYWNS1m29+LMtVseqaVCm//DO8e0knYCL3O+QTDV++3xe0g
eNvtcI8y3n5yqRF1dOMBcgJ4qkQPtBsR4yusJ3shue4hmkmNfk6uABNgyFEHS9PZ1HXF8dHaPLgr
d41xAUqUZJqmTEiLAkhHlAXyXuqqXycsiFimZdjErgHk69JVixnBr//tqQJdJMXuJ5SXpwUc8idu
r/FHz17GVwv5L9HHk+Cd2VpRaP30mAYC2MEm50JA2+7OjgLrJJbjmM4z01lEbB2bHyms+0+14Ll+
To4n9/sM3oaOdsbvGNDcTQJzQt33j/t6o5nz9LOweCNjcCEEzOkNCNjTrd8YmF17IWixs38rXUF5
QVnYbLb3zagzjzOgykkZv21Lwgg2Cui0Ny1aIzDQcfM9ItUaLYvWl7hgADhj2lfNu57z3ZTp2TSz
JNBKTGCIHuXr/x5T5Rgf2/bGy53zFnKJxXeLSDWssaUTENUjjmRb8nxiXt1hVZHTOht3H1uS8x0F
5I2NIpKCc1lspD4ox4M0jRrqdFLHRsZ8AycL7L/jV4lRCppkLNDOjfDiXBXqm5n+Q3WOB7jamLto
Pt5cFDhEM+g4vpjFj3q8PJlYeHcJLLAM6OMuhvIfaBswW9EbYik9T1T5NdUpUzjG2E9hhwafHzu7
Hroim76wdR5Gg9+BCfGT28rlt97LeHGt5rjLDiL3Xl5LoR3bG17nLVpskLj0TlJuacvKLaRNKkXX
v3oHZAWRb4F66Ji8tg9fElZ5iJmxgw3eHwewAGZScitzHjM3wNaOco4hgIm08fXVBFr4og7ab7rM
X/KbRtsHjVO7oRVXOqrI5ziCmOoIgTf6OBnjBoPCkZUofSyBaWtt0UWXicWNzV6jhJRwwksKNXSI
FaSrn00uMjitghJkB2Y/EKjnWQl+dpzT0sBvfmDTk7tfDNVJqWLpMHVQRVjNXO99cnxB9CpjvPU6
Z/A4jvaXnPaiYxwFeRvS8eLbRjNWkn+WsffDJJhunnN3EO+/MZs5o5W3mCqRT/WJ3zlP02EabF6t
VlCbBq3sD0E+RxljUQ1qSLujt/t8n6whyxF77qy0sBP+5ALENiXE0aKWlzx+wsyfLJbLjNPt8byu
/3FSx3wVdmIOS90WE0Gn8FgQGHUqvav9lRxpIPxC6lE0TqF96ifIElxykHrHdC4rf/uligp6vxfh
qP2W4jodOWKJykEhPE/anr711Bgz68lLuvhrCzW7MClKkXC+YR5gASDEJOL6CCMIikIl+WKCtwCA
DWqAF+NkHggqAskiYMUUkiAs8EsjQ4UpeTOStVCVxajBOAknj9qzBwmP0IOy7WYMIVdIX+xflfIv
a5uwF5kDINi4Umge5heCbkVZIvz+Zle/dRuvCGMsCDQc2OIFiHMeUgMWVC8VICxFC/IRY/ecmLkN
+4YBq78z/fJojyd1dQdTstCs7sD8KnP3K09DFBpMl+5zTNeMC6Vhuk4/DiFzGq1aR+6f8CUtrrmB
x6w0GPq5yRcBEtTQbX4eDIzmq1GzciV33Eo2nHkwIGQE1aGkwSebYop2LxgJNgnPQOQmfZBj+6Ns
JxN/vXEYyXLiL4ESyqpJfLaYkT5RMf16RrLPuMAC9cTscYJ4771ayOReRlsAQ30NkpbBqVO0F7xc
ZhWvfkY05vGidyVKQkYtkmUZObkzenqas+Gx64hCTHA8groEb9FwRbbE3oKknHxVTa9sewjzzF5z
bR57sVS1Y1zmhfuldReskMKLNBcg0w6aPPFR4UC5pHFnorgmU7JTcFycrghJf+n5mLAoZ40kU8hm
Gh6PhBPWahys+sy697ZHo1XTr7cGSPwXw++1g2bxyWiLYiDNib60Ht3CwSvemYxAkS07N5L5RDtg
1MbKE+7aAixlcMmhfsiIEpwT4kVk0UAze/4y3ckNAD65LUZaXr+dPRW7dhNj7AEH3UC2R6NF7jY9
AbTDBVPwDAIhz3R7L7cjZQsoEob43DmXwt+E3UsS3BpR5x1CuTIq2wa46XPX5WC4uVDn+KYPlnch
5PZIEEYjwX05AgwaqMJOk4R5RhRy0ulaRuNhJPPTg+hRgtrdZHWIutUw+GM5aFayK0ZQwyBKKL4P
OSuSNWYEPZMW1+2DBA1wqMkBwaCVA9ZNxsYe6NLTpbpM2mF4ayuVvvrAP3+L7LLjIzltYjD1kbO5
h8CmG7Au/TEY8ViOW+MJl0MKYNn0EbDQ9okTDJFas077qAm7A/rJLrayjtW6xwDSTSP/PPuCRHMh
WWwbrAPj2YtsFX1rAtmFMGVO6DJKnYaXD2MZr3NLgCZ3jx7fwZz3OP33kq8lrOC1NH4w44NBH5ts
Y54oMz914bvB/hZgTElCPJ2KjyH8PdcSL7VXw8KVqjAjzjzlfAyDCFDqoK+LsMzQGpBOvhfoFon5
Ivy/mm7vdIYSLa04a+4e5bxLz800r6cXa32ELAtTn569DTzDBsRjQvCkKftTK4Od11jWLuwWjsH6
KRp0FdU0UeTpUrIw2U5ZEPvEYBh6JWD+NBnQenjBa7Df49jI5WGbQjJqXT0pyB8tFoPZmfvjmvtW
/ZjvT+sjlH1JP2WwxnK+OwGQK5HsjAkYlPGRkqfPhbOh1qOp89yFbt68fYPuhhGcE2HDhjMgj2GU
HlxGAUhF261hi7e/52yzI5rPYquko993c8bxhV+VXQjTs/j9HYwsmHUjNfPE1Hz+rIumnzzLHAO7
gmMzZ5o6IWPYMpP/k1QxD71gKAzQP7RJyJc5UjgkmOB1Ta8CL8TtIv+swaBSQTTsVoAneN/PQ+dF
iWYXlcJ2yPm8Bne3q7KarC3EDT3c3Dv/PeEO9/PW7QxAmExXYCD7l2AWEAomh8vaQtV6GgvqI6xl
HuKpdgUVu7STb4InIlt4P2QObjwfPEpcZtXepETFVmQlMQVSCZYKI3j+l9nssovMYTHj/xiwl2IZ
+T3O4CUGQjPOsCYBpSrq28gL2wCNjor4J2+V5tqTDjht9lVHH4DlJMtwcbjUQMEHJtOqNenS8l8+
DbL+Rq0deJGPr4tfv7fwJHThY2ahI+kExId6WlFV/87y/c66Jh93p/YMQUfEKR0iRY1aAH6FOTs6
7uJdTeTenM+AOQSGuE1hBy1aZZWtHXMJxG5LUPruwY2NetjrHUvZ9ssSfm7blrZ5sAwjrXuKOsGU
quZryHIG95ys4iOMW/NWSaOZRFDD+6lnRk0j/BlJhGTS4au8uUE7tbxRvv7Yb9/K/Tz33jgzksQr
Ay0kN/zEvzu+zK+MY5pbnyHUz+07FhgcVjBgVXMTVbmafquL71kwqdDEbVvjGhd5tkY3mgUiPH61
pHWpyMw1G8Qy2Pu4wy7jjVMjcRBIKSgzsQcZcBlH16rIEkiJzzMAWMgfLQEqZnaL3VUERpHhjGCi
GE1gDfV1Y67DyMNrBYDdwWAmWTbCIfY2XDwgHAEF9pxcTZGSYi5Z1UCu8F4Gbp0251QiVSOs0HGK
qDA/S++T0Lm10jDK/MmBI+tP+RsH/MgO31MBJwWwYQM1t5TdSi5hEaaGNxKWQ7EBZu3iyQ2YH+8O
m9nDmKJfoipFsEYKmmm5azZRDW8XVEXmRtMK+LUuZgl15Xonv6izXDyhdk7T+XdlOykFRZ7YYBz7
wWbsmWRHUOqvFS1LWw2B59NIoR7QMRgm8QjmisTSgXBxfR7xH1UMLKZfcliUOreMEKpCL+eklxi8
h8RkWDtMDvGXXTWS7d+RvK99OA4Vsv/b+MMN/BArjEzMRKLW8g2oET9dHH+JCvZB4Zu5Q1QAOKU9
N1pJ8e2c1iOv+X71aTMH4wu2DQR24YYvZo+GRgS6Jcy0ch+1PUxTkR3l8dk8VYArZD3yTdBwdeyi
R5wJ0qAkC2fL8w1RIU3wiACAJyTlKdG+O5HL9hgQrTDthEWOmO5I5wPSy7gKGX84niZguFniZbyi
P1WhsTExfjYM6cwIBo8qc+O6skttEpImO4lk39pDhiDIV631ducVDFimjv1LhHRQsIHUb8L+b0ND
U0Iw58kB26PjBm3j5UJNWIF3l/gUrMuME1E99+QsTZeT1f+ilHRNLHHTOxGXhwB1M0j9ApxAB/Ov
iSooCmMtWaDfogza+9qmSivGbt+FwNWFSCfKNPhezsCYpVZdxELz5Hx0G4UcPQ9xE99hizba0Jm6
p7pWZnPzRbmQYpGurVQd3OcqZ85u/I3MqvJgdrwZXyYSBnDWM4SkfhtNgaXwUMLmIbotH1qYCD0u
d+y2mGIQX15WnmlntnsfgehWe9gf4lVzqZVlZm5whpRX6rtluUX6lumvuVo2i6YHIJfxAO4LkUSI
TjKENrxu0yq+yygpVOYWdD6ZE/F5h1VezHuJjEfUwzE3+ma9h20vyXanqXzHl7w8so6OdrW/P8dV
oVueXW0BPGvJPPhDJxBhhsLMXl73f1tI8/Aw6srG+v/fvQkXJ3pnxY2FLzPf9VStrvaxqOiCvner
PgLQ87pOYbwwadzGf1sr0Cgj1Oxpvs/IaOMcYovsORVD4A5843xUQUCgIC9XRGXJIHTknF24nU5S
flBY9lWAHlG7Mef0ypYj9k7TPeSmx7OMZPLTvxVJsC+xcHfTxkej4BpDSt6fWzYQ5zpVaXRBHLmv
wXUy2CSxBKnwcGfFqvyjxlFjuHDaJ60w/6oRPBTWS5+SpZii/21WtNWA3+WHQS/AVKRkX8R6fXnN
ds1g7X8iuEzHbGQouNRKD/d5QdNs6xPTes23VyTuOkRPaQznn+1B9Vtns3juadi7VHv6e/AUDaqS
PFn65dzc1vVVajTA8Afw77jwXKxOXzYfxmZ0vLu42P4AqwoJdFXdokKvLPGgNnptac78z8q7R0nF
c/F5AGIfIMdHDYVAnrUgl3+wYAtG3UTZauQDiJfjVFO8BgZ8OdnNrDlwgH4YcbVGQklumjMDAUft
zwU2e/Yz4yMG51GvEDflzKzIhqsOTx9Cj+mzPPVmzyldcoy5SqP0IAP2VMpTqr7ip49f85msXfBv
dflBvvnHE7PZcAQ6ZZL0WQ9DchKrXXPx/DS9lMQrQWIXcxH8kkhgMX2eVH2OkGBHqW2jorZcZ08M
/Pv6Sq0VkgWFByeRhSGtQqTUGHvfA52PhxIAzGpxQPYsKXs/39dAg3cimc2ftYVI8QN+j2fx/9Fr
xXfH65MNOXBhgLPbvQasMYBoPiATCPigP96DaOdp6BEA0g8SsXNE89SHxT2BovHDnmjC4RpaOIs5
sarofyXR5MaUEmkSBEUj2YVIn05xhtE6Z9QYLndz8AAbIHEnPWAC/RfWLu5AAdyfGluEF6IneFkc
qLHB3P4cn2ztm5rwu+6mQ/vp830Im7WXQu0a3OiKNWmEj9txR3qdO8CeYmutX68lyVBcem5ylFCf
AaazpAcQjRzngnjNHWsXAbqdlrmmpf/GB1fcN/cpwWxbcrDA/KtYy4OYiDzAhVwq8Iv9jhsrstoK
U2yfiTjw8nz1Jh8QQPil2fVeZC4bQuAtoTeX2aDTMj1BmG2YUYOYWeq6FyX7T++iQmZp4fW7vVaO
z/I1Y4Nq4zvBC13578/QLTx71oe7h4i5BhUA+1dXKIZo53NyGEmdI7RnQAiRIyieWemdUV7qDs6D
mSfkR/7z0fqhqIAA/aiCg0f6hpYD7BHbWNn13UoKLir9Cbj1fN18bHrcw6RDDJLfLk3vdFk14Lkn
sTImiuvLBvKAiY1/L1SzKxY0sk2tEmGz5X86MfeAfNxXVsRSTCHt8EFMLp3Q2WNuqDmv2KrqlTZa
alKRuRUd2QZTCs1DSW35iUNeD/mEtBvkil1mBXSrqdxlsWZyZOdVrnqcOiPMh7FZC9iS/dbpR/4M
q5LD7/u6rdHyNs2eXmLAQG07uPwGyCmk3oR7A1dVydiI9FGqAeRlqA0eIdy3L8V1IJFKCDMwVZiN
wZVCj+zYfKD1rpMufLe0I09YOXtNVEkfAx7t3E3XmuG/I+pePAGPTDy54zFRPsDjYjOh0qAN0USn
Irc/CQyGhcY4h4FGgNjBOpqtfQHQMuhtpOPv+/3kvk5pGGteVJb4XaOFiibjbLHhJsku/NE/fkL1
4x60IJzpLJpny/XsOGKdcarJoTdUbxW3vI4Cswk3y1Qjo6a9aTfnAQs1U/Xy5tt6E28YduAnQmCB
uub5+OpJsedJyKdcfAdwMaTFwf9cRu6JMUdPYXzhxB6+jcg3Lfi1LDyeo1bLMVpJLf28O3Js17qv
v/0kCpzHre5nDWmUaKlzi6VGDQpENKGEysIxX6KzJhAbnGDatFFKXCsFZyJjibhjXyDj3tzyUxxQ
FqmSy6aSPw76DeK6F+mdwN7CCRJ0h3tOTPl0gwnjQ5t6d+l4Ve9LEjR9TJYcsUVse2pKWAWF0fTK
BsZfYW3rjYhaV0yif8Er5UUDe4rLsjsHGZRCPJMlhGisd5isBCyA128B9Ld1s0DA2Te/K+VwXaqM
IkYhu3X00EFr0uAKe+LWqiR5fPYD9JG/GE3yN9V26aSg+RVKnsW3xl/R8wRaoHDAYhZcDdimrLnx
U0EYLmUU2hr+RvKtj0QBYv6tSg9YtFcwx/gtfgjCmF02qzLPE1BTFPSBQzdj1io/NQtxqkeLlwAP
AGTzT5SgpBwl+BGgHmc0hwlw5Eg4KzPNnuM+wC7eooygbLQ3E4NKRI5R9+JsXmte7LQPiCyMK/07
BRTFNoQ9yekt1i8cHQoM/f2hQCzNlA8lpavi40RNlANmVrBHCaLSBfaQ/OkgPE8ZNkOQsAm1hdbl
qK1t03NlZFIlEHaYuZTYtGG/taju87sFZb/WsNPfBZ/oFsBdINpgsQ8gwvopM6/ybBptkforkVbF
hQ3ql0wE6PyHUfxbVebg+KehhFXjOf2AZVvBGRf83xjoghdMyQwMfjpTjwgHOjuPW213bkZwixbT
f11xpVbnAU7+EcnXx8a1pjUY671dcIOFExmZy7+pHacMjhXUpA2KusFy1xoigUQj1G8VY6ia6uBc
gVbKxQGKNWBNfKwdIo4/d0E/IVcXTFW5ZW6zUgqKpw2sNSPmmb6PWP782RWhIIWi2IuDMzYMCwZM
DjqPlebGxjzOXPq/Y7vGpK/E7Q8g1yIpYnKFCpa5J9YtAGS17E2ow6SzfaxpqQZV2cbI77hb+tQl
NUHj1ZZtpHnS+pd68uh+DWXnhkMzGky/huWfDuW8K5kLetidQzzrrExrhANg/aYihhR+/fZ7vN6f
Qbm1OUbkm4IWOyt/jziuYjM1/UTs7sPPIX1/Dwtf0X52Jt9M+/P2Fw4Dkdul3nyLfj5B/wieNqqN
yYobCD4L7q3hGM1/IuCxhSqO2V4u8eobYrgp+gzzCi3ji54M3GEV79PiHVFwftTt1DgL9fA4i/UB
PE9Wrn3ga+vk2N59uMT6r9oJKoKDB9N/sPYe23NBVZWrPgTJFsEsUMaGDFGI8N65XBkFSYd05Xjh
ceW9nD0q3+kWqkZKKNNq+PWryI1FoXDwsTjWbN8uZZKM3MkERglV1/EI2tMXdvHyOO+jUyZ9qfLU
PNv358gd7g7bNje9DXQ7pf8k8GP6EXnmE7o4MuokFXC9i3NszGQ4kVLrOWmpbTvpG72PiSP+z6a1
mo50cglde6HsCarbNPUNtuHUlu54tJocDY2u0n7XFiHyOieqfNcflDoE09RayNogyewVvDatIocC
rByFrNKbWLET9UfQtI31L1UIWb4W/66sCXaez6VtxV5EzMx9d2Yg2zVuDFTZFmmOjww/JWlfDB+a
fH/sC+w9jf16NmDzSiswyI9p5xfrdgSFomzt0Q8LuBk709q2i/st0gxb/WHrji/HRD7OJVw2QZ17
y+wkYDY9rZNEXGlp2bYC76SwZAlgMnkzgTAiP8jXZhlDsPPodaRiVT1A3bnmZe7Vzj8Efge4WF4I
90cT/gTPhB+X292Iw3eXGaQymc67ksbl6GiIP5Qz4FVH5ohsIVWb7WeyvMsZqPIbtLkeorR7bxxK
b4p2vTa+CJilwenkURGFPFLSuXaXvKG1+4ghzuU7q65SlqRHIiuqVzr4ZDOCo6N0qpe8R1hCeSXg
EcNQ23H/sYiB5EkqzpJXTCjwtaBA3W90MhYty9YHhFFNxM7JoOJuxVel0srtP4DKdWHgaua07Hln
4ZxRc6rL8NAM8eU6+DfqCil9ZkHvzKamVt+y03/hz1Id6GlZxDWdNvVjxeizpmfpgxKyLk+1Ctyb
twbdWe0VXJH3yVnOz+JGV8YFpujpBwgr6qxSjTQSFF2RNUhU+istz/SXaoVPl+GF2Kl3acMIJKD9
h8zqcR+Tm14HppJH8QcBC4JGdqHIUF3DjdBeA75ZI94LHhrLLL8taKNh+rowej9oivVCXZ+Y/l85
gS2xJz7hxxtWCg2B6PTYfyLo2uZOEOwkJyjbIIGbbw1H2gnKDIgWuCCyCgpOU0CiJg4eDQlIDYka
TGywhkBqPjbQxmjm1CEnESfBQAIl/qbWm4McR5Xq3U8WatL4d42oBdjYaUad4UOImva1KcY+uB1m
mMPXL3j2iIY9fD1NaSb5ULgShhC+J6GDrI78N+ttcPmjh8Fszrx6lcZn9EIlq8Mtzb3xb9fw4DLs
nIBv/7wxCNNaerS5fZBFfH2J0N6ODDIX9rFYfktAMTQnslT2OhRRLAWDLqbobrlr+TMneiK4FMjb
WywbRp0RIM9HUcJyFJytWEh+GiC4lWTByLLsRmuFro1GaRHkRS1sF+VK8Iu8V2N1eQLvJbFAHSSv
tgmANgAZ0MVuDfmO8ZNr3C9vI+NgaGexIxbMtbjkWTZ3wTrBjUzmjPqK/FQwdV/GEbRwuC72JX4g
d1vlnB38zE/OJgkoVmkhVGQIDn7kvNihvsgMmWygwmhyN14qQ09Rb4wA3iXSKnr0s6eiZfEYyPtA
JuT5frtyPUW0BdiIGjS++oVPPUAh+zdnl0DQ1wqKR62tjkIVlwcv/YN296AwXAQvDjvTzXAtvQd1
CihCBSMGCKbMsby6woEZfgubhKBAzwtx2FrsvSecZMq9/A7NnAIqPdW3qIfLP2ZwynjUG5VeKQ9g
CnDGEmXV73+MS4dRJNoOkMMxl3aOGZ4qmCoV9EE6Morhkanu+UTFNzOem0Jyp64BRrkk1P44O3oF
oKPBdyroP9M2qzG0pokpj0ONvqdSSkdfVv7gVk47L1vkr/RohG+aHCVlQP/4usDNtwXCKNYXFyvF
UbeHy0RgsHG+NcBkppeq9Wf8dXMg1kA46K0LGp1ijWxvGXlJBwvRGtrMH1+SOhfzU7XXIwHFLqid
fuAz2czCtk8GWFRG505j/Lkb//SNgG1+eNxQ6fPkqmpr+RiBtPgFDNSqwaIBRo8QY4E1l5dkf1NS
3BAUiaeTkKUGFnhjxhgleokIyneZxCiKjkH0XmXlsIxbQps+j41uBdhjLrNntdNdTbtaHoCScN0Y
Wq+f2ecwGzcfxNyp6rfmLQBmHL00+DEzf0VQeq1wJMsta5I9Rus6WlwuymUMRBYlzynfk/OGcFtc
nX8x+/E0jmF0xCVJ8GF+OVycFmi4QQjDzMFe1YGQlv5jeIkWj9kAPRyH3PRg85X8Tw/ImLoKi57r
8iQQ2ZJ8gISTZ5nhr10dXYO12fRjHGVxYG1Y00eC0YbqCOoLIYhJkQStMoeeXX7haSkuFnsKkNI2
tS2bHuhpWkPyrj9iv+2Vi1wTkwoXqQn5O3L5HikAuxavNylA7hvgxgJmlIT6mu73I4thpcsqxXnD
rYiV1EWjWFt25D0YycFB1836QphBzZd7ixwYcEFFEQJMMdZXWMMGigc5pF/0XPzT4KKAyfojY2Qm
rte2T+uUr3AFcgjDrX7OdTgmha9K0jRW9imBVP1/A1lQuyS+1227SB/xUJnEHt3t8trpVf2y2VKk
ejLtETXUehapbLKrEqYPx5Q8868Pj+EHARfWO+ZsKOsc+AQ2wUj2bz5n2tKXKfVWyEmZwtkUmgLC
vrvcpNWlhDI3AM3aFCEomOi+q54Ir1trCdTgRPaumRNXrKNti7sG4BQlAgW0G3CTgpny7vSm0Fnz
xo74eW1tgurGv6PAqa6Tl/OYOsCFLj6WRB66kVDXbMT/rEgEZOYQBeArpIHgqgW/SZCUJlkwEtdz
yaq5dIhTM8uW6r8QerH1Xxom2gKkJ3BF3vP+OxYVoC+pBC87VwyIbGuS09FVxs9I+0aKh6le4R53
Zey4UUvB3jibkhHOSb31Ymilcd0vtC5Cir71O0KJic4jMGy7b2/Rap6Th+VMiF2ChLHdcbGKskhC
K/2NyQNTDrnm0Ywygn7vgcT/S9EbkHXzmAbgtEHUZ7EeQwTypdph9gUO/759kADsowTVhmDXfQVl
hsckBhirwnqdJzUzIU+8wLLrVYHvPAQefbTzPlN0vJ8soNcxKTAThuC/VJnySHwExiO5zGmRznZl
aRT0kPdscj1/TosMC5hJA0TdfRF3KYaRYxJnypuiDFr/a8EwAYrvO6Ne21mkbh5uKLGByaFKzW8N
ro9EZTIF+sZTXoaFSX2450myLnioTvHfOV22K+imLPxRs+7WP6kezvZP00zZcTYxoCoy+FOAXR1J
lLPIMhBY6OxL7orSs+j5MfO5VmEhrCeNr6feXRodSjwNBzKl1o9kUL7/QbJk4rcotYl2p5gnpsdJ
Ua3siZeh/ShGxdY+Wte/kJEAdr29JfGEtj4RHKKyyzK9D3jDU+5yaqNsE/3LhXVtY1KN+T9ayMhI
CVR9BCZO6ey1VhF4bruQxf1Ye0jbyKTK1itVlBU2Q8q6zv1EdLeytZ7YhZel0fWgoRwFZyqyRRUp
//A5ADiMPSUtPBBtfLWw/DxNODBv62Rc3ya67PBH5Cm4SbwGbtp2ybfCI8ZZ9og/cTJMJ1C0N9eK
apM14SvrIC/2GOf9Chx39JJ3pxP3xqL8Z1mV2BDZC2kxBmNvIlrc5tsXXnu9gCihftOO2xvD3NF3
skqU1Nf2n7SH1pXHuyjioxp/v7g+X22FW2s4lY1uCO9SDXUA8uB2d5HJRhdnncc7MnDm0ybZqLU+
lW2472GqjSG3X8aFGfQpTQhaSrTCR0IKM75lGSLU6C0dpjmP0X9wn/bCngCirASX2WY2BWURN8FY
UR3RRaRW2lnwCzoMOS13YtaKm1VysMtoOlk/YmzcW6MjHroKMYlRNETBE0XhVeJVp90CvH6O9g4a
2BXqd8M+upvixeyGbqOaTm69SWFucEcgE+pUhRPipqLWruGwF8eK8y+Yhry4MWKZ0E3f5RZmB2Dk
lRH8P3ImfbXL8dWiM90+0W3adWxCGjS5l1FuM88DXL+t22exbCp/k318uF1U9FbsNBAFxdIMVVIa
mgLOkjQMv1x5gOsgbT53AqXhbWG9l33QaTzUnAJzrZOXnzhxQJDb+HoBodYzNBGFMooriWou/gB+
OS2UvqYFFw9/B4d7RIyssNUkOxHkE+YRNekudIj0yu/lCqqG2atMaSvfQLicN0gKuVyywgdqSTAr
P6TzgqxLpBEzezUFhY8GSfu1t2UqMNoKhn65jDmly55429TCqs+L6EVIk9HAuY0PNmMWPjIU5+vn
wpULgbdl9lhYvPAm4IdcqJnchMDHTjbCjkA4DxRowZWliUK5W9ajjv8dtQhoL59GdqYkwGT9xnks
HEcC/RxO+hUZg1IryH+noD9+QPUumZTZ97QxKsM39qVwEoaZZQd87pdI/pZP+ftSkvFOWy3EHpRf
H0ro2iUe7AWD7ZSUrAIF5YN280/fEEHylhebGb32iRDdr/0ivhzy8Vhkrvl4CI+GxSF7jV4ct9eE
80LWb7QbSDttYfONnlUORyBmfyi7NfMN+k7mXP+oVmQnI0yVqqoK71kEgZMpoz/5HiEnN5ac7Z2E
njzv8vIGo0DOnGk32rX9u1R1nbjGpUhlEOKyY2taAuj0mXD9FPkhWo0akjlLY2OO6IoSuIypNGcm
uYLDEfgsgQ2udPwO70/V5S3VBxaUXtrMShA1c5SCgiPLblcHWTC8Mq3LtOfJkxSB0MNRHmPauvez
RXLq+mJNlqEXhLi7QIDSq7nMXb0T2ARH0FwGax0TNEO7t5k4P9HsFA7niDGegQ+5oVd2uU6dJH4U
x3EyNE+3m/XZ68IeN58kJLNuELm3t0k3NTtfWaD1lfl/SmzwaWcpuMFTrCz18LNAXIpPRWmHgsAu
X5dvE5B8y8TPdv7QN9ViVF+5ymcgxtbCWV0MyJgz19YU6VcX+cxoBh28L5cIHf/lVn/IumQw9BSo
oGtiJHElNqEfgyitcqqX4jiUttM8o+ZvmzN9D4KgmqLM4QPj0MrVze1ab4+EULFpuPhq76psDRIt
tdShok8nakFL2HtMSuHYY3oQ9ZZ55gwaBK+QG6imhUSJXmy3swkvM6Muqbcios6nOZezfe6pnvYA
oCaWlC5a2OBRCLMC+N/tX2MmyFPYwQn3HEF3TS3rW+XaHWEdElGSooTOJcA2wUOigu5S0Pi8EDXS
KGxiBvvDT3XvMiNoCyYDSddLRiqhAGQ77akbqwFCsZG1KM4iSxxB/nYeQbLWoBem3nZ9+s0Cy/8N
XPwyxqM/r1y3y6IYLWHOCAJmP+L8um1Q/u7fM/WWCL3Q3LbzkLfW+JBTf/CoZyfjvIBFdMyvLEA1
6WudRIaXNby7VWvGGPPKTbtpDuFaq0kZZGxutDoBf8IlkflqyZ6D5bOYm/Qng7p8sRQQkbr0Jy+K
ZcNgtJpz5VJ1JmpZcVgqouFFS2FfKU41T5xau3u0wevAS60bnzrgM/NO1MBXPRUP7RKWKf+V8PMw
NG3/yk4dDWn0+57f9lIaDLN+Vgi4zohWSDuun9D+BMd3NqmUMIr3l+aECAB8QyiweMPfJsUuJgv+
tl8d7uqYjQPisG79ccBX1VDRbohnVhTfBFm5Mkq0VuZ70y6mQhtsEnBROP++E9m8qdNglo00tj8W
32uI10noLsFxR90J6KSGFkYagY4+9Dn13VMuKEbi/g2iDEgZhxWvsF5CwLSbMLLCPf7TTD1CRHcR
WgUl/MAJCV1QjinO2tGxfaMOf4zr5IJShc2/qG0gAVSMqaAEgnKOyP0l2FE4d3yW0bZ1ciLzmx/D
y2ZkmAmRQKcmUS2y2SnDdzkMFngpjZpEHsTGjExAczl0yPv8+CI7buGu+wYXGg4cHbXhsYQW5k3a
gebgFJuetHC848vaL7mdu2T2Il+ur+z16wQpjkRa21jrMSP94BfE7NfNrwmn2NAe9O6yKTxDXNDE
soWx+QUrM0KeWVOvNdS/ppFFdN9PRgIz6iC97fXYxcKqUOvYY2JFc4w4DeYVWYRHlfpYdRZ2rpUz
lBQ3sLEB/QeujPyZwWqSdRZK0QuYnKY14GvnnXUU37rWYzuxnz9Obwn/zDRcGGaFTbegJ1cfJTCI
yAESNAO9kRDXVZiPpNvcLIaT0i1U1BePEzT7fqwBhhhwe2EVeOy+fBYtF4cG4Pd8hu90QjRojpPw
r5jir277wWtk5tE4vmk6oineXcfSWh/H/1cpGzLfgHuvbEd3O19WVC1qBHPIKPJRMBPfoxIndBZQ
VWh4k8/NW+zFYxxHKsfOLKvz23/TCiUEcN2cbcUuYMtHhQChNKbUcLUQQi/LauDCxd2kBKxlr87z
FM4HXsc371N8ejwnw+YSTNbKOMqUGaHZIqBvAa2yVnCzJxwiORqoVCizoJjGjjvmUT817Sx77kSQ
HIUmmEXpoqMp2PI5HMeOqlHwK8YkQ6+sSz0C0U9avSRFPBvtH7+GhPxr0XB9FhkPbOAnbSLkfUdO
ApEWWIft7TNfIpxP7PZ7r4xOtqEo/R5FtySC1ZTJdR4GQJJ+yO2+3vJ/9CZAhU1H/IvTasuGigaA
fd44BKVp5FjWSzoex7rzDI4npOzElgJ2biKAEb3gR19+MHTrtD2NxhmEKY9F0G9JLY1dEKZ4+TNA
3635HaAFodg56bjH6RRC3aYO4TPk20ZlTsMAqY2Yq/HaTJDPowxD3rjkhTxlffMbqKXHcoCx1nmE
kVbHk18t+SSGmyg/pXpGlJvbtnnn2h6Y9VI9czYEUVUfTP6WJByn0RjS0f4hMZcVybMlGV8IIEgz
8YMB5EvAUB4/Zktq32Q0Yet7vTQ5EaR+yPktC/hkpb4p4txJbFjfQhsAq9kcbpwaZWWSKGCE1eiY
DCm4H0CBv/ruYnTEapYqMlFnLj81qKnlx+J5ZB0VNjynJl+jQAf/vJT57xNTmtfd0ok+KseHiVps
0mEup7jOeLqOIjko9IMWsUmTxO0ie9OU4aiun106p6dVSQcO4XW2MjSESluGQAWP+kR60WqE1BAE
h8kjvs0hXPfnBeespPpW5yOGzD9PzIJwghnmw3fzgOj1g7gHlD6L+Uzx2b1ggtmtCsbZ5cmh/btR
NvqvcvDTkvSgE8zYgvsUnq1SGwlO3wozdbQMNWgzBaeqHaoZ58r8juhBD+bZ52Gp2f7QdF94zFMP
AWHSvBsWZmfK4BI+MwMpYGZwt2AvoZugdjTvnz7sJ+Rr6CB3H8LRTfVvjzruCBBXHtSBWCSOawnR
D2BqKiMVUa2eJe5BXU/zru8nAJtVopMMI2EYMGvW7aqZR3hGwbG/C3OIRSBQFt+3s5P0q/9vZ3NT
6Bp/2qGWdGwzXw3BtSnqlp/WdwEiZNr0FbXTUZ4xIjb5J02bJHTpKZeDoP1kWVsLvrdGwSTxgqZg
duM15V79EpSucx/yBQQcfxpfIqzhe1ikblKHBeWvBjt1J7k7iAEHPb1Vs80YPUsa/c7a6cT2VM5c
kXKSGqbAIpb9hxtHX0mUGUsCAgtQ8+7pxgxPpHJIvywFBW2PMSZvzxdw2UH+SF1HxwmejcfOQiwU
t4J1fjwWZ7jm2isP4uNxNn8GJUhIZzuDJapRVdgeYyaBScaabVyXgmi4/Q92n9SArNzbPdEcpLiq
xN3yhci+VWP+wNf+UO+xiCzP6QexhsRbsjce7ugNezchb62EHEMT/O5/bn3TW2EAkCEcZNg6rGjr
35cqPJHcS59RpBScpSM1PCmOX/9vvmN22t4ck9s8OhMHnfv/ohCwB/BTkH0wuMNkVXasx10/Ecr/
x9RkahfxjFbboCE69xFCi2r1FElyJkPoBTSVaeZkEVJ63wlFfgADUzEhFUwBFA+BFWCDb9ITtVDR
IJYbrcMn9GoH54U++zo3uB8D+estOtGSWSf82HE2yL1uOTegZy23wEYQ95DcAxtf/meg4n776GQ3
6faZrT65lgJCSKdOCsxq8BYwx2DtHxJesVPNofSOCoyx9SUntvUcIfx0kiyio62xyiqWd1EMzkin
VjD7jK9n6NREiqA6/xRX6xsRYAj3NCK1uFDwFYC8nV8t95rA6CQOFybRR30uqzxOkVIEfu3PUhhh
Os5WfceSQzSW0wWNpMsgohtsm43ZTcOxrw8YWg7tkayOiMpCbyLajT8U9+CT/p3Td7NyQSyW+s2S
BRstUA5IGaDDx1haiDxelht56LmI/KtI7g/EwGPr4xGQBr+Sf4ZdNHa5Ol9G8til4+bjhW5vLk0y
5ovrCvv9AkJpSdPD04DrBQx525qCk0t2Wcx166XFuyY5sep750fTxK+dv8GFagkgdSIsIKeaEgCG
AHuRVcfrc7o/CvuOXMG6rznjq231940UK3FxvLOyzZ6O1Zgav5dF5GQkfeZy1NGw1AjL2ocRz+PO
uko9cpwKfy79hCy6IF+8sAeV1ADeRwdyF8c+LwJb9JoBEpfQ6MWP/xZQciiUjIrxP7eBMJ6F9uEW
uJis0FMGjojeccsMd9rgg1ukNc1Xo/lebuOAOI3DE0ycDTeUmzUcpfyuxylhHjgUo0ofH1KWoiTR
VZGXBMwhfRY6Th7P3OY06q7udist3J1O9BsikRug0treiUl8S8hL4lC4Dnp26Q+otqMpXLvijpk6
fsEv+tpH8yJ3OahMXM9OTfIrTxurfXrPcltkQBHCPP9FxQP2Of/p+C8jkD0YI2nfOUFpBL7XpgxL
mzUShjaqmc31KkI39j3yScC5sZgp90BdPxRYExlQitpRJvM0d+bFeZTYVIH/w5m0emeWOTdbSdok
gZdRTXVsD2HaIZ8xVKhNXejkui6bEDWUM2krbcnXzixWTfCCRDjv/sXX3+elxJmvIub2ut5beOqF
hhOG44bqedCzsoL4hjSkqt3/mkv1ogu3/okVGZcVpVcbL0m2+/3SQ1cdWGMCDlKXm7/+2dc48Vg1
A9QTDFpg9MpIh7I81QLibELF5yyVfLbejOIWCfo8wWHLv9XH5WsfNBD6+jVW5G6eVRpCXRHra300
5ayGB76CWOUosXm8XYuMCpFEHhN7z6cYZfsMInqgMzpowMT1y/4q5WBaKctpsYkgSXWjyRNZDfPI
Z7rK6yENb5PlmF+OAN5d56iOGWx0qE8kSBj8RRxYPl0/KT5/OXHszsjTjJxBA+XeGldyW7tx/lsW
vyCDihQ7Z/Zq9OlfuR9ez4lw6Tgh3Qv1pIuVhfdNVgZkuwwYQ9YCUUntnGJxS46KywhLzCdCf9IC
Hs86B+ri2+r+Ous4dZrmfp4LbisueSm33dmwxmLBQRfBp6SYWmMqQWn2K7A4unWhEl7wkejMOCTW
Bb1HkslrJXvfmL31i8Me2an7yWHtxsWNXdidtE1bE0QF3ia7JX8VvwTuQieztv6970D3rgHGhqAA
0E9GumuyEVIrp1cSBgekNVrx/C0TMY+p99TO28qKFPlPHpSaumggJeZCv8BaWwxDCrU6KfWmMUtP
C4WpjY6DqOZ5Tx2tvGarf1Q0B4t4bf5tyb3S1d7aUsk1tlolRzaa+Om8VSvn7uMCTlTJmzPlvXcy
JlhIk5TYNOl6CnhkgW6cTL00720w1EKxrn7iF84Zm8/QJxPxnvIrBjf4o7QlZuGd/fPphWh9vCPe
mscpsuaDTokMia7OAGOSKfonhVtYbH9qdftxdogaO0KgnF6/T0BVhBkhokcGTBCDTD6SWm3A9xiI
Sd6NDtYdeR3rTzY8mNdE6HSnnt9s/xDqhuocE4yya9bymGA1ERIu3f3zOhhqeOleuT33SD1X5Mm0
0LyRPOae16pZ51zncnIfT8LE3azZhVtwn6mZLviIsOFve8N7rjscN/r6EpudxZ+jf3UctvIpaNEh
S9bMMUOXxjtJFvFqoOZYwsLVXOYnrpZ+aozcLo+xTJJUH0MG7q43gwg3cqsBkbEd+2KXruP/uzRS
mFB7CQGpxyp6mv9U/l+Nh91LtpDhz8YGzDkcgrFVt2+J594ujZAwDoGfgBlyC4ijJHcQi0ZUWV2K
NL2nrgNe2yoikPpl+PBtHqDXNH9a1OAZ4YifF+aVtCrVRXiR1MvAWNhHSaSUtx41yN+xuwZkJqrg
6VSDj9f4x9jhVssrIb59yJBg3cUBBmoQWCwlvczWa8Ocy2I7ZL3ijhWpLAj4d8sIEc150pRU81bn
W5nyhH9e3yehOVZO84uxThPkZNM81Z+Bg1sX8fXtizIResatQjRzRMqjaVMdwTok20UmmKanr+CM
rJCTyUfuVBfQayQ87+uBlazjFS4MG0wQaq64bnOj0HjzvtoZcqGtDkja8DIizxwlGQHtQw4Gsd6f
0KjeH3QJmyvP/iMAMPtZMSQ5rzdkaBkL1MZ7uqkYnEuHIpjvCCvloceLblkbomtsP8zdjgnv/VVc
K4ellYxBuUckhPb3WyKGXAJ67NEq+ejmlHsW6HQvwJbRhYXz1h7LRqszYmVU7O0o0Lb0ObcBSLDR
tzM7XcLr2WWgnskZMZnU/+j/Wi3b5f5of+F/2xkRPewoxxCosjizlLJQzsQo9gdDDuJ8Vc7WqT5u
HrHB3G6i+S9AgtMw2/QDBPSQF87XExzuaZe9ThYGNM+UtWVDE1/my7M9qOwZYkBNzgb8GGOwjRu5
3bK1j29tnaikU4pwBdRFUeRuGpuuVoCa8WW6mJ26VQxMjdoGmDEddAemRvDHZf8EuCBc2GvHgtNz
ljLW2Trmv0yryAhO152od/iVA6vYlbBPVTttTaMEXPtRYraiP7z0qZaEDVj/gSsEOzHPpufSbTka
GcYNY4FDN0GTz/TwaQ97jtiUUaBeAZndLePH8QstcNV7MZ1bjjO83rPjY1UcfsIsrw8Z2l/S34U8
ti0GtBWqu9O707rB7oOiL9rMOQ2p/r0t4lcHWrfmRG5GX79qP8tS51R9zEQSMMP1BGvmfVL8sud0
+uiME1lYGtcfXIk/MFTxk3ZNMXfiiaJS1/mpcCZjuRDjBK1Cc+osC732KCyjq9SW7xG6CDESqKo4
sDJbA4LW+UaUrWkdaS28blIWd687JSmRsXo0a33aHT/gWMrdnJ3jrJ7EmWjSMVj8fFosu6xY1D+E
zBueFTijhAYivHKI0+uw2Wwl1VHmEgXtcfS1MSf69C1qagJArnd65IAmRvRFsVu7Am/Wz244mkox
JiUn0AUVyUtPFEM0l31jlZZ33bWoPgbwgxFOZiVJVU3s2z10EhymlMO48pGJKsL8W7jDyPjfFxRw
n2wGnVfLlqtmc7bfrp3ttTpzl/QPpQN/6/8SxPNgG9J2xPjeXf297mTVZMzvc+nsVhRKZL6GYdih
1vNAJxyr44HdILiAwFuisMKyz3iHLYriTfSxUGXxr31dZrIVoIITIEkZD+IX5kJxWq6PQF8R55UD
UeXzPbHPKLRV7mibY19hPChEjA6mP0SGWgRbczRNOrUldP18JogQ+5TaOj+kgC45c1YQNbzidSiK
dbG7jXKclLHAGDMKikNNPcItgR6MXYL8MyohNQwtbTDiPYwOi23fLR242a5SRJ841Biprm2L4V5y
+W/f/5cPbpJjB+zeT/VL1BOX7+vmeITzhK6zYRWk64Mp53hPkI1hNn8XRJof9+wTVXvtEUBsOphe
UFQ0pA3TiocnWhy+b5hx2VqRn6k0Xrax6P7wT1NLFrSePIX00HMTGTuk5LU44ocYPnF9De6vXfv5
O7we1582kE5V5WvznvqY2aq1Pf1/W9O+o9zvUtwfvo9AxYZ3aNbJrMpSLQKDc/s/Nl1DaTL+ozft
SyM3NraBlVaTRDO1NnAD96ZDMkr9736RkFzk11JU+vH/yUtC2ekycgEfO3Q0etXS4CFW1ZgxajFJ
VY9Osnm1tTh0MJwZmdZ1Q6gjBbMFFY0JkGmBiCkpOXxHOoOuillaM78mSa8X8XKxSjME1SaeOX3l
/SMyogPWSR9+p1SA35Wq6+1EwceL30Se39woWSpq+pYmQSmY7AEXcJcvswo4g8pZtoysyPYMxvzK
/qmi/p7bFpk2mLGlOcW3SZOprqY8xE+259SJ4kDyVlusURRp7qpFjJF3LStBKqtFsWM9f6WhdS6y
MjI9hX/nZzRIOWOzFXWHnBP0UHtiN+gKb278JP8uu7XBmXxoa8wxco1upCXwTkrcOt8qJKFjBDEm
VB/pNdGg2H5To9L7oOVzh3WOk571Y5wMJLmEKmVaX9X9mxkVB+bSFLWSSs3S3jS8Bkrzh++hCWqW
NFKlmOm2VumH62xgmp+EEDtZJdTDuOddfTamiu6JUEggN3jQ4OGcb7DRPfis7BAbTmasJKNE2N+0
ni004U2uWxEMKIW91NochBGO2YTiPm7QFT2Oo2jgdOE4O4t2hHdU1nrBAabUhmVQzsHHPAH1W2cq
tC2w5G6X99wlfs5aejPhW0xMBuEurcJFgcfOQX5cW28xb2ytRKt8m1Be2dP7iQfFi+KpLMi5GcdU
aKAQXhNDrqWyXzqg/uPx9Sc+zavvSI/D1kWxWPvVcTMcJssg2HxrYHT+0ycUuuIA/GeqmC0IkfNM
fl8jsTvTkgLndxE0s1loRlBy1iLTi8dq6SycQItvkLxI31PmP6oSQreL8ARAM3dLzWoCAGnZ5Quk
oZXkD17uWV5M/aWGiMl8Jq63zkJgmiVt9V7K8esUei20lH+0v3CRe2yTFSION8mberAt5AQ157dq
UgTvJtr5aF2RDASrHicwFuJgIaibCml2C2bA7058H7r6nP3YgqAqCNAT2SujCkV7y6rn3U7RmBDy
K6DE9O8/lVdPE0z2SUtz9HdCRRNRtFcDHdV0Qux6dDivbQp9n4S/3JRbjZAHSoKSur03u3mZalNv
hL0Ax+VGzelXSud/lX90oZqO5qpJDrBkB3SK+gc+4nUHHXFAG/7qamBHnySBRgQluNJnQX/WrXzW
6fcyRa6g7xm6kc7BxJEV7f/1d744h17JjEWqBykH97ziqDCY6X/05oug2Byzu2sRlcp2YGC/l+Do
COzF8Y7ujkoqUrAhUsMElX+xRhlsZg17rEeo8eB/hl0QUAIUCvIB0bF91jPHelK6AQKFUK7fXtPJ
CQ/G+5mdo/3YvosTRxICiTHVX7++SfFzVLno0sLvSasumySStXNMHUTh3ECe7ZBpeso6KpFt8+g2
lFny2g//d75N8+1aWw/w7eUUH/j34HdcbmlVM1VjsyprcVMrXqMTRx2qdmsln83JlwS1WYC9pQKA
AlpMnm0eqQwBjNjwyKJBpUyVml9jltQ/P3c1T2RlQlADGINOlmoNhJvH9bm6isM6syvVe7+m+XZ+
x+YxtzCx95Y/NN2JZTQg/tN1dqaSXaYoQW58VFOMCaAecNfNhRjDSY4AtiDMjuPyyqxSWLETsusl
XehVaBx4NqmSbVpYE7sWCNi6ljLmPnA3I+jkfnSDg9doPWqppmW3YF4J5fC0DrxG9kw4G57xRxeC
/h070gYWM/E6BLDypuf29IQyFh9/kMqSIF/EozsHJHgwy9Vf/3OZ2L6HboTNcURAmzwqUau68+vM
zZ39jdS4efpZOhlAGitdeMDdeBk6JRhI/NrAtHK9TL8WiAtNve/5H1qUmQGhm1Ek5FhkI8ghIA0e
PJmV9yvpYalTIKTmNwlkDrQNfMTXZEsbtaUyJWpNYGs/Op4m7DC73jYImQnNi/2xF82VxsxN6dyx
zZpbsoLeaQonSr5xRn7eaWHjru/TXmiYgQU4j48kWL2L+BWOQK4ccg4MgA5eXwdQ/Z3UCSP/DncG
WO5nbP1L7g9dlO6HV/nIy3scFajBJN7Ix3rBHm8mf/b30SK4kI/33c6hZZ9utQ/srNZmdB9VkNU2
Wzhl2KmuQQ1WS1hP0hGy1BmjAJRIHhwPIVuwDl5RsHWQBgMx49+MjKk2H6q8JBBbTYEqugeGDIiX
hwJ6RptVZPvOPX2s8yFQ5n3KjxtFZpYNdnbZA4u7KYuh25opBrkgaJM/PapHQcDi/G4738mQJT8j
6wsVlujcMQwjugy73G4gf6ANaVRI/Jlp1a1nE6rR7KUENwi3TipOBkaq4p3uplyhf1poMpoG16ZR
FOEBRV7zQtSLsW0pxs5ECAHZIGP5M0QcdkE7GmPUc6nKopnD1HXPoVL/WVQn7Xx35uruOt23Ba+v
YMJ2MBnkiVuh4Jw3/G6H5M4xAj3Wn4kj041gUMgUh1urQgm4eLijKulpHTow/24Vt61hQvIyTTNm
DfZMAB8rWAi3fPS9zce6BysbcVOY1kmnZIl5wzajDqFsrG5rR56BtP5ACnlac1ovz+UWaU8xUGLV
Hha/N3cDN2iLjzVmxtYDBVM1VhsmXj/LkTLnttbra0EfZmLQQi2HFXhtKKlabsVWUY2DPvru9VC/
sWI3vAnlytTxMuWoCerLawkUXuyPGSd06KrjogBG0FSoTsO72CVQgGqzUazFBAL9HXundAXCoUl0
9JkAxPvJq1jzbmdhvCQEwN8SP7d6Ah52ijn3NvKKlUS3JV2XGhevS6w/6C+PP7+eZfZSkZbn7elE
UxjC2LM65epJHSWIfna/GQTxpw4AVCXiXhJ6Q9PT3WXh0B8v7otad83OXGegontD92vppN0B/qYM
C2BGHkq+Kz1F5HH7EzVOqYK8659Ej9O6iVmk2uHXrZ1puU7SAXX0JH3bVYWiqSlej+vXtkfSL3OF
RqdCy7ZyfqUnOKPjti3O8//Ecnaf2HO6/emd9O8kTNkNSS12YpI3Ew/rzBgfIfPPXDpWlpGmj0B9
7yExan7HVgj57BTd8ABv7gPPFMwl1qxxBXE0bmryXFZhDik2DcNFXmAo7mOWvI23Mbxy0muHCiYX
mPPVmPtx0i2I44ajJFnAQBwalQKKJIs0b6LBVWSgL+ZbHVeZeJpiGB/vdF9D4X1nq1GJAc9f0hpK
8RZBRj8Gtf+3vT2LV9plJLff9JAjqQycEiMrZM4a+ZxNu44sHp1dVGT4wARMmMyShuHjKP4B77wB
zCK9NfR0Jx1+B6kPIzVjEQcap5V6k/10IKh5kwL6unxmbl/93NoPJxa+JwNnDesEL0cN0fhrSxg+
ia544XnGWxtGVQu/LO96ReThNrU/6ALsC7wcXth/vZd1klbXEswxLUhG5yqcv40/jy/MB3J6SJev
0IK3y9GXTcMiMM7EN78TTdlqMXrbixAjJwzh6yASgT6CZANRWDrYoE4gVBhrHmHNLoLTiggIbf2E
e0ZC/9aEQX31hhNNobHvfJr9/Uyt+sR66XyqcXKNUz1yce0l3cDk6G4mEow52AaBCKKZOzIdOvvM
1mGfKedz1B1z/9FN/fvcif6poMRDjv4lkyMwlapzJ6fmzWGyAfvfv7UvFo1ts6zUMSIVsscE753u
WESHfdfXa1eKyrUJ1BJ/CsIu0PavIXcaRaLsRGDpwiN9kcFd9LYXrJI24fsPYeAx3sZ9VxjCzd4a
OV+eKTjTfXVqN4NsgVCkKWnfJLHkSuX3YspI3/WDgNhQ/mIB1xEOPB8cIhzShtRp4HpkoJHlku0E
tTvbbh750/QqMD62U/BDpkYZt3yNVBzRVNEAzDtzy9flfcoMvRGpX3Tz/8bc6vNVrJIb8ZtMZVKx
COkghqvLqTPA0QnZWLr55anSXE2O5cSQi6z4VIroVaXo/p1jovtiG6rUPmAWqW7L0Fjcsi6VPMNs
/V0rgdIuLrktaFPmLKOusgssUP5BNzL/+hC15rDpiQA72Ae/Dyovc8xLEVjkwwvKTJgUzyXqlj8q
wqu+k8xfb4IZ2oJPl2qlZEvaiCm7WqTJj/ykw81NG/FmN6Zox9lalOUK2SbuTrtlzX9gXUHbFQBI
0pTMAtgOoyMAEstAjwG0AfEoE071kFQGYYXhm02lIU1xhKAX2xmGU4zOBd0+agN506eq4iih/bgS
OHfpxld85Rh505VcAdtQwy/wIS6s5UQCUYiH5dza1NJ3LNQXjqi2SVd0f7bKJexaw+OpUMX9uAvL
YPKDXI2hLD63jUxKElDe9LJtlkTINMQ/0Rbh0UFpdftnAFuqBAoeqEiG/QtoXEdyEd0uAcoOW9og
AOrn8lPxWreSe75qLy+EsILQtYQ0j4MTGi7PkAhtpfOe9o6m+jIDQkSHXmePlvYutJMskKYjfnxI
BS9DIhfHj1SU7BYTS1sbjcV9toM91hMuaVRaYtO4EN8lnChMKa7/2da0iDcI9TxosSb0rqkomp0I
GIQVRoT/xybpPDi3K0vVPr2g43q2EO2lxgLK955yR6XPVunwR8KLH8kHrR3RToEbD7Qh+6sMnhqx
2Lc4MlRINu/hzh9B6cjgfbz+QPrwXC0dnARIQP1t64kZizpU1xKJG9X3b/unYIGe4xfmZWtj6Ohm
8LbEesRMzQClIYcdxyNT5+sObP3zE2S6UB1/yYCrkiywEB1grQGjowHVi8A7N0qTl28PFuNxVXpv
szEfCjfnLW8p26XfPO9L/BNv9+KfuHEdf34PkMDEFZcsaDqgw9VN6LvDSUzhaygVG/rpoPcfyI73
hEsRoc6WudphW4upY/goJ7pvSec887fKz5ljS6mH5z59HeA7KK8o1esYrMlUHXs1JBlbxQ1S6Eeg
YkyL9BIgS469KBcM1QVJuNvMZ4EAL0X32NMkesHa0f7skWH56iD7nEsSVEML8yiU2Prm4zV1VT+6
qHAQjkmkTSFr5JGgMmkZ7LxvugIXp7zAiR3goEi/M97QnmTmJ+rShduFGzxhS3oEEEtG0yLLilNm
iO7mVG2HyYH1bOfxLSwr/ZqmoxAgzk2HbsA+hc+sES3R0jEM1c5g8qBz5xdf+ndnO0OZkGhd8Zeg
SDFyFwjzEMm2LYzNxodGgfiGuoT5s6HKIzbitQ5Bp3rkWbtG7iYTC15F2VnpzNRTxJ2po27kXEI3
v+PWPBBl2GotHESK8xgW8NsRUZrE3sCTItqiztIqraUvOI7afStmEkjLJG4MqFdK922QbnY3g6/I
gAUz11eLNL244Jlxx3tmheFejjYCXiB70jgHBUhrVwH4Da3QaSlWc2IyV57o6RtaiTSpoXwlCmlX
sXed202smBKgVJSjVrCCGYMuurkFnbAx/lvXjU9MsnQmcwLNFUP8Sia2jre5SU+zk/d4oF2qXcl5
q2cHMOalmYAoIBpMs5a9LeZjVObMdpjJgpak5sdfp5GsYSzs9nDcRhSd0e6yrFQeWJ4eZQEdb6Sa
UwFzT+ntEmCYgg+la56zlcX0mDHsKpmR59j7MvHU/Wk/rMVc1OhtXA5nElBU/LXtRa4n2NLZZx++
PeuGMNMisfdXwEy9OlR6h301qTy0UBgwD1q8JVtozpEvNua/8x9ohNqsk+202QorKc/U91A1pUaD
pLScmsxSlBc9CxvVNoi+NBuSsfI+Wksc7P9Bisd6jevxs1ghk0Wftfr1XX9Y7HA8yecinSdMq7rv
XoCxkedXd05BT382T2ZgbpIjwt1787/BD0H0MDUK8VZu8ZnvQpaFbKEAAJzzM5+nLaYXrxmbefax
78Kjyl0p7M9mc2z9XJYdg5r8TEwnV54a/9Tmd76LYEeWLb0TVGjvfoJ98pmPaOBVnS0v7ZxwOuqv
gY7NikDu0sWRoCqUtHg9y14+NQ2neuFFk54WkU9W4imNcnUW3AFj1TGk2V7jEyjgXM7mQ52h4mem
CYPup7PsMiW4/IoK3btfkUBZXADnvmA3+IhzSoOGFw9vx3KpnITuE5RShFvBsmbdVETrmGy9SrNf
8YAl0nTFloNDJGYfDn7qUcannU8y5oYWJSI2wbI6Y8m4/Vkxs3MA4rbDYoQ29pmAiC/5ZcM/fhVy
62RTTp+IVhud5rk4OqKNrOezm23wMmfP2kb10i5re1Er9DmKag9BD2T3NKFfF6jyBuV9KZg0ngNk
201aBQwD8fWneJ93Gf1Ladk/reDo+ib0sBQhetaCCS95g871DmfKJYplLoD/4Bb5tFK8Wxo31gSa
DDKq84ZY2dI7dtklsLVFt/SwsvUUOAlLodNbQoAXYqcASfYEnUftkGXSkGPPJUaY3kjQhVl5tnyQ
wC8HQwQEPEOSIE2lsr8nh/uVvpoRwxcQWD/xWGue21R/WtTYVwxQnfptdeH8puDs2CjGSY4hyYxU
GyYgeDSvaZkd/ixYXhN+qPKNCggx8Uv2nIXyI1omrfubnBkmcN4qRK+OU8PrKdA9fahDzxU/olmc
a1BakAZEKe55+ODf9MqE42xE/051buSo2qt8AUUAtGN9TGiFYM7gvcM/wWlZrpwZPZfEvjEj111W
Vj6m+7F4po7kg8n3DCUOlQR7rSBKmgM7X+mMDtYeiywg50iyfc1b0gBg01v1lr2QMNcwT9apMd4I
0//M4Wrl0sZjF00a4z97peR0I7qyHISe/Iz7Nc//jNsMeRkOSaT7HvkGGeTyWRShIASPYK3ZAg/c
pg49uQdrH9fMtyJsrueSRSf8SdWCJOBhyNuPeDb3gFhyhvfhy+e/qbSafZPm6r3dtpYN2XlVuQy2
2JT2mB4fogHDztnjmVoHZd7uJMX+mY4roEwWzMbVNmzkMXz12q1LmD+HdxApI0LQH12Dzc+uyN6c
VrH6lZiCZCzJ4ZeGwYgUq7JQiob6j9gdkBS9ibQJejDDbpD7ybXU3LR/uOEmpTRtIH3CTBuCX7Gh
mg8VXrkxS+yuEfrO+EyW4XSSqzzSZ84hD0OV5lPJmTq9JEGD45V40eEwY1kOZ+XHtukrLefd7frU
Lnf//VTWB3o2KjizYbEU6h+mHNluYX/4p9CAkjDkYYZZZK2zLwxTiIvG2hkSbCfKnBVk5kZ6ieRz
2x1jPbGJ3jTkwQ/gyxVHFEflVs6bnWL2Z38NQIcBr7Qxqhm4ZgUe7Kg19hLQTWXv4Nop5h0YY8s1
+auG2LUNk9CXnNPgeQFRswuKCCHBdt1so9PY7JEt2UVK4BBB8sD84TLkIsQFJKDhSBqLWtJFUcFY
rQ2Ax75Ud+Hc7jG3GQSG93qdr2WGEEeRZWMKGX9J/oVFJOjmH2nOj5fpGKhSPg2Tbp9SxHiPT4QZ
p2i+HoONn017r5PIZufpRgqijoTXhhB5LgNBYlMaKDrKDNkK5VwUaw9ozQPqvTvzHYA+pRl42CsL
FWLH6wuYAEw0AsbcbgpAd4SttvGGijZquCq2/sAE7oVrw6b8J7DHyQzmrKfmHCkJmSENPrqDV3wE
TgblRb1pP7RTfQSJt3OKkvE8JV4CTStQGC+0dEhXZDfgc8wSWl+5mP5Mt/FTurOgSsNqpgJmdOs4
JyQ/hnFxmbAcyht/cz9lVl8w5IHsTjmdIWxLQmmV7n+Ol3rPzSUv0ZIpWVYuxKooyohJ6Jie+jBw
swWUzZmBkIbFXUhUKrgcgrjDJRvVHTCAkXvEibLADLFkhkxPZxzTdcYo0hQldWTKpAmiHbcNjGrs
qj21/+JJHLiyRPB4tPXz7Dm4X3GMcHhkMANp6uXKD1je/FgBHq4pmVFI41MhfTxp+PJs5KHK7rGX
pnMgbDn4nTZHWXWHIEDyu6KsyYq8dYckCc6rqzKqjLklZ/+zvxGpaqdRPz9LY+PUB+lgcYWzHx5a
HgvaYy6ALCg+KrSEO1AivUaVroa7FEBJgpSV9FkwJ2Pa5MFNwHY6OrE2R8bZuJE9OSusWVAUP63z
rWplDyeyL642qPNkRupHHQvVyU00agyUXZuUSpqbT5NsuCyVmOYnNQT1rQGNhPf+PJOy4/k55z7H
X/wygliKv70b3k3Q+yBXaDLEzlyBfjUpb7etAqIMCXcdgfHfvBkNpCGBB2HtiOYyLJaaVwXyDAM8
94Fl3c7l3NOj1oJX7zH7yUcl/k2QodIqbvGJlf+Ojbu3V1HOgilVQy0rHqLibF1B7Fq/dicMSCgT
mULMxGQ4aOEc3SRBYDbmcLXuBchBYhqKhC0Q5h4X/qN5qm3WKzO+Co+abGXBMAztasgudsI6iu9M
deQYTNeP7XGAcR9Ee+90wXT2l7fHkynI1bUTBYawY5TjoJaQNIRAQvnZBdQ4voii2L53H2Q89sNm
gwMDtN/YDXE70Y1HIBjnqXpaUTu9nMBi649IQNBU9UnwvICYikDXk9bs9NED1osei44irBacfawg
Pet1FNfEV7QosPRd1QwIaLZ+J8sURlY5vZB8CKedREaTtlSpIppz2Oi+1x5EUeqEsTPhu9ZOG9vf
B+PuPd72c0fRHRDY24S5B16VdTADgdn1aRrx9rBk7+fZ4cW24TmYMMtps8fSKnmTOWsWhdiCubGW
h9l16lmGaMxTC2hzn1c28z2e0aa0gbYtvNvQ4S6gKtsIaGrwe2MiGA1sz+Kmbf3XWd0inrH/c8WW
TB3lxvqfS8LqJNmBKm55E66KrNGv18qBfohzhdTHwxQ5tFK/FEVqhXKAYAr4hQU0SI7OxfYistEI
e3yxBiQY0vHFyFNT5h0wDVVEFP6kRmLL0EJ/gijzD01rxQspGjOGbH5oJi2kXWPp/liEWxCB95GL
sqJ4xeUridXy4hnExSemYlOga43nJT3PBroVv7NMMB9mt9SIdr4wlzbsvO0DsnFMRqA9A+Q8ePXo
tsUy6dNrCMLGfob9+uMzkMwmXPSNTiSO62JajsPOaGYAgS/LjC9qxDRE7vbkeUU5F2sDiUxV0QVb
RCt8KwiWGRstzcnuEH7cjjQnDCifcEgcE45wSlekvIRZGIlCfZKEADmMago0Vjidb/0iLXrOC8J8
1PtsJ/PUiTpJFyeYjObNKeaiOgaJF85bpRX1rpYzqQuC/dyWFAUSaymAVPrhYulVFaIMtgLDutGl
atXBT98Sk+GNLeQJvVo2O/mvR574lU7u+F0F5lruIZuCISBCNwVRqTQv0RE8dEXi16nyPOKhsn5B
4JixuAQlyaDBSE9zgpFtxJYMD557NRtE15R+jm37c+XObHr4vJMRuDR9pOLfVMX/GnTZxmh1uHhE
97bZUuAmHWfkJaoKO3pnMsLLz3kdSssdvLRAYQdYZCXhBsPhSHT3kIUINiZ+mrbaZnhWUDZIoX+p
3axWc7U3yYxJYK6+R4iwvsWrA96zPS2UU4bovIQkj2CzvusrOrRKYD+ZF8CmA8BWmwfaxpEMbZOM
9VKsfYXXHen7ZYiXxzXoySgd1b+rfsCSbG2pyL9KVyh0QIwrlgbYtmdxYTX/mYQwhVux6JkghYu1
nl4BmndsFwwf/f5t918tqb3O7rw6flP/pHjDLl/1el+um/JK15VJpRys3WpuvgPFpAJV8lS3G2uL
w54JiYlbVijuCr2MskYOKra1pnOyybRRiKKCZ2kpFrlA4ukggr/AWag+AkHQyrF9IuXoQ8Uyk8xZ
2bB9sNEBdaokxXfwUtLpQSF2jC9wJpvMiF8IoxpsapgGLAGmvpUkKfhFOKzdQrpxY98IjH/19D5D
ZtdZf0TFRDvhF+GYSWQg2zXJ/JTFsTB2bozkZPe9wGsMMXTWmV7wdqbtdEOm5PTSbEVVL00k4h3H
PtjNqnebjr53c/cQxYrhE+DW21WPQ2JOabrJmyOZeX8c8vtn/Xnc//hFghdgRyeRZhRxRtvpn8VN
HwGafG60ZK5XogTQOfa4dWticXOIcafh1MovvH+N2OBL9pitFXFim//KUaSsq3oZQV4tLI/d28+K
Hnp2d+jSimQV/hdl4P57WRydphgtPdK5YnC3uZ88tRb2W827kesQeFjNp8izxsukoA1lgERYdWqn
JuQuQBsywrMZHro8JDO4BA/v6MKTGc7Qr7qx+xuonmjwg+rl6cXSgKYef8Vzo8bVMOeYAAZRPuaO
xPMl1ViLS7YXOgU0g+r6ztrrnTiblIC4vfFpb9SqRPa6Uy1qrgMaNjOQ+0U6k4x73ZrbLT8L4Iuu
CkLJQ0GDfwxaBlqqpgeMptaoLezr+bpb8uTBR6QY2F3gCgn40+DcxwjoOg2GylGVMo3r4vBIQ5xw
fUbcYhpRc/n0Hl/dwxEw6O57ZoxhKdUb0rJL8EWUdhY/IDRbfEKlDbPf1lmIlH1n6zh/meCORGQb
XiP+SH06gtqYT4lOohSG2kxzYkKYla1qfxqo3zpxYkrHOU7l8ZT+qCEcjmvNGx5+BRRsLw/GWjMF
pDEbCYZHwPQlXRU14dYG2u7r7YCbYvHyx563wGlEXaw+ow+Hl7I4JK2s9gXFq2nvQY0/YhsBiHtl
ppPmYwxcTC7d8o8dqFGDzw2umSpFI1bIDdgDKme6ZmcpMF7WikYf+o9L9JvYkMS0Fe1D02LZtYio
hV/9jGfSEjPz6wTnJIAgRwNUazwE0P7TZrjARZdwoFTffTk/l2+04svifFSeezVxVbUYoFVz3RJp
SBgtIy+lp77PG6PZGDTkOhFnFAslWSscj/djFKo0OrB/hFtscff5lkccQoe2wdC88IwnnfRJm8RZ
tHzuNV2KklEoQnn9EfuKcl2xAgKOeUJ+SFDZ4O6aKZxomoos1e1mjuQZP4F64jH44+mleqISD0ZF
y/Ym7yHfLyX55Vs+8Qn5v2kRAl+qxiBfEmwiDm+Oo1goOGRPHCxPGHwstvCyfsNaOrQJOer+Y5gw
qmpS75MlB/Mu8mQjq0O1opj7PnidzGPx+1BtUM4M0ElAcwJLPtFOJS9/uDZQrfwlZlFSuVjhcGrL
ofkGDnp3TjoaE9Biw7wwIKyfjqA5LAni1egv/0bDbnj6PzcwN0yY57Or8d/1uQZrlXgG/koRnzGB
JMfkCxIilJsegShQILA7hVDZ1lYlj4ffIm01gsoGJlhWbYEO26A7WOgQVgNPyEGeJZCnlV44SpoD
XqjBA15QW0XkljEs3uVnZQt5KebuJAHWZkpKuz8he9+yunmAQrURBbbu8HtChKUp4OGcw4YzrEu0
uk16Us/t2Pa3JwjsbGrTvm8safbeydJ3DRkZJSIYIRVYOUCc8HzrfYJ9Kk2hChOCyXjoui+DtqDR
DPiIQYg8sTRn0yUScmvPnuHiNyXI1ZxxpILp5loFWohdBupsfWyhWDLEthwc3r1YsDMiGORtlXto
GLiFdWP3JUII1Z80WIYBg6mAMdUzG6pvn1HZRUgnqty6eLG7W6fa/Qy/fS7ivo8RU9T6BkcctRbc
ysTkd8+mZ/s4fMOXiJcBNnfW4sE2bhwf89G0HFidVmGY/+FObmtAdsBuJU5LFITBGZoNN426DeLC
WRhffDkK/08le2piPalRCulTY4YLqpf1EoNaVRBJuEcbwxgFYUqrd/gCM8dWNtoDqX2SOyK2Xg6v
19ixVA6x9WO8vTqVJaFYGRVJ8mif1ON43CR+EKq/7n2IG1iIoPkFWtIZyNoBF5Llc+a50TsyRS8Z
Iv/2yBsP5uXN9ahO12RhLF6kS9pDwx4d0YNLfgs/LmtKRHU8tepnQch8ammt+HrFI+H7GLHfKN0O
xPadjMTWsz/SzBQLCqDBEG5rHFJFzl3i1Jm54L5oCxhDEtSf2uNkiE5kYmIEGe5NFbmLbdEMoq/E
idg1EWOL3L9DQjcDc+2VgtPA++aOf/DkcNmAizmnZqyWz5FOhxgERaAtatvQhYNmf6SdEA+ffDAg
TiPKxAnOMc0O8g16IMMt7uh6L6evf3owpTMV5lBNadUPWvhBvUfhV0kIpSv7VEV1EJ+mbXwAVFi+
zDD+yC0PEiZ9YXf8nmLBtvktq7VQ7a+3Q1iOTAKlIQ5jsoz4etIdFrTDw5FZK3bGfHmnNIDbiepy
/BKoRM6C/65Liw9ZkLhO7Pac83L4oVue98eOW3xYIE8szybPLrMkhtE97N+ULgJ4qg2uSAncS4sp
Uzd/y8o/iBqmkBF84pPuCyNYcWeb7U/jCGh8ljVu8QCbhCDy1EjmgHC+PLGuOZLLn6RL/OxocmJC
7NcR3wDSsGPwSzVhxRGljuatDWY7aQjkTw09Y3UMgSe8WKdMzLwsk9F4oIROJTLPryOJkSed4soO
lNWfD3syvqCG3y2jL4F08dtznwCY5YCY6CF6od3O2lKVOcCch5UkD6YUpLxbzrve2waeyfOyBmm9
V9Bo7r7A42PS061C3FUV9pdY4CSwN8DsVTQe+Pk+m3swt51a/eySTdUEJ6/G+fbUiuq+P/W3opf9
1tPICsnQAkVyk12+xMZ7OPUWHXv8M36r6tmDiMlQFJV19bqj1YIn1Xv6L1LOSGO6lXeNzLcHxjpM
ZH4tPU4wZtyGOkbtkF3xKKIEpwRDVcuBNwToUyF5MT/MHreNecwoFwxOtwa/TIRmWsHPEtjwtU/5
GliJ51YqYFmRd/DiqseKukK78opa3OxxOHCoN1jltKRK2jLdh/JMaUiorm+0T7aW+C3oPTWedA+N
9YqHJMh5bCmBmzDs1zzIWjAJOCi/OP1DccVJFrfkMUM0tzWjs6+JTjMWi6BOQbFFMffoADYu2Ca0
wig3zgR6lnCFDTiLLd70gVjIUM0m51/hjiK56p9VPYCB8VKUOOkO5uikXtYdDp7t5XrYjTSQuseg
UALsswjuVwmF8QC2M8DpraCmUsyLrvNKPNlPFFzTlAgMrpjEsF+G6LF7pnHLDmsgagJ5IUnEVg/6
ztsHhQRV6U50CYQxZn5C1oY4L07YmBu1f2URyOBFO7RYgfn7U0I/9wBkdE56nDfoY03X9+xMOqXf
/+a+G7o1RT5VNpyiXf1bnI4fRTn1fSLfQn6a8Oj3wPh/wgxlu8WlSeZmU9gQxBwnucxCDAbFRtse
utafC/4KdZE4XtpMpwJ+HbCVe/mbdvaeZa3DbCFn2/i0STA7Hl0DD68ZuNsWI3a3qj/gDwYeHQX2
9r0ZfeXfk2AHClNdfm9IJFXx6GTFFknSBt/3Yalbv6FqvtWWDHHWXyajIhR14QXehqTWa49w4s0p
j7cX5jVZsm1RnmednEB8yJ8PYvK3I+08tAt4jnYfj2f7+1oFtd/zZoF4NcS5WVMyQJAc1HqE5RPc
cb55/Y28Ig3ETiSp0lGzIkjBv8+/56eH3CDrpOgJ794gjJn0wigGiXA7JKfbqn5jj9ngKR/WLlph
MueT7QnRk41R7rKm02s9L9K1e0QtcgiEWnr4nAWuuyKRY7LJrS4EhqcgjLkaXejU14MUCsccNvZg
UmpFB8+kaQEX6ABgHvS/m6ytJVbgDkRb723k5aRpOz0KQd1jviGHf+EE1gLcvjPj7j//+QDRlF0d
G40lXTw+a/igFSDVJd4frc+QgqMDZuXU9CJfFYh+8Lfq7BgHfltOhbYcUG+XRNbNcXDaicd4jokC
W8BYNv+6VGFzduP7XEFd894te74L5tHvbUQKzxvSMVsuo2fKGc4UIB5eEiHZcQpfsZUCkNK0vJs9
bUw752k8D3UhWCmXNXrGj/drJp+E6HQExGyWtZvCGZFZN7A8SLsBFt+eDmFRUzXc9NoKeP44DRy0
SvY8J18E3igj8TGotxZWp8wDZ7g8tW2y9O8OLHYD3tCyn0BK4/Lu+1SYKZq3fVDgCLgvWGWrrmvh
VRfKKvJMTMh1prDvMwRXBCxktInep2fKGwcYG39a1EeNSzR+WxYa98cFcadaQaFEpwCQmknTnUhu
zyvX83mCU3H1XZirjnlRzJvyIjX6OpxiET6lsUtYjQ0im6ArXS2wbG1/4FPbfUxCPJgNjJYo+dym
BhfY1oDYDyFmPAGGQezSXOGzHP8Hp10MPfcsMH0Xbza+Rzj7MUfsK7ns/pwV4OdP26Erkx+qtUW3
SR5k6eyZmgjkCsXFRSVzFn6KiYa7nik3UGn+B9917/8RWTXGMWxgF/5y8myCs4vJTzgHoy5doE2p
K0a2P3o1L0/uIFV6NXRGd5JUSzQIigFSkH+pHImNtT3EeUePmk1ZOZ7XdWq05/YaMXQkq23iMbRR
2PZlhrnZKj+kWhYJD6M0V1zfwMRe0yDZt8ANpshECVpQ2yHH5oUIXXgcYsQcnIZZfkks2Oa8GZ0H
BE7F8uAo2nVjtm7nehkOrk6hAitdx3agHL0/Anaa5FFcCIa+Ue1DANYWXMGfnbqNcnH/pApjsc0W
jsODUVueAFzXpaoNarC6rlQTE55BEtImxsZNR7TNWCNA6wmo3Zd8EB+znxyjx4Do15UyFkCpQRTo
gBW5FQCQrK09pV0VEjEM3fvepENeLzwLzC27QEOb/HFGn0o/z6ltbMiy9QxoVPL1d4mIWvVq6hVb
cVkhujYsvVTKfocUPdDQKMGeoqbs/V5l/8TMOyc5tDDM2w14b7YHjzJvGtf9Ag2iUK4HlYs8n9sn
x+sIcVLmvHpMnXkCvUhed/pO2NQ+Ar7cUpfZ5w4ECwkpQjzbE5S3Y1DgZSYHTl51HVfp5AKzcwDp
T/PuYUaMTwCLEXAs4DsnFScQIY+zOuW6jomyhyuTJBvwEcP3wIzg4dfsOtdrLpsXN9bGNP3kfyou
XK1bh4iogzRmClthCvhvE8RmIF9hW2eOWZw1cAt9Zhq+/fCSRc9XFzDv4M9JCPGGVq2cvoY8BhUO
dwj+zYR69cmbo8+dVrUG8jx363c/hAIGqwSCoYNOQ1XXrYvE9sJmpZQ7mHva3/DNJjwiWe52Pg1Z
dyhNthOjfZ/aAQQoqqiA1f9PPpxonf+HHg67fBBoR8xxK0YuOCM3RFN0gKz8+uADtlKDglPBXfbY
clDJDlKKfYTnOxSwJq2L7lAm3f3xb86driv0BgPdeZqRpCdnonFQZ6smTpOPdcn1Srs8z5UCN/Dz
JqDNvItbPQ8SbIkXgxQhmudzoRa/jqHT7clTQFUsZT+2h9AIxB83kD79aaIkcSOhq4aYcBuQv78F
UO2RSC1Dt4AeWE6PS+kDRuFTcb2X7EmEoGw7+KE08A/zw3lDn51RO8//lesccwlo/kl3fN9oxBhP
T1bPg8+r72NyBLrFXzqV5if4EEu7uP0bL5dORhWwYp6whPc5rnjpeV/e35XZwDsX3/PKHE/cae7Q
MqrWcpkDl+CNTomEfmIOzym2GWO2QAcJaiEJhyVZ95X4gtB8U8vxRkLls6/FtphVgUdWZqYmqH8L
7AQU4FNahZZysN1iCWejVmCGNa1KbvT16Gc6tHTpyChByF6DR1fyOfNbRGM87Nt84AYN7NpoqUEW
XEiQxXaTKfCF7YMbTL0wYhmaTydjrhasGNLJL0QGUnhBIHEuEe99kHETJ+9XtqXgTPts7o7S6MSi
FrB3XpalOxsXVX6PjOL0e7XrfUfDxIhuQ3uCwpHmSTzYxD0DOh47CC+K3SNkbBnZ/8D35UTeX9aH
q0ov+cdqBheiiqZmxUBAWGW+WsQjVMlg6yLPk16hd06TjnShB5E9eDo868Ad3qNGcH42ykHWsD5X
grn7vWD+KTXeuSTzLQw909UKgDjUyh4K7d+2/Wc4o9Rw6X1zYvd8jGajSpWEBmj9JCg2rtq7bUr7
TveihW4SE6WuSJ/DGDyXhVE4AyxPvMjCcKyaQKQW0OmALinIeKnsqLiYUX3V9vjVFGwm3Tq+WeyP
wtSGA6vkXDX3qAgHrz1YztFsQeyRmKAt5IjzyCDw8PI/P+VSY6y3aLDJrl81g30mCSN9Du/WWgNc
jSEWu/aKX3TRZV3swtWM5JFfK52whNe0wXa4hLjmg3VvvHBZGf5cx22u7Lo4DRsehjYgunXpuzql
kmGdGqQ/VvSlK+U0LUG7bL2799YGFWFayWwqTHSnBmDulfUInLGI//rXwOId5wIGvV8MqJdJl2Z2
eomrJmoOnD3OLYKc5OHTwuPXvdPCZH1LIMj8CQvCzOGdam181W/CBuUEx2D9cFW/oNIcokYXLE68
VLDaSngvLoO0gl8g2rO+0P9mX/3RvjBel1pW+KfETZHlmTDbkeETVrFba/nCP+RBT+mdJv/4frez
Yue5RxXa3JsVM+R5MF2A2ZD+wBhEJKip0QieSYgWo5GKoNThbE/jOQ+OOlsAOigTqR244hc30RYY
KplflPOmhrGRLAHpBD9O4OYGBw/DrtHPXNvsm25PtbUpf0gXmKfxBKw++Iv6GiQaxrDvQhNVAOBS
XCL3gx681x/vRJ0ojIZ6fF/LQXdu4x1YhOOcvi6Dpn1CjyRWP2tJs/JGlLhGuTfiGNM/sw02H9Xv
wlgKdB+5EywgTv9N/DKBr5Qk60sFu/yCq5pHQ9tT0ENofNBspzxDaKeELZrYjRcQJ522hhmjuJx3
j40ttMiYKAGg4IrPA6AuJoQnZQ01FG/qe2ZpBj89W82FASd0CBdBPdLMacJwkaPqefrtBABBaPFN
uUKAaisz21BTKXL0thE5ee5DEpFeyABtWfDIm7T3OHX5pe7jrqo26QZ9Seu3TyUR/89iWypQ3tvo
y28VdeQ31t3UjJlJsR0ltJe0Aen/shz/EQHArf5fVK0XmXzePNDBzkiCw33u/RLC7gatgCo+dhyS
gDIipmOAHkbH8u5NmVJAnJYYvcoeyddCSen6ke5AK0+B2JBE9LHQYhwhbOH9r8BUHCylu6YwrBRV
mf29wGyKSfI+qUxrDPm1WTOtxoqVudrYvf9GpkMA6KOvRb8I/SBDXKBcMiHWIjjNmmZnkDJh7tPf
5RfrWkcxAhgdrIxpDGMguOpOyTumvJPUdSuB3zYykTkUAzQ0xJ5Cqb91WPi9aSgwgCJgYDcOiwPx
cFr8+O9zdQKjQgXFxlL6IwG37W34QboIKMb0hDL8syUG0DrOk9l/AN7Y5O0xe22M/5bICqMa2fKM
CxOXlSskq1MLtRqhtM1NwjKhxuOfBaK5RF33Vu4XtflDrVu6jhxbf1WFKZxhShcFnstjd/3tINaa
mN6QjKpAirpHdnON4CPxjVYEvCvKIwnpZTe1b52dE9pggrx4skhsfhVY2RaZm9v3yPBLhGUf3p4p
u34r35QLjqTKHR6wkR8eEz5BJ6aThaqrjr9QwvkraV6EHtzWWAB7mIWKDZypFIgJ/hm9Ur/HL3PK
bOSVOfbPYwZ31Ua9W66dk/oVeMnpduS9iDINVJR1V6Sc8tkvB1fmgWW9UlYLgZ/+yFB/RiXTRC46
72dVRJDlPT2RVz+4lKkIM1ozwWx2vZ/o6fiuRFexup0DR7C/oPu+rcq7zaUiKdSuRtfcUSASPaNO
WEn5JU5C28vd185thgPZ6sCEf9HdFyO1H2aEbg7ztrpgssQc9Ml3EvT3ej6Mq8+8i5kzG9naaU/k
EYv1Lh8ZlkkHLzaiXLzeG4Iat8rgN8pmqc9+ZULGN7ho1/VPMRLTRNVCNq4dVbX6+auJfvZfbmZv
6dd6wrE5gN6wg+KaZAvz7tORRla6rwHCkE2E17O80c9XRPJ+tYkdcGL4FsarNvDD4aWUZ57x4t/Y
OeZ2bPPoZ3UoHwDbLffkQPDYnteLBzOvc3fYiIiM1Ud1TJu7dQ6VgyB1bJue/Jql8oP4Krbvp1df
xRXh6QZGqGLjf/0zYW74QR9hypVLZCLpWwpCMdCenFPrv50XhRkmTBjG18A/Y+NNmjWFbyos+Kns
pLbczEhUgLhTGtqZBE4/KdwW+XmByb6XjdVxNCP8+wmhi8aqT1Wvj1yhXqGfa3FRuEo0FJTjt0Wh
X3j3fEqjQ2tKfjL0JxQmEod+X07q9tC1+LVDgceeTA9IYnO/i25r9aS4Ly4lDp+Zr+wfeOgvkGLJ
U+N35XnE0Qy6nb5UqySVFAFBmiclmvUSus74qGA3EvIVHQ0h3Oafurj4jB/LMK1wTaEDmwmBNHV3
647HhAXo/FnWFPIbohuQ9DJcnAtmeTqRSU7eS8OFz1efv6T4nWlbQ2mixICUKsQ4Be6TfxHJdnOg
cnUiFuxY6qLe6JXIDkUEtrLn1D063xiTAwJKZ2GnEbmrrrtWIJ+48z6qZx0t9BD8o3cDh58XVxjp
LnU4cTIGInWDO4UZuTWQZ62NH93mu7ilQyLBqMQSlMXGs2gzKRmrzWZYncAKWXvv2C104xuq5Ay1
oZcDiidWOYHpS2xPfsp0/Gb38legKd0iT/mWoXCX/w4sxFws/eujH/1yFLFCxH3DQGNXQ6wnWCp/
AEsmH2nJcp+DHelNhicdOyhFOHCxC6Be7mrdXLtSBgAm6mF+QgoP92d4cVqvtMYzzo6Hynvzf2Nv
a3Hr0Jpb2Gl9fWUD64E9le0B3UzmNThY8Py09oNtNkywDDN1RPlzeN69gf7qhykBV3lOF6IcmGMF
r1SnVpYm9tvq/eS8hovPKcVdcMJ7lwRIBhmAMe3sHPPdX3Or/n+oKrSj14G6QUxVwQ7P0lRSnGYw
2Yz2+apS3tPzlT3PFSCn+Z+EYQIlRUPaKR4dCwa+IojtR1Ishxo+OULcMvJK6Cyr9Q45esIPTSyk
N9Zlyzsp3B3ogtYUysilTzhQkz/qs24KTIgjqLuQlaZY9RgrElAEafgHZc9OVG3uUtbr+pX2rPlY
5BXUi2N1If9ElMCazh0iYTP/QRU5qNVD1jIlqRaRtP/jKWIN64PPv+kdFKkHKHYY1jdeunT3WFBj
XRc2X40flgqn87/uwhO+CV3t8M8f9qvwj4G720T90uHJMLwh7KA2DvUvDVd0sAn7Syw4r20/2jl6
kdVGHQ2bcDQAsAKKyoVDhE6RmGsLtNFlaxELkjE6G+bjfkPOr9JUzFNs4zKhdg3sWXiVWGsnJfko
mBT7HWYUADNnJWwDJ+MmPx7gIrscDDXNVdqsj2eeAtSAXaj1wuE46N45U0MOTVGmh71kBB47d+FU
OVuRd+5RzYF+EV06F/70qpgEF3xzwig3v0vP8YdECGs/ZM4vGPO8c1u6lWkdlvZvkvoucLHsHLn9
FLN124dk/hNPARFy688ly5cZdyZV6IBvtCb1pGnWL6IlnUS+yJiRPP9AoE1Oydqt64vLQR+plYcK
+54kz5D5ElB5RPlH8qQD19huthickYorPv1SuVshCrIL8mwR0ADm2vi1KS8kAjiq88ll9ol+QSEW
wbk6BTDcR+O9tnwvpslxS/rxdIzpmV7M+dCBR9AjfczIl4ol0fER8It60dq9XQ1tIPNAN56zwFy1
VzMcc7WLb3aNULxaxpWc04PO0T4h4ndQwJ/Et4/VMJHxsM5wBMX+9xxTZHZXclC18m1Ezm6m9OEV
t4YS3d4ZRkmhaMK98DF9BiK/D6tbNRuQg+lcDGc5/yUpCo3ZAbjxTPzkK6Im0aXokEsT7+s7KUvM
mVA9p+uqS/GxySVMlC/4BXYWCZgd1a7cBuQhaKPRy7zJ1YGsjr4FMx3RWhLUJLJKvEKLYvVrMVeX
16269HqF2LyeXEYI/JAuCNyy2TB3MiM9lhkciN+xpBLOzM/HccRzZlMHiZe40h8X9l2PV5sYD/1P
fXR4MstPadaN0yVfuaF60o1goLvrny2EZ31R5HaxxyMF/2j+/DGeMxYNVTL0RCUOsw5Na3H5uvBQ
HhZTVPHJsmrDdUAc2s396TKH1+r+tYsnbDXOq73/ufnadsvKGDm/r6cGDuqyW37PhICtKBXNc1Sf
kRwS5a7ReyQrLyHlDdTCYXY0yN72wIgMa3FWdLqCvCN7pmkC94c+xKzYLFB1B0yDy9C4yhDC0WU3
8UMw0/5v4Z/CVrC1L6F6aINLt2SdfqOtPj9sECLsbmR17R2+Zq9ZIryHRR6ZNPDIUgCRSfmGkoqm
YnujUBP9yqcoapGE63R6lFOvgnHrxYDfp0L96r9ZpU66gpnK8A1mReCJK5WxmYvPXiDZOWjsHN+8
CzbydzDWd1rYTLyXhCmJGZ9lWKJlONA/5fhVOwd8y5oelGQbcqcRbufiL06iqcfB/Uu07EYNf2vU
Uj1Hkhv+umFAxzl/LuxsT2w/NfdLfOBQEA4PQtnMSzBcofXoCpZH5usrAtyh6T4i3KtspdxR8m8U
waulvEUra6Um0ouk7clLSOOaQaNVRiSQS3frDYaq0Ofd9Dwcm2VNk9+EUDS/yebzT+8VJfDd0tAS
GZYXGgNO7LSJng77pTIBxpJswhNm/Swvx8ulupj1R0oBiEsw7/NrxWCaiTf8PjhjsegvVV+Upf/O
gqn4WSCjVtwLJpmQMNLr+Vl4hLWqakT+KCtyvwt+ze/uwTg0+OKkcbLn7OQVENq4xtSgDVCtwBac
XYwralqp8DsQ3hllgBJDsi5u/b6tvZQQY9SSABXrnncp/FZr0h79DhA1ruqO0yEOye9EkEfUIobc
RVrO79RoIRZ0l/Ooy7QWRiU8PvJd7GZ41sCgNjUixk61OgzsKdwxxrOdJ7vhdlh6LNPhu+Rmkz1d
aG63f6y4q0Zz3CdKagW6oZI6JEzwwOKx33EdYdcyFsCQg88XTkxI8zdvzAv7Tz4MPiqg88bvQ45Y
O5aPMbtF4xkDUDnp+k/t7xBQdLxnd8pixjDmXnz5AseoAOWGyaN7RNFdFMPimfbfyd/ub9/ZLlob
nODnfXJbqJ8scTJObBqZwbVtCnHov3gi4678qPZG2nCmSc9H1KbOthWQQ+PJ+2ws0HDBmMJGCFA0
fYIWw38V9o9aRmJYdykP0G01yocpZ9/bo9rhe5M88nPIdK2GDGLjH5/aG+25VyPbkxhO1GSqiffT
OGifv4rw+9bZlYaGQ6lZSW3Y94eFUwABBwJjxsJDIgnRB3yaW5QwaQ0qgF6/svgNGZAwtq3qrTo4
kky/+rgd3UL7DjJ1Bwf8o8q9aedm5tELjTaE91Y4QZpFwIf2DTSuL+1YSEoUPgoJveRRZ7a6/Pt6
IqmBx3G+20g5rjFWyqFZUG6xPlDFGetnlWK2yLbscD5smworyieW6Vdwk28xECTsPl8PKOhT9X3h
ZcuIAqGdUQ+JA97B3VnF6E56JwzOedYdcW2D2iD+WUaVxibS1ZSfA4LiZmNbS2VXHUHiwVBbnKWw
i5Xy1rOOuSq8i0B+LCiJwUXna+U71ETemvMua5Ut+CBxyxgpyjB4cxE1OXijA4G46QFHRAm/GThD
gN4ZZUzqKif6HHut2JZlsNEHAsdNm7skNAYb78g4pf7U46zIqsy6gWw1PdqoUfv+RnzerPIYe470
qarMCP0KNcVy/0LjtI/vv2DiaStWqdQCgZX9dZ65/28mlAz8N3nmY9safk6Yw3YRR1xeXCuYn2Zs
IIAGVT9emVWEkf1UifVeHSM3l+nnNsj+spssrseZnR/ks1+x4MzmjT+esRmV6GpG58tfo31Vw1Ig
ACjPDzzNZisdxmiszrKXfrQ8gxH7Um+LWT+Vo+zZZlClXXtHne0sMiuT4NnkAv4y1oL2/89HAai+
f8K05ZhiOtgnlkcIv1pOK54OXDrVKWFWTDkyz4sNzlTNAeiBIykaRUUnhkDNIgsOej8+x8SGsyZe
BdFH7Bu3NVanmVUeFA25ty7/khsQ0abA7n2/prJ+ZqvyqVw8mI6GApUt+bIzGTa5UfkvBqs3Qx7p
lanuNwqfeOArqI+ajjndx0cD2Evn/ENCkw0hRH8gsED3FbIiwwhQRlimqk71dzrxRExZPNt0REuT
28pXwq7J2xtj+moyjFEk1zG4R3uhYXdmFTACa2HHg4hv6Dj74T6BbQBPgy/8KNTGnRCjS1nri1Ri
Bq3lIU1UWj5Wpl7csD3W3Q4BZY9QALaJeqDKWMlys/xyyRicSwxrBzXiWYnhi/FlHNG01/49F6Ej
0GbbU/Fr0NrYqi90icVIedM3C+fhy2ooNE3AuxUopZeaYT4QtHUX0S2KgvHtrn9PrA7q8rr9H7pl
KDbjAc0+jpcxuDFmrhX1A0Bn5PprzHQDqKLOIYOv8zlO4U8tWb0ZjlcVPt2hd7OE8om6rGt1I6s7
r+F9LY7O8mWVkcxj58Q5pCtcTYcHd8pu6Ld3qGt4Liy2oLuPSB96xT2e8OG5x03SoMTXiE1brIQS
qht+rLDzaQPOxrhQ2KjiBZcstwSw1FSk6b44iPawjL7JbHUvXgM3nl2E2Jsfo9IydSl87yt4nJWV
VSkO9pHHiK+ON/+SyaVkkQzDEgYpRR07Xt7PTb0Xp+v5Xzcx/R7quYaVNrIL1N09Q8eltVgWjr5f
WWJ3Y8ZrzcIfPhw1TLT6cnR54mY2O83TdD13bpIcQau7eWaYhvV2+r+obL0mRd7NqwkSAbtIPoxg
ocAmhJniOOsyEmgBeXBrzGRk7MXqu3ZXsTmQhBlc8t5ZzB4xv7mXnCXADoF8YwEtvu6t+FEMF1BX
YlG8eoVjnJ5T9bsmtx53zqVAJ/sy18RPecU4z2YTj87/3kPLg3k2bTJX9ySRlMBX3iERfScFwYS+
TEW3ZFjXxXeRaowJVzZZbCywKlgjIRDs0RxERP4J9WnVRCcuFSg9qXZicFzZhNMujteoa4vfdamU
Sz45Kb8LlvkOB+I/CLkxurQJLFAG9QzVaOwtFpxH8YhHB4eciL2O3FIEODnAytNhZraFIb1yhEY6
U4pr1wJ1yUt5w1xZS+RoLA8kXDNQNFLUmGq5JGJpXvykY49bq7VqfCYnQMGjNi3M31jhMJ0cKgSi
erPd+jZ3sJ2T+0yZySHJnBYGkl8G6G0l6H3SM87DvEFl6DzLAEhM8rYH4VbkxO+O32kSpNi8mHRH
zedyqgEG/Wc6o/i18l/uAAch8rHqYnGrQsWJv2wF+mpVKua2i3NGUR7b98ElXecPFUyzWgZUrsDc
TqZOqq1VCD1oG3WPgoxiPhHrorL4QrhlmCJ6NlixDsvHL3KQNWz89OLlDLpGE6SO4guEwJvSJ8Sc
WuZunPhkx1nIpk9zkxlUxjaj4Q5O+WNhnDIBI3soNhq4ynM2yh4zZBFJGptOb1ad7+V4dPQyKwx2
ntL1y2j4St5yh80DO1hknsEVdacUbEl1IjRD75ermmpPqFpqBi3lsrYi5BoCqtpJnjIVNDktpUqz
cdSZRh5GcdQRiF23W8VJNCr8YnIrzAXVNZiBr9iL4pvl5TTw7UmUX3BEEUHxl5NWFnYNcGOFrSCA
895ClPoeNy8foCggViAh69tCWutuF6TK6zCxCNXCg5eK5mhTpZ3gjteB9HNoxKQW9mCmf65E8sUb
X8MFnHHtCnMq0T0Hgeu8+32uWkaPaP0YrzTFOXNGn0wb1rRDSvSRCfv75Anma3nlmAPJeH7fIA93
cFh9m1ZaChwqZxA4BQtGESzO1FZq1JNrL1a2EfvepJim27B9OyY6lD/+yeTS3Qj5Xgp587sqMyci
tp3rAimRboRSu2/3CwilNKB2msI2ZdIyS9DFbXtPKPF76fPYEaUfcSCdqhMOjf/+tcPMho214VJo
5T7CINtoRRVEoSjONIqvUwzpPHvKsa/JwO1OHP2ORkmyfunIKhavGr/zhtNx7uiOv/zR/X88Dig9
Ec51usRTi7CBqNvMXKaPUoHS8aeAtms89u90SZdITY94Qtb018RuNSRZwWu0rjyYjLxkatRzOhd9
Z5DWKsVPFJnAYXpMMgeOp/BjBpqYfthJrwyu/Zv6yHB+gZC07FdhZadBESfmF3DvfX10/KVMWVTr
gqWf/uD376Jn+ORCAJCK9M19n/ro7f+2wGALktGLSMfbUM2156aOYWE5Yeu1C3m+IRzIhGeZB5ir
kFdTyYaiAVedYNvBqOVTxpCVQAsLaAZyoJWKrMauTPqatYV7SQGWqjxTFAFh8nS0v59SRvmklWj5
Br4Yyf8M1yxBorDsYymhPmBe5KUJuRsN3DWIqcWuO2wrO14rhprXlxStZW3+gxSGtyVLWWItbUhS
rVtZbUQvlKKosdpLlGhr2dsdVYDI4Gqx5SeaXtDYbmRqj2cni5hZZ9d5w20eYsr5/Z08Y7Hc13Tx
orxLmeiXRXf/O3R7SYMei2dIY9q790mdjKlNeCEw4DGNgTPrsWBqcz33QGwusD/Bs/XCSRnh7c/4
hmIfUrWjEuub9viM6Mqu+ehxl06C1fdLuodsGQXaQvR+MhYq9mgWi92GNGA6YFvlDTrMmFYzGtWD
sde6wzxAhsjsaDLEe+WjAhEljphu3n6/b6hldOyN9lD7dwQgzmJT7tlJNeeHlH4aQw0l1DVvd6ig
PUxF8OHadRHm/7idOE6SnScs5+/IcwVj+yv1jwVlw3guPFfc4dlzGk4jcNeqgqj3Bs6qYpuVLdfl
yVblD3VLWfbrDw8nsmPO71ku55j2B/LcHN2bt1eD1N38tub0rSfGR8rKSJgtGKM9B00JSSNSZ3HI
bfiGvPmCowIgMDYW9RI2OrMmi2GdugKuWqqg/JkbXYkEPb8cOV3W8npJIisUKGEwDuZVwQZPrNrL
NQ8Vyzm2hRi1aNwWaK6hLLBsJanWxzFGwHEfpedsi9CNGNdwxppXsYxLLJhjL/JGyJyANhHY/Lv3
gw2DInF2ANKiPOb+mybTJ/3whFa/K6W4O5YlVgj8tB1u9weBo478nrjIb/FxDorldX77wHGK2I3v
qQk8Cy6J4B9AbEOMqOdYcsYRBGGFoR9ripYyIQ35xQ2lhNWzvOER2CCx9cLYQCTjbG1Vy+FxuOtG
XZSOaixrIkCYsqhcx5VpgN4TzOVwzN6rtni7IRj6Brl4bM7EyZWmJ3hp+Ae4XbpKBj8Qx3xA/SxS
8uo6fyafzz6thSR0+lbfQSvrqGevzZJCXn8KBLZMKs+P/7lpvMD3j0QG0YlPLuhhdEFTr9mz30mI
aKJIMrGlk80uuDgo85ibWIz+b/KzakTBte+IGsuUXf9+/5HhIES2FClG6boh5ggVv2FFF7wSuMgw
2I6X9akO6zpPcUWZ7o2BGuDbhOqb3iYcuM+jslf3WEzZv0UuKQTMHYYxep7rkt3Jiogsa6fglro9
fYDF4Yn8gBh5SI3CIBghE46R1mchosMEmSbDHpqXXf79bwsdVE/xf2S9bxCtKedslTno2tmn01rt
TcQTj3yF1dE83CrhG9IVgV9u3caU0QijsB2BR8mTMp4pEtpCOOfmPpIPti9G4prU0kyNuhcs6Dqa
Ug+HlYxC0u7kWChFd1y5ot9Hu7wCLsz6Gb6nF6XYKeeKelN6Ts8x9fuxMgmCzSqDvwtIQAlcGZzf
w1P+jE+3jLzUU6N+ZDw+8Ql8l9CFtvKHzsCpHbbzodf5R7dXffsQ4g8Ji+dy4TkOKa+RM9nfbvqw
Ntf09PkLXY8PSEDGOSXj3FBLpjufgpWlKsOxV97AOMZ/zgn5M4X2B2s7tZ4MWBvYLSc3DfAdwLha
paDsmHWdPo9jHZpbjQt6mVqDrcrbDlr7pzTdiIZ6ea1mw+DZS0wEVFNeeDj7LoYKY5Ufbj598MyA
XpN6cmOH0lCCMErJW60VNNKNrYGFY96TmVpcdtBwqbJCCngd0X3dKp/U7vxyZjmOMkR3QOUZ8AL0
8grpQQeBA849x/xQFTd721SkSC967G5LHRvUW2uySpaOMf3SMBf0SWVqtYsY+7yTqMC6BEySMN6L
4Awpa307vFEcoeFVJ8qT+KmsYvdXrYlDq7ZsI26Tolp5bfQdeodE46avmSjnvpKxwpiCeCQJs7GG
m9Wwr2C0xmYGI4YVuewnbZXmCd6ZqvBcJkssKeDZOq/4bU9UXIlOdn0Q0gsfIRzCJSiK8GbgH52Y
LI4JF96OXFjcPvTQApe791BBR8R7J9D2191VLseMmLRk77M3PYpyNRsTcyDeHxm71PhbiHCXKpI4
kMBAO1MWJrk1il5Np4fQLTT4+i8R4iI5Ay/YKV4okslRWqWZr6qgdXBl4l4f3xvHqvG8I+/xw+tt
XKLjsNqwBkykVR8150cZTwnIYld8zUwjffeHrpMjWySLRRXho1gWzZfwXoKA2hFAiVzTcYFGhlt9
kRZ+EVcjGGobaM58bSN1PoIazWfjK8QabHdYCvXm5XcWt3FnlUx9F7yCMrz0+6n15XmVDx6dX4bo
U1L4RIask6svzRXCUO5FPv4b4lYFWSLxmjDTrkd8UmtgQgvDpzmEYiJDyYTStm36S0Ku/ijjCUV6
ap6yTHWk03j8vluFBL/WtuCz5oVBw6NBdbqhYUeM9pWDMbwgGuO8g/ZKyk+eacWjKM4Q9Iogtrmi
ZM0UvkN/oR9X41yYCI/25/J5RZT572ioQPG9aDl2ESvmbNo+xNmjtPlQCjv1BemtyQEi6fyEiLBE
HXnJFIQVdQhZEdqamizATWltzveP+ZBk8Hg1oJMwJTdFZMb9wSf+nCPtHK/Wpp7iN+h6sgf0jeik
cUMs33JKFcnVgx30qBNMdnT/UJceQIFIEzv0/qE73xNFqpt4TALbjTskNCOfPGCOYWYGrEHOxJ/q
BY4v08KjTSPGXKtsmZji3Z0sRURQcQCVZgnF7+SIeXHze3Wzu6cuU/Ace06xEVQNiwXTVBv4LePp
586Y76jKce44v2JPUFMJcEZjY5FI5k63uB48m3j+G2zuGDdSqm1lFRWlRPvefLmPzgcvl5HglDqC
I8RLuYbX9WlPmr7tq96jYMupG5ik7SOxrk1yn0l7XAoxKCu628hP/Q+irL6gQIbrcY/KclyQ0OWP
xw7XKyqOqZgHzAX108t+xSEdtDsXO7Z4wiOX6DWBh3Bob7T8OSDHRUbjZh41XvtKTXQ18azGqtvM
ITZpZpptv6Y9HKH5QXwmsw0vW6XP8Pow+5UsSHX4jkGrs+4jhbir0z1XNvelOpsWxZxZZJ1q8XHZ
5IjXQHj/48epKQceVU/qScbWJckKOehjIpoI1KstAaO3GQ/H0RYkQM2U+hY3kON0s6YIyEdmgvKv
1csXSeQm8k0xYQ6BIpPbcPIfFK8ZH/0N488YNJi/Uei7nlwkhiDN/TBqq3pYQ3UFQHn+lfZNYs1S
+/jkK9MuFSmklhmJyZn9osdlEfFFpU1PH/ydijae83MaXuuUN1dfi2W1QrYWTkJ1exXq6A04v47F
rIMYv6SnDrjeuvpfaMPc0D/KLgQicRdXfzvWR6enmOS1yuaqITapdEqAKFxWXbcmuQmQw3OYAWb6
PBffB25pUZIvJALTZSQSWHhecDCJSC+OjYDsS9To5W3xWilsmt8dYXqnq5vCEBTLxRbsBemyzj7m
v0RuobLkPxyH4nuZHRrkrWk2xB+NsxQ59nAzkxxrppN7/JAgEnFKDQShlDnHOHXN2hKLFC1jqUgv
zxrTuZXL2e1qXLFEVNkJAWfFTJINYjprEwhGZ5nHzVCOs7Lh+V//mTLuug+p5KoUhOlTfE2tHpsb
yJARaUsSwXe6Lkjl6nFXD6YFcNmNX1ZQkrMMBDQqdAS0Zlg+nTksiXr1k7SAR+/WbkWya3+qCIa5
dGfhAIusgb4kA7PR7CxlF8DoX33jT5pmFXUf2IyW9PckGaFa5uZtS5pkb2fWmhzYiME5zAWCVVqN
fFPjpdKJcQ3/Sf1kf1CiY244AlZoKcQoffDcj7a7/Alw23q5zed0TmbuMV8/tKTEqyaURmUKpmPF
PcwCoBeCb8jyfdbA/UmP74L1tNzRI02CDpWv+fxXvrVcytRC1HXgHOUYqSoj3SIhfEN0xW+MujMk
P3//aT4T4hWkT79EO7nGpL7/grouYOPP2n+RCAm2oc/ZjKblU0L3JX147bLVpf/xIty+hFt1H433
2UC4gMgTDQD2ZsR0ykG/KHnasL0+xnfOaCQPbau+7nNdl1kzKyK3F39SXOcMkffVPKE53BwgAWBJ
mFVZnheIv5GwcuTtZwPyR+siTjHsn6GIVFN6ItQGJtuu2BSuDdn33Ydq2OIYEWSmbwRAG2eUFUQ8
/sgOn8B3VzbS6urBEwGrDAlm7TGy8a2l94xiowrSYmBX/je2R8O+RE6nU901A81blPaORQWnAxYt
VvWvjfVBQoaOQhLJ89lTEJr05BzHCW5s97EiOaOwAdgG973hQPYnBbnNHf/vWtjuxOJjdqj/T7XW
tC5VNJDOVhCBogCszI47B6l6+hl0fXFkvBSuMAI7r/59V17G+xgZK7tvV5os9lCBH2E8d15W+ZBI
lcLXjKWs8JIKQHQHeYCdhbKi5jRFJr73OLoCnIwc4nCt7bZzaywfC+bO32J+DtqUvfy9CAWjSvQR
PjxS8x1Q/+m9hggBQAtGC/V8zpaYIQplbcDzhlQlTnNcrZkDw9NvNNDOm812YkGCIf16kUdqraOT
ScHeIHADyt2HFzmYcPdMCCEMGIsoO+jxZDjkPPkdFZBGl/mZVWhbUdsFGBp5ojSFFdOAzMVMljse
LOzPM0goC1lUV7oZWzqtyx2nzdjgkQwpINBL3BPHJseeKrmdmj3ZumzYQfugAY88qiZv5GoAcmyO
21VnhEwJcnWYbnx4JWr/ncrwDqcrSlUQ98JLOcqQtSVqybxEh6BmhxidcKIAJkq0N729VGZbj2GD
ox46/a1JlA5og99VeSRLVnO55JjKU/dbvvnjoj37E/r3YFAmakHqGQfCzNiObtD3Pgo4rldfaMzH
y4AdiR9mZ1C745pMOcuM9iuDG6n3XUnt0IQXgTCArJktu6MZfhzdRD6d7ELqho+m3DcP2FHLxuW1
QV4upnpZgJdHcNH8Z/Sn2vH73LcnXqkSmUgfeKovZt121AoO7P15Mc4eM6pZZHmMgybVWhsxUrDN
qgrimEUwdnwY2xY/VLb412Jz6F4bRzDDCz3tdi97kXHppyrJljy5soBL3FYKRFNTDTn2mu40D0K/
XFAoxFj3h5k3LqPP3UK5MX5CHl4Upm5ywVKJkJ74UQDqinsqF+UXfjRJnoQ/SpZWl24IshiJQex0
cBlTzHn920C4sA3/6GpHSHLaGPMdlp6puhlxkVW5o3GH/E2tXVOBFt0VAOEu2tU1ntI95lPzk5uB
BnvYd0joAq1nMdzZpkoM8n2bC/Rqsj9SsXwnpLmb/z+DTgD9HER+LrLVGtuXZqjOL7g9PUFthHFB
TiaR8esBJhp+7z9l2QxDKzeQlq3WueD7Bx/6IJrX4pMOfTJ5IbpPqSYzdpE7RORJLYOZFf8HdGKV
14V16oU1mf/2nQwMT1nxjscT1slxaZobr1wJlIZ07KVf1Lj4tNwOR1ud3k+DZKd1Gp7Ke78hf141
6HyxOyannbXq8Eg+E31hWm9dJ4Htag8WjOqCtMgBxk0+N7EKKQBcRDHL80eMUbqcCDfFjt6ITMJz
bfcKQWghW7dm/NV0woN8EDXiepxI9L6gehLBNHjbVSl/pJ8dfhIp2m/Hn0NDSqJ8xvPFGGzPf/KO
eZAJkSQmJlpuE1UvP9OZqJX4j96AkuwIdF7yE1e9MuizgjOfTgyQ/0hxryc5w6PdZehlza9wU3wa
4Dt2D/wp4oLPsJwxpL8Vw4eQ6bqgI0vULNf1SXJeb8kczdnGuG6JmJljwmRmQN8eOnSF1z18yAro
jG/OIN3elAsANoC66THfIWWlXbR2VGeiR1ew9pLpNjXJnoD7jtWc5bAV6V1Jh++TN119KHsvjBRV
/3iAPgI0Is+uXh3wHvFGw9BM3wUOztzuCvS1yWY/MT2/GMFl0JcHiW/tDRIWM9KMRbuY8TGkGE8d
2QL4j9xn6SGLNCD0KqGU6Pwx/eKUl2HZALp13mpLpbxRKUNY4SoLpqr23Tg3KB5yAj7DBAfsKpBX
t/INXC3FjKpHxHEdEtgfSLv3Bsi2+K4mCaxYyt7u7pnxZWoSYYaTMplxUVJcVuErHKvJLimpnc8/
3FyRYJH41aFcr2n7bo1fXHo1Mz1wp5kbv5dSAjMCWe0arnMP/3tmnkDcl1e/1bPHcDQ4aUhuMHmn
coxZZlGwl6qa7+uTcFma0iVN5QXNwmYbO5pC1INxwzrC0kBVTD2zEciq0Ma11fu3uM38KWychK5j
Dptj1sO98iWkTMCjuh2vsSlJ+np0eJPzOaqaBN8qQIR1mpN5oarUg8+KN26l1cZhbHgnAKA3XwQp
iXfqKRu/4vtZnGIpjSIGdnETRzUe6iWdNqZ4LkSDabD2h/p3M4Hm8ZHgjMOIKJp5wL3AqXkrqud6
LIV5E2wxZ83oqnyADQKwQcAmF3SAHiRrlABJG7qNQdbOs360kR6YDRXK3N6EH+4NU5TdqiPSFid6
qY+OquvEZDWfYSNPSGXFQZZiL0ch8sYiJ0GGxL5nU3Av4ILO4sMDTg+p3oLB0gOyDHGLSjNKamZu
SptKkxjsTe3tsRhkRhOI2xwEPVXzKYhRqwgwbiINT8O+6icMy+/OXNMeLthUT05yQewmDR7pPp42
juXp1xv64d4Ubx1wM7/LVLxhxFqCYZ3X6/SeQpEi05kXyVXIFxTQ1L8FetCit1hI6jzIbs3rqEzL
eh6Yew7cXJ1TjDvU/XYnUGlyCTKRiNRsp5TkP7f6Js9IckWGbv6o9h2z67J4zHooPwfjItZ7v1bl
R5Xz0hExWSHzOe7mR07vQ4X43gaI70/i/VQ+Sg4KGA7dVe4RKX6nOz538w5/tQISkzKIw6SCBZoR
PPeIo+X1M4EaQVvYKIXfRsO5WzgDe5LwapNRBroteVzJfQQVkkucfzw0KQ/tTgZ+YWmGxFLlSuja
tmjQWazvR27JNpXKbbY1HkalyjqXp5k3dwl+pGDKVQhjyPdUKrHbDAZpurIQIlta+rFeLI8osg/O
hXYcxROvbDnOipAorRNsrDoo63qBKp1pT/NKtd6GlTaOK2IWvOfJMb4H73Q27Tkm4KAG2sNkP8dY
RsEyt+2Szsbjg/phxwF6+FegdgpGjQNoS+fbYYGioO6CzQUWqhDup2/SzkA15ureScimhYGIRIRL
CU1ItEkjatCUtFP+tbYJBLeAeVV04fguQoFAznZAq8+BdpgWuyNOlnh+FOtCwH0+8oLuM+YouVlQ
GS4nz8tWWsxZgdtB3HIvCucaI8yE5EoqYpmFw6gGMot0zkaRwWg7LwOgvlpzrxJxoJU3EONs6ul4
UqXlPKgUGHUfpEUAu4RaFqwGdwTX2Jx8I3eZXm6Lp3qglNMEKCWkpRWA9xx5R+IcQdiPLUjCN4oN
PqjDi5NvD14yD3J1KFSrNkzmVSE2ahLQyaf3guQsRPcO7fPisYk4e5mCSuL+hvDmI83v4P6gOKvb
Xwp1XWOslEIXi4ZNDXnf3Km0EbauvZU7xi+/yPTpEB4B8Wa+HHbiq/AdG7QQcggpQogWQL/60gD7
IhiIVdpadG3q+znAUIhrjgT2WtMDgN4xwtnpEAr43DT2lhX2qexX58OOxd41twR504OLYn5hhn4B
T2j+1XF6FLcA+uQ5j+mGh68YcG4PAI/bSn3FoQcilxo52mPIFaPtt19VlthTmIC97Be69pql0xhy
hj8XXcBtOUxg5u9NKzEiFX4y+8QGq5jgVEcCyXftRI39Ud4vI6f/m56OOE6DjEl4gFccZz9VviqE
d/UMZGqJHovAmjuGeakOEd0b3GvjR2wZm5z98HjaCxMOt+vKdUSYDapwHWPXKx9K+9vzLsB77Ho6
ZbwX/Az7N3eLmY9X6na9ylASDjkyxPXUxsdI9BUNwrayS5L5Vjv3vNf0u+SsaPq4gy1qbsR6vNqi
vWM/E3L0TjFTDsRJn2JCPkCQB7j9aWayDkcUP5VZlx372KqGnkDvML/3bqea18gQL7uqH2fuLnmB
Iy4wpN7SfdI3tRw8JF9627NmOJ8VEu7XZr9Xp0tnaZEW5y48c+02tjEgnWvR7lZtJG+OIVuGtapW
R6o1+m3YSXl/k1wK4q7JJUmFOVvgs5PgojrknFJPKCaAUPkpIps3DurwkiUz+N+Ukw+FNfuVPG+V
t0cpmm0vRD59WVVWx/H35Fb7cZVMxxK9iZOBqaMXAHLV7018cVi7drXOkbHQIeU6iVgl+Ccvqvih
KMpyfTabbCBLDCcTqpua02RggQEwZw/t1SSYZeN2ZMPJ4khBezsZ2IUsRqzAVW7mZz5ZdJGeXhku
jJaxW6dzA+fDjqgfjb0V/w/2iO9hjaJXTDcxD8cSWsrhWcbDHVo1VM18Gjo2nHeEemur92nXodNr
MWgDWNocQ5hFCVd7sspnW6qEoEQAuMiPwHqPdA3bbgFHy6Aetreokw8WUPKn7BzRFtgWOjbhlmR8
WPqmL6ttCTnU+orfTty3Af/z4Yj+spPp7+kPYUtVN13JSySbbrnt3ocoZEZnCKhVOKWX9Dw4r+b0
KmY0Alm7IZ2Y9cSGwj5ofOk9Anw62hKOZ3YmB7jAqq4w1AdHWQst4rHcT8s8Mz8LzADTHwxYYUTt
MW5zpTGShMJ7OfBtK3qLuwhOCvPvM6xIblesoRVd8+lScE+xVmJ7G453We2CViEnY3k6YZyVC/Au
WZUXdz1bTYbk0G+06J2vvYwFeXS2YKqesq7cdBJv/pf27C7rm3Td1VIs4YD8VW5xa8hBDhP68li8
8v+inNqq5FIbzgqi2pVyOyyy63VxtmZQlgePiVr0uWezRTFcrwyr4TFEy/GaMpCXKV8FOa/pCtRX
9Fpq4w9trIXnDpsOV5uAmhT5e7rD9T2TeVI8/uREVNt5u/BSjCsaJ/+VqED+H+4Us6Dqb1AWHcG3
1h6pDE9EozRD7ZPRqzzCFTMGr0x3S154U8hfkkrw6s8D7EV27GrrVpEVN3XLAeMW3BCi9Q57SeKr
ECY5oQoY5luLyqgor7Kbtk+9hYbUGFJsQWEykJDfTIRboBKEpL4mH02af44I9OscWrML3mgxTX53
hiCJOUvAo9Ku8ekBFbMZ9rlUtm/mr/suqy3kSuSC/El6jLMLNbuy9aLGRolP5RFxKAct8PlP61/9
P9yEO8hjaCQ28MVleLF3fC0dB6oCm2vCpS5FQ8C5E9tAQEXwrGnDer2P579y/XqDsP6XQyYaTt7O
dZxCo9/e71C/U+HZEQftuyw5CDiE+/qV2ZqQM0Qiyy61DKI1ci/eZl8fW/rWaMiUvWw4w57InJt/
PoeEiohzWawNuHmi3TsMvcthIkq0JlmGL0Kon28tUMjkYracSS6rZSol3et2MlsLYQzeZRlgd+5Y
3RO5MyteRzFm5xCRS82miG9kmzw30EYrbD8St113LxoWomvlzPnL9jZZH9qaM0/LiNTJhQ9MXzo1
6HOLFBsxIVZq+b7S8OCxYhC8hlEoyJvNhUByHe/JivqXo7Uf0PglJA4LRsrj5pqeG93BjTHTKiPf
BUL5h0QZFfJaRxpt454OtiV/gZBGoomX1sIdglV1xQDigCH3OYlTJKw66HccVgJvG+3jTAmltU33
DIb5siO0gCh1vJhD449c2pFauS/bblwyfgWEfuDrKwfKk5gUIZJgujcfp5HNtggc+0w2bkBnR2dE
yFPBccYrxkAIca6K283bBMAzASuGP+lWQ3Fw0wK+GIS1lsZdsKn36p5OLS9kwIbnJri+77sDQjAf
O1hCSkhgT9nKNiBm8UOWBCVRGHjgynFYj5McqpRt4LSnFpqfBI2pMyjkSWj7/Qm4V46JsdFCrhyg
dcWZYtnVD+q0vinkZdx3Qg3ORKQUvOyRb5H53dLce47HoZ+YJhYsU8J/ZQAT7icbkji0iFcjWT98
Q7mU8p9xoM2e9lGabSt+Dgjeni/bB7zf1oEK5jrp4Fsgpmb30q2M8MawXTo3ets5DKsworZaw07X
DghlGE4aquViR4UWARawbF3qZaxS3QICEmA9GddxlUnRvS61bLMTz41GClwZ/ICDHzczkvMWdh/q
mK4WEVRGtfvL686ixx5qo2DR8JT7y9Ekbx71DlU3B9nqjfGp5cUo6/bVoee9P+0fFTx9RP77wzJW
9pV4n0scfk43+S50dppRzGbiwO35tOXxVc0i4F2Ab1dAKyU+znPZsJa9G92NS47Y+dHy15gZ6n+B
CYKxocAtKdWdYxkaVeu3j73NCx2nV7R0xFtn1g+S65WHOK6cR+Ej4pAJnHHZEthTpPwcXhPQoeQ+
N9mW2f6hap9DP75bQxJRICJO56uS+D2wKBCXnm/+ZoP6LP2yTSH9YevmycHRBo0IBDVOLUgsBYYX
fnCPMNrBbqbgUXw+jh3Ism1USbNx+aiyIiEcWpTBDjFNmWqIyNgGtHnnQXlQCraYtg1Z4w58Bo66
PPXaOb2Ugjb5pUAwrLja8bMuG4T10qRrC49qXs16MEPcKPhe090yP0Vmj7SzHX+Dns7DlMaMnkOM
7QeuT02Gy+kSFQuAkaRAle+QX8/OCKM4LUfA/Lr8o3qLhA/C4hYHsY7ntJFP2aOwCkSQCpu87IjY
SdbaGNIuh9hNh5UpxecxQXNpf0uqqtyBuyKomiiaCnaeg4RjwNJbvQ66Tb3hEvG/xW2syitDB7Ba
jPLbfsOzj7K0xOqhx9BJ+wpbgowfeWMki803rN2oMhGMAH24rl0rbTE9Wpg9dgVMvKuP1f4/RdWh
43Pj8Djvg1/dFrW8BTxnKFs84HNptSe6lkt4WzqKPT36In1Fo78RYW3aW75oKowDOISVe6UxQF+2
AZEXomqmQsq9qbVrxUXI+4iVukdv9HuBQ8BeH53c9HaH8TTsqZiHVKnEV84K8KaAEBojhsJtYCzT
W55UUjJsNj/ZwNO0g01f92XuqRWDtMJIsi3x+O/KaOxxypG23nDHgmTQFD0eKsozYFvSSAH+FvAn
Q0DJGJEsxBFzs2puhE2zQpNQWYOFRDzbxPBU1JKD5NK6d/PwE0eYD6fvcG9YCLmar6sWgYXS745j
ZmH5GENNBGAu6vWJPG8lP9ex0dTD2GnVWNcyp71Y/HL/e1irulGV9JVyglvK+aQTTMjMFjfTVA+r
rjNN5jb0Ko+1h8jnUcYZ8Pv6MpO3LUb0qqNFlWoYip1mDyQ3iIHh/73qioVa+y3mSaofVgFb0azL
HZqQXXXWviZQ1mIVagG5ezuQjnNFtdgep3RjC+dB4SOJmBlBBylln8uzKD6fSdzwRAhOBrSt8fMP
e8zV9uW+xAu5EXePfTLeyRWDn96Us+UanJ+tZ47L2i83aaF2lnj6Ex4venmTshL9vI1ywWxDRycp
RgJ12XDqGZoq9aGDM72gAe/2j4QKHuUDaBn9/DJWrlKstRNlxCA2DcfXYT4+7dubio84pY80UCnN
ATccFYv3zmQMlxQAz6xCzRHh8y6Qqgipwh9/H4/0LW+y3oZcL9rkLJIqVNgbEhHQF25FmhB8+cRy
36ZYAwli0fNWQ9WBb+8UW/m3Qd1ccakzXen3/6VwcE8FNZRJB9u6ljvqG0MeEr2uhySPEj3GQupG
ROSP9f711CfVNny+V/FfRXnUA0DTXxrPLDDXrCiP0j6CkzKJfhBNe2DXecspLjCNodNMPg9aOHpL
jmMGCKEx19/QzoY+CSCPfZY4ZEgKfr9d+RyYnNynKkIS1bioEz28KGv9Vjhk/VX8kJ0PM1olN2WH
pEQOxsldQxvVaR+1qvP0mc0u5+wGhCWIAVBs/pq6cbuZi9o4rr6a50jRw7RYWcmMmas3Lrfsi+Io
5I6rBCAGzG8M8J6ta3Fv5YttE5QzfYQO9gofUeUQWm2c/GNPRdX0hoC3M9uraEa2qRyHGJaq2zPN
Iy+IO5Auv/eEHNZJuOEBkTZcYVg+dGfbys4AFHaCcf1Syak/3BKmsKDie6J9FY052p6wfAvSERUY
5gfGisWXLYHA31Dpm16l+aCXorNCCe517wfiIMPYarBfouVcYpzcSMlJ7C+cGXUiDknrVj/ljlKF
pr9NV1S+PyNLvDKewWsta9WLeE9wR216QoRmdm9fDpu+iCXHLjwYccAuND4yfMYNaFFSO3LFdsso
9Gwafg36U5HpyAf3OQp0LGTDgagkKgDUZ+Ujnet1VbYCe6Xag1KRj84PJ8fgJVsXI/q5xF17SU5L
nJowiZo5XTqg1yTmNv0KLNFNSfVk8TlQYgo7mkmpEW83o8mSt7dbQE6nZAZzeI5lJxvuX33WFBY8
MvUQHaN/dL3c2Kovo03n+U9VbkB1JOUz6OJZEoyRCYJBNnaGIp6WQ7NYMtSRr2+i1RjaQtGABcuA
rM3zATvEZWmso/6Bh9CDcurQOeCPh8UjWx9aGOliW4hOMq0hrwHTDrWWvTadPI+Rny6aremnJExW
tRswzFVaIEyoqz8Al9knZQCPQT5eAxcUac/Yrh+Gxd8xBt0SCYk+61SI2DNdRnEgn/WCY35GZ7wr
gMUyRNE8Sa4nx88BPSA2rU/6/PF2NWBaO/zfmqiYBw4GQPFFal4nblB7ZeZMrjolEexyEa2zBrCR
shlNAeN5VANlce9ko1RleNVqxDbc00g3TT0F3Gx+x1Jb7kNUlHYchcxHYmqzhskteo3gJMl+XMcz
MdUDsb56joD8hTyXeLBNtsp3GQSckbZzjrgEeVqjP01+LvcdIPqvbcAVphQG9GtzNnCBPjOJwk4p
0Mcq513NU6XvPMTWIhSqwDSoVPrtBQMkO63ndoKCbX4TDlAP8H91+SlNhCt27GJmUn4IJCGRD1sp
/Frr1sesNjUviWI4Eot/YAuYu9nP4GpGG+YJWkfLtrneLAq0PJRVz3lQNgBX/dn3XVwPjdqIVQoZ
EGK4UITjjl3eY3LUxlqFriTp21GCs2rZvck5oXW+ynC34xt8w3UC7RCvz2NCdjhRTTDIWxEzm54M
+comwdh+gZcqL59OeOvKljKXCycicBYFb4SO208ZxPGg8DEnVy5R7RyPH6tCqqv2thdoPTyok78I
cLo/wMvTiuoUR/IzS8gQ021izBEgf+rm4Ve7GqR3zi/40/eIRjd+NESwX0HlNZzL5zzwiYJPmOMg
r62zlu3IvSG1Bl/PZbGVCqmGdyFhAUcNwIAs3c1fQmZcVb3Rl9tjdAwMOyCXnTZmGleQDeLlnh4t
7okXTIt/wp+dbNoW2b1/bvrXZFw7i/VIM4TkrRhnJM76sc6iyGlE3RKfzXn4HfJEc2wq4PAkB3yi
oPtLh2t10RRCtsb6OdKJfBsKuk2hNJjZPwTeqpABUyvv3elkAXl3cc2bPEN+EFkKNXradIoeqJLJ
kUhSdNFVJ0d9NOwzKIgt+Z1rURy+UKkFhr/H6O6WyTxoZJudhEaSwMuXZTluKcmYgME/UwfpwkZA
0+mgbOAqSRICsJ7cVtfV6Gq3+p7chjBlivfFt0Rw6hrGyl8FDGd9LUikGVAVli2jLUVvtQO5GUN9
7/+yqUr4sOo4YlKtSHLpGIKcJwjhI2THKCK2dtJG3wPXThATix+23dfqnCJBBVszQtryT7nvVt3n
JrofCNoRsrZRVeoqbpd0xNqxyUo+qCRcjTiYBOm/FxuaDYt4bOlGGHQJyCvVsbTPcfued8kDQ2fT
w5Yy2vz52Eynzq3YHJSxtOb/PUX/90YklBs3DeTJNt/dNm/SfzWl3O23q+brRl9kNTAo6I/lhqkh
wSoBy8UKZs73zeDds/Hclgi3IR0sIgrYy5ZauB3CspINuPFHEhOQeAGL45hw6wl+6b0+g0h3eE5g
dIX7OAD34qBw5wEBfalusxWOIgB21su1ZzFdKneUnkOYJbZJJysPNaW5qhyrubEt4vBIUH6XcAP7
rRytttzFHiYN4sGT8U63eqYx5UXArm9C6nKLrJO3yvsiVldff1iSgu3jz5WzoddU6mYwthbLGQbk
tWEPDjYAq7gmzSibzsRheCUEE40NhW4ul7kocenxUDIy9A9o1LnJyXsVem1UiEt2Gv5i5uNgEEV3
MSaiVmgArJsIEmP8X/2/P2N8pzCwQoM6u8NII9Q54pFGmxJ0ArBWV+bFkI2MkVeKXQ+rIXjehIz2
aUyx/bgtO2/hcsFyzPewfTbWQBFPct2iau8jfZ2ej7fsQ5AB5fBNssMqoEUAke9Vp1tXSBlByw1L
ObMhHLWzhQR7h4jJxItxKGLphiufLxPSe8GdCzorc/rxzQAd38SVGNVd1TMDlOoBTlhfhGf/s5Fs
M5K8Y8dPsZYQ0NC0PuyPzFaaHDSoYbqovbQcrEp8hzNP4mQyYY3d+EPw57Opo0JyPrGB/Nw8BN9/
AUjEQcV+IpWv+z9/U8KHeFdK9ZDM8FrB54c5mvvvRxyNdVqcrm6xmi4mYYtzcFm2l9vyb8gvjyUp
FJq5/JAMDpz52WXlKTYa8jbaYiRVjc1V/+g40wKG+LN2QtKZiU9KSwZyub41KYoSQ+VpQAtua0ed
ggK03cJZS/OFgRnoTanKHcRcZrjl85+Cp1rFJJkZY/5LD0NTIpEyZ9nz4BgAmifu1R7YAKmbYKSe
OqIbGi3Js2lEL79Naou09OLFqHncwqF66BufaAFo+Dr8UcbnNxDoDB2iBE+5iDDmM9Gy+vX35iHP
Y7s47MaT6SLK1L+cZeMDofdxFIvxBtjv7La5yd/J5a6gDt1hyAhYWPbZ5rgIL+OGLNT/R5ctJEy8
lnHqOZcTIjhLKRNKmkvX2ROFW2N9lxHo24wJZ2U8lt5iY195hyWU3LfUqnBPcuU9P/rk8/Iv8NdS
hRMic02eT4EBj5Dr+o5BXGWwyz54pGa8SnlTZJ5xc5udtoCxTKY52Lnm96jCbJ1fWAYNoLozz5S5
LH1rZ5QvdGGUK1TssxsuLU5U6TrpUtTCfpQEKvzO22xkaLhb9vwdNjHgaUQeVWrPpbToFflNnJVH
2Yw9TytxLrAPflkCo3MOcwfZlo/b+9b4nGJAx5U9xj3v1jVozLmmzm5T2TqnwfV5Us0eHMH6VALD
MVBcgSOOzgNk+j3JY42vEZXTh1MC6Q8B5OFXmycc8mtQ1kRESWUmyG/9bZdVrBC1Y8LRSqlitWaY
1KLWidNWtsHnIkN7PK+i0JSPJCsxDkdIKR7yCqpN9Oqz9INGO5jJHZkjcGsWnUSaS08v0JGPsyl3
k9Pu2QZXo1Xj5sy6rnJDq8LKiac/UavWTIgRaSU0qUBgXWkXKvNGRd1RSjQmjYgcbwDQVuNsak6y
ycN/stviKoNSZQf1QwByGg24uemvtvhNuC+CkP4KmXpJUGdJVzYK9ah59PwmPqk2DkxGHz8WZp5U
Erk9ttnlDUKUZVorplAP4mevmAf5pkKko1ylzAlFrmh19fZGfjk5Rh7WkhIb+c8IQqlcDGzjCYbd
iMdpPhYiI3VLXmMq6CJiPQkHxk5kfaq4Hh3G0qs+xS/5Es9pvN6m69jIyncQ/tMAMKPYm9k7poCI
kE3YX3Q5F7IEl0YOnLHvfl0qQwbYTM9KG7IbS3jEFhIT/KaGP3innshsv8QfsVRjQmI5K9uwOrWo
Ut3oGHBNMA6D62jDl4uprOFzhD0YbBfhnZitJ/OTwNb9W9pMNIJk3AJijk7rclCB0MGsL5cV6unf
HXL09iEW86CHoTm1RYjIAgzwlGNi1zEoGmPqEYTVpCH49rr8uBbAe5HWasxm4M00Nr9b8fVdUc7t
8Lnxiw7PmTn/ntHjIljwiI2SBFmLeVWXQKJDFcXBxnabQrGCbXqaVZazPREVtV8ep8gRcMLAMbMm
9o3pG834iRKdTr4lz+H2QFhr5TAsIx9th833WM2eBMu6aVJKKs/sLkPJeGHg+Jl7AWTNFERLJVvI
9+lKicB3FVgQE6VyOcHPLtR9ruFh3NXvQaYqrrVhHrRveIYBhe6TJUt2dUSkif7PWq/LjHigy7a5
23upN/ntt0vku9PtGbA0wH+TXSWG2Su23N5gVFT+fw55LdcZpG/pLTooQww8SnI5k8SjeRhHdJtO
yRiyGr8rHI+73HDusD+Zh3wK2PS7XH4vMVSdGjAsXtEL5XvDQoxLo0roXhaJhTzgpeWbUltddsBO
6wLwSP9ZHiL78v1vZpPBngQZR7tkEu7ZKBUcMyeiphGAh2vA3ROluAizoobFIjeZ6I3oIzL3FcY3
Wnxz8h/Ns1D0JvIing70jAYKW1aRIFhA8QSECWQUNlEN86B9ZColAVs5xjQ4RCjNrnLlzIiafev9
VrrO8xQIgamGNeDaXIf0O65azYHCLSHKy89m0b0v3TnNt3c+Hjo2zxQoo92mGx4LlFxMQrUpygwy
XrJk1Y3YUqaoj2NzJxscdg93sJMJDCYiwKrGlapBbitXVcJFMtUjqu3u+/EonkcdlPWI5v9yxYOc
ih8x5AvIc3vxQedPjBFajm+nOH+KgTVU1kBzdrZCN+3vsmbehe0SqP+bwg9IMoN3KC+9AQ+OMEwF
yue+aPuZnnw64xqopblLccZdwonrCsW4BUQIp9gT01/oAo8rbWe/9y8YZlfGBhSvodTQjtl0Kkz+
Edx3LOnBclEBlYxRrq6fin2icagRXsESEmnfYwMGh1vHnELgRwU8XutDb0+U5cqmIIXnddtjgzy+
PTeEZsPw5P9UoawLClDWvgdHpY1ciBoAqhMG1LNbhQIcAM4hqJJCwy5D1WXusR98MYu4vWAEZEoG
01FnEEkPMQV7jUKtsQWjXxfqypx1BxM3i7VS4HJpf8YzofmKRAHfrBauZCsTi1duF0qS/8oowfIR
AVeraWRVcBRsUIhhNCZ+9efZTNgNhiA6O3OUUVAah1hKectQpiLCThCnmdPuFH+TFmja/6qKQFCb
+X0fIgvRX3ea+JkyZnjssIFbs+3ml3RcHI5c5Rb87H5gojBiejWhw+DiJTUdjf9K0RyMJY31Zc4A
Kc8gcmptKEcgr+Lg/gDGmLREL85NIEo63r8NEktdQ3ohZ7s0G8FaxfbOl5Iu+9O2lqil0NIwWCQY
KBNG68m7bLJsFzPhhDU2702JIK2hQIsHsywLMSTPYHc/5iNZXTxzYn5qBPyJZRR1TuP3mODJAzi5
jwew+ZhOd4u/3Jm7IZGzAlNlyMPIHgGl4AjZMvO32ClG1r8rGY1wjKmm9ebZgbpd153qfylGKQ47
W8ohi+vjZdWGLL++WySoIc8pKITpoKy8UB80AsSQOx3A2sbbT+WFizlf9Rd8zBD1+VN61M6EQW8b
FMwgNj9cQF7LjmgaEGK6I+FanPzsnIqxzeazdGQDsYZqDL+iA+8dlbcSuE8m2eXVya/srwPLRjNw
RKimO6L/3WxGrae6YTxQfOYzxZWApDsCqMbSameuN5vHaN1KOBv/A0F3OATq9r8VsyCBvURcTCyz
69Gx3x0Z2Jf4uXWEXie5LQHNllGZB+V5J/TGGlgvvTwbnneixtLiPS91GhUtx1scLWPvZ2Cnzvcd
jaRkV72LHL3lzLzpoOxRCnMClSeEPMWLYkXsb8OBFCcj3UoPjVxbhLJxP4MliFj9DvjNZaLyeexh
h308K9a5zpwxDi9wliw6gGNOeJhBXOMSe8i6Xi1FeRBq3yqb/Xx36wowUDGglzvqN4zamSTZXtFW
hUTUhWhVq6xXfXD1HQrOmlhTfD8y+kSencz7SKSbRiBaKm4cskyXZGPwk3b4G71IbWHyross0nER
Se0jXfyO68ZIHuNYNQP7DaBV44wdtKNymugvCrTB959Ts9ePIwbWdDqK5eHlBTav3jZtoPkJriGm
SPQFdcWGmD39VYBWNPSNi+pT3oKPymY6xjbEyNitIpqmDJbkt5V2kwI4AwBqayVNOQWQKxc8JmjR
SjBa2aOVp4R1mGzV+pCfu43Yp/doZR5ZmbcLd6uA64oRql+9kk/D3S9xsqQtzjva/jdnucdDwexG
AdMK/p75YxJFWNkaqVZOoJoCZKr6RfNhZKg0bBhTofww86JFt3M8i/R51TKNj+FTN4sos9hCTN8r
2VX7jLznZ7oJ6TqqTzT5/RGQ/3gGOwe/GbcWRXDpF7PuvElA2MO2k8zAuE4fyOIgD0GlU0T8wgU2
pvlVyQhFsJM3KWQQ25dXAOZozBLwtEBhgLwBFIWH5Hpz2fMEiTMKY4zwctt8F0Z4eIDKoN/222A2
a9NMC7dZrjA4UaFH3jbn/PjJ1+C1DHeaSDaLWz5yADLJ9P0VhiasUTNKYYDvEIwPeztIr5Mhv42w
bYFSssdjSpxA0exHaweaft4xVihlh/UDJz4OGtquIfQbNc0xKC0wNGy2F3a+oi2CJ8ckjskUNKLR
Kw4f2xL0J0YmlhjJjWOukLXP+quSfemgBYfHoMKh3SsWLork+H+L8JK+u9ODFHhzLWsLMb0ntzan
oa+Wy5KNoyC+6c3Nk+O+wZeXZXInmjG0tyauuGz5Dyu89UZLUOtsR91PPZEN6zWg3gDwchs7qrTR
IoBbHI0Cee9NTLh5MhR5P44z8gBxYZWt+Dq24CEi0tScBqBBurJI7OtfMQR5we5t5RXToHPCo0jR
VppCZilBtw1E/3HiwUqMWvQ7M0+q5yb3hQI9Xf5Zw5rFd200fKSlH+yJ0xuxJ7FunCkT+77V9qOG
2DTeHPG8h9nm7065uvmVEitO91yRwqX3lPAkzf9dBZIuRKFVIRArjVopsuY+ccD3haUnbLP2bPji
WX2nGpHnAW+U137hiKODl7WQK5TfdKURGwmP+Dj9F7y+827F7nr0SuEsYXj9jH/ly0sLxbf833X/
Qqu84hZUHe2d7SmiVVX9nbygd7w1fxmLjK9gVYLkt1WDpFqukgkPkJflWgT3o8qTCUcL+0kZfsHA
Bi/iuAbv3NG5SSRlbrUTF/b6JjFK0XUXMGny48TCFcD7W+ylXhzni3CiXB2uAcQ3BK4OTGn/0prK
hpt/QvAs05S4z8p2bMiKegMmtDngj4YWt0LqrhHzJkdcZUOO/XEQqYsbXHBG1Kk6IIs4hI87pdbL
JQlOE2purjqjNrZrLjkMP8e+w8MI0WxFY8/hmzmL3NbUHF6VwYd5PYeQbNvGBq5o9wmx7gcWgkgU
chXh0Mg7ippW0lAAVszzxgBnAs/TUKQnKRW0GwxVPJevELwquP69UPit/idRb4e3YR7O/zkdJecI
oPtqKhP86X1vJ8juTIhwWdGmaxn+TRlQDiZO+8DrLesPR0vIoeJ0+lykDP6OumSu73AjTybe9KLD
1PKdZuWVUGDra+R9HnWWrDxveylhodScAovCJB//whprANP9I9XPqMMosd4zHEcBFUtmWEw5qwQt
wh3k0gs7nT311AoVIJeYNIus309aoRZMe3WzQkqmatfcAiTEcylgWANyGGG59zdvwDwnFYcJzz49
XTeCo3l/4MVuRlseTYzCJgsCvqiAgeZesB5lLet3N0yr3cLHo91R+uCyQ8cOVbaTfnm0NVtSvN0A
64BbhEXyokNcL4MmFD1mOzFI0Eka+M15Bb4GdU1KGX3FzzqbA5N2CDdjebVSh/UQJyZIU6H7TMqx
vH9O/EJXk2zLFvhuNg9NLCb8RV+x2srsW5CcTgOatoUyQ6O0KM+EqKvhkLQL9NcG0Kah+BzMJipC
7z8rdeN/nBquJUNEd2yU9uqeeBxZ7jSYaMrqN82TP4u+LVdkgAR5em9dCBo5N1+AlXqbL2w2mA9K
yORG4C6Fb9RkBP/d05wVuKoHD0/dIxw4/+9uPQ4c6WlyD8sn3JeOj6UkDTtCWWDuhoZ6xrf4cwuD
q5lOUtetvZnmEexZb9sFhLSnk5woYTcqQoR5uRsBIZaTxkEJko7Bl4/rFRfC7uqeQedrnpb86tEr
UiOUd3UECc4+dg8UkTki1w+W6FnYIbvt3BU/799C0OW/XicvjS8NZ/8JIFTCH8ImIuc1C7mIrh4u
Y4wrL34dtKt4fRf87Vr0aIikvpIDcsWLiKghokO31snP4peKMtaF124Zm0j+o0GsxpozcY84RBux
2wr0Ohm6N96i7yReFNu7wtjACX1+gmFkh4P0OlczMX7I21GeCetjD+T6acDBbLLSFVrNzPC7N3sk
UZ4rnnNnIahoKXaUqHyIE9//dL4hfygIm9f4opBhHoUJS4MhhElACon85GKjqAt7zBlV31PdlPAl
Ss2f3Ayx9GTH3TYDuFYBBGdPCX8p7bEpC+CqSg4+h30afvTHrhav90QqscVGijtXsB3SKys9qfwy
dA1nFGgSFEVJvC6dZcoYStNDwPrYp0F/TWWtLEJ63e31xtPS7Ri8DcWi6D/XZbB3mTjzcSzzsz19
Mnv2Xb/RwCMwOk8tnrQk7Kt+lDM2Etex3kYMqLI2jNmxQgSgFYLKTqO3FW16zHuG8t8xXsQNP0L0
YOAooh/RhUvWRsubmVDhuZ9OGXWv+lfz2KdbT5ro2W30GfBrugh2s07WaQMjOfsNxrLLEbWjc2vn
bW4z7lxUF9V8yGPoHiB5KNDuT2Mno3UlRAWRZ/xCLnOFl0DxjQKpqtxP24i4TL2rd0BKPiFfyhfl
mnTjXx5J/XfzrKQei/xOT4OV/1/xwpIJstE1ULIVPi4C9jrUMCtx+3/9Y1a7ZixZ/aOxhWga63Sf
j+47+wJgQ05HGLhfwWktf0JTQn0f+xjwyyNfarXzfyAaGSYH/l5kmmMzwFDc2VnKk5icTBmUbk2B
QHAEWXhJFow2+Qs8HuYjKRsWI3FBENa27Np+1GZX43pbiSDsbuADODmonnz5FPF6Xs3afvbXdFdW
NG+sEFn3mN1U3D4bC19MRLYvsMxyl/6dR2+sjDJ/UOBrZyerye2Z6HKm/0lP5eIzPWiCLvQe5+Ie
wuJWKWCMTqJOrpU5Jlv1hghp9aoJNgaC7R0n47kJtlbmZOgV/sINgxs2K6dwZnLpkGU09sr0B16P
ZKktJMz1QJ1yKZYe3Y6W8CKG8KQMlYDODwyO/SfEeLFEGX9igOo6cX/1kEPmUqLfr4vzLiY0CI5f
9rnIf6iMwQDftaTvPV6bflekJs2w+qhHBAItC3bZykzj9mUBP06MXLg32on1dND7WP2a6Lk4MvVd
IFwlnHB5hAUrjyuOCnjsq00CIACwWBIIV2748NXjVJwj41DXwK+WT2gW3zw/lwv/Vqj89LrLbQsp
iT7Pv6KTWipL9F/lsJXFVyCBOQuPM4ZQ5kExSzEfWxB+dUNtD/jk5HPKPZB3rdDB7PFcRgychOZ8
IeHnrHh8OyWuZR0DiIGEk+UujYLuSkSpcXYOVOi+oaXHLi+NV6lG81yuECMlNAkk4DTk789sN2Jx
ZguITg8ivhiAPRXuc0MBymQQf6WwHk0zC6e/KPRNAriTYgFdQXmYmmE/q3/BZVjRtKBz7F2ccF95
oXwD1kAqN5hzsJJFpV6e0BGxl35h7ZoPwFzoeO4vh+nvqUbE4i89iY7xc8rqa3phdMd9xT56+QkL
MwUMR/iXwMaoSW2TB8zFQ4zpZB+ZnHUKSqo6Z5+Eg/t9Zt4rOcwTOiUorjjGXVofhYcY/S0YNWhI
hTMnBvDzhwGL6E9jW4fmegrINA0rIaI6mDEJDEN5swg9aY3Fdtzn//alXNIS9nBsuMerzJNvLZ4q
smRiEa5okgRpTuAo6Wf8KkbwMXT4/+uisIj1kUXb+Wf0Wliy5RanGjG9G21KsYy8h3v2na1bWFSS
LfX4JJbR7zBKV7ieI1QR0zTS26NUfaxiABPg1g+auyvY26mdFTI7GfbfPl1KTeXhX4Y+YkwZ5d1P
lxpP4LBsoGPyxkZ82JpPbQa4q5ajm+YbkrjIvcQyha/7HLQN6uc2IacOW19gKN7mIWPeRjFqO+Tj
cALBqjjkkKfFARqQEeHuTtYFvs0JCxI7SbXUpiJo/PKu0EvgMt/NUUsaP38tE2uasNN3CykZa2F6
HkenYjJd4lYxys84t5PPZAYJByicwM/QJUgROZuwEDNUClHJpasNUu4D/dmWN8LCjo+CnNvB8Q16
G79GukMRHzFkihID6RyBtEDzIRFWwEkptlX59ZKNhuRP6zjzKhpHuUq9hLnma6GoHK26zcCMi/r0
BbbL+u5Bs979tJWamK9X+CKWFNaI4zOVTKzL4Ad5u4Q2VmQjA93XAD7MWtQskoCRkzYCKBSA67k4
lmPB9LwyNu3mNDJTA72wMDhrBlryZp2yz3fFeuYRia2/L715bMKfz7tYNjWsTedEVCxV7GDBqyv8
WrKRMZi9klYqeTY5FsRCqhNbIx4VC9c39NdHGUFtTZ9NngyADhOlCZf2vZGQaVgTLukLJiYUFVdq
EZ1OyQ1/eKqwxNmT6D2906TxqOwh/tAHd2+ncqx7QmCNeTFU7g7+aeg2bt4OsZc0aef4OR0VcFfr
Zvmjd5MDHMJ5Nlvu2x1VDiC3biJ3LsIIpdIjqNsbPQ+a8ToI1V/DZw0faBEIIGiJ7uxHEIf5lggP
x2e21iLWmGMJdMwjLG98oZvmUR85nW+8u2HUh1mHFtSnp5sSltENrKPHGQukBlBv08A+votprrnb
FkeXZHYikNWMnmoNcaW3AONwjjuteRAs/U0g3XE1H3wZGuI0fVAMlr52N3/dV9wJCVUpJXJNNpY5
X+9cSZVME5xYCAWwq3qY2AvUAy+vtbC8iwtor23PwRtdEBZFlgM0kN9OJjNaFvT0iGYnaDHuDh6U
GWv7TvfNv0xqNPiXWYtSChYVsKcRqpI/mNeDDJjox8wZJ00r0VGq3bykSHDOomyrqQaubaQXBYww
UAYkvIuzrNIhdbPSnGFsV0UsMQbVeJLaWkWuO8G5u7j0wFB1DTKHVk7Ew4uGkiGoZND/X22uMNG0
ui8gdaamuEUrsgMObXtBt5VSKeG5P+I5lG8DHoNWO2AQ1gYv82gFrTR/2jsjSbvxWShKRpuLJ4Hg
BWryRtYJFIp1Gnzy02oijJOAdXNLsvEF+YamFJ+/vxzJklKZr+I1Lge3NZ7N1LYAccknNuw9kjTX
Hv6CHtTm22c2pGAIm2EaGyeETeS4gPij+FzHcRUtimHT8VH9mtB8zxpWRvBSFMH2gBZUK5JZe4YL
IzDu9wHalDaTmRVtbcpDBocjbPneJtDrX7Zl8EFDGJuRvKUdIHlp8PIE2GmmF2q+zbyPMWMpKAKI
X81H7HHihnLhsGuN/BQ0dE8s6AC2qzKwq7lO7tt+EOzjYN5jJyQIE5duXZJTFstCsZRLiE/SjHNu
/1lSPZvOUp5USEleyROXUgybBb7uFW9aaAnUUWrFsyGaG4rrifH41NnCl+Lq69oKosq1jaoGOsG5
4pDgiGwVbt8XhxtRlIF2L3mREWSaQ9D0yC1Z/wmSTDe5dYrjYIL+fYD/ze8hVNmq1uTGayQFm51d
O3JTVAUcyHW5nPjlc3j+TjyUZPcIpC07gJ7ZpFzEACEmd61lhx7k4zUv4QVIsHAKpXeHJ9INqFwD
lVim3RBEMDDF8QDi61sJo6zFRs7Fuzege17MmB6k0uETrm+poUcqz+ky8zUHeKWb5mWQLJkNn6zx
Hd1SdzF8OqFfq5HtqlCAf2DX3o/nONd87MwWDsZ6++0zK72WGIVbgZjMM6CUlhGFimyD5xh4qRoC
xZ6/2cwKtk94yMyyLihrmCvlMhwVNc4BpdXHfT4pKxVvSTDP11YMwna0evp/eKJ1XTx1iV3BUwTz
VbuYS0crMtf3FNBSrG3fy6g86X97337sh5+uE5vbFXBPeMtd1R5nGfQPc9c0Y13vmTrfDCupea04
MXNQS7WznIbH6JgqPF1OrjpSnmGWr1WOlPEb/DmiLyAI78RooWP8eWxTe/2zstSWopnH85gjxu4/
t2QZVpNMyMRYKb1BdLxOhaksXVr00vB3mwWjflRSYuKJuuh03wa6A/Umbq2xznfPWSl34U2hSx53
H3TgtkU5nmI+Z7J+9PIfOep0tw2F634gEjTLdG1Zf07Vz9nFe/owmh97+FxszUZPS1rEk7YXflrD
blZn1Cwpjx3zIoUp8YBvopLCB/Lvy+tjHFVqS0wz/f0BcPwV1E0ChVWlBVzVH9TiGGwxnTkIdaaH
FZSyKnK4sNC3uz1HsbDNYovH0KtjPMFUM/sP31BnvVs6wCS/Wybtf2ngjjYZXvSFk1MnH/KqzEzp
luSU5ALLXea5GX7TFcrppBTD2O5SFMG29c4ZLi0tLh9Hu4yrbFxZF1s2aytwURvTFkm4QiSLof7C
JJQm8GYnEmTEeEoI3B8Qnsr2S59oWWSrbG1nSBbYrWWYoOakO4NEQkzA1Cu0pfwAK7q8xDZGmeAA
X0pGtKME2ysfurXKy1jUYjYQvarbBm3f/oMQrKkH7+zY9CHJPxRhZyU+SDpPc6g80OtIo6fnLy7h
52EVs+qpd3dAMe58pWeE+dScQaBc8Vf6w6dP5ylvCGvoweWgngTxoAKSIUcOMSuCdNwXJ+CCOxGF
Jg9ycfXczI6i1x7NP582R+jGmhI+XVjSfZfHi57DVe42+x/v7j2GV7qB0QhwU5OXgGg2y2REVnZ7
RFAyAi5N/Oglftt1xsWg/6MaVwAqVgIDOOa9wkoVfrBXpoyvrHDryo5wxWVK75HmW5X3iTyS5ozP
sMWeD58lYv/gkbih/0Ggh828xqM06rW677Z9p8X7lpE6D0xTK8h6dl51kQi/Kf6Fdxgc+9ZfO3bW
/m1TnkxiBKhIND4vQiYLeM0xgEoq+1RBX6mEMvEsl7L1hpWVd28gzj2UwU6qixFZDrUkLFcp/56T
hFGR+QLf5JBUrNtZrzUMUOqJ7YW2sdfXYjo+923HJ3wF4EGvton1tPoMBL8wbZziJgcHBZK+BYqp
3V4WmN9Jt+2xJ2MFot3XF2JCN1GhwIM7BGR0Jx8V5IaYmRXCoAHP60on+k9EUqT5gywnn3/HOWz0
OqtPGUJOs/yxSwQ5qbldWwMHmXupG0jBJ7jttonXRy1zTB+FA51LwfMdDg0GWDPpnTswmHZPTfN/
oYM/IWg6DfIR9Vce+NQfY7g0Zjbit0t6vG4XR1SN7TVyOS7+dEz4+LKqSMWtS6mpScotH1G8eQyB
iaftydSVw3dS34Ki5oC70d9iEs4t+MgSUDpDCTNdydHxdWY+0HUNAxSpIKUY0w/H80MUxi3U/bnc
n+80Wf+LtPGy0YD7T6IHWQE71NzqbO26/7H5e8A9heBe3thTnZtOe1PO93LcmgG0nS1NiV3YpgIB
Lem/52syVgJYbO8fxg/GwdckevnzIrg+lWjfKg6aK45RnlMlWRDjWBD0UtVAwYYIJdCSOM6JSG/L
e1QpJQQfigR0jJ1BFNv16AiUDLIB2RgtS8UjDd9HzFIfcGg4Z+ElVqfGeOMwNCv66uiatN+1yMJj
F52Pek7QpizWrwQ6DB00VifukZWpNJ1LEFQY61qLYT1a4+x4KnIuFuUqggvspmqsadkvoQijRWbQ
BQqS6DKM8eA6bjX9Vo6IhrdMLqBypcJ+aVJorEQ8JXq0GA/j5O9yq749Nz72t7YynY0wHyADwouJ
GK6i6cim8CRdcfac61aEdUIWcIpsuu1XTA1DALOrg8ogFeDx0jt+IxN3CJzwIbp9vPdyBNCEjtvb
JeRurkvsEmcvYHi6RlH4lPFRpDgxNRQM3bgmRV2IbfBR7GF7lJddz2WukXWj0lsdgD5b9a5vFCXO
wDXEltvCKyZVD32/duXRYrm6UfqYyWUWweEBnTKUVcfJKv/OVLDlRzf/5up45gtcYJr/ib+qk9of
3nJ3EZoUx8/t4/88YG/+wGisV6k6QMgNpapauHI8gzR2yBWJZ/AlIYT/ulHnIpxPxmqOLPrraJo1
oUwf6rCpqey8mue1UKwwMWOlkdO7SclZ5xkea6mNoHdR7unIqtXNIzwnM+MNUgkodGKRqXAw3oM2
KX89JD4F9Kwn7aP2CEptPut3xBWBLH2luZqee3zyZJRuIgX04f5PdVMDWbuxvFFWDkxWuMXzZg12
NZ5XJAgXXpXca1o83JAFeCf37P6bmfDQjVqTd/hbl5vW4D/HRrxey5r2iy2a+taLRCt4fKAzt15F
xDeI2ZBB6NCTXxU4gxp8W1k0MBDifmE7w6SAghboVDZ8mAtzYeV20g0IHDwa2Zg2Cy9I0waTb4NI
cqIMMQHUkNEg9Q+2Fa8ARuxdPK9Ya7CRBzvvVzzOUmNEwVe7fQJUhpiTqMYvrvs+DV/5oUIeOUFF
QD8bBLkQOxJ0inRa4pTpUYp69Py25VBl80qKkNbSTXtP/XVJUBnOK2Yx21wcFz778oltoCn69RX1
w/01IlCg5zbX5snxvGopt86h5XH2bQ/xKRRe52ELes9vIaTqsBAJR9cR8K35H2Kwyhv8eQLHiC5J
Yh5wfGC06mr2EdaRic0LX+H8y58xc5mmiS+igHgUZSfpt86gVTs8EXVaz8NQDJ9tQQLV6OPXvIs+
Q3vuJ27mu/bnVKo63wTgx62ZNFAghhCCpctvnNl/WC/VnkfOa4yGzx8lmc1nhZVWCzA5j1B937Bu
qXdtbNfrnlVursxUx3h4eir2SLQfPTfKLl78JZKUAcQuw2dqiTAyhhZ9MINQNTHidzS4zgC8Xfan
YwgyDnRsyZKJGsnZ2rolnTn0QET3h6DZBMcP2AiB3s8WPietmRNwOPIKfID4m+ooznEkTHFM6+5u
tXprsBSwX2/W+IzubFDhEM0w/4LHEJXznXK7QwVLRdWTBuXg+2nqsrnevcb7g6MsHkTV4kgi6I/7
5i33M59gwpDFalQKhcurwACSGv94IqrOnHsjpoedz5kOPtUd79oTlLG+kHKYi4qkW6ZbIFlfCZ42
sT+jaU7u5QR1CFfGihRaXn/H4qXFwwtk9LWlRlDzo5H3AeBwzKwzOEebFqYWmgB+SBJmtNZh+a2o
Hefy8g7AsC+FgvwrGnz64QJjZe1ORe/Ktm3Mio8zHf+ezN8TUoJC76UUWTiHH1ZvbopQbVjo+O8V
vH48Ok06V1LolE7ofO5T4aDZBJ89v7OdsDRFEd76VVqUI//tF++pUR71UjsuQSv0xUHYh065eujd
mMiOW1hGI/H1PDF8T2EH4iJ3pnXbGtPv53R8zBrmZyRS0FLbF0F5il8gRNNPY90VMvVHlRapUJpu
KugupuYbffTgZ0Ok+g2HrLQmigd/SRtl4wF8hIjq44lGawhXURYDSYPopj8/h2KMyk1c86EcHXLD
KtkRg6+jwy1hvvsK/83u9S0c74Qfl/YOYurmKh0oIHKekKcT93FixKP0kDe6pQAKZJj0SIIcsanL
VmWsk3Dg85KKvHKwZ75gCQFoA7XJb6q4cu6snmFk+zq1MArAVLkodW/yGG6UkQ0URJ+KVDsRqyFo
+RDAA6gnIaNVNHgRFu8j5dz8B9DYXaJzIPQ8uCHiIrbkAI5Y6bnl5iBi4SzP6OB26A/PZRWUfeTb
7Egshwn7taUygWgLvADYoUrwR+yFcDu5ymMlKI4lwZic+wXOv42R1MaCQ57Lg9graNI6HVw7eXDx
kFOjC9VsJIKeFCqHfU/6ffPhhpz5MVj7LDdPsxcRs1OrH3xrKwlIEFQFihGlr0Pm99UwPQH/KNuA
SldBuxaOTwjjTaOoTLmldRzqhM1KqV+cvd+3kjTsS3no8eWDzqBN0vdHRO4JQuf1+ksEFAO5BbdE
ITVquWj4oOV3jrk/mjYzvNC0Iaayc3KzFugubUf5Vci/KuCM4yE3DJfFm9s5F3NaLRjlRRe492xB
VDRARYHUpG1D5/i+hgxl+Y7fPa5U6kc+/0+GZv68IB2W0nEVnetzNLZJaPHap9KF6Nh/mqeMvZrH
G2kJaz/srzYH/Q2DgduJd3tHoF2f8X5byxzk+0NZQiAwXcPLcphcySQcepFXA/FzKdkKnYsi0mc0
n9jHUQbt7uqOyg1VNoQsr60vL9G7xXRIs8u9ciRax3ygv0jjcYEizh1ysL7eNyo+kNuA3ZVuDb1p
fR8P7RWf7jnyuctmny0biqME9e82lPN4K0tFGOaYF3VJ63aB6Wm/d2NF4b97jxW+hFnoBnNGcnOC
NbAz6/9BVV9qArdCFMbhfacnQVyml9QOCyLMRjwwiVtMuMgykZ9he+3Yh8ZuJg3Q0gtMvE7A/jGb
/nsTunpKlz61IUYHtjk1M4doY2SALzz/LrjOzSSkwv4NkkxrPjNKRi+DRKiaRb26uO/ZC+/j3Px8
VJMkxGcWF5J4lGhmIrtDArhROLg7zMOgriZfbJJq8SerdfwEWPGoC962kJmZ3xWbNB6cupIZTGVE
E4c8bz6XmIpuJNO1FTYjSRrCrr1pbqJ/IXO1yu1OyF5NGQKii57B+oTtobtMZ4Ai+DxDrN/67VsR
Ze7yATw6idOzZW3ElyIPLsEjvwrz7K9kEoI61MR2xwcsa2mRftx5oWeVPRU5ibfxcdfs8ooA8yYT
0O/AEevwBsO12kSo2DaPpMcuuczruVUyxivNyM+ZBKugJKVjLLXhiYI8VbiRMQVCpYqLaf0+e3tf
bWbrqUiCx7htfGs4YUsQ7/aFV73gADnYcSVF1GEz1OhmIt7Rg3M99Q8MUC4TxgAUliYarARoK8Yq
ED9N8/ivmjNu9sZNtLTT666OF1YkeqUNwcygWVPiAx3zoRKBRCRr6FnvZs+kKhuIsWbzKs++cZjz
dMwEAO0sVXjJ11UMiplYXnO5xee5Fb4fHXaTU2IxQpr9u874bS+KAiZw/8e+jHNRWWbkYSh2LWuu
J2dnhP4uLfrZ1VBf0B3GU/4KGnd7MiYm/jm3iI9dpFcCWBktcjcFMcMy/sTgsK0rzveMctOmTbyn
ZDn4b8GknT2/MWlKmOwqNvoGf4R2SlKjXTTjSrdVwIQHWjIYYZZ9Z1pgWZQVv62MkXr4nQxZuCI2
Nph79Uy2JjbCN4f/TrtiRY8keKShNvT97cs19dmk3wEPW52qBZ9qldsl6xBwvbHv56eZgyQRT9Md
rSu4CJFLUGR0iEnZH9F3CW+sLDoaEbclRgmNRyvTO2RiY6CFkrKpj/zJUpLaxdymBewRSONEfszK
8T77lc1Pr22Xs60Zqcv3t94vbhpfx/JhjzSOkpmUcBC+U4BS2wkgHKpyZVPi5t8JEMdvzJ02SVVZ
V7vljInE5Ucm4aM+32CILpmR73SAUXJbWmauxRpj/qCvtUadSmFXytJnXQs3RD0vBg6ordmeKXvu
mBPKHW2TQ6ZF4JWe/ZIeKxy6+ClXhvK4NJ9f6gLhLUmBGGcAgGkikbBY6qZ5MxQlnhIKP2Rd2skP
8i27Nk+ZWHNMVmWbaimOivkgRaxq1J+P3rCyehao4buXfYPUNfQ8FKc4sYXpZjgE6H1U8pDJlxnO
98xrHfWTkDl/gsBSZ5foqxzlFXVV+Kc72oXULefU1gLvbMkIWuBm8EoctzedHMHQMvv6j1ciQxIG
N211UVoP06nAn5/BJd10RLUV+JDGWDqbhii/Mc9gI11xpwXyNAoMbVkDBB24+F+js01UImWpQRQ7
I5yf64yZqEVhnc5tRivAoC3AFBfQLFxIoAteJ7JNTNBTF8kMj3Qh2GwUVt9ow8mXOznlfrJ2grlo
Y7oOjQ5LC/XGonz+T222krtDIbXigqSXu2BgUY7m5G/LxE1eLg+CpfG1cmH9uPsvzhp6GKdU/6ug
Xv+jri+e+X0aisgcr8o74BrvS4ypCSIFez0g1GvQF8WsUc8GULDPhbBvbSqcZNBpaZmlRzlk8V25
+iiJJAfaLhUVHTnQc33LXFDOvyplb5aZMgOVquulnTqhMdEiS8KuNbSyJHIitSeExCSwHCP65hiQ
IFk7IdVst8Z5ci4iiDguDZuTP8fbNH+KuNoG9grfhmLRxLRjmBZ3l11ChO/p4s8COo7/14rI/JNA
se5gSaYd/6KNn3T4fnJmt0qs1Jfs+4GHEP3dgI0L2MNV8IKxW12e78xIBwgnm63bLe+enjb6rp2X
zcJq+m5MjqeYcRIVjQfYTge2oZ8uxKT74J5irX2PM+kW7UjGsoQSO5B+CH20PIUJvtVVvnAiIgKi
st5ihRzQFTfusvRouMfL3QJGMTQD3WbKNuN8TiwpVSwoOCZzwJ/1oi3oLH2GMKYs5aFzAvtTp3Eo
K5K966r2D/N5hnjsFvoguoGsQ2EYHeby9/l3eXNGsBJohEkR2TwzlLqut/X2XvhXN/aBb2pnglk9
OZwA+Kz+6d2T2uxp0P00q+qxTjrUwh8y40PNut/yp+F2CrOjfydK7lex1G9lygTwcbfW2dh7LlRG
6qlHxc1/3KP0ultEUZcrI5T5SYATgNNzf5+OQdcJ4e6ziwlLNyYaPEqBz5vT4BdwJvMlJX9mPtLg
uCPVyE9bwiLxqcrVQUgHxg5Rmo6TQe6/7FjIAxY0eBSAnasic5Le3vBAKwKH7eCeP/j8XBL4qKVF
vhol2EJVW3e7KPbmoLTFBvlxTQ2799vHEyl+yZ/ihEIS/noHQJLtSbKMtK/K9lVaxktNRGcn8kBH
eY4k6WdoZOQ4Ntj1M5jivdvNdmRGYGfQVGZoggC25MS8CkuvqcflcFhWhe5dABKX7dQ13kkAVlhk
koaQM3/T06NANPEAmf/PYneJBvPSonZ2t16iUAgj0sG+MM+Ky4aG6ZfkCX2Cy47Y0/nXeDosEr0A
SZLzYxLIOJIoERiAhBDonpWwuXFJF8QBo+lOr3J/OjW6VO8nykFs8xGF7ejWA4wuqFZ9Yb5a111H
WurkKc2tbV+kg+0W9qLPavplwSsrlrCUMr7X+gvjVqTSbnu5scDLBRmNvGxKm5TWWtm4p0Oe/Kly
5urIkjKajfDhR6HE5rEcgGzVOCL8/2P62AQFbkAazpDlyr6laX9pCH77SLq7JwJjyW2QP6E/ruVs
9o6xvG/6nDE842d5wpXmUlhAG00TJsiGVDv3ePJZ5LNCXG0479qesq/ZeDMFxe2GJVksGfg0oUl7
0rhaakYYn/eLLWB/vtXpw0rtRnjXmjvqJ2eYIJv2gl4tTAzMnlS9DCQ/ydkwGAnkNB4iyyyokrk5
QSdnVohf1OX/o5bhjkpauAh3+eTMTbb9IFBPBFI5u2ox7+BFmS6ZMVeZlyFbtPw/rzkaHiW1cKWq
HP1gxBpyqv2SuCoCZyXXSIIsLqW5+lI+HKk+cVJ6gvdFZEsXPMz9wBQ6pbFxs9+u+4bn2syIctNk
2xBjhD5Cl1aROsI29lFdRm8ElSuzZVTtuQTJd3uBSxX0+J25hknkMWm2veyduSRNK2TV9EZKs8k6
gMRqE8+mBXx+nvTm0WPeMz4GPhgm7QJLAV6k0jn6ptBS+dWtD8ZyRWGEmIXMVK/5lOGlg7+XQ69O
1u14am6K1/UhGH7zaLWNJOc7C7C+Sg6Nu/nPQ6EwqYSHfaK0rTL34fDp9DOrWJ8bxilMECbZ4gyO
RD0kRdc6inL8SSeYZFQ8h05OHy6OI76pfJoXl428cc2ueAv4842JBdwthRf1S1rf5csMIAlYF0Tl
mMiRGxIQgg5xG8xWVYJp899m3CIWdW3CK+nWw2ZSzK8fGhsQ3ZClZIG+MyVPoBOo0T8myledQqxf
LExOSUFAkCyiZ9zEvjtYpQojc0N1GoDTU+mZpSTP87NgOTgScy0KnOGm48Iyiiex0Rzq67wIpKqE
HKfb7deq09h3dCZKJmFCM5SQJNLKABrc94IW+VVoctaiFqQ3hslKSiQ7E881I1mYxa0rw/BR9r6O
dnB4w1COEReFN6+T4CnK2Yklz1p2gM/T2kr3l4XqgLLUtCMXaRdDGaKTuQm/LljaKnOezUTBQhra
l/gfS0aXFM/o2WdeGWwdnQKtVCaxj9vd6dv/CYM1X3Ilnv47mYPe6oaAdhJK/dgMQ/de4Oiidp5t
ZkDHt81jnKnrUhj0B5PedkoAo1VSZO54pBbKnHjSh3k9RQqf63ceNrSem6QHrKMZOnX7BCJdtidP
Qq3egLBwtrCVQpEpmzaYkcQKhU/bIyIylkqVo+1RH9z6d38gE26chOoH8/YAgurXqPHCJp/Ae1ea
EU9VSxrlAQBtJeitx8Uf6vW4Hlk7c06Ih75eC+2u6X+QmqEliydOXkw8HysgpOxpC97JJg8/qwrz
2+t2RbkoqvLPgBLrjmT0Fxc8v8YtLYSbuFdokFnn9jsox9apK4ERHZ4jDR3hgc/fy/U2nzS5kALZ
obgCpsrPE4dnZaSdjkbdXayre/IqxQl9KnN6GpmbG5C2kNol0hWzzYic2bUW2g0ANmZvhrnLdFrI
+JRFaFkjSTEI0LQ1/H6STEwecU7vBipZoxeUbc3NxnON0K2cWLxejkbcDelooWk5/rut7aC0mayu
e/5HYflBf2rSkkRUfxv+YjM/eq9Jpi2oLn7DJ4gEKYmX+aP5QIMSK+mABR8YP2gotzoQkYiRWz/T
fkDVF8WGJ1tn6enu+LZ7uHkDKsejnK8OiSXr9lbTT9rHpndhq4/tg4pPPuAp7Q//TTC3dTgPLtkN
hy43qPt+0dHH980KBi3V47+Zw70qsbtIZQx5GXPWdZHiY0X1UWJ19wihhFSpdoAx77bmmP68o/e5
kxbgdVLWCP6PyY8Use/6JLREKn4mZuIA95ZaFPta4F/BfTxYs1zJhHVFpFzXx4fWQbU9RgjfJHns
Fq/JBprIoHp4Kn1Qqjo2BzUuE3jipaMYypOuHrlTmr/PhgtpMDqRUod18z8F+7USqmYR+pFmS3Rl
SbDkv9szBY/ZqMh55X4OUpl8Ix9HqikzL1HEIHtg/ktriLz8RRvIj7Iu2bAKOUEVMs/fbcGYyvmU
+Ul3tEspOt8Nz8J412psuUeY5zrn9dpuHK5zEjzar8qX1xydXjU6eh+I3UT4vPdSM8Agm8teVptP
wx9wuizzbxmUI2w2+8+P7Q+YjRT+zgFkjlyONvEZHCloXuDWtiBXtBTpzwDtwmCgZmKt00Q3w/q8
gYwhTvf1zZE1kpoa34kpWdf9719qEJtZ/pnG9jWAPUN44IxmWWjbli1zhsiLirujrqSv7+NmwPaH
85SLFOa3c8R1p6C2QvQXdmHFlB7paLzEw2u3aMHCmez3hqiqYuyCkzOc8ggGUd0EDBD+fF5k5Tiv
ATI+hmR25veg22LK9gMcgBBn+iR2t2/pUy/OrdrA1BNf99r2LD4fHR/vEA1zc6IGEPx/mk+9l4Yc
PX21sik5hb9iyouZHfzCzlwCPQuv6b6WozdxozBRVYpgWNIk7Nni31yMI7enH/8xNijTJERi33a/
MqqQwmBaOAcOnPRbBJfBBhXAfvReLaXljhOgZTQoLMPWwe0ak/dNzR3i70+YpRhJ+GW5+baGE2EO
IZcrLi+rv/lznHhOZBtfuBnWfcKhHOdIxqt3ltk60rrkhF1w7KDNu0V1VtW4Ld+gG1b6OX1EKNLP
eIderZ+MbS2gpB+KPPzipCGDL4g+bCCz2TAEt17IjLlcS0MAiKbx4EmmKF72/OiCAE9paJkQRmWN
Kpg+tbOAB916KXSNY0f4hH/0fK1ju1CBpJZlinHNjohZMZQQxL5rcBFfYxgkNWTd9ok4x8CTfq+C
hprdfQfjvpmRQMPZ/8up80a/oH76k90HUTMiuT8gwHz1icuYggPIKH2qlrA25sv1qBj1pJdeVJ4I
dBqAR4r7UNMxv0/9xltz5xvqvljBpc8bNJUahJt635PJRZ1ZOaaGSQwFpgOFruzFWAvHbJg6LVjV
pspNrjWrucK5UJBgg2JtfR/lWhHaryLk52y7IA6DJp8Kadjevrvv9JcKwQj3F7VeNfWtlAdj22Y4
uFR0mBlst/XoFn0JJQ26fFX66QkNa7PcIbUGuF+cP4s5GSGUtvMtHslmytV/YInifVtXMzJ4gwU2
sAD8sKbSCKLCGdXcZex2gZy3dDaT3LGaLTCK7b8SQ75xQiZEfniGEyv61vqcVuVomPVW+vURSakI
FNujv6gJBJ0NhoOnLkv5I6oxrPheFIjaCJ+ZbIzJo2LmnR63ZIX6F+TIktP2JKdhH76ZDKM1hwo1
Ech38gKWD+dHsg8APPuZhFslce8UrneVHsAIkt0JQK6eNkHdO8Ms7fj5ULjShZPuiTEy/5QI/Da3
56jkhPMSOBjvCMgtxgFH+Rp5GzmchGJKtAY6ub/3VHKM86SjQjvh5FUUbMr3U8oJZr+vb7HzDZ4g
D5MhYOGt2m3qOsKt4kCh4J68WULgXYrdQftDSuSCVqUu2bS4eTzl7/J5tEWKSmEH9u3dkqukzgDD
tM73SD2rTf6NG++peXOe1tYHyxa3Qu+PuWs+cZsGW8Bt5ozm/Rk4sFfbngKINOt983DB4YQAFHgN
UqI3BNRklS074tO9lUhK1TdTlcPUU9iZ8EYdCyuJCDz5N9r9Tttd/bbZGhTesKYXlfVESn68xN/N
/A/V8AtGpd63VpNZ2EQw7aa+UW2EacLpBUuRE9HM5jVoiMtxj3PNJ/RyZHZxLi8AKhOenckx4PXp
XLZqUXHoHsBhBipmFPL7e2+Vc7YZJeWdBCQGy1xdJNGWDIaV03z8U2f+HBxkiYMWSE+f5PEJoVw3
Or2KdQZHMMjVE7f1KPrX9PxQ9KDnHN74GKqGlAix/Ko+z1DIMPZ6BMLixd8vjNKMLR37u9IgzXvZ
st+uc9Gyuk7GWQPfw4cc5eV5nOYLZxa8pQL6+teD31rrppIEKt7zZtztgCTs01lYALn7ex+NKemQ
06bjY7JJ3DDaYhK8pnQmEZGwhU/9OIdtaEoY5LH5jvFBhtogYSyFH9vmnJsPcFGWrJRAqU5fQ6Sk
2YZX9gRoaq0QqkqA49j2X7IPfsL94RkWbns+2CNrGTypUrUy/kh3ldhgO65dVkiaSSINddkpgseJ
xc2jHaFosjTP2OSPckQ5OO+D4PNv939v2EgKLz34r7J7RuhNwaWS+4V8MVPSNITgL36Xt6KdA+vG
Yy45e6QHqPR2Y5d+KFmvAiLgwhAoffy/3CbFgB++C+4GlMicFSJ20JLjsSnmoewKZhbFCVrZLS0c
+GR3gAfbknKM7s/L+ThfcxpBUmkLJ+FTgZXm9f1HZOp5MOQqUonc3n6nzb2rK30bbpV0IpTdRaIw
bq/2ZoyGmabKhP2QbsoHoHaknLaSkQdfGjKmH2+XGyJkbx1O29CH+Ueuo1Rg7VSnbx879SNq3GnS
g7nfqItLdVgW1hN4WlGeRaQOxSWZ5dldBzJ7DDm+0NwDr0V/rplmLjjkVqYmD96rEUZB85wlFulj
wTE8l236n8MlxnbAEvR0HcKDBt/DJZ9cSYNrbEf7fwFbvo0o85fklZ71LjxJTo4AMlbIw8RNYsxg
GcTv7+Rgk2swgQk5G94WGscx3CpUSSyAiJzW+reefFNzSFMPbJIVhNoxfppSP6OWS+FIXsgDrqk5
zqks8Y2gH7EDBYlsd9y8u4Sdgp52ppTAfP0WjGy7LZSnqKA2BD9NVLyM8gqw8+YzY3Xfpt2s7PCx
VaCo4gK/edDAgqRpu8/nMhjUcZOSGOQZdaGlxUs771YuEpHDf3+gMTPrBx84DPbaoMqL0rfp4KSq
3msLWnEr4BckQZEpNu5LVVoxVP7MyEX+Gks+u6olval2Mr3hg8qA2vxzW+kK4XP4r5yccmlWslzw
3IKOAkJsDPLwmv/nwlfhpMwgHz8g8CT7ynbvuqHd9fX2s48Kk0GITUtIjflnSu9S6t5flv+f20EJ
fq8uCaAc8UG/H/0EDLaKhKIgO+I5fqzgJ/yQUmFL+IrjwGVnTQEln0kN7oz90Vl8mzz4bh7rHPDW
IU9hqIxRzf+ug4U6UyC6diZUj9PRzslykTuYxyxsPUtCtPghMacESJqP1SNiEfNzcNYw0EUI2ncm
UsnHLaSz7sr9rXR+FDZNKdjQNTptjayKQ9uL7Vi9Bri09SHDdSQYoB76PGJ7VT3WBXkVG0FNg3ol
m5w1uRmAW/CGasUUTYg9lavDy1eTpzrYdpEbBFPrRSzzcT2Og37bv2jVIubV2YFiD23e/3jBU6d6
pRplV7pRAML+yhKVNKpyTB7FpmLJE+Ekc70EdcvkqTetrqe0DDA82rsZl9s84ZBBRVcY75ZJ+CEL
Is5KkQoW8CU37BZd9EhkQuuE8QqES5zhf2X5Gzuc5GMzSXUjQ3DauaSF3Zk87HMb9qPYAsW877QK
ZNrV9FX4qqKybD4VyvifI6sCYfIUmWU+JOhRkX9ewT5bLo7OIiLVVZ45F3x8bAUjYPSn1V5TIJrR
OfV64grChN7PMayIC9YS5CskVyAtAzgi0vQnmJGvfmKuNP1yG3nX+QOwrIDQa2UPhjH1jEvctHfX
lMn0RKKbGRCxJfm80vDsy2ch5ergwMNjXDBmlI+/Sds14vDBuaVPPsqj4yODKG679FS1Dp8wy8st
JhNRewoVvALksbcMGs1iHp0MYsDP7K9EPLTZpOO/IbF2rob+tTLL42xA5tj8V+BhlFusjIorFhyc
dWIhzxW7mjOjmaWuQUhW9hcCRc4RL0nhj5sJ0Nx3pWCxW+NpoDD+d3vWlmGCyqhpHRHNmGnZ4RMD
eLzE2LwXGT6fwWIodewM6J7mXQch5wsEbnd09EzSdtTvuCMnybNckEdYUwzwBylm0OaS95ZdJ97S
5qNcdj/zkAkVsrHysTHa0BOf+SJl3ZRZc73jixirUJemtiRyiSkso7qMes4C7fjL6calaPZUScE2
t5XqgDo83iYeeq12lBUVpIyHQRdYOWCgiaQVpZo7sBoIxAYhrywA1kpGMD6pYvheAch5kb3deDQh
rAwsKvRxVGuAMMIqa7SYHY4kOdorifaNSdNWUo7vqOPxWSZuVAo+yixycZd0ikPHas+SuQq3gbkL
3NyY3EI3YuzhaWQkgJawjQF6goh8wc2oUHSP/lo0Efp21rhBzOurscQsAXCfb+FL6afda4rn7H3y
4wyjY1zBUbMURZ0vBhBNyv5kDUJ9XhPXyWmmxytyPAq6PUKlBN0zTc3e+kehSKEu5izeouSd0cx2
PXiExoQHAsb7HInK4g4Lut819VNDHa4WQ3loEygaBP2GYhYOcYifyWQwlSAH4f4rHIoxGtSLVP50
fuF7KiCioYFwibb4w2jAKmFuoAopq3CdZtcgZD5ahcQHc/lvkp0GYGVQa95dA3bU8SXuokMD88J3
b2Gvus/j70faHIGhViGqLYDZj1IDqd8pGVmTvDl0oGkXcytYc2cd+lZXBuBCNSypP3Utn7oX4Z4A
dX+2tssHcpY0cPnNIZFrQa+ZuOU4OkQebWZ14w8BvdqSdWWONr2jtwVKbytDZqnyVzGnD4sdGs4U
5Psi0geIUmUfO/XN9CTfiAvOLpw2ovw1GVD84bPt0fiFdrztRwBd4d9HSxacoUiSN3ce/bDJmfkR
hC35gljJGeuZ9McTad8JEcYuYYSaw7rJKJcUBrtga70fHx1mZy7O2sHhyB6t0c+9+eTYoszNGf5X
wmwi8Z9mWfzrg5/ZBOSszJR6Rz43eSn3YlsL4I1mWh+YP0QrLRYhUZaEN7FKmaeP2jjKIb5eFiWB
RUS8w62kyuFR+selNjdB2M/XrKMrF2CzoGcQRjKQUQhrr6+5TdCVzValf+iUgUK39CatMGyHowoO
4wK6zVoGIgmVYhbKBDygmtfPvtLLn3LNLUjgcmQFLSOKPucl1vZbcu8P5Dj8Y/9+8wBMvzyfgUMt
o96ql86+TfTuRiPzMkNwdQWFJem5ylabi2fpLETaQnqrEktHH0E6Nqp0W4Gpy0VE1tDKFJ+JXvAg
W9vrB1+YMyI59pf+ec7KO4p1zkOhSaLSqOfZhvLOR7Bozy1HsnRQ7D/NC2reco1diqNV1pxBuXwh
6XPtGjv7XVPNqw8mOdktjAhImqtPBOiWr+l8Imp6cHl8k8sxHa+bD71hR2Gfa1FKaEgIVWkHFx+8
WJf7R/VuHTqRObTS0EcFiMTyCfwj8kPYMHB04RprX4IO2y2wViRqb8s4EYfFZqs0YKV9giRV6Nbq
NwRhd2UHtRlNfkshXTQ42gpmxAU/pNRvWor7Hxj2c1kxvu0W39L1iLYS+B40vIcg/7mxqP20gqDD
eQc5OPeuRrotvUoTOPzEnawPzmK9mxYjDKkbNwNOF37dFzzlpfE1xuf8jLJTew3qLcqfySG34/Ae
Zfe07tcoSo4RkOLUH309D+27GDGfPMtEflLtSyW6k51gUT4/rBuxL30NFKxsMjXKPUg99thIN+Pm
u2pPqMh09rjgfqAxk8k+CtUUAbxag5kTePEX/RiMP6maI+VWCUNoTIbMjfYuR7CFBljHFI6ts3ls
923TPJsDRL+nsNb2gHro+Z/Y51BigvDwY7YFQZuuQ3+aQOnCUoZiSxOjVvAAXqiQQhMPgGTmD2MO
kfUXJkLCBLPwYFxNiS7BDKQH8pvn255FwJ5TDjwHlgvzE+jx15uGYDuibDX7niEvNa1fhjtcMvbs
ozbzcsEWIhvG35okAV/XyAloISeTTbULqJ8b2PvkeDc7nsqcntSPhVrv9UJx3+kyQiMHuW1ymIQf
NcBkNJU9nrktaAF3RAjA125g1HjKeuPh4cxL4AMPVK97rRGQicq5gNp1xj6b12OMEvpTDl9LsmK9
mg8toxucnuq7b21n4WGEQav9wx1STuPXROBCexE0tbPHBVThyOkCRIQLzBidM7kirSLK4LsD0fH4
pehS2lU/aCsknOGpGYdUJQ3BumpSKu2dmiG12wAiotiXfjVr2jvfLucyyRnrKPVwsC6iz0XuWofv
eDQWXYNsvpAjmW2S7jjvHJASeAa67F7Kk0KTrCcwzTeXgjXSsFOfafz+RrxPd0nLqY/mQt/AS3Em
cYY5HgQv4RdFMaUfhUEjky/N193A3MsKnELNzjhhiKUQrmByuvhQkopR3S607oUNt+gbs0hdFSfZ
eFLk0t8D88qTWuIHzyGFgjWB8LzCJSFl4v2kgA2+ffC+rM4z2yKa3VHZ/99cNaD05KVTxTNF24Po
MekP22TPjCsikf5+ReNtZGoN3Cggna4XyHrR0zGZeHcPZWERXeYtIGaxfQWTe/D+L2nRqGlm52il
wxcbTGhU/y9xTQ+iA1bJazJXvjCSOD+GfVyhxxy3rYx1qFctGB/0gDWubHXdn/DciNRjW0yttAXx
RhEJhTSmp0kj9SibyeO8CzeR1ZvvX+Gtl8d7mnn3Nrd/u4TEIywY1wAU8qu2f7MYavhjPtMjAz2e
ZPoMqD2KLuLlWck2+p3XapUG+Fo/l4jHMQn8yTxlHyAk3J6W+cm2067rjMwIx4uwEWmRQx12zvq+
8W3KMC15IGowwHxR6uqUZpp/C9R7SM55TFYX1XO0FTqslnXf1456sPNvOjhmWZFePI1bhYMvQewG
KvYhlvUuyn8InXPSm1/KvxThCbYfNpcHJZ1orrOoRymW2WfOvM+R1Qve8fDgCmt2Dx/C9V8YLSGn
UqsztBqbRAdVR5P2gkOYSRuP09y8JFysxfpJX5RrGtedaKnzQw7qAh3zBN0ewsnw/hZxGl3Q7jr3
rHRU7B/q1XiJ4aScAvqdpWM5Hlwf5DfOAGCs1wQJnCSu6XnjYhjKp19+mRXuiXXpG/A0duoRJQtI
wOcPvXefVCHJSjhgIIXhI8LCBlLJ3bixhGdR2x2Mc+TmQ1pP3TvqKuAZuSUhwNCMBVpckODeQwQp
xX97+B2HKliLQaxoLel1WtIZqIt0/xtLz+bG1JJF+GMoWtn+nP+fuJPQuTk7D5gXbwROloVZAWmI
VnJFzg6kaPhc73x8CyxQhYkfdID1L3gNEX5fkoMZm/828waBN/u+0zQOZGRfKa3jq5nxXhXWHhR7
UUWYkiqEcJcELqWLi+ufZTtFyzy9AVGcyL7ULpV5oWJWGd9Ui0OkE576mwg8MI/mIPu9+0Ch+Wng
OZGFbl84Dp0Vfq5MS2WU1Ahr0YTKEakwmNKjwOLEOB9Wu3wcEhDyufzloVRr7uo5PkOGSZX8i9yf
xPxEryDCwogBDNOjLrZyqW9LG1XkFhpOW4Jgg5REIulZ3NYRrhNhaB5pPxsE74urhL9I0A1MWtW/
fY2LpDDsbFhQ2O9leEVEPA86NRpjGjqXSFhyfuxHsv+cKK+fZ85G9ArN156wrGi0E9ZZvk08nv8l
nuhRRRqxbeDdsBoETkJZWdspJhxKUpEPhekEILCvyyZ6ZLzOQTmQaUxyn74LZyh9cFb6CtEtluTX
Mqb9uhP+rHiAqasF90FT7hyFEjMuNAs+cg2GxweelAyEQHZRrBtDKr6QqVLe+XLxxro2koC3ZU0v
IdJ/MUxKHxGoj9goC/t0LCYDP9jeDH0OdjSnT1RELOVaz70nNuDYaZNcJf53Dpix7oHBskM6QfTu
Cj1omyudJwNPNlxSrARhyDjbHfo9eMbgK08SeKEOApK1Bij1v19RNr80QWVXPRs0J7TShGsJGTUC
fnbkXE88Kvpy4ynnNusS4pbL0YWKNbH4+oDm8wRx/4Qg6AyFazmzvdshO88QLdhpqwPZ+uVhMzUe
Fo4gxkDJH86Pmx5HN8Ab2S//ByirhheOuqae2X219WP0O7YEu7dFgkOMrNkDHEVSNn2UT24nExRX
Gqz8rJGM+dx453Nmjjy2GF45T9AeXaRZb+bm5ic4/b9FZIbgcFpFoLm800zooGLrVB7ZkHSES3sZ
0q5HLRq05O5iSMpN+s3JKYA6R9NJOcTxlrCfQLajMEg+3W56Loi84Wgnivb/14yeZQeEnxqxpts8
PLhy5Bdyj8EJlVWkHV6joWdttEA2s9iVoK98GkmRe1vltnd0+Ie8hdi3mClZc653nWRsDaGvUlhH
ixNRWgULaRV5YfyOi1lR4GY+g5vWNRdrxem0VJQH24WUpK/MxsBcRZCstFxEqbevcKansxoCdbGv
2SAbQVtaUBeRSil8po0ke0LIAZVBQvkp3ucWDdOm6HgSeYqBteIClk5X9TP70xjiMUQ1/AmUD6ar
OK3FsKT5s13EkuUpqiA9cvn5XV0dsN7aF7fYRtUZfQQYOpw2hb9Rdj/8RIgX1EZqv7tFES19LabN
STwv/4JILeeXJfBeNp7BklWtUJHaGOTfz6kIN9vbHTTsD9kzLvgC6ZivzSYKhbF7VAotfgZs5Psr
pgs8VCC+T92fLaute3fmgiiHCEDGoemF+X3BWOKIEHSuuhYkrpJ+jHeh39YGatK132zmcJumaas5
gKYt5Qr8r4mJoHbjbF+VxYZWxxad6nfHDJULQJC+MhEoXsOHcMIpQR4xmp38aA6WreNJtdjz3X5y
uuo7FVTK/KLL3Pf476BgAyhzJWmvLWKGHCF8XAAVDNBwV2FDMk+OZeu8+Q9U+vq5F17IpUU9cDm7
Sq16ICvsT5Ye8zuOv/D3dEmO+Xc8o3aNCqiF/avV6vwVsJ2gVdElJ1sOGOn1UkLd6UkgbbHpM0Kz
WNum8jZyPa0uYrZKWJneOi/2nyVXxgB8SDluMDvivleJNJ9InpwypXZ2vIl56PnAeqv7wwPmj1I5
H4W5Ie0INqCv/zxCZ/6SJhU1lTF7NNiqOv572RKmuvXRg1DpIGTXbLcJ37azArn66K1jAobIM85k
EXJFhGIkohpPrkJyPItha/g+gsTG6ZSYE7DdrPvybC72Abc8bObXmnKy/pRKiupZRQWnTaZg29yE
Dpppp+bzDGX13MZkV+vlRn8NksBC+SZz3u/9kjcMTDQv2MHOLvY5BIqqgtfvW0/oPpquBcCMFjG5
EzskRMgs32Oj/sLtab8S7kcmCtY+uA3qQBg9ZRMKrBMfh87v+r0tQC4TNV93/+3JJFZhuqEtn3Ad
rT9mDJNKeavqz+/vNd4vQtleAHeaZOe/alZzCLlHpVIGKn/zXhMOIbqmu/ZXB2i1qeAFc8nYsKbP
AtJwKWtDxk68n3ttCROOhVJnrxBPRC3mNsvN5X44o+4ZzwnnGfrMbbHbFySEdCJ1SHBBZePdxMTa
l5Duf7B0L2wUwcqB5YjkRU+X93lnKl0Ma5mjRXYArakCcGAJ03K5DYDaflAGx26LteHf/WmY8Skz
F7u68l0nb3A8Wh/WjYCU2wWz36Y1hG9vmp3DTbabcpx+e4V0smcK5+6R6BjK+fwkN5rQgaUQf7iF
/VQ54F0ryz3V7C2wW+hiIUS26Q/FPviKuS8qfUnmYQswCLWdl3pCzmbKGRfyla1jwkRbeSAk5+CK
q87BCcAPGB4+Qr0fLj0Fbj3PrVkJusLAg3cwe4cw7evGsZfN1yCrcPeAu2fqlgKCImxwUhSDcgmq
Gt2JwlzwBkMVDDzqFoP1y9xrbX+28bcFw07e3goHuFNrTVjjKgMop0UN0kYKE3+C1bieJWHspxdB
IO0jPlEk6E/vE7IamW1NbHp9nnBQcqml9xYt07x5ToX9sF+Lpho9k79x8gvSpSgrQRlamfQwRUUW
PZ2MGpm753+rBfE+es34r9mUD0bgPKAqtx28M0veoUMV3R4lAQDP86oz16kSZxDr+cEdDzDXEo63
fUIZKUZjnhbncbcCFXLYmFjiePqKun3mBD7IeOJ/nCiIRqn6xAR4CFrJwAmkLv8/AHOg0hMidrR0
IL9ocH6L1CQFwEtxIWVa2+3PvESqd0FpZd6+1lL6gVQaaljuZ1PTTjcqWLwpcqMXqFfwoWL4yo+3
z/oLJmwDwgALhLUzUpzzoI7Jo7DO3K0ZzzFg6GdGGn57HnVW9qAhPPugdJRuUOYdz6m+e3JZ71Em
lksBBcpNPLxqhXTZaj14+90jnNSWjWOCubqSIZH0K7A1rZM9LkZk9LOHOC1swx0oM5iDhUHIKuuW
fMeZ0jhfiVFBYmFv4zWZOuyOp7EnORvfNe3ZqeLhE/rmqVxOA6v7XiDB2k+IvSxbeGAqAzLoq1nI
u6D+60idE8Z7gVdi1hopgpktKRhAxjUpr5zQ+YRZL3X4Ldy1Xw7TBwdb1YgB4kJAFHObMCRIYMDo
mQX/uhLnkeRdrIca/aBI+Wj9vnig54FTMURDARS6PHnHcaMOA3oAeMml3TP2vLI4+kejwQvPubOg
hoGFyrQiPPuyRRpWUxKy9FOMLDScoVN2dK1FiSa7vNK37UZ4dLtMs2KRrQBimAfw8JheZQDlReTq
sjjbAAPpUqGo2Ypy1qp/vY62/9TuDuZDJ8xVhD1exOWpxLUUvQSUOz9sNKgY+ZI1awELNRslDDtL
R7hWr7nb0qpthzSAzhGqWq3q5aYcH2kvrwYyvDvidXpa7rWmtcUVGMg2byww4gXJeLJ7U5mRsmTL
josBUoqPxXHEVf6B3GmKUqsCZ4zF57OKnHIDefPlJF0DtKVPn932OL4A0QRnUJEqqNiGx0VGR4P4
49tU81M0lpo2a9onE94HgZqprSYdNg0fu3XBU3pIzSEUtGSdR+wLdVF3+nYluo7wSbgCySGjjcBU
9XpyJ2r8l5j0vDVCn5EEPEH/U39ZvP9fy253vExUA46Mki4KqVx6q1htdYlPqv5iAzE46uriE/XS
qCm0JH/XLHR63nk7BsBMWnHvPkV50+ZT3RxN149davKeayUkD+lAk8eslWBJ9SW/Ghw/YTHJvKED
vjML+8qfCXwhOFmKGDmRdHuo/QAL/T/HiTPy6MMvp+JVToXpcSFkAMhxAD56Cbg8RwwXaia9G2sh
O5o+bWHqzzQG4C+7R62iZyDta4lTj8wKbLOs/sp9Zc58kBZ+OT8rimYLXQ74+XAN7t/YGwo8RR4m
3iaEpT9SRany7+utTY9zxgv0jnnzfmvY8xhUIdvB1537DJBHoic+w+1ROhQm2UbJ2UoIYB6Z+OVy
oVOHo+Zhy0ZjCRfQ81IP5lB0VPAWl6aknsxsrJz5qoW6lWKkP70Va0KSaPKoPfx/gSQmR2fxJR3x
ubNeGSVUZrQtnip153fDIz6lRGJDG/pZwiIlagSi5qX/0OO/muc2KTxpiG8+tGDtTPy6n79xUXxZ
2ebXAeIJ0BdR/Bm4FJbz+NTKmF24rH+79m2K+oXIAYhdNb3IQlbqWfVx3UmLvXnc2xwaBBA9Ihup
XZKP8WnMboYJJ3xdfvAPDgCfd5F7zp2WAoy6H14PnAmkV9+HMbrbh1Bc62POk21cZarI9UOyMOMe
fXrkHk8C4RKO2G+Y8txOV+fhxSax7GxLaiDpKjGIwBdPbukKc4e4vnBT9f5a30IFZ6kA4qQZvRky
w1QvsUcGKxEi3QaNR4xKnlloktU9M1G6oSJDoAgowoiq8E2uhoBKn411CsUiWPVyo0zoMTx0B7a9
3qcUhsP/VNxuJ3WtjfL0KgeuD6w20FsTZVf6l9F+/jwyMXeYfbaK2OEhgA2PPyXycDCJDSDhRv6p
wx5YIaHFbKe36y15ZfZ/hSG8jGWEcGjM4lB1/6Miz1Tcp+aCa8kx+BmHFYSFiSoTMAvBdvPdaOAv
K+JMakaAPx2Bn2/V0uEUN5WuC7d3wrIBQCJXmUbZtV7NImFE28g78b7iausv0Gis73K++HHsxpdO
lXf9Z0Vqfwj+zomcp/KSAy8HwPCsLDa7ThyhzIDfXpoTRN26LJPEya1vR7nkDEvP3KzXBAdyw+pg
AhqNUivsbkpJW0fnAeBbFOETtsNMee9HR+utOoTKv6u+Ys8FiHLO4WMI5Auwu1AI3ZhtsTp7YKMu
BAuGtCBeIoSHB5v2O/1nCohFwEtbzPI/KJ71g6lXaZLdS9vWN/k9jQBpWnd4FNEtGqSud2w5ZfTB
EmSyQ/d3/nkVkPzKRaTtIelxOH2Do1HitKCjz0M+/3oJajt2V7uOR84PEEv6yMDEtBU5O7haRELU
KqqkXNXDhNIQJobRd2TLoyjdfkdrGz+DWp3ojbA7ahAJqp1YfJUjq7xc9KDsLZkNTN915KT6b9Vq
sFa3f+yw0quimFwU4wmUB6soIKkotZmIMS2QURBI/VTrnoD1TMoknK6exRpF9cog8B8U+90A9gF8
kw8FODslACLc2uNaPFs+WYbRpCyITemDinHueP+d7xli8qDv0ewSzJXrYSralXteDmHRErH1+EuR
0DzlfBkf7V+ps76RQvGrl7BFuxOtfxiUJQecekcZEIqRqNdlVzvolN0mC4wjBb6IBuwExu9RbbGc
GIeN+D8W53VnyA5o97xI4UL7Fe+Ijo6Ez8XpVetcsWnrHmPzkf+RN4Do+8+n/+RQmgV/RDQSBhWq
52AYyYaCfAxxCTIx7NTljlCu09iS17T8xng31aOZPxVlLa1UqBItg4vLzSSNuvJeW4N4b5x+ZKe/
ujNna+61mS/WDk7Ql3CKboWrIifqKRheI4Auy5KoPeajjtSCMbNjB4LCbrawHyx56SrDduuCTU0k
idqjxXLfszpJy8yVv4AuItDiIaCcSbt9HYYK02IN0oxKht7NjzV3XknVyUnss2vSYN0T6B+Hd5SV
nqDg0qDRu8jr0nn9Qiv2Q3wau+ZeIGExQ3J0akn6wWeXRHnaMYBvggkEcYqn4kjCwl+LQIFFfpg8
f/9ZjTK8x5fDJleRnfTUPRSL18N9J5hugOvzGMyTQX40pHBSU3pWdS3Len9a4Sf3HCizJjxff9qP
G2VY1hkejLEyqm8d8piqDfOwOtoMyvnG1PHxqODkIW8Kees3B3TbjAM8c5dOG5KFWfvUlIgSfFfS
E9EUjXuQs8HQnPNqbHkMjnpWwa/uchbCwY53HDtA30flkGTPHAXRzvemtKAEW2zeg6Bm9pIjki3E
yeAWl53nOsqZ0w5pLRVTRPLftgtEq1rDUEhkIx1jVlfPcK7FtnwivJhgN5ebO30ljVcIMTCzATLb
lKjs/P7DkqsSA9jVudrwt9Fu+ZytuMyT6u9EX831mdEuOL8KVblZMQWB0TGWvqrXVYLLzGFIMPsd
wBMEj7RSjaqIsq+kH3tXpD27FGkD+0iDr3YFBGMCg4pwyWuvjXB1K2ZBjvbOyfvz8clH7E5+Wfsv
+2c/e8Bg3tDNNDEy1YfyDAr9J7iCaPmyu50k98+r4vquR7aaYspaqFmTD50v9y+DLAfy6Ws95vra
wmwGKEmfgKRCN1RcwRc8i7Fd2UzrKIGxdq88dwc5yPBz5kCH6eBH8Qp3mHf2BmLjRV3FgEsagFHI
oEfGo833RLcczKIgjwzCsGe+3Sh0DBs8m8qsOkAd7OaF+z2qyvl6LjudFURn2WoW6ryhn0DXrnHu
0YHhRgAP0FOIUxeSYPviM/WWUWrdr3lLDuA4mN90dJXX1bEBlAt3maOAt5Jyg0ahw/tvSD7xMDLH
+XUnr4KHBvKQAhE+5oX6RvzI68Fic7y2yRCAXWn+10Qclkm8hoSt07KnQbUKTi+fpVt2UWWr8lM7
CqVFSKqvfK+0JK5gY5Ad3WR6raaYjVgAe1FzNXCN5oruwOCLRfN2kdYEIbFrmlpnBRvQSJCCPS7U
3I6V3XDW301heLCViQ7SZnMCZzLExrbrqh1vtmp+11/ffmlNEQWGqwqRlxSBrOHoBQE8mKfsxr34
B2/MKiJF/pUMeSmxk2aAum5idQoPZF1zBhrTUzDLj2VSZmKMu3O92czuUzS2zswSVu10w3Uz03mC
E4pu6fIpAiVspgVxdmnGm1U/dy48SZ3OwNghK8o5hBv5Q1z7p8j3oV+CqQQ/a0S0kA3gnp+lz5j/
YwG/jljXTUl8jRKHuWTSuPSPVxy3RnD2rytYO8Z0qD4wBWyVznMvvvu6x2yCirJeh3xjfALWrX5o
kwDScW1Bg4WpPhPFURqfB1+8jfJNoHYguAPA5sTHrmNCY76o0JqOECyqDgsn5KI6S6sn2CjU87ee
Fscw3o3PHTIpenbRGE7DIGAd73pB2NcFuQMpvNvO4fui0BWZtHkjsPea59dxCNRsaBmoxmLYuGue
O7T/+NWqFaCHfvKEcnlH2FSby9bgJVQrve0uYafb299vdn9jbPQ6O8+H3v+AFuw0ZPP8Y1BXpJXk
x2J0b7tEKjrJZV6NUHQQwEfObiLuFRepThZZTc3qB37UPZmUuek8JksOGzCQXNPLlUS+ACe9hORo
F4J1jjcaF5yhZ/Vp6UchUNU2vKG2Isu+1Eo1jVWmj+MPqoh/HZSZ7SsSoF6CwLAFNWW85LqCAwh7
J/WC4+GMGw6n6jGx9Le0Ebwe44BOYgO9GpaHCD6jBT2LdmNxwTCQ/skx3UOsr/HvTLl7zgIl/sZw
BadeTmRryYf7g/w4uGrL03ycmh6tdItnGsFehjWtsVSDaY3XVorkiPdvYryS8kN1SjWiBK1z+Eo4
Yo/PZp4tBMaVylHZ3ngaIUgf+ji26dRWFkaViPUkS8CgLcgoZ4qKs4wRtLSZpNux2ysWgrbrQ/DD
Qe3VwMnvGcrtLJU2bo7gHibK9hZ3vd4EWTAI3ZOfLWDe5PckrbcexlRQLpkeeaxuaV8ivd2LvH4a
ECOF7B7fGp2xok32TBRPUutIuLyVGqt2CV30Nz1icxFDSo7L74PbIMP4HViEynoCVYZoYxr/usw0
KJQncW7j2v0inqhvMbs9vJumVVtdcz3Jx4LLeImWClKun81Ffohkezy4WqRnc4A1uQ388bz2O9t3
dUpsdJ7Eq3SLiqRQlao+OZexaD2qRX3zyK2fyfIB6DsyNYmPgcXOb9layl2mfbDAjyaGBphF5e72
+YQ9hWSh2aCT0vU6DWdA71JeIZbI/B4s3wqnw5LRD908sYl3XDvbuM+e/6KwP/T1A3syDZ1qei8f
XhuPD8/738Ds7JcaLU650CcSnHZjV7JnZHkA1iLxYOs6VQ9NX8UpVutURWFnPESBzvFpKliyvwMt
h3W5DyROh/kBZXumUtgxUOLQQLkvID0TusOwM+WXhNBzNQOh3Udpq0bW0WDiSQjAw4Vpott9k+le
4L3+y+hdTVMq4IH3n/+ue7/nv0nGM/tK8ECkO92VMnQbV1TDwpcYCtBYaQZT8YgAWUxS8RfaeCMS
Iy2903qXZpNKvoJ6zx0e+B3fRAFcIVQlzwBJL+W5wkWtUZEeKH783LTQJAGounB+ZcJNxbmMwpQV
wkcF76QLLYXD2Wu/2JW7y6HR5I+SohGpLWE6HdobV9acci9n5Hj69yHPE4W6yN2Tvawxxev4JGfA
7+3vvTQeuC5n/Zww+l0DAUOHcb6R0OodWrLIxj09XrdVwYjI3hjSfst978jlfZmGuE246j+pu6X7
ac/i7tm8JzYHSs+bGI+rODWFet8mo1cdaU16LMn4TOG5iM2CpSGgA5bNN0OEfEHJUv9xR9MYDRk8
HDcMKHwXBJ0t0fhtUQaEw9T4R3t5ObFWYm38KCUpJbTw3hWURs6fbW/rfUvgfpdPmTbymBKlYCyg
rtpVQwdA2qtIlne/coptIKNWGoatUw06YVzd+rwiACs1B+gKo0IzWIVVP92nRq9XVRsLBwOzCbK3
8R6mblVj3zP6IYPVQY+Y5/x2oJ00oilRVJsqQR6ayHchbqhneWz3WV0PYWThxKiBWVDKqdscu1j3
ZAdZTbGoIbVkc+AhnZMFWEPNM4MGJxVqMIHxgAAQyOFp8zGOV6J+FjmbDHXqAoYLVbcUR3km6ZmH
jwJ+pwO2OfBw9FG9KRZRY0o9A3qtrhKzmlxl2MjtoUMQvGdWdW1Q6M1xs5mGW8rxupK8dTGL8caj
0LoWQKTIo6DE5o4SBhfl+mY4oEUa0XojX5G22PZOpklCNl4vbHIidIeDZSDGbO/UTzyzVDW9aJ0u
CgtpNc1W7Dy5hwpMjjWnqQLqPS0wlNrJBTx+V/xaEWRwrcxEFYpl7jlGJnCvV4bwj9grxf94u34i
KvxVG3BAly7fcoO3AituDRvZ9B5HNKox6ueYlDHd0PIlyyPl4nWKNoIcvLPYQF0EasNhtX37nOe/
G16tcehberAVauoy7VKH9UVoTuyNlcLuuZY/o3RrTJF/e5QkKJM3yRTMwc6JFUCMRpW1LeFJzQQ9
wk65KSl0Nzn+lT9IkEBpRgqJMj201WLFzC0jk5uMKHvcCeSxunVBKlfWMZ3EWLyCDs87FPin3IHl
Nh645XG5LpdbxzKB9C7d7BripDjmSszkfo7Vy6/L28EXZuJFmhMeIMgG05WoBS36upoOSRzqKRVs
8UAgYMyIt9KiDFq7YCgE+/uIXrg/Bpm6KvN20YvCBuAbAhgMIaS2N388NAhLinOHbbkmUTI/ljhZ
nJgeEX9/esDXqnwqoq3UKPdTtM+pKKycZCVZAEYblQlQCIydz1oUFREoXkpC9++92K3cYMYE7917
RGSyHlWa+f2wYVg7QiRUVJZ9wmVyAv9C05lgqslGeIE6U+iua5kG64W5u9OZ92/KiYbxh6nvHIcE
a8JHFTyFL9ng4vgowYM7MhUkzlZIJkLK/Wb5uchVmYQ8Wt4J/02dINzMt3XqVs5eSvV3sLYUs8TK
OqDMnFl2lDVe/c4aWyOaAYOQu+LWsr/JzAipwV+wPp147q7AAL0JBHi/LRsIaM7phtXe4gq/ZMVp
3g4OvUmWovTZ4kNLRlUxDm7l0AdJFXFR8QbN0C+TKk7gxGop1D4QSU0X5ltLSUr+FGcU5hx/WwQG
LPRzcHf8WqhA7U5bksIy6pTFvkk38qThX2PLYwNYRUDzCD12mXtlhA52VdDxgFtg1+lG69vCArTQ
D8SRlVEjmXpppbQGtYFUtm1AJbZqLJdXSqzr05VH4uRBuvChSNahjhFBrRy4X7/PzRmQx/i42LNA
RDMrNckRORwV9S7np/2qz8DM+DpDUF7fWf4QTJzcSVK8+qokYG0NxZZkzN7Rgu9VtpOUk7RSFS5s
+V0CYTBFBCNgPkqBJ24CPjARhNI0WKunyl7UF1dkgfCI0XCY/gjLi7oBeWT3o3IJtpKmzW8/2E/S
17oc1hKDOBJSr5BRvI8yGbCMB3J3DySKU+jRQhdWDctB11aJdpb5/Kv7JKv9ehQvbQufWd1StFmB
WFHWp9KtB3ztF+jt6H4PTGxv94qqCoGvuOCYrBksT86L6LhlDdd+9MPXvTd7kD2LzvnsyIzR7kGz
VfrPV5+AvUOthnNLQ+Fx4aWHWgyF/qtl5bNeGawgFKX+UiE+JamzHenY4TF1dTBysr0IvCEV7jDi
55IJR+P+cB3n6hUAuXxDaVgWo4WwzWNENUKP25EFPJPTvvN5x+O7SH21tmluXak2L3kBp7RYsrLd
YVsHJ9/Tit20GtPGWpGELf3au6LAF127GodHyYUj0FRBbT1G6bzBrvvr2nOd+nn7H+A3e1XaRa/B
s4q4ZMe++Ud9CbMXPD+elllewDq8fQn9HX94nufr9tTskbiVioIEdQB+WXVfJwdy4OdAGQ8ZpOKw
Tj1NCNiMJwskVreH0If46iK53jnIGLOKO+a8UWQvzM28AHWnF1ubxN6Vh0PISunafLtvezHLMwkO
erHsYb9RgQRvX9arcNWziPXaoctyEtnvx0smVpNn4/+G7fKkiZx16y9lDyRPXTUNBE1S99SdoDkm
dQjrcum58DCfRbvhEYATSweuq7Hs0pWpy3ECHXh0Stg1IAVwtaQhaxfbk/lPHggSv46YcLsVMtDn
00nvPTAY9SDYTxtWKxz9I9rTvjZJky/699M2m9laZCmd1hoPkuv19aivQxqbmAgK4D2SBuwJAG7Y
hrtqSavYkiSTchapV1ptbOsrr3gOxcIn+v1eE/nnPYXrMIq3MMukL59HEA+qy0mxgOh/QE7l3FHg
yNVuqmFjo9z9AWJwe3vZnzahiAQYhuAAPj2lWCdOctszQJYzbH5UWcC4JM51Qr4B5EJl8XdEa26G
NZm3m2gRyMi2ThVJuRkoGOb7Hn7pIgum8wTI525pbqRyU3q1Dy7WqRkiqW7GANSV7BqJTuhi2J4s
NBXsp7lopKojbkXzTG8MF0TJNOruntDW1K7H4DbdGVevZIA8IwohLO/SISfO5Ub95Zw8+taINibr
K7FEOkS7eOmtg8AJEvg8xLiIC9hdWc0Q9q56pB5G1TonVLfwzhqSVng1EPmL/7FQ5NSKYr0bklF6
hln19Zhmgewv/9jIjM0JW4UKDY1On8EfWTkZWBCfFpZKDqVTOb5XTe11wHRCiscwkorjvv5m2R7k
6zIQTePXKfnI4irGNCbnbR+0MkhSYlUqrSdHC4i6aQaIRgJjbXGTUoxEjQN9wBv+zcuyIi34mqqO
Ggb49BgvjQe8HpLN2OFwtePIc6rDA0PR/a2MGLEnm4wWjN2yTsgl8XE2jee8FxKVjjX28BHyZ2Kr
kY4dRgp5I9+YCP6RvyQY8e6ysgS8Yrm1tztTLoqLxnYamvKcs/4EUjpodb4qc/lVVA/pJrQL4t/s
YTIov0Sq/9l+plo+VHFPEHrZ+O4qWOjpX9JUsexni9OLiSVUSX2Xd58iQoKXjRhECQV/OMsb0YnS
aSIQ0yitpjuFEXnecqLNtoBStZKqPuHBovutmgd8ZnWkVr/giJjLG+eTWPFtoX7aXnY5jCgKH6lm
xzLIMWNvu1zBu2WSrfgjkq8FcY3j6+AEh1Vpnp4m9GytSjpnkLzDJ2fLqdsRN/gFwkjs7och9v/B
eS58dELTgtsd3dVa0oCNkrmx3kIQNNVD7Gh6Bia9aUKzM3k6CCXC3Zns2CvCqIuYq0VD8TZpa5nF
c3K4+E3NT5JvwgeHzJE4F/aVp1RJquF0ydIB0WfMc4s/Vau4qXPDnizsSDX5qA8uhgWIL5XCqghj
R6iLH+nzMB7z9Q2Tm6brMEgkLvV35pYQ5M7t7s4eIH7b+Or5olfXj76pIeSxp/I69aQ1Zy2bjJjs
2LRejvdscvuYkIZ762NVzXreTgK7acWbu6vWQBrIUEdS4Vp/67b+WSKhW1kf2RU+n4h2EwDfHpX/
1wjIreY5gy8DztXft0RDb4uTCJHF7Z8caf/BJI0y8q/Dg7iDwVmWfkF0HSOYb2PBth3lrR3F5Uco
Yg2oRLizlyhbixry8exrDsiOdXivyJMdR4HtaxXSu5Ulbfj1gGpVPDPS6Jdoxx4fq4AQM0dVwpxB
M5zhZXk/3l1DxxPGovEpbzrGon1L5Tmg69nY6lVT/TG7xeSn483YWNyHoVHH4lNZqxa0dpwW69hh
HkSejwq3se2+VB9Dq41VByeRrdtvp6FVnfdy/S133XPV9OZ/yTBRN9dhPKIdiRhnPB2TlZh2Vmui
HFoOJgSrdEs54Dc1diPUFMHO45vD4ia39HlW0sehOphmYV+39jQNzF4EwdJW2KxD29jsC38qFj5a
43zwrF1o1rsKrNmv52s2XsfUcu+hlDDJ56Jxc3Y9Y3+nHr66nK2sArdDtaA53j82t3fRa+STQ33G
D/Res2nZ1Qkh5uz6CypGFA0zZtO1m4fJqvB5Vq9drFwLFngqWOs5SVbHg1ge/VsdQyLoypsyC2Jx
JfrGu15pFkUId2VyoxkbdhEUhzzw/fM+SJ6VHikgAK/GgoJv3LUKThZV4zbOr/8Iaf6IbRsbFq0r
d6ZN9E8cG2P7XoJFBQFk9kEOVXa+zF2sp5isiFCy62upzB6mFbD86jUrKPIBJDRAbAcT1222FDw8
oB4p54hSL6RTKhVjYMs3X3xIEjQ5yWNW7wK31DnWRPZg/kEZiz4jSZDhXGhF2X6OX1nAn1hOL+XI
AC2O85n6q4LJDNoh57OS4OAVhlByZSFGXt5IKHXb8d+yj601mQ4D0J+bfJWrB+hp5l2mRkrIUqW9
K/EzU19b4jjVpxkkv2xaFGcE7BqgshYIz/5OOyE3d2HKC23Jnak6BwhfxWEjeNE4Wba3MirJjUzp
sKBufhMP/BYXOvy23WQaM8sgr1fjv6gRpCU0VzUY8ipvn6Wzd1Wm+cRzwYgDs09lUEnRKD7KuTbE
9iZIcpw4zs55UV3txO76ZavRKoM5veBL6xWhcrv2dg0bhASeUxdfavcZCgmk8aGJcKjbLuPL5ZvM
xtgBIScmTAkHLcmVPLcOOIxNUuJRV7WvDdKKXNDD6OYUbdmo3YEBHzg07qrQl32Qy2AHt2YZbMj6
+fwU6rYFdSjwv8oZl+HkVbE5O0Egvd7mj/1JrscxeFU63gC2UX2+QsNTe3/iMcd5bwvVD/bU831k
G8qtm+Sj41p0bUj+bTAZ/K8nqrlzmHRXgOOdgVwo4vJBoaDMowmnS+Oes93VV/lbUmUx+D7bwXuA
lgUWDOaXEcuiZOOEXEDwnacya9udPlYz5umb7245Mm4KQEP/8EHX559IPO9KHmvO09X5/gjOv+bs
R/sx9+q77LnhMg4g7Z4jv5LkLwNADSChm85uw+Ug/lgareINEQgEiErydRJjGV3OZbsvi5hCgfJe
vMH4IwTgu33vR2E9smycH9uROjZBXFip/dRIqy2kUa0oDIoafqFSh5y+G6CeO/naN63Z+wYaWjXO
dzJeG3VOGh+me0Zpgn+CZTQINp8l5LhCDAssHszx0Ax5F+7F28nrCWGhUCAehh+TrQNauwZitqPW
edqyk2ghueX65287Sv9NUlfZaLwUznJ90JcO8Pu1qrWY+dxyezYvlt3La3IDdbh2GZ+ybPUbRPqZ
Jry4S79RkXvvomZHjPwa+jk7Iodm/v2Icm/D+Wi8f3xNtraQTi77dbBUxt0/1wulzQsUu6AEk2ic
TNHALtlIrQs+Xq5SaORZSpQ/W2FE5mJL+V0+HT6lX/FBIfOqiI6YUn0xt/8+LbLPUB3/F3hdHpSk
JxQbKSHnbKPBVPeKuvi1lgnJMczpBArZ2Bz9+09gEkrwxyeNq7YqoJFkyb06zjfIpwvkMgmjUWxn
pmBhYxlDU8vytpA2y8lcEpFdOSTlIcuf5VZbcdUNnEJN8OpF7xgqpgGvb4ormG875aJ1BjeL7fRH
6O48XV3FDodNilQpinyi/g2OODnOnssh2fbh6aB4gtmx2S1/L8W/0oAGiRaoArWhXclj+6FfoW2o
inA8t8khQjEBhVA229UFRfVEf0+IRp1dsI+h1GT/h6vvjcNdEma756G/+eBbi7+cvzePp5Ya3XFq
bCUCoc1nbQlI379B7btU6uC9MDESAgjOHsRNZVzeX6mZd9VnrYj9ZpPf+GZduYLkhrsUmNAWv729
YMHzKNb7cLEtRoGsa6zQobe8NP0Ea7OrQdnUT3wrxGLG2KJTOOzioIzNH+cnjcuXxrzsM2Lw3bn5
zFDAyfR0xJVrn1vjkbW9uu1wPIWkTWPmXsTumf9IJv8dDwitpSR3Kp5CzwA4fX5uJORGJCtSXC6n
fu1YVQoZ1XKcTmysJyHXuNvBNKUFn0O38vyWe1apyLdFT7fx8DsM1YAV9lb9P8qTxgL7tPQ90BzH
S3dz9vZCt177uk5d3CJHsTJC0P8DrQPIJxaxJ3hAmayrUopgRITVuVUxi7U6xww2eS6Q2x+UcUDL
Bu7hec6DVpwvEH2yGiOAn7pfP83K9AXhQnrD9heWsz8HzuPLAOuPCJjNznbVfgW9cscEwmw3fc91
wpF9g8nzhILxG/mdtBcXdgxUHsv45bnLKtNTJWB7oHOK3t/rQp8yy67B6Bh3+uiA3nWBp6pKF+X7
0wwto4dCzFsPWC+8W9zTiKWv6OV6gjmcS7vfgiHT73tZAcK4Mr8dordYbs7vUetoIgFCINLTC1bZ
6zBNUpymL3Pa3EOJ7QAnKSOq/nNqBxZO8Gcs9NKF5iyf2Nau5gbjzNEtvUKvZBT1xwYdPRV92ggl
nrDbdrEK+s+QHRY0ahJ3P934X7wmYIp+R3geIR5diWtmOJTNVOXfRpy17Nn+H1xx6tnwMrYaDgwn
DbO0odanVMGI4wUjJgQNqrFMMl7MkMO9RqgqI/mMMW9eLlgCiVSLtxbJbkRaVljq/jTwTOaj4YEn
0e0PkY5968kI9KFMVh1SLenWm/BicbVJsICYuwK7IrrmoxVCQafyw2dege9vHQaPCiZlqVSWojF5
uGzRGJYK033CEKMohpyDq9ciF6Tl4uYR4eV+mEqe6rXTxIpD6StMTSCK9trXnlxmqYnXcdEnqDyp
SeqmRbv1aOijxLR4jsJQybLIvs7LK5P+Yk6QvCPu+F7Mhwgg9kaL/yXB1+s/YqHrUYYOffuJtlDo
XOY1ErUofS1XqhHlq+RkgQUwNKoBlRKH3t5jdmyKCh98OCtpPp241ucb/C+/hS3k0aU8TqnOFYtf
zj9GuSdPFzPJwCqmknj/r4XiFG9zg8mmt+xdom4pm8DkCszIU9OOZoIdjXVoeEQ3crYu3mHahy0+
xEVTpXjb72mWlJ4AH1+uvSNMrnmt8dkVehJDnZ9sqz/4oeQsl7wzng8c1503W7P1slOjhcDQ2SwY
vcTf8CRj4Nahe+H35qgk49dHtFgxX1cbDau9p0vbXhQXylOWJOdMIPG66IafzKtg3OggHqPFs9IB
aqbKEb6fVks7QXbk9BuqDO6OjcJxeYgs0+kE3EmMhpBLbvu3N+1/WoS5Dfh9829vmHIueSsU4oHr
zQ/4XOuP7zgFxWZMzpOdFU7f+CoULAHOcIh/0rsJY2lucmXeplILOBa9dxzrmQrPZJW/2NQUrUJt
IlZiapaiGK3PBDCvkgxa5xo5ZQbACSArV761hVhvN7EUzLxcZykBJdGsd7YGlyrN0y4C9dEg4A7k
Bd7bvQom1w9d4kUYinYXMACnE7W+6Rmb1sr1GeZ/E4SyuSMGKT07Z/CFezxp56htmBAuSzHaX6h8
cH+xT8senyCnE5QX74AAj1k4rqnwZ9BkruU3QNynYytpiBuLBq1JZ66CUQ+TcRXiC7Gz5gcuEVBW
0B2JViH38aEN8wVqoRkAuHLwRxVY6f4O8hOcQJYm5z4WFs9dtn+DlE4XORdSQbLaivKaR1Dy+KgL
q/D3LidFdu957EwixZDVknCQJuKuWKz46Fr2DzVglNxdvny9nDuEKqQRtgZ0g1O/AQUVzwBQR7En
XUhvzL1YVXULT/5fIj5qqjdKyDN0/Uwz3p14IjoimPSZ+8CuMAEzFAfuE+hh9YOnll1gDnaCrEpw
G49+g+4LjVvbCs7CAmBzgZzMyyxnB0Cu2Dxm+fTMGynxYPoE9zGsWNEzeZOcNueMzq1OYsvGytVw
f/MqtnFLX9/1pDUkWgvLLq0p+4TTSxqQW7hFc0AYq+KI24u+H2SSeFSVpZia1FY3/LG+ywMndp6u
xJ9NTBc9JIUTaPKRx746LN+cYhoGp2ZON0xb6cj1IC2t1zFwfuu6wGGbiH2BF+Qjaf66021kjS3D
mpso6M3pTnH4eGzIXVrxOCNn/gOvxPGFFBjquIhfp7ddAHK5arL6dZY8TSj2/yfPThcBDe/kYvMR
+b6wUZGM2hXhMbuqmqkSBt7/EinVQH3NdOBepNqCsWuYsxKw195s5mnvfpKvGDeg0nUdDQYD1qVU
Mm+lmfN1+E9ax2SXXu2jk3fkQlxcB6PpdaNdjWlKKzCZ+ZjwjKz8j2Eq5jWnNj85zD6+Hm0B/XF2
7PbttqhJN97CiKUtsj4DWqJm76iObzBQ8Tls281SkJxi8osNvNR+kLURQyyxYXBZLCG/82dClwKw
OgzAh5qcijLFI1Cn071LdAd0rOA8ZlJABDePj8ViRa1/iYea/nRLuMuU0oaKomFFt4ZXJAR7EYo0
rj+pYbrSyq6KAY5iVplbUR2mrvKzz4Z5cO8TGFHBr/YZCxBfk7KMxnkyIqrNUbuSyjZl03cJthdc
wQjC2bzBdJacI3kLGOt2kE7Vfr/7bBNWOAEgIR8deyPZbWA0E6NC7s6k5watuKKYFdGNHKd5dTpo
f4yy23H2Zx5exfOcVifdBsI70NgEHeZxE+CKrdLFNT5uSHLS95GPVS+/DyZ45FadiOcnFbB+LBIP
rFUsLhgkvfX574YNx8UGg90bRbJj9xTLRm1WrQ9q1+1fGPSiP8NLJC8pSD7GJcOSlR/HPPPj3OY0
taFzcO1mXTwV9HmcEcjaaD+ujt2ac8x8EuszDcLdlSYyXVadMwONkX/DL6vedRRNwu9w0IE1+V4u
48oOltS4cpvd7GkBt4GCtdLr9767CV15k6SLRlQfpf9UXXY2pUWjfWtoK+nR2996v99tx9S8xh7P
YDbQlgI7djm7U3Bc6u/6Uvdohn65t1v782bJ2pCpBF8/7iuneewgDOT7kO+YjzBtEcEaElEOO6C3
JPKjIIGZnRc1tK26QvkJMnlihQCOoRG1bqaBgMv1yejl/AmBUMFqBee3Zm9K3xxUC1Icd5jlFVi6
01LGBM6/36w+CC/8qOZXMWsZ5qTGc9pUsB8om0lyGxtQD11A+kjBIe1f1TwIDZa9N/G8PQ+F0AyR
c0b1VI/dsHxNb5ADUbMxadJHbBUenizJP67ne16yVufj9oYfRZuCojXMO5sE07Bt3VAdtplAi+WI
oQ9ECs4t/833aQ51D92Tks3M1owKQ1yQaVKJZzvL6gSp9m7QHdWmEkQhlhOy+mY7d0qoIo6xRynw
QE+bt5yJqnBNNAWcCQSthhT0jhFWKYGt7KK77ApRVUitoc1w4MF1slBJ4YL/bxPp+BtjCy8k/ARk
EOJjLDPcDGl0U6pR0vJOKl2fCND1X7EP6YIZKXcyiliyJxbq+AE3zqOyKShnIvyaJhAX+DVlxgGL
1xmq74/VJY58H3+oGPFqXGC2tG8kqHWJE6EvNf3AMvTA8YwOnAuTduqiALrbx8ogPWwisp2syBsP
X7PU/VzSUM//9YURkH07d5L2nemiXm5ULzBuBmjDgenamsXSiS2hRwVoJPurAjlMmo3PlixCHOKg
qAZdFWyAuaMV89hToJQJCfkBoTcstwfyHrwKHlmb64YYDIElYks55RDD0dWE5YNUndbXT/dhJlpi
9XRrkvjlSgO0O0hm1L3ejNMeNmhe0QxcXsnJfqjglnpbzBhT6I3E6GTZpytridA8JF1GyAs7BwQ2
sHSVnEzZAMKDbG9yQJczKCRVkFVhmEKGZxjUocsh3ZUNfQtntLzPwkUsQFZmY2HdWDHsB13J27vu
/lta1YoceADptYATrNL1lfe9nYwAeYOk9RAILNOHAsj04r68jvTK4ZnZHA+0Fj+KyN0cqJU3FORM
0VYsFtqajCd7NA6lI4KneGYRqmLc3aTeTM8SI7DRBG0fxJ9EJR1IqJ5dJB6f91h+/KhNTFUbPy1F
d9mR6xtx+Ek1qsSpP3y5CgkenoFXT488kFCMLARtykLuza0DKtSTsJfSg7Enssr9YgEj0E0c+LX9
gSBepBQrobS+vmN3MWwtLif1bsfXn96AakxlGCsoGOSSUSqx5ahIv/UJQ6mCsogTBUwUEW3PNPAF
8Vrx2EbIfm47M7WcJh2442baMQoWZMWq1pMv3ObDTQf//AFy2E+KWYXmpBB5RY0SdD4CUR4qJN0x
bJCtFBVcfWqq2XoWDfGx91MhNrjDukJh1yjS/DZs+hYH6yWVgtwY6/G4zLxyyCQiX/jKYCUZDrJ2
7VfzoUa7RY8c0N+qR19qb/t75Pf1cBdrNN+ssyKdCXH+wXcFSwAVt3hs3XtceWVdBuTDuBhD4DVR
fDobRUMuRh6xAc3kSBJY9Y42v+cmXuswH3SsH4uHZjwf3273ZjZAicQ68uHv3MptB4b4pYFJwTpv
mznJYNnQTYTpu35ssmLU/UivYKRk3PSNyJchQhQpYI7DGB5w3MDWKCgxv9oSc4DkGTqMboqm8N4C
Gz+37mzdF1n3GY3TuDlO2+0wtbEejsocmdj5O5EnRwcBernlp4A3dO1CiOn8Sd7zx+nSN+DBfjgs
MF9f0oSUqQ71ihXAga0WgX/Jij1xN8OpijXGl6Qjwlee9C1DHk/WJi/MUXO3SQjQmqrJX+PmmLXA
+BkHDGU345NoSmaabW0YNU2/IAoMYdK+bkr7wwlhNkhdyD3mf1ZhIXWXKxbMeiW/6es/3bn/C1ja
208OUq2GV4iNKDq53yHw8NsRmyI96NU03aXQkRFR07uu/WRw20nicN/YaNWbTnPheMpfyt4q9D7H
WqUi26b65Y0RGQap3puiYLDCCbIpf+uhkbK4Rh60ENE4/sJFzU4CuerOLUSCCtfnsNX4futsKThN
/SbBah7xvIk8VIDdDIXTJ2gt9c7mh5446T8ezkQVqdLEmjc/eSnqeEj7ZT0lkPAVFT0LWceHDuPV
qks90LDso2PbIkv9RoI1ywTwKRLRvNUtEKGG/vlbTNgomYlAT6BeU0kqZJ9J2atCMR2eRSdLDl6a
aCkJQU0BrnOSBY95fvTsLIdPk6WXXiT2RZk08ksKl5PtdOzYc/+AZY9TIsv/CT0S2fhWM8/w/6Fm
/Zh0as/YEFJ4k7Tfxso6PJhozNJVXCskT9YZagffGTYL+XEDrNvGhHt8BPh1qQRXwtVTSuc6aaXL
tAUQowzdes2le2DwpRi6IUBCh9aIOniluye8CbSrlUnJcSUFUf4uanS6CnInA/KEGNxAylSBIcAr
DqMsgciFiC0DwYZ6GgoUVkTY58zgEIXeLY8aZyH9QKE1tF0Tv3Zi6sTQj/0oPSHYaWncYIlA5Cmo
9BeLuqGfjfa4M+R7MXUfwoQOAuuiSdILi8t4QrqTFJ0/3MDwwX4ZMIfC9XsDiVlxQNiXKrX6jYsY
KqgGe2m3vx3iylALnhD8Ba+9rDeMUKWp1tWB68SllAsZdbHgtvzG9J3NZIOVfIGuUWoUJ3yKSCUA
J9ZY1/dZkXXKyp8eEPD6/wHDiSgcBBpribTCurEYxYc2jp0qLegJ+hAPlmj1JiQUBlZ163EvQt/8
/WJGZR3pjRcehnz4SCwugcn6p9olgSutk5Tc+WWDGsICeyJtDIHiVOb9pAxh3U6qWxLkiC4qDpXz
DYYayy8OOv5Z5ip9LvKPFRraTua6vmfDY0ANoL/UOTZ2DGdR4xjUwDIQUmSPobYGaScyn0YCO08O
SH2JtwQfGoMfXBy1iFsqiRWAAwmnU7zlbiwdUNspUJHakIObF3v91+g34TkRhSiK0075Ix3E/VcS
GV8nrs35IMjzLPZFGautcn4M3gSCSndHjJ3xED+5U0N5G3XvOzWB4ISlkIsjrHfnhBCkvkTTjlqe
qz6bx0EBrweVUgsv5XvMlFgehPnyruywc2+xmKNdewHtOYqELs2a9CP/9xf7UXI4zpb88x89ThSi
SJrEfV/D2x2FTr9Aa5q1Q36ZZuHoYhqM/sqWPHQM+GjxMlcALFO+lIa1qccd8NoK/EcveQfIdFro
Bb6n7QdHL3Jagfdoxmgc6ciGFfTV8DWrq5nU3fAWYELoa97j/lOwPTU18OIh4fhbPq7Wk5+HSM4+
c+qLAanA2Te6rYY2HsJLFXPL0OOhIUausQYZPWbyN3J/hA0OTaM+LNr3HhwVot6ZlZYNI86C2GRR
4c7EJTSMxobmKpskCC9bj2uwIRYpWLahUab1GbEpdYlI+0zeEP4tVlrr/dvziaddEL3rE/PLTZnk
uNFsn4nqewWUuOeypLSQ8NPlpWAlp8kwde9riOYXf6Zg6ghiKca5GP6a6ZYDWhl4RkgXYITCmCTu
4bNaepAnhNOSiLcQNn91epPnYKPX0q0dEBsdmVmwCwpZLy355ghsbUTMpUQfIi4kaKZ8j47DWkmq
7RpOKvl0GsoYq+ipkOQYQDEZlhP0OwmK3O0TvGq1NWZj32CLZYgKKb+uNfru81XglLeYeF2fisw5
3hKccrIbxqW+GVgwtIt80hlmKpdgg7+N8uGJvwy9YKGzMw4nJUuVfSr9N7GDoVvgIeBty7q2tZsH
ExLYieFpy1FfgPdRkzRW3N3O0hu3r6A/jekGbkyNxsAQGvzZMP4mlvfAKL7gQ0SL+gDNCw5T72lj
miUMUJXz6T2XxBtgENLo++xK2lBCI5Xb3oQouxfjIj0AyYw2qC7IOIFPfArq2+ffczVAtc2p9TVV
7VGWqZV13Dqh1KM+PNZLnMWfKHXo6JuOStNY1FlTlmuamTAJLsT9lu0/HZCFk4z/b9Md0gqv+Z9/
LlLezToYogZAkLe5unMF4xJYJG0fnUp3yC53+zLlUlbmI0zxIamh8hW5y01z3wtnEp7mKeK/wKD1
y1YoZQWJpintkx0TkcQ4lsr4kJUuiwQRSxlB0eXABOXLW/dmDNiwBiXFBwz2Em1nL1TU+ALK0NNl
U8I7vbr7MLNRUaJwbUz9seCXnTWlKFtlS1D/7KBWBvQNgoVCl3+XfcouKohMMftTRFTe8xj7cva2
iWhm1iwHNLUqkJVuCyFhkvd/gWVRhfKhrOXRQSi7rp5kPRP7mZ6Tmtga0irhqji1nlhdhd85YHCF
40ICaqnxDH8Yq/iBThacl3bv2bVh6NlHdLFZXHuXdWAbFvj2WDo1Mr3KLwb90Eh2wQcfKC7NFSiQ
5xDZUxSJ0Emwsb3P7l7dfrFt3jUtt2PqiWWIpNcgaqahBeNJdhuLaaAWuVNFOAN1WkJ/5TeZYnJ4
rZCMheZRgXyHp6x2Cqju8zOAyV2L7J+/8WXQ66VPnTkDKINfhpCU70JoRp6WtGp4b9U/fEjnwJOO
wTmCqdqDd/atiFY+rnTpK7KLCbfOs5pGbCmgRstp36AKCrsT9HKFO+PsEcDS3nAXbpWjsqMrSujX
11k1yg8uA1Agp/L6i9pWxg/re8vYhftdceEEArjZe0CgaWuYxU8gnMaw6rdIClqmfWWCKbHZY/Yj
zbnlcdZ1B38VfbjYI3hOv9jVQ19OntFd+WmcTdgcr7h+8KxGaJqkfX8vaaVn+aMO7QUs4tWHjjxi
o1CDa2vsjSt9hRYdDvNQpdx6x9eB5wg8TGEiwYLFigfiYlgHwHWZhqomJrH2pM7OhqDUAmuZGRt1
mAX1XGDfUkafKGH2Y+KUZSkKJjyvJvOjEUzG9gzQWX5o2RaHgJaBtdfzZlft++adyBJVXD9ZwaU6
PxYRejFWrqnPfypc50MW6vuhpmha8aOEkAHmSEB/GoZlIIIiMK0as6KV8o5o1yoeNr36QtcQcVnR
IItqeXw6fkDGyGQ5cEwa8O16LVtl7vdbwhpZbRTwfa3XdkzFdSNjdCvZYdrPbmlt9rwg++gwmcKL
tOc5mKyZDJi5f0anNSq2aehrItsdx+jB+ukDM7ngj2DOl2lXipD6YbR7MsyqSze4KVhabrlY3pOu
YGrmmGdehEQJK/IQooZp4LhiLFZL4GR2OJ3lZZ5CmOyBqCqf2DRToDj3yEvYme7UNCIz0lCSek85
1d1pfbBySvrHx/RxUzqes/LV17nEJTToArjGhuu19PufzPcV+mFwo4QlXBqNCHQs0aX5ML1/ZW0h
vEDU73GH5AdPpRy4t0ZkJjBJ70DabnvmjEMVSQvbv8qFnOrESqNmlI+KNmFLRF/jkh0Gv2DYtWax
9EK7MKoCsJDsuVJhIw4ZPzYe1WwEYGPftrFsbuPgCGnqCP+QkoM4HeRlWDkiqd0NzA2k7IUV7Xr1
Ti6tumH4G42uHbKgFZ6ZEjIJtgVYsrVm4+J9h5qLC5O2u2C4HnxXyDFT2jan+MskDL/LzKFkYyXA
i4pOEckwgxHMO8/7TbjxLtEH+t+e28YrWkcQp4R1UsPcPMdXHy25KGq1ZeYYnVPWvO6czPKWVrfo
6nhF60nS84I0MZGXKMMulNWK00vvQxsDt41x9wa5/BwzX+lopx35LKuG4ro5oHO96eBrHC4w25XZ
z5pI78VRrr6B7ZoBkp8YfaDUEhcM88vgOBvEbIwTLBfBtqXyVXmz42sgpeeGW0l6Iac+2xak/gcm
XNhUglfQstSEYB074K1KBoLDxvb2p+gWiW68ONrxiQtHPGYywFyWn3zglHS7ZB3g4ZZ+MHnemPJU
9lsjCJ0lmp6wSJJkEa0YWvSKz1THD7tutSahJLdWUGjpnhwqhoI4Hndt93v8cl23Hu5RUbOwKxnq
RwokCOdYmhNUpmloSPwhyQ6NKO2ap6d0kiNBZ4ulRl4brGekwYk60KLZbw13MZj3PV/G4PYYw+CL
ITNfYHWYslfR2Y+1y9dsxsayC+WtV9E+dd/Ps5IlkqdsM3Hksv736ZaE4Ncf9PzrbxmBytWskBEX
dYeD+7VR/DTh0O8V7FtNkebJknGTYLfpZ0NKHrgWqz9tM0ksBkM80vyM/eFeCvl6hkbovSBIPBsS
8jvdWKnv9ciFkbJp7/EmZupCdRanFtL+KF222zj9FONDdo/AClgfwfmqEEZ/kNeKtWXsXM+y8Q3r
+BjZMvQg/IU01BYJQq7gls0Yu/6TkSr7KZDERL7bLJaYeIuYI5TmQgWiZLyFDHUg6kGVwABUh9yV
TCdlDoOZst0+byklF0fWBA4weX6UFuTDxeUWyzKGWMjpmFYuJbjlvY3yRL8oDV7Rf7zst7fFYLDO
a3IDpw8nfOfLmLTehG7miSWdoUGIFDKngdmZfqR78Balmx2esMHakVjUgXW2rT69feqoZ8tb9YyV
BhyVy9DaWWwHmLIzquGGy/MLCsxIfnFi8rKkznbjBRgA3w8kpW8dN3Qd8XP0fWR7NOhkzaKRkG4S
sOar1+BW+O6TJzW4TR6KQ0DDn0rSEddYgM9P27oyjzKIk5D7MU9IwY91V7Xg0U+gyIUyDAVesH7q
PPhqvP2QgVD9cwX9VHZm57WZ0ivjCS1Ip7A3N7Ztk9oRQ0l3GWRW731y2DZfNJbCnTG5SM0GukaU
6+GVCMBvM07mR97F8cySHe/juo1MMYOOfilJ9YtEPBWC/2fBch7UrFMsIOXZmk1S3rpgUgmHWel9
xDLQmG6C/GdYbyG0mv+iGV524XbTR+rEPJ9Tcq4fDPge4x85zRTupWs4g0l3wLTsL5wx3pcvExZq
H0YGDlpK+Y+SkZnLBatoBaFkFGC2fJpWf0T0yMwhJhJrQv5cLoFtSmIs/F4+3O1f+ioCokXJpuQu
YeYrYDmAWmrAEUd7NlePMdjjgnEFbs8cgAYIoPqBRk2THiXgFtR4YW5t4tvjp5+mB0xJRCj7Cpud
OQPAPu0wE/c7JxumcOd8FmcZqNfhdUiaQ9AQu/LXkqpD/KvblKQyytWmr3gezhv9MhEKNUaVgQkj
RhzNCvnWgWf89egFzBeCG0qgzu9yG+wnvbKxZKNnlhe+vfeH9/Fe4eIUGHfYxf3wV5tlMx3/T6vE
fbXMEYHagSSTckIslY3uiJpDjqWplmOFFCdRz115F3Q90yh0C3TDYgpGjXB3p6TZPSFY3Gg0AINH
57I8Im/vqMRotkCUvweJDs/hw3F3CEdinYNzsR+HUgix8GCx0NnyHto9tih9C8CpLXsTUeav4oa0
YNKq7Yd00Xk/b5udv72TPsinh41YmiZk5kCUaXOl4G5BhPtjQXW6kaJvHDY+MI4gd47/owL8wXzt
pnTyoQdMWg7IsRdVMswxNZul+0j+IMyJxVu+9i+GjYo5dHPD8QPm/P5SMQ4MoHR0iIF9b4GwJffY
RMPmN8/pncRKGe9GymZZrU5/iTqynT4ZbTI/w4vzvpQzisgJisJm/7Um4NDZqmRLE8FdeAl+az2F
aV5Oy/o6jLdOFE/rdwPYHod8SfWDkLBQH75tXONBWoQmpW9j920RzmyGsbto9t7wrzKLzut2YrCt
1JgkjuXIWyHKQ/6f2aFt1njW31UiUj8JxxjFQjkuSekNoEYUZJCYMaOnk8+7WpvSmI3qtOgTRYAq
maiPE0VyMIUmnNEcE3ZNJqXoxEdKoNZsYMWRLKgSiJ6R7Dg3JZuR/ofDenSV5Mf/cQ882VQl9o29
w+kdh5GBweth7WgcmSiywxVmF4hn2s+/Itb/6VpEDAyHFGxfBd4Y6TOMNZ3yaRsb9r4BJSR+qYP4
JZ4cPert52Bjk197IrCTFntjQx8iD54M9P85ffgOqWkLbcTbs23x66TAJ+GO/1H1KXgZfhxfeT4j
7QQG9Q1ORw1AbAaRTd/jGa/+ODzQbOi/02WZvvDKDbW03lo8UWhvXy3wvVCZP8dv1zc+pPQhoCmQ
Xu1V7P7x8UDcZr0L9MAoBcgS+YSFtpwjZ3FZasm11hwwbVpv5VVIZzZBrBJJ2M1PgSr+CfVa5B21
YRWvEfl1sn4cXNg8/eA3LcGPadddpJ/UbGyWBAtt/mw1g0lcv0oqegeMah1NiXww/IFpEOfEbmqD
DAzyuo8skgqcmBMNZdm1yHDWhQp70lVux705BNK7pr56x24bakeX9L2V1fWRshB7bIf+kNM4onPW
vLOp5G8zenfLt07CC02r69iFUZZfwF7Gpm8JbTJ6af2fhj73Q47KBNYMFD8gIEnw0yQTAy/MeOv5
M+IukkfQHlMBaK3MuFbEc7yMDhAWYYx2WuO2GKUv0zYxCWeZ0mYii1xwIZ1AgH+Jw7cnOpeZtcAl
TT7bf7UE4huaey20DDS6WPkJ1Yu9k0aZYlGRT/rxHcj7qw1ENBfXHpIqAWywH9zRVnPNjq4ATvcR
TyfSNbvAkErd0KE1EQ62HCQhSli7AfznpVO9vCK0rtJ+51/1OuMw6sDGWGlY8hqwgeAa4Spquwdg
YajMHdEq6xEVgFRhKzPqU+fGPYXBEQ1UZDJCeHnOxxMtxXz8KwEw+R4kPRUOKLin/Rr/5FIxEapD
2Axxfx2DnRajrxBkB6w/oH2jnVsMeGNEjWE77aSZu5IkfpEuexiOqF7Wl2jt+XpUBWKSYkVwI1C/
2lfsrKnqMXLZqnT73xgV9BKT+9Ay7UOgggXqj/OXNY5sScr+jY+cf7acgTST+V9BQF5FeH3iYFF4
OkmfhEmnWV+JYo+Ve3ulc4JE9ZI3yTjSf4D5qNzHOGmX/fosArX+o8fSZtCKQrSUXbe6gQajiF7m
rOY16/JXavTVmU60xwzd0ofSequQ5ibc8s+4F7MT0qX9Kr2p03W8A899dfFyarLKg9sB3Ghfah2Y
ljPwvOhQDKP90kP//+EpXqa6QJc3izF45aiOFEPTJFgmE3cVTg6/8aDMb2sSD9GWL4BUUvzKgoMO
NfYcmgU0/SXB+thlnDzOE9/i6Liq+pJjvHT17Fnm2I6155BUtQB+hCu/iWYefe/5FPgnS9AiHsIH
C0Z7BlQOne/d8w46hggamSAci08LLLJ8vrtY47V1H6XROfPu3Nb6Zod6rfJkiSIO8cSsGjYlfvjU
mDX+xhYNmbT64j64irZyDjxhwU1/lFCIqe5P5EmEneYnD8VxhhU+iNGxsAkNxb3jL6UVCLj0izoa
TKu/EQJWGvu4lk7glt5XxiHht6F8T78GjKDsoBbM8NvzsCo+vsJ7wXmGLAu/rMn+USpG+sY65Mdw
cRjP+lI3QAFBxFLyQBBp0ENH5zvZ3lv/RNOepv3JvhqR6B4N55IUAvLqbpDQbZ2hv63tiBDL1Hn4
lJD4H0ZU3dOKPpTqcHsFMJR/VX6mN+L0kdNAmEPRXCSNNnMt0LitSi5UMjzRjF3GvMHelJuHbyYr
QG0sbiLz5oG2WOdSMdyg5fPNNbSlb+KNheujEqhN87vGouuW2WEhRdZrEb8oK5qzeLqB+Jwrl1iw
73gS7nMAWSfok5QtIhUH8uaW4c3EMcqs9PxY73xo1MVt7ds74166TgAsijqgQBpZNr4JHXDdumrt
zFd98NRA64lShhWPFmF+bxsg8N4S8mqI1E/lK/iJdPM/QS+hxXiFAirCESFB1EwVOaZK3k/jz+Z7
oGwWK+8tqoAEeurU0siIVSZrDy1zOe/4zPwwq8ZIIdowaE+nMtfPJBEkUVdacR4V2uf7Vj90gfG0
cX5vp5XFVVBe4HLtQW7DtThkvI6rPUwFJtjqwiyfIZYJ5OsUZx59s8LbFSJJTNkogdCtTRcIcefB
hfAYuPiVhHKSKrY+zU9xg88He49JPhbUj2Se5541+JRS7oImUBmOldfE3alyxYIASErWJ8muHRsD
NgAaQJq5LQFBeYqBD1vhBRXtKtFzyLuk+0tUqS0NgYuxUjeE53+6FCBrpIGxsNsnTSJX9NBMxLWC
fUmQn3Bbz6YdeC9owan6ZzGmSkPGf4EH2BVPdcGnzJuctSlo19NCPBSlPH70pi+HSzQzP2JLsJDU
xQmKGNRN+obR7D4r3d7TvN9MLHGmUonjHcOkxSPNxbTyxVKuPZ7oPKoSPazFPzR8z3e6F5QhnxOB
WuBKe0p4Ia8B6P8FnsEJnBRCsQMFXj5lNOe8ewNjacR3oKuIUKDiHmmOu8H2GPr382/HQiJGrDxr
GMFqbTjVCB9hEuqiH1NsS1rDsO7A4+n8uAso97BOp2iqVw5pycSoPg3m/Eet7wonWDwtJhAKlJkZ
rOhVLG7QS4EtLWK4ntuvat2rfTxKfF3+iqAZISZowkXTnL5bPlos1dJL0llkkSMlAKp9wMZArX3M
wuIWmLJxeOdZd+k37eFmFEWmXK3no8v568veDWfbxHufVeNTaqK8JK+ROwIjEVUKbrzq+A7bPwO7
1uAaZSezOsyBiJMoglDOwFyu8Wd/02GxVOl6hf3Lw5AOiFccz81IJdK35NSV4n1Xw45o63wsIW/+
U6az+WaVGcr+ActTGfNJdWVuIjlhtg0oqy7IK/CkzY6FmI9Qy2JaZH0G1KRn8PUomxIZ/rJptDGC
rxyK2MQYJnn/E7KaPZe89mdzKPvb8tSuDZbYkekanG+eFpLiZnIicdN9ks3QYyIZo7vnaBp+YYz5
sKY9CJRF6pP4qFtestMK9cRRk0vTZuHOQOSBLB5U+pUKtbkl5i9BNFytHQ9c8pnaZhEiHeqLxjmQ
OLAb3TY7t+mVeG8UfveCHyph4ktkqOlJ/mf7hcXPSAVLlG9I9tV5Zr0lgJQ6+49bx3qCFQPcKkHB
y1qXGApKEErJeRoYnsG7DKHsA9C+4HtK5f50SAkMMHnUxryjwljMoCQa47LuAIysKb7FiRoqwqxO
Dcc1A6lEofB2yjpTlkXyyv1sheZhATgmAXseEvQ4s556wBBvGZGSjTd6gSoPOPXFLyGMwBG7KslW
MQZV4lBFBZ8pBq/bzlXZ6SP5nlcXKGowjAxChN7K/KO7T5TZ7psq6ahECOPs0IpMPjZuQmau0fx4
U9iCODg1soaDwjKaVP3LGKSjEx3b1TdifJsCLosojUrBVmcH9JwK8Ks9pG6R4ginS287LkV/QpuE
KhIkmW2wMn+UOaFszhT+yAErQc29PsKMUfn6AukOEwsDzY3UzC3Drh0rsyjCtH3fpH8qNBvTmLky
x6ERpvcZLK65WcBnMd/uLXMM1K5c5l/KVrTyZziOeHzTOzg1NYRdQt6HI8M4Su9qM8C1SL2/9IKF
8njSOaUwgzyYFI25r2MYqSaxLSir1tM4nReuu6/OHKJ/BDEfaeC3n+Y6Ugf8mTiPGeqK6HV1v8P+
I0ErJDLHedof0QRgVedQINRQTMcK3sm0eP47Q/PH6COt2kaVqds2Gl4ADErT6knw7gTF/rWhj3C+
cEAmg+88OujD8X47LpuKed85+uIXqx7Ea1E+z6uZgO/GCR26+5WFNBO7/1Yi2lXz+DM6F8NwraRc
eCKmqiPaSbnS+8VfG2RIFYu87uBreTe7Yv5XBJVkYNFUs1XfCkHkj48NZUqiO0z6VWiLwAAAF2M5
4suG79PyM6rURxUC9EcOmiF6LYOXk0PCyt9afc7C8iUNZmjxdzY0TZChQNWDoTG3G9afK+DjpRE1
E6nzd4/jepwGrVwVOzhOPaLYHwMm16dTU9zhoY4cJSV9EYvO9vom+7t7bO46vinPoV9UtvOLHZXJ
xovs6tUbP85Y+QML9HCQ9d0KIXRnW7QyGzPwMOVM54XumBIRYmLypMy3EsVfjcJaWU+y0lN4Jpts
ckoejE7iDKw79riVbWMQ7vTYcip5SwSczgxRuRK+tr2ZAakJx6+wOvKEXBcmJrtJCrlYcb0TOa2N
va55lR4ipu0Whq0SgpJorocmEtOP6YHxgMKzLq6vfr3mWvef94bvac1eeJMOHp/7kUocZNUX2NQb
kwVMiHn5k9haDK6q7cQOaxl6NuGQPykBsCbhKNAkkGsdVr85dt74d10dLJlxtWhCJrQwDDxvrKlP
L+LH06lB0dXxGnotP6BMgzjQGVPBlznq11Jpt9LPhbvn7LZdFB341S1LVtngQU64BxkUJaTOsmme
QSTku/hoa9Uwhnw9qXxYPMCc1XNDh42wS2Tz2p0fDf0flLY+VQXubawlFYrhA8qyn3FlYCMvIqXd
AyADQ0C5eBmnqbvAfBsWS+OyPpBFNz48yqscQi4oG5roURL/L1Deg2xT3Bct6pw+/RBAEblrZ6bZ
XyrOxFC39eRGmnNPxfKe7LTt46kcmi/1OBWIfGzWNizfUcPVfSNSg9XpgMfMXupAyPbdzpcIj9lK
1gxdUJbp7/2BZTFjKILhUqUCZO0Ab/ioGYspnOAfiQHJ767KcMic+N7zhg6wyTIYYecSd2OZTLWZ
q+PLYcZkw53Okv58kd8MfjghjX4BudXh2EQ1BYcVGZ3gfQLYobGIjd6cFu91EBQs06Z8F543EB3l
kNoXgl6FYr7xu5485GXRZDZjT9PMnf7mnCoA64seo8O2u5UB/Y6WKK5csFh1tWAs82YjXklMppc2
woVVrXDXVtQ3PrQg8hey7f9p3QWimLD44Ux3ogo3OZn/8dpkIMeq7LQF7lr9kkfaQ48NUKe0776J
/05A15iJ1MG9OCtvoVbhVgyIxCvH2GmYsbk9TOPoNMbsClDkqudf7SRTjudfJHwEjElvsWHo6ITv
crmGIshqlp71oZbCZVclxDA7+fxhjBG4rVQBBGVl3GgHS6ZQ8a9kr+IHPWTWdK7J5hQ3YfBQTOND
76VyrgzjkEdVkkzVzd7GHKKjoDTdna9hSR7EaxnOUzg5CNBNOmwbCWAfKsSEbMu6B8I7YWMp0kXX
2zaWAm3Xzo7FMwiHMSibZbxR4ZbD3OmteP2uLnFAyarVYs9l/aLm/ni2YSVNpPYnxj0+B0Or1D0A
yTfRvJuviziSMTaSAjDPzGYY9Wf9SVF1TUKESPcMCHf/QBqrxx2MmXfJ8OInYz9hcg6CXCuihSvk
pCImIddotT26wiRphjPiBIz7AoCxf01Eob4De+hz6U13JLbQKCngvtLUUq3C3WDRdEjjsDGsmmmP
1/HzdbXr8dgbFqt4KoucmkQAHowGSCu0u9pyNvtV+R8RMAYyNHbXKLg5lxPHdY/7GUrYcmjS+nka
R7xs5ZPemAavwt4IxR6zILkyMMcIq9+cn4Yo5EOHScnjtif4EbdAq46rTTCYlD9EZpCvUoK18IKM
Hh1xkCrjnBsIFqlJYPRXxZ5xE3k5ZfAhsXqE/F++Z8c+uQxT5XrDFQ2dDMPu7jx/D0TGofVuRzvr
ZcSW6rtjeHjHesA/kv17+7uh3hivORPODRBvNpbe2DJh6DRLLqGPD2Jyg5EMURyixVqW0g4cQNIl
xnzrnFCvr1iI4y532khLaruIJRGyheGVvb0gCKXWHjqU2WZ66cY4JJtKM0iQ+lPvA5HipLxTXtP9
9tfXIucCFU/5RzedCG96YtTZEWD4boioMFDpLY+8MfVQEde+x6j9IHVJD7aFU2ebQJanDJCquGvy
2OSH6pP3YbN0paEfvT2e1MVqe3I9uCuJuaLsVmibWgLxzLQF5GAOtF76ybX0+VQzw7WpQAvYoQFk
mAAYf9/pJT9wS7V1WCkhiHi31X5LBYuSvNOR5qAW7Y1leP8OeljGXZD/ojs1+C/aXf8czXJTtohj
6/ekQoDjs7xPxKPJ8nefpc1t/TEX6giGvNIvgvZn49s5gUaH5ARitcZylK26D3AWSLw+egVp475D
WZt4OvYq11u7fdxcBvTjfVIcVbeao4OgmBrYhh+ZJbwGPptVnP5Q4b19rSc8wBA6O7hYKXy+mtZJ
jaopumUu8YTuPvnBxYxss4Z3UJ2QBn+4iuWaHDAYAbIBUh/ksXrcvtDUjeC02scj61OZ7UQY+A2Y
gxxvWJNYbN3VMfdnlbsfzTfcCH0Suo4pOwYjVzhrr/exjBqRpKRU3+qknI6ifhC2Yh6b8GTLagSe
kWq4Nyqp79NvSD0Wdswh7pBk+U7orJRJ3aIUrMlCDvaX6T7hcxt2T6+HwsflLC5RNF2wHC6lnRRI
u6bC1gpMoLNLHe/QSht8aCUU3bXKALWul2B7UwU6sBw4zx6yuTpwmk0hRWn0BsR0szJEL9SOWqfK
tVepAMZUSOmkNG0Mjyvj732LDeVQ4mlL6ADp83HS7tPfItZUnIADMjJkzznPFIRyHdyKN89PXITX
2NgAgLs36Q/7xHJLBH6Uapb/2dDaUugbLRlbjQsz7ulqflJfd5nUVIgvxM3nGvfbbd8uvn69jT1M
cigHTQST/iCr/2KKu1Sp5o2Z2ma/c4xRTVMIQ8wQaUFDwwUrKy3OF0+dK4A+amTmEkIhDalWFPqG
wnXSIvdfVMy62Pot0oE+lYea8q/tttzpqjSd1qdVSeeE04LXhi2BMjdOBAPBKVNohF9l+9O4Loa7
DJxAGSAaJ30BuSr+VyqPdSHaJS7K/isLXdLwtzUVBlnPziZ0eEEa6SmcKrL0uilb5aw/QEcVHlop
BwvxwRPtJ5EJZM5olwCh+HGZBxZXSL7ta7rA8e0tTf4238HrbCQNIl25Dt4HwSz/D6b15kzbGrFR
UTNA3jkn980AzPtoidMxE6SAVmVCkhaXXyE4OVPPFskzgfgFrxbmcvPbJLJ4jyXreo0p3QbOUdLl
GbprHpOhIfWjRIbf80Ql3vE3RM1XXKXF7WNFhb//CHm+gKiwZmUl10L/qCwbL2dKGuRJvDWqvS0t
P5xK/LLmTZKYIOuiHtyi4kcABLBdjo8gzr1ihBQNhD0X0vwOQroxtio9VlJAgBmtatqDCMVGKpp0
0EJXEepJFQfQWQIQx1y8VOxrLgX3VUVi/0sg+ptbHSJnVTF0tovEs50rBz9t6StJJdn2x4o3jW3I
x+d0Yuc7WIK5JUrQIKd6FkkjRujAP/sjnQLvdcIX+Ougg07lJ2C5gcJD7dzka5/LboUmg+uiVTC3
ItRI6BYlhmCJdE3Ptgt+B09g7Lcbp3GTeqI0XFHIMm/etJr/0LUwF6wvAbIUWGmaQdc9ocVedmLO
jCXMf2SDhnKi1B4ta+RY22YFlPqu+YQi5lIqdhyvZXRqPozQ3yl2mb5KSLlId0HCNuiBqFtsD+fB
W4s5T+YiAx8ZgDgIwmxEBWHc0bUymf+l+2nn3h+Pd8ySO2y2EK592jYybESBLHEPaxAFWRY6NTI9
W4AHAPq987DrXWuXoPxnemQU8NNt1A0mw+qwaCO1C3SKBKAIKyaXZFCz+hxyUqvx2mqF2yTElMWq
6Kx+GICyxB+b7bJn+BNKJNMxQeESZb6BhNE1EZP89aobW6Pr/wGI3dtBOSr29Fmrczju8SePCjwJ
vViYuMRBIqsr3HheWxYVreYpAMl6s0zgKJhsVY9GZxhowDbA8RnzhELTzZBYVmfzcDxd+Dnuec/H
TRdX/cVcRMQ5aclWgVtWqX23BxNyVyfweeAfNYAR7CgYwLGNVFqaxER9DOMgvPqVuBhXPel/m+0h
ux1+VZd/7eaLLWikTkpDOvX6BUAIXGXFcL2QXgG47g2bxv2PxtLyV1l7iyQMz1MWnYg1qdynuFqe
4n1gXkdn2icoKiR4MR+dRzUjZr6+pVOOkLMe4QxuRyWn+rT2jdhISDy/fIqeLpsbC56XsS5I7bWI
Q/+BD0jLLizwH0nH6amVDvdiBB6E+2+IbTSoZe0oc3Y13jG0qMAbNl9pyjdsfvZHfV4MpVsSI9JY
4TNVwTmJXsWgwBmlxumajAKbfA4EchWfTJfx9wOD6+dnn6KtyCfb+R3tEoIyZZTasU8wjOgow/nd
UdqC2FolpBjzJdhw2HznW0RRs+H4PwtrStPqYA7YU8IS+L09zQTRRVWGSsBKT0Fw0D4mga8OiQsb
UUjtY1HNhu2ZdJu6XfKhu7CKfHI4Aq3+67fPV4fQzwP3oGwlvHu+SKHym8A9TE9mgfvStC6rIUSo
h8dGk9HQHhtcy14dZ6Vyclde9QMi8yZByCqHylPyPycgLiE9n2jxEh4kYNue6XH0zwR9/yX8Up2X
GAbvpl29sN3lYMYSyvzuUQ1nAcKXONRIO7yoU8ceHGpeV8A9G9RwXVsm+ohR456gk2UEQ7jmqz9S
qhCoEnuZU+u0KUG/ff6Ksl1mvcyqCHuM3kuqsll7mh4+xzFIePkBRtkiKBwUu67Et+Dnjn98Ag8l
Y499b4bvcQZoYe912Z0ZSGmURRZFHGv8F3aVBR1DPMWlBciudrVjoclOW2Rzs4pzBVBObsr+T3WT
GRt1PGA1YKTyVQ2HMF8x2LsvNOmXQ+wE5gliLLhnyknlwTwkmFTOiDJpR5rnxrfh1mNaODLGTofE
6bEbHYTsNYxwR9HeJ6cQommdM7mezOAqgjrR6C/NOPqhmy46Pa9gAIG+XSo/O5egYL/0zBG11bAL
bmOeVsX+6zetdOuWIeI/gC2k9mZtu8bUb9myh58Sf56uzcKaHutshvgauM09xHI72odHK5Wmer41
iXMCc/iuKNe9iT31x2LqKMDDlgOmL/UQ6rkVsqPG/O7W6oAHnDYQM/TEGySeiwAEKFGTJNxw9f6D
nwf0LpEw2YIsipaeY6pTMV/hh2GJgY9mXD/ldWiaYjVErIbaqsiQNvpg1Z6N9ngiFPHJqhSP5VNv
XV3NtvyIxcguyfcee4yOwgWdTXq+S2bVNeQmg7X7zmfFxVXqOJWKOD/JxVN80yVyB0lJvwq5XFaF
evJcIEgCrITFhb2KcIWOZ6jN0NEyI+JxsgKI560ztaABrwi9Q4PAnPYOjWmob7LKHzn6DhcVEpgD
cYsoVd/Hy006R8PFtWpvmUo0W8J/iD05NaTzh1P74SEXsRpYpKb7GB5TaY3o9j6YjqH9KNBxAAUu
bBpU9g5ctaRYbVrzNrxg6n+w318btOFtsb+4uVhODUs0kM6/wRF2HSsEx9pQSG6Sa2A6800EURQv
NzbzzyGbdmf9R291WP5Y2LP7Rxuwi1DK0On327OGDnPccJIUN/IzV/jDz8JXTNarXOTTeFk11NuP
3Z/bN/Fyatb+ZGVPHvpuDR846BHAlqtfpW7/BrNZ4d9wO+s3H7i4XMPGENgur522Lba7ZivvAT2b
PBxxokCic/rkhvpPK4RKd4wZcD3nVR37v2NzSwTFj4k9jLy0lOAOkd/oFk9+hMDhM28H36s3lECy
iKEcLv1zDutDj/PiwmhMURV6EVPqZqPEEeH5X2jw4zWc2qydqDuzfhv304DMNSEGdU8dJHFR5Sv0
jRq9sic9BJKy+O3vfoQVFcROR88orllG5YZT3QUKaFDeWnHDmatbKdiwNqAMKkiKzDglUwocz3vd
Z7aj+yWV4Pxs1mkCNRovvUHXSLkzG2mEl5+yj5Ocl0GHprdByCRjbW95jg6m/sAQ/WHv/fLLGkVq
kXhyKPSaV3w1EOgk1Tt1gCLchPRHsYD/bBTg9PrziaoiVdm167ThnNs8FhyhDds5M0nudjFw53RF
FV2a7ZliGupu4AGKQwkXpqlSyJvJXOleKJWupdb6t1GkhfEWsIP6BBRSG+d8X4aSbStcav9JjXY1
cyjtUuw5X+KcCfs1qJ6hInJ6BFYZTd4ME8kUz1Xhey7bcFEbEWBuVLEU14WyIkPODTqG0ltDTmoz
rNP4klh+ZfLDlb8SH6bsqHCdT1eGEa3KaBI7RITnjMNg7C8X0fOUMnsa6hh5b65wsIKW7RqC3qOj
LrWv7/n9DStCcwzKwOdQs59Ewq02HdNf1fXVUXfk21U+3OGKp+qRQKT3B0DOcxJ2tELuUIKJMP6c
Wj/j8w3dVDqecoz/A6Gjjpxr3tD3OVa/cTb4157gtFvDbjdVPHXV0PbLJPzmn7wLUoea1kJQ3m+N
1zqFt3BGdeE4C9iofSBiAV5GvE89JSyWQFSr8Qp/WcPhHXjqXqcMGf3nQkkt2kBySmRtYDVoOcij
BP/tXB426p7h3rtd1UObbCMHLFtXkPDqXBJn20sHoUdmHvWxfqzPsgjLnFDOZM8qHMG0S9hCb8qs
CJiKAfjNcsJ4WkbWUdqxqmgmCtIOqiG2IqZ9tBYnO6s3m9K825RVfuI718McVkziMZF4Nmq5z3pT
NNcOkDdfULNrPmb7RWruncuMaXcKpdqil433SusmJZXs2dluMTOr8SGQIds97f8s8FQ7ijXwDO3T
mRQsoQH9XcFzkrRiFSfch7Rp/b2w2ny+Brw8nEmusY2ZL5HFGiH9YCt8wsc083NOFHlTeiJkX81U
6eq170hziBvoAa64zJS2CCOth9wBGGcbQT3uqxAy1WJ4d0npMPTPdWvpV2Vaay5JMB2t3J8ezsY7
kHW8+ScO6bIReknYL/r0AyRiBPS9DhPUA7abJiEPpvVyABbf19AyaB4+k+OH+7CmSq+nVpF+WYnb
WH7UOYrfgyb/Xd+oebheWvCphlkASq8qWX8WzSfLRlyM2sLJE/1F+egWCON7WmeHRl3o0VdLGPAL
omF098ptRtPcDEpYdKeesShoF0SPj3ig7VfbD/awFvsWWx2YGzK/QNOgBaLNpDlpNM3JB6XuLhMc
1TC7sD+QCuS3xgCu2JxaBGamd2moRe9EPxVuC86D/JTrY5dwoqNdfw7YlEuxAYgzNrnqnkauUgl1
4Zu4K6ekFIDHsP45tzAIzWDSVT6ptJIHFASE2R9QdMulXPlXVQ7s4mhL/RDdyFg418AatObtWzaQ
1awT4LLDAA6WQmh1Bh7PSwPOR/xn1X0TmREvAI239y0np4q+G7TV2qq0BiQb75IAAS2heX08Go96
2XPVbdkYhzCp/47diubNc9f+k4tjprB/FW5M1sL2E1Ua7HuVT9PUg8fKToLo7pUVBEtcE4hCfS07
gwTNiOkTxmFXAoMIpkISzKIbMGyZjxQOdOuIxleJUu/IJ9olsGmAkqGetIzE6tW0eTAP8kcZ2ICy
5SJG+uTZm2euF7LUralk3bHO7SgEgkYtZ7imSRSKilXhR7aky/kGMKpttEsCldH6HRMk3rqur6Lh
Va39JuMWuYHSsFiPuH5AUhK+TqX8ye43W6PfFzV8AY5IfMuGb45w0rkirUkx4hK1yHhdmAEqgdT5
NM0jWrf/EuK15bZs8R7CTHOxLgxyspw7E9By895beiQrK60h3ywNCIUemlnUvNJROq48v/AYa8J/
4LWYIAAJYW7Bsv/l0vrlt8N1zAR1IqpQpAlMYGCpnh3ET56taubGrv7xDV3U5Xk7HCgiON4x6kyF
RKGM9I0hmfEl+HhVZAn0KHQIRZl1tOwKGzX+SMnRcfZ3TSF/LLr+WCfFjnPr15x8CZ3ksp0h9j+d
OPf+JA5Ffc2HGpqwJJGQ5vprzLISp/MXlPGmTHohz71Z0sYX5AWha2Hatr8jvXA+zHStWUENdNUb
BifibtOZgfTkl82FvTGhhhjX+Muhx/mGTedEz8mLp92MDmnJmQYMwxylInzuKCZJ5+HT2Y9hPHRQ
VWyV3z9Q5ChV5FV8k4KQS38MKs1Y0RxC8kzvBCoWOmKJVjUe+63TQJSFGruHx3T9pG/uOVosss79
kmWLyQ1+bk4ulxkPVfpo6J0PXKIlwCT2Cza/J9E4Nb64vFlIIDAS/qeRq5PN6rjPGH0du/cuzGi5
EsNWFobJ1KQRsY8LjQGxgTbkza6ZkWd2P0tbnYHRPxXf9pY6QqbbswH/NSLJb7NzhGueFfTVw75Z
3Ty/DYBGL5ua6bF6j3+IEpLewV9MxNbmz8II9mGF4vZ8RJpSc9Fk4swuw2Q2Lz0oRyOhkMPqwvMS
2HnfJFOOBwpqzV7huyKKU/8i77Awc7qTjHh3jcEi0dvBpxkwGmfvguHfJVUL/icKj+uFrdDzUzWf
nBqsOd/tor3J1Aqhn7T/yDl3f3sGHNBLhf/7hq9nlC+8nfB4//dPJnZfKin0zhanGIxMVx/WliQV
WzkgZKRrSFXr1vFUVc3mRWz3foUKZH6hD+j8P6DP0UFISWMs/BGklpQrjsaWg63JIeqMKCaL2CLM
J9tac7NQTnJPtlCLswFDZOzrv+FW6rYzBiTGLClVatZJsbMQfj+5swKQgWy+vv5j+jknlFpg/+Ey
NKEmUUK4U06enyxcA8P5QCjPKPpD5PCaqZMb3yNdaT1FQo/xjhz2SLfO30ihXxJi9+SyFo17VoHC
Umi/sxE+W+1I+9OfxJGcqnH6Vjy0gt2+QLCkJUQQ5n7iP1Y3UNmCxSnn5AwMAuuU6ysUi/zi0cF/
prUE8ljscdGQzlylaFk5v1i/aGmZfPU3pLV0aRipzq+CJw03WRAJbk0OaEGs5TnFoxYVtDNhe37Y
y7Qf+DhO8cQOV4bT7tkEaGgdwGYUQHu9SsIdBmCAYai4GxJPnNFa7cmsSLrt4hXmC8T1myjAOP8y
RjT/y5ChTy5veJAsbOulsMznzdnS/HYMdWqgRlGk1MXNIv1fePRfAXZ1Ipwko8Ik3OlYPdVBop4l
m+32kedr802ghiBmJK1X12G7Egce8GBfJwZ2zg4u3/YsGqyxO8vJVfqu6UcoQuv4Rs1A+z/PrtgG
jR9jYRVOT6rlxxnQeXzRDB0Fj2auXKo3gHbOnZ/Nkf46q93s2wpw9zQV72yNVC5cUxDScsaNsNsU
H0D9wtIHB5IRRSYjhT/wCh8ro3JMzoTrTRYd5iaYwseC+8iSZ+ibVmGlL22EhwxxqqbbBlQngATA
96m6Rh1XSX+DNF/85o8ldl7qBciu50fK5VoWJzvBdox8ykQ1oZJpnYDoaL0qqI1ilCWuUzg/alOy
7bBm/HaxNjm9owSxmnq0QqQ3fI7z02bYM5bK/IHlQYkUk1so4xmPrU19wKneLh9uXk7DlScWBIr9
PPpLjgQ4BtE6taT9zG35s5Eif358By/uy0uQMrkq/NexAQM7ObPz+gpxdzBwAMLuSO4Xzu9e24X4
hT/yleTMzvNzvmEH8zkTYfBxRQkd7lgr3jPCB39E3iB6CJUGVQ1IMv0U2UzDoRr2VkDpTTYygj4u
4JQgLKkQ/182lBoYJ5yyvnaxsOIvyRG7NVT7QUjjIJ229QNs9g3wQiuUT+OlrRCVF8TACBxPRQmP
FaAP9yY9lVEJSJ9gX7Oo6HwPxEL4E9K4YQgzQXkRG9Tn5u8Xda+nZp5zRisUZKtLfWlvFl+t1pgO
4QiL8lJAIs4rnjNdLlxXOB64XqD7dwSTJn95ufK4Vi1n9IzWmVCUZ5yFMY+7/edYMP2tF+jJ+yW8
Jdq2oOXd/yd/7TMUFNKzmjdGRLt2ZMUZbV6cYltWR44ZcQDFNS27u30uRGJkJIUSNIpOT52qMn3q
nWqfxCHnheTcfuw0Ni68iqiMTkTk4scr5vt4cEg4pZVUXDH7erQIeINakN+p0aDvvPh8bYBl7UfE
tUHWGk1N50vu5XFnspgBIKsam6wF3eqk73QB9HwFDVne/iB/1Cw2A2Yc0JLBRQHHDWWcegWRHX64
cweEEVBuQdfgX1QCkC5Rpw5IBGfjkTvuoNv7hokgxujGf/ZAV7CVzgxu4tr54BTB0oWEekvTcG8E
OhsJKE99Mh8y+1qQSNDB3ogctbpfmybfeLNxgLCRqypSFCkLq6Qefp9uDohsORUar/ggDQCf+zpP
QM/fEPdDFykXEefGRaedVvGhF3jzIvWnDj5a04g3JfHxY8Sivd9ir04/r2QDFN9Wb8cuQinfK0MA
o7Ow8nTfIzs78CbXMEbrGI7BZ3/g5YBs7PQmkQqAs5rsoBSFULORUqiLVDh/ZRS8mUpOzhDVoMHo
ZlhiSh/X7fnNEg4TK5Fr4hy4WZTgYwk4Zy3MVJ04Q9021fuEb4Kz2ZspIK6UnGYXymtbMcvLTR3l
IyDuMnuyrXsAT9ANMaQ44nhAVr8FUsAuX1GiCmA0NOycFbCJsrMVfAobckalpQY5szMlNWtPIOb9
VoaP7Dxp9ZlMD0K7R2tQx3gCoRQxjrEHAsrCFB1/efKc5Z9XqMMLrVA8hK2QRPkDKwdMMO29574b
BWmCgidsNP49xgLeRFbV9e8U3juoaHF7noOZccFfe4nq3N1/cDJ7u1d2U10PIuKn85DgYDExfa7W
KOd3fzC6Q02R+kUpf8Ztbg+rxgoxtLJL4BwkR8l7cwiM5pzyzTvzL6/ZVAsvenRGXEJ7OYtZnFe8
ydMGqWZqrPxaXbupqboOpKb3DbB9UO3Ahkb3gFNO+jLsOLf532gd3q5PdlbdkQwcOCBiQgjhYrAU
RYdcSeJThoeAikHa2LcQ9Qj/8kmk11tGR+fteW0HjQk8p8BI+5YE929wFb+Guz2XkcmzCYkKSOOy
SbSPKPugq+dbieYQVCPhJigeqt3Vct+DrLFX/4fWkPJWKXWm/hbqHo3JjD4tzoB/nX5zLiJJJROX
llTYLpb7YygI9w75QYCh9CPzUCnMDDPyGoALlT3MoIyKNr24e1lh5zILuGJhYmtLVHpoog8kThcy
CFZsi3hC37B+zBCjWgg9Zm+TkqaSOH8sjRKk/2TJpTgxGy+sHEcZEEPpilMCRQsh+lDkRodcgeuN
wjTq2vQ/lmkrLsbbV6lPzvoF0ZEtgEtNTmOjYOO09ekFCh5Zl2W60vpdiV0Ih/of+lYQNHgJFaWV
gleN6yb8uONp0ybSfkEx+wl1MdKqcBVe6pqLQ8qdIyZzdU9pEdjTu0jSU62s7aocbNAEhnu5q8D/
2wnJ/Aqof0Rs1R+w8SCA+QZgcFcvyTxA0sBlXXTuBxux+DVcWWMkM10g0xtKBgkwbErlRDxinG/I
QQxMz6AN/4RxbhRiKVQtzwRsfG7HuluBfh9yC5uZdoaRQdZ06O9khCj3f/2T7FhqLBBssZJKgn0U
Z7Dg/dAmY+Bo+PnUdrn6QcJ1Xest9Ml82TSJJV7FMdD479DTl54x0px+I4rIwyj0LDyydb5tFt5t
EWNZ30YoFqhcWKKPB0cdZFmdfd38ojAzYZK3wSbk6CVH0FQPZ7TgKwH4s966WYXR+ysq4OnXN4Tm
Y+ZDt8d/qMXbav009iG7WeNm9AQSvH5L7/FzjGWaeVSgvDufw/hPgNQiMNjRtaMoc6GG3Dw4isJN
wUzI1pyIPN2cLP+UorDyb0EV12JaGZjnjUMgyIwLLcCfA9y5fKtVSlHph4IQ45quJ/h8hEkzEDKV
GOgRftrr3DUh3Qe2tGfwuCNquwm7uUaNBxgUFF29DodZk49zJYJlZRe1rH72HXJ1KiZTMTbIVBWi
M5c5e99s7HR5NOyBK1XXGeeVAF3r0n7P3LGpisnPTC0Xfjpm+zU0w1mPLWy9CP7MZmYxcoDR+oGu
3PlUM9NZnO/WWTl6EJ0ko3Blweu3thQrte+1/Wn5puQ/V1bstkAFCE5tGP82ut3QgbOlIcl+CHpC
LuIQEoQMEmt19roWiEtcdO4yrt4IV+KH6oVaKALxzOqh5+MuvXhH53ec2wgvBLPOiSBJaid89+Mr
0H/dpuH95d8vpo2KYtQHpxlp8lBT0z/Nrd5t9Rdu7T4lgl83XTXGbRQUPLGoH6DZE8cG7cD3Tv4R
h91sXdGtXWiFylq5hJYOy6QIGhA5OSLyUdZa7/ytq9pQW37NBc28czUPInz5Yu3n5Lbti5Xq3UVu
95lFlbPjqbPzqChJ2vOyQgJTaahBwSI0chKtmkvI5IKmrdYvx+Xyn0n9NQgePxhGlSuOJYA78ba9
3Kc9ipiESZ/q+YFXhEWUQcI4zHvxZ6i6QcVeDAEk8iyy+CciKvwv4sm9tw7dWzUcZCVDzlFACfcB
6cUZAmsL1Am+v+P1cqZleVQ8ATq0nxUPtZnGLDb/dLIzuKg3wOuXRtmMUnbsGAxhhtKQEObTLkxg
ipjPRAq75ueb/hVjIxnoxUSIL3R6nYEqSFI6QC/mXC+vnPKq4U1YRBwO3eCTczWRtuueyMqrbDoV
GDkChob6/TbnCbSeoidVElwXuaBoxVSPFTVaeT7KKxR4qdq+Y2brCchjkblRu694/i+9iWhktc/8
kUL1The0NyYoUxedhyUDFbdYU2upa0DoVHOrb1GwWhDDejHEmDgDXNLiWIeLJ2oh7RpsM2WoQl6w
+Fl5kdCx1TVedRSsBRX2hBixourCTzGydnKzRy6KuShSNIoMSmqoT2rkyS3DQnaoAzPNjea113Eu
Eow/RVtPtCflidMv0qEf/Lw7ZPUV0/6nys7HEBX8sD6GNvC7SUz0JSX5rpqnCxlBcFHsIoZ/MgFI
GtDZGl8Nzh7zQxDCD+vS6walhsc6OcCks4x1UCZgo47Pfa/BY1XGvgGmm34/GbATPT4b921zO0gL
xoHq4tT4Z1NlENjuRFy1hV9Y2gYVnMCqe+ZPxK11LfiJ+2U0nj5A0KnQR2KVs9Vh59r20zyxqc5J
TV85QSDY88EKWwBuNhcWhyowqQGRnzE+Nu47D0Dg6CpBp6N3uSAFhFiOFO8HUImEaPYAGnOddOuj
nvxi5yeOhMe+pD3V4IxhOITCq1sNFf4LPpX+yAsWKHaZespu78kR0ivU4/gzUbaxj2A+GWorJOkZ
UEKAXiFbw4GvV4FiTmQedgp4BhUzhIUWPTxPPryZbpmpWYCTsRB5kPIzdLALrTuY9hwAHvgpfrIk
D3ma1gk6e2EqCt+vT59a1gh//lcKcX4JzupMnFaRa5Y3SOZvHFCc3p2UaUsmbJm15Gfp0abgiU2h
qmk2tqamQb3UPD4T5obV6GFIE3Ei2Ud1+LFhuQU5QDCtfOAHEMyDhpus3y90AwESn1XUGPv73Zf1
1FE+t7YMp4pz5m/61oIJJgoZqb24p8syDt/OFZLlQbDJ8ew3SP6W18viUE3GMhM/z5oYX6oFwz7Q
3BIWB8TjTq+9zNGaOjcACWHj4pPRcMVJdyZYF29/QBTDfuy61mU7Qcj0N8Ivafql4mcJilSYbHSz
PqF1yIYrXQkx0DveGAjwLjNH8e4eTRSfr5viwD7YXO9O9cJd9qkbicKGnAPuyvLsSBzVR6zdDU1y
2j49nf4Y3V+ndHy0wEfpJhLAm0fK5vpD8B/yClr+fF50mLe2JK3HCYwIAn8ETvey+jc0bPOJuNQx
CXb+2CDcR9o05V92lM6fA/gaLGjzdtpztYdu/ryLAwu/nVJa3y9MFv9/AK23Rr6+m9UFK4algSzx
4c0UY1VCWfi57lRA6Hg50NTf0JM8tpMIGCoY+ZGv6sgkYJ0PUhkXDwrctAOw9og6cofVwhSe1es3
Y0NHPsN1nHn9EoT1oOE7LR2SqBDZhuCaF6d+cWMosFnP93yHSUSbMJKC7YdMmGO7AEWUrkEEkmTH
Uz8g/49fSI1Cn5NYf68nfsR3xxcVUt1OZ0C+cxkk7GuzPdRcGOB2qihPwWBrwuCgyMJx/rI/GRxt
WB+jAgLsaly4rF8CztP+JMdb7+zFEcnQX73Jm37xRMOTnilRbI4d2OH069BsluXjqW9NKeATOltn
dpwBJ1xv7fRlMzAZg/lyBG+rkSxw6MFdqtliB5JXdFlYieeFDJDwseMx6EfLCI7sME07J45xXxrz
Frpenl3nRIxz7LQjflUx8c/h7LP3B/zNdTgLyQK3qQGoZ6Yia7evlEZaqwYLZeHqqd/2BfNBcQBk
lfHEk5LfJtSCdFz228h1fTu2n2/7Mu/nLRXJx13ImPJ1YsUijAwOGrvaeHu8rwyxJ4+wkfgJmGiM
mW0urBbq9VIYPb2ZmEv6j3x6nHEZNPvNQTRdAWH3f7Ojj3HOENTH8QsKmhAzmGc8z4sF2txLmNxg
Or21UqyQhp5vNqHetuDWgxTof0Z0kVFEbpN9XsTtJCZDR30oD9h1G/orj0pQJJaGaVxYPMdpUeK0
F21ANVIjij7ySUEbG8SLD//zQxzthwneim77+Wl3/VetDRiYFChhtkuBCh6oYGqJb5bUYskc0gVb
zTgbucS7nAs2Rn1/HO8d1yYwqKJaI00RIhyR4BHalB50NijCF6R+Ez+8QeQI675vtrts5TGpv+UF
PqzNhBQrRI90xiVQptf6owJgMvTrdQRcs0o1wSbawywGmvmhu/jiq0Q2JkvI7gP3sDfumHizqTy6
WUqsKW3Co7wvVEYh9m6zZgD0BEeEipeejyvcc8O34iv5qi+KlyK4noGMBMnuIE0xrwcV87gMEZ2w
HNrZhJdz8p5w0YCBUyMpNlWIfQAR6pyFDyvfh7uyzdiGm3AQtUfo2vEYodZ5DCTH3L0h/IS4oMvn
+yDBYjZeXlxt8bF+eQ7iZ8/fMk0iCJm6+R36FE3Mgae2kPYYKuO7kpcbCWurjuM9DZh19UXoA5oV
Ql8agXGdAvmGDq7YcImd+cLxYXakE6bnXJYy6A04FoCZhIVt9BffiiQq2wPYpJNtcMALBAdP6zVC
sEidpkee0kDvVF/wdPvp52/r7yvlycu/lT6A4EdSFFKJujNtOrjz0FthvtXV5+zefG2+1kyylXmH
molVYWlE5QOrI9JQZ5SRfEEegiugyFHz2dCSHQSdRMofSXvIu/2eiss5rrURLusZ2VCpbQr6Vsj1
PUX7H3oSOVL4x2AnEp7UeW3+5scj1BBabWJMtKF/1UHfFgGZ/MM10O/+tDx+crsC71naOaJMEf31
UGQC0rt04Ky3Y17M1vl5I5U/V65KFFMg+AX6R95bBzlYIJpC8oWBRSu/fPL7yKtcKO9clNu2FjtM
mUBHwt2/EPB7ZOOYvyY7grTBTpUNe6FT2TEa3FCBScU/puyQN0L1CXrmuYiEPSj01PswRRVv2hl4
Z75B0aO2R92wpOxHK3AgheR6wy6Fjs4VqTAJtvdauycjhhBsqI18Eijn3f+fgoINMdcLld336b06
XO39sysr1nbNdiNuhk8hQKiY0pg09Q35JqA42eM9KeSsWKrCF8LxAWek874Mi+9GLYa3UHWnJqwV
zjCIRR6j+P6hOZVkRUdfPjSOniuQL6gC10aCGb7LIoQPXGo/TQYMm23uYYEQnqqSV/UufhSnTNid
Wz5736gwLgduFfPSWABL5GrI/ivin9QaZnLxcYSacf3pKPJY+qlhgQlDAHi8BlqGb2BexRqSqSPB
qhGOBQ7x9MTVk9qIWBvPC/YA9UoSKOfEpOKR3w/uB2Y2EzVTk0hSdEzrujvhPJaraGbj+RgBOMSu
AP9GNK3+uQqoLBbttWc/wQ8axVfp5mwpBil8i2qxYgXy7ZNaCtngtEsXOiVrn0MX8ctfeEibdftk
5M6WYvJqud+4BHe3EtpGJ73MRu9gIPY0T4Iut8mWP8q+o4N+rFwwhwO5+2PkcDoNtLo0ZfAVSaTR
1V/JOmv9CrUgK3dr+w7meXQ7NC+9ZWS6w+v8/6km16v0vhKQ/BtD7lUAg494Kgenew37A6U47vaw
dPcVLzutI1nGQGOTJR4MCD6k2iB5VQy2BcdlheZUwlmFnMqqcyTNOjb+3PuWMV/yEDuYIUFevMxp
Cj7XN/QFDch6CeWB3kTqFkRMoJ8/hllfnDV1J2JsVoWStLqzOmgTsJ01/6m2lEP837pGZyMrUHGg
Y4TNONEXgrIYCpWfNfDcvX+wJfMGucN+4B8ZWtS5msCWBjnsYcmjNEF/Wai23FrBtYFIL4WNMD3r
rKKVSY5DqBuYr5snbTQjfLaZICMP2MAnfH8Q6vwn4PMkbHFsbSnD6g2b/CegVpBz1xoikgwDcLwj
uvEKccCrQBEJBToKcAbSb5U5Fv9klrJDEisupWbZ0T9YQ4DOlWJLavlcHXsQ6ivAaMieij4nDVKy
Df2glIQo9c+y3snvZvn0TU1RO9N2rnLoZK1x5esxKbF0PuB4fqjh7L7/ky1+YR0mku3K8++256sN
3Rso0NHYha549ehfIUTbSap+5zfxvsr9bo6SeBBcV3gZn40KIRWVyzRQO795s5w7z3vW9NutQa6k
8wTg6I84K+IgALwMC5dMA5h/6AwrF11j4P709AL4ioMyI11r6/qG2h3FsUU+IHqOdHfIXlBpPL+r
D/pzLtsolcnGXShIQFgS+FaNJw06Nb5lIRMk8Fkst0uUCnI8K0hxGI+/1uIPyd+bL5uaySTDepZX
UZSIZD20o+MMCpshaEo92QvJVHcK5P/zBwwRGBshWmvBP0arA2GCKuAyTiwOcOITbAaY2mni+BgS
Zlp4LUs0Vy7VKvvEAQ2HSgsnmiR//iv/JJUeEvqB5VyGDpT+tZS7AO+H5reW9KMgKcPnGaU+tWb5
YJfZ4HMYFJP0Mm2k4bZDiUxz+oNaA8BLSYsVf4J5704uxBQ+p/vra5phrXuacQCZ8DaqXTRzuUW5
eUv+5jUfU+koi4FGu0Bd3UF9qNUliuIULeyvTMRUPOpn8KPmFSHSS4ank3ObVELko/ml70/diLZp
AEa31IzFdiBJIDGUcQCLe1B+CEZhCUo6HnaE7ULnwRQmLAbJE3wAIYBuNaytwE/e0QrGT2BN7CTb
PH9Jxa5iwMxubtEiOtp18QSHnunspV6je5liBPS5Es90yY7pcCpvPTbUowRGHWLm9HHe2WvlsT9u
FgVvUD8yg/9l2rNCEJnpNnCGMw2IFlmvML+MzrM1F9GntXNkvLXliaQkUiS7NkQdgN8i5LZ37S/v
TkryuqhN4SJ5y5qQIFKKc/W49w3+JVaio4xHVDTRiZ7+fvUvFDNKQ9l15t2wYUtOI8MOrVTpHYPe
ND3OwmEiSHoUDV7b14TD+fRf0ebrmWjLss8zXNvaSSnAhj6TecHH/dy9NJscGN7ptXvqQ8T+1UBw
J9jPQ+yZY/U1RaoNwxegAQHBvwHq3KBazRji/9XnRQhp/J35CaqPssXDyfNJ4EJweRvKBAueKf+Y
T8TpMTADk5UXEoK8nk4oftLSHz9EkTUv12rnYlyOk3Lm4yLhHqn7+jTsIFKUBQrbi3wZJ1LIhSiU
nbMvkollUsi+zSvaoYs0vOgNx069koqcZYb8N6Hd5Uz9tjKz9qZ72rpEb2TcZCpe8tmssgVHLBny
Pu8uiLsGZzK0xyTclZn5qB1ZMBMLPCXeh8y6GsBdkUjOY/ZxL59JMMr1cC9BqSV37mLfO2Fz1vAb
wC4tSSM6gyXeDfLaE71m4/iZ/qvHglbSauK1dM03kMruPzdn/o/xSjwWcQhDKZNL0iYNc7hXPbEK
OItg7oI/W1MVAhThnJJAMrzYAPGUR43A0t2YL2jFjBR4igR5A+hjp7dZiFosOxcu5/vHP4nTyTCY
YGs80ySyZ1YSu159HEmxm/J44VLApjtOqbL6Y3E78vq+abJ62vOM1cl5qYJKdTK1ba9y7Sbx6vft
qldns9SfOZH61L3cJ/9qa5fo6DlbwG6V+8hsizh5lQF8rmq1R7BlghaqMwY4zhnjQ7Wra38Lptdr
BUl8QzEhdMvqKPSFD0OJdNn9x5fq1N0zppZLXmq5JUMHz5xYfEzRlAK39/pn3pY7VUuAbrWaxWAh
QkZ38Gy33mHRot/SZ/QMZuizfJRLuluyjOxp42PwwHWD0gxe/oYWZ1Yz19/9k4JuaWoYNuwc5J9v
e5/fsrV7xy//y3y4kpHE5vDg2mkLxIlzcIa8V1XRKF6otRDJTb1YSShOSnmzGA/V/VLbAwCVBmMQ
yJkngmxm0UEvAW+oHNDAFSo4SNBD6vPlKEJUE3wzFDNDGMb/yMJU27K8reLKkt9iPK1WCA+qoeo2
yBQcKIVYVLhW1POEF47Vz4vJql8RGBjSv+GCAiKM9NnNqlzOoBgVH3WUPwExPpKt90QCxmeFTtm9
HRABypFemZYXOeUwLqYAncpATwBuIbCFD7YQeoqBLyCIMaOb4PCVhnCQeti5t2Bw0TO69GjnEeJd
rhJaegLIeEZd5n7ALo8+fMr/XBcXTmqaYkkkuuR7x+5H1wVsOpIHqqDEUf9N83p8x4MBshVKiC2t
K2H87/luzPVdMpoCZVfgKNdtJf4B79o5GgyhCGfeuAM/eb56n7moQ2Nyk25O/GaJ5dCC06C2Yfs8
VJx9Px1icRsp7ZxPcvhIsKrqD9A8jzHQxpBhhNGEv0uOoHRzTcyKDFaArfoDD4Yi4iak7y/9GdwV
gjIglCVRviB60tuvrmcW4zRml71viIfwd82qydQfG8p5CHVnYRG8kvRM4rq302CUtq+IfIveCN/4
hN1XYhV7ZF9XpfKfiKEfWtYdjZNOMSPR2TFFKwb6tfk9BtFVaBi76u98uSdgKk4T+UUb9iSTgbf7
mhOfqgSj8UE2SvEP+8Z2+1k+Lg1IunDFi86SpOFON7KIVAVugs/WE398UEnzp0F9TCAyIq5/h6Lm
xriJwh0CVhnWiS9Lc4ghLDxgQ/rAc2GR0HSMAafKqDEDn/gGi7wNeipSp6+gBZOM2Zfv8ItRHGnb
R81ijQ3qsssP1C9Jp6r2HRVoIDUsvviTmHhgiDVTESmqT26GGhtF3V/UHFycfU/HH5HmsL3hVdPs
h2ZyaiJaruVnSPGh/pqhAX5MUBBjCwxGx2UKR+eoMahcK+V+Q2EhAVngi2qwHeXyepuxPLPFbc+j
NrCipH264EM70xsQmEpntzAnMSe7kj0EQqYflLH+dR7Z5EeA6Eg31ln9uob9vUnKiLobOcvOzV2K
e9pYBmxs6eUlEEgj/2pcRCTbzksR+6dl2WVHxAeR7i7pzqV8z8MBhZS6Gh2v240C27E8mYzQUzpB
UR/wofXn30SvhG32kyor1+obUJus+tiw0dODuhrtuztcl/jUHWBVDrKJ+tc1RSKJEXLP+3dVdz4r
89uy/CkL2/ZNlvuM62uK++UfdlPrmaZrFPzGywcrI01XxrWMTq6deiphBHhhUGqX/ls83cfGf1Ii
BjMD5ClkGdWyTUDzMPUiLx78St4ZQSraeQTC6mCrIUJri0E1rfzzVpEcUowRF16YYEbWfgKfoEE5
UXiqigu6M0UcOVgw+9ShMXU75Mm/6bA7PQwa4JQloV+6FRvreA4hej/O2DQpjnBA4EaPCG9kLq8i
OkjbhIsGNELyTlEmUYb57EHRMm1uk3Lt9JUi17jEC05mPxat8ZMBqpsgDyFW6cHAANFW4KF4Bu5t
cPCPgUPLtf78non43T8XhaTiXxWbvVlxxRCf0hlpN/DNtY8twpj52wbjk243eBHRVXjqjD/BRSQU
5atzawjnB+HG9oVYcnUbZm0kHWT30+OoHTlxHfJJ+EGQdbchpcoy9JAeEV+xJHH5rmLLWZDq9aUH
wNQdfhC5goEJvax4QUaIByi5XHQjeXRJY3N2MbqA9IbI8jz2wNuCNsZwyah080VeJx6gTB07iBiU
A3ZkEbBDG7h8y6IVBg7Pwh5YdLi3dYG3VAvHCkZUfeYpRPoZ7PaJtILnkZJttCJc4uvGCisKeuMv
ej37Nz3RoBT1MgQrkAlTrj9ABVrkfc7/zQ+Z03wYBiiMV40qSyem6gKvIIlJK+vkj40tQ+H9pRFN
w30yu5QMgeKkqW7GipqoGArlVKl5Gku0e8+fkNph/dGWqSyuGfoo79/qfbpgl+ToR6X2bNQX333P
kSLoJ3BOScjclGg3Ldu7SsmBMiGDbUN++k8ZroPN9+c5/s0FJSr30cSipPnMqszuP4wCLqSdZp7f
zu6DVlbd4c1DUWV1rKf0u8RcBIwPTiZdgeJcjELhRkVm33K+eBMkw946YK4J33sxIfAi7ohd85/J
qpX4+8Opjz+aQ/fC0v9x/0quMCrWqSIhHCzbVf3pcbAjywLkCkZvzD07iVGv5bFta2ZRwbFIAFHI
GCOM0iPRd3jUJbFYYLFyWhPOqVEOd59AYfzbryUD3torE+6t7/Vdr2BAph7wYp9ddhmNVZNHTPD2
/ukwf7Rq80+J8WBw8xUriyqWieHfu+0Tj9HwB9AHvHElGNmFDcqHf0PJepSEWXkPfCfG7HNML9tH
O3XeWdJIbCN4GB49VupTknz170r+sMgeDWvNmCIFoieCBNsTtZq0wL/ep3YXoBOEb2q+insf6Pee
k7/aPugZfQfac98HvAu6M6iq0EilTsA40gLrH+q36rhBY189PUPS/FJU1ZQLwSJK1ZZnJHEfGal4
1QJOCJ6Y8bYsqH7x+OIWbhOWu2C93jV27zHRqbNVoTct2O1SQhsncx2E6PMUBgcTBY8tXXH7oQhw
X/iW96nM7vjKRqwq8L0Eh/T1cfrCV4yF2vYZYWUCVtn0PKJuR3Ph5ewwu79aV3jb6jmvIl5v4ctN
OQ0UbgtB1OkdfUEBZxFNdvi2QdoPi6YiA4SaCpBM+sn9DMzXql/4avfueJ7PLKkWMJcAOSUMxZNF
02vbY5sRwpSfqqSy3trVb6sZkQ/5xdi2t4iAi3F4oQ4E86F+256/nqn7kUw6byHdyOjVmK3qjHip
frkEa9XnidkwZg/O3GTrWZ4y13f51ZC0K5FhAmFVstC3dzG1hMqjlmBAyOC7W+imMqPgIOxH7zr/
btXa/lMPLaw13foQtjK2aFoR7iGoeC6r8jQiVv0PSnXQ3hmFKxY1ICRrk7yasyZh1KB7jhiDa9PO
ESgNF/0FSBdWQDi5sEk7Ps5EiQVpup+M+iFNezYYGigPGw0kVkKayAqSdKLTljbkqdFFh5Cfvcsn
elJqJiYvTopMQjuQKzjFD8B2A/P+GAqz2A0eflo+aLMQLC9vLf5J3wMtZuAYcVlFrDe/hSKjB1og
qZyK7jkCgEP/mc6CfDWpUGHRe/GbmEAbW2ewtHAcdUgjxdAYHDUA0Cel7SM47HxPSZ36I0QnQ2DF
1X9yEtrIQs+mXk2cnam7d8s3xjitowS2CDiHE+LQDMIPzzkNYBVyDKZ4mVleVIr4r1QBjmzpv52A
lRY3oKqVhaeYoGdiFkWL1rcDzYDtUM9xlBtCkT8rw6OpdGu8+eYKKZkgA8OLpoTcYP0IJsK0yXoM
X+hvLE3+Tx4hth5I5j+aATHzb/kB7sYgwz7xRPCQqpwPogDKAqeihg66LiVYIcEwWn+2GawcRJ8i
OJqDnfEkeWiIv30amkrIuE8zotLBGfMfYPkbugWSCa0EFaT07WBtbn8F5PWqSL1Wixey72Dv+cE7
5p8SwR+PGl4Nx353JmHbheApDCcRB1B6LLyaWLRmEXBKOodTJZKnIuQEbqPpZvGBaqEzsl8Nox6K
NdAu7riAJg28njBQ3s/yS71DrYfbeBk+ImfW5j7RZ7v4KQbFvbhCS+5wnzjbAN09Au6ib1ACgr/o
CUSnE+cxdo1fWKe7A/6qYzAGKh+0YfcpGO4XoXTJniBmYjhs1v01XHAm0PD/aycQS4XpowSHXae9
kxVh1LWvQL2JvB68/Sy7dHXEpKYNfdJ4b4YY1s0ZQqaigVqkhUfs2vWw0JVtulHWpE4Rrkeef1hz
ImnpS/cQnPkMmt6YnNs6eGTI6zo4Ma3O4eTaDB4iPtwTjbrR204SLQlPt2DwqsfZPy2CLxsUceG2
7W1taeYhBFd1uU2CNPbDoAkK/wIwWqhwbTgPiXmJVtoAEKAMhl0nRbbnTBASlkP/upLDZAWadAZd
FwvKs/3hqazxdDusvsfeNeyH/ArOdWIeMqVDo4vXNm/GQ5Rysk3dQxIScCbJ/P0SruTiclloTJcM
UXDaHxCcrV6VDHnWSymYrLrmFdkolVfFpTaRFKKVFb2gjOOZm7ePMuv78U6pOjzQ9kPcFjHHBntK
SOlAdB83tbKzNAxa8JpaX7QiY2l0w/0fJe1Yx9ck5nFCNP3uYaNG6iniwRD/ixh21tgZw53XoFuO
XBeIElk6+v6vKNZq4y4aW7DqcZg6qvYHTy9YVFKiZGwZUZ3G7C1Eq/A+7ZNy7HkwtdICPk494hAt
Lqb5rfol7S8wSMHzJ+yUY+qMWXE6gFMxeH7CjusWQCpfThPs51Z51ZbiYp77IwD1HYuB8EWhd+CC
d6tlnDF05Onn6hglFLw1F3xa/Sw5lSj42XPqDHzyFCEHUhJ2GyMJi0Jvn9nnUXSJh/v8KOQV1Vo/
ep4XgG7F8wI0gNTepwFaeJ4rfh3tvIiOyMZ6YFnHepoJeTv79uFcSeoyLCM1DuWV5l9TnhwlBIJS
Bi64qm2FN6oWk4CRNmPFJUMUZocqNUdRxt7SWIhI8qr0jm/DFXsL1cLYuwcNCtbd5JGezCjZgvHG
wPMc3DnOMXcbAa7/WiZB15KeMKII5Hx127TsTexxa/UDxzPfnT/AzgiPiWtCe2D74jyB65qUDn3X
lGN9F3MvQ9HzcKZofSiKXSfCStTmTmDGGRybba4y563oxSazZ06n/xrXL1wNrSs4BcnMI93m3L+j
uhG9XAUMmiElfUAmW/7m7skiJ9+LDqGEM71fyFpD1W0Z/+SiahNz1gu1NpcKg3Ra6JUDbnsx42zl
FKwnvSB9eaZ+SlkY9EG9YLRRN+r0HxCQRzUltQTq4zat7KbNPwys0LmSGGQOUvoxsZFA4KmkUOya
Q42n4Pn2P4d0gFx2X9xnkhEYYk48cB1sTzUO8sJyCOFKvFFAPoghEFHVb9ORenogRTBOJeKbdW7+
VLYY62SFygqCW9bfSpGiTKiH7JhNklNfCUNySQXxYcSvydBf9bJNLPgF18Uwzpl57LLf5G88EAvT
Kdpa33Rcy5egpGbyqbGhLOqrd0ArZPkBVJTj7VrTSEsws0uzL5IMUAKAyYvo4yTzsMlZ9svB1hCl
HZaM5CgsHpJ9y1A4K3Ts7pLSKMO3N5TomkCbiaj5N4azwSzoEWT3jLGMTLwIT4aPCIqGlqhJmgSO
+SQxwSrj0wm/q3ar+p+iZZsZ0Nwsun0tHUAtQvF5i9+YUqh0pmCj1AUhISak3s1Fh9qWYk2TxYaL
WkODp2rMR0GoGIeh06o4qRMVVWSKHrrqMNdKRRkzQlRMXVcfU8NF8nw76yMlCXJmWw1v2E2sYKOz
Cca/r3weI2wfH0dIj9cJc/jvRObK05688DyxRdH2Rc0aok28ZLpCSy6xmUcFGfNN82d26C59BlPD
xIKaQd+89mWNCMjctAzTpCopTUxgyp+mOAJCxslEDpysc/djoTcax0vlqaMj2SeSYFopOWEDMqtn
eaynMykh4oSzDzVBrQj6e2AG6f/gWCl3KMuUyiXo4BE6wV1rbYCmeFqOOY1+tXMlrYXnlIiXeWg5
bVQVqs3jmC5hfkoT/T0Dq5VP2XPojeuzLamGSxwgmmLtQen7GQcX5SfUo3f9YkFiiWvqgrk/XMiJ
VvjLyrcuMAmFnNL8WS3QlbBrvcHAWOdW7Rn+72LU4mClJLkPID3qKN+98bHRtoF5VcMeMFPvVe/p
To7V/gy9IdbNpvmCGbUCscFnWc6j+2wkoOGkIxohW+urFcoq622ahfWykTmPqegYuuqgcdW84UeQ
3DEzgeQzkwy201sjKoaByPy18OGYuA/VpX6qH+okjuYhublR6IaKLWsSsOCdHhPBmuuodFwxkW13
33dIDQ1ILY3AO9xHNFhaSVnwD155nxS4ScMGnrgT+o3XNxoXsZcyb7EjghI/UbIJlOSh1jdLSBNx
KtOvzIrCzzob9N+v1fRTtinyS8niNdj76QCd5lSxbppJNOYy1DW2QOuT8aqmnzTgOs/eyCALPgZt
UOqtlhrcl/StO1UctObAcN60IZCO7c35JHXSe09erGvxAkusAJlqsZkYohBTzlAM7Yxs2YSuVcm6
bZUogkT10tQ5kdNEbh51RiqyhEtHuItIBxFWtJjA9UYW0X672gCK07vZQU05tsu1Nf5IU6CJVQF0
rZwpsApnEWvuGXmXkjMsBcEQWDNyFWwCmkz2yZDeoJFQbP6y5IraUK7GquCXKam+GQaRjTNKSAt2
5CMD9Dh9dDFyrbJQU9u02bSzoYjzoyV8Lbtt1U+YBA2OeSHj8rQtgjq8ECNr6vYYIXQ2J7iJ9O3D
KBIWHQhFWlcA1HhZ2GD5pPTBf4FJzvVVaTBpkYY85c70793AsbM6hix4hmyJ+yqMhrtj4xQaORYl
R+npPxSLj1VpEI2ve91mOHMeBTwezxlE1gy88b0zuNUtBA/NuuWFFFv0M14gMKgdnw2PHEd9VN/S
xnXel7de65zL5+swfKaEL10uPcMvJxVvAArrcnRYnWy+X56RQrRjp/qhGUEEAI/Tq+y+0CIvGyrv
ZwGXRf0FmnSJrxIF4ENtsDyXAqIWmpQWZf52YpsB9/ii47Oy9BtSooWWu1eH2vlssHJMuPaPy5JK
G0jJvLcu0FwyEf4FOPPSjdzXjPRwR4qoeutsC9s2wxDGnTLNW1z/5c1n5KOg9g+2LCJDAFcIZRUo
Bi0tWRyGx0cxaxP8yfqwI4+84a0XKPt3DqVkdNHo0Kw8+z8AeWyIJsfl8RtERA3aqZV5U65sw2FA
RYNKacPecFye/iuvvUXqkR/CH2fZUQ9i/NLLhDHcw5DEFSS4DPj6Vo9JjuItZgs8Nduoyz6a5mwB
bqpjlV77dcVDS2xV3fDHFqpw+QZztJQuH7efzzp2uEdu/9dCRz4bCd/BZJeg+ptmJ/Wezv7jirE5
7Lrc523JOxBo53EFyroRpyUT0v0VnRnPxARLrB0tmXDNEX0/rk3oUGQ9Y1Xvm1SyAnIgo7HfUgwe
mZ8X8fupm9jisCLOXHN+2UWqSgs1tOhKflek6716Vswgvein9mNieJYFPFZxQiqV8y0jaeb5anve
S38nifgLmeEMJYXPGR4eF1oSQOo1jpeKSZXmRkGqP655IbEF+PkbG4TZRQrQhAtx/0gcxxBW5t5f
8UwGJrXlfNAaBvjZamtkhT6Vj5kbt4eR2cj+EL3UdEJPfE/poeWK6IW/tjpaJDLRl6xILhmBrXhv
fF4oLbvZK4sK76bJ523S0sZCR0BciG+riGJDRCTEOUxgh3+Ct1OKpkO4+AbwJsqm9OhNNFKY+fUE
pUAP9nwO34WteCEASWfSzCQmEOX5MKeUxW1cQ2gf8mxFrS8CR8wzbutFXU5rkMe/zwBDhI3+BaiU
zjAZemMndD1axZZ5bvPehVdyb5tAisooQ71flYx1YaaRBIpr2xaJ+znBCyH4CPDIuxWkDz6q3YTu
oNcfQPd89M/X9GiMPIx26QyCtGfo76A1AMFpJLznXh0CEoAFHRDd3UA76et9pasMuav6wveLHEx6
bQ0sAM51Xda4SSMSpdqoiEFuvv6V3JaE/Tm0gU8lnAl6E3rnhsmCBtWS09nc8WIBWXqHA5tf9vB7
n7bHyWLf2Vg9E9ws07my6BXDwORGUL7dzZsB9pn261Oa2zmwr9tVuKNGzppYbL72P6WTFPt4usCz
gbr46P8DJAtCcoJftE6RE/9ufuzLU5fz9K2l8qgmyEfS23hUP/e7wTKqcUwFvhc5Wm95+pqUCkCB
VK7gWjTKxc2BTq2gCw54/rmTvyqBqZv0aMaWuwkxMPRrjuPBKaMTq68YMtT6jJSkunj3UYHYX77u
AJSfxUVGFwRaheE8EaIQVcKP7RqIIQQqDU1mMDXgjwW2InZs9uykrr2EwZ8WfoKIEjL9IDFDKv5E
VOid04jZrrK+BC076fL3yDQ/1a2uocURQh2zAYJMPvs5yI0eXpQADhz0RwB+kBX0eQWF0cQDWY6w
kTt2Pa73GqxtoliAj5vP13NNN2zs+9wZVWolDERI7XSoheYs5Vr5SxpFKgmRWHfoqYZ/FbB4BnLs
8YY60LVjHXKyLDBxJ0X+v/0kyfb8v8NsNayiOWR9wdny5lGc7VkRe2TboYk3v1vr8wUyA68nD0Wu
kjmmTvyFLuCSsp8WESg37qoBCw+NpGpMH8TSBdDDp2mq3NdXtD5MmskIh/5CeQtnMCrW2AQNoHjl
5XAgQTkowSut3Vjwq4sLM7bGd6X8lnY4U3dSz/eWSHd7v+w3sO5kQYGtY0E++dr5ao9tYqH3GPNy
URbrp2/H1HPEXbn1Jtw//UAOLnhnhQFLONfXOl2a4OCM374wTJYWOeaQNAVW90ocMRSneAAlGiwF
WTNfIHyCAyKAshNz1IgvtBA3EQnE0nqGaFfKCOuwIp0oMZdIg+xgiH8by+hgqk9L17SUnl/k/hCw
4Qzz2ibzPN3Oj2UUJQLxwcHVdP3Wj/vdSemu2JQnonnHsrUuFT+WLUZpKkKLUTeRGpxlV1ShKO3F
6yW535vjjVH+bhYS5Y6dyHjUDAaSw0TDuqkpkEBSr6FVLkt7A86hzYpTUChXY8Yihsx2nRwjdmNh
uU4CN+BoDo/EUqTg2yqd+jcXNUZS4omxlSsYGs7XLQ1+KjgHXdNBgLCFni9jpKHk4xHKThy+gLEU
1RbddUUHr0zg0nreMttGT4zUqMbZO6GPC12UBhdUB+vYmmRtsmKXEnvaTsQcSNoWGX/drWSgmILo
hpEAPJGrIBCLcpq7o0scdZRSmOLPo22CwDoolQG6J+7ZlBQbOEQma4E9BV7SBLZFQSIcCkEhXCAA
jeDncufJ2cprCCeK9QYGa/3I6iutxPduKgKHRUoGtduHtCzGWK2G4sjht1NEEQwc+tFGCE5lPZQe
WvNugbg/Dp6dndpuyCRlxDUDak3aHgeKDcHbriUX69J6+kcaWDinCibyHm2ff14bbm9xRyBGgkUF
Vf55lSMfBzfYbvBC4EbCDocQv4nQNOqxDkw9xiTiz2QJZRXEdzeCJZn4ys91aRnLPQS2Fs3Twk7V
UD2VJRlmIdYJ8wxgjPOdtfag95k0qrMrSMcdAuNTkIYtsihTR1w5nj6qYdP3CXJTOCGxUCybme+A
uzRNFH5eOi02OOu3uPCWk2eddULTwpSPt6HX+dNeFj7Uh1jPaLEMym8nokNqMLJp0qA3AFqHSPz9
0Z5//HTWa5TpboN4jFZHEc5DQcqzzTTedABO+ejkOYQNi097qxdqJwNlWnFUYS+TyzbwdbhHIkI1
CtB52OraMti6TxAsmUL2IYgLrTTgX4NDa6+QAPf4eJSMbi53yYv8AnaQVg620jjTPRcmG92MsAma
nkbKGwgJKnjMKtbPATw9O6K8WllvoZsC5UbEHwCLA9xaLTbz3huuHfM59m0VLzKUOnZajugl/u1c
rqGzkNQdLIecWbWMJfo5Y9nuBZikiiObsLjJxIhHP7YmwycBcvybHR6bHrGGrYgaZLaBY/ZIWaAu
DuNiBkKlGgiPKaVfme8sGPRNTUJkpJGouc318XUAIER52CLV9JS//hYCrkOjNHBRHFl92oypq8SK
RI1wLsfpe1AWwO5H6cwruvmmnsGQbM+voaYf40+CsjIsaeOXAqVLerbmJTR5v2q4GnrgzF1uq32j
tKwPTxx0I776SZyQ9acsRuvSL0gQRqL4+RrzAXQyBZxZtB4BnY4FEjY4z9zm70LG+LV6a/RV5ISl
QJnmBv6arVPoQjKKy4KHCpS86alKwFdP+FZNIz959493jKQSGv3NaH1H1Ut14fYGrQ7CviQU9+e6
WdFPfusgqOWmnS2i4Rg9QyXLt1k9hF84zPB9cA3NCQllHJR0WlC6BhM7ENne14fjT8c1Zao59gnM
4ScQ7hCMNblVdn1wqe6OKret5LwnK++DroZJAp47S5CO8EU+gu6l1INTxyq9Asi4sWYdqVQvKOYr
gHnjtSVDjlkDvPE/bPOAwc3R02EcP+10WgKO1zk8YU976LWWxzbR8ZbX4ZKIYVsUedW9DxCvKHbA
4Y6A5zSskwmyp/QDKT5iJef283DPzXVH6FmlFRVdatQCsUCBt1ausqp8TmehXEJblgnnsUPMsCTD
1E6AXeGNSobbi3J+lCH1By013iTh0CkGyHy0/DnJGwROjK9Y+ngk8MWYP9h48eSatfdziGkn1GE9
xsRNo24nyGHqfNWQPkd2X0RNfUNcvDWDwKsOe/cb9wsUO9c44YXcwlAayJSKAz0inUc5fZNKex1I
At1P1YEiuVn5+3z9Zh99ctP7426NLwGWvFJwAJXH5i/WlLTL+K0P3BSACC5XRd4dFoSmmyqjUyPj
OirYyY3nqL9F5+vGnqt9FA84oMMZEeyC+8+3V3W/iQom49ZDimHq552PV4iq/ESwAWEDgE4TTHVs
eEX/RxYZpHhlthu9d6fbEIp6XAMEk9o2TVTQlG3Lxb0iWdHp/hrFiM1Nl944lR9lF9VPm7hEmMo1
qdpZoDtwNU+5xXxk/FGNr2WKFYhWgLsHXjaLenbHsFVWEQTk4tYfnBvSIfzoL77x5Pmoj+5t4rGX
8nCyPQf454DuZdr4wqI8jSXI0Hjo5KLRzgv98Ld8/kSndAX9L0s7U/DisL5NwaXqy+ol05heXn9O
sQnq/rFDbZR9bMN50LTfZktOJHZEGlKv2JiuL8MkfCDxX2gC2TwW3xI3z19X9vlB/G7/zSlPhWEV
B60RNoo8tWD6Ba9bJmxtmXrr/ZE+eOKvaiieJUyEzEoiJCiM4PnqaOD/Tip7ZaZOs5KyRvf5ynHW
vzq0gDABSIceW+eQD5B2RuDg+xmUcGMoiZrZuqMW++wm8wYChhyFDzurBvzsVUd1ZmabU5iqV1oQ
tJ/c8gux9UQhwaJPP7gRwuI+FpvGKgGFujbmHz73QhzVkpnTGKgUL5xheDo+BrHwQu721ERPKZK/
MzVwd690q0N2yo0yKfExqgaFTPobILIpdE0lgOsD7bKjyAnvEi8duQaaWoPoXaZvfi9/E6kX8nw/
8ExxDRvS1+xzX++UJDq3qM4/2Gx4npfiUnHNx0y5rAQ2p6TRivZDtyJ5ROf3xh/HUsFUKJe4R0zB
VwFpdyodAWa+TiAAKeqK5f+dPMhJd1OudhPOPxSIAuwTqwg70FynEqHNBBXag+2MMqxdvF29bVEF
DD+hNPRRiyrbaMpHExVQvvv/3vA1WT7hmc5/6LQgsruizOedjmgCHXvD8F5codE1VtqfDoyjnsC6
H8rFRuRa78JBIrhMph9xbaN1ec7i3p+zMEByLO2MAkJccDzjHBnMUmirW9gx7/iHO33ttzCGtKZn
aSgM2f8APwo/kjtvAkxHRXS6KIdAp4avHH6Cp1t7AeScfUZOHZfbkXLjpeIKlAK1kuQu+AOVtrmb
3Eg6RCtkgDV3NSeTSL5RES1jM9mklAWyBCwJmeFoitW8iG7wAQmOa3Rg6PBGVRBcortDjY84480f
Reu2s+AZNTS/wpY30kbPdomhMO13deOM3opEidtafx6iVN6eUnbkvybSiYCTj5qkm5CU/IKi7YeZ
VUfnnxQlDqF/3/bTan+WcwqYMG6BR8r+yXolRDGqW+UXPlIONLwsXWDjfgT50tn8eoVRjuayL6D3
NBwsSgm9TbKOqiCT6kEzhx+jvxPYmLQHgv74JX4NyDzt9N0ZPu/Se+snnqg8nJwa+pVnpDY8VOhO
ttZ20fBFebMTmVPcQFALoBp9uEEFlMtOKzgtVDhjdMzVEWBdRL6V8E9qfUQp42L6NQFpwvO85c17
cEwfXlxM9VK3Gv0BHwB0yvbXtoaPJbSgGmWdBD/eUKeRP5sHA0aqv3midMQoyMejNLsma1kCiNmi
fCOOrauIncGTOFCS7sblIgtplTa4CiSAHK/MYuhxD4oTLefreI9SXvm6637r184NsG0D/OLqpeHR
0QQSOxHVnbGCRCXkXvocCv/3d13CxuJA69VtWbN2bbLWA5rpREGhABrLiEntBk18z7N7yjQkWri6
WsRWz63BW+54y4cbzufNB4PPuTbqmLexezE3kM9u/+BRKyrWaUzcu91B2VB6TJpHRRSlt5tZGnML
K0PPNGLWWidxEZmkH+nwfSScFACcOnKdx5sz4oRj0CeTo/e+GPdxs9C/L9J94i0SEfIJufbG+o+C
Fw9lkvHYi+NSSHmFCz7+4myaDiVQghwUQWevugT6CiNevNrIUgEP+IkqyTVRTNGNmIAgwNM/SVFW
uEmGPDDQBQxZyPjB67mAlEGeVmIpKL/BKTZKE5KStgwL5iVkRyH4v9l8B2yLn6NulnW4JGXu8Hpi
xIBI2w7sOf+9Yhc8bGLe8QSrjGZi/m5Q4BynhbZ8vZfpNMjcA9KstSoU1ZNogHZ8unJdb47Lozrw
rzNfKcngYJFc9LB51oVFt65X8+Ya/UZJm2b8jqvvrpYpGxed+1yy/xNXxk+ZWEJVeuBGGggPHb/S
arvMPSgRsKDsiHvuzU+bUis6gfm6FcpWwL4/Z+hG0oDKo0SXIe7N721omuNKZyJxMHH/3I0+hBSI
5JHJveMmotn1lkVYj1cZXQcNbN8dNU/POF8StkiOigo22xzHen4uaonTcp4eHDdqKFoorTxSeSGA
ZJTaJivU+0YILf+6XBQ8hG8c+FmIoC7CU8KH8vCNh16Mgz5y4LKD3uUbnGJ8RzqLEm9fAvbkhLX0
MxuAj236inJO5d123wc8FZ6o7tZPAkLqkNXyTcXeke3vk0RI8RwCPOSjT6KhQ+/FJM6yoF9UrWjM
HIgCHkR+xv5VnTSE3eGuFhmfW4GJljFsaje7DBBxZ47FaYOJNWVwsFDMYwhX3j5hN8U5QmRMI/OI
zHZCb7bOIKBjy64mTDhnKi0bHB/INQf/2yMXbgDuEeC4ydHKDiZm449bV4wkPUmBAhVo5pSMyt0m
e2a+eKOrw7V9396xrpBe9mOWj+NZxny88BeMGy/5m7uDnkiWzARjXHSGTB8m/Tg8oKBWVYlkbIxI
l/Cp+dUQGNMiyZvM0aFhifyXYcpUTLVHqum2gsJPfaPt1K6fQgVtCor3oA2XGMyTUm9zEuISsF/5
fZffBRfgeIWwQ96RYx73GjIkY8HihW4Pdvnzo7jmEZcoPQi9Pte8r3ZB7gtDvmlv3qeyoCNn8F85
46VnDhRhLQSFXx/O4huElm3w6npQzh3ouVy95REgKjBZJOiuXRII5zgcBZG9ilKVRcksow2b3rRS
QaOElG6x7U7HNvzqtineTULYmoPRPNnJkWuvAM/X5PS0q3JQM5eS1Quq6+1+qUPB0hi67BUTNpqS
MID7KXuHB5bJXppBTCWD+G9vs0DYZ3SjO+Tko1b4r/HQC4GLyTf0Zkxe9Q1cqo/omZtcuDgEbPws
6FhuMr8Iuv2bEuNfhvPZB6DUPoz0dy0sQvtwiHwsEstzdETI2RFV4R3jsmMj0gT5XR8kVmbN26zN
ihchFuXUSkkh+cUTAQz7v00cb6EjP2JQ/gXz2wBzCHhWlk+RHBvIK138PS9wXJbaA1cPs30F8yDJ
o0qBEXQOtD+5xjIYd3F+fE+UhYaQ4/1qpvQ4vuim0ux0qPjzr2px8HQBiy//INjnorFvzIRHV8oo
0Yaki5Gjc7/PjYeu/u2da3B70Bn4lCCK7l3vbU8PjNjppniqNYkSBxvgJzUU8dmtEr5Vrl/0Xxts
TQUTEw35PKp1DI3fASjzvJv9aY6INKyb2vOr3kVDIcVMD+kLpwHE7qipMVAIYNmmgMfVWwwrqvtz
Gr6agGYqr3L8M91okoZKlqkQXH+dAj9Ilt3I6YU+xK63sXQk78jXTEkrXAoz5dDl20jUYUc57bDY
GjUK2mOPAILDHmq8dHO0WZW2xcBCKkQEN07HeR462+fcBc3znDTwuJmivdDnEQvj4mRo9J5BnqNb
q3F1DHUe5JXzvZkz6QgFBs2uN+GAb+5FBbeNuzhZDFhSLwA7dPAwbzA2WXjkZD6qzWv2RnBUyuXQ
rXVthTm9gxZhLNjhW3Ox3U+u//56QvHQJ2U4PKqMJhWcUFUrrPW4w8qp5mdtk6cDyrrxit+Mf42i
r+ZqGS2pq09Sqm/GE8svS/iG9gw0xxeyKtwB48HT8gybjdwTye1XrmswHitxrrygt7HOVgRbqM5e
D4pyTa1W4tYI+fprRJ5KPyfUGi4p5U6qSjBBIkKlBMDwacOnxWEpzdvS4bUhojwluHgY26YG1KBG
w4EHv9SW6pItqSolMjFSnyG7CswIpj1MEbUP/DkPRj7FhwVBH1vJbvGQIsCGze1l1afEOubqAFLo
tTLBaijblb45y8+yG1gP2VJC+nA0WLn6zBUphS1ButotIIj8S2K1CsICpmpMQb9ACcT6k3rcUh27
IkE+LYZKXicIHV1tTA3/7YkrMkQzO+tel3nKahBCV2za8yPXl67mOCb8H1jM5bk1VRO90pdDWaas
XG4HONxFWGy7EySXCTNhK5GHD6nSrdzVgOysEhgLZqY+s55ah6fQjOEYKsJjfj8lAHmPSIH7oYZ5
/ev9+y4NiakjlElDImQjQLiXxtLo23AjQMIgmPku7DmOxqRFQxEynpaQGSDc2455rm5bCQ1ESWDE
xd6guJjTxcdWO/rhyDS9+syGLBoVsfJFiuHFscOsP4U1ZrtqD8jlNRWFzt37AGurcQ6E90BcJKXI
m4poZRZPgI8gglj57ldzsHIfSa45AK5tchEhrGAgxC//verPYoSsTynoeyDhDp8+dZh9eP5C91r/
dXAHP+R7pb2tgpjS9UUnh/ibDn5lUcEptOr93emWSJZDdaybbP10Ml9D3F/l+Zjl+iv7GndqAhnZ
7e8CiKEYQYSdMOLJPnz4G1SamQtG9SmSxROhULlSGoi/yFkzsA8E2tLs7UFyAHbn7L33pi2TShlX
YQ9qZza5/Bye1Qn3LFX+qItotyqfrbODM+kWjP8lJHqn7sCZAXAE0NX9kyQ1CkoymBoQarhHR6ky
Fu1DxiiXvp4kBtHh5nsyPOSYRqz+ukFETI49iCpgKIhp1mVuWwszGMsidRGTKdvkArBHN3sElSUP
T9EbP9AKZBRklDAFOhK5PGj1eYzBNCvUCgRVpz8+CMdYuBwbMd6Q82s63hiqVF3ZMn4u6DWFNUEt
a8M3gQi+8iTCWDYWUKh1dx2DghZ1jlfwXkp7REEljlOnC0TG9Yz33YHrPHTYIE9EY/TGgfGLM59i
ZMvk7KKwrr06ORIGYYvvg/szCMqZ+SbsqDICF5fDJ5qtU9dRlgsi+ejgT/aO/y/n7rZadKTKplzf
KpDxz6yJxpnymAqANKiU02fA/15sdFAj3lbn3Yh+39om/R40t3NF0lvp8nU5jFH8JQyR1tTtkUhO
bVZBDieECf9ULzUlGbeBMXganEoWMn1NHPvM86+dKQxMM3qhyughzzO+SCA/nk28+ZuHLuyI1E6X
43FhkLgHOhkSj086NgXnBTgMNohzw5V46Uv7z6Y62A28Gwbx/hjjVlSWhwcBiyZ9OJh8ja7M5WAm
a/RXt+yr7V+unb9al65bgyuKVtvabUGHdte77EEfKbgNd4IdrhVApYJ0p/Xj+egJSP/aoUTdwzrw
/ve48blczw9D1IImdVWbRlFkh8Zg5WcqjyK/KiHIeE8ygKXZbazqLkrdtGP/xWnxpjV+9nB9b4zA
FszpyA+YcwuEArSb6ETw6CU7Ii+5+gHkIUw2WAGlxEGly5w7N2zOvuszt1mr5HcBELSCfScxP6YK
pAFjbT99ouxooqBbXbZ3LPdEyFqhH/MhJUaFOT3W5/AmkhnZaG3Xz/8W5QTS3kbP+e/SVcpkL9gT
/R/HkH7+Rgmf11DM6ZWhYLG2h4RtXuYaK/pX6Y8hYyxSXkkKMU01e8mfzvxhcgajvY3JRROxDEB+
KoRzKpN0qTjJdS1lzrCL++QRthaZEl7ZVW6rmYJbXQChHqcMyVRzV8hR8rQAcxChtBzdV//GyxkA
wiRMZmPjTTBx87taEe1NVI/2Q66jB7N5p7O57KWxh+vM5Tgg+84ytaZ41XnwH84/Jvep0/pCVLBI
talvPUYXODgQAk0yB5GAoiBQD9VwyoJdfQfJ4vU5FFwxHwRKDG/xEB+evYu/Gbk0RkHvNviVypIA
fNuCc3cldtqINQgpe3eLaLzlGdT0ir1siKENXk0D1/upbo5KVpbT3iI6brGxBtvwI1lwT6EGT/FJ
laxeiymXkZOCj8AINZF1x3lki2vpXirL01+G6tEjl6ASxLkooKa+ruHHAT9ybiVLAAEad+5vXo2Q
PAgBDI44K+dxIIxECzdJiLbzJlKuT3mqYhrUAXD8KzcP8I3N4CyJttBdAr0CHh3LcTVO18wfbF1y
mDD6o/worEo2GUDV6byYoPaPPgd8blytp4CzCf/j3Gl3wi4mpRni/PdUSsgI+OAgvyHYdCr0ujjl
fE8vG9gIDgeQXlj+pR+fPkL+vPtYNCnx2L4m0IVDxFRR2ml09ica+WlDH3U1WqbOEK8wy1oOaaT3
ltcYxgrRn5o0wyXg4MlKGN71ZkbFrBqS2DtzNmkQEsY8BChO/8SPG5UoBR84JCQA15H1JacXd79l
6IzEv0dMiDXh+qi/W3yvTBboQt/xXjvTaMCyS4w9XmKqQdmup7P8xhELzSWaTks8R/Wd8bSEUDSe
Pbopc4vDV8EA7kjl6WgV8IOKXFJsN12ndJA/CuRJt9DGa6qaHaS1LuZ3pskNMwq4ZLVKYRZQOvkh
Smv6fT8EQla0bH7ziIrhjurR+umttsE6br3fiWFGXBXB55ojztUsfifBF2aXU2HbsC6raxfL+6U+
igLHPblFrknWpJEumVbsD+i//25tKEpdhPmpf41EsTo+wxnznwfzkus8UqVcbf5XDSI+caoAleJ9
12VHgecObPsQUs7qxqipxIBhqx+FVX3dP9Kv6o3myLYWuRKBV9/biuEf52tJpee+yMRR6pb0K2Im
9m0U/k3klvuveZlDe1K/Aiduq+ewKa5A5JQmw5tzm/R/nCou8cpJr0N6Fu1crzZpMKAsgNi7d//R
PaQ6fPqVskWoKFSN4krZH2ukGVWNOZWGDYZ0pqgcHmXTxMoTPngVmDzMWiVlo6a2a/W50BQe76Gd
fFuszC0oehNaLjJyVEhKcOC/j76NjVwrhbJ4l90zt+XVVsuTWybNaRahCfCCRCLrMCEHEzNZU6zm
zTkCXkNjQWemZ59MNQOi/QEFvdMLfI012nBMQlulQPZ6+2kv1edpUpqKLHjo7TJ3DX6Rbm1VFmfn
wWeDn/J2gWI9wV/Jm+fuZXB+OdlPxPK7KpTTTOip1JepGkxI5+jCSaOmBZeMPfbVwt8AYvWxKL7Q
h45p7vycoWl3fWmN2O5FPtmAzc4LJmNyx9OYAqnauAqw2RdGSz4MRGtqKwPdk1ruRkb1wnDtNhc9
88JqJL4OS6P4uJJgea69xMGi2KR/7enyugPMEJeQ7UiitoFitxcbX3jr25hp+XaUuevRPj78IO+p
fxKqpWJbM97Wyag3G/Nhx66bR+/VWqSh6F+if/OWSeXJ1/iaMLrzuqAodruajaW3WS0UdKqFO4gz
C27GPvRkImdQQKBqNZjiNBhGn7Jsm2PMpr5gfC5fEhQ5I7ov3KlYS0PX5iT+puOyNQBNKYaiPhbO
epMsztEofqY99p10d62PSEBUl/YWsg/oPyy0n35t94rfFvJB03VccHXnEU8gtL80ybamsJMU5bfD
u84Bp0y0FA7w9GdZH4FhxcySZ4rWqLZaexb5/iwVaUYkM9yRii3ZJOEWYDJI4sF85IGosZLS/HDB
w7rXLw4fLwr1ij6WdOwydUvzl/QfwZ2/DkjBHkNYJAjBtpRWRWpLtj4p2Qk8LMyk9iQutRivDgB3
qoqf9KMsKz4Tceyf604+Mc1ptxea7AQaNJwLK8QkqaZkq9yEoS9mOKfR0Sg3kMY2pnHbRTdwtmbK
dFQ3PK1OcO51AHyZmm3SUOsFLYfDkMUnrppYHJN4RKYiIm2S8h8V7jIHO1bU0x6x24VfwXMoc+nR
VrH6s+ptfPSGftCC+n6Swt3rPXvUe5Ffuu0ibRygoqeiuOR0bD5KMfRBYK+dEgV8M9EfroKEr9zh
NeoZ4eQvduTXl16yaRhl5FcfpMTy93F15r8vvg59+dsQdKtvq/8xyOTde42+RyUQ0xcvjnNkmHIW
djp4sX7BExe8bLl7bp0wey1+P5c2yOB7hNTqnzzTUecL5bGPAQFmenZZE1/eYpHB9MwLD2FX2MSw
bh7b9SZA9pmIS/gg+cJAZM0EQEP8xCszFeaBLwaIDecM7saaDMvB7IqRA3I7LxOZEAf2oZhKpK+P
VexuT4+ZyUQIRdOnJO5eE8a0Ao/UztBweOhfoDOem3CNDBG1nDq2m8NQbWMssTaU5VbXwW7PYoV2
mmNnUrtUblMchoUkBkmeKCieaEZ75CysgV8UCsbEdNKkWNCuE6AVDwoL1V6lX3hyKbwx9pFq9Rmi
/xDONskXzy2U0fMhpqhxT/SQkSs19slYIxvjU5UpANg68NhwYTqnf8fWIjGE3kFip9cZYyAq2ZIJ
bZGvBVIibMoL+lSbckobeuRc3H93TqUeyBpx2QfWVI4uPTpOm0GSztZybyXUf/aO5wB0I9FTiBVy
gWPt3W7yopOUMw24xJJifsTVIBItnPCGpwpYPfavfOGFRjvHt0NipveXTMEWV3uP7DzPE1eNA6fY
5DmJQtpXSxd0VDiYaGycUOLj0ccjLvaKIaAOP6KIG7+ulVG+vUlD1WDUQegq2R9xE2kfEThOdLQA
UnR012OJ2/pA9+yzcI68o2+S4Z7UrozNJqRTg61fJ2q6OEkUyIJs/Ur0W6jRTQbs/rq+mfTaj9ir
Md2ZzcAMKozr3IuOfskXJ8/OdhYkpOEL3X3QrGK6hfJQNRadpEdGHEzyYmwMEoBYgkL7EjD7IOyX
yy2siu/j1rf42dJuB9sB/MOocxk050I+L/ZBmr9GEptQBgcHcs/3PE6mTWNb1HzYgmnytKNhLwiz
+ISsr5t5JpBO0ALdTl48FyIYIaBrqdDxPoOp32HMF0QLdxn0xbda8f8rL0va78/SNZG806NlzVD9
imD4o2g1LdvG1VvuALzNVsluww7sIw64Tl3SGdahMp2ShnXv85zsLCI/dNKR5b7Wup2/RXpXvT+X
provmbgPdjlyjZX7/XQOF/0AM0Y0zn8hghuhggNOCpuufntFCpWsXzXkDC1QHbSkyohtZ9Tvs8LX
bWoFR/zswNZYxuIuDxhVmKuP/D7RSykHVueskrlGEQhLMncP5QEf02i8GGrzcRIaCi4wWXPTtLVI
xKbkcvld41sevmCdD0QrYVhzSMz0gBT0v7XZBz/wLw06rEX2jnSUrG8qZL0xRWzymG5iohynT1ss
qDu42kzDE4cp9sz2nW2cf1ADUmC1IFxtjbe9aO90ctMiIkNLQa2B5ZZj7QLv03njdGw/Slimmmsh
ykUVJNj96rHPqZW6li7ktKuEkPe/WZVfQvE0gbRGXRv7uMphdPq4+Y/dmKzLiqZqLt3a6ZAe1uBA
GYlgsRjWz/YCgwMt01rUGa9mz+gxFCj82e9WAakWECY9umtida5n2Mr9iIDCryXHR7cP7bA7JGwA
T+qKQwoY36ZF9isfY/ad7SLtJh6aP6aMl3OGquYDRyasUC6TBH9G/Rlh3d0O6cITbCRihYAlpRGv
ZtFQFFMIt5GnjonuGC1J6aZQmF4N6tYoQFaQRnR1/dDyrP9WqLORtDXr7ztsfJmCpu6tcvZNdfjK
4CSbDiTbiTG/McIBrrcSQgy8SWeOF3NgMTk818FYMlO2y+C+XLF+Sgw7THQdTDZ9j1tKGavqBI3X
4E/L6YpJ61Jt4DgiqSek0+BrzjlnrSDRQsybajb985SuiUBtyTnyPidWJn+mFMN+unsRTFg2YRpI
1xoHUim0H8uPQo8w6dD8+K0/ExqnV1RxTwlPhr4pY+TsQhV/6h/nRSwziCxYZ0t7KOcmh7XIYTEd
Uc9bCqUK/oOQ6WdmeN4g46K67h2iX8oM6HY6X9AxR1Z1EjbDaN1l/EHUuSZGPrUSkm+N6D6VWAEo
GQVdM625WlzavcT07oLmhWytU9KMa8TZ+eUCnVIwKIi7m5Bga1ZT8U05kWG6OpcpyvCjiX2cM8ak
xSPyWbbgN0GuI74CMA1xSlHWmHzHOCyR1JUK3JoUvRUPCajE/lkKtKtSS27vI/MBdcSryjFdnLU4
wp3z4xiIKz7oL26xjpCwIXlvSsuh0UKpog/pCiMYW723U+GmyYF/vUMFbzHs0k4De6Pn8VEwzKsz
nRHvNrimilhOYTL/5MW4JmXI3Pe2CRl0wSlSoutzSuga3Nh87+4M6gzeVASKkoVm3VVetA2RdLqA
h7PWVdzQEGzI4aHRK6lZ+okklq5Rz4Py+rxOtptjO3C2r7MxHND4xXzxB9mKTYY0ChgLHhmyWmZT
0CkepILY1oRJ0URnD0l0PsrC6A9CeS4JheC6Md1N5/gUwEi1WkdZ+MTzJ2pia1UpfuYcIRuPaNYW
7cP639HFLeFwMVd1bLkXPPIGi0WnTdHhtsdynX6pc0cjlsKX4kO/E39V4AMg5yitDJ0A461RIXjy
qCiY3Yfv9sD5USyfB2QyIJ6vuhWZ8mqsx9puzxnjriw3mPl//W57gzwSYAIeABlcFOIfGoQ0vS/I
qNE7LudMN+mXckaIpWNANZ/7hF4r0Ox+jwX6DNCQMcMhmihRPgSfeQIosZp7vByp3+Vzv9iJdoEw
zE3mKJyUE389eZHHbcz6Wl5pTBCd5Y/yGRr/taf58eCOw/yNk8X5N7KdYKDgsagjv5Pw3xM62qFV
qK9TT9z6Ll4y93OcFnOsvM7duPQ5wbyMwXJmGTwdXjTHbD+v4pFkmZ62kELdnyqcVv3j+UhxC54t
ukDJR8/MtWIXXTZrCP49Ee3LONxZxX+dY26jIh75mm7XvV61SBVrBt/4wWH0+CGpYkwzos9TZnVM
1VoI3doNz2n8sHwJ4XwtlocTO5jxXecsWHqE+Ejo0B3jFojW7v3b4ExFK0EdaI4lObVYhOMMKQHA
fGJbNeelrNMevpbprkvZ8YKdNr0lUEwwE2EZChSnjEv4G5rIkbtXjgSsq8UEhAOC7UWPs28kQQ0W
UGnVnNFX3c/4i1hdNjeQQOEyf6J+Vwc0fpVGDrPathojYSW2Nxi4byqU5wDx1pjH5y36rp8QzJzv
1WfMBIy4nPpRky5fBLnGumDUXe5HZXIED6tL1ZKIhFT+N7PEcqMVBJzEPOdEp1KcOanr2DHjGoc6
PlY9qsRZcEo2KD5qUzUv9Dm/uEIDDq37NLqtLcYE/E/sVCDKmksF9fyo6Ky0dnDeahD64+hnLMVY
44XCslKSwBW5HW9q91j/IHrXfzGBZ5PH5d96dj40IQt13hN5xx2JcI2R7Y0z5W2ioPuxGj1OjPxw
3EGyFkThJMjMk7kNa51lYrAxZIQzPWDXqTFO5m5LfDDZ97NuGd4RvzIC0r+9Q1tUtMowv+gshVL6
He7vovx0DpwEsl1yQUppRh48Y0GAX74PV6SjNPkFLWWrQRLEAES7DjG7c1LqGxxVqvr7shU3SRfC
dGwerqPo2Pve3UdSXpJhS0DAAWq8mgtF6U/MkbJbyOCWfkDSX4GTWotiKmhjT/b0PRxWfPTMu6c2
nX9IzersILpYhyWreTaJMJE/ZuO8AxSoZYMTloGLiFdG7B91dkQ85I/hh9Vg66c6mkTXayDTRgwY
dxW2V6UXbRoCh8V9pHDPTnWIt/rz+aE0XdrWAbEdfhFeqOFFRYBekMCGovFazdUy6SjQrbXIDcPj
reBvM2gpir7ydsaSHe4kAhNgNWzmMrvDKOUvaywtPRmyyvCtcxzmBPHWrlq9kM9MzyUEuHaWMAPL
oTmjNLqzlPX0CG0uCQKKbhQ8Ns3h0vxhhXCqWv5qD29mblw4+7e3J1Obo8MVk+qbGj79KZcgA3K2
z7UDHCKl61+12V0AH8MTmpnSI23LDy3EPKi+lnQy5pG0POgRrBtaSMR+QzQmj3HJSqJr3bdxrrRO
ksXyMUtpzLaqVIrKvF5rX1n0Weuqu3oRsuB/uX12g+1z3Gft7MD9cFA4UCQajRT6FjEl70ZQygV1
kLt6kCR1RRsmgEZ1TbhFsFQRI7LsPPfw4xZg+5RbzFlkUppiJuoHCUaDcV9wcoxTJMWzbMtENeKu
Y9BIkOqjpRKBjYFslO46XPobp7buJFuRjlYbMHtukCc5ToE221wN4oO3w0v6Ib+mdcDz3i8kTCo1
qxd4Yf1miCgegakqQy7e736I2rpioHrEYTHM1APy/5gRvivbCk/r9LqWHaQnaJE+RrCIeROqri8w
g8NTFhWqp8Epv923LRrrXKeEUUnYjrMrtmVo1krR3yPFFdUW9OrG9MiLrmH11vHq+aD5/DDpU8iD
nEGvaMXZkrslttxsKmFSZybo+3HSiHC9tKlbQX4LVTG2iahP2fkrrU3H3mB0i7kkKbTyF+9XjQ3P
d+EVXYSQbAN7LtxFvJsiZi/F1y0dBO/lO3Fux23Hz/hrN46Ug86kbRd3j3o66xEWIN/zEvEm6xJc
5Baimq4vznRsgO2HgGP64p8GPKBtv1YopUaasKwlamPhwqpUsey2twiuE0R1edqk/VYhB+Z20+RZ
JjYsQGGAg7emrk1D8yYwqb6mv9zq2M4iRu15pquFHJHUIxKxTFXRR/Uj9J3I09+oPDWdRghDubfU
hM6uapAB3GrTov9R5/A6ZaguKWRJxceKjqFb2kF6RdgHcPT3HmQBfYVTpCVurcC4KRJastO5UGBR
w1u9L198HEXXTlS913oeFXsQaBH/mCqk9OoOUbWRtQ0ZLx98n4GIJP1O0C9leaFPmtJDqC8y6MTh
+EVM2FsZp/XVfxjvhjyZsq0y56NnPgGKdGNkEGncATu9YEaDepiSAK1LOWpmctBNtWldbfJfWyxT
3Q/mGLlIhEKhG2bEWPLetmf1UmH151iAhJ7XTsznVvAnmk89tbEFTxJdvVAaaxNzNtvEqrsZXdBK
pK9tV5nArF7j6xgEAhmytQST4xYWkNKGDbZM9PdH8ER/iUdUYUvn9vptxmT/c6b2B1DN2Gw9+xAl
nn0RQpa4kHvle0BKjvi5EdrwrPG3+wWUy6hxn8a1i1RVJ4BK6Mh5UDGXRoiVywhqU1k+Qlg1xlgq
jmj74JwB4DlwrbD1yiCYg2MijhC01z64xSjOj+ZV89BSZk863Oyztg6eLQw+GbrCkX08Mnt5Yc+6
B/bwV+Pds3Cv/Q9E92wKX9We3L4GC6pBu+ELM3mUC5yUeOdjlycHyPvZkHzxJm7T8p9Ch6UugzHf
itZSzt9ARkdC+1fuMXQWiTLZh+TuCnd/e3N3TWmu0RUYiGlGPaI2bYCAASIm6LobyvZB5WARkarH
BULEgJwbnDQN/CVvqxe1ZniPvVdQuyzWr/wPfA5FdYtrC4zF3dZFh0yjxO8K8o0662Q983d3/cVK
FnbZT3iLB6Y3/4EDuB2FpR8GPJzbfczZok8NWDnqDW6vBQk8DLbSxyCntYvBN+MLg3VJ5GUhm9A6
gUk+3097E9SvmJy8SyrsimBIco1sYhxanyzzk1mnCFO/xa6W/qQPOjYidP9dsKzo8roY4UUZ1ZPN
q1eUA5b+dpGtzsV5iCS7v/Ryn60XG911Tck8U6IYBbRuFAdMyMEJKBVCrbvYg64f32MEoq8istCS
qKsHIAyqDIIGadKu2rgkHr+iaeYB9G/HMz9j1BcDr4Y7dI5qIB+lNy/UEfjoGE3pJNVvPzxTS51V
bUFG5Z5cRV+t07ONzjGzNi4hwlLzOcE4F0pU65+JmlqPABFDU8kHSJUFJhj8CfzonCQs3jNiLmFu
N/eXNqUkc9+oXD1OeMN8u1yeY4w8tTh+bcQVrvTOWK4qQDySdNU6I7S+klR/pIluTRyLl663mIVk
q6FY5MzrNCN75wEEBKy1UDLi6w6/pSb0rLcEEEo6DC4hm8sJJLnHCF0L+OultfiugY4lyUVy501B
bEA8bJBC/+GMGe15l+jc6VnzRZ1nx4NvaN44byr3ME5fruYKCTqJi8PPh6oaprbUNyaUkZiR2Q+e
QjI9yeotEfb4ozwlqNPdat1oaW3qvcsLZeXrmB5AbP0/ohRjmU1P3grMrqvxJdzDbI05cl19F+AC
6VenAe76+/szAIMWbHRkfJV8W5l4j4BTAb98PISykhi0M6cWKtlgp8n/vpEkSEZp946lx9QgVcGH
/CkgIy9KWJ2BbCu0TwUbw7n+40ZqC3/TLiA4k88+cOP0cO/wyvSajtdwX54/7G84KU0HZgqzmnaM
DPr3uKTZXshB0lPDrqY7Sptmz24m5s5jQh2btERl3FslQtoxCRYIz5DxHiEq4yLmXITjwiOFCP5t
OX0bWegxOCOGYjvYyJJFWffTtwOtIhhkGsYG8HeAabokC53UT2tPtS9KlvcULfFibiE5ztqoS6hd
r+wB6j3m2Fc5I/koLOKqKZYRn0E6+pg7Kp0MqXTtSo6wkVD0TP/ur2Ep780kqc+Pvcmfl7vs8KKK
PsdlDEAvh0UDC/gUqGVd9T4Yuvajjo3kKd6jxu0IsBJEnWwfD4un90y8YJt/HKS6QC4b+2AGoz4Z
qwfwVS+jkPDswqX3bio3LtJYjwoZw1+GQSGHXuF0XcpuwnQ4r7NYK2k7zQls4/M60YlK3TZbkQCz
C57YY5BzuqfqJdUI2Zt8JrJ09CJ9ZnHvm+kynEPtN+jFLFfWaoonitIjLAeJ033zRSQGmdT9IpAe
MnPKMo0hVVMv27dYsqcXhPHA/BvFY7n0S0vazs2WFL7UhdR1sm9s3QrB/zhdHTckc7ZAjGb9PRxQ
+lRZoyXwCtLtJwYDxXex465i563I9KxKLWAwNEd0E3EqI+Gy7lQYPxOVr/jJ1tWb+TpDVkRERt+D
nW+vnehOdQ3fkn/9pEoAi0uFnEL72D694GuW09fVhcu7tQ0Z24Uh65cLtdeYckmaAdW1NdQbsMqu
lj6fU2wN6V9FecSrvYBWxcTSRv+g5vXO5z2Y8/hjXBLzO2mYYWwnKf+ilfvnK9V5xNbWwv7/rgUM
OLF1jhAlKpAIsUWg7UlJ5Xq8kCGCjlWz28x9QuAfUYK5vHtLTwcmwahzrDkA5wztWoKD7OqaqOt9
viV0fuITZMaluLrbev0b1HAbAT9c2PfpJhBnruQleQBl2sTM8gkUKdU3dLlRbyi7W5GbhblMBSuI
kCTTF/K98DPmt1+j/D5gTe+CBnB2Iw1PsHcGL4CfOllC0r1u5u/S72YYv6fXNNis6okqr0YDkw4F
1OonhW+1aBzgRapcqctaPni1qa8gDjbydtfN6J2pZ5TT8KzQ9388dOXQTTzTMbSjR+Pf6zK+sD6C
KGmPbyNE05xdseNOB1r4QPusErfpCbRvuLDl019ZHXDI0uf3v0RXAqdvYuPI+X3Q+ZQKBFuHYWUh
DIeBWa3s5xMlSEKn3Sj/ZIwaEt0OlLc+8aQBsgfvdyW5HESSli39mpd9ZeF7HxrgFJZmUpP3aJYr
wekxWK3iuPbgi2QoZk0API1Wy8DTzHhUaHK4oqCTh8rKi7/EGafAXdecq8N2FbrjAwyOznaVwNlL
QlkMeFIoeRnIt5usGkhBMbAOxdQGNqkGA6PaH8Dj8O7/qzHi6n5/QvQX3NwVh/ZBPa9ObUFgJ5cA
N3dX2wYJFhzLVhjLSJWo5W4p2AqJcTSKH9/aFKOXIyWZpD7PIAbq21M6mih8wwO3Ul6iygsF3pKS
GV7LheNX3qxERmbyLEv8DuY7hjdbDMaPz88eC2/4PRKyVuAe8umSSZvFcGUjnXFHz5x9A8MTsR8b
E/kZgAniyWCKPdX2W/Mvw+VtM1ebCCKCwcy16rq7OqPGSmrSS97AWepIMxL8Gw2chJHjjGlpv6YE
NlgXrcsLSDjHeGLVheadJn7ELVaUkwlfo+pEAIbQ2FzzUhAKPMHTvSmnjQRWP0xrdsQgWnbq8qdI
0tzYC5F0KvoDWqgjC+/COpeu6Dr8hJN/y+uPYaVqnPFbIHWaUjvSxkeYN6lzX/t0ZuwQ7YQG/yxs
pkRgsnMTIMhX6fz+rUXB80Jfx8RamyUN3VTaOg95HdDfiq/dqxomsiHUTU/98pyBrKbn45wRjJAi
3UNJ8zfID1VBnQh9Mgc3basQJPRnhoHpMbIpu7WJAwH3utP0P22tBYU3M0KEfUbb5WrNwVj3oIlu
+NKniRQ3WG/ag7p91jptINt1p/s+zPrT8uC9Z+Ekcl+19FlzfH/kjpxHT/qdSL9ti/ImJRtHz9hG
kzuKHJmsDfusozK6YZEm+hrkrCHdWpzrkXESkA2/Jq2JjOI/qDg3zRXcbiVYCCrFJ5pzlizTjtOf
CgdJRE88syUOe2VcPeJJUMvfrL5bOX2il+smP3hA84c5GBgDuFLH6tYG2eWAbQUulVgS/SyoL2ZW
x9pZV1XOsHrSze9aeANIeMJLOX5Dogh8UbJg2MyrNwD6Tw7Ibmj2kVFDpBBFOpqfXmZEgXnVqczT
oF6geLbMf7PByl8WvIKyCC5l7gPKwTo0lm8371iKZLUvChm1hDc72B4V3tiHS9zx1hGZazyqAnZv
wI8Z7xYLQNfqxQBkOOuy3ToprF8BIw9U+tjWDj0/814yVhD/WNe6kkGtALku+irPtNhhwvisTGwU
7CGuX8QR5XNbpqenekwhNMMXJcBdpOkSjln3Ki+vTpapntCknZi4Vg2dEqHF+ibXz3zPO6hDtzes
QfXUI1mggTShjPhgE+GfcUgi98DXk2AdD4PjaWvlFvKEQgEooJbkaiKpcpD7Y0SFbMDocoVyp0nn
U64E1cnuInQ2qvIOQL2erq+ZQYkQ5THn29mrDLnt1cAR0RFFhMcO/yRCdDhHaKQDJRWreCF+TyMl
2zqEEkG2pbVgkBuLEdD0sHVoF1kBHLgcGv6Ihx1vux2HPiLiPHEviwJVfUNr+q6cy9BgH+jmxLcP
oNk6rKzcLQC18kezRWArvaJ35IGzcgJ4gCuLiDsmrZXPnvAHUhiwLIbRnXy7jCWT6R6g/dXCfcI7
bd1lieZNhWPDNjiyB0+4Jeool5s+ZFr2xrGFxbqaepBn0+8O7a+tQ1E6OucRRGzfJSLYJc4dNI1N
8PkvLzUrf9xEJ1aCCsWH3/mCP/mGVDLFGb9LG/jjVIaZSnbk64B0nZ/EjX6ebMhkYfQ5O2ot4TTd
RcRYVjpjI6neCxep1GbqdiaPgHSj9Y8hAsL2vNiiDKMiGuAvpLtrwnJIDsQjHtJWf9ygYUW3D6w7
V6ckhXDbDcnZDVxk5RGOX6lQRcYFtTxDSqJn0JDaQEGe/Ge4RV2j97Jo5d/UGdpM4Fe//+xWrpRp
nxJAkW3ea1GAM7fnYbl1jatVMESh5O8iIMsl8EPkrlHI2xjJV5RZUvPa1gwCLH7gBeIrV2PgXrH/
f/DGuiAWarmVT2X3yPxoaFtmJwxT24I9lRV736VsFM/hc01aPI11UG9PdzRkY9J+CHiuULdxCO0s
7ydTdMN4oSaGG7i1bxgIWV5CFtFT3p2O9IawCn+LxFbavvw0j1+m04WXrpo0Az4OHnTThrNjYiVk
3ahVpEo0e9jhRXhwAMwqmA4OH8NT613wArQmzHfAG3BTEjohSfcjTE4EoKhEaPHSlPChkeZ6GvLw
ZLGALJB9WxgOL+E+wz5tCs12R6nJ6985WkRkg13cOxOWjAFeXmHnyrCuJ6yLR47Gg8Q5Ep8GhTW+
2+s3PkXBArFsykhGaliDfM6IUu6w/uKh91S+bHV5gKH/foNpbu1bbsvAtyekeJEcTHBjqzT5409B
/nX+X/spyej44TdPqQtSJVn0NiDIsCxqky3O+BOcDdj7/HDMYDwu2nw7b4lmEN3Rt0Fu54tZfQQb
s0rlfgaGXS4h7P2f56ReBKHws82vFLTu2d//TI7NMPWI5tUtVWapARtgAQ3bVEdVv2oNJ3EraYqp
+ygiXr1KC+q3tQyWhINqX2uAGn87W3jMFKl8QgJqeCBfNkw53cBi1swqWW8UyJj5dICAqeJZ8xwL
74MxpsoCPs+E7bYGgrsYAsHuw2/I4JhmfarWyNPabi77HctLH2P/2b3nsmt3Y16B45QhhNilqDkW
EF8BxVQ7aAZjS0BnovMFgr9ozU9xViVws4reJzd3mRezOoUe06wrYevSInSye28seWtQTLFn9jji
CpocPryUVSrf5hAxsDF/j0ag49m1rDzwesMjo7v8zkwqNXowOC/bKwwwEOXaXcqMDNBtPnMq6UBZ
OKoYKboCFQ/YOrD31GOqo3wbk0V/oSxKMXO4dmXzJ1A7lQJspFnG2uJR4DC4wfU5c7mZ9OKqUFLA
nQAZbK8y7oUFwipmfyTmjzokdtyIWl09FTtvZOavPtzKryyoCLOPp/ij6PUTi1M6rPibIFY98G0M
BpSB0hbJ1uh6+DWoPGrYPJfOnzMbfdaF1w3cyJdxUkV2ym9qJtZF5O5nm6d+Z85nFsetF2nXej2D
TcQIB+VdqwOiE4WxDiZndU2BkIG0Gk3X18cdsHNOOsJ7MbOoWlYeLF01vrozF1pP3mA1moM7JEvh
zn6HII8zA3ugeLFA5TYsAw7G50DRLMC92Rm4kKEjIVcIFXTRz3QuAssqFetCVQZCUse2WhPWoyxX
kSm6Hz9Qwj0FXhAFs/zE9PK9nOZ9h5oWQgmFl479mCycX/9uTqn2Qv8C8pfN64Zr9Gqp9aRub4sJ
0MudiRMMQI7FOxboAJSvkd1QCU5vjKyHcSgcXTMMIoe6ULrDnK5MGcNpEugeJ/4WZ68c6rBspGfy
4H9bN/19vO7GMOyD/DpZlDwwggvntlFiBs3n6mcGyZbQWsSwcimDIGByU4biI3ieqJyKIeC/64rh
eiGQJsTe6vnQhaNyaRX74U9CP6vBJhrX7uNkvgpMWhuroa/TDcGp5FpRFb2CAN1qpTIkajkk0ndD
wbTrSFn87Po/qKRiyc0bMYc4NO9qY69ZKS+xl1nA3Sv9uHH/ZYOKydsAC0pfnyM+wUdqzdaEwXH5
aa8Uv6wjy2dszKMv6YuKi92xe0U3bcZLHZgLUs+8dMfXjUGMmpPSaUYIdTtbJ3gdO8TgC+7hEyu7
pwinSXkhuAs08L9lJwzzmniVANoQ84dGKwE/5QDIcDs406H5ZcqY3ZbHCV/xXXrmKnwCiLea4X8Y
1wnnoU66LUTE76bYwoFiNJcISEcgf9PfEnzZUUrmBSDOWlh+Pa79x7p43HoHhVKLhKmpzPkCW56h
8mVDNvCA/SYY/KQGMSjlQY0a1G55TRRfCYQfutynAbIItCp1kB0+vOLw1tdELXb7mYULW97p5xot
dYRZbo/zCuVNxXO1a9LR9e6PdyQ/tfu3gRLrGfyjG2+QuqTv7hcg8qzOnvXg0OIf16NIebJxeANs
F2wqsSicugHyeivofT05IkERtaaCWeoN5CYVwM+AO7SULIuVkaS1ctnGLkxyJKtPelAAvv8GxzCN
0vFDJj/gndRHTkWe7X0LInGMyDbDtGh/zi58TMtovuuPRhKLARRYH3xtHSghpE87cUSoS7uzY8J3
4CBQtCjHVeuJNgWx4W6h/cEFDFyQF6QzQQlYyioQdG6sikKWLQwDhVOB1I5SYhk7gRRyrUWdG6dw
fO4QHE5qbcb+1BOCZy6W6f2WrS37R3jNoiGWDqpC2S3Xnbk0opnzMItwqxXJWeklpcVdjGuiPzVH
vxZap16cEocbNHOuj27KM1A7BD/eRXytzxcqqjcULzdclMpLzlQUEC2fi7cuF+pYsnKg6sGd2fyu
Y/Ab+UDkMwkDuOwhBeMn4aIgM0Rp598WgKwhqLNe6UNm9NtSk7jcTBVcA/qcBHIafig4ncQsu1Or
1a52LkZk4VJR0qgvORleSgbLILyn0wWarcnOoKsKBLeKteM1X0EIBWSZl4ReAtefYywMp1fhYSSN
y0naNg2itCmsdxmo3E67GkOBm5SIS40joAe99PU2JpnPejuUwmYmeW6lkdamTZavhhNiinWIRrjO
IYK95cdpBKXocr3PDFubFc+Za887TEwrlBmSQ13VdHY8z8J7E/vboSVUzNn6uOgj02GXOX2sFePU
zriyzHRePta4D5bq5kOGJeJ8DIIzWIwUUJnj2aOzVlllpy4R1bw9uWmq0Oh0bmjmREvj1Rljouuc
C61L84koL1zm5RzJ672N6J0vGBKLdAnw+7l5ucrBQgw7ZlfnyQRGKUX5auPBwXWcTbFsDJgL9vxv
uA/zMCoi6G38K+N1+Py1cKel8L/eamLbRKo+/FARxqLluJjs76Qr+vqWeiN4tItIrPAH0e9JYrFY
w8BLai+DRKBquc7pPKKZUqohZ80JmTDYdXTfZega7OKhK9Wh50iTh+vNaNPjeBAarcwY9xeSF+2m
OcFweoCEaI5C6VKKhkB00eWT63XoMPt5SDlrO9/1kpfC57cSRhds9RkkCn/QvU4qwXTSjhXGdRmi
TmB7YW5gUJuDdCrHtaFayEbAax/qgfF4MWKA64NGpb/FeBQt8szJVNN/T7rnn7j0Vt5f8frvof3r
yCHz6TYQh2LBb2JrdA0hEU5rurDEOiZ0d1i6aonqqSfYsidUgVHT9MNJrzXmL+jCLdqOCodDsm3A
apC3wNqlUksL7VuNfpdqGHLyMBJaq5UgJu3w0LBwAr/Qi+Z8X+m5kiulgEPIAyW9lfSVIn4FMmjn
ZTBh48jx2FK5vhNhuY088rx4q+3JubWymRetIhzUfPu0zv5k+JzUCg5tlBifR4dyFgOiiDlFxbIN
cmvkhZrIubfmiZt3DwPKD+P+2yKGeP60sPt8wjZNTX9AXYB5klujMGugnP5UDt7x7RLUExQKB/0k
YhLVvke7NRq444NislwV1dX+aFbHKOk+9dWZrDQt3olHza8DF6YDW3ZEyQujPamPmWfMuHuYhz4y
40gFaN69Tx+xPTHQpRDa5Hm1ZgF0/pig6NKcN0ZawUu2pY8oArFSbYX6ypQ2dcUqVUBM6NRUn+L2
3RQFpW5/EwXr4br/Kb8NTG+NzngniZ5C6sKw9WpWefAmz5ajAqRRrS0/IXKybPSwTarYlFkogPU3
Qcv6jHO4fuYiCefrN3rdgjNPJxpY0QBKU+6dErHh8Kx+veeFvn8l1eV+wZ1lZrwQVaJGbi9vQZzl
bnLaQtTLkGG8o88jlAXEFIBwH82GxPAaQj35xwcMV0Q+p8INAlkgAZ6tiEo8PrtNtqmuN+/fVTcJ
kavIP6kr3cfBZ5lr7Eiln8oSE/30SrvDYxgs0atYFgNcMgNxwBj4FmxMhqputDfBzNqn8ebE2n+x
2fUa6pBfoC3bH80amDtiep7UDWZfJlWxkd+9FfADUDHUyLesn4eHPqSEl/QHaavCjfLmYqccq8Vo
ksN9k0P8dT0F9rdfateMmaHftR0K1E3Wd2O7l5vyQvqyKSfjXHfuhGBWRwDuC6bfsBTjSvuPr1WL
P/RQNb1pKJao5h7oxTjE7Ik6u8DMlWHbPB+AXIePWTJM740OYDhL/NfvhPx8h2ixd+N+CXP8Wb4k
3mPT+hsJtfv0cQj53BJ8O+uFfE6Q/ECxWRofTSC1hPflvPGle1HF/vvLgJ1N+EOK0Gf3n+hqWTjG
g1HecbbpFMXy3Fc3V3ReV669IOBsNRV2WckBcURltnve/Qp7J4+ITZCnKPAlKPT17lVpqlD6U6dI
7Dx/X10wX8zQlEjtam75E/FoCB+VIsLAWhfUWtAMFiDR11ceM0GV2FHEca9bxIC+83xFugMeqY6U
gQLUMDTTkAI//BIPtiyFl7+l4hh7WgrrFlQhfZLFklixBMoYpkVPZnujmDDDb73lr3pZBfL4kbF4
HJWcbMcvWWPTs4uMYbav3WgaMzEnnMBTFKaKqxCaAT8/N/a+7oyAUkCYEHE1KgCnqv0lsI47Qrm5
GObycUJT5p1ZxREHFjwVI86dXA7h1iP4PlVuqxMrDUERBLaMsGG7A9rPB7bAtTwQx3y5NhMERhTv
N0GFJN6sZrbgmcVXYyxe3dDH3sssKZzfhLWmntb/lsokXmzGvpdznxqrm+dPiqMUHncXCfwjLt/R
wjzCh8cIr7aPppggGH/tTrUr2CbiyUra30eo8qZcBhoH3iuCmnxQ2DyFtr5YhT38BBSLP2vPXK45
ICdr8UUOc0DWe+sYctoIgrjvHdD5RyUkUm7D72ICdxd1+GWpYq4hOceBdblb7WGckxxwwTbLf/U5
HDmmyCCA8KZD5AIwIbsQovfzLTg2yScKlBgs41H4BWZDkX3nHc6ihPBlQQAA54SU/48cRC7yJa2F
fzM15qcCn+045UW9w744lbiYWtXcqCoYIYKF36BJSDpCz8CJAUi+zBjWalHdH025fr8HeeipzrwW
XD8cmlzsC+IVZ3pIvP7ORRUo8DOsaNp+s3B+VjJ+1oKR3/6QLcTR4aQAxLrgdp1icIqXGXOTQEfr
18kWGHn9zco2PsLo7nFdPbYbL1wMr/KSLjARqrnu/8gBw4ccOKVeL8ubLuw32pfice8lsPtYDqDt
nwAtEt7+1pMomMMTZGTelY/ltW991x5Xi3equ7DdauOHVGYttRUCNqK33chWxpdz1ZtSWsV+mD8y
rhwrIjQetiOCU0EGoM9U4YBhknGC5T7EJKcybAGyINsUMwaYYUoGGon0c6O2qKGne/un63ufRXn2
eoxpDeND+m6OIF8MLV2gXHWXEFYULIWO5vIVEqw1XlnnPJRwLthkDov2QJ7hYGyZ7f+yqUFJ6Rt9
HgOEEdCLv999od6XHA+WV7zRI3M2DaFrDHAdYdLPOlxf8P+5IBIY4ZjKtnf8r3HGnORBnzy+0zlF
dVqTqPssiv57DfSgllWzPz6xJPK+IgNR9C2YTBnv+nOHlNzx1ELXzLnEQriS0BZ64kDjZtqCuhta
6D3XJH7a0jLbM4I+y2llbyNVV1Mog7DTWLIzAyx86p7/ny9W1/q4XdopNMij3RSNjm3bID4kvYpc
+wuLLIlo6iOFp+7our0st8+FkhD+D695EogB3+syZ4k2XixkKbmlpT0ctN16+CkYOJUaBnOEYZru
AzXGWWWEbMTd6hAe4aPNlO/KXVkiMpMEMok5L4USRyRR4DGlnC2453t+q198wqWas0eZTFp9o3KU
aaDykETWl3whWiJrVgah3OK7jRO8swin8axqBvjg5/LHqfmZGcXlwBSq0fhvaD4kjvlR/fCvNXHm
7PfdcV/xr30TV8WyN8cq9qWyUEzapzW3FDDrdZ04+g/eOLSpGEMSK2G1j3oIK8/ytyuU5hYVx64M
+12Hz36v21zkl3PgCIcWM5R5g3uHBTv13lLcHGonzPcMijrdc5SX7zNSIyqQYMTN02B8o7A11Caz
pA3ISKa4eiWM6WPc76DulNnzX1c1PCUGVB04yMjutMK9vEHBgG3+aAOLXMQL4zTprXGrzzNgqhDT
ghBZ4/i8rCTc0YATmA49lRyJnhri4jm8SZ3JjHv+oV1YEqC9V2mTvBQKz/0SBjcoUQAD8Pbpm9qa
FU1MBgEVJ0ueed6Slz+jYrUxmc6FN4g7B0dXptDeSPfNpDkJfRGcMr0lj1BpYlOOcKEeiQ8UlxfA
zJBCyJULtCasp4jRb62YKavomk75Trbgw6ocb7HOcLQxH0iTciDvtFnxzJqJ5cCDGTxKbwHhbim3
+da2rmvgEX+Ue4L3nft5uD0eKg1c+fYUw+Pku9cYYWo04MkQIOtSu2DrB518iXM9NrsEYypqdqA5
RTh5dFH4dp9ydDjBO6TztcYEJLhynaXYZq87s4u/uNvpR54UJP5RHWpf3MdIwkraKejQLldUwPXw
YBjeJ4ISTbreKIaO3TlSVoEDNUalGcAKn+faYwQ1ISAeML0L0Lhj8lSsvGSJpppTJETIqrpRo1dZ
/xYK6SyJAQJpjTUsiwHjxOvcw2Lqlh7MSgHNL46tHwhsXMVYMkbgSZqkNkA4ZhdEIc4S1HVwgrmu
zOlqXXLb3PAJ4CDF6VGNutxVp69cw0CY+2cnPctK/COjSJg/uUACFJg6ww2mfC0gLEkYjdXAuCDA
wt6hqP2xfCQe5TQFSDW+kpuBNhmWzHweaK/C51D7XZWI3J9OMKiWkj9OejUg3lMmksndZaqi2zpr
UDId0YXzLm+f1xJmtH/sjxxrRbrsxk5JDda9+4CUeT88gKx6JxMIaE1P1pEFHeDk6xs41IKX343N
GhN3XJMzluCeEdf2JOxN0MbsMbXEcPoKIIDBnvxEKzJF8lFRMdWBhZRhExpT4EnZWI3GCyHVx2c+
nXcxzzddanybUW3SzkrSE8ffl+hh5dutQ/JsR4dshouOXmv0EZK3CuPCpQvg/aoswXzCiFbNv8Xn
snF/5Mf6luI+bdIarJoL64zP1sbqlU6kQlX/6p+oBJ9z8GamM160cVpzTZu5saT1a7m/ozHEmyxE
uZMnjouCSxkBR5B85FLLrxcN0bFHtHsvPcENngmZJfnRJtt+Aldqpnd/YKtzH7T5kPrA3cFd2GFT
uWPU5BvnjxwrR6tdWvgUPFERPXP9bjgQxj4PpHnvhc8eXOSGBUW5bl+Q8CZ8dQHQeJ+9tTsBf+Lu
aG99VHs9qqQO4/OMa3pwkHqscHOXWJQvG22ECmcWB3gheT5a3+g/bEagJjJT4zIUJnFNac0SBcbM
77JvVCdy/xPYehmlI2bFTOPFChXyI7tf12T6Nj6HqkXPHY94hgYB7iYvgMW2MFa350nN/SP8Cgik
lVLuhoG+Bs3XsDVg9HG2R0UaBODh9Wx5PrJrVoh7YQtRa1EK7CGkG45QCfbDG6kXwyok2+p6wmBw
n0ZMqrUDKkwqf/7sTAKZdWPtibXY+zfpaS8jJ8kE4ac75gjNaS5RIdwaYHd7giZC2MJJtdEyY6K4
aCzV3HiFYssxhV7WJq8kkBZfoYlhzaepoTR2b822zNSwWuazKvJtUTHn4i28Xmczlx9HSCW0wnnH
LVo2P+BCCIergqqjPyHn46vvXX8hJhRFDaBtkFEf6kbu+EIywiQv9IK0AdMpSjWQM9qNaNBpg4Y/
gApb+Jt+EzwpNKjHUrDt151pFgAqAqUUQdrb6GELwsQepbN89XtDRLA6kD3azXI3HyQKotUlPsOK
IpYtDCUGKrKHijuuT7Lbtiz8dg5Ux2dkK5Hk+NlIzag54cpWAg3ZrSM1HdLpv9fKqDCdcQdyqrh1
417DY3qEfE5Aj5PirJUJaEUq/w+TFInZu2OSQ/SzY7t1c9t++iNn2st96ZiPs5QHERJJB6XS/K+x
TlueJtmyStyks5wBoAjDVnizHEqhGSH7K33F5tGHMWh/0KZlqx8c5HaqXwTh+hB9w/V2FkUMREcP
ySyNR9jH+cJQEF4NcaEiFuefrd7qeQam3/CX5kOq2y26zJLBSR+EtZ6l9XpISJSYMTZnLzOyx00U
myQ2RDdQTmCWDfumxDKaevb4DEyjpe60qOicRcuyUxoum19lh6Pizoz8U0kiPGV51d1WMn3kI0Pa
VQNjz3/Uh/swe/snfMvHNHyuZXdkz6HrgZQZnKLtuOknhfxjfMDisSA29jD48bxBtTFnAIfO3e1c
75M9dSt3dyZUJLNm8ZobeEIrk/U5WS2KH8bq37mSuxpy6lj5PoyCVOFL/H6MhIBoDBnQ5Qzzow9H
/RkI95BIZuV3/WKjVpAUa913+dpIZfqu6woOMXMxdaIUIlgjMlHOMLaBQvwyu6LuTRntCmDvfE1u
B7KpjL3amSHAGDdxmC0EPyCIRLZoHVrIyS5ZtF0Q7DIXXnUxs24QqvWgxeP1nUT56RS4pt9Hzbcu
5Qy70cYJuBizVutLwCoFrSPIF1GJlrUc5I6ktzqPtL0GI18OGribqrIfjvtq9gccsfWdgDS+K1uk
lnq4xIO/US7KqLnWs5xQJP5bNJn3O/5oT5W4aHEBt6eJ3+baBH03HytRjcldaT9jgKKytHB0sa6c
Pux6Hd78xHxT8oHQIWJal60vKdiESaR1UeCRnS6t6NmgAVZR8BIt/WAdAYdNrlYcungbBQJnFFMg
F/mmLNz3Dp6Bes2x4Wvmh/emlR5B8hQBzu+7nGHFwOM+N5W8wTJdLJ2fKTFxILgNh4Hq4CbXgHxL
3e+R2SfFcpSP2AoLf1z12GZWf9UY2ledqhB8F1wGqzYol3qx228h1hiLgupk3xeTh5QOJU83UAJk
luixcng45Y/YSmLdc+vV37MZJKtsQTKkQmk4BDwrFAwAJPB6RipIl30IePzw03NhthIfpuHJzf+f
M81HKnkPio1Kw7bvEYMEoplBfxcfOhNRRk41imXAwlk5OVGRGBgphXjuGmDEas5ycaKRhQdhMnsD
iXUv40BKO+bK5w/LbgGJDfwNjgzFNWDYpU/wRl47bErMUgWY+kKzY1Z4Fbzvo3mZfv0Z8h4V1RrU
FnMm8NqmJOBABr9zUz1NMgxFqs5SlyLLZsnRstBS24N+XYqfV8SJwjIu7gcUOIc5YD4PvO0z7ijI
7lCjGY+aDV6XgAKlIQOSz1AjSOmK3DqxoKx/SHOiDofrwzyWq7BypGPWOyt/+niGDx8DBAQ7JygP
16yULYFHy5Rd26Bsdg82Dqiq7PO28pCxUnjOzevivr20YsX8NTHqwk/LpixJD6iYt5hfGfW8YmIn
wh9V0nrkxC69ocHBJNbhjBeepth2IuvXB0heh+/JR/FgNbHnWTO9pNT+0gQH7dK6/eTD0uqWUZxZ
UCkaGmHJNgHZlQ/uzU/xIr2eUFVVwQbECXM7gZGoSnVZsLafxsmLCwvwDSRChIqqmry8mi/CVTbB
cl1u1uQdT2g8X2QYlSkFEtTWDAV7QWe87MPWYKm3Jwm38zuVZk2XpIQjacl9OuWaSiTLy54QM+E4
2Skgsn4jngKL9su7nAO56hSwVFa/NVtmqLD9/2AEWpimX81PSuqycREHAVvSSsc+Ag8JjQUiJeMf
wJb3Ax+B4319Tpr6aQGLeg6H2oqK2AEse8zFRaL02FnKQtSGR037i6xUomdjNJU3oPK8kEQwdsVn
z3ebo8tSTsfvPJNnLZxMBNq64S/VHNrZDbgfzZ7p6tcwhWbO71ZlfMEHbmCzJjwrUX66ZmBxHmUj
tU5YHsF9NllVKwEylrEHeMWZRJG3I+w5IK5/cXZurx+IIDVSEZEChSSMX7i15P0KePgvX/30UfMZ
D/+qcClu1vsP9yF3mZbwNZlkp613HcxrzsSPdBf3Tuo1SIQpnNAy6mUjiYjfbHD/z4SKwontGUZH
7jsP4RoMFShfe+8yU+YuzslzaQSnrtS74S0EJpnVIkXsX1avb5rj9btmEYlvmyhPgAI1E0kk959R
uTqNi9bpsuyqEHsR4p8KGhUpmgqHqhwMOe0OeYooEuaqpKFBkk8h259IbF8f5sOfS1uzfBTzknwn
B9h4WfE1il/E9Ocu4gz/5VlPBbnaI0Zcfb2Xoi9+TxJXwC4daW/QYvs6+DULm/fzyoIyUR6l1Exp
tJ6bBOWH4KmVhVPhhl8WR9BouZ0+x2cUhanU7HBKSajQAk7akcst808+fxVJg4V8+BiCSNDMQ6sp
VrpZgkK9LIKOOTQODK8PsAicyE1FSU7pgNLOg41f+XGIRLWcNBJrm3Z2i2UEcaAqoXKR6Y4rpgaK
U3sEcxiuSu/Dnx3Cc4J8WIVHt0M7vzyod8lAmR/BMLmmEq/fQLC/tdi36ngW4H9t5wQsek60tStw
gDIj0Q3W83LuETjLDyMyBb3QcOvm0QGQiFoFH0lW3CyotzlpAGmLX+BkM7nXptNqr2LnKWkJPxw2
ZCLxrLoP46Tm1vx/KtYvIrqVzrwiLdmJIlKteQHus6bmNgp4HfQa9GrwflPP3CUJZGy/7UcCxEv3
butQtRf22VWhPJ6iIm6ruOJ1UsLzE811nxD7SG4J/3GsLd4IqLL6WbTs8AvQxTufYe256zadT3FM
lEEh+DVYR5Cll3OC2Ttj+ieLjd8VrfbDLwO/eBY50ZAAg542uyXc5zTL8Clqb7aZrkGnl2DHd+qm
OlRHTWHZxB/eyfU5ekJXBcqH/pqF7uZpFrecj2YfjnXpBkSjOzLZvKuNJz20ZuoFFJDFKq1S5nuC
wr6IaKBWCzqVnz8nLjK5TsMG4Ac4f7UX4AOc0EuD+24GKnJRgsBifnfwtt5mqjOZCSZQUnFjXn6F
faMzzgBZAcIdQaKUj5c6YeL15hsMvuhXwVZjyOCfYDdBV1Bz7Gwjh+atkRur5bdddvjsWSuAO2G9
lEaldZ1Ckse3U5K/oYG2G+a29FPEAbcgT36F0lNQ3Ah9xBb/ia9RdWpgbbq5bpUMWQ4ge4uuxmtc
KcGj5cjXAZ5BkAinWM/iSYiWxNnAdSGV7dDiRr54QcyCx64WJOLIg7tAdnixxNPCAtsvEGAhSk+9
uzV4l4/Ph5zhqCUz68TopdlcMiZP8f1sPVx3Lavdl6BS5koOtj8/NTjauAMX0VTLX2BQjzp7h+7K
VL5Vahoz+fYLqJYweg+MOYw+MsUw4Ra2dPTXWH2+PbAe1SYc5jrjkqkqKSslbQMbw9WeaGJtS4h8
WtRzpK7EFSGD11HgFzAlyKJbnOAeCGT91JiOoz2FU5zifnvWa6X3vTd/kZKpib4mC9rY0oROBUsU
m+weHcjviAyhHgM2Q91+0P9tbMXVu/KBquXb4T2f/p3DXv8b/5qkGjgN7JDQYnRqeCY2LBMSqQbO
eFFqmhEQKPYsl+Cb87DkzWuAmnWfyjWL67QHOXAsyucTbpGV0Bor+FIttAebDM+bFkny2i5xZLsO
WbyYKWSFXWZin+cRJ5ABALQDS7zJ9q7b0c+KO32hxXFAs0M664SV3jUs8P5J3WGVcSuzIjaXh4s/
lQzsT538uTg5lbQDRo8eYo/raXuWKme3J/yL940Ar21j/afC1TmBKPw+exVsHf/5KH4Qzeo00SGl
qh9p1ChzhtMySOUcgmNusVBURbPyO0wAbekFfUgdt/5b/mqpnqrY52Eh5mLdccjSfpArjepaxAuZ
0wgA1OnESYI1N7i+81rTOvt5tW7zCr+fWX8yXAFXD1zkq1kaC9ZPOy5GX5yJbCPiLAdmQsUdbi6H
qdK0oGLuttrhECOIe6eyW/H7bPvec4wTpSbgknMOk1A9dGVnpxXIIisJCoRZnmOcj3pmHsuNAlHe
o7uSFWNFltcQlKzamByVz57UnTQGFNSYc4A+c53O2GMV/Au9z3PhHEIzMoMYzL4HIACYvv9lTFOm
LXuFSOFOtkMj8k5RIEsWMgmCnlSdfqJTzhPLWH/7dXr4gSsti/0b1mk4WCXbxprElgXA1ATI5Njl
lzKSh8Ovx9hLtmbHrQnSN2ngZi/rdnrdymbX3AuRcvMwRd16KR+RFEDIdBu0/IQdKTDFf5Vg3jaX
BaI/mUL1VsBDNhLnXqBYZ+qNNS+gIHxGHmhXxivva0EzQ2PVt/OW5FkEHnJCfSsb7RxbzRe7CyqC
CE8sSrzN0Kz17OIO9ybD/XmDHl7mpmNRgwouDM4AHGv52NMgXJlY74nBvqLQ1b9OCr/pKybf1I2F
E+p2sbPUjfpVHpLSAb8c8AgSjuPMOP9LSO81gS+JNO2zyUOg+Wskxi2/4/7aus0GQLcZMjgN5Snf
6qFW+4DQaLR1hg+TQrpyaMGLwGE1vU9Kg56KHx4m9FPlSCiyc/pLsonyjI8DUUTyLn5XjHu5lcAW
ZOM4v4DSKjSuAA6W3SExKCpqdRrLu4AxMRoCRJiSfC/5wAApNjnir5sFYcgn5h1oq4dJ22tSINvY
bJpwfmLWzyhFt0vbaGlZLppChcKvnMUpfH4GVoHCUvzxOtb7TxIrR0wUBIOaJK8uxbn9mhtHUjdN
7EII/75SnQ8Dws2/7s4sVwjOCELb5V64Hjrtg0LYlgZNYwdaUupLjqR0VB8N5XDnLj6yiM2DI+Wn
WiJBLWQssurerSMIcB3lmYqgmjaW/nQO4Tjn+kopG+3i7TX2KMaSKbzUjdBcDdJHAQ0MuijnoXx0
3Xk5l+/ALzINCdAyPJKKMWkHfCpC53cFPQG7jZQIpnjqgILM/ujaVSQhltVWLAwx6/MOyu4i2QjW
d5zB6lRUm2+jK//8wjFkg/AovAxCpCnl6NVIR9Ze8WmDaPKbcgwwzWf6vEVe1Swfi2EGx/+XoEMI
9kckbigLli4ioGhkySHtuCZUO+nSIHHfNvT3MdsCt/YpxqwL/jQMgz6u8zdgWwD8g/GN7qP4pcZo
CiieE5Drf0pbfsDi4uySsujPAJG1UDpndcFqAaOrLPzmRa20EU4P5KVHXLZt4VfqaT80vvwtrO1W
HfjnLMMm1zgKLbaB2rOFwx8t0YNEZRDlNQgq0ab2srCEafMn3EVHgeipfDfcH2JqXaslmh+y7T90
iN40sCnO/PlXQ+Vq8F5Z0f2+ejoNueyYOSSwBrnKjDcC0Tn7Ek/h+ARkMVsaF/wYz9My9NKry3aB
7DAqMDcsO/eG3wY61vf7psCGWAJcgMG5rz8llmb4nThl6wXyfJ/MC4RqlEK6kAKG0yl25Duf9NVd
jZTftdubKhKvQlIUFE2AbbZVBAnLEdzguD61lVQ7K3YlFJEDfRv689dXzA5+cYM13E0rV4yPuht1
DEsJf6XyLxZfKwcrgpCmMYsLajM8YXUyyw59pNI2M1xRz2szy5PFN97B9EB3b1V2kQsb9opjLHdW
HAwn4abLmR9Vt49gDoiSJySlfyr4Ig3BcKWocc0aEX7MHZbkJ4IBRfzAgVCw7p9aUxrxKreF3BYk
huO3MwcoGs5sWGKTH9Pf97bArHzLUUKO7NBeyJAyIQ0mSqKJOQFKmmT3t3wy0xwTiryhc5NKW+aX
RoW4lSibTPYzJJUAnrklccKNOBwe3L7bwEDLEeH2BSgy/CGXjWMUjJIKwwNNLULs6ufd1QEyk8uk
pX+6bEzl1ibwwV06AzqPnwPNhuRzl7nguDPQFglr756lm8zB2ruRfupKfEw9iiKAIvjB1XO/nrR7
AepbFwSUztw2UsBN7qyDwiMrjsbSDbHjl5zJ3jlQP1bTLfac23QksDcrkx5LLFZ0jlaeU6UWm4ID
f2rkjbnDjs08lla0I27MMlvMF0exq+GFZQxBVilKTqL1JVBbkR53dljYFTtcyygI97DJ3EgTIylN
XyufQ+wvUJk/xCF0hj/PqDoRCIP16C086uQjn5T6mouyNRBQMMeJ35MvgNIVLLdvdhTISKk/vKnM
lwW+s3NeKgeAcd8uC5AVWmlt0aGAZVUkzGosLabEP7pvYv8bpkIXwY3fPOZauYIZkPl9sQ2y8NVo
RvCvSg+q4MQX/yFcVBxf4hMR0xYyo0XZfZrwrRFjvEup6SebHE4QRfthi+arckyVtOJHbXDKk///
zuaabw5kAOTfoHP3Dsc1qAMViqQhjtDpAOrmPb4piJnfHqvZqMbyV3mCFvJDgyERox1q/ahE+3Ds
kgcATTgfZxFo++U6S4qW4ufqnETzXJQK1FEdFsNVtBNEXpDLMe0sZCZq7r4/xgMiVtozOqBkRE6o
e6X8P8RU5BbVboTkDtANEijw0RBSNxuXrh7hCZUaZT0JC39G7aMAF4GHyokPDZnu+ZIemHPnxIdy
uzNSgXq0qljlXUKM0xzBif0+JcUmxvmCt0S4W3ic1QeVOw0SIjX9ooXtyewqsQ0nDHnJZL1OFh/O
mZuEStZ8krWCiu9rQlGIpN4GU6EbBjpTfX9H4XZPPMfQn3px9Q9GQ/qEVPOXyQuueSPsvrmhpSCT
9eLQUL8MpLxTnREgfqA8yuJ0MdA0eHtDGlDF5cmZrcBRioX3Uht9kAPmC7Y/3zB4cKBwTNyIfmXv
x87oRO6y6IuLhOK5dHrgbeEQC6sIN0n7HSTfkv71I5ZfVNSscVTeP6eZ37laTe3t/S8JYMZVQsbJ
x6tNP6HwrbMO+9RfMwa6kBKfK52mHszYivCkj12OPmh6jpGR016BMkSZ0HUFYh1ylP72FhjLkdre
mCdfOY/dTBo98Vy2OdMS5KTTGu5BnpPRYX+J6IdjVBCpv4B7R1P0FHj0tSRaATAISzSH5QPIdyx/
EaxImcwu/o+uUi4unyYKM4bcfCeDZcy/0WbQKoHMexm3tj696MHryPhBzxM6x7eEewBHEUQZF+i7
9GtOIe8F6aOMnJhScdS/O1zpOSZfzvNVMp4PdLpir71A6nWtPaHb0A0PPtMCdgfaFSWoqaD0x3H6
vcyiJkSpPIFHA/0eLKd8D1FRyi3ULQbij0YaLriSrL7eb4F4kJPAYVG9BW8SxHdxRjW/mAp3QyP0
ng0ERMovBtcWUQJ8FMMAL39x0aQ6Ms1N6clmvvuqcgKZgcUwwHdit4q2HZM1g0R6McWf46Xy1OWm
7tlwR9g52LD68/PKafreThGtKFrl/nknDgZXnMHYwaEz2DKabu2cGCR+Uq6XY3HCxBLtwjZlxblt
tt6sdZFH7WH10isw1t/8h+hrCYm24Lw1UGOozyjP8dM1p0XnZmzXiMXf+FdkC3emKgI9ONDuB7xf
ppzu5BM2/DgL8eflyu/Au4FR3xQV4KsiXIVUHVfY3Qaj1lp1/FB3wisZhTYYz2o4Fhu3PHUk2uzK
vB5fNINmAZgsUVL2w6peGowADceFjzjd+ti+lMePzEpqNuHPYPToFnM3dLJmVVBM6wC5t99Ywve9
J7PGGqgNxZiQ/lDSoRqtxn5AewblxQdYQr9sq3tjdrx5ahKVwRPiTCcNNNCVC04BD/7hsjLums50
cbO6LUmnNSObcmmSMrk5THg4EdSzuyKP9mewi1YO/+a31SH+3g5kRh+AADYdzgCKPRHHtFWi3vsR
ArXgv9O56lOGn5UIV0espYM/xtlrthodc4wCBJ6D4LwnMpY/jfqG1JHRLD62uAxaeaLI8nJcx1vc
sygXsRqloyZUM4WAfxXrHA4brgeauUcqVbiWXAlEvTHoovuFqUzDFx9JZZRVc6yboncMJxH1V9cf
JKYPIajJgIjy5hkYJh75LnVLgkLgjYVxFffAC2tMFu91p4nD8sAGexzQa3I3z29zIgQdsbk/woHX
YwXz255qIVGX/VmWmje7Xcmnu7GKGFqkYGMfq5ZMpoOPxIj35JcA3TxifbVArpSmJ+7tFEk8pfH9
FqcbVWDz4MBsb1Sf8AHTHYqIuw1QH4ZKCn9mYWRuxT2Fgta2fEP0QtJZfBfle0g4SGxUcfPjrg0V
ThYM5pkEqvqFkmZD/LuKzEVsXhk0HMJyXpb4WL/qrsM4N5O+1Ea4rHHeY78pO5T78tfiN2JomBMi
Bw7/09zXiO/Az+Op/UO81jSAPGYLkJLfjfRGBkr+5e1H1ABwsTL3mRxTh9FBWvUbQVxra3VS3wDc
LXlCjsv0umbuzvuX1kZltlxtlaFI8xeQfsaJ4qteYd1ZrPisamYXu8ZSXTAuLmVZIOYXrx2Sv3Pw
RYWLHFl8LDNAFi0O4Lk0gkeokTY1v7Fj40KQ+KyzXLWZoJBft704a02bnFvY8ANZME7WZiWL+aNF
1DZn4wpyIRQzvwUjdt5TpJCov0ku0YlbBynLmbf5plOGaeQe8oIDZFLz8kunDTq2VR8k+47iBCuX
ScjM5z4jk4/QOfKKzeTFZZj+eyG4tEaeBX6LwZ0NqgWYZ7tusxNPHh5QLTWGcncqK/JcdjEN1E9M
0J2mR7Hvhw3QSRI0x0qYymibevOLAIieeDaDWkmFsPkojXm5NcJmoL000cNfXUIL8//5evbjTOVF
/sw7Rz+YpxTuoDmDqdvKhvL9JnW2fNBSDYZtttA5TroTxLE00LukveAZRuskpiHx0dBkXcRPvanH
4sWp/HPNVb7sKMAzers/cDsLUdqF1hOFM89zgFn6YqkdevywQXC5asrA+8p15sIqUfx2BI5/ZzGE
J+6EYj8Zms10eS8LgimVQk8P6A2wy5cYbpL5QWwX/MICsgsw7a25bJw7Xkvp+3KTlERUwwzmbe0C
p9/s33mGOa8V4kocH0XluAe+k+BVEnWJMiZusNryqByDD79kXNG7Shd5hxeyWb/rdomuR516pd/K
+h5LYWYXbvstc2XOYzeWHkgjDKns6mxZDHyDOKyNIaJhqGuCaOjvQpbusO9jdbYCCjL2xybeCtTX
ZctycTZ9ihOx3050KQFhbrBRk/fA80IMUOX+B8HX9De/ZUN1phVyjwvf/4vSAfu5aLr9LnFd1DeQ
pNucnWMqFcNVW6EIFMkMkrxXc0didS6XDeDMHkXWpFl+8pM+GYeBWIettD7IQ3H66rKHbFnSAcbZ
vOYwhhmNVqaXjfvOF7y0twdOxA7isP0sUQWc5nuaoqo5SmdTXJ6XC2DZ12MuNCsOTXvgzqQ16PN7
xtOMjvBvJ0wqf9MgKw0Jg3dmLCfm4zGiOV+BXq+OAUWlNeiLgb48Ot5X3NSsc49sizQM9aKFfUSk
MzICQFwgJntKl7N0sgmnnhYUejKjBs1zGbwinHTp8YZzCvkB4BnXBqk3+ezUo4m0JRMf8VEkqWT3
F5ezbbWQ5kWLjv7PQk1BvvE6+F+k5wUOWXKDd7b3ZpVffNxY3q+aDdtQR3lAuqHPNb9Fxuwtbl2v
QuEmgFElTGbii8MXCyzUr9pRYGTgAg70NTuo9bXCft3AkM6yjI6fttp/757MN4NyhEZFkZk1PXHM
8FoN5AewsN6yoLXDDxMQL4x8Pn3LTIkKYZYN87VZQ1JOsh7HNT1esJ20kaKgKMDenWG//7iHhiM9
7ZYjlgP/xQldU0Nr/aYo/Nu359IBd4r+kzleIwrYb8IeENTh3RavoHObB917F9s9hczelPzHUDTL
/vVw14ML5VHjTgaIYit9CW2DD5Ms7tF0RPMoSP23dbGV/dXoh6mIb0izuUpfV1RmbrW9q7PrFnrE
wHXPbiQsPeq1X4FnXKbaGHF0x3x7fXAv5UIpZqVmeU95NF5ZQ+mOA8JcRdIliZy3JNuRUS8S3ftr
Cwpfp3cNdiUgJtGCzAnkeDTNUMj1tCT2DVtYLnan6FHtWdGe30AeQJjjOVVpF6xDgqMcPF37pAnI
whp2Umc3nPTUgly4p8Zen6/DcpBaaC7ozXWUlSFWKN0XZJwVA/EmF+Y2luH8ZSNnNf3nnquGQPEh
8W6O7UAhqRXwTuzygk2tISgWZLTjRy2z4yhJ8jbvvOdB+MsIGVRt91ELvsnWQ/61TPSQMbZFC3za
4cYNU5fwalfkrQpw+xc78gIoJ6msvHzWZA2hIItPPfGfPv3BVgJbOENj4NfZ7xWkt53ivU8XTNtY
/kPvTtiq00QvTNLQ1CpQBeJOiQdH6svSKBfYrsVcbJiB57b8m8DAa2Fv5Co6xsoXAaVJKXL2BxSm
rt9sM99RcTUb7/We9jt4c1NAh75Fza0rtIz3EMyt8OoXOB9ha38Nm0Ga8ENpYAYWwob71G0RtZgp
+y7Q1ajImkKKiFfhTUECKxgUiMkc7jXTnm8DS0ZyFtVk6rsOYJ+vGyeevG65kCtWZ2F1m94j0WcN
qWTPUELetqkozZMGzhU64OGyRcpvrVJYtYTCwqTkYn2oqJiKMFhQU5AcGn9TplWDxHzWYRJLH1hx
Rs8QPx3Rm+mNSqOlV3Y6hgRqz7VGt36hAedzFyfxOtuxjl4eWYhxgpKrx6uh3RqEvoOkXQg5UElt
J27l+2J3FJjzFtlw0LyAJoDbXEWPojzV1/sgA3UjyYg6G+Dcgf6Xfo3CsLFIAbCYkOf+F3sjHGBA
GTnCe4YTggVIvnxgJZ88E+i8Wwn29bi0fVMDFxU+4diJS06Z3/j/uzLr0SotlRogmOE9hNSky4+b
g4w9APtsX7z1UWXiejJV0BJ7dbNm6VgzBVLFzDlcjf91eWTmZZ/Srn2nh2EnKTB/tPwqqqBZ24Se
tv5HM86T6AAt+zVIn7rHevJQEemQf+OxJ1cvY6Pq0V9jgvLyp39uRyfd/QD+KfcVH+Fye4f42ej5
3j82U7JcaR5KxdnvElzhbEXrxq63V+U8I03RgqJvyufnwkCejzCC878lTXY3fclwy7hcW+Jc9kPa
8SlxYK8t8McG74tW05Ht0Jim170Okd5c0k5trjJTG6quwEjbbzyNc5QeEhlVyoVZi1IfdkgdoAw4
5RwY8oG/ucH7LBz/rC8UptkRWzM02LpY7/AOvMkPVVI6qxmhKkMtU60Nqom/gZhtTdszJ+YWVo5c
KAvPjiUNMjm8NWzqxQu9BgxZLVfVewBElK+MZ2eE2UyyCD6EK4rYbOuSEQtVmFiNuWRlAwzuvDQX
9DoKMuyeIibIddTAbt0viB0Boz3J70jqW0eVTResXexEOOqlvfd9uVIJJcnThekX26xLwXRkwj8o
+OctntIRfP7ah/98pCOFneo79badCNgHpXUbI+eGiUNHiwWr19TStDaEsrP7IciR10nSI10z0+oz
b9nmq2wic/uN0TuZcCGdzJSkrOzjhhmd5hWGfnNeP3hWkoK7DwWbMCfwg9Y08h5O2FcG1wCd9Dub
eDn4n16l/0iz0Q8LHoawRfCTQof9mXZCJKXrh65GFxcHD5AXYCpjbBIxLF0Q+QC5OnHM2RND+v2L
chnfg/W6YrnkRz3nXddrIttbzVa1YLUtvzukwzxqKHeOvNlebLMg3nE0JV76V8KoCF3WnBlWkQz/
YJkP8uQsG6ICmaq0cd1hAEJxq9EYmZd9vQtveY14w947IQt/cbf3QcZWDJZsF9F/GTGuiCcI6p8Z
C9izla0QYIO5G7W0tB/tN7qUcMDsmgQaXnXiXJKaNkpTW2d+2J1eZNvIaAjGAdE9cZyRtyhYbGsj
zxqya1e9jseGnH+sEZWskruJgcTfO+uwR7z5KXEj2VMSoEVsfVG9cpdGG9b9wHEQ8HtSRBJyox11
MWGFsjEz4R0BCiPnoc1VCwoMKGL+s9yxAMIS9sU6nyy4Yqojv5jAM4wyDi4qcJo+ajwBrqqczpQJ
shKiR/nbrPadXCQ0O58plnTTAPNF6IkCroqP2CBy6K7OaBTq7eqSOoYd9yZKEzEin8wgwokv43dG
I+3MuFG//S3SCB8Fc03AqsmzZtcTQhjzIHMuN+s7NYWm/Y2xN4TZXKdypWDGclxY8hXCP/QfUd+7
s3Ulphdex5GBy25yrJR8QUOZ5+GuEo4xTuL3qZOm8mzJlLKPSafrvDwjnT1Vxwvnu+wfbXmxt0IH
n3WFv7xKW0AF5UlSZuYj/Kg8yG1k5HUkhUmySntlXurKElmr5o48kBQd9q8Z+a9wrZ75CrF1jg5j
lpXZjIvIXNXWJPAjYx5gV1Y4qSCfesuB0uw9BYT9SE5NRYBOyqIAAJ+YTJpQeg9/IEAuWI4vjjFh
jQDSJvQ0Fj8vpTYuuKb1tL7ZOaRuGHuSic1NDS23IjwSi0c1Df2MdjrBy7llPMzKIJ/h5oMelXGY
oJtwepi2bxoFXJ3u6MBvQypHgKUOPZfk257WOhLobBgho6e8awm7mVH0guvWt9/6YMBGlgZH2uOA
m3chapDAh9NMI99Ury9z0QSnA1h0Nkw8RTRvotmQzujUBNALC9XjWyi1rOEggxKSUdgcqDDPTE3X
KAJ2CF82wgdJxforpzBi7tH+yRU6vXiDpl9+gWszixkKY1g75Mus2x9wNeDRoOJ5Rr53yW4MhV6x
gRLCs5qw/tLrPjJ09YTexfmBUZkRPCfaL9VgebHmVtL0PzbGxUAm7Rya/9dph9zIt2d11loI64jc
06j+ZEI+pZgsSJLETBbyde0Flre+yPYfYpcKxKq1filGD08vOau6gofPWggdItu2WX0JbLT25Syx
LeFHdhFnaXM4ghp8ycym7xpt+dIC0kigN9mBMSU1hjn2t46tYI4Evcs7eTg/5rP9ETFONPYGcoiA
TlTn5LR+eRsyPgDlp37At2zIHPjONwhMALqnjgUgH7ZlMU8Y5efF2kZG+IvspevxqHDX5OMaG2sR
QEtaE0YAR4Teao18gDv72unQQ4xHVgRucW4zL+NSRIHcCaK5ZW4QsGbDZCOfm5G9coeRexjY//E8
i/ihClT3yZENBVZnR7F05tifFdI4w2IHu6Aevul+g9XDQVrgH+uWYpT8t/A3EA1ZFw/nHh4/uf5d
6zSQ6rNLRQ/EKINxxtGICLOeENrUILpWUMr9CFc22W3olOZPcDQ9iFafr/9tdB0eKfv7pS7+x0uF
iUl9WHsOw0vSlwPfVqs9NvTHKdIWbH0HCL5xOrBTWcHVL+MVZa//Tg1GVYN9+wlvMupO+qg/cBNr
WNKeacoAMELmcej5eM6256c46NPUR4JPFxdaAHMedjaBSiwVXXZJn2BnfjaHnnlBKTWc4Ke4MbK2
6Z345+vxBd8rF6/3YM72+ID2gPj+wd+qoM8BWFNp66z32W19Dicy6ovDqgfKpa0plgz7Zi/uZU+m
hrR83JU+PcVo1zeJBXSA1dYNS8ojEGHxnBmI4e0Z9QTRm7kK+1v7hWkClQT1kq4Axk7IuJnDaSox
ymRYP1HJ/l/I+wYePpVNqttDrI2aQ9EAceaxGZzK0kgjozLpi/prwvRiaIEaxeIWzH5uzC4GCSMY
mlDC4owNmhQrrTjTLHOjcpc62QMxFHsHU5tO4X0mWDIpM+biUTa64sx9V72wFaIAsXVwBtiieUJM
bHv7m2JgImCd1jXe05geahqFnHT4yWIgoIXWqS47OHv7RSTGQJAwA6slh0eIR3FSKG/baAmRwebC
cbsAu0pO41CKisKlLC6J2yDAG2mM/26Kr8l0LNGh3TYz3yHek5UppgDVcRdxlmbeM3L5EiJa0DXW
LYrIo1/9b+PHlz8T++vM+zLnCWpd3PDItUvrKMl0r0Bvld01tyvuwxot5HffFuUAIMjWnNiUyo4s
ik9SLOgwevD1JnqVaOsG93xh7wZJ+Rc44R/L2s9TMgHjKAG+Atlunuoc0LopKAULXOYVfOtpGd/6
GHlyhGI2fg+W6kR1e0qPAVW1wA61EJXGt6vFb46H+bKspF6XSzH7mndvUPFel+4zpjRDv8GSPkgy
dWVtFUG5oMJx8k5TA47E4GsXJQJlk8ZLCza+3jTiRM8xz7qSUEODC74jtfZoHgwcchN5TFmX0wOL
+SdmuJ5n1u4c6//pcpYAi9i/aFmC3wEb0lnXbGvf3SBMH/OeU8/eejt6a+/q88yFGMoPAmlVrk9M
Ik1WdCo+jwo2LZtrpjKbJBmNKn9jMIj3gHUlH5TdITTe4Um7teElSDKXp0iB6PWgp5vTIUMMSL2U
vNB5jr1wILUBRY/gdO5BveDZmpMbM1Ct3i3BRKdtYk0jJKNewfNfCovTPIUNrQ9mnxLCQEQ1azUL
XSkSIRsaEGaVeQUWxoQg9lvDGuOYS2hM/fpFQZ/hJFoLp/79iy6vQGS5FSn0dK3tiHFm5LhQ/GTE
95Rg1NADTOsl+Kk2sdKUvT+l/HrdQHNL+E5ZMsa831qcjU75WQ9ALIUwREm9CikYC8VFikCI4dDh
EaSRE7Gf1U/6ad6v6VIJNpBu2A+TOJSZe3nzW8bdh5GI+rEEe1WC8YBZuz3oftgyEOnSrhF2cLrh
c7BX8zx6jttWvKCAVMcQg1XuOX022zPQbU6arb8UTMIxyhlafX86PAnQ9oOcaUuU9i1mZIRhnQGU
tp2cOq7NvkJiWN+LsuLZo4qBBHZekHX4C2ofAOSl05/Q/uNeZWrT9zg5VJg2w8/izAVd0vxGGkzC
n1/AROzbw2dymRPYUNS6J3iuASdc+8p2eZTcKvVW0tH9AdLK1FwKsdUlL8Dq0wsZoPVFE7umeAmJ
68WTUg18BFLa8wuEGsqKZ9cCN1jEwCB3S0yGtuZOknTMcHvQkVKMOakiHC3sb7BuysSnCQtPAani
YXH8/J5Y+QNmeb72imUUb4w+ASgyOJbTLzfXPJC6OheIIWCsT7Abxw7yxYeiO+sVbdCHQDcpOGhk
d+07Y+JCpkQYtzOwnC3Gh/G+xE3j9Zxm7F6HYQ8QlT7vnOGzruw3PZmrx9euLXGVTJx5U/lMqqRo
+cwczQP1wk+h62IrZC6zMEB4LV7TiChm6EzU72799ohhG9Lh2Jd+AoqAEsX/luGdG1akIQAVUS92
QnNsbKORYsJbK+IfoawWsoyk42CdfFe9nWYNcgfOsLd/s86rjodvRzMOP7z8X3OSve0fRc1fFBl2
prVzK89SjFhGkVNrsijBQIHtBWetqU7t/CJAjBvZRRpOiH1vIxS2RjtLOMpqg8p1Bgt+GOFOnhce
pYcxuqKVqoKJeuoYVnegyLeP31Bg7IfyFcjgDH2il6sAlZ6dwJi1lWe4ROq3IeVCQvjuQoF0sNvA
niYlwYDuvkXcnavihNJU2nOF0kRpXZot0RgrH3a4eOMSbP4ouu4bk54F+KaRSBMNNYVi1Vf+r8bE
DxNXe8I1YO0/wuxsF4Cll44uWnWYD8TAJ8K2LZo0jvt6rANDrKLbaJOwKT9FABLkksdwnhztirVd
BfuciU6alQlIFlEcv8rUPbGWYIQF7AbIBoJpS6POGEi8qbGK8hITAyCAw7usy+eG6d5HEZ1+fNFN
3Uy3PkNzJxjRGIOCpSLkyMF7wCEiF5aJf9vNUfObQpw7XwYcIg4BFbpcVjvAfpzso+C+D9SvpSKF
0o66W/QeORJguXFADI0mcaomRvYZ4zefjPlXihhwH3W65711dDn8IwetGWPL6WScQDuFhiyRSHvi
8+Y8LGnr3SMmk/NBWkREGqyQSVjgWH/t7uOXFU+Iqsu5htEa9uxCopIMc1ES5aEUIXMBFlXSslyH
dNmQ/RqR//P3JEfLFx8oynMJ22hg5SDp8nU/Xch95HSRWB0JQTPN90AcCdQJ1R/+JZKo1RTIQPzs
UU2S/LFzyoBkRSXcrAahF3/buijcRDuhKRqxo3BfcHbFh5BJG59SVHNXsXZtWgsKxABbsNgWfij5
DZ6ljDkV7dcYTlEZK7lxVFIxEAHkf+IEKDcfm5c7nAn92B3kCmU7HFdgpmOewvXt/4YrAqn6ETHN
iB/2a18W4BRxGbin1Uk1w+mikMRE2kh71RK6TmzmsSHEgziAI6aifXB7KHuegddWLqGvCYn+N6DK
PcUBVOUZSktmPyt+34B7H+cxtMGgvmQ1y4bBG7mhRFg7BBxkT2JTSmdk8IKYk7DeGvdVGoJZ51EK
GVOd3DOKhCxbzJUXsSph2LLkGmC1KE+F0SpTSLFm3NDhJniPU/YhhKF4LUp1EmamQiiRLwoL4uVA
Vaf3fYleMiwfacy1WnjGcUbf4Tt5fP7aOcipSz1FjIbV5m/0oWjtX60Msk5HhjXJkhUjgcolG1Us
6DBRDtcoTkeu7Jfakceu4urShZrqL3ZKCCV/m0GMJaOg/Srlc8ENl4ohqx1cchYC46Ds7hN/rKDo
A7uKuySw+z9PiKfgxKVGaYocwraNDRuMLyte58E00yOJfGmU6GvMlzbN1QvdBzBHK/Lf3t8KDRys
zfB/i7H/rGiUs73aspvtONFinmdqE+VU+oXXyDQkX+K8mxqCT3FId0Jt5ruGjDljnr80m+U7Cb5i
tLBHZYowY7cGvd49Md72mkz+dTz4c3EVTfGtfBORZNLK+xS371kBSKKB3cs6x29lazsJCzHObZgd
TNVlZdWQmNwkGm++1pPgpcvkHRSh0PAnD+YSBIGVBDtwS4UVAxX/rhY+FV+FNa47lIIG77cp42Fw
pRGHIBy0iuaYvothyKVycrah2L20k0K23F5W5WpTW4C3RsAUZ0om50A0paBX4pOK2XypgF4YyTAq
pofBWKZ7eEJm5elrVb+QYWw7pkzwP11JfmeRpagSyLiYao5sYE2TtV1PVjkptYeE9Mlitwnlyg2L
U0I2LV/F0BioMgOw3QWeojm8yiV/kNVqYnsSFHvK0J2YfeAxXfjhjLFWCnVcqjmBF3z4JgUdHb3e
XP+d8JM13RY4YW+ZNKqYNrygOSoHRFGydgI0WJK2x/M+VUZmBaZPpbBUfpRZKInmAdKS+7nUrqW1
ccmjtHF9udcUB7RRJoZhU/8p+MuoCeabXglkqIvR9Fe1T8knX9lLIss8aOoksKIfRI3rct0JMRPS
kizbGdKXBusyinUFgSugrvLsVZNCHR2tw+3aXkPB0N2WND8ZdxuQ18X0ARzBMLurtVdDhKSNJCeT
zc5atw8CDlMgtebHIu7DhNJgxpIvsn/NwmgR7AvKa+UQ59t9XovOFmeZgjZDQuNQRMm4mGENq6US
q9eQUlmOv2q1VFFN0Hl6daVBMaAEgISE9Jthn7OwcGIQ2FMUgr6dwSUX3Bh3Gb/0fEQ8Gb5sjU83
63O2zBI3cwSfqDtbvaguPPfuw5IOj1QMdrVoa9EvN440Ax9p+YK4T78QUWhcPvRphomjg2HSsiNX
GTYKpgvL0p654fLbw6ncfqAlbmerRFdIU8hPJuTmFbSB0hGgLRaNC86uGVavDaQOGkOUmbfegGHn
0/5n3xiLhP1VU57N6G93mJoMNcEfof3MViyM+wuFEFYqPwjEw/KXH6ydcTt/whgwYXkYMjR3h1cS
0GsvG2lq1osFLYTosg5ysEc7AG1jYYCCzZY7HZrm6wA1+eI1lBoGpmOkyhcaDz6gdjUieXBferd4
/k/+FQGu+vzcyY2cmFN2CJglU5aa5ksS4WM8fdg/PUw8vk4QvhJY/tnSQV5GP9OLIb51Z4rYiHfM
jWFxZk8HLWN5zDPGwJye8XxTlxSa6TgTjSSTs6JKnsjq5/SFid3VahvjBoqqJ/8filPhOGSfV/Yf
jkY670xsAXAnmOEA3u+0pi15BpSp/ueOovlqp7Mfs64yLeDoQybh5hCPmlZqnIpjLH7kJzm/Qx8h
pTctzYdN9obLO1HwwslesHSOA4L62ZsitpVZidj8Hu3yMz+btjnalqCaqu0dOhHwQi6BvTnNHJQu
CCdVkxOzTE60k2CmDFAHhPpStjoFqpsTv54X8XknviICrhS5XF6l/L6TqttjXAMt2IUpssVXDbcD
grlAJ96U+i9I3tkPb8eEYLwOyaItdJXvJkHT61sHX+96LZD+j2+ri+gq6dCOJdlV3YroMkTmtyf7
gBErNvaXvnf3Hg9f5bb/668MwuK9ONH30B9OOlSAFaE8a+53aOrBuBiNfFzcJ8YBehkUU3B2VmbF
BeZAiOw5RqTMwCPWPs70MB0zIupMAwKHjbDPCtaHJe6usJfvgX/SHYrOC7Fs1KLNRM0GhzeBka2R
+LTzLAe3V28gYqZlq6mQ+hIsbLXpsdKDwjqAaXSMfmRSBSs3SFPfkws51dsk57s31LSizLzUrbhE
dJsOy1ToItd8LHrV3b2WM5fmZjlR1wkeKKrUjOtD3HySK8kq95ayqqSRyguOUDS+BjBDA/CMrYzi
9eno1mgJCqr7wN5iDlxlwjSdg8RxupO83peqe89zOKjR/9R2uhQ0fCoI8jGgtK2addlSELhS24jv
atpi1Yfgs2u2MjNdQTRDTU3SSWCa0w0/x2/485jSWjmdPfKNRNy3mXJwWYByH0pQQk7LMXihP+I4
lKaHY+Xsc5ahM5S4v+TfQ7vBf2k09vN9oWVwuzUPCSQ03r2wIThfJNIQMoii1kgntLBXdY2dz6XN
WkPj2w09H0dySnO2H7CNPr0jzRKVhqOiviBdh7Xmuby6yYr1xzNGRlwr/nN/h8mwpnmYPeozfvxG
i+y18VSptoU0I9vCcgfAU5Vh1YVco9rhWRsp5MpsAgoDP97eaC+oP+i4crHezi53scN4Ivu2nVKL
KAfuzYozj4qvsdwRrV/0dT2gK9vjHN0rf4/MW4Ln2m1AFOMjhbI5ZJVUw0ACuipEZXWpyj/jqSLW
NeZ3ZqSqi/KUI2ccirCuZvKmqRf4cCaLj4bRLBl1ylUEQ++uwSsqgcodFS6Q6czhumdBYVEG8Y3f
PTVW02E5y/VaQWHeeKx5eodOolM9Mj205q5Ytb5YX2Vttf7VPkMSSxfN+9Fk5Iy2Krk0oWU+xJ7f
ksaxH6AznnGn5yQl5SVJpLkyI8OykZtPyuO/zsIePyfiL8GhG8zjWWZMAXkmkM0AVrCnMAcFfnV9
Si+DIHto9eJd1/ekDvRYQeM7g7GP0mprVqaGF2J6R21k6sEjnhrTvyLCU1TlYvoz/2W8Lg2kcAbk
Gtk4TaGrKAr/nt5B/Hdn7jXpDmkPJoNDCwm3S2qAdsmWWJ1v2IoK43R6o51mViTVg0Jk19KyOVFw
IAz3CBueQShrBsGJui4WzKk34t6P/QiXzpO+AQY+2Zu3tcVpE+rj08Xxg6LcyHrC5TSxzeNHjh3t
iF32YMDLEwytQaIobjFI19xIS5OVKw9pWTGoqXvbC6oZ3/+WBSMzUT9sq/t6Ne1DefOLdH2T+hEl
OsSXTnG2c4Nee3b4B1CKpr9wi1m3syJwnyvp8EEJIScPI+xPCK3GQ27Q0nsO7CrvfZ7PwPvwwfEL
/7VWk0+IO9LZoWp9QdrEj670ZNuRrUabKDYGeXCytI/wQjnFRB29UDvnAX4BizOQK5N3KcRZkg40
5NGGgkwWsg8qHoDcRWWly6a4u7c+xW+c7rDDGnFN/wuiUsP4PwyaOJcvTdzczmsswwYPsZG1IKKx
z8wxMkDo8pGBGGtyJSqG+neRbJGZss4SyhRT/cn5j6lsOobwfJxrdogb9pd5cUm+Vpi424VsE/4q
0wOx9c3671I0UUMWesSm43sXZLHeIveHYfraB44eJcQaD2wSBgHxbCg4GV1QdXK1gvJAfcr0Rky1
LXOb++XwLXsr/h+XLzs6Px3QWpTT8bsw2WlAxAm6E9VJEr57TpuhjRqrqMc6t2T4PClzzfuXP9pm
IGtqRKEpGITsTEEy+SjlNUBaRkQJOT5p6kb9QMgmKkHqy2hS5KqFDHRcmi5EThRZNUjtLEFRnv80
XpRrzCe4EFyuPm4ncotjWFbyw8LdBB30uawlKC94+xURCSTnG7q0XUirZItFrDX6AQWYgY07AZmz
yuNMgpxex0PEbOwwjeD0OxBuTYn+9n3krCy0s6xvA21TY5HWOYDUkTzq1r1WIO6St1IJppY1ya+A
Mdwn4Ypq0Mo1AdlKW3hzG73iMLa99nwDLpkbCm32AxH5NYlzWs8SFL5wVQadkYFZ7IGwLaz1Svdm
tLPw0j/vqxmbHCuWRdZ+iqmfCGlrIS568DneLkWeMQaA8OWUVYULS/Vr0zW5ufCGfmsFCLfnuaTf
XMQ1CEm79hdoncw8YqianwPI/movYsNPqlfR7l1c7YHO/DGQ/FHTB7fo9vKmNde0Fa4yHa0olG7B
15kflOE/cRAhAdKq3s8kV2MahaaJlO7C7lR4GIXWL6UuPyeYi/Jm1NWrKi3XF4tg0zqKFqoEasKi
7uNJPUoMe5NBncwvh8vauok6JfDnigvrEjiK4Xw+bw77gYu9nY8UJemjpNjDUPvCeUvgewcqHA0S
afNX7+6oKKoa0WA2jU7bjvyjn1VriKLOe0gCv3WYKWlVUdkv88tIYmVSS18lCjUXeg9ktHavcSh4
WuwJklhyXhQYjudRIm3CpXVC9el0sUCeqRchq7Jm5uqQhK6iSlp2uLRXTngNvo+Rk3pw4AYA7vKt
/n7Kpac4/7p9x0GDDrwvXj3B+D89MLTBfcGvc4S7GAzHTmK7n0C5G2KheM7tJl94tM7JA+oAiwKI
jOSvd/poQIzxT8UV+zsVvZfIgVZfXJlD8u3zee4q8iVpamZSEZNZTM+BozEe7EqsIxJjhCltI8OP
8UF/FedRJmWjvnb+VqHZapJNz/ttKfsWmzG5JB1+K6GGF9ITN0AU/QI+X3cEOJt72i4J1i6bh5gR
pukdsZorsQSmCLQ7mYvwPzjJaLF0vlHJmWwFMlvM+B1c1KLwgqPwF6QjF6cMc5Wjgbgycz7VrJsS
HSFb/EHsNMuswUG2nXby8Xx3QTwSFQBFzaukwv2Hw4tmRQUSA174k5qZ/clfnbZG41tlFrOq49ZW
bBj603437KDds/whe0pSInc0T4L3P0IlUP7GejntN9JD/kpNOkJiHObJ7WAl5kA85zWeT3Wo5FVk
6pV72PHit9W1ff72pWgU9sXs1MTz5JhRUFsco44UoZRoj5I+knQVda2PE1iww1qclTl6aANS9w4d
nFDJzUEyrIl2DQAF3fXfUQYGuSQEBj6wR43xQMMBv+lnN7t3S5NJg/h/Y/ACqUr57d4HOISxjVHs
Qo10q7jxe/H8SFbhwH7TiOKu0pIlnXsbIwn296aUrrIoo7w9QmqAsONF5Gvm5/VdylEamS7VKPNn
PM5ItEE3OPnTn4vUv9xXz8FWfkyDnh+q6thwQK9OzG3kQz9qHF67+T3tBk5+V/K3bj06LEZP0sT8
naOCScXpokrIN6J9/fIojiSeJSIeLuvvcaJgSOfgXNvq/FibyB1LUVuVM9rchQpiQEH4WvJS1ACU
Ov5Jtvc+XfDvjlHreFfahEvFEFEapy6nV/2oPHVBlqqr+Yyu5r7gSj2gWd8rtrGNws5AowUsgVzg
uvb52DhUjUs3l90ODCITn3RBcoogwkAnsnZAKCcSTa1UNHWwvw6aw14vkKVSS7JNfgkQSzOwS3K4
G1h0tqRdSdj1obBzeuOb8JTueDdGchxIIZrx9dTEFBWqwaW37l764N6p6eU0ym5f+f4T+lnCNMV8
ytHyGoQjrY64uQJvBlQTVV13hZHRTtEEoHE3v9fflpEDzDQQQgPTiXE59H1+gRBqtTK6Zu7onXC7
9WacNMZJ8KrULEvMXDKHatbo41cvEwktuNV/LzdgfDw7ABafPawYncpO9l+IK7jaWdERuwHwGpA9
t0iudYR4Q5e42MrQM57YoLT7QfCuiGFWOTh7QAtVs9H4ihU9wF8OGgOXcI1//Y3dx5dlmZ/R67xn
UKBsAuR9g4TU895eEsCQZgnRrOhNoLsDcMWNE2B6VL7+xhOdK+S5DtnYyVLBiXpY9gfKydu+AQoQ
JvvcpOzu4Qm+28Pdh9ap2iCB4rCGF0mR3QsOJf1nbC1F3IvNg5haGbz5hzJ7ijHDYz1L+8Kj/3lH
u7rhN+39cV7QD/YJzB3t49MeBSZzqmBBQbPKGm0yaZqS5due3NPfob2akzWVBfhXBj3hR11RntG6
H3wUc/l4TZCGsFX4UTVdjsK7oZi9EzlBCeKiVBFtn0gLRfATp9m/p3VNqih80e4fLUL0VsNu1EVF
iNiJkSfSAqUNI5G1mFa3KgIPdNJggvIOG2p4dZF0kd15+sz9ISlf/jvPoRhZLbioWOqvuUn9RmgC
ZFFcuUdBnjriDBLCOSkKADtJRuQkFGgloxPpulI+8KPvsa/sfqtImxIBdoYje+RcxeYaWlQjJry+
s2sanOkJhPqHlFqT+lDsKDPbYyGk6hF9IqaON6XmFzrLHcjNNExeVMvL+irNWawom6IJ1C+LPK1C
R77iCz1Lr6ruV2O/daiWdqS/epLxo9oybmfSIQTURpDbYTfoXYQsBz9iYV13g9Jj5meMVISRAeDq
ADXAlKizj6vG9olNzGDWIPvCA6tZvXjyu1JSPoG7xI/7xE1CybAOiw+QDyIp41xJajLelUslSAKw
JRlCPZ0f38ATtgGLwdNVfToGQ/h8ygjVJPKEwcifg61cSpaMdE2wzwZeh+IeOYDIP/Z95qVAUSdL
xtSHqz6OqYgmWEe1ww3o2X4UhufSJ64a5ojhqrd9rLadRSKj6dLC68/2FqdmXYqGo6LsDohx9IUl
TbD4ytcr7fge0ceF972UROFUgj/jhg3qnvRtWzUERliawa2G/pALrMgYu+g1kOKOJh+Q3JqIAhav
TvwzY1SDH7+z5qxbI4FnwG+9gL/lZy/r2AEUS7L6E6BlUzfRKp8KjmyzBpe8WwLPcN44u4OA7u4N
j//LATIbXSdCPKUqE376wFXBopu/ugYRn0B+RJT6Dx8cPc94NN4t8qkt7UV0Z2J0q0sFIWuJ0UA/
2dtvRUGQyrvkFQiDUx7d9ULXYUIbB+QKQIV6wcRqpofNlRqOFBu8g6jQMWTbSpxFLLWFDFdu0ItE
Y36jlFvTv9M7tl+3iDs6k+z5KW8iHSmFOPd0X2JFbFW5rXrmmJC4pqUGJnyKCxconaQOyo44jGRy
IpRMBgxpDo30l/i0sTUZIr81lIV921mcVfHzf/hdCFESc/+F2tXSgGErz6J63qWOameBgIWn1cgH
i/npgJpxhHXSY8/u4qGmikQUC/3YLutYqgEAMpWMWkSaVnAx8xSg4y1wlJ/SF1PEd3bfMiJcZFI/
zWfrI5uVvNcWpDC8/t6JvmZBj7Nz0lCIqOvvSM8grfW+oDJ3wf+lNTCoWPbCUXDP30O8PGD6kigU
4WwdOPI5MbeRSo70t2QJKgMKWvGmq9Dfmsjh6AxZlzdbsRCipdsaZRQFeMMYQ/KxrYycSujgpapo
hzAwcdUJbauNXFCw3SnVOjWxVrnZS/mWVHyioz3FL9vMM4IxVZMpz7FWDnjS6NDCMC6rww/4/D1I
l9lGVTX6Uc+Jg0xaacFRZgjEFq0IFpAmoA02Puig7cvuIIv/VRq3lMLDNV+0OtxogdLcELihxzMt
0S0/nfQK+M3LK8nvBZ5BprLp4lQBEJgVvY7uAVsbypdUgY8V8mtYIKups+bnE2v2KxOBDM4nJcZ8
T+xp/DGk7E4RCo11Akos1HqgUwV9IADgTb/f2isqer9C/2uQjkIQa6/zMlGVAGhuYlKITQ1f5FIb
C55jShVu1H9BebnV+iGr4QI3eWvMhQzn3FgnHAUESn+F6ogWs3sI71bp5+2NjvqF5aoSTDddf8MN
g1hoSxfrrwG+4AcTX8+LE1zwBCjAXbZviHcUraSsMi7M6MJGlrRuzbBnX2QzFy29n8lUODyB3/H/
58l6vMe3qbZOOCmmKeqPREFvrNeAkn0+KdNGJB8LQlq+dfOFh8Qcb2Viz+WGtC7nRTZDoKEKbWS2
pxt+7DNrWhs5eQjfQK33Qfzmaoa6gDvLqc/xv2FaOQb+9tA/3GLcwv/sYZvyfo9vqbUHCW9wv15c
pR0TJy8aoOx3WxyZIZ7/7rIzEtQr2lXVN/51BBdP5x32pBLP6L1i43oTFTmZ5DkId5s6GJcRPFPy
ENLCiHWXB6dgoAiCXAiXy46PDQDk18i5aBYfzeo47uzJpfEsLizhtCGW30Qx77kTUuvqkhFDPy11
Zk+knt7/O8ruA+q0nFVb8WHuovNAKYfIjiRrN4q6l4qfGGn1sahO4RtZw87OZVSK9Q01MSMIkZin
j4y29flM+JrXRp6dnYOtbueGVJelzIiqLRV5HWyKmr/KDCAjaTC/NGqGLtw8xTouELmj+1p5a2Y+
Sxo7YqkK6t1vh26QC/oZr0xG0GG2PWULvakgatU8d0qxTCV3P50ewy+3yciOnV6nbTKcD233u6H8
qpze2x+V1a5TyE7GkHgT8aLsuaWDBUYHBkm6TcRMPejC5FXjCt+pYX/OtW2PKbYz0quGs8w8aBr8
yHvX1NGW838D3cFRCya3EIoHymXTbLdH0RewUfRCNbMM0l3NcNyaBH+4bqFm8Asz7SNeIKC01off
Tzec479EZUuRfdgCSC3IcpqCAbMcpyUMuRES4a64bNr8rj/lQdmc8ycQSngGPQ0HNgyvNyj6681o
rQ+UPzqfQy2P/TLKRDWF/iluJmNk5OFx6z3LJQ/QP2zJm0YbL79Z2eMl7uUT1fyPD9ewq/wUWfrm
wt12wMLihBBZ8z8knPHEjOFUymimh/8NZJYsFAfKkZJu4KA4XxxrcvJuefrXyUsccxBF1MIl4sdV
ehgEFdb5HUPq5hvNCv1Z4kShd0jdhMdNbcfrLBpjaWn9ljQFfL0ZaensVve0V5ydNcZgk2IF47cH
6foHBFRPfcuPupfb9SDUAsW/RccQTuNUcEc5Xw/Mnscd490YH9bL1HBtDPiahrBy2tj/rp1s5CvJ
A2As9ZMqiqi77h2sB7dh9sLVem82O5zfqBtNG9GbdiC0kIfBEGbL3musN14eVNQ7rFB39e8KoPTu
xH+ftT9hKyuYGVANCbtyMYJrGIQFJ40XLblP26VEeTnhGHp2mr5esWBqVJ9XxzMy2w1d9UZhdkEp
78x5d8YDfQv8OOIbdLGc9HT4wcvAfs2c+e2Oz0DkPPZYxtad+6ly7fjKH0k27b0iHvbWtvnEH2bw
Pk5KMFWki5toKKJnBgnoTgxv+W940IFr+g+23f/prCvoYZAcq/6d2dgj95KWgZGlBp4abeV7Y274
BonuWPw/UMXkBP9HfQF9ZPv5iRR8S870pEZiv0Gv68x6KMM39uvkZuBpJ9p61OrwCc0DCgX7rC7h
JsHqi6yZS71HcaHb9lsm4mpXtqaqdpRHvJ6VVr467AJXooKcXv/kx1jskM2GwfH33ASbzlIP5AtY
ombvC6BLJlRhHzlFmFWBFbQqSoTTH7IZKgq0SucFN5E21tuf5VLqr/PmTCAit+p3Vvhmc+/9dQpD
9pEjY38ffCj2Jl8Kbkgx9G2BV/XS6g2a7Bi5o4AhI3f/dOVHv3P5h7HdpN7dfs1QyaXLf481biYi
p+h75x+Ei9mtr9ZFeMAYDnRT2uHlfdob0TpVb/w6s/PVi4PYwO3vyCiM/ERJEBglt+/LvyS7Dxpt
g2w/iEfcKdPftHxajP8EftBTD3QZW7oFLr3ODd1GYohPPaetOHTkuHzDW0KxrOthk+koYNfRk524
6KJydTw7aOqExBqnfUMXn6rEM+DofjC1t2EIKUhNIJHmeFUC68rI8EqT+TwZiMrHPn//qBdkAlzU
bUAW5Wi259CVhc6rQy2rMI/Dt5J178vTR3dUzF5GEisVskZ+FKXjs7NIXVn3W5uDD+O0H3S7ygVR
JRWmlAGEL/ltonB9iepAWx5kQJrHJvfMOd3A7VPURTmrAmLF/VEABmrck0SqBkb8zabEv716sld6
z290pePaN8Yq0pe7k4N5SI+jqyYi8OGfqDc5NAUBI/ao0tvklTN5aqAXJl/68J7RYKWqJ6FuV5IB
v4D4wx9tlUTwdNUU0i+inZrRQOZf5LQCc/fWKA6H2c3Hm2ZE5qM4dbNFQhW+QfbI4ImhMr3/zwX6
KLe0wnpGZGOvY8n5mG6bP0Kk7c6E4RisOQkXer63BPdsSRVXB/AtDk1p4MqBBJJaS0agQQ20a+xE
p/jQx8/eKoMVnMRZlzxkqtKKHjsjZMcwSaiZUcqGA3ZKwa6ee+7jDTdE1Hnmt4DOAGDAOAulnsuI
40Y4M63BSZRZuPREqoDLHGIRRb6/TzVtfM2i4336QBBJ/V6q0/2De8MEKBy/q0BZqRfCp+BPhTWH
K9jiDLH8mkd0wv7CHrd39E3dtUCPWTMrcUZmmVL1g6VuxKM28se+kIwwlejeAEB6N+fIcK6ffizN
1qRuCuIWVZaQWZHEXsUaNSV6GHj+y6NGXKPuEIiwXHUjhmcL1gLsqPlpTpJx20m5tksfipvVIVJu
rlP8lt3dC4GdsQSLpJzQ2c9UXPGVeH5VfbLzDykQVeKkv88QKZ7Ma/gcV2Ef9Fynmizl+lSFMkRB
NsEyEWOjaYpSWVY1swtBq+vtFGrdgo4w+bBYbujcRHqen3fWVKOXypXvZrEaQWhVpyNIB5aptDhU
VrAjjpHAIvBDtsIE9fgdLDcKgm+cMEREnKcwcMDcdHKq6Zt9sDiluZ6ZtvlX8louI7LFkfsx8G/A
iSXeBWtkjNft+or4Q0sVQwX5hdrResh7gqC3ffeUcRWPzzULxfqx2ga+RYi/c61Mq9CvE7PMzTSn
ubRkYSfktb8N+vkHLt4mOXqKHeZzOSysx6v4CyUrk/QeD24tNGsEHnMrvDjPsw/VaBB53K13SLUh
PNDfmvclCkhtWthzLMzlzoFplrqY+mn690KoPn/PiuD4/sFycDYOTOZxt8Xx6hKVPJZzFbgH7Tyz
lzj4fbZBkmuAzURgZI/RAq6p/zVbK//Kh6/xJqIrEJw2HllZ+32WW8HfNhcYg3cVs3EKNl5wpneO
ghu8sEH/I0wa5Und9khIi/Qfrw9HHrIPPQC7qrnlsGSgNWYuu2++uu+RMIU//ojH4bl8eo9URupw
DQx2JZ8JqafK/Gj6vMlVR04Ii3fR5EyChe9WibEP5Thu2q1bX+BOe13bO9/k+OjOHyV/bVCu6kIs
WR1q//Ao6omGDbNWjNB2b4jHAvsKMXUyQI0uyH20E8xYoOiUMU6alJCbxOmJpKY74/uUNYoc+hpb
kh7j2o15WIfhl62yEANnIxYehJKdN6m2zkZcM81oEqQiEY/MsEIWrY8jWOEUZDb71PibT5JIJ3/g
krgLs+GW03x5gIgnzVX2UcoRPuSe7xZzaGJEfZ/+Ho936rnr8WCMwq8Xf9bTm7cOQfgLFXopvIQK
Msnkbu6MUtryI5CNV5AyKTDHcgxKlIrp2mdSpialu14HipB4tj7IfQiHm5ECxDjV40YNlK2ly/kw
FyTxZOzDL3HYilspnahfCSC19Pp0MrienJ8D/SF8mG2zztBuqoPfpsoMX9+Xzo3GLGXjOvzuJSUA
HZOHzyXOE1kNDhxzjXfavNsfLX/CGK/G33YBrXqykRg8gGNivRcoX3b9IkSoMO1ANarJuGmGF4CP
syOC3JS8koHryI02n8hmcBEPtZV8rWAkwXHxUf5NPertxX3T1PkZGxwK5IorbQoosWmhX3q+NTlE
37Wur0+v8GflJqxIVKvUT6pIRS9I23Q2qLRQRo4W253r1YDCSlPgIkwKHiQAoH4SzvAVN4L+ig/C
5UPJ3xkI6EiLp11A1fD6R/eqJ53t8piLIzXizD4G5O2I7EBk95TJfugb/As1qd/6OUP496JsGTAB
SoMRQzOp9n2Rrm3HEY4TQEskcZW57NZrTF6UPzNdu998iny1r0ENw6MUsp7HBroD57Y9vL/0qLsf
tyisNuiFIEI+vFe58RB8e1FaFi/KraZiBqoecPJAW1qY5cMUslVQEgzY/yzaV0HWYTnUliWW/KZb
BTpJ/gDpXUyLSnQf0cVy4n8o80hEHpzxjTU1ci2pooPp8mW/TPeoGq9wspYymuLlrpcoVfYredtJ
z1gXWKc03Dg5zFlM8xgW3umAivuVK/oAvLRKkVzcGgUbvjUx5CnYAnk1xxoMXgq6MS9FdpelX9MF
A3JwtBy/q576u7QRGkstEonfTRC85OiCwXg03yvfS03NxXOq26aG0MSfW4qOChOCWDvJFGh7jPcN
CPwDeXKE7NRaAqQxcMrBz7Fi2FetgyU49ra2l0JGJ50khWAM9rT6oTCG08Aq9NEyxImXcZJaaKra
A05kywymq1wpULWBfHXUlX7TIDEYrCfBsPibDn7Fzm889jfjASnPcD9+CoWMFItFBB3RYLOKmSFD
puSNp8UQ+LtomdnPnitRk7fTgytbCqMfInfs71j+4u878VpTRQO5nAdDcJ6FSW1LyTSS5Rs+HfhG
j0bIV6zrHzfWy/7AnHWkL/vpx+GoMTSeDv4Fgc/bqZF0gODkl4ubKjZK10BA5bwixZ19xutecOhJ
VdWpLG8MN19uqGxiY3aPJRD4O/zZ8hax69oryrDGfhCM/NB2A25qRF3YmzZgQu8pg3EFiqEh4DW4
ZrX47xT21jX3dR/3lZivhYZKgJgIz2NAn+g0qc6DczRvRzssQ5dRlGzJYpU7cdmWT/31FUgm87TB
r4E68dYfJ4aCzEYNwCAYM8/1QJRzEDdHxCEXY/WfGtDYT1Uof/tHIJs15Ci49fcIk/hcs/Y0En8p
KL5e7DXxFqu2hkMp9RmccM677SWYTF8q6JytoFCY13U8VxY/w2XMhiPHdUtI7/fmlk6GF3/m9LbY
8kW7xJIv/qxxTxkKQ3j6UPPXs5IqCiY22Dfijfq+SDunHlbNFYA3DXM2D1uyHsoZa4rBUaqLmDH3
1ptqeBfoSTSEC1F39r21dNUjoMK7cCQuIkZgEUAp27qXDHPwkwlAB+pqQnPpt8UfCGZNajCv5CEX
fw1Duto2xzwZ1mQCeKIevLYcfZQdQIN4mphskiAh7qHRMCszdQuVzGEAkc47VwakCi3qCi6Lk3jH
BlqL/4JFBeDrCD9EGxJhh1+Dl8tvBnI2enaI2VWqQiv+Gh5tagEBpKFss65vuDx1diYQszGuCmCM
g53sy+Xlr1S1AADLq89JbU3gxVQ7vDCrQ/pC+tM8f76UJZ4oGule/2UMJSD0dyabhFV9DCe/Vhfw
D1zBhapWP1prKgJ+Bizb6yMehE8QcqX6GHvtmeSfRHRMmUsHM8dPFbClvQqBO2hyT22hH/iwuNss
NOY0k4kVhhS2HZSFXkoHwWFAiiFM1a0JzUFvs2s4L8N64wKfG55KJyz6u3ng/hWnz370MJ6W8fC4
BUhvk/J7rzGCexmLT1wwbDi6NLjVyyXbeDb1oIKznYUxOvaPUT4cj3EyczDell1no5LRGuY8/5at
0NWhWocp3GJkCW99U+KkEMmSIzRDmmaLOZld4/VkjOzZQ0lSF1hUVx+QmxVR6tSjjDnXTmIBQ/Yi
x0ib2h5D60xAzS/o94a/x3sTEkLxlftcdQjZdZCE+2yvr0KYZyHycvHXAZtEpbVZ+l3uYtZ1V1Ap
LmPVCprdWow12Ga+bPknu6wUFLnL2t9HjU8dRLqVsQAh6xgn02fwOJg83C1rS4stkN5eAnqEr2wn
JY5OXr1jVOv3HbYkCECpE6a+yKItZfNK82iJCy590ogNCKdBfa5odfO6JvpoZrTu1NziZwmL7TJh
czskRk80setDxsz2svK495uER3za8cOxItuOjt/WzmPW4wRQgzCZm95yIjSmwetWZfMFQuf9gX9R
1c7iduFq69hMKSSf+4uDxdslqcpH4J9GnYl0jb8EGizz9QppQIY9nV91o+qh5EWlJjHdbQ79nHAH
BH3DWL4y4fX7XwC2G/kZFaXBan6ZNmh5Z5n9A5amC/dqv4WVUrGiZNyvVvjyYKAyxFmBely4A4NN
iECyNdhTpvirxvl+0qvAzwkgasNJs3cKnwgNomwqxY1LGDipziMrPeEDPlRHvtBA8qZUkZ00Yu5T
3T1JMnr7/mUxscEgH2oCZdYcw37EUYt3JgoQJ8gNIJl/giKDbxWl71Aa9x7MLYcxsIkXuNdVVeOa
lxMrfe5ofBD/4wg1rwkE6sPslqzW3fAtIPE/OI18KXPuQvD1TD4gl0yp/JDAPwp13/RPzEwq0kc0
CFE6esGyJTo5B0ErXRqYJ28vxqCQNxnTMShLw1j2ce2iaxKdkRI2sx1PPwdNH3puQjqC0pI0rS5+
BSK+MGoyksA+p83/kZ/U5qwVK3RlsIWoKeiaOHid0Bgj4gWbGdpFav2uH6APisA4gjOru+ntL8Zj
hh/nyYNnbWvp6+Ch75Jn+Eyr0THiKcI4Bu3y/nwiLIXEj7Mf3OYojLd+jK1pGmVWF1cbjEjtsuC9
IaraExTZg1mcZvM8envOdkplpvBXf7P1O7vDdHQ/QKfglz39/DuaqxJHlhNV1rPVcm/QVBfsoAEH
6HXc7tvT9Kg7IdH92ChTnK2AQZb3m46EDyrsdd8tkUEEVhet5iMqksYHVBjabramiTOHtGBHjFsJ
9HejwV4DoU7UP7N25YENvketCjVM8nnRnwk7BQGcDVgdOAH85834x3KF53DpfBaZnCkYu17GtBOD
qnJ/XMZctUPykG47nqOFGujHTgzqQwTa8HdfZvZ3G/P+kc4YL1C/FWUTIs3kAnO5rRBvygo/nHFk
XElyLTaO7cbP3yo6VsSCwvHkbIi6GkdNetfDB7iLRMwXrpj3hS3y127Bv/AqIZU4KUDaKizFH/A3
HPOIkxqBqi4t36hur6AgdGzqpoBu6LUeMSpStdPh8pEg09kJvvNDadUFIhuv/4Twn3LCGmTIUgBw
ylNciSyG/jGfLFN5YYaBHNn6tWCgz1pN5Y38qkj4k6RDUjb2aT72mB0gX6z7OTSJaU2W1nJJlQcV
p6GrjuLKbivUbAQS51P+P2ux2wEgPNgI7IC/1o3Yg+Kgg4g2W1zkQ067h0966vIPmYDNZVphN8vo
+oSO33EhfhvxWJuy0I9FEC3LeqzSkY5j1p7dlT2wNZqvq+kFkU7oIVuK/I7N9eQ8za+39vwNfV2d
zb2esVa9kp14LzO7+zmCvX5xJ1kNG3FYT76bD/mSxHTbor6Y60HiNg9bz6u2iWW4txVrQHVrm9aj
PAH6sdV8fdN2q9NXLvsyENZxXqMQeB94qRGyqlblzp8sbdqDTEzVjROqR5DspCxlHg9r9IVgYeov
Vu8QU6nDxQvMVMbpe/1+KwC6IGzYGfqoX4QooM3BFZTuL5InyTPCHuQZB5Gtgw18MmakZ1wo/Ih6
HPChSRVRl961z+tfaYazPRo6cckK+IfBHOfAXPxJPvoMoNHYbGBPstTq0ejbwFdX6AiYGUxgccZ9
LlHIycJAfczNpAW64mlUQxaN63zBlbAANqqpdm/4P32C5vmJBUJ62yQSCk+jFlNv5yagCNa+1OOB
JsUNxx+454B8hSXUeIuRf6ewYRnGrYrYGVL2Qd2SQl7g2C/SgO8OeuARrIFGtM6O7E77mMCtQc60
zvs+6vTAJNsFq/JMBhx0JvJjtg95yOdu8orktEe0rxdfnKrv9pAJVybbDC/mANVANy6gNyRec5TJ
CR6htmy+G5iRcgr5BMYIafcZwLorPjdpyU4RbqaUxIjaslMhmFhLC5LlBQTETRZu2isGPb6z7zC9
JvS/TSAqYzHfmWi3di3+h7qBUIRzuzNLucMGiYyftYdARFugsh2NbjoZO4Un7bThdTpPdK84bdj/
fof/Bfo3UuLXh9FsiYum8VseLKHLHrhUPGL4MzhI/z71qbTtqj8ZHc+uBIHSxYsbXmxMmJKfRJx4
++9qnWPqEm7VF3GlAciWEbKufTFLZb4ZjP0aBsoRyuGTWWp2TW4vnhbAn3I6SVK+kaAnOULRKEKo
PMtSSJC1nEaqtFC9AwgbSXR1f1FwcIAGntOpqczVGnRPdNvvqy4FKbH1fIxne0bbor0s4UbvJzyU
YmmxlRfzL+GQi4BmtybZz18bJ2oeXP4BmbuOCS/75qLdmrd/kKdfeGqSnvLH6POMK0oorQ+0wnkW
NrEc7Dk/ONgwXYRBylotIHArQjvFQhmuf4swrECtzJU0iUwJC8gresHiwDKGZ0kU65vag9GvR13y
dfs6DmyfLQdZjm1KUMrHPDfiB/VM145EZlHXwLkoCP1JfrzGTY5MvJDxZssdCwmfARGeecE2cLoo
XvYT2QIBde361XTF+teZW+IwPWk6N3LRAGWTup74Ge63JOFdWKkIL/Y5n/2/IRtuj7AW9DuoZvzD
uNjT5x9+qesBfoJT/KSPrj3ZmHqjPggcoo/4bqaK7gVuekX+bv0mLEkQQvmNkQep7bAq/aTSyJ/4
jxUmo97lcVWMquYWtJnttwXoe+ZJ5fmspDWK7ltFIph9YVnAck/9ubCRnmuHL0kpK1pbtAgaR2q3
48RCdxho0ztx03zipo/N5tfS2Y7C5FhfJskETn61UIAOVyhhHixN5mB0IG80n2fweW1oqRhQIke7
SakYnukW5xjkhxmM/8rqmdRK7OJTc3n/V/cXu1hqCdBMHeakz2gwJHzQCbYpKbf5jrDcQphVO8QU
HWk+quOhV5aJrQf4NQoXeFVXtXSIaP0M1vrq6Rg55RzgiP1sINHqc48cMgJ2IBkAyd0wZ095Pcd1
fCFdYlK8QW8cCoHWpVJrHT4BlYitiIvToKxZ926MLgNFz51lJukEID0/Gnd/27b79SP5meUhrq43
zMBmFT+oWkkJf60sf9Wg+Y1e5z3jbgoiO1crILhG807yAiP7xpeRSDQdzXA4gAcbkVjQIjmUWFj1
+H4qIwi8m2V2d1ErKP6JxsM9gY5hmn9HwJ907j+LAu9UH88CE8gBre5T4VOT2DNbBkzg3vLmJh9q
fDQDwJ0KBzb9x+bROJwl1Q0H+PaWIaJUdynLrDHfXlIvYN/0DRR67y03i3u9OvT4PzARkfcrlORV
GkZrAtF8jAOw4ZAxtnHTsyP1C2LbmE7fttCFkbB7OBsFLJR1PQVqq53NifECTRr9663+cM0MrMMv
C0r/r6Lk3QOh8n2fpOaYDZHJy1t4a3lN6UvJ9pbd33HL2h1iroR2Jzsw2K9DFaTRkhmr3AGMush5
ghbvEqErQ1fVw6NWdjuiydwY9zHBCahp371wDL+391LSXAxAUfFQsOdP8iiFoT9heuVxO9M4UJ9c
2tcFgyH/Vd+CLoFCTlTwztPmlP2qIgt5x5kI7biZOG87I2HtjkFIueY04s0PRO8VfXDVwJvd9HtQ
lGYutjn8Qmg3GWVZOM2E0m13wlzguj3+Q0MNrlaQhTjtwGDiqQVfXK4FIUskh8jJ1i5hCVMQUy7o
hlOxatIDAbHsS9D6YY116D4CqePltggBDfyAwUgRiaPFgyGVZvKTbzTtVEOjDeyG+YWY5YKgkhuh
eI5oeBFwJmLHg2okynCCutHSx7X0uiPbsGeqxDi7OZZXB7yMO5+fQYP+6Uas7w6/Iuurk51xp+HB
kT6WFS43m2Zn5tkIFr6t/VWY0PL4nc7jrbiEwxBzXrGlkNlRZSEebU7wNzuKuN3dQ20XzRINYgNG
v20eTIli9wt6DJSMrapadCKydrVai44YiTBmd+q15lXaL8FTKICfsalWMMrs7WjtRiV/EzHHBvCg
n1s5IEEp+RE99mlCvsPcVwJeASZRqdW90DAgHEiRJA9BuBffadoJH6l+VoAp7gzlCn3nZkSZqNOo
lkWvBUW5390Otcy2bRI37GILG+oGQxUoFOgGHnDscXC1C5ntJCHHySbKyTb/6IGCarq0ri1gWFIH
CnrtG0rt6QYVxFBaAKSEde0dKWz4JaPu7qlVI2Kz9rHhPvEzZ62QPYXGVo+FtVthGUhmCWHxHHEP
D8WwAHVIbs8PhcGn/MTj0YjRkkl4OHDicCg3reKr2mG0XSc0YIkUfDPF73SAR914XLkSeotqLMfZ
m6jjDM0rdD47L0APPhe5DwgK1d3Y1J0HE8kl3T3hwh8MsuSpLnEubu0HAmYDrh1NgDc2lGIRD58/
B3QnF9UXiEaNnsLoSRwcx4yiUGC8a3bBQEgZ5yWovsyQkUd4Wf2d41vTd1OBFeaQdq+xgHVO3GhN
TcAu1ZKvtuHFP8FmrGMV5GLQK6MFDEyOIyFwybzkL9Wgc+UpCTPEKmBayRYEFi9obFrrKaGP0pNk
nLcZLE1U32mPvEOPXHIygvMxGWJ9gJER+8nnrnjLlmKtlKDG3Z0DazVWl63GcleoE+ekRYq9eVWF
zKRyMlppmiOKCqKnWxtoLr4qpqat0KkDIBRDx9LgjTrZlXxuUx0MUKcSDfk157LDnxgPqA6oCdOh
oB7eAJGBDB5CschvzYg8lvZXvC0R658L9kGXDfW+1nahmk+K9GMTfBiKpV+1Kgqx7P99WHucnOOp
kw/1s2FxxPe95sZUpZakvV7pKfMGE1i078CjvFdtNDH8M9wBxgOqZywFHSopuoLnDPuEy1IwFNzE
sKhGXfel81vyjU+sZQZ38vpJ5Sr4NUt48ejBnl098M8F58U5wo1zFddUPRGOLra/5GEpNchfQBUE
x+L9H4z9Vauxah5PRY0rJbAA4KH0slkTsmV2N/f/MHfYKMi61ofhCMD/kdxEX52g9qIKhZT4O4c1
2gbI6m4Do1bAqPMtJZDb+P9WXyQwS6BCrnWbg4oruV3CMbEAfJhFts4M5PLUy7bKwGVKzjft/gVi
WLQBOoYAoDvJcPpNYz2vYvVfhzlFByzabkT+lYwI3SOnhdCBBjCsc0VE05Xjti82bWmw9+yfL23p
p1CdQWgAMXdfDkcLMbTFeiwsXxqd2wtbCw4XGGyJgXElMuLS9Oo4KQu0xuj9At8UWvkF15IT7wUS
ltOoTsZBZBjcOuurRdEBDQNXPoprues2P+s1BQ7v3GT+DazpwyZsFpOAyLyQAICMv2mGEIEdMk7B
jbgmdL4UVzfvtQYwkN3Lsj0plal6/IJHlfmSsy699ed6Fv8fVhEYSU42l8ceEjkDzrmdsE8kFvKq
jLUnrRVPaLQCvRSbFAPImBVot9cLcoeO8EhGINC0si+eG1nv9/uiHFpT/5olwsWaX5rht8qqoIW8
mlu3nL0Ea7fH3xgD1HqBISW4Wf+lJBXelN+kArltcNN+shap7+GpU6wRXA/gXE1m+FLFWSrwkvaW
vQKHnvcjewIHdesc2u5ax4KD5zqrGtKIAGyHtgKpAwptStMH1YtK9BuaN61wI9wFf4D5MxatrHm8
y+yoQcryM/KPB9dz8dO4DFXHsMJwSv/2dZOWRgG9bmVlx6OFdCqXRMwrgWEp22k1wBqLWCrpWF4Q
oOmFoGElHU/4SViZVWqvs0F8didOfka/NEMkLdk5ntRfoxoAG6fnJbVcwiV40R3mK3VD9zDy5GQt
fSttuQb36RdrYxlsE5XpE9YXbP3nllNXKKZ9KUWo0pUIXZqgWTn+6Se/dXCO6mMk4zJTrKH6GTXk
Gu2SPdnzH8KhBLcFrPw8svzT4dgXBHjZODpMNjpECct3NvYlUevAnnRfmduQhcF3FVC2i/f8a3F6
zX6XKCJwc+FXcefEfbYEVlb6ht/y2KZkuY30M1L/KvbXaPIxx21ZAudagodveXmCrPKhyW2iwpWP
1Lh7ELzSD2ROE7iIO1yjfamom69Uh6S8TgSW71wrjHvDUBpBPBkcMTN+Ih4Zrzbjl6QvOkRIAt+d
5XziMUPx0K0qmHGrDaQjrgNcgEVJwPFrTr097eUJsi2P8Nm5VhWvC3YEgGWaVhFimp3JemJ/lijP
a4KOk3zFdm/M5BbdLB09kuVZGcWFKjV98YpklnrLSgy35qFjnUoorfMGUvqeX7kFQHQQzHPWzSQQ
9fwaIk9oV+Zr0ScYYbe7MIZ4q2+0hsdMYFI63dsMiFI44wE6wFpCellQupYWEFTuhaADMxfh2me7
+i3ismKAwleATcdNZYKjPxtLea3wWsSUD1s5Q26mkJEo3101GxYEfISxnm0g3n7VVcBsm4YmlUgc
KgHSjZqTlLKy9zvoZxv949h2c9Xh3pYmDRgL1LBqRMZN+29Zr2pWQ4yuw9ahcZ5+Jj696Dpy0CxY
+72fpbVY+me4Tmu8vKZNsq/Y4Bg9qRch+DeoEDhJyc7pQMfbT1J0YL8vqdAiKVIBU5fzhk5xJKjk
Ga+W1CfGygdSI0bifWMxT7EqH+Wkg3NXyoEWV2kkO3Qiobey4868EKzbnuSOVRcBGeB3ery5fkJc
PD4svCJz1/fTxCj2PiwE1Im9f2kb2QXnqHOh6ohTUNqTaHQsW+LnQI8s/OqXBG29LfMy6XG3CE6F
ap8bE0R5lKbxQNZbDHXFv4vW8G15lB0neIhRpG/i4+5jmPwCgU82MQrVGknwyyJr3lKGz38TCiKo
GWDitf5syeF/iIsQzUsEVpIy6YdhcTzxiCpUrF1v28dImCpKVPTAfWKsJXPo2ohCbaRFYbWMoqvp
oYexLy4jJqh5vN/ZJk2nTwnntyDUMP54otC8wiCDxnMBNtfeODaDYDeiSyST2i8v2rnOi08UQrAp
HYzBcw5YXJyI6T1Y4QaLJ1kIczojq8fEugUAP0fR2w0MNNApq1EDQttGf5VC2TdLRcuGvEEnKKAm
Uvx50vKV+rIHcG1RXk0N715p1jUMmZvBKFvwYzxYG8TnAanvyulIIB4dwJqcWjj3l5wss1uGLTNS
M7s9dwJ4N49CMQ+c/OB+QpqiymNCOJhgduQ5KxeeqS2SJvfX90EEU8MBcPhCZXYFggS+YctwMV7p
ojllsEFCaNIuOjxbcDFlRNuilyYcjRMKUbLwAcn4sBYbndGKG78Y5ZLTwAnJBJrrzTafXcfbCJGH
XYyrzewgO5KVO53oo4IXIgCOpAIT27wrrVIULA6pRKvCpyn8LPn14HrqFAHSqO5xfVsRTYyM9G2y
7y7b6txzGpvjSppbUy7zvxQwhLzaHHnG03ST16egqi1OWBV7/E64365GzhquNsIoIrx8lExWarmH
ERIj6XZdNEw/9CzaAMS51dPBZpB2w1sy8loVmD/BAy597dhJRMvy6K4qmEljn7dIgJElbKB+0EI7
dlDwS2QqRiH8iAa2fjUZ26vbqVxNTkF1tE1K/mKMEXRED8pows4eUDmG2NVcZxTqJxh6GK687CBo
BuQoXXLkcQ6uwoRiame70BLVzZvdf73IOP/rlzitrgEPSe2V+xFTBVX/eEEDYYscv9iYNwc+nK8v
BsuxRjfy4oEle8e5seRTmyvWFN15v7OecfInj1w2FVCoVAPUjuGGa4cTrk8nUvgU6+eIoMdVBjxj
q0oPt4c7ndcRv4B8QYjjqb63/EXlLIKTbb9A1QSn2fmYxshI5KnprMlJUZQIDShZh5f/d0gwKxtN
JyFNwodGbjqE5BkRYeGKa6hhZj5Mhgm/KSXWPfC32LAaVlQOu3VI9M8tO3reip41coijSrbyKJWr
LUvKUdj5KvHc3cBT6PjMky//4pKQWkl34PeQDzOTf7kKg3cn4RXIUgcxtUEGYE/p4Hvu+RF4ZatV
OKu3Pj3vcJ4EEQz7y8d31QFitOsCBQIPCOOHfASSi0IjdqfyDU/WbeajPZUQh0u0MQOFdAFmMTVD
ZkPcS8rKm6fFAsQg0MExCfyn6+8TwrI1b8Hj0fIxQ4tXUU6cMRtBjq/ikZLibLd3kSX77PisKBnG
nma90P4ygQEoUMCCivuFGAS2epWF+Y0EG02fs+KFTauldtsX3MrcUu8rtgyCV0tFdC73+DxhVCd1
ma9Xc9xMR7a4FoqEKiL0GVPxD5iJ9DtzLy56JTPMRqRA1EFyqP5kKwIDUCtuNxqgEPJHBgB99f+f
qcm8cMkYBvjXNWta+SlKHWtWcaxljyJUmfHqSya3TsCfENAUX1uRvn4stKH9s4bXi2qRlMZvN7Yd
vUyy6OsyMmP9mnY4v/B5rAgFiiGeGyaBfzgm8tZMnKns4n+AcYfTxzilN3FlEBrSQzy0rMiq74+1
T41hmY8tsnsQJgHpzxn4MS5hATUVoR8JmFx2BDTTkhB+l7eBBy7ck9zATPkOxB755EgMMvwgaadF
xDH00BAROTwzdy+/76y4MWXDINCr2IFNhoVYGXmmYM0jFZjqL8SmZJC/PakL1xqi6BbZkWLOeOAJ
VicyIxl7UEM/FUhGRuFxd4eqDwWLyZ1R6SsSC1cFbZOSQlwRKMyhh8uoxT+D9wP6YMPj5WUY5ieO
A5sbty3P3K2Ms4iM5QWWLhshhj1R8WCu1KVwIDYGRt/E65HzW8MjBx8qnLvpYJ5yBoOT4+3glAec
L2vbNoxdBSmmkygC2c2STqeNsI8bH/QJB3CvLlDz+U0MfqTsDrniWdHgPoLZs52vUvmV9Vhy9dVj
l+tndHRCedAW2tfJ0IXQX5INcawvt26pJsKIvhBSuMEAuWggjFILDI/MMGARb2QB4VwUO5j2M2pp
gewZSMsn7Ot7qMgvTgdk0JAaJmrRpt909EBqyfStFL8SbEeyR7hpVYqTlNcwpE77/MLQL7CN3tZE
V09v/xBIsLvbynanzmvm/GhlN6uVROMP1I1tLTfXTTqA3fVCZQ2j03Y0F8U4+Pnt7hZt5sRrDEof
sI77gpBE+tEPICIMRq0V8Mb6Vzq/i65v0W5wfcN2byH3lBDWvK7u6BcLCsSuq/cE+4l7C7rmK38h
ifNVfX+DKYJZJoKAcSliQoeu0jlQUcp4aKWqlmSHVm7sIZnOs8YqeTa3lpBqnm0ajosnWGVXe7BY
1MhRFAyGq95zcA/2LMn8smkgR6sCKGk2zJznb9obxCuo6VRyQgKPt53hQF71OZAGQAjM/gmAB1He
BnCJni5iiZh8nhBSY/zGdWd4vc8fwb8E8+KzehK7QHdUAB8tiKpOfGCI9aVsAWa3tbaX1qrHfxDV
CqNuo55hpF+joRNcqwZ2CsaPfCE7zMNfHJz39ApzAPufUb2NkAINuiQjUzX8k6ZtcRbHLhnugx/e
HN/RgiDHmMW311GVdYUUwG8i7qglPplFNse9OVzdm8MHJvxUEU/Dl0da233sih8C18EzHTZtvtVM
+nywjDfZ1eNXMX/K0G6wLQ2TOHcayrooxl2jMJs+krYTib7uIxQC0Uy1pmEm+XKdA0PGcEQAhS4l
rc6tlqyyxz4GjPKk2IFVo15oFOlinvKC7cHthRg5vR2TKCLYBCev0l0ASb8jjAuvnaYBVw8cQjfE
03/D6iTwpFUmjxnPJTfKFEfmdvGmHGEfvjdqswIjCeIHr2L3fzGYpFZ49YAQttnYMr7kqKeK6iQT
/GItdS1liZSyEgty9AZrDcoP0kU2T0NEtzN4j1oZHF4CYwZ+qTJrxTaeBBsWuaXrm4aXdqgGUw6O
H0zihO3hnD10+e6v2G9xkkquaWlxsQbIKSalmzKyd2BTGfYeWjSAwAeOvSJoPHRd6XVC68gferyX
dnaDI2tz8qNebTztwqHIoR0TGOiW6ztrsa69JjxL5wVZcivYugPoFcMziAqEP1zXB1RgkKCvJS55
PoGhlhvVMS19f1qX+tTySIwdsgMZYps3DCSS0yec+nD8GcaB2l7UzuqlBTeA7EL54X9UsdohVZJz
kTD6gAEj3ZGMAypHdq7NYQkN+VG+BuYh5zpNBsl4oYYHH3HKTinl1DfGlIqlXdL6EZVca3pViyEP
cuyYTjx5px6iMLs4nLuXzh5RD5MBt5Od3RRiL/7psOH0QkAy0t75jx33q7IXSH8zISsn9tImuFTl
yj6gK5MqMKmN01bnHCpCVNONwnAzMOLgdtCF8PhnFmKYggsv+umqYrYwgRKmeAfzf+EDAegLeQbP
OmKuWxfphUi5YIOw5e43457M3SfezfwDjTNlIEeTveCyuIACgtNb1J0sZuNJkEbyAG1v0nIemaM3
WVvW92Thszh21PLhryrbrnmvTyouzNnQwE//9Jw9B3niRsJ4hDlv01SoNs6EgeP9yWIMc5KwNG8D
PM0DgjRLwCt+CHVUgF4SCBQW/zJ3n4hFLd0xwhjBI7jR2R6/AEkMP2n2pulRvvJnaa1o96o0xtog
OgdK/6xVox+UHhRqK+xFklMVItum77b3tikJQF1nRdFjtME0ooyPe9cvWAlK2e1k1zIQQL2/4n1F
lxNEe+Z3v1DfOF+BL2Ou/txu4+xiYoYNo4COn1x9ibeJhvwH3Mm33UefHwtE81Cd4CmT4SkMAC+O
7VtrnqeNojF5WF2IeqLmTTaSVbs5hhn9Me8h2uHOtGvB+XufMJmwiacOFiGWUZObcfhZCZghj5mo
C/y1CFBqJhxldfpqLbEsgv+tOSIcYWtJ9j0fqukymny6xBgO8neo+x6hCOqqd0rJQzAIkKoalqjy
jxKY6XvULyu/WMxVYEV+OwiO1iThOdold+GUFGEtaoU8tEVhKcw9RliYEMCZ33hsa+qhStJgqM8Q
vO0vuDbj6uRveb45O8ON/kX1jPHq+qOTsu83EIv2ifLmhUmFhtcfzpdFADgcqVjJSl0EZC852w2+
W5zaJJqXca8gGrj0yhPI7z+2FB6txZ7GxO6S6vC93PAMOdD2thK3QqM8wDH4AuhBTEYsKcfJOQw+
9CN5B71xgLBNEWMNING6UFrj2jpi8+NTFezDFQZZtEUD0xgCvmSkysiAKOki3XaTqMdy0koTo9nd
tjGJb0OLEGlhLyXC5Yj+PKC6CmS7an/FIh+hCePuIO5rebFL/++cjJQM6toAMQLYqctu8cK1FmnW
bntx2fNhhLxJjEvLfz+p5ppHG9kzb3cakzFfWA6jCzu0rqvNqR6bOyjnZQXqYOzQuivM+VNWFfQ+
3aZzoPEKNmYKDLwpdumGXBNw6TALM7/poJP2aldRYQG6/whmvQ3Jc4+U0Ex2qnffr3OSXfxIY9v+
IzvMVaJr5uEJYsZ6ZacyrvMAI18w7pMKIcbHAPpoBtde25w4n6tEpCx21e3LYcPuwaNLfs7P8DW4
m+do7YsSa9jLKHo/VH3TEG6aPVdcigp+vqVY+LDJZ0AyEtqBDzdTOLuTAkcLyoQC1iRReQ+1Bj7M
XCehXwUtDKdnwzGlWMfhmHczcS0GK8dVMD5otZ3X1axiHnt9BxXNp0EzDYtE5+COvrkisAz8iOGy
cYZeQIyxolhGDmEWlfXNEP6go2RjVcqd6oyVHs3Az3n1qYrLdnypO1LGM1e9dS57c+Gra4HUBAvd
cc5IGTimWmoUFYwZTfUrsCEGqtsaca1pU52jm6IxGQHVs0Ch70s7n9iy2XFLZCfF1WL0UJJGpKzK
EQiGpVcnp1eyGnxQTkqDNyS169gkCE9allMX6clrHrqXiozLlzUJb7mZDcHFTqAftk+ljOL6MqPm
qp2AVNWZMhJ8KnNTfa6efeBWZ+xoBRzNcxTXI44+g4pz+SPHfRhomFAXaR2tRAa+dqK7yaBcobZP
fhgDuDL7xyKNAzaFevIpxHKuVPpKina3UQ9RiZVy7jJiaO2odCSun/nQyMsx8MLQoacOVI8wC0MF
l3P+NYdVDq76FntC9Q3dnDa9Wr46ZR+xBfR/1z1unVdVF68gdZMzhUw9UArWx07s0g2CsY+mTaCr
lUa9XcFCtirMuq8eiHAY2BNxflYv9IRwfg/ep2ZCRkSXpyIF8jOCTEn/Yhe0pYzDPonrnUoUDDxl
K/EG71Hpo5SQ62MowCVim23AlVs8g1W8+jWS+0Mjj5OkABqrJPI+8NnUUxemKknllv2UFddx3goQ
My4PYirjrD3ok2zWz0z0l49qRS1B1ZajLJ0PuwAkOqRWdraR37QPdrUwcC5Qp/+IlSXwvWl7zVG7
Kuzl2aM2uq70+UypRVJAHD0SJ4NTqNC2zxVwp0icDCwf4UhfoOtf5ZMnTNjBZmnKQ6BRC8ZOz2MD
1DpkFHO2caItbBshyKONqdxOgvkbiZZUlFE4aYwagKMF0ARXkhPw9Rvz3Dr9b2bqN0ZHbExD6fDy
2/goWa2NA2Yu5CNasvKTDgb4CkSW4qrAnoZVtPAdMQcUUYv0j1bAQ2Z6AE2M7x1ApiSHlycKAwzd
nzx0xShxLl02AUw0gyITTxMbGwD1f9r4dNfziniC/QTFGNOAWbfZlBhYsyClWjROmNF4Ut9+1Eo8
mWWV3tk+yJxwjnLckFF98iVugKLZS48inOcHRe4TCUpzvpW3Cd9qvmosEJrK8Ji1AbMPDWzt9iQR
q6ZrvHYySjMyvYbLeFUeQDxdMPzmq5zaLFMBJfMvhS/RIorejAHInZ/Polv1iq30IPpBIV/p2LGA
UrKx54UbzZeEAV6T26lt/qI0UCHsQkKyvTSjjeIJp2J060pZjlGhh0oJV51avsTkZ+RUh78WN/U/
oj5kbkX0EuaBHr7vXWZkoO2/++RlCE/0DJROympG6m8UrZsH71Sw/lkdQHdV+8RO0OhFSgnG9iiP
9c3nIoQGUNa/jUGtIl8QXHaO2cGtPfZC0/tyljnTLchr2AIjf5pNA8ee1Bl3W11/2sBn2ya6H9bw
dgbx5/tlwdvMEY3XnfjezQmXet7FL27UCZrHEKmDnQHCt5gHSqRvN2jMqBIX+sTdD4qaWQNvSCnR
5cwUeRQpMwKPw+ExxH0P8w1uNNXAOY6qNql0myzHqMnQs7LgxOFkTSlpUq2V89CzgTl7awK9sEkw
3dYh4aSvxfEWcrtI69FyNymB50gtF5ZH0YeAWmwTE/fitdhIjI0iK3Kz2kVZU2tc6ksjSCNgt7kK
0OjUbvNUwuJO8tvZAAxiegqjcVlh+p9npNOSK5EOWpl5InV/KTkmbPG5RrKNI4fw/6jUBVqTcUfv
oPj3Lb+puKvq1TkEqauhhKIvprZGxZJ7ph4dtyA/I2lylrIqXEUKahDY8+TMSqw+aVirTyjT5f83
mUVWIMbx7MFaBXsKQXfYQn1nq+rqGXE7aBGOQgshcueAjgqD1gHu7mpIvT8XMcJ1RqM4h1aWpr4F
OHw1aV2aRaj4odYi8MfH/QEt4kSOQ7+uaeOnachtTJYPkTnH2N6OQF/QyBPZ4x5vn436zPYRL/h3
k+aNv2qp7qXudnPfn6j0uSSVoRnfUiEtiDvx6xgjGkrMxVFhl5yfT8dtrgKkqu5swVCokZLiYhTW
VAnwUFDD272TbA9reJVIkWBdvCUOCWHSpLXxtfRCJ21r9/roLRTK1comXPdbtca8XnK359P7ZBK+
FROsAi8/A72dGhE1Hj1Fg9OaLZUxgXdtuLavrISWVF+iQrmF/7V2yAmO3K8CXC7g0l7WWAhoUQVf
75ns7CKLRiv5pwab36EEY/ckGmH46hPRV0XA3Cu72GEZlg7b3riFKXEydbw/buVtmh1ijGHmsmOR
Am6AyASDzh6489o+UxcQhi68bZGXLM2boHh1y+8VjwiQCluQt/AoRSXV4EbN64+zgNwEOyDYyldb
M2k5buUzA8V6q5TKaRwlzx6ajvFG1Uoiuv7U0Jws0nGXgNjpyKBYiDWja6QPwayMy09pqrHHoyH2
94LWBsao2uCow4D/Z/a4n7En/S90VDipD4w0MpNACHv6LbTVxPxtLX9IVhOb2hbryzfOSUpeFArW
DiGfQDbK8E9ASYTDeUm2pFfpBY/1V9b0wYooqPcMAEQD9Q7tex+y02qBhJNZuN/dp6ctmCRUXqxn
4RCGrp7CBhOematrXLgbUa3w2UV23+LIoXlkfb+qQQzQgnnop3XgCON6ULQ1WCW37g/Jro00jCmF
Zt4DXyQH45/m3B7MlDm/ZxcaCm/By7bMeyb6pFzldOGG58877cAjJzPQiFJ3lKI4ub/rabEAOXME
jyNZEqUVvHVhr8rJXMSdBYi4VX7BGRU6Sf7I7Px4z5DjNwWaWI4az6e7JTzYg8vfUBjjqcaCijOf
sRdtYl/i6vwdpyW75WO+ltM+Qbfz1co9TpkByA7LVDIBKQoeyi6k2UqH2Dn5jnBIabFQKEqHgfcR
3CCZkUaJqB4gfcBgRLcZnXOlC4qjiWBCjkyIMeJznH9gSGXtZbfoXz4RS716+1DWk/9kWCS01ObP
hvVADQpxMR3lI5DlLhqtJKzrHWwyyDScUHxMiMZTYkZ911CFwmEas8tZuHfm+t1u/YGUcH04l0Nj
w2SJyLMj+O+Lm5+H/0x1ucKPKFfTj0E/p1l9F6Ys5UZFscihBUhG1Cxw1UQIP3SWRTkf/8yXcm/P
xy11xHgVhQDqskMGViR81Z5nkO9Lt0XukNqOf6JtkdnBkEah76RsrNNORhyAymS8JGr0Uewqc0qB
KZhNNt/USWydvWo9cuResT59PI/RP5bksABNiXHbZCV9qclJNo2ZA2hv7lQFQd6ZaarhW+8A7bGU
5dG2/z5v/WOry9pGNb4rUGH4LzgyLv53CiQOko/n7JmtAPM5k9NGqJMKwCs8rRW8Ktadd3ADpu7N
r5CL5aB9OF5jxQ+Rt4E1iHjKqQrcL/pDeZiZaNAijh7E5Gzs/ut3vvVFI0DWwHgPcFoYabNDCZuZ
TRlckh5ZAxtfAFDXmtjZ90BCVNtFpkDUQhHFgu6aAjQQpRH7BNU+MeA7tkF+2rjvHkMUY4A8Z17n
6zysknp07vvEaoLL3X8B774UhwDLlDzWJYGx7KJ1BYRx6gxunRN854XRU/EphkVoygxLlRocXzA2
yo5IBxVYKtRDPSInT3SiD8Le2koDDkJbaaIkpaBT2w752nSali6hJ49/QWP62hw3WLq0fsJrVIiA
UkIZ7sTR/VJnUDqVnReDo2d5iop0yC56o4B26lQj86NR1ZnaD1zlyRirf8eit8XEJhChPtN+IMky
6l9rMIDzV40HULMSlT+StyO9fy29Y785+Hy/f+vK6nhgmNfOLpxhZFZNE86EprZklLFXPAC1YXqf
pqHCGIrCb8z3WToYrC/88r7m30Z1PXhX7KGhaQ+aORTma6mV41Ftq4NH7KxnjVJ5vPbRKPz8n5iV
dCGOLBe7Yfa8G9GNUoOqIwsElOzG0Pb53h5YqbkMLqp3ZS5pOFJgkKE4WUq6DlaV09IJNkZeFYxv
E367Gtse6y4c4PrZbPVUeMTXWfXnwEHxafK57IpXC6BTYCIIPbZI9PWrENmDjgi5BO1Kgol7trwc
u2aKV3dpcWC9QjaNvoHBRRbyiH0tkLEySsrnKqkqvhclGMzUO8rH+MWTzI7ehCPoE5U2nbwU9s7W
og5TwFvudMOItt2hXyOA/TE2/ze+VTE8ukys8qaOVsNQ7MdtHcEg8Q+/mumRovGqa2nSgdd6GbNy
nfylR98ElKk0rgwTeVmtz95BoPBmhxMalbgpK7jGkcnqvb0TUMXZqr8AwW0z4pl3wgT7LZKMQKDp
sBg+YEmj3skM7m4aDVmIscs4+3mtlGGJTH18qK5LaMmfNGlA7hapJsDKqml0ty/EfIa0ghjN/ASv
q7kD71f/bB6khOKxWcAdhbAaQ2hK7GiTZPWuCZu8dKUXWfr0CQLwvYhHzxfidj32Cjhhlsg8KOwd
IjSWPXm85FMmFRhwiT5jPNqXlLFYPrSZKTwofCY3wbQdKr4seintEY0iKrF6FggpfpVTu1mXnPSd
EQtW8PzroqszyAy81cEkrbUO1900e+Oybv8JiakTvypTU26hC9YNr2eLIppNrfY1tztO9W5jNz8o
8tmpAl0ujN+uAludmIJO1W4Wj9EWuEuDdt6/I8/NM+3KTLbCf5ZTRMR4MK/UZ42UYjwfEOSeaBTw
5sVxemjvRkIsduQTjduvP8pAX7Lvaomja1CjdAbHQ3sYyVmy6YRqqSzncxaVlqGV+mby4exrljBP
cqnCBIF695lthK5pNqK7ddNNWXlyFPjd24vA2TGJqMSpebis1GIBQoknYLD4ZHKOb0aPYtD4DyXa
6wQq9I76HjEL3LmxTFE4F8daoYdbKpqjpenvw/M7QyhYSvlshStEPOlqo604qkEE3az+eN3n5ofp
b3ljW7DbjbHDiUWgfhxezjlEIrXAMc43nvXhhhxzQLses0x4kNjj8d3yfky4D+INZAoglfIjSlFL
GDQ+rxda5Mv3RlIQr5Ck7//LHeJ1Kn+TF45qf08EweQ/oIQsUVYDAOtvzY2jZNwC6PRgbsO8RuQX
W4vP9u8B7cobQHxVBTA1P5k2uhz/clPmNsCeipVaLHyIYYUKrcBbK7l/Mcw88vQgOwfCqBcbwcGG
l2iuN8CkceBRcbfh3H2JfsXMq4hMftpY1srz1hPsOvZkS5o30XdBwUbcsrI0AArrY7WME2W8AFVK
GtyM2UDSJBHzTnptvL4Q63cuMbgoiqta7ayfYNMsqOZqTd//pG3pwDEPQhN7YHgBKlNhJ7fcQBj5
xapZAlQs17iTyzTUAXkARppN2IMiGRM6VafA9qy2y96B2HSXzMM86EXdLrnMa5IZ25TX+sOzEE0m
D/olk4pDpCaoY7wdCLIfuKdyZIujzdFPCPIsNcgMy8X8/DDlElyJHTLVTZsBCWm85C4Fez2L3C3s
q9t72AJp+Btv/zHSlJTqZBHhgg8qBFupdrzyRbrB8MgC5Aah4XnVUdJSWs3IPrBZMegNnNNqGTd5
WAuGEPxFBM7izuQCx5htH9GWVHJPPo57VXsFhdZ0MxcuNpcMr3fddWEQhq543pfc0av2/hU1Wo+N
v2vjDygdOg65QpfYywQnVVLQGfznKF77FV6awNwq8j/epo+7fJCjUWEB0oHRtjZUCpnrbNsnLqjG
is1eUi+heCKEBa4XsaXKAo20qHIjhAbhXQ4+/UXSnrQ+9zTd/HAH7N4qv/UllzvtVFLUl/JmI4v9
CJ3HST9uUKURn0rZhVPthRTye/B+9CmPgWsDQMk3uDd2/u+rsI4IkbKI0zZyR6Zkgv44piFPhQcj
amwzoXaLCnkdoT4fpOXz/F9KckkhmG+2Lmxjh+ymf7b3mSV1L3QuwkriyiMfnyWPhqInrsxCsvoz
6j1gkTTwHPHXlnyEhdt+ZIEV6Owye04F149Qzn2lfLYUh/ZkK8V6w5QEUW2I7yrw/BYRULtqbLft
uCEH7ebh5bjP7Nyusvx9uDJA0d8CehOIfSmcYTRYsACRz9x2X1U09eq3KMORaq68Sqki4HxE7nTT
SlFDaTPLIvSIDD1FuG9xukEzJKF26+1Y9PVHlXI1ZG6aNwdGsSY4GF+CDWaX0xE/+foEY2SEAvzv
bpK0SVMud1lFvKFyJSw3G3k452SwpAbm5h5+xFdN1iC+x/3JQ9KDEBxS51uotuzkz4imMmhvTHSk
HpTln3HUynLIC7K1IEOcu31F8LRvOZ9h3tgVIyG8MeawWX5a5d4MDgBjvCmSfx5JXamHroyaPtne
5hK+SGbrhpVfQatqYhJ/fXyvOzuE15Xy47XgGzkXG0mBeL9leffUR8b+oi5pZIJpmgrGneV4dFTW
WPG3DTpV7JlKGGh+slUsQ/Oj0mUPy+SWZdRI9NynnMzfiQ+2/3gSs0NyGkEU92E6cfGASkajrk1M
QoPmb1n4qJYGeZZOrmNE7weBB4TRhFtxh1b4bkDPQKDFPLH8/sz3G+Bqy1lAH5SOuCP8JWX+RyFp
zZBVod6MASJkhWrfKDbl3a7wiWvv0RRjYyzwCAx/60CAUMr8bBlUTQ2oEW2QD0V5p66KDJCEUcTE
ELTL0u9FPFI+EKVOgFIabH8y8WJ3tsDLXs185R7E3ztTnCabn31ZIjd3pUxshBbTI8JJhL8brcdk
FdaJD1GZRst3pUOgf938/wWllEy1L6+h7lUqSzEHlm+D+caDm5FNiKkuWQksA5DXK8MitEPtwJgb
Pev55g0+wiVsXmCw6RAWVXxzfTgAbDnpdLczBcHhjj9Ugb9bSSH/sS8/6xVofwbXn006MhAdvISA
sSFvAv4HkRdwwJeqtwha16fSTSoihMLIHa1iY0YebCD7PW7k72UttVbTCqCDq4Ogya9S+yoWkAMM
vTQrDScBmfb6rVLGSXq5xfX9MyqWcDfimKhnmEK2JtLzStAUZflv9/ZJfSRg0Ehljj4NwrP8b+zi
/LLagtuUhEEqngZokcgx2olfQrUDzo9rW3XAnfCFhouYg/qJ+O/09ciMzugdJO7+AvjaF2gsLJ22
m9The7kG6xybMG965j8UC3nQiIx4qztzvXyO3b1Z+GO31o7XD4KCkBvf6WH9fDys2vEiZMz02K0n
3IXhtfyddBbV5azPkwaLjIAtXOTjEPObQ5FdnBMaD1nYKJBSwV2f0BhyvTQV9xRoFc+5vRND2Yq6
RtMZSOJ/0rxpMHwiMIOu3LWOQc0mKgymrqrsKiFY9h+FFcfuLuhiZvBkHAHQ5wWYbFTRCiCnU8ii
katvUSQ8w0ocMVWITUC3iT3Pi6WU2ztsbfkvQ8gcDEE95rWB+EEcso5DmF4a/tJsjgn8t9kit3P4
217WEt5Q5BrqQLgLGmHqwBFbIpeJv1VdMAn1NZj/sY05jByOup5stVznNrW8L+X712SC4RsGtzL6
Qk3pLMTcNzkJpdjLjBEiRu83cCR+k/xWs0Fo/rjrczFsOKNq2AMf08BdC2vU6gDJ3dJAeQhJW1Yj
A8g5wNrdqg3mZY0972YqFQuxrsiNUGR17/mQJVX3GYyAAv4msKc8qvMvme9n29sEd+wsEKcoeqfb
5U0fetxsbYGXY3cqBrvkhSoHVHk3REJk6woYjAbXXDYi0xW8rDjRgB3MB5CxUJx607n6ZFnCs+fh
+CDzn8nbV258vBLCjj/V3PJQL8B/lGvlaW0ndnTc9iySwmg055x9DMEFBTq/7vuZby5zC1Z2ycIe
NvEn5vMhAdNzbCFAmqfmXj2VO3ruH1yPt2lfNPwEQtm2OGlAk6HmwL8Spmj95GVVAkUMz2f3oAOc
e49bGYYLkm7F+RTl3gGjbR4N+rqZDL4w9UbJSbObLunSqffiJOgPtAnbYLddHGhjzh+lx/XxDxNl
LzenF/xzA7l5C3EQUlmz6fwfzq+2PReOFbjX6h/DeQQzIhfQjjWoFc8IMXhP5l3EVP1iKcu2YAOs
uSuE1m+dnIc82UkSJo+8xelSBDLg4z0CTi2ltn5kbqHr8v3xEgSSQvlHvqME0dM734NMTSZPgLtF
Vv8WMIMrGNCMQGjonFErcse2FottgrFIQCz8ma4uCXm7JrhqSztviXSWhq84GlL9EKEPe3j79Zoc
lUe056CNEF+bYHVLCAyrWdyV8JGyZDrAIgeZNUXNVHJaVnmCv1xtJRkxr1Z4ZsF0Th9OR2q5B9/m
0YC92/fk64n53IvRS9XakdkXZIazIcv5bIh82la15etumGXX4bHXcu9Wyr743PkPCPv3ZoNqkOz/
ENrFNpC92Mo4RXv+yYvt5fVHNs6laODTpXUQb126EIvEvyj2BhnoGBXBPRxij08Pus+tJdNtiN/g
2NIY+cbibOP1LY+voABdqXmZgPBRCB/Ax/fZTvlXeNj2V9/ZoAfiYipFRvwi3kIQYveQJOqh1fDl
2WmCX2iaAFhyWwI1DsY9nkzBoq0yvzN4wMTbuf0/tdtFWvxYs9CGpFpo+4bf2Yji5pSPKsl+4sni
CVmRt4GLFId/08FnZz0B6ZmWtcX/+GvkNAnBV6+sHjMOiuZQR48rKc6UQ+XFXiUEEqVPvihaV4Vp
UJ5zNZvxfCfX9JD0ziGO1TRMZltoijLictMGKmasYvyWuzZ5mz6V793KjCPeaG+GbO56KFUKlzWM
H4FPXDpoQC9HJ3hCs9rQM7eTSga+6w8B4sX9zRnVZku8VodEaWJY8eUzFzIu3o1z4Ecd0cvZK4UL
y+1+othJOXI/5oLBemvWfiIqHTqKt7IC1CicOUHAbRpSQOPosJbgVbVSjS3bM+4V0qBflk+vhKAb
0006AgBKpGHLd0wqDGPWfkeYCM88fzgSPtz9Tqs1jQsuXrRGSjYrYLbBbVf6/eZpYKM4d4RTmFMs
e0AQZqQzZnfC8r/Ix/DUa2/CR1AbYh275zRu15i5yIDpW8MFpaQNFSGSMaBIbSttCC1n2zvvOffL
+ZR8ZvHU5eIL9D/3rUynj32CUpR7sUVvb8B+UJE6XXqi9NWC8NRm+SjWJhcyVBFvvuulxseR4st0
mK3XzbiPv6qYZL9qTssNRfrxO8xVuSh42uWlwuLM39GISg3MQBM6OPoh9xe1uPFenspxxomTizmF
rA4aAy1mLO0JiZugwm8c8xo3eTUKSiyGyUWM7iZVdAIPACLvS22GctVb7Pp4geKZqRsc3rKQoP/y
tycCzjuD9CBBsRPcZSyMkdeMDDEHilApxb5ORjeXHPZ+Pm0naP0ccBuYLEEEmKzi+30Qwf5EXuhU
equcjNAn2KA37dUuSd9UxHFg3KdkdxMPb69drKhiMSVgSGTdgB6/ZeI/HDMb317X6G6RJCg6THF7
8LtH/Bf5tv2YhGGg+p3lMXidUkD7H7rXV2763gQ64uAzcBs+0Rej6ND/LZKEq02sPLpRUmOQYeOo
vioTX/UxaKfjXcseieNL0KsO5d4xANxJBQJUfqFuBfpoEBmOxLSetjkbtpthr9rRdEN7K/6a/sHL
LoA/abDoMyKR4O9KTZQYBVTW6iy5mRE+yyb8GvG80rRMAhmofomfasoPNfZZaLHY0JjRuv9Sp95h
MykAMj1GIZwLaHD160QXgAsjDOGdc0zXG/gTM3nD+IDRt5B29a2fhOzu6/dayvD6TMZK7v7ID2vs
uMSWpPCBX++LhAnOV1AP3Fi1y4hc3l76TlaNHjN9v78piGKUjGJAzAx7rMqi3O5F4ErHpB7R9DZ8
xXedarYBuJAIft0Gqh2gtiJ2aIxBlVRFoy+q1iTNQVaAP1lFZMEVpbVx/SG7IqJSYMiRGai41NLI
s1p/PCdI5vjaQ51JMVtKn2aLPsGi/ALhjjgc7sp/FAVj6uuK84oCBMLOffcr8ZkgRlTrOoXOET1r
a3NWFHEPmViHpRHmmrUll+nFruAVAkTtae+4EAoLBESrmEJkFeKD8NpLsJNgQzsittMQNjiw6Dpf
y5tPRXFJZB9056CDuENc3OO4ZVI4bfVKEQSsPHmy9FoktUmhyz2WOl5ejI2sf4ENs8bHFjPJHtdw
RIMO6sQ2wtvj+EmVrHyQfaNZff4swZJXESUaWbZKvDvYLGb6C3nCrUg+vkeH3hRHpOrFx7DEo7WL
rF6uQuVyrfjHpEFIsrYu6DmfqR2tZHqvVvOliYiGQ7NgYD30hEg1mvj8swYSF1fRlY8Ehjnz7TUQ
es0vSSkJGERPs7dg5c90jCoNaVv7NpMu6Qc3ZoQLItVyY2zWFH5+BijcUtKF9Mudlz/4tNRs7SSI
ruMC2QySrwYxxM3dt6uMcbA4gKsqr6KD1OjMagVsWE8P0aWCIWl7lRdG+vE5YaIb11xdhqwPlpcd
13CrDsk2Fmf5eylSGixZ5ENtPPEYk6D9FdUP4o/3eXeFN2mAuPYNYmlXMWjCFXmogIYqO+H7sDAv
T4KMzVra52fouWbpNb0sP6Dzy9SmJbO2884Uzc6+A9YkNhgbRQXYsHsIgkiNuF4NOcs4mxCN081w
aREBD5b20slkvqHEQCx6UIvAL8czAD3xkhxp0FQc8cadOdi3oybUGgCWuEhHscWCl0kBKs7JLs0W
II7rUD03GjMQtO+W9WR3jTzwGnh/edDeyirhr/DWedDXw2x5N0xqzSqbeSVqVERGMSjm+O9ROFV3
++31irlW/hmt+2wyERCTFuBcwqeD7o5izrvQdDUCmc51q59eYuNsiFsBHeX7DFY1FB+mpAAFtY3h
iY+yvh2bdcSFxZJwMRhEz/MVpUa31Xusu6TFQoWbUyl8xjsC7CWXI9SQfZ7KyxgjImciMa5bk0MU
9ZRIOLSdYxYEEAp7+mEJ5hcAIId3BYoRvfpQEzKKcIymTszIQ/wp7nOY3l2wFl4MytrEvylctrKM
nRCDsgsdfwA0ecolYsm1dsMGFFk2W5MEwhOhC6dxzUSTJlUtN3fHMqgdrBna//5jB0FKlAEiaPnc
QjNwkzwspYmis00nRGDUVAhVbSakdAnu+B3N/GU7QP1OPU846c32XC+VilX9Q/ddbIyMpe02y4Lz
1ALXPXMGsQu4mm16b3jqSRXO3bp/za0yh3UAUZZQhLORck5Eey0QUaChB5JoAbJu/ARVsHWrhwHE
HemH+PbmBejUW3hbwhxIuB3AFhKVHhER207bwj3fxGCN66BJOGyl2IKDyOeVjBmCEXEQ3M8qiyI/
5xifAhqxFbnrJnpDV7qP3cD27nTJpszANAgckKqlW7V0kmNxrI4wD2DIkqBFrT4qDJvCcDTvH+xG
WIXBT8z9j4v9T7UaPbX2IKGm9XZBKEZd5qmDHwJmSWU3v7Txa6W/BImCNysdUMihrLchSR/qvpAN
kKDBgsYmjLBMoARW+6gT5xTg4O7pAw4pV4C6DMaXyuRTGUfG/m64RXtm5r0kCm99IuYtiUP21l+S
TA4aIQ1M7udtmrbgbaAcTe0XX/NnwfEUDeL50hnH0J/JzJ+esEMSy4Db5FnkxnhrYhSLk649eo21
VLuq8N14Griz9/z4oS3hOfAWUdHvepeXV6a6cnVR8aUcg3DgEZ88pVHush34SclthLcxfMVQCe98
CeFWjMB6LKJu5/TBYiX85kq9ro++4jXaSLq1htzfviCn5cyNrTJxRPxCHrVhT2xQomBQ5Q+FtQkq
njRDduNrnv9C7xFM1Fv3Vhwdgu7U6v9EiCh1mxhVkXZ7Sc1gX3V6m/7/gl8FGmrEqCWP/mjlHNTe
j8MCZTjUfQVknqfLyt2HldMB/RboYIgSAFcOMas0Y3rsiuY/r008M5grCn4mxNA24icbm/jsfPxI
2YqutI+RIXf0UzhlqNtjWc65u8XNSyFErx5s6aQUzpIjFwed2QSmIchYhOSUr+CvJdMvUAwxJuK6
xd9Un5wpdew8Scuy6kOQkSwSF85RzY8tN3mYsTPzkauigdC5Tna9cIUyDQ54LYG+vEx3WeuLXBvo
MowiIh6qVL626HYEexCxXUiUZRZkuzpYjrYiBBzQzBu19awXlo9OtUtrff9VVHhkigpkNjIbgsaC
B8VXLuKXvGaWjb0w/FjOW78EGXP1UmXZc0ZU9B+yFY1k5MHi+GIfWU1dtuqbUMe9CyMy3H56PCfZ
r7+wTVdGWi+d6kkNvKUISfwrVzBjdE2vn2RRxm0Q5eQOkWSB5OCz+33X+FS6YFHhR6umGd9Az1o/
noSgn3PQBZjETI+gMjNlXyPA6MJHXCTU+YQWiMh/4jcpdbBjVTNAcaWBzrPRngOtQTltv/4QlUfW
7Nv2XR6xpTxSqCETTZnhlbrCs9FG4efOEVVZBaazx/+Yq1/rHTFH7O8ll3Ovu9MAk52OSlQ9DdwG
C0vDrSMVVaVR40Hw18j0CnL+AElToWXLIoIzP5WIKDcvLk8+HmMvM761l7DldwH1k2AfCq5rHRor
KcmHJsZbl2blHzv9OClaiy0DxKleflUl9oua7K23AsHp6wVJii/vA1+Bo6dO1I8e5PbgvSGdX7JR
QKKrd+FMPflLxy2dqkQx2xavRpnoK3oXUE/MDAqRuWXfaReSPig8yGOif5K0X8nc96pfF4ygEa52
cAehf2+3JHv5TylXFlLf5EyeRXg1fqd9WC0d7YhRi6C1dgVeT8EMd3I3mLtpNxoiDGbz+M2Q+kaB
7VAaSZqV3fcvJyEogRUWDezyjIjR2pjtJWzrG7w9g7b61Mk+qO0PRT+ZmPFuY1bGVQXfMntzwbxY
ztLZwrZM6x8GsBOK0d3kFCU85aUYjpCh3OnUmc6TNuP0wm0fmEVT+dUUFvWIqAuq3ebsq7FPsFNj
jjAjyL8QwvbssR86RXvyDM4JDERNijEmzN4bzoFX/yNDZtvBNVQyB1RXI42Vh94XU8jLw4fDdsJ2
UghdaUAMLeh8538UU85xNcWvyLinZYCzcLTZIRjIl+mbhplkTFtK1IH97pL8UB3ORNcvwKcQS0l0
RgH9dvC7b/r4TbDdRbWqNimTkcGl51X5zKqQs3LIwbOfTQ43bPCwWpd7bQe0H9QlQ2syh+Ls6m/P
KCdanDkaFVxrsQp3mqQks2O0qfOUI7W2IldVm4M/MsvHR5Hmjw1xprGfLH77E+go1UJrsfccN8W0
phuDsmevQ48bxF6USyMgVaUQseyeWdK+TC6bh8XCIWzWPg69isFXGaBf2fvgUzUFsd72t+Y1wt5t
f0rDHwMRgLbNVlagG38ypEJ2YmAdwkt4FmltypiKf+mHR4te0liZCngvAAbDtIRPO/AYLoHuRAkv
5O8mPTfGLpE7wZ1ngJmtBzeBpfJhsg6zuXDlrNwk7/MN8+gK+Z/QEM1L5gMW67ifhCzgm+La8wWT
ljkDrvRaXXASEfM3WORK0DeCdTIUwQJu5vpw3NbXhRVDL80sm5PgGj6H/7UA72qS20qqMThZmZGy
TzqaPMkoC/rv1ykVj4KGnqaKYIIqSg5YmI7wPNKa8j7efAJJ4JmlAdUNTcx3ob11Hm3qTRggMeL0
qbKy3hvA8fdIy2W62NPOP+SHznF1vmK9yyR1SprPW1rGvKuHzcG51h/2kPkdUM91BXTgp+YfHD6B
wZ6zfaT2/kxav4+CDw41kqp7A5zSDT5gDh5US3IRaScjoQCMq2QjsWrsrMuGqXJQKXVhRRT+qvDt
yZ/DsRPYUwPAkev0g0cxaT+h6g8C3HK7E7mwgqyxu5jaqA1iux2DpxEagv0BjAcqOxTTD0Ui7mY3
zsU9Y5al2Iz4iqz9rnJVoEcV19ZOpGDlcT7W+umMCkBXxgpDpnSSnOa5Gyol6AAqoxHwFvta7Tao
n6IBPwA/h+SYVuFzhtOdxYJcmmiTszbKUbgVcl/w/aq9xqlldg+ZURVMEQXs7DigzNbH4X14F/Az
8xbkqU4Iuzz36AMtDyb3F5HiGUa0nNeBF0UpL4j/yGGSQwFW/Jr4pfMrnVEmlZmMmh74NbqXY3QG
jGoFXjgXMJGP9V3N6qM6cS//Azg9oY8lkQPiZ6cgY2qHKbIDkuZb2bwly5PmYpg1w9kHLEQ2oFBS
BZBVj2eJHqPbdGUimUUxRzeJLjhQtTrfNr3DuYoKdAKB1kCnawbOZn3ipu9ibE45yWEBnGR+Jbhz
wUUpgBHsT3usb+l+AgIdf3qVVEDHn6KNvsvq8FEEErvimlbCcWXUaFTdGbyyOCr+WRycXrdsw61Q
zb9BwxxeO9q0Wh7IlAau7K9v36mXhTTeFgSMvlKBBFKH+wMXUwXee23MQv/pmGqOxKhPTbGmxEiL
yr2bqo03smpv1Jl73v/hASX4GdKy2tT8PMHVJHRDF2pOzYYkcOARqR9+fOoYqPIZG1FmLsa+Rkpr
8UT3NnHVRQa3ARicQ7OWSJTah3CNlusKsfmTOcfnwmG+1TBQ3AW40vTtty3POZBKyT7rWxZTgGgU
9ci71I9Cyb5H/BLPebuRmcI91FqpcUl6+S65STbwRH9CLpyHkIKJOA20KvCB+PGYQsHn5Kk8Vr55
D7viACz8ldhGi6+zQhgbsprP1+SK8aKXroaB1kVWksMBIkMNNpit98objx7KU3wvFT8AG2O2MpdH
WsjM0+9A0Ztx4H5jnK63IIUpgkxgjCuwznHn1d6q8SLJk+b30dQlinhG+8XHlOhcqno7VbeGqw14
z9vTO/wwZSAqeFhDJHfusWWhJDnpKQ9yV4Ul7lEgBHksj6HaO4eludawmaV71mPzbEiCpVvB93Vj
p4l0UuoTaK+bwG5JNqndtsJwrb0y334j7DqrAbhdq8QHap+YVOfYXq/Zzh5TWpEbXs8w6x1WMwaM
cRHn/XIMZXO3B5EHLPVnBt0zL64C2s34r4kKgQZxTvnUcrNmo+JM2NLNuv6+k+poqsusah1kLEp3
O+qP8ze7hrkPYr9g5b9ifN8rQd0/zTOfdSYwoR9rEG8VMxYaUmC5/Cn8OJyPeAobTgqd+9DvBdwq
rMlhpVhGAyWTI+mtxc0b1DNJhWwnncli7wBOEdex9/tTYYlll7MKqUVKZ9fIsQ1hAS2AjaMum5gG
TGsBwoP2SEx6MOYNemMKNW6KovDCgvN38Fw9OYkRQ+oYabrwM+LY+NGnJaBJ2CsnR7LtiX5VHQ4s
19ITK+7G1g4GFxFN/Tyz+m3r7hDqF0DBnqxKljzhD8J+E18LPkfCVItF1Ub3/sxPmgUsV18CAfva
GkbJtFgMsVpRtQrjTn8i5jS+KUZb3QjhvtUXCwUNDe+LPe+xKCNr4Onfq2GCdGO31wwpdCd7BUTs
NKG2400UnoPGK1IOt7f22r/+PZ8rBu3ojpg1ba5vL9r2Dj3D+umCOEZ/eKxAJ2sxO3QP7dqTNTnO
3BCSJ8ksm6yeQdiH8I0bwFDm0ew7gc/dZ8wgiFZreUohX5dR/85p3V0gG6QRvsaK6OflQ5iAzrcL
ZCQSJWj+ExSZTRNA7FYlJjo6cAvHlkfE1WKNVszVhu+Kp5q+j7/lfp0XXwm98AN5BmpZ6MWnpRNL
/1D7JhiFAB5aGOE6N3JtbKUyGegIEu4+ahe3KHNhNvqLAwGzeR27IWT7w1tyu5Bvr9Mjm7PxGRz3
P86wRgcHsUPVbUToDRrR4n7hclvFs6NWGllq/cd2dLnte5YqNLXNsqqRpLwRt3Y7rHlsc17QKrtO
N+JKx+aNTorpbq6QSzDjKBRahacmhFjxlaBuPr0GTL92d9tTp7agjHJ1AnQrfiC7MQHF2sllqWw4
oXuuw0eLu9zVpZGu39pRkAB/Lb1hkMpwJgNvvNmiDtHcjOtdOoomB/LDU9NMTzGbNcm6lZdt10ZV
wd1MYlWTCMxg5fKaf+wbu061gSgcqyVJ5T4y25OAfgMD0uqJnTpOb098q2ZfjAV92QgCcoMECEwp
N0yGPDql05UpX25lmvMqC0sH/9OHe9Oh0/NCm/5zN0z7eNhTyN7mnIR0kBPDCtW+TXZ7zOHJk76a
XH/V3I14YhoaP/vmwzmLH4Ug1dSjJMSESk84yvqwa9NC35Q8BUquXhF14/+EQY/UtHr98LT/f8Ni
F03jDVx/RgVFMfg8WrDhM36Kj2nhPjKyyqdyVZaXHhbXH8DGdekxghZQB4qd3/rzuwQ5Ia1gxnyZ
HMAve4ulwnYCfJcn00TajS0Szj6rUCwDFa+BA4OHMyDP6iuefQTGwL3beQqbf1p5sSC9qNCzswn2
4V6Wsl0F64P8qSWgwfMPWDwIaeOzASkkWbFQaPG3hNxS9kOfJ5HthKj1gYrBdAfWPUTCkcneN43X
kRgVJaoYQHTMgPMdKddaK3Lg8drf8ICgMWAKoQZ3FzP0cHgPhvssgOR87fentpLXTptlsGP+IBoA
QkYeagR2gSAZClUyt6nxr6rMFVMBhddbMWuUGY6+tAZcBAz+8sdQnwK0+qhvip0viWIYbxKETz4C
lrI4HNslwWyf4IUc48oWFiXiDAmflQZnd+rIhiSNnfGsN4ppZgmRT/CO8nOeNK6wBz58NGNgQYTw
0GOwaVRfT09Hi4pcEOEOVdvGMh94gcdJEigBAa2BCTa4BLIm48YMMnO6qF/d9ZxdOsXMXA69WZhz
fSIacDaOBSsZ4IKV3bdsr+upvdyJeqI/u9kdJphU++x3qDw1MA2Ts5uQ3gV9oTaDiUSXXMGIvByb
5D6ujJNloZdmr7dYjHDP5a0ACFwEwt2ADd2fZDV3TBxjs8GhXH1LKriF7tjZSVc2lDUpS8JK/RcX
kzr1/WAy+RMl785vrCuuPGBYjzHLyBH58/oFUPapooMRL7y6D4n97EZ5x+nzfxX9pDmVIDGhFVIe
EnLvBiIZJuPh687ctZIXcVQ3LEpC9GJfJdxFP7KqW+CsHeB9TsmHngyEkMrLr9e7s3lsS8TxWHWM
d03Skuv9VTfDt9Mx7Wf+oKc19D5Z4HPry92gO757wgyxQJVx2MNxuqB2BD6D1B4a9xgfaZpl82SW
QzcvdB/VhmbENSgifLU66GxYUtjdsiwSmWNjQEX4bPHnUZH8gM0XcJlztaLUWfjaLI9DJPe78lq0
K2Bj1skBJ5thh7FqfKMrPH2vTPO5ZiRX9X2DLC0jOhpHt0tcfP/JkbWFbxjnFO3LlFBkioKZtJb8
Sfj1b+0O0OS5gER1eZVKJ8ck+wBDFWAUoNF4lHo2E6rBnffJc9Wht60ADRg/+Ze7aCBnVApPBkKF
gJlP452nUR8Q1t8/dxbep7zKh3r0+l1JVxrYiGz62V4AlJ1E/XKWuQcaO4ValI2QSvmQO0mGf2il
h2XTFAd8uZn2Ncc4KzTH1zQikH71/owfTvCAb9QIifBSqHnvjGuRQQi3syB8B9HnEqzWk103CQiR
T8aRs/HQ3yRR9R/C4mKOrivqDEjvFQ7t5qsoVntDo1DqeMA+XN8G6im9ZGhujBjJPJ8Y6rBhT0F5
Ng5ofYWYiBHTk8uDq30pkgANX0S9Qbhbi1QeDtln4eyYuMuw6s/mgOpT/ariKnEA8OTPTISgKntT
njQB3WFhMTbr+WNLVmWLEacMU+JTpGU3tkq45XIeTnaLapZVnIyRhxXOIsFGWvS+5hkhbEvgaxbE
j6JkQlx72MWIRkwJaKTZRG3aF+38IMZE+kWlkcQOonPwh+xMODIKFwodmg2k0m8ellrxLj8eFTQw
29fQaTanDrs4BtUkYdbyjENGSh2VJqjGWw/JcWm3yzZJ3sUGGyRb05UsmAuSkGONe/v8Rtit2Tzh
5ao/sFe9srwE6aNco4hPtYW2PclNE5q9RfOMvPhggMKyDJLS/1HlPyqTSeAg5CAUEFc0KobL1kjS
oUDfHxYt3o0mYrw3FP4+vj6Ih4B6v8xpfPbOYxSYMBr2YCoUQ/TvtDMpS6L4YK7gwSZbyOBZmX4x
n+7yGR7S0AgX5OdWBON5NBuodm+IqLG9UWS6frz8hXwtLNubQ7PCthIGXzrpWMYVTiBPuhea73vE
5UQkmZVD+ByMfsKxaPvHHtVgDiz0ZXD/+++ZWXpuFloRLYxzOboVSaoMedJhbUtH7UY3VzsPMabq
MtBQO9QeKMWp8rm8trlZXl/gCW4a7nNnTNgpL3u82N8esv4V0snqXdWZ4WF4XuU/MuIKpSiign26
1tGloULQYpwOMOSENKY8WadMg63FQ4lW2kGPCeOghgqPCQy0uW/BBhjYLceht9S6ZAjUIM2nDhp/
u52LY772VZQicmjGPsNBKQmmXP6efZLLBjRDBR8fU4z5bBj/qLyQ0aNseOnz4KAYykaLz/ecRqKv
8xJG/eSna+AtH95h+vO2oYOMFsRPyxf6GreeOvrDABEQAd9yS0li/4qnIBtC5XU8WPT+Zm1P02BV
KBsrsOoItURM24Mka0kCMbCM7s+qg1ZPyQjZ/nKrZIEmdfzsNBuJC6ELtkGbjxh1jXjRCkyOhDx2
3zYru+vv4gfDcDWrXDRg7g5qdaRwuUjlTJIVjRjSk4Y6fvHTKEnRV1PSqcK2L5msVf7YvxQ4EgLM
S3F0xO7X7i/lPWfbiyWG8IUOTWk43yqJAjqMD5xAF603+XKsUaxrbSQCTqJWs4X/8/PordYPaUvO
fyAi+9EAZgMs3KTdGVXEuvWRq2KIITg2ZUanmcmg8tNK5wzBjBFrlTLou7M66CyrXiPD1JH2O7xl
jAEIbu9aBHGGfn3CWQUMEvDTSXwvO0yWEmrOuy1RPsBM6vjeicfd0OWpi53SO4w6ztSXPjWVdQ28
IbFIZgLoDolj5hXe4tJzhUgJsMcRQlGt2I2xtWE3YiYBYuErTGt35yKM3YnQyAq52Il9f84v+J9Q
1nos/+vYAxICK3Y0fOJAkf6fvOFKWaGkygA7fGfyN0OMiWBJQf84900nUIz65cJUb0gtnN7QWw5g
2O+DxMosYohE+Y58ITW0Xqr1tVXcA3eUCqLR0k4hhgWMY5BT0nx4iCuj7H8kJeAf5clQKjjZoeBT
piTnJ4KK9hq1JFFnUmq5/6IRdbqoJ5m0J/Hcu6FvieggePSZTTJkC4go20UtnArsS2r/6iqtANYb
JnyNhOi/Zs8nsFoxeeri38Rswe9Xp/eCW2RdRmbVyR2rgocB0/LPMNy7d3Vcp+m4nK7SvexEVmjH
FvflO8FaA6/mLFBYmeeQYPYLvstEbW5jqJdRk1qvJMq+W+i5CmfuCdUTq2FcvXOgKSLwIfrJvfCx
RyIw20goLGhvY/vBwCsQe0O+sj3ToSc64v+qmE+D/gA2tGFHxU0ItWSxV0GhnPl5sNHfXvj1ZR9J
Voy1Dhfd6l+AKKDBQINPyNZ0TW9aPFrlWnNmNdHsN7mQENY0me6DpEFhJffIEJnSL4CS+dpXcKuz
zcdsrgilcYxaPrNMJilKG9L4tjON3QOfRUoINaBtYCihENvl+/r8zGLmZpiJv9lCYBXKr686hb6L
MTVS2ygeaAiqwBgBDi7GlqD67DMiC2lcvrn3Yuy1lKKsQwgx0+cTCQhWwgtZk9dMp23fHPz6kNw5
uq0GkHgPOF/nfmh6WFscWoXn8/huhK/S6PP1uT3dfy+IOrKtBY+YtO6xPrVzDSxTCkyMV1G3w+PF
UOMKh1dbCqbEJOrmitr2CJG3V+VUWZ6IqL4Zrzz4Y8HfBBZJ1JB+HFjljG0S4vBDfYtuQ3+B+h0l
ZMS2zODUlBRrw4+o3IS8oAn5zNFr5OGKyC+UJWQd5VHgM4giFspYUEPV+ZvmIqIfy/VyNZ6UC9LR
ahG4rKHadirAUzkknoF0ossjAbD8fS6dSKH9L5gSPz07JU9DQv6URbvrEN/KPAponLAudWLPNmTr
G48kaxbLaohbGA0h0EfRx8JggX1k/sHrFa14sL0VBYpKw1Di5E+oumZNoJaD88uFwtn7zMRrV9aI
F7LvuiwJjbTy2BRuc7DS9YO2MPyyl4zXq1m5WV88wHh0qicYvreBytvtPhe5NLdW6xSYXMf8PEXu
spqvvIwvAzNiZbzNDtHwJz4YAErHNNxxcVAPeXsCZuCsidLih78jNrzZ20Ay8apBiVXqT2QonDgt
t88Vc4RxhXreV1gwvyTqstSkh6aXbKi+ASiSR1cb+FNUpkG/3KDg63oP5CWUq3HebNjoUkK4x3AY
hL5mca0gWCVZ8nMT6e4W/dvo+9TPdF41UugfZCrPXgaOxDrF5r1LE/niNdzhljW3dJh3ccRJyBDr
LERpqBLe3VNMKnRTYER6Z+4Hr6W2huSq96eQ3sQHoDug9snXs/aN5O4yPNII2v/tDqWozVsA11dc
W8k/tEENjfSXPr2Ag0rzJ1zjPSHLdIAtpjVn6YjrvSXU+Tks8hpO4PbTLU5bPcBg5rrvf0HN8yU6
TuKlGGIA2zZJcSuZkB4Vuj4h/MIZwIEG98tWJ0aEnT4ldSgWA1VKYXbTQKudDbVTn5n2zbbB3zvB
QotjPxp2dRVH64ESQvPbkmSzrc1DgkErmqVkBsqE267HeXSA+9o7PZ+5SIWCloh5w2I3WnOqLTPf
L0ENtmLjh2NRI7sb97F0zOhTktczJTVHmfg9ARi4/Em6t2JREcZNK0SC/yiZYyAkdtkTX/3pQZRJ
sAiy9QcCvpS2DlfvnPCo3c5dCbbyx9+OMY2sZ+/Ijc5fmtAa4AxoVZ9n+o+NAmMmVKl/MJeW4uNq
q54IroO9V9/ZRPo1et3SnpDwzLuMBrBTilB3WgLu+BiRXk8z2Lwh6HfhBKUOhcey0h8EO+YAi2rR
9Te41k1kYOXMq0HumWmZWLGtdXE6e8rLA+ZyjJobZdUIrf4lTieRjzSjBlhVLkMnvP+iKWm4xKPV
o+fjzKQtwyrOpi033FtkCDbrIa4BBlL+P7chtjNsloDbIQu2xnmvYv6AxGMIY4lKDA3ljHCVf+AK
vsVchaTKyQU0Qxg4X0MOE174aYWdUbBxRlmSYgUTpLOFM26GB/Wf+z7mPlWbC+BhZP0JuRNJ0iv5
QFKa9LoVZtXVdKfqb6lawiBDi+3R1CX+b4GMgDiXKmo5UOgslm1WBWr+Rvnf6iBq4rHAdHpfi+C4
ANGbxRv0q/8tLz+ZMD+wi7vUQr6jkhXNMlXUXuEAg10ZW3QUJ12oKWw4BqDtfMDIiGzhBwzcN8QA
ccMZ9DkppggBs9NwyO8MTfD4zQT/YyuCjrMiqU/XO9wP8929ADkMCoAK9iPURJ2QARos2zuHz+e2
4JDgFZEIlRkNOcFL1vw8iuNPwniaiXZF1Eppdm2Gop91cJ3oD81hN5rtqqjifcBawEDxYijmvn0T
U15H8uwH9D+JytaISbW7Mk6xA70F2B1NDZ5mdHFNGrTN7U18TKyYUrpqfDfwqBTxta/FASrVHntY
8U+tATMeDKrWqSFJPCIiXARSEX7gvoO1xT/AqlU7DqIeBrfQKl5le+m+8AdXOBoBhWr7RB/GhLab
pMas3Rr/YNrjE6vx9HG4IQtkz3F5/2aDgpkYTtNUPkKtsO2bji2JANZ4E3XW/OyeUKSD+OJEvjkV
cRmn+nQkmqQyDdJ0NFgGeAmkmvjlqWCMlbsJLKHrFCPkzvhAJ6mJevX1xjlvwwaWcfMw3I/uaIOz
+y/ZHPRtMMZsA/dOIxpuoAPr+qsqtpXpFpOHOZW8a1uVDAYMyvUm4CpZxdP+7AX7UHnsagC03CMK
1tAeFw9Ip6ZTbSWnRkyhJjIxb9s45gxn28YhjRtgW9vmU1P1rPvasl/PkmsLrd6uSVTIFTzzPbHA
sS0pE55rn1qebbbojRT5PuCnE2xSfe1/VHdVwaHjONqC+2leC2+iJJn8iGw1W/NqQUJ76Nuu8QMQ
NwKIPyBKqzCK+qLtU2eiPOlQngF/qYMonIMwXCK5T7CpelN62QMHSk85/O4xMHsZXWtwZQMjxGEv
2GTCEJhjqxQ9jpgCs0NNrKGdlsa6ZH2eO/gkufBoY5mv8wusiVKo0yJjnpLsqWTo82UzUfckPcLT
CVY0raUSS9MEkqcKzxvl7zHzWmwmFuFiMQxFCEyYCI+gl6e9c1830U/GNLZgY3gTmyg0y8LCmK+2
Dx/uHo5AMTMSzhq2To3u3meqhqfMhMzlYHmBa77qHJMmWBlXsYWZlh0lm3c4iV3kpw6FReZY24ab
2qgamUBiV4J0X5wlN2XeprdmaLrJkvraT9Osq+c/e+r8ktcAhzmOwL3KRc7fX3lkoZcbpjPvSq/B
0QrLyJWSwzCZNOr8fd7Fx/A3JK0JfZZzztKKGKaE6jDL0vtu9JU8tYz6ydIcArQjoHBlBrPDq7I+
h3RA92cEviZXhnmwa4jNu4Xxk2PIoxZB2BmsTKMlvzyK69DQK3kmUmfSvlS1HPFQfbVxBgEO6q/9
L00cCg/p0n97TYrLDJQDcYzQSZu6Ll84rk0jzWmycupRBfRfwRqxlM/z1Cq9cfMPXzbyIFKNN9v5
xttg/sbLLO4uETkcbN7NLRZALOD2fzZiOfhTxP61C+8EBk/AmuT2NlcAVwkR6BZ+vcQI4p39q4ZI
nYjSsk7C3k/p6InxWiyidhnDHXqlAtPdQrfARNGd2JxtT+AHfNQGFi424SDSFfga5jbC8P81fjDm
mgdbiBVIvRmrfwuyrRf8Z1zQVNXdxb3tKv2b6URKPbaz9iP4P6ILcTNNLeiYz5hEdH14oFdvug5B
LFkkdp4excmv4yWDOGOAGtPdqMw/UZLwfMN3V4uPxuE+d8AkHIPZdgq4il6Trhp8vPmwhGg3K3VS
oLOEYeEQj01vc04bzVdwHEh5VlMq4ao4URucaYiryGZEBJQmHn3XICkRjiO1hW8/fo6/au+1XaSZ
39sTK0x4qlMM8HZCqp4viqmvl/TUhFTtJuFrrOZQtw6dchd2nZV8nhryc8NnXiVl8ltBwT/07B6h
Y9y0nEs/cmYyuIAHWmN6hJZ67Th+dISpcWxuXXrLqVk9tAs7kVyXwgDoTJxOjzDpu2awGNtFH8ho
7cR5HYV+gv0KFT0AEkDujHJcwUUVmktgpOamEduk0+RPRhibXIaogLNaiRUhuRUNZX6pwPXI9Xu/
JDVMPWB8A7XLLWDkv6xV9bsFdF0reo/P5d21f48ZhlJZizKN72tCQJyXHctpMCoJCWMryhJLTSNq
wtr5ZFapJ6FGo3mWGsExG0x3GaL90y4sP4sEelpmNIReImEw9qr8kXbrRlorOV2UzvWVAQd2+Ato
JMNO4nggesukQom5QB7Kz6RlYDLh9b+Ruh/Ab8gHMjXkUlOfxNPDxnpP/zdSIrdj2q/3M3LnWCxO
Lo7TJiY9bxPKeypktSlDVImNaanvxX+jFEloDC57NRplax8FmB5qpYWCxCkyJm6RhZAMojU5bxEq
RxhqSpAFR4mqy2XOVEpQ9+ztUZSxrTafV1Abe3GrJkqPOj/+zbJ9W7t0hWon0Faqbgq6QIAkin+i
fD8EWHz+nbXTwsgYcuraQVg5CGsqu0EOj9W+GUVXCdVyu0eht3/c/xqyiuIHvqI7wCxYmkZyPDV8
9EMgEV272GPTJi8oHoccJ74hSeS63ZF3eZYPlxtWR+GXN2JEDWEE2PwhMaWub7yWtZAa/SSWcgbP
97dKaPP/zaJskreOZuwUVMVFLHwMbV+HbVzSZVkQfov5d7OX5Jt6wZ28fZLyulMrIyv6Eb0712oC
vL38tagLHmoKj7UaEBn6k+e+5LrndGDKJzI4zah7o+YlpH5DUVjl1omnTK/5Aglv1oyZsLLMrukE
rtt5gP71q968raYXUiePu09OLVbKrPsxePNiL20qPXPcGwGGcH3xHlMIzqomTebILnmbY6m80w+b
dbgQzZBNA3GK5b8tWkg/8Nqdxmv2TVsPFm7Ht0ftUpNBikyaRPzLITGIkcREOUHUZJDVA/eH05sw
JdyR1UUrAFV+0ipbEcCBl8Y25Qtl/ntDic/3Av4XUXi7gJtxY9leMb6NdEZPqzIy/2rqsBETDMyj
25rewmTA44XedL3kHHkip1FXTc9uAoVyhlygSEBN5Hx8Gt2eIsrocK7+nAVvEU5bpWvI6lTfyYdx
/deDoMChtju240mTmnRySm8F4hHrPqBVUbmqcqmiVhgdIaArS1xDzKUNWDojjrTdMnjIoC+OEuGM
hWnALvV67ppHTxFHZB1o9OwKW55tYtEVH7eiN/fehP2sdq16dURSRpxhYMYYsThKAcvZ5tOVKsZ4
uLhdKSysAqXZwIOvVIhZpPv5lwsyTayUDX8u8J8JqWAMbJL/fGLoNH302VOxdClRxY8KNYvd02Xn
P7RWASQ0ysM7sL/SJAKFv3JYBxuSrJdmtnR3vGw08Z48feinN8TnhuWLvgUsIV5mTfLfcMxc6Ls6
WA0HfWIksh7GUERHL5ld6t5Cv1Qkzd9v5xHYyizg2HPU6YXtQJaz7HrlCUHwlmShnzSTUtNgyrA1
LSTAhZBiP83H+a2drBm9jtzkNYwatHQg6Ec9sqtufVz2InP8eWIeJbN1obqJ57jouXMV0OKW+dtB
XqPyp8/B/7E6hIphsZPL5d9e/cygk00U4izA15yP6FLLy7mR+2DP42lSbEyGbnFpwUHIHfIGR76/
O5rADHcZhy5bFIEMc+5LKQWUb4N9j8kBh4YPA3ZboAuDoEs5tE5SSQG0+3d8j4OGkXXRZ9MJT1CO
nwLw3gZGVl1HWRqRreJD6/qr4kCc57aULclGTR7SomO6/JYpDzYwvgZGpVxGHnjdrTGcWfcGIwLL
3CiOzCE67F1yTkgovUkSNeXe7qhOolA+TcLCn7hpV4HRzl9KUV5p9zBf+81J6nr4F46cxPvF2/LY
KVRhg7X0jmrnzR1WxP4Fxv3OWRwL8hCreOVMOPz2NoPmLYAKs6Gzqi+OOdwpOILlT0ysw4VD6yXB
6k0dXtIcEIoAJxu+3yLxXsv9fYXVDnEkGQJ9vxftsGfcdbeUm9b16ewdDz0NDY3aBEmb5/zTKI29
fe4Qwtd5NkF8cD+Hbo8nEh23ItFRG4IQg7iA3TL8CDA+ooWm4P1JiLeUUyUPlXTP6+DBOQEna31N
Ur22P5DL0Et1lXY026F2hf1rgOMgIT7wuSXIBC/GDI95rmLEiv0c5dpScIct6P+DZ7jQk2yBTnqp
mOOQgD/uZkcPOXbimbNK3+tT25bXivx8ShvYvEv+7eoMO9IBGFfocjl9WA533pBsPk0pH1apLvRA
+CWcqk1mI6idrIh7803+6/yZkCwY9CoWsyor59BmVoIyiE4kokMpV9WRL65mnd7DBXZ0hyLeJNjP
MBCTODT41gmnVTnH0eQQEPASy80VNkfujM3CAtxwI42mvMH6NvhuHUxCO1Ty3v68/8GR9vrx4SHl
9eie1UKZmLFxi+NqJ3A15PWYL8SGraZBMLlDxtDY1c6VqWuBdXNPvMC/L/ONecjJbHs8CcqFcmCg
DHv2PhQATHb24Ze9meYF+v7WOaNq2QSXUDGSaX9cOUUxU9/umEqmevdClgRxnOwx8BJvS0/mWDse
guWT47A3hbb+Qciht6p7tUHctkb/rgOE4iqnPbHnFcpgU8NR89r4wRIwXN0HH+X9B4ulzn+8syXD
YHmANkWjArjuXJflvuaTq/J4iPvvACtMTKSgqSggmO5Fn8g51Mlr65SaD6/cQM9RgKM3JgBOh5vE
9liGFi/hATCy0tn3B+8eBogFdg0tyEukoAlzYCa1VLTVcxaXc4G1hjgfolscnTGAesoZg+cn4rLD
CO+U1CeHq0VAxy8Yca4fI3bANHVlyacozJT5WtypIIzKtV56oK3P61nykH7yqk1l6+nKR5FNEsXG
1lR58o41t1XhgVVKffQYSJKmJNlGU4G8+6itT7RgNPTpLHtcwvC1PyxUK3m1x5FWys1/n1riJS+L
gkDWSL8igtyo3lzxIbR/XolVDmZAIcPvaUz5ZttS99Y49QpS5BisgJZm1ziFMDGWw7qQbpcyvB+T
3FPptFSGlO9PHovUTWvYEzsY0H03Omc0qDpwoq7kBCVqbli8BTV8ilrSP+g4+2dBzUOiAgNgIeob
ofiN3HyOOqWWHsrwFyPJt0L7DEwcMoIkYQG7K/wSD0edU1Hiw9LSZFHXDOTdWtU4bzCuUJNC76ZB
zzFp2cNwkSk4P2Lg0XPmzJIQxOeZWEHQpAyid2ybRL8bhfwDPJN53IFzVvVwKPYsUfjTwYceqyaI
7nAF4oLAGT9tjz7mePH0AC+XBMYkg8B8Z4phGY7xF2p2jE5bs86M/R1QxcuKBL6lYeard5xO27zs
cijPEPIHPPKbJOIeWMQGF7xJ5DBi5OOj6q0uVInxfZ2nZAG9hPZTeUBCDHo3Gqgwc2JfsEgs557e
pXnAAt+/lelWzEL+f3WHVBijAVab5Rq34itz4a9bQ+1IvJhahEysD1+2ZWkBBNUrAbdgqznvr2QU
FjY/h4lm9/Goir2e7KlfOXJFaSBFhRTvkb8R5BdqjYj+kpbESFwQJZ6Hj4zJk7xVVJ6Ek/bkq976
E+eLs9aOnRaARcqJitJniFp5z4UD8CjdH97hc6/u3ZFUU5AHyUSBdK/0GHztUv1DNjsTaspIUYGj
Ja1QfmStCT4fdA8xFbUiBW280jdIybsBB/h1ryc2kFLjH5tROHXoHuppsbAVWpS2zn2mI0sVLjj9
NCjaWiptIa+2ZMRl9fKPC0WfiTs7vhatxqc0TuHGmCS79SkXTe4bRd8ouTtV4uR/yXhmYf0QEPeX
4JzK/DJXrTOkAG7rfQHGaB3z95QzKiCP0dTXThI/PSODa9gJcSbw1dR9LrbBWzwStHrKJfWHLu+Y
aKc8IcSaiOK6j+PMNGAZLT7jBGQO5K1DaiwRj9u6sTxT0kK1K7GM2DOI/tEsBOJAVf/CZtv64ZpU
/13rlptS3CaV1aNiZAS9rDcACKf4m5f5lqcOnlus9M0eSDpVO38eCvWgyIOQbuNoH86mkIPyzNq5
beRWfxQYgI0rXuinrNKVf4WQFXFFD8EbXl9xZ2hvxtbsbvKSiYAl7MCzg0zp9a9PlmsMErzueFSi
YDKmAfQEjTMH99uM3jRE4s7Clghr2iAKUY6sYIsNg5KPyAHzYofiGITocXK2pysIJGUwbdi0CHAp
kHw2KT0Xfp7L9OgMFr6/ivLIIM1ChKA+tjKVvMd5w5pMQkhnXa07DD5US3IhQzcScF2ms4gMwNlv
17QJvBktVugdtRuTHEN6nVboqov9h2hDY+DdnNvKKLPKHGRK1/gJOlydf1CvEYFIj/zgnGUkpCpZ
FL0hjRHemBLV+21fEMBDtLa5+C1MlqJuE6aDXc6l0NULp8wLeUa+qERPNlY5RZQbOfa21ajmp1VP
McvRVYyZDOpmbbztyU9WeObdo1DicRAnRuUyfeeUNG1OLzqYMyNOHlWUP1vIfHAiUjuzC0VxxmXR
6ZONR69sFq0MNvkWohbcpKYiril8NRNhx7x30mig5bXUIV48PB6fjpJlW0vWV3ougJCBu8me1ot9
Qxj4dIAaGbu846TtGwKAHLB6gyPM5cMjA6psicyqWliUPDsFmChHWMf53cKFDNMIELkJVCwxVd7s
dpSVbi4TNL0gA9hGqcNcZJo438KpwNdB5yuea9jf39m+2QTksZIshmMrTSSA236QtwtpLw0PfPYC
8aVsCn/Dd3JsbEY/I9s7/6vmbTFlBXZMPP0eiuC7t9V1MlhAynHRlz3toqrvan71nCJZZNbW0+5v
fhhRdlmpkbue4pdBjpW/hWGQvnQxA1uMcDwlRWqSsSOmwivbvZVmQIJsLjbtUbTJnQNGigAkPn2Z
bIBPtC4o3Dhw3XEodu7FksVH7z36Hf8lmcs9VqLEkPTshhLd62QccYYeie8RiE721SLTKTqORV3k
r7excqrCVdu5PiATDyocFnNmFn9E8r+PfA7bTSWhtD0z3toiejg72y1mEUj0AFDavwdvkPp3mChD
IsQ1N/s9FXiR+J5o/hJiH6+ZEa+xM0McNuug3cwrW84q4tP7aXt+Qu9NelMg5TmwIEOzsyHDjfmv
PCitHe3A4cBVgoWgUyXuPskWWmKzdJW9ORhi28w154aaPzd8/RN0YWhB777CdsMKRqMJYhKGt8Hj
16l9Q2zC4pkJj/EFLVuLsVbkyyG876gRcL4yjX7lqjorXJvxmrtzCGDbawWRzdaRnX03/KejhuEk
YbzOtL1HZdUdjaaLUjajQtOl8gmToALq+rrOYttIva3NlxuAl5AeLFB6SfOzr8kxCRj5n738T12G
lsbUnxN0uhQI27Xjs78P3quethCPmCQkqq0Hf7XvXFlRwWra5CRq5KYY2Srezg9i8qozZJ4ax9mX
pMXN5qNdChdFo+PrRQ8+g6cMGDRc792fyS3Qm6aajd+F144fZsPaQZXYvhOdOm3wrpx6D8uf1Q3J
+ubM9o689lJum6l9XQsREUJkmu0Bx/S4rxOXJYotpBLlk5ECV1tsljTD01rFgbU1quocb90H1qFL
gcWPx0O/DpLn6uV1pVh//G985Id8AKY6lzjK+m6nU1FCeBIlMHCSjROL+T1DvwTrrxTGqJQo3Pq0
3K7kXRd4+ucGb2b4bfru7x6WkywxZfsV8lwtj4D3+HDJV49oFM5NLC0Dzx9tGfjEHm+LCMLzofPi
suQihnR3zbzLMQzzD1eF+AkDUl+HS+HjuYVtutyLIoFkkLXFu1Vg/rtSh3+yfHdqkFmzFvOYvDSO
QRdlmVkc7GM9kbZwcQtlwrvyIB1PK37iP04xt8l+0R9zRyB/hK5uT8TM+mM99wXgMJGjpgpaIRfc
6FyHQLQ0p8khm8X9oShexdkTK6FkOaRFUOM3C/b84j8R6uw8iSbMkkMXsx5CDfcqH9O5shkvprlT
QzzB9rsRrqt9SkQgSVtYDSotcHmYv7V2YSXRgtGENjxQuwoGEIgGvnWH1V9Xmw16Y9UBD7xXECf3
HSCF0MKAwaQNFyhofOBJTHG+/GWHwtvkqwrmAWtvnWuFY8M77cJcSB99Dr/SX/XSWR6mNo+M8/W5
3PKv50UuEjusz2Z6MwzJ12nUlwjF1u6ugePWMrXC9Odmr00+qCL1IzPOfdefjTrdFk6/dv64KYQy
kmHHR6oI5VA0el46cM+g1dnM4UVmFCwPWL5Bk8Pq3XuoiyQhrDCJi8rD0OdjnpnQCqXPC50p/rJD
sp8Os8QP0LZnCYz3MzJ2T0g8a3unUBuA7CHREOVGatiQNDOS44ag+3AKDcTKmrZ7ZXN2sPvCiOqD
NH7D0MyBFi6Fpv91Jxe87LKc6mI2cUPBRaGhNykEPQPyYsVcDSGBqvjI5oQ853WiUMfcTtDJkvYy
ER1c6YRNWI00YyNEB3wDDanfDc5Jpu4Uszfi/453U3R+idW5LAwi0oLWMyWYSGP6TDkbd3ISrWxR
1zZ8x6CUxQe4q0kx3p3iJQDCto2H8Q+wRl6VIm/BDnkazb2zYw4nVrhqEBalr6tRhsWqnfMeoBvx
oVmC0jmmbzp+S2LRSoZKkW1BbJWDbDhHK28X3lrdABSSXExQCzQ8z3G8MtrvXwxuC/AqHfM32aQA
58v8GV/NOEct2p3MA36nnU+jfRXYVxebPYYE9F/IZc8TvOonNlySrWxG/LU7DgppkrtIPNCfTNBB
MK83IIgGA0y0SN8JEZARdWx3V90x2bgOW1jFtqI+rOdSlgoJLB7D7I7/g4BNI/vhiHoEcRaAsf//
B0zpzxX5YLqvwY+ukM656R01QJROsfSpsE6309wE8TJR1M5HmlojqE2j+eow6LqNMd+EwPpcbZS8
bstZaJvuqNY3qFUmBKOsabvA4J92sx449YyFjXDusk49vewmkNIlbtso9CWJa6SOqfgtR/bCBFoK
scNkvJ9hOdT2ScrPUmypeca5oHhwRClkM+CsporYIVBeK9ikUPAEAvfysNdeMYouItgXMHjZEj2f
Lx4G6SYZg7x4FgsEE0KGy1LlVa3FgeZhjD9r3Fg2f5gd14b38oPnt+jX688bspNtOGr0PsUD0L9I
I7f5rvtYlVhm0EXFNH9/fU7/PyJeUFpOibePYgqz7HxgQAwf4e3XLl73gUAv1qgDyOwAEyHolf+1
4oPTCg8jDvhNTzdNFr7lxes749cTeyfBEBTJ3SE8PKWC3xDWtQj4+5V+htNSmRtlAYyPt9i9kULV
6ddZBy7rDaLzhqppSODOzJcr0aOfE58AG7jgglUdq6vPlySgaBhvjUuZG4/mb0J6csQaNBZw4eId
Y15mtwK1SNVAs7kKfyQUqn5knerCbZMsic4iSH+lRrRtq00IhyKLSKV6cEgofPVvO1IQq1zmB8N9
5+hiQKWxYLWamw33jHeDUnKlppz7z6Qn9VkxaZtAua4jGbYcn2aSbRmL/JyKwinGn1Z1pjLYFxXJ
SzjdjypoDMJ8Z1vG4A63QSxwn4CwIuFzHQjiTLhhL9C4pJfsKG11OGJPFyUjYK1o2PgxkUcwNO4V
U6TjK+NLilEFU6wH1kVFJJtIHxa9SA1g4iFIjniefIEhs4M3Q6yZMxSCDhB+gt+75Rrt3pdfxvkz
p1+V+JpNPLMkaZFbYtuJiXJA8OJJj1+FACPY/VyntbAFuOl5qtJnzLrNSn15ZaxzIXTzNWn0utu2
hs2IOQjXMwQM9o4N2wDJJCn9Fl0L9RH85FxIwHrUzexfH29g936MsA+An/wj+vmvvy4hOD2hzSe+
BHW/eSZIlJdMudKY4L3Ce/tm+NxAm8yqbsojOJv96r6uD4UVHVhrrzgImSXx0IWlhsqXGv1XuVUE
sKCIUGALcLy9dQpKQHwrT6dd9FBri2kVU0TlOMoRcOYqx9QO0BAefutahVS/ACVUulWA/0vlO2xg
lYdVNvNwur8MYdfi17apv9FU76aCkCx63sOUeYtbFnbnuAX2LrTemEV7Udanj9m0/i/xraBxIq8A
YcToKxh+GVaDCbMN+X4m7IB2xx4csfXf5DlIv+Z4efwaQQNzNsQ3bEUgK6LUDM21x5JrvNPpu6XD
BwJGFyG44bQGxNRA32U0OAspsVUryZ7tW9QsiuzZlN9YHNjCKSy+SHq4deEdVkxFXJNK0hgscm2V
7MOxWUbwT0XSRHvxe2jp20/auwLyWdbOdMfRmoToSEA6XYUWTJc+ob0mS4132vm1WWVUSQeQsdQi
Qv0VIRfMDDx7beID0x/rlo3mcp55u0qPl2TBOgcvJAQmpYpQb2KPaMu/OFq83T0uMyj5hAFcTtoQ
HBLrLrmVLk81xbUBBMrLmqtqKMXbUJQnxRHdNvtiClCzbyTcmEz+tIjauY7g8rC3ouBNdYpI24Mh
7TkJhUf38DTDG4koXFzXskb09ZTrDhwhuJfrM8vFo2/5tduRzdgmtasTjlswyO3LzfljEQQBSCN/
4iS2WaSyQFOWIUhGY7pc5vrxXLfEtQg9rd6oRhuqBksjM9yx43Q+b1gsSEcjceMYBzJs92gpNFHI
C3YJ3w/PUFBH2RhJJnxYpfs4M2Nc3V1+pGX43aI+QYnzUdh8TNBEQR9HcJVgsGjuV4Dhs7R+Up2C
vuATqJkfTAsVvYaZMThVwAKRD0HWjcwCptri/4Ytu6NMAZpoAK5b+/VGaCSb+cEnRE/Uk52uEi6X
8Z7/Co3nMt3gmh7/Ng/X4goRJuhAcNsDIUAEwU+mqxZza2mn8pswnosACBVQitkBfeg9hdU6HST0
yOGhw1rZ9HuVd+zp8PApiySS8XiUkwIaQYUofWSQWnGCwQ/AW+ADTjJctGWcooCDREhrHis1X5gl
s3TYly8iAxblRcvkSETJrKAjwuKzMIGgAEAbxO55r2GUGyJkl7L6WghPuILB9s6BjEvOaacBE7ai
SU+3Xa8YCdd4cqJwaOLWG62fzVZ+kHFcO9WTvaPRQYbLbL7hH+Hnl50zGCCYikcBYmylbilKsTiV
WCuxIuXk53NZkdcu8cW6bslkCDoy8IPVogvMqKYATitU4vy4wbgOdyljHZ4oJc53jJ8VXyobP3tb
AsBJ43p78WRzA1ATe6CCXIpBovj3ss/OXFfIwDW6sofT5p2P50ydbb5xWIK3tFK8BHdblfZFsyhw
CwQbY5fkOCTDuarHw3YbTR6cBhkjBwSLxAgJiZDV7CTTq6q5oK3naNYp5WQeTAD2TZvBk1Fe4oZr
zEgUh15gpts9rCyYsgLsItNGB9adcQoRkpErGe6bryL+DFnnkcDVGanWWuJRtqldl5JJGxiAmRFn
AsXJ8NPx/q1Spf3RA/SWjKSg3nrQoOOh772HHpHPqCb1LZvogxMSI1grNeQ7OmR2aS81Elz3/MiZ
73a+kk3gfwTLXfmP5dPMKpTmDja2HA10/ICTYQ7kyrPcSOGrowSLgdjylOELVpQvv7nJ1OkbVdLV
QrriwPWk7N5BqkN46ZtkX4srbJeF63wl/9CbkXizhx/S4kmnB1L23kw09aOfhIAv4x5I89jVETln
kz2ke2/MmXaTTviKV5t0KZYvugPXf41Q2Th74syDT+RlfyOR2fpKHbpB9Ge9EC2g6jZVor3SIrwL
Jj1qTL47vSyqyWB+D9vKtJiNFiIkqVn/MGJaW7+KATb8uWGr3wNN2FQlKhNqHxryKmRDggXxPjF7
drJWCVmTDZ6nqNNpMpF6ZG+hCDMbAEx5a7XQ+KjjHYaTOeQ6Cj+k6LvoEv5/7AC6swE8hOa7ZyFD
hPbuGa/AwXohs1NPRAIDwsznuvXcJHcyt8C7t7Kd9EBjXu5Oyo3ZLwuwAXJ8xqcPZ96vVhgdNKM+
OYbohzTg/P5fucx1FgMhPoOkFVKMfhEF/yLJjph0B3qKVjA26fhH0doaDtCTN4YiZJbV+tdff9fG
9Vu+LtYF0yFVYG/N4zcjjHb35iyP51amtg/y2nzaGfy0+J+vslBb4Zjf42uQOL6+P48ESKOzrosO
jZTzQ1N2aHVwPLY03hx72bavlZIGQyGsdrWolGi9TsYLsnwrvqawbvdEce5o/g62N6G5CRknT7y1
Kg85ysFA+GWMEKnscWn2C++kOVg2r+ZXyhI7Y05HQwx9ZyjSEGPObdRYsKDNl8NtMC8ESqBT0+6m
z0wRv2iKv88jUn8Z+xxAWnbaOYCjnPkzIZkx/w8Epn299Ut+gSwXJy8l1c/7/12EV0Q+FVr2UhQD
RSkxr8oKU3hg3vSNt9JeY7f2OOwxU8EEuWZ+epIJRoxaW7wln5/Zk0rC/K85HWV+IyuzEBjOPSzO
DveOcydFxzfzV83U4p+hH0cDYNn1xTkCrSXE5IexnjeqR9gmixNy9XOS0IEQIFLjYakXmIrbzWCk
c9BpUdIYQsz1JW7YVFunq0p+BDpmCA8liPIigyDqBdcAs0w9zTxfOwt+ct551YagObEhaYHtqb8Q
rScBzsfguoNAZIqw8aUk+mh/ZpB5bSVZQKWPSo0QiPth95M9RuQ7JFH+eCc6wWv+i9Rw/b4mbjYX
DlmunME2TlICA87BPRbAsm8zDgiscJMP2oLcwMzK1283K2shqH2+fNz/jc1oQM1K4SYSzZkuiLyL
RhYaHXRLGxq131HsJu4NjcmbYfL+1q+wZAUc5aEDxnKFQ3DZeGVEYeNCqS7uQgmyNwCWXh2C7lfD
4E4Lg1tskX3u3WTaV+/7IYjcSpqvw59VLP+QspVSGY0Uk9hs9lcIm1LJXryJg8y3i9t97npYqYUf
oeWEbp/ArDzllgtIq/IhMgn90d66ld0XLDhLs9o+0UpPIz2a293cmOpkZ1LmC0GDbrD+9NslEFvp
P9TyYEP4iwhfL47hpUR8imNuTFGygSGbA+jDiC2g1lfd4IEUQMkKXr5sx4V24tLF9gkI7u+ZrWs2
keSRNXlvXNpbSpMJpZZrDtkjH+TXkoauyEHdU8kGpqvx8rITmRyRpZbA7UYEdNO7PDlEso2obGhm
Pq47OkjhzPsxfAUHPj2bjI6gekxTX+GpNA1jX4VVyr4jlBKQz1glgz7lqx4CgTr2iVisQAoffPhv
HbBd0sZyaSm4mI+VlK95Oo6wfHwVhBHzvmerz3WoZEd0SVs0lqwg3PezFhXWUp0NtRfZLF64s11m
TdpdpfY8EEmzhMWen1rON/XnjL++0Q59LykMYbczH/cFt7mUpZ/wscdZsY08Qa6SdbumwUEIu8VD
XDKXvrVD7VFbqpn+3bgAWK+yb15b4wTTa6rMyKrJ3uLP6jxWPMDahJsbZBc9h/Y3BaXXRB1k+us7
QQK9Pr0BEMd/43opNQ+UsEWAFSsADmhpEX7oRAGO2cfhZbo6P+TEDr0iDwA6bRB0DxGjbQnDZ+TT
W1/qW1G+QdKdbB1RePQY89w4Kbi9yBq2iazZZdqyt22tF9keJhrX7K5m2+8k/CjaiyN5LymWp9hr
OvBlOHS7ScCFq+RBtBNzx2rzq8dloi75bZOfUNA7deccUUs9mF7RY8Q25ot5O8uo7PiwHFUH/inc
2uONOy09RjNFanZvUcyrobd7pssCojt4FEc0j5vjwANO9QKGP0nAXqfr1yWLBf+9kyaA3WA2Xnzu
soQn89Yj2To9EWT1WYy3CoCGyG6zTs1KPO3DOqR2mFom6PPLeTl31m6dPjtKv39s0b6Gxhe4+Trg
2soSVa8LPvumFPl0zRWHaPyPfCp+QUqjdQJixEoChKzy/aUqoJMlhokFVNlbLmcDpluzD8LkAfnw
SDkKZwGEQFAbg7YTdH0WdWN4PjeDEh7uEMSXM6D+tp6/OXH1J63xNHWKaxQqXMsvtHmrw5hXSZ0r
iJieYtqxgZ5752pmkc8zGlB09mR8nSYmnFh1nd/mZgESoGi315++Oe2BZRPK89iBpviIahLpz9m5
f5tFAKRR+lj5TMN9YQngRmtC2ogu0cPSeuWMdz8hP5r5Nb4WN1pMD3G8PaqtsDZ18Tdcj2iznlEp
hiva+CexuXUv8/BWGrb/xcLxSe4KL2hMBAN1TtHzKL1YzvsymCucVnicYaMagMDfwO2mHY4Ve8+y
UzOWvcK/58r7rv68D/uYCHPVixKb2soz2gxxUBeD6Vuy0lg5pgmtfx2g6rtE4k+/uKyhgsKmYdhQ
vzVDeNzWabkCmVPFHjs0nvXBoz7TiQtIwKBLvqduSeCrbqQH6R/qBNwHyeyf++pgo4AvIaQwYNLD
XCmFqUG+ExVfMdXc7Op3SiYuvgUFRokSkqreFF2KmcfJFJrf+oVSMzJDeSVNnjS6QMRcRQ7jOuxB
xRnLBKMIAPRJY9c6YtpGpQsSqBTukEBeTo3kq2c6Q9JShvvpXeEa1rmqeZdsfhc2POwsYdNDvPdj
+38htR9MaZ7WVbLVBM8arl61+EvLMITzAIF1G5rXqe9vt738YrlO9+aXjidqgHoUxcLs1nfE26nD
88fECMlGMGI3sRLur35byQdIkqbRxP2BUSZDsR1z2FCEV2Me84AyRMCOsNzev+6tiwklcgb0B5Jz
A04oru092GtPSFTZUDibPFk7WrP5mfV4C4FLA2s3H0Dv8tQsdVRjuihL9MNnk8wwYF5iyTdhmlmO
ZoalZoLSXypCEufjLwlm8MOVmmGqLTQKNZz+QdgFp67fx0zyjRoKsx2jJW/EXfUMzTTxdhZX3FXj
VjVDoQ2VQBaIEaI/Sz5v37DR3Nv9u/7LrZ/LABmeIV1a1ENsebjp/ArV/LBLHbFsAomHofhDs1yJ
QPG+FuRujHMwMZFOQL5jMbtowBPVoFMzBxhsB8OI23/vzHOIhGe/uj94E06vPXwKBHPT4wjUhDIi
eohW61NEmLHmA11H87aBmvq1/t1jfp7oCeNZ19LZe9KpDDbua0eNq6ix+ThkNIzsbbIXAddzXfdW
3ck4jZZzI0t+EEJYCnvwIfPmx4cdYPPSjk0IWyhTGtR6QylMSWhrPzxUmfg3BEGMcpxWZyErwv57
3n3WYFOzhVendA2wbnOjYH6HB3I4+xLtOW2yZqR0ram5ef3Rf3WuWTInPdYxKENQOW9GQ27iaee1
viiBsR8+f5UxHvN3pW3fNgcGGzGD8jn08gDl4+bG3cDuKZTujBI66UQ7NL//inxBKGa6RC+czSGV
dabd4gUbtBhZbOeMe4GQ1heHFtxvj46tDBtmQ+w4YVWZYwoGOlyGG+zCqh0Ji7Ppk/1kNiv1tF23
gdGXq6vitLejgnC/PtRc1gk+ggFZSxHogtLyKS1lK1wrl/Ngz72KzR2Poh/kctZKc0Wuu7p0Vn5z
N0UwM92F9f3yvG7kn49LtyQbLPeEHt1u9S6O33ZJPOOCnMWtcUQCu9J/Zkkzkap6foSa0NqAbfce
CzP2IjRnw0/dTQp1FM6Bbt0gQvAYexM1SUOeW2gJtx/rjJP9IeN/aQYfFlLmB4p7uNwM/2ho8l8K
7XjI9ObmyPMY3oBt2cO/UKEuSA7R4TSb0THKMoFJU1D56YfLR3KxNMnVzM1DlnxJR2IqocwnE8B0
KtomDIA2b8iTEw5uqQzYgZ4ZAJy1f54faVJetzf81ta63pqlgzlpNL7Dv7JFF1j3hDahwUsNNEmK
aYiVVz1BX5ow6qN6gEsb8FKruRmVgya7ZEvzhkhHsAij9vgHMVdHZ/DPHqbt21gNts9f6phx5jdO
42wActunRc7ODD1tgLffAc4XXRxaBEwgVK02Vxof2JveCPjs8RvVEweqG0CcZTOBf85vXuXZIPKc
ne/eFlgim4AoQ44hG9Te2yvqh0y+4/UTClFxVfdT6TLqdu5DbB/EwOHJXYuVEZd8LSMOFCbzjNH3
6wgNGMdJDMz9Yg+JUOCaGTO2008zJjOcj4aqxGN7qnTC8EN+DD4y/nyXZhi5kxJFjI6qGfGhqd9c
0qTDoy9VETcbu8tUlFw635Z8ktDP7Mf0Q4b6G6Q++9pYKpfXj/+S2SK8dubiR27mZjaSySklWdiB
MBt6CtLXa4phO1/0WuKvETsOsWQeQBZkl0GGEXIQnGbjneE152GY6fY7LD4Bnrh8SrEO+OCQEGnO
uAWFWk27f4EItOizfwKdMSq3peMK2dWuVIKbiEsgF6vfgqZkYf+dQJ6oVOsUUyLqF0syt3PcDol1
QeM4I3W+iZB/eFErscuYXYcXbUrWUpF4lRhTngBS6GkuYOlr3AjJIOZefoIHF1XZnC1ahFmPUQn0
v/eAG0Au1lSARws6+VB01YnYHfeF3u6rVZKQAVR9C1NAbu2kep0Wn2C9gMoIn9sScTkDviwEGTiM
rsOO3a3buhinqXS5OPz+JgU76+t48Eg+i8cH/p2HUvXQDJn3fn3AwKaxGmnXYlXcRdVmhcsPmpsf
uqFbCGySoxTRbW90KYH6Y/FJw222cEVbOJwfpuReu+6f+RDjG/Koe8aUQjipWvBF3qxNsPBZB8AX
8sVEpPR753lV7yAZFk5R6Fev3Xmhrc+aPC7gQnlm7wj/9ikemiv92QPPR2ogNoXTvcvVnTjpmgxv
KD2hNoyWnycdy36bRbT9aNnJ9T/LfXCxR+MIHYnJH2LF/LRlroTiNVIH3VgF6z2iDzeAZmnDtt7f
2OG0uT+zIVNNo/5r2X2DmHFXY1l1qcaWMgelXujz3ZigkBPGcjk1ob3+WJXmkJ1GkVAuF+rHXCzt
ENebrZk74aG0bx+/+JvX68bS6VgN1oZjue4YuIEuMr82Gh4CpYCOBxfY5N6k3LTFi3GVZfuZSyGF
UvhibgPok/AvMwM9NMnfYQdYssz8WEUP2nb2rKAgmFcnlbxz8Ob98p1tb7dp6NZQjqMx3c6BjX/x
+tcr6PsSx06kitZ8IgMWJ4CbbV4aa0pQVUlZ7E/TEFJ2vaVl2XU5FidYPMNsJ1vc71bqDclGy5dT
YyfO8TGSPhiyGSiZFs9xbkk6DCE3evsb5vw4+COggN90bE/P0dupmZbEw/zvK3lTRFYADdgkUnVi
TjIMtwTP32DBqwRr4tpqwGdIn7Q1gRZmdvhSaGJHGT3B4bcXvLVnNac20PT6FD5gf5xpKJOV7EW1
ld0NOHkI9ooNWqzwXFuTkFMeUWwNG9BWyCkBGME/IMI/j9mAzMfj0EC3+rlb8ZwiscgCS++z4jJQ
wQWXjJ6av5QlRrz/rPmCNn5+5cxsNQjeJukr37I5DbyXz3e9hX/GxGaLQ3JmmUe5Y+P6vTaNwhii
HvM1L4NOdTUc1ol1CdaV7L4JBzN48fkLhBH9DBrAmXAZzNRNoZ+4WKoxe1d75PybJqs5TBCl13jS
hBZxGCvlduM8g56IAR1TK0D9aR/Xd5uRNdhgqWtwRuuMftNuaSy5XIPG1aCt7P+CRJm0eVyqbt4s
I2rvI40OWFBaSOPKLgF+FNC5zjG8EpdvAq4guT1ZuHS6v62V2E9wB16OlosHI3PuZhDN0Xloy/Nr
8FgG3kV9tDCZKfpk2TrNn9as64I0U8hBztO4Q+KvEIA5tLD5rChWBq4qLBayBJp1g5ENy14LXWmq
LWaPn3zW+mVkXaP1Fq6mfMQvY8H2jAnpu6X/cA51tj3dQNQqU8kU+jCvipO4MX4eoKIcWJsPnbJX
qJ4eZhNhVNVGdR2LxUYnDN+asNppEXDnCQSA45zSeVA7ZhADGCBXE6nGhcOiCFocz19+qwz2UUZ7
DsH19JTSRNxY4p6HEiS5aUdO6Fp5Pt0ghMV3OYJiG3Z16CJ7dMMQpbdILH0ViUQj8FHZtiLdKJgI
G35pfeYryr8x4C6yJ4TsLcOAq8oUDS5RUNdKP+T55mwiC7uVCxsKZ1iW11MTvOggESsiZOXgdAgg
FPbrpbamx/OI6z7Qn1UzpP8TXL0SN0bhJ/5crk6JC18maPfqyaA87g7YkUsUmyGf4dYlVaAc1JTL
skp57Y5r5XGptiFuZ8LjRoIF62xn9I+dpG87OjKcjNBvkhnSOPIK6y7Kwpu2VZ6DqYZND7yGEz8c
JLnuVf6aXBqHifLZbDC+PJOqc2+l+8WJIMsJGra2+c8OU3hpAxIGjJWKqfTYxfVFbttvWe1cVdvW
hXmq0RVoPGWnLrS7qM4nG/Iz7A/6S/Cwbj6H9gvTbiLiQuLmb/TkYnDPf4zwVuC5CD2qRnILfuni
p6v48YqBYAlFXBi7NfYe/Qt/DkeCAoyXD6FD+SnnZ9JyPrOHDNIuS6C9NCD8/Qy9swsQYhp8Rg6p
tVHLhTrHbUPbOFPijI9mlOCX3gXdPRSJh+FCx4NaNyLF6RNV3sdeZGmdPh6lpy3qx1X5PFRVsO8a
Wfrkw8OvcRpMQprJ97tTzhSHNaO4uLI/yK8LuHEarXiJofmZ84nSuVoxgW0WfDZOSc0HMPMiwofN
M69jCUP83RSWvEJABr+1Fu5agqfXCpBO7o1s6emyUlMXex2q+rxnvkrQYzo3ybz+DbwgsxP1PGMt
loKcZGHcE+92TBq8+G20vt9p/livcDByDbXVYTxyfo8DlSyrIYPSPNYumnH80++P6maSM1rBlbS/
kOqHaPx1+yf3HjmkPuhgJnVjtu/SHttvWmWffBM5+woK3KoQGq+qX0DcNPc++IgS2DXooDeERoen
k79hX0uCkFZjpftloalbaaG6uevwaoBizRKcmhC2AlCb+QLAZEhBH57w2hgJmrEJOauqYy3QNnxz
W2WYCa/rERSD3kwYzXIhNWx+dIyaDPK3wCYMnBwdNFFPAl/5Uc6Y9WHWGSUTGVFXfMZzMSMV/LcQ
oNUNurpY3DF7K7UBjDVNofTJUr2EIBaGOeebwnxH360eUnKJgWIThP2vxyTg2ooC8y2aq0uYz676
avz/p1Zl5/uT5SR44ZW8of06KUP4vQfR8dmVZCO80diuxBQvJbqfYNRZikqWRuS5ycWRK9hl3U5t
DTKT2K66JUc3e5JMPhvBUCLOssvKaFqWV/r/+CcNzA732CLV0uljUhO25xPes81f7Ax1PwXzPr9U
fH1pYJ0bRnxNqKKlcvnkeAZ1ylPkbtd5XvKUekpc1D8UJnkpsV9vwUPeMAGA+UXrkpudB9OledtT
sjUP20ADBzywMb/pWW+zxnPCMME5bYfEhuIerYb2qcgpJX3PVxS/i5K37hChY0TW+WbEZvX46f/w
8xtZa9KAFfHnBIcMW5tsjI4HeNroaJMnV/hqBd/Ih6rbp6A3s9CmbKxWl/mUK4Lxz19hkHmkHK56
AmDXRQdj1xyszRsxoijmcxFdsc7kwapx9YE9G4UvsMdo6FV4VYdxvadbK82ukcCtvtbSlUFrXCMV
FlKKuScMpRCwy5vTReSS6POXqM2E3Q7Ag0+P7fhWiuOESXaWN7S/Is389qtjc4h8zxxjhHLnC9QA
0cKeg9yO5uRocFl5BvD46Rj+Pcd2cxzbLUU/lVxtpUKY/UdAIoooWwWzimmv0f53/+DfxBC9h9z8
1mHG7OB+v+/DvXfWWFji/+b2P7l5SM1Fl6uNPzaTLhlVSfk1dyhPOZQ6+g+DtWqVMlGW2zdRapE6
zFHoPW8VtHHSYvfc57etQyzvZe2tBkij/wnoe+KxYLgciO6//NKR2ZYvCJreYr9TLNa2G7DiXriO
DIGQ8V1IGYoJnjtC/gXLFyTt2e+lucZloxJCqZJ0xIEzjY7vrPIZNu3H22SqVXy4chVpIX9Cs+Zw
jqsCC7lbmzz1Bfp8Py86IgXXSO3JTk9bpv+YVhe0jiCWaBR6yxNF6u7cTL6yxv81NEFC3dVVmAmR
oZ6JkGTksLhqIyVjHtklpQR4QDFLTrOLcFDqHrsANjkm9sNpNdZc0G65synCAHm8Cy+tflP/nlKB
7owiepsSJsmZ/VjdXhpoNH8XqwyWEYn5xjeSdnGXeIPtpH2RSh8TsksXyHuKi7V9OX61w5uH1Bha
cxDXa1VDLBrUj8gt7+wPXNotRdSuNh1YWY7m+Lllu6unbQV0w+PmueZbc67hMxJBo1hUQmgaljEs
TQU+FLsSUI8VwR69PjravylnGzEmErrGOfG84lEZGbsCywTKI6BkF8NKCkejGYomuqLuTOIpt/sb
1AaSqrAYDuXn9hliifJ1yWHd4c+aTALPfvD9IjNARNbMTaUeTFr4DRarJv1Rdp9GLVYVgwDLb2Wj
BEl0PycGCVL/Dsc85nJcPM7FPWVo+cPl0H6Pd8i76vNaV8oTjl5PPASQEzX5mfUkayV0YfcPs7GE
Z4PbaVRlLJBa//V3XeYwwIUZk2TUWwU7mPO4+rG7qAWQPUnh05PETkyk7bbxYJxEQs6qoQhRbjJd
uSGSaoA/BM6miZqcfOhxeGXsqpdlSf4nvyX1eN9moophsxeMc18Mxm996jpaGfTkT5TmfsooDJrI
FrQCW3qRfquCQ4viQttmeXxISbopRQYcXADb8H7A1a44AWGDKgxV1ED1LmyZxJhkX5E/Lnl+65r3
FRQ99wUysE8rfTUxPjbYM+44lPn/7PLbfGfGr67tH2c8Zr+cGj20NKm5LOoqr8naitQUcqHHh83k
1mA9+233V4N4gGjuVwy52EGupVTLGryotoo92jdnf7Pxytvm5nhUZwMORthEQAgbrQ72/dU0oBmJ
TbPXpoe42WOlTVrMnlVpP8JbPQibv320gdr6Ws64oZlAhvM4TCz49MfEHz1KeWod36EcyfSLpqix
pixK5De/LT3SfUqh3Q6RvbhDEI9L4A5I8CHfyqVioor4xElsLDTFBRgsAsj31wTqT1jknYJdtf21
PEKLD9NnjnRmzfcVI0zNiU0KL+a0eEmPz8OIFGsLpOzQCXHHUYMYdCNz1kOnz/gBEizUXLthxejS
Fcfvr+3Fk4VailWL8Y11kWlup17v+gfOyKIJnspO8ZBI6pbKQXEPKu0K9Puc722Lwa3rkE/k8jQA
5XDuhfUlhikK1xOHhoJKxURT4TwS8XtbcaQtA55uLO5Gy0t8lWSWVSFSw0YbsUl7HhKB0NTFZSRE
zx1sw+yQs/J2K0dusg/oxuoSLDSjY/WmFmIgUdIITrAwzzQdfLOBEONNX21WzLIfsRA+u5WtnQli
qewjxk23aHkcTVqWSUL3T44cN1+vQ4xmlgYG6nLaN6sb34lPB4nr/oeky50J765oSWZA1N1+xTdH
O7lOAtzIw0NX06HiPE0cXynwrC1P+oPm9yvfwWEhepY5GKSDB7a5uqGHDvE7S2Nge/+EsHMxvjFT
Tbs9vW4aFjw23tigSz+tke0qlUydLVI5pOWbDgKK1NtkUACMMV7LxaIsacZd7OSd5MOM3Ec4Ujl9
J1/RMHJSvJ+vLiqoXpuQYJqLoIb4uUwHiVAx5nrau/3lVNntRwudig80rE4ntQOIz7UO0ivq6Ujr
gOyS4OHHBDi94FD9iXCFIJQP2sr/lQvAV6GDL7lS0cHUaDDn6+L/7fqC4NIiduV7dGEx5mBsom/h
ymBbopsuIp1ZBjaDHpYYSxWc3T2WYRxEbfUgbDtEtva0LLKYvpqYYT37gybp/hIctgg6aLqNY2Yh
G/+BzKgTvozvRqiPeOqCtE4yZe+cNs8Wry+PHxb8e/pFG5g/AwZFynkjGl3cRRSqpnPpdKXpY9GR
rIaPNbfqinDWWkudypY1dOqeEmpBJOBQfnONYzprFo9fkGc9+x4b3QppYy3TgJxxEX0l3zW6OYSe
Vn2IpGqKdwKAE0sMsEZLevCnINLZxxpqLiPoizoRgDTf26n4DNzbFP5n4pEjFMtH/yJJekqCbmNu
ER7q9n54+rAbB4dP14fedyzlHYltNSY4ZiA9H+yfSieNEZCNA5/2BBjifdHi9cpgmG21DNaXEiW8
arCZ+tTOBVuuFrb5nm1La43zRe28fkAcerOTa+ZhypT0OYEoM74n9g7vfIVNci0CzgYInYUmY0fD
TuUvvNfxHCC77BVtEXWxQW5vpeg2za4L7lHqZAQTLTgp7YHMPbdv2814YXdkvInjwxDVHseL/VQ8
C+527J6MZdxjRgw4IWbKqi3c+aYw16AFVyjtExHnEUHSn2ZGP1Oomt7lluPlTY1oOfb8YuRVS/wF
DPQAizK550e1DXu4maPrOFRk3Z5jS/wcOk0ZuJ8hVI9dGu7Cgh08uqiTWa8CSJhJ2PE3e6y3bVv1
+oR4BxkkfUE4zTzIkSC/GLPl+3b0dqP+kWMiC/mnoRplUJbrofsgrbOI4bdkq/0D525ZAt88tQLU
X/ySxRdbXjLzZoT03huN6CNCQHWMyH6pK5+PnLOEH4oB1LYhbM4QCvRdiV/8AlMVhVkun8v2C3ia
ldzbprTuPzs9v18+5kS/fZUy+2uHB1ziNay6o7lpC5I9LJo5hvA92qsyfwLRbsH7Yhr93owNGCQF
GpbDUMfFPg8XRg75BTyURdjJFujm8KlkOtKm1tVtA9UxDeGbyeXJBsG7jOaEFsw1VLUVURMpBbwS
vd2czAthIpVEjOhA+Uf53+MUxpHGY44ibc4UeMJ1QfhSBDWlVcvz3kJ8+bhfzzlc1MJBlWTBxW+V
0srV2wmrWX5ODWTn5XhbdTL2ulG/UGx9T3XQoIf7zXVebp81MrnGd/ryAN4hx8kVv4HPf+B7Cqja
8uWiKf8hlDq/ZEnZvy0E7QpYzwkYoQtfHL1U9/aLnPCvjM3qsEEd2gTfSjNw+5k7pkzQv6mDrgJy
L3rUJGOzmHWjMkSgKj4vOiJL6Dvgl6dXjJx9VA8e/esqptW8ucUVrq6ML/t7/E7clCUeDF8Idwxv
uloaEblqqemIdA1lMyYaJt7ayVOA3uCQ/R3vS4B5VLDOt6SO10wDO/IWEj95KqBOXrDF20bsN2qk
lsXSZqQsa81wME7FwTphhCkaDoEx/IvLHkpiyDmxNUsRuE2jOW5aqj2/dQ8uw17lKsKKgZxYcdZB
JPwRyttnbHCAUlFOpjvu7MWgbPATS9LWw5P3Qt2IaCtPOS/0nnvDO/aowzitndbpg/t0+5f/y1rV
It9VGhX8g9sy0aNJIZHOaOhQY8wluQ4HyN7qWeiB9bykfRgCrEEBb5lX5XMXu8vWxPW+a/Y/m9iu
Oi+r34SX7r0Agfl8I4RnePqJxka8Rdli+tUiR1+7pz+BgPXc1FvWuwlquyAfJjwGL5l+OQ1Vk/Mj
hT/H8LTsnQcP9YIYJaNWND1Kdr9HU/SER3a/3JAih5y2thTkFh5Lyr6bHaYB+fKqklgsIvBvBA6B
DCAM3q+SQ6QfSbtPhbv91Q796L0XJgVL+NXD28yPG/F/k+djyxg4ARgwpWK6EqRR7pNULFPXCxPG
T9HeOHcEEwdA3nxlQw5U/pzjJ9/ESP3vXSGLWHm0ZJXlyHfhzwv8SdJGJVyuKpaPwwTnlvBVOBqW
6D31RzltKEtY4RQaUaZqR8kmKjN0TQLw0yVzezyDA12/qcZaVGdGA6/ZF5e4MceiMG+diI7UTEwT
Fni731aAAQ6bnvru0esO84jdGbotz2qrQHfbaNbv2En2m2kIMcVvYQrWvcgb6ic00qmJAdNehQId
A0UCZBqYzIVqQPnPqwtn1uRAv95gF6gDfOhfXQDdfE1PTvgyZQKp3Z5JlQYKlkraAhr092vLFT3V
83OhV6Vg4et7g9mLYUIs1XS6WEYOdl8plIxgGyu/tP9xSI9qbpvOu+QHDDr/1bCvGKwfVSM5D3Pm
6m0vEeAvpx04xp6UeODChU/r39fCcj3F6BKjwtXgbRucFyCMhb2/ClrzPSq4OyuDBEyLYjXN+Cst
+t+/dsjqN/VlWco5ZGrySOXMYx0miZX+zO0oLxX9Qzz1ieTwZjESx3f+5i2uJ6L/y/sh/6q2Afh8
yt3otHUAeoJnrFs0wnJm6edGAigp1X0X2Z1F66Zlc9JXq2KmApwAb6PQHVohiJKw9scaWacnq3oW
EtdBb3mGAUXfhoZsIcOk9BNO0Wy8ACfY6MTQx5gQqdS8uDGVjCmmhMGsdyAKhLioHdJy0qWwi3tD
WFlDYIXm9W4f+PTtRTdUg000IloruVEkLTNocrfen1kjUHljYroIgN1SXvvHnuI34Anz/UdOIALy
srh29ZcYz10wYQvjlzSbs3+r5LchMtnkimES5fA+fEI2RMTyVaJwaNeFTzlMkVBbVX077HEZBTD6
uNEZSdDYib4WuE2OH5LhPoZOR5bVVpRlrtzRQPhP+Rs3Gybp7FezmRW/Mh1eSRDOhHXt0bWtDTyK
YgagRrZkoPlEelHfYGa4LfVOsvrHJpe/t+rOx/yqeOxrFfezoao4PvpEgSxyah7cZvqoiNmSCNDa
R4uTlkYFr3JmBKEllgAhXyQHOeBa4d5iyd2c1A/SO1f3+bNBmTa3Y3tMCFacZ0qBA7UN1pkwI5oV
+6b/TAB50ZhNFN59lxRB1WYEYghRQ5OyUN/5TclAQ0QmQrho66ua+GawNrIPMc6d4yMEzW4PHArd
2Tw0mXR75t33RiXCD/aeF4p2txMLcv076xrgtdaZmmhNYuQmcgkWpQXYvypBLWUxf6yZSceJRSh9
dnz+2Yv5w9YykcIdzT95NZFx9+xSx2pt5AfqU8PXwbif6eeVRlTRwfv+YXE3Yj6eQg//bc95a4qP
ooHCpoFMiBv/86s6KqM5qRO+xtAWVLenFBMcABc8ckdwoRT1Bxpo4PnHvUClPLzBZVpmfthFfWDp
CZP1A7NSHEwq/VX+r+H/fu+j/aA9szGU9+mb2WeFmAxs6Sgl5jmLTnwQFgf3HwT2avbzIXvlPFyX
Kde7PEa91rOM9YR9HPETMjjuifsYHAj7kVYZ+JUg8CAvzhNwn7imlTj0s0mLExIoOZBGiwTAR01D
uZ9z6QMu9e4wtlhgQdED/VI2/Rb/Qc6lTQfb+z1tZp6TiDMDCXPrVi3So4dCbNeBAQS1mFVG0pRt
184qbmOm0+CubeY+qSSMu6xrnyxn7dSILOom1qBMo7LU8U/hioXkAegmDv5H8Syiky8yzFlE1JWL
d9HLBoQyhnSopN/0APGwqj+sHPfmnkT+6SR2ooHoo1J8BOB07F5oA2aAP7FaJ3SO+jNd0YW0te1b
vXXEaqPmFAPfexSJRd6wFBVP0oXpmPEom+sw9jHbncXRjcl7dTOkXQ8lOhuaKQHWsps/TaZWi6Fz
VD5SHivMbENzE30rcc8LQMLuaSK9npKrq2c+Ou7v4gxVi461aGS9UdWw3ccfmZXhRQwCrFuCGMfj
cFeKPwt4j2Sxx+CzD6vKbKFINlt4XeEuKxUcbARaMzy1mHGYEcyqujCxXMuYjSWTc72zXqH6uvJr
feo/Yo2Nx6XGLfMp5jY24tl0gThnDKSnstK0LE7a4e8ZV8oQr9+Kc209a8GC7Gn2k08E0L68F2pY
gsS72n2vRLakakLGper5HxTtlMYWgM0KIxVLCH5aD+eAFl1Dz7IwRF9jFuX3AlvFJUAdAGspBnn3
JFKfJBSqQIjwlTibSmB6paIqyPA6taqEwyQ/qki6SB/oyXqYCTsduzDkIOE/AxMX5tVuSHfwfzE4
1cXRTrA0BkOwKkRIdy96RTFo0O7ZJE7dgvLNubkD9V4kpC4Z9zpORC5uywci46ww1Z1jQoZq32yF
JNY5FMq7a9cSGfAhsDCEvHTVv9QvDfz24NTQVdmIP49J7icdBkI6wJfvpf6TiADd/cptv9QWx0La
FFX+587RuGZR3mi+1N7TFzSMRTwiHiMN9P4K0a2bg7P9o5QCjE9FM/CDZ/v3E40DW842e698lD5+
UzvYbrhHPBnzjZDU8HR4APzJ+yY/crMlm2TsDZS6n+lzl1GXQ2mPrOHO1lZ4pU0ZGwCjsrZUBH/7
wbp92mqToRquDlJTs1NRurptxdbZpPBFY6b1Z1hyZ52dc1Dn67XLqvY+OyvcvtvGjkuiCHF8XcwC
uwmDuw9Tfgg00LGwgppC9AsKfXTZ1Ov7J3ivOAoMVZnkeJYkGRb6bCRMF+t5hZb7G8gDdlbd2X6M
68TKl1Ew8OBX3JLcgtZPqaefngKu2n+YVhtgMmXNgVkeSvhjHosBpg13qgudAhRTz3f9/Zw2BMcs
awc3ZeWL1SGUUAkQrcSMka1W55iYCfRadigEJThIGJDEIdjY74AigEb5LIPxzTrPp1zDImfBhSxW
EwpMNvyLzVS4FVHXTw92hG5I53jBZUsET5+Ff36apjBX7ewggutIU2q2VOA+6JkJ/JyiXf+I3unW
Q5YFPThLgPw09h+5nkOJ6mKC0hzIZEo3VX2Y6cqegNAbwDOkNzHCCjtSrEMt6hteqnUervtWeDv/
fSj12eO6RqMAcq9LjYMKzXxrVuoj1MGW1U1FdEXLN3OjpOyhqQ0qChi/rjTcOYIFhptxVHiOm+sQ
43hcAKlnfHA3+cVJv+0n9rU6Ei10pHEk/m5qu1+ZYXpRWWqY3OHkZSfQURVNnEatDoDdcIL06AWa
1+fzvna2E8htJTLAw9HDXC95U2/yZhDBl2K1j9meuy3JSMSWkU+BeHhIyi/o6C38iVzaHsSgYTWz
BxJAye73lgQYt1nu+w2SDeelgOyk0oEuNmM0xXFKjqIxTiHuP13hxhnYk+vesE9hKP4zJ8buW+JL
l7y03VO5ms5p4GyRDpqqFcLXgycYosYSMhSIdBq4N5CUSbSUh4tTkyn2Nu2nOm+zvwgyky8zYbhC
lIjNdmOB0cT7VeURykeDmnTZ+0DngFcfG5JnEODn9tl+yGDNf57vbsxC6g6ZBYXET5vS2d6k+ZZl
BSMiOkvZo2QVTDoJ5MRPq9XRhSKYlWtdg4BFHeQqlGnpDDjagbnirAEHUgprw6y8/DPYKHWasaaE
MAjiUUp2qXOlujZxjERb/xd+pf35L2JUVXyLOCjcq9wsyih8Em6Jv1BLYBdHAaSp5DVy1kuR79oT
/NnnSHF/yeAqXExJ3CkPTaEU5VR6xKN0fLbAFqHjChvb8RhLs4chBHi4HxPojSKIEYaaLw/ViyS7
vFqSYcioDE//BV1nMdLMTG0dxuXe6fUzHq9c1eyjEo/8g5gVXida7w+eS9Je7TikLQN4uYLsTkYa
yBY+H/ZksSw9gOnB3qk61MvWhWMGM+0HnC9/NocyuKEKxhbaovZjO9u5RLTXPjkDiNeHDUF6X7aS
4raismi/bY1RyawOJcTRGNq8quim9TbOinM3kcBFX1E51559hs98SHct9B9zB5dpZzHC13oZD3pb
0JgpZ4X8xDL8/1nTN7iQ5HKo286XJXaKXWzwJYr87q4vPR3Bw9CBH/wddpwErlnscQf0attK5/dl
A9ePWroFTQ2g28BryHLy0K1lZwFGbwsOdkM/8I5QNgSIkA4itHw+oH1ElMOGMp2qFpeuvsg+R96R
sLbY8o1d1EPko55VxtfXUyE+xllrRCAe16nrtXaE+bfPFuahkdLqs57/8sEMjTTJ65ROdFTXgMjE
9FnmTQ7MzzolKqWp6qpqNEAutXdWMM52AqIe/abznWahH7wjcmGmDPB1z16tygevhp34cimS5Zy7
NYes2ce4iICQV+r+DG0aXceQoNdaPhp1GDgob9OjOIaD3ylSGNWgck44YdJ1U/vl8gzDIS5whhiF
0a9r+lovZX56byzNyQyJ5O8JixA5ozO44RGVj3ryDKXMDs1Cz8K61wV8GHVHQdWZ/JrnUHzcwxOV
OqjUu1V3+0l96Z0Q/wL//uAD2QniTXPBq/cNBMjOCgHbm5gnSIP2pxmMV9/KBt+xW+e/Mn3955XB
NUrQII6BIFWU7S8d6qlf7Ngydum99qCV9DPkwqSuIp6za9GcKpQmgAHGiqHVsaZeuMiUaRO1G6Ug
IUR0BeS4EPZIr2jg4mpEkRXOFwRN/PdN0IhU+dPacFtgn8yaCV9O5dwBcV4Fyf7WkubGKZU4vaRA
neyP0nDDgdsefBc5zM0yx7mi2dEPgn9SqxfU/yWEYyyUhhoLIA6YKv8E5jwIYQCR3u1V2BAZof7M
2D75qGJx/NwEkN15FidXH1FRF36eJVp8xLeQId6Pk1god6Z2ywOtamcrq8E/ak0+1uW1ae5bnih4
24V7D7mJRTNZb24F8wwqlcSZOCLvzJRBGuTESB8a1T968GtOjR/itwkpbI4zYLPEjC0pLbzccLk3
CCzBieoUPktEmN+hljKICYZJ9KfpYv9VMpr57UagfwuPFpBv3HtVICKLJ2KrxFBmlB3K3TIdSJ+G
aJmh2JtQCMyk59ADBYkEyvJ+YXAzjM8USrh+CrGfQkPHgsmvw+3ammDRR9dEs3gwpPmysfIUolqk
x3RAsV7bJC6uw4Ei6QucH9OcCrPmVQ+/kf7YdqLMkAU4ILyGFCO+LqNQjdeL5SW4zWuXMsRo7GVn
mR4UDIqOzPup5sUDdNuzx3mtY8/vHAZMequ79aEcZkBynwAtgFQusGwIZRSoZ1p/0Voxv8tEbZcX
uZiuoy1ZiPpJgvmufTyetoPLwEaZdyjBTjQgIw9x421N0EPPTvuA2Qyjl7q1mp5s3FjMebSt5Rsq
aURhBGf9XPTDM0iDTynKGmchgXb1aJe6vXnqckfLkdImsCFxPJydvA4GSaSO7SsSpLx/X+OXV9l0
reKBwRyurLpkLnGRcpQ63chvZTVqxBjiQxp3rfdc0DAZkebWx8mcjUeFSAptwThdaLxcLDxoGx5O
F+PEGOTGUmsIRCkLrV50BQj/Ha/mKfYl0i0+tHkvz5eD3TAuvWJ9BTq/iRx1/46chV8xEwKSY2ho
oywU7rBMp10lHjbZ3vwJ2YGn8uvSrIpxBmdcLCGb4SVuP6CkyYeQK1N0AF9Sw70Esiv87ZEFhf0B
i58Oqmy52LpDA1kYvCF0MK+7WVABk2hs11Eg7wbv0CUVg0DSnwj2/B2jCaIHEnKXjOGNWj6eR8yL
vQn66I1kKuae7AWaya3wUL6LJOLBgDZ3A+i7f01uDDeoDlu0rLFFI7RnpXhgIgB5SE44x6MQOgUc
h/QgYJarCkg6tfVrws0rZydnWof09HGck2cxwqh+iFtoQYD1W6x6TMFaiQUcng70W4rrWQ0ALAPC
CV3BdnhB12OMSNH7sZNaThy+KasX0sepNIL7t9Nj5Wjn+Bsnf9Z+ID8gqGOixkrfXQVwUw92U+69
gljDM+h46CJ+mKGVEjT5clbARfe+tTNXn36w6chvuVb5kCD1eMYM3i2LQn5AxYtd2/N2OU8dC+op
rKLX7w0W87PCaTnudQSyGQ2dzagT8mlh4wpkvgxavhJ5hcYRMRmhQ3PTM7mpRfAbMn8Pq6KFare4
ibdiL4GZ6XLgJDMqYSRdmL0EgQMYl0uPcSisoz1hmupJhkfeMDnayXvtV0h3jl9SJvxOFwyOkgBy
CxuyxI2PrgVzjkXZn3mUqbltga5s5INIelQkUfLkszW4MZIznj9DJB+zx+E4mkwM+V7t3QE0ObBD
jYYAAME37/gG+geuTCbdbx2B9wjAVFLQIQ46EVs6DVNJTXGXo05++yRt0CiOXRMRzxL3Z/Eve/I4
W8yoMAOqBeVTpkjbebp9eWSDIXxrxMj/TtrsytR8xPIJ0wk7VsS4Bdm25M1OzyKdWYy0gt4LPmRi
7kPnwT23t8sWfX7TC8Dhlqd2y7xr7wJ/z4yEbO2YFfq+AEF6vqy9xypPHqeumpsfQB9D6SWT/R17
k1qepI7umVO18YIw475EQwW3dJQ6PkIKjv0dg7QvwlDr09xLf11JgbbvowPL6XYvPHBiWz8fyexW
Lr+x2lVT5BlTDjIEXyHpV5dDYKUUSSYujjU9KXrqqM7q44ADKTM3HfDvOoFjO4baVptp/0nB/cSy
1/1WCSXiuSFY5aoaY9QZeOhjvQNO1JmsNU9nFsH52H6cO/++m8wiaLKKuFiqtmRQIksWIKWOs5hl
uGEOa7dseNBWM7wBvMI7GS989QK7sPe3vQwx5nSO0aDli2ZyxCvu0mHurjJ0cbreppt+pRtRBibC
vhdBb6tEon0XSnM7vVkn5aYSCTYYfEiwSscQJccpYiKgozDmRg1QCPS0xvbCMQuLkmhU0YNleFJy
KcJUPa74HsaYTzv9hk8agz9BFvrfcpp6KtIPwjyBQxp2ibONj1RFlf0l6hKaEznF6bMUkhk5YD65
Hpci6CP18O9w9aokxme/DEh/F48g1ki3GZledpboCfLFqaa3uB76eg6FtJkHbx+8XxgOt7OXNbAg
7r1Ln9jtmla7GUth9fGH3O5yfEvnp8NW61Tv6NLeiprZIjvhc6B+s9c1TfC77eNxOhkOtkTQ9rG8
1NwBZKz4jb+r4ucdZiSzEPXxBVs6BaKyp2GM7DFCh2kwZwgZzbnanB/s3Tde6adMvLdzrVO+7l2H
kH5dGJp3OUBXVFrFJLoirWbo4QHYCf9XrXtAJbQrPTjmaISBnGku2E7BvAqZZ+e/m8qXUSwWTINJ
SaavfE0e8mfLfa/aHWZjf2k1EYtuhv4IHqfNiW9mLSNsITn0vxwZBY5HgUf70pg6VNHWYpWdrvrY
YK3gBNiVIKpYSmEP8Wg+AV1wZw1qvqQyYS4GgifblbAjq9QWx6HmulNmZyvvuf5VXJepRYQnKX0p
cC7liLdb3U/fCoZDXEhpooesQ+n+vTXwKzsZ22g5M/V5GiPEOqGYxkWBR/kIeIPb2NmpTwntsvEG
j9jd6drlZRsZK2bo3ZuM7JsV7jEGk5q9jSi9o4quL9w7d5oT80bqiCFbVM6BXbgMnJw9WRCn3nVO
p98v50sCh9C22ACVnNB7p5PLGxZB/YKQv9e2Myguitqv3hQLzxhl3wscpfLtKu4ZUEvVqE++NslL
b3/U8222mCcmL1tcJSXA0cwV1/0IlG2FaUwjAyK5bDLXho/2z5CDWECG3gDmPE8sRQOxDuS7XSmH
aaCfInGZbx5A+sDtJVNKTJq9Wl31OX39d7byAYnNahL32pLcz8jUowrz+0MJ1oEKqR8ZdMYXqWFv
MINQgM2h0A/TmTu655NqeYaDqO5SzrPBZfU/qdXoPudeYI/UKDygF0iBGu+2Ayd9wxcg3s+HTQyr
9Jl3upQ+64l+RvA7nGHX6UHdO1GTIL38mJ2N/jhmtXR9/4JLnR+DUarWAuV5rNFCeL6Et1xS09eV
Tw2tnPKDahAXmwYNeIX/RANlwonKyvF5jG1yVPcknDPgO5yAPzSFm9e2mWGlzjkWOvxR8mG7ugNH
MMH6d7i93HJgODHW+9NcGDTcPQwnL54riXGjupMQYV4aiBIu7sQ2yJSjiXGQN+zxKWJKtb3z3mr7
RqhtnT2dvC7p0BTSnymugFTT+BxuWnYkXMEoGDc+kEDpr26y7GlLPskyVBxw27tIshyUnnWyl7Wb
dy7gqgR6bBEG07aaNN+AEd7EYPSDoktJmOnqYBCUO/djj595BGbqIgwh6u9d1qEJ1FF2aOMMxWXr
5lMoIMzOux0HbBQ9t69KvSKDxLKvEp1XhNs/1Uv/wCvAauWnoChQDKDOc99aaPxIywXvhoTw67yV
ZWZdgP/QQ8lJbDmax9wtZdIjhM9ZwnB6UqiTij8aaFMnWnVrIRrqXs9lj2xmP4OPsabjnAipOUQ8
fzlpbi7hN11YS49M4kHZOSo4wThG1J/4Jod9I7PvzH1pl0A6nRLBSvEBdKMuubJqRYhrSbB3hRhB
ICl32Aemx5k67agQF5msFfccKirVZp8yGtpBFlSgurn45q5/zmCrbk2wBfVwvDbe66LRRzoiHcrv
lJcaYBAql9kUIiJznXVFxi0dKN/BHJpZ1sInK7j3MhI38py9eLeIZBpA0GYV7SSLx/ZiCeuKwoVG
hW1C6rGRs3/ff3avxXAef/zcRfkkY1hp/v4fGRhOcrpgEeI5628O2z4F7DJzRg7DFU2Lk6J408M2
AgCrLr9V/qkdGnsRhXoz3L0fm8+AQIv8o2JwUer6RUReOgOpewpflKGwBtcGOR2u+Ad4YYev3AtV
akyveJhCPvkFTyxQt6y4/lX/HdgMknErzqxdujYx+rJlDHYPb0KGDTBFRr6HhbZNICnH46PmtofB
AZzSr7KktMuGfPq7ph9uhwSCKauuOWbAMfO2wW3sHQXqNJ0a5qXvNjRMVnav3myfOT4pICtgmcls
WbPCoVNZPtuxkgE3LZCbFdIOCGkDvDuMRilNoJ9ORnCa0s8CpVQEgm0wGD60welX5ayoyMDQ9hoR
NXIZNsLwpkJ2p6s33LDIHBsDJpJTkylvpbErkVMx8S2ltcUXNEBlNBAchzE9XqHJGSfOLcewIYmX
zgE7wM1sX1Q6bVd07f5AQ84lQWo1ZyXBBvw6NiW48oNPUr03b6RCyqH+nJFcE1yDUMuuoaz3VN6w
LSoCBa7bP8RlvfToq585rAHPOVDrzBllfUsUyZ2qdllL4n091dusbx/sxZSbbT5Ww0qITtJFWaX+
2u624Wv3hRItw9+iPkmtYcfkH9Wmti/0ProyarzJ8ev6EHm92fflClvFbNWcoywV5TxtDlJlVbo0
f+NP/wNZQQIRVVp9jBL11lpCA6cqpNBFQyLdk16y07o8rhlE1WHq30TegxP9/Lre+wfS2xDuMz1Z
DfOXRWPn1GSBlcK03l213fQ3Fwrlc4KrAr1xh3WFn3FiZJIipB0A4xK/iTinvqIpwpkndK7RknCG
j+9UvSvvg+kpK5W1fIxoAnEyUF9b/sjOtHdIkzKhEJ61HmNgeDES8sE1uRIFKUHr2PTQc5sLQFgB
DFpNPcXRelIVwL9ck6BP6bzPArriFyzetGVOr50kHJqHR1Eof1sEjzk8FyRNTxAEMe0BknR5QBIK
SHvHX0PeyTmHTahlxYU6asBLVRzQu6WNS07cL7mnUAJQQZRNN2RHYXA5N9Ll3svx9/xOwatYyiDh
xHodY9/NH3vhFQ758zLmkEb0w9/Le+n4HyqpaOHJSr/Vp4LgM7TOq5hel7e3tCD2D8REfE450B+s
RqFdA1/HRrfm8h87fbCOZZJlff67uCJPlkniunVG9JRjZH2umoQZFnspkGpuFHjIt0N/gxKe1Vjz
d2z+A/GT7jaECDWgHkeP6OCd/2cPI5fBcFjcn4jONCFudBJw6DGnyPyFzK4GnD/tpyUmfhCEJqi5
48BQ515StktC/0a/u+VjWizefROZlMIxrys5WzLYcPwMI8Q8kfBPGA/MWT815KlEDsDaDT8yLlU1
OnSpL5Y2T5lwnSl1TN8ipm8U6RDO/OKVuTUgYPCUDVg6kqJjnskmWcvPwav4wMVO2meQuMzJjS5Z
DPRrJF0izm+C85KtIUNUE0kfTmDrxjSSd6H3bDBWMSPEm2oKtzDvLs+1Qr7S4KU7ZH7Thh4rzLqg
yqahjv76iVYsFNuI+NLwsCs4lk/7/430wY5x2DSU7uBRTfXJp6NMIqdTRdchSSH4Xpfqs2C1spTU
L/oovAMydaIrRdObd0b2If/reWbKXHQsxHfp7dYonzc2qUxI9XxTruib6c6/ZQj2eO+Uh3o77/lZ
tTWdzQWDAd/S6Fctc2oyM7Bhy6I6ZhfaRLFQrVeXjbaCyZ1HdxzZpc48YGUAJmLYLapfrRuyGC9a
rZwgiU6mESwRR4qtQw8GQomGGJVOPLSXW5i8XjRjOHzJRnp1ZPQhdZq9DEe/FzHTGNtYANYWonkb
GBeUDe89GI6zT+xqa3RIAR0L6V6+yJ1Dx6YeNxurm/G+USqsKUKRX2PFX9dNkYoQGS/8/8qDfRTl
9eGPtjgFn7ap7qiwkSYqKT0kkgdT7UaNbQugWYXroO1RmAuPjjMgT28DZmWNChFpcc3BWkSVJuti
qJ3e65tVrXbj9Xy7KVx67462BRxVXtd90uF3YqtNS7jDxvci9pspv8ylBdQe3L3sBjXAsWGKf47S
OrBrUv4u+B2qBH/DX8Pa2MYT7vW1xeqGXLjuyN/E2I4AGyvupbXTEq3ks+0/30GUnYTiLzIYQi3x
aef5/eAY9+P0PwhDSmKyxvd1DVjtp4fymVsSQ+9jDCokURhhByP41B55fdLq0CbfjUWNm0NEyp4e
+9W4EXAcCQeYXtLvT3Ia5+SsMdHq4xorTHf5HIde+ax6gVbqSEE8VXoiJrVhmKLuMre8AzdmV+6n
S2BuaV8BbVQpnXb+ue49rwsLDinT8mEAecWlolYMZMw5TPYQKqOIg4HSb+hETav391PWuXrwUp0a
mJJVjmHGviHJndJAwcVB3YFLfA48tEEGId+zYV6b0VlyW/9Gv21qa0RRRJIBJ1BWFniavKImm2GY
IdyhwaTJxE4AjSaYtT2Chxy5LJZmdUqGm9KZdy3is9DoBO9ExF3MtuZQAXkMs1/VVQ3OphDe8mqF
QQWtV1NZq021H0s0QKlaY2MS4lLD3HWnRkKJtUmPPH8U1mS4YC7IKMcmloKn18WNvaxBhV1L6CWr
DTWi6k9jCtN/I2F4Z5Kan6E3nTVrrr1ESHwcSaUg3UKfzbPT7JKGUVCOVI07VB98aLCOFYvx2x+T
8rqQe8t9em5zLqtbbZf+di/5NHu1COaHhz7o8PGPfqYulyharvynCjCI8OhelH3O74Ejmyr9Pknj
bx4yk0JN0pAQdLEg0hkiLIFaa4V33Tym3pegExMgvdinBMQ423/ldTob+qDcJ9ftGose6cGWUNyK
j9wSDV52pTngzjfMnGFt9CY7IiPWWR4NM8jpMwMiGnYzXQDS7v8Kgw1L0xsO0LRuPB7gdY5kd4C6
/Y485i6bbSPqnTACNRdYC4i4svC74b8acVO21mPV5iNxhcvb4W2N78w35WQKg1ES5ZuDEORcviOF
5l57n3nj1UstyEkPPM3PXImrtKqjZxFjqxrCrEumRiL7AN4b9Ift+aoy9rtrVuLpdjUd9f1RWdZ5
fjX9nPl/dHFNLeHBJtyisxWNx8e4fGybMQS/d5FUfOur0hm8jGNLsjaXCpJLIVIW+67Q7UebKKn/
waIsYCgRLdrk3uio5PIio37mOZ6DIPOs9gia7OJQTx/W9T2rj+EhpLKlvYpIXU3pJZSMJ/BDLwCo
/j8eOg67tpS2ZjTpOaLIX5q4Qk0pMgEPIZzgVJDNxNsnqrCeLkzPEkQt/RsJL7F9GCIh2/LQit/v
9zKJVH1scRSUoL5pZdoQJ9z25180C+3VgKa295e5J+nNxUDruSRhG5hFIHS9vX/Nh3gNaB2pdQE9
xQi2u1Ukq1h3w8G/W8jrk0U5WS/86Up4l79KiWRZiMrjiUNX2Toz0Gdvliopu+3udIJxL7T9TyS+
3p/ltniGgUYSwwCzEZ5cCu4+T1XxHyTJ7PQ3r911LobX4cCFbxjqqs5UJ20u8huqgso9hC6UFX5M
gsR2jEWepoFlCYcZX2vIsChiNL4WsDnPVOqNt3U5iOtbIXH2ksBOwqdq674zXbAZFcnKi4J1vLEW
EcM0kejeupjx9dIgfKmJusxOQu1dl1dLIBcs5J074QsnZDI9r3RXUf6O1Nf2czH5I53c4sI4MGIF
uc9D6Yk4uR6U5SJDRdzTQ8ErKgwsBb4dZDEQtenMTSglrUfL7MgzldQeQfNxFOJAV3/JC6tzaa3M
b0GL+u09sXLhqrcrrYdlKNNoLploOc89Qnw2tl7h9FgQOmG5pqG2VUu00Qd+n4Dofwd5Wfo6XWQG
nqaxoQklQXTfMLBur7Ywj5vUsKV/iG0KnUYExYUA5hO/6As/z/ylwYhItopKvcF53xGG8K3yDNYe
6FabytZB/hwDqP/VtIhYGzX4sXjhec1r0BNjzyeLpTNMivs+7M2L4kd+P9ZawiiWUINsvsENsxZ7
IRGfdsxFQyKu+sKz91Cg4djk1wCLMqrUOe7m3R0m+onz7fEz/YdzugLUFZoHeLP5TTUWfqE+1MX9
47yxkdqFIzMWhptE8EIf18cwb1+YVWiIOLilcYjnekF3Qrf9f8AjOh+0aN3nD0bk7fmuon57j2kS
cF8SpjjSgoxXNN5/vrn6IGdh/FT+xjOUihEhV1Gq3A7tn+5xuNltUSvOqOXF0++iFGhV7ccwy54R
DzVbt8OZtBx6FgvGPooLTr7Bw0PKEfVG6VF3L0BR9Wp2gH/oFsptBsmA1oToJt/HyVy8BQL+iM1O
vQh27MV58xLTzQGRnRPakbytuO7plM/9/2owjI4XnuAwRXJoipoVODWL1//u5bsatLJj0bfvAYiH
Ie3Btdx795874Lyk74Itp/dZYOPpTvbm4J8+fmpv/0tg2TannkfbjQjA2C9/mGMyJvbW4f3VcS86
WzigZae8ug5MD149R2j0z9lfMTL2UVeVQUiQmwk5HqvH862+ZaHA8h/Q5RS0KmQnJWQSVQ8XoIPC
wr+HQSCvsIbbv3Z31Q8yayPN/U8z/MWQnL8bR+rvjv3LdZnJPCzvTDXU7b26v5620A7NsUYfEuHw
/KSkfhD0yA98pReomVw8ROviGxY8eIEjb2c/OjV/eFCohkwkJA+gGlbVKG/EG1qZp/Hgw4OAJ/ke
g9MGYOA8Wd6mXajkjFZXMbwyT7S/W6DerE2RucK6HWlYr0J94WN6hTlip71DoCJUvM8Pxn/KJKgk
AeUlQlQeJlsTHuY5MIbJr+WW37FFbb7wQ99YxQrFYqlUfdBL9VRiT1b5q9L2rUATx0OLb3hB35+p
Qnnqvnq5ZKRWcHBRuur56hmYpwZxBBMFUp5HvXWI2KUpwv0ljLki+yQiJdGoiDKPLCz8Zu9xyyVW
u4ZI1T6rUbROPmI/q6hCGuaRroy20RRa3DJ8WOZg5WqKLM+Pdczacar1o7cqUQlQFBQqA0DGa0lF
BeSUXK1NyUyg89/eCMJqJfWMZ5EsLR0h0WlWzj6F1Vo5oUVzTmdfCb6cuJDTuoYb6u9h8tCx9KG1
gepe7kHOndvy8/83TEx7HrcUpNOzPZam0FvTAQWSXyRFXhGvrUujEqE/MvK+yq9qSUeOnPJxQLtg
wLl03In5Q2iMnv29OAQXaV8QqUF89/61E69fvghU5F2yhjvlcCqX8tUDuQXUG/VTQQT86Pf/zYjz
SiIee8T25pQRchLQWSq6rqSriB6G2ef8wwc2F4SwMqtpBGXLel/r7w1EJUsAV0UdjjG/lIk0yf5Z
X4a8K8AQe05EVkhMH+GIqnssMQg97z27SIuu6+XThVWhT5lcQ/JWFa2luBkuVzZpPIbsSYHTpbpX
VujhskcoIbWy/RKp10PWepnQSajPbusPsOufPUI6Y0VZAnhgLzYiAEjGLhw1RYLnCbpmtuELYEmE
IBz+1oDBGVDu8ZpyRqqO6XYuiSp5yv9ujdFKlrW1zYYqh0vWww7FobR/6kBIYLwQT93c3ZmJ9kCJ
Zjyawo2MNj+Db8cfzFNk3aFAEwcvDdUSvhyU5AbhqVlasoQ1QPYRH7TkEyZRaj1aj7ZFPfPOQ0Dw
sHHuK4ac4zx+jSf97JmG16b4v6QRvOJYkx++U4NszimTvKyat4HeMxXhKzCMqH3aKW9RhY5UmG5T
dX5ziVoTKWDTA5+J6vikmeFFPg/uQVQJ1qc46VtekN5luKHpQmqmGVeEqYMWFrBbpoRIkFocbBSi
iWKv/w/a1zRXDNYTRFW2e47QqGFmp1zy1irtzLlVV8g0Kv/DAmr1bNNO6/M/X6dqAKmPB+JF1Z99
/YLmUseRXbQu5YgtK9ojq4C6hnxE/PcsMPI/hlYqZFqUqIgQRBlwDgcQ9YnkdqR5OEOGistJOqcs
DrqjRDtDaxZ9selSJyUiad0BH4gxF/QE04hmQNm4VvZoZhY0lfkAa+RL/fare7Y+8Y3efW8aNe0B
VMPTWz0fqPcBYy/mt/cQx2HtEGHAp7/HOqDAbB4euRGyL9LG1op8pAdQr4tWTksXvjRDiqgL69wo
UUOMQFjNM8E5AvKwqXTmRfNTctc3ziz5MZDceci2QjB2ENQ7cmLT9B/bc0k3CZZB+mTAYacn7Qz5
czutJ0RvT2ar6uS3VyF99A0dVjqJJjLI4Ia/8uBLVCaE+KAwZIVBmNW6thKyUnk78e9KH0mku040
wD5s0FciKTC3E2+b75XWdLDT70vVT4WwitI0k/xoVpvOo5QT0SYJ5OHCGZUiXOsN2+06beG1TolQ
SQQ7hvC1k+Z+LIvKemFwpWzLqaKVXPxuyfND6zONGNidTJHp7QRgj0DTrCZCzOo0wmoZHfS6e5y4
UkMKkfO8JjSyCXuUHDcn0HoPKXlrY7kv+cgPqDsxxus0JDUyQyyEqHr1HU+w1puyhV1LpNs7NNL8
5Y3jbU+wiE3EiiicV1aQc27k45wbMuha1SS75Tspz/dTZG9CjeX7sWn6+Bk/mMEF+dHBx48VK9kX
mevRoHCzssXY7X3vK/KzsWDbVokppbUyalGiuqaxaTw45Wm75t4VJUD7/+TIpC9dcWttsjXp210f
RtnRdBRLiV6/DXbED7h44IHq3Ii7KkN20QdymvfcZyNeX+tDAod1og1sMZNvhRaxjjpTnLZU+APj
wbZKNoOPngxRPgcX2o/hlyXGFlnhPKkX1A2CcGuwvoKml+tFVvR2AU2qe77cJ2PWhbbSS1/5TTFS
4RY37iEfdVG/EeNOQbIovQ5qL25k6lEuBP0qDGhOcFQL1jStzsTQ9nedoOIlh3LE4INvmR2hHm8a
CfBS7jUxJBLzkexDGEAAZnIJM8W+lx5bcMg/6GwiCRtTfkFd602efeB77CJy4RJumYF7rUNjkWhh
aLIdp+k0PxWmea9O2ycjP2/o5LxY6sye/kAr5cD8wwnqOjZg+cE9acRPVUUZtFaTDqd6I61ZJDwc
sKMCODfTcVPjMh8O4gSRYxRrvixqqRQnGo1+m+l3Zk1471BkpTveKio4GRTqCE4wEXJ8oDLAhyFq
Bg0qxkRxKbFPxcXLX0ixEsqIO0kRJMZMQVtJg9eweaYJBnB/Ns/0MfC43Clti+2rsGlfe+IfsJty
DILLLohOFjQVVaGD9tCj8iftJC0Tkcg3LMCJWBb1FYJnkOeW7vpJ8ol8/p/ykwgQsaOD2mheGFdK
r65cbtQTg3ZyXiIfk3btN20MwVcLwNQP9NPWXDSA/qyR3l+mk71ST/CJfrk1onWiWXVnywlN7V7e
xAhmmAEkCf/fdo7WAccCTph8hiZuzNx2FYWpT+jaZwsz1DdFXB9AhjK/R+a9xKQaJ1f2bJLVid8S
dqfSqyT/3TzZnUpjWws3Rhoth9FSZc99w2Btowe9AfBFQ3l2vbxpr9qJeF1i58RmvuIRecCfqP17
N0R8TnGtTg8QTdI1SQxEz19BKU3qIgYz3deC0hCAOX8GT7+iwkec+MsnX4oN9LrbsDnGAUsu4/17
irLL13i8AHuI8P/8pSU+nOXabbqjkEFWTjk/sPutKHG97MMfgY8vVKUc6XYyFHFYcGATAgkW47Vu
7yCilkArHODQjWKZf137r9lpvUMwJEVwhubvcUWxLmDuoyfSib96L4/a+V9eXMl0oKe+xzA8qLq0
46YiVhkqjOh1CWxho/i6YU1vc0IPHK0Kfcl6OxqArQ5FoCuEUxIf5/TFfs/g92lu2xlowLlZtEd8
xAcI5zWIVAKNdupysbuBdbbQy4AIPkrLq7jkXbR7IY53MEUapGn80578qkRyJJLoyUxNa0N3N91c
4FPX5lMcXbHV2snx4yeAKa5ZGmnRdNJhPebq01MXtuhZI5kuAV3AE6EFnpNSc4DNGsD8jtpUKMiz
L+WFEVZgB5LEf3GcRGsdQQLSmVqh3TMTZcsbzPvzFG4QwZXpHLYIfUg/93ipXHaVy+9C4QeaSnqe
jM7BKC1K3sFy595/Vsq/GaI98n3nJ14gWAQ5ARMI6heSXQ+aBjHyTEaf27A2yDZP2toogQho34P/
X5FQUh84DILNueIBk2uADNEyybblHfN95nJiSyMH/buzuiJFsVytadfjQ+CeCF8ieHSvedKYbCC2
7hxl3IzEqrv2DCE1oKEJ38C+LZmhGrmONvjpAOcz/KBn+UvQz2GzabKFUI+31cs0eZr3e4ISb13V
WSldYMRLMwY1dS+naYXc1+Cp3ZPfY22ZTkKeR8WWoBCek+aC5t/sJ75igNHeAmn9zidz9Wh2A+0Y
X1SfsoZA77VLIkFQobsBHpNU3/QDjP1p2k9FMtiB+Ik7i8Ejf2UCG/GjqBYhpwfdmxpksFYkbO9d
7G/bxBL8NSBFfvHbWmecDz8abKQiS1dAqrEBK83BaNuFBRWjUXrCfFcsIDodfxK0Vs4erhqzC4/3
5NAM+UhwoJCbdtpbn+674NjbQ4k4P9geaHEAaDFMAlpk+X3WXmPdNm0F74Vjv02DtT8a90QJ0tYW
Xe0pDNdjkjpzzMZ0n4s3NCZsKFMSCbvg0qRk5tFpP3vkqfylIGdCd9EBWJ3CDREoqynA5fgyKWqZ
rpXJGUfK4EGeo6j9JdPcW19fgS/OyYAKsuqmpt/rVOInEKRqd89dU6O9J2ic+7t/jwI2vWFBwNYo
UNRYNGnDbhq587obwN07I+Mng2EbqxRL/5y1tMJv6XSwRcbUXQ3u8zGRIij291OpMPm7VeR4cNuL
tiVELIa6UU86YXxhyY0zpfF6aLvYygVctesTOgpiKth3qGnTFddRqS2KFZyG3gksFK3taBj0QVm8
NVqjpE+IPhUHU60cZ9+BAzm7AvjG7KWMgwFNEl2MVJAra7vcAUEQwl5Ei6Npw9BOhwhqUz5BXfrb
ueONsT8mQ/C0oWwjbGfCRABi7sBG8QSg1vmxdOgG33c/J1Kmg5Yy/OKFuCKgZ/46yusTHcLNc1Cx
7sSLqgzrEY5Hqtkj3oWjr1B54ZngaRg62MOJszbS+UuP47cCe1uPkLVsFiG2WuCotto64uSsHJin
f0MV5bjchEokJ0m+3ylaiAqeaeV5afOj0hZEt4ZSop2PCu4E5bQ9C8X1EB/lNnrjgzGdh3VVF098
vY5uZlL36Ii6w4f8MzJUtHEVhqiYh7H+4JteVtkkr/sE1EU294nt5QsmbjgtBzXb3/N7tvMD8v3u
Kt0txSMfmi2bbEQsZL+EaYj5deVBdgbf2hWrlrnujqWDPDxVB5xpSCTMYI3fYl1aTCzlCkVWdcGr
srp0X9tiJsL2NHMUKMkLwdDOANhuI93Tz/TG41usDTc/qxETFLKVN/Pp2kg647fZ9JpSntBUp3Gm
eiFuoKUuqU7zh3lwW0sqKwyw8j8bVoAYO3qVF8dfYdVhtQhUjMkaxN8bcboVf9m+qqD/w61S/PHm
vifusaCED3hmzb63pc9AyuGKEH0UG8yjVslYbMRH/Bsy/wrMl2DTNibbmdh3wCwoEMRExNfgUzdW
lj3c+xAVL+12HCAFax+2HM7cdQszVT7EyxLyCVChTlzVxLd7xgKaPxX603HSy9bJkBvAEScaJ0iO
e2Y7O835gbsrlN2rve0Jw+QeOgeY109S0b43YQXPdy5I4awZ550qhRQIP6ynIugIQoHiJxRt4r4k
lX00AVDD3HBiFW/R5BrlAKZQbPl/WwQXx4FDOuJRYnMeMrWr9+i963fymxqq8YtO6Upxp3TDKkwe
5ew579GzZf6GfbTqjE3jc4d/1h/tq0edEtc3Qa42WfgaKXLhX19OhqSaJq4KuZVhjrYng572OUa1
a6+53GKISoIeAlDfQgSQoAg4xFpO4Wo8EoILLk5SRQcXREoLo+ectCePfHdDRTmz6EPBrYvVn/gt
3PIQRfwcqO0GooPTlCbSSOL+d1HzDkjsNdJ6eG7DGsrixXi+GqjxR0UT11OnOnyBYbRAv9NyoEY5
SY1lBj7X6gpEwELFgMGoU15Bk68ctH3NlSMI9cgBWWMDxyP/70s9JySX5QO5ehRZTTLwr5H51Up+
v1DXHbTm1kQgHC/oP5SzweVr24bQdg3NzGWfBVISRot1pH0G8hk/nWPP2QzaQfCW/byVF5a4ZaMH
EEZvPBGqhfTeRehQnbGWI/AC3kVA4nz8cv6btdWBNITMrYzZ+NJHxIy3/lH2iOXEByb+3anBpBVd
h9jBk+Twya46A8dZ+UN302PwN2TkpfMpF0SdxldxNjU6CcGOi5/RgIGFpXjOPn8xRdAXANXFjr6x
iP9IvHjeBmjuichTMffcXQb+MKoCXEjhtQRKMEgMJFF1+8qT+9zQeqLQkeiCBUOnnJNySWYH0SQy
hje1KP2hPI4nrJLww/Jx1V5HXWqxK1WlZe1vYtU+IVOiIRm1hp8m++kRL0nqZ101U1FpfD/pz8+f
4zmDWJYWspLAH1wmFznBa2c5aSHmF2H9Fc074RlQ+Cx+ci3sIDKlTKo1MZVDMo0BEfGlXVvc1sBJ
nlRES1dRN0CzdR71jfVAkzJuDpMsWndjawC+xgKb9Cnj5KYyFQluJxLUcxEmQBtZSyPoPR1g9kt7
dxHa4t3atZbh2cg4XacX8TY1wNYemVaEMCrhEeGG3CisjhTJgnmmyCRZ9aCOMnQc8YQ7+zZN/OAn
NQ4fb1KfFkg6h/AhhGXpxqN7jPbHL2VP658yxWUZDomlG77FbXq0K13D7/W6snpscsK2LIFkT+mc
KTN0Kocxn2XFgImpeW0C15nlLiFZgSmM5QZgXTZe4vPzMKxzDNzIUM3q3QO8zJA+Fbs8WWq415o8
yMyHKdMco85Df3sXyq8LGSpDmAXxerSiYS6zz8ruh8O0QUBmKy5EFTHa8J9moR8rdK8A7+XRP/Q1
UOLfP3vLty4VsrjbLJyMT+2T+SL3MPhEQxZx3h9e5gnFBgKSoJFRjIW1P9C/g8zptnZolKeDqdBf
IGXjWJs72eniRpWDQF4LbAjvQEe1jE8XQ+cuv3qJZO6fSRYOM2PS0927JkDVzFWzmxQEkk4VRpLQ
MHjQiwuAPxzKKb8/NpTLMFxXq5AS9IniUY1cDQnBnxhBSZvCECpq9h1JO5D4SYTi7rEqg6pRbzWM
GuojJggwDnZlJW6KG/AmmjMcKmbgv7iUC+0YikB6xBfumCQwYHjhSTGfzaKZ6rsRm3E8Vnm7iOW2
b0I0Vdu1leryZAss22Zd55zDDvc8uUmTG+1jPcUzLZuo20MMQzNi42niKwlcdJ+YJ3SjJfsL3i34
WGavBMTh+PkQ090363e+QdirlT/nRp8/CRuQBhGabcPaCGREVn9bEodHCUKCBbuaJX8W+66w85VQ
iIz1GpU5OUAorOMv66BvKPedbfZiZiujXQ/tfD/vkMNrtWRtSdAvJXiexUzKKhwGlNLi6XmmTMn/
fMsKiUevHZuC5csHeOaUjOCeqZk69P+WhFmt22jwJO3FBXeFWVDOAI6kJzc2l5GQBbs96m99xCTp
83hpK9IFcliLdubTFn0FpSH9hih6loZfadYyzGevLXMD2Zln7UMYrqCFxdXpSPijiKBeTxVh2isE
GpuPEg8YaRx2xioUCcC3ffM1OgP3G9VCUVXkyA5fCN8Z2DSzXTA621hqkpz7ztQ+EFxF3HzXACJi
p09T1MqRmrX5zgWccj/WOmuwqrPdadieHdmDJ/L8pdVyoZkqrNkdkh4f0+WhaTQR86r0K3W3rLzn
dO1svMQ2Rx64yuHqfjRJC13xAGyTXaUGufCWpfO9Q+pkzR0HeAcRgFwSVY10SbTlxzB+tc4q2YZA
c6nV0sMyjq1a3iFs2/+imijOVWBjmh/cdmTCCXYQxVdKdDm7oMS4ctbYamBWVSRwiRlaqinkt+lW
Qj02isCPjJlfemGkM4Z2qPZoZRsHUB891HsosHDQZ5KECX/7mljJaWo/TW02/xMUt5TWxmQ82FG0
qD/Pv1iT/xNTvm2VS2YX9v0Lc1M1+LtOecWoVpg+uVKVRbR9HF7QDDZ6NsK8ztpVVzwhBkE9Ucwx
6P9p28Oj/YmfbAdAovkkcD3a6uQQikrC2mI9FBLCG4n7isWyv8PVbRmhg1FlFCxZwOdtp0EXYIVo
vu+6CD9HC7Ls3V89ISHs0q81GE88Ibtr4MPVhzD8axuc1/UEeZKBLT1F65vH/TTqwxcdE6s0jd6g
EP3TiwRkKsF/1BumfH2BzWrPLwEOE7wvZUwtnK35J+CXFFaNS1PCvZZkJxl8O9qWie9lgZo47IQ+
BF+bKNqLZlUuQiP5XOfJGyMK4t/PejQ9oK1Mggkv2y1N+I1/jeOMCAePjmsEPEYIXyXhH6lRtvB7
/U49tJDLS9RVLu2d1kemrB2pVoT/gjEYqsbc89ZK31IyqOKVEZoZYLUq+1iZhrS8DiR/zAAs5+dY
3erPpEpGt3pzZm9m18T31CizOSua8PauqnyY/r1cSzXO8/sp3x/o4+2WOy5kA6ymAlMbaj+aaVjJ
7pBgqVOyRsPmqUUGf2mt+/LMhMxJSI3lsonVRdlaXQfEgfzLuz2/5j2ojW3Ftm//xPsKfd65cgc0
9vr4UdSAhSOD7WRXMC6er5YXJ9SdpP20CqMmj39tuTHOajDTyhZ/51OrllAjTLTlO6C7+TOmwXWq
/0Fja2R9zRO/uevyJRQqPZ9l+dIgXTsFH1fajrgEpgaakCKJHYNsunzTeUZe17mEYDVSHYtqFWeD
+xTWhGJGR8h2dcCTTZOYAof3I8lw4fzEs3Z/Dcb4jobnW+BLUmqplDzByCsP+gQeHc6pu0NccaMN
7vYxwBId7XczvK2dVVHtH6zoRSEBXuKxwpZj1hlT1qpOZgsTIns2Vn5x6oFIdtejVz189Bp+oL66
AG9Gk8TZy4PfqZW3PZ5AmXP4VB1B8eAbLqpKoCFd3FxZClvL9Hy3WZlyPTEbqIQQwkporKUQE711
7cMzhqxn0rJQ/EL+oRd1f6B7ApYog5L691oMRJeniC6EEm3i/a/a9oyoYCO/SYlSSZV5nUQwpYWW
soY2wugbuB8E8vdwloayCmn30ZeR+1kF36MKp/xxdSo9WqL0FI+zTOuNJ0MnGFz3YbmTTbh/st7h
DAgaWrVB9VapvfS2ojUD7RjebTzZpxn0CN1Gj19yoWj1OCMbwLiMjBkY8lUxUN1pNKhtGEYEwbhc
b6UGVEiqtX2T7zlRrfraJTdjOeiA3x4IQ/SoKeUka27bt0xkYNfMVPcsxPiBpnwlZaZDi86fTG0q
EWv4vlmAf9+iWQxf8dQKn50FfNvEiaIOTbGSsoHzCqBdKnMQihrHN+Ic7L0QvKT80e5OtokJ2usT
c7r4t4KrzLOaud7HIDYeS4xjbMdY/xW/A6cWPXOIvoZowLqQrRQ498v2iwgBzNVExNV6BtBVhEyE
YHzB52XuvIIcrMyfkpejyeas7N1oc9EdfsOKX89c+P+iPpagY2P0AMkqW3HLmFEGv4huHiWlFGA2
PTc/peyPz4qK2nxh7uHpPa7EbYFgB/H0EfC5mvzKDuyFJrQdBR4Ob0XrBfQgzioAwIBoBXGxWVsb
IJuRfIxaL6OLE6ngMk9cnSSzxMfvI2jg6YAaQjgL3ftlwenDXeJu24IE8tRYufSMMlbLwg/Vgyro
2G0uZevXz5wj1dXwd2whnSNbBiW2QIL7VEmx8Qpi607kJK8J9OimmpSJ2AmhjwRdVttbsb0x3o6T
0Y0SrhCuPl/QL7S+TnyNAgP2l/AZ5RMt4A9b6nzF9rULOSF+27EaLmlxW/rNqWsSfo7YY6bm48jJ
CYV6TajFZMSeJM6bfS+p/9dwvE85a8D3AJt9asJxQ968VjyFFn4KVzrOpvBBA5i96mXX140fL86P
Uddot9ry2W4aXun1/duJxuunJMeKZ0vkbxHQTiKUX2n++3h+q9gR6CBC54qnJykB/CgWtH9Inp2Z
dlzmHg4vkwomqtwQ5lRk9zHy8CbGcE9aWkSnC6fPNI0umF26AYihCmVtYVbxLSpECzx16QaonWCM
cBlbvkHv+eEsDVtFApnFz9t7WWlhJduT5B9qxHdX3NSOFUUORKRugFzrGkQ6oMtNap4V+Sm9J7HU
R55O/dEMAzS+vl8bp2WZ2sNTXzAa93Fr6CNKNb51STpjQ4fTF0rG3NgmrkShMeX7z6dOLxmu7MIX
3Kd2jNpNJqXw8GZWYyN+RzeHay9bTVGm3PVZaQwKfSLTrMZJN2k+RL4gBoRv4ejVxE30TPzgsou5
sdU44NpehohTZcOLaX67xBCqiD2tppOqtjNfuzFzGbKMVtEDwR6kGoA2VOxjUWpJpB3miC+JdliO
iryM3E0Bu96yh79epYxP3ZaoRes0A2fgv4BkOMWhi96UQYL5lmCIFPZpG+zRuiIHp/s5tComx6+H
vTLuW/FIUo7w1D/tIeRABqkHkAHZTsouhqgRGttf3XxvCJvTYYb13YK2Dj0PomqEdGfYazhQ/3FP
mtPelZsIuY1ER5jiY2QR1gLPAayGbkQd5xpWKxEBZvxIPQ/G1QqEl5f4UuXrOm4YgXFt8ppR5tW1
IU5qF24TDZAhWq5rH7b4engtl4kmzSlasicELs+4trxGfOctv1vlHSr17PJtSKq87qn6QUUKMh6T
DAeHs4uDcyzaY2rQn1Zmr/M0C1Lf2EQi3VU5VY7BLvwiNGRzf7aAbJJeqGvnudkUs0fKoeDL0d50
/757vy+Ns06d9YAUWRWdnanscBFhCOSrjsWtfYQs0llJJfP96WXrQlMn52gJir6h63nGy1X3ve0z
kQjOzJf+eu0UPBiuSIORbOE4IIDdLQE3tcElcYdNOchkRX+qiNABvafd0rQgUJTRwlUPqf3NYJIq
IzaOyp8Sr+Ln5LNYiQ8sO9c9IsV3VVboOmo6EvDNT20HwGRtSi+6J1CoANZOxYFIkPJ0sAiiPnwb
GmTh4WwAITCfn7/0kd2hjIlR70q9e+X0CIgz+27DpfHrpyGgkcsImdZCz6ou1FTa4w/ZB9DifqAR
+w8WvvZgrt0tfN0Qs2JFgVt2VugyAu+oRLU70v4BUikekhmgU2XPZhI12Gkm32Zv91rWXRB/zCOr
uzhCvQjoJKf1ZMSlbedlFhpZcEgRJ2JbIE+3s32Fj0GHAc04k6OMIM/0ZAXtbe5f2pyV2nIifZZ5
rG4my7HLKvPADl1bdLekkaqJDtm7BEhkfk3jQMlqjN2FbIXSIiLS2dj4iZH7Ys9FkOeBC2O1l+5m
lgMDrJXpzyhH1/GVeDjPLfajqTjeO2cZih71uBkVtq1l/e8ApZKppTL52jp1hCtnJj2v9gdpApiZ
49JrCaMsGC+TwBKOLSCxhUqQyNhRh5D+pclkGoTh6QF6GE7DELDp1kydwjGV0OoH+f4O3pSV49Rb
Ohi3HQKD/zqONpUGic+64lEQVkgfvGC873mtciO8dm5A/SvGrh8eG9x6O6bZOwGBpVKwaIrsQpS+
0mfJzF/Xkmtami52pB3asmem06Ds/DEey48kIU/J8tVJd7+sq50IxAlvgVUK/rSRuvIUgyXYu7z6
MCklNYtkwGgNmOYWgjTOeAHsnaX9jKiU1fFEQsr/ujfyC12y72uxOlym0WLXKr3/QJjFhb3vSHiv
dA+nydu+Kdjpieet/+7P7qcZZzdnYxT6tOfZnX8ca/N0IOUk26uKiy13nWHf66OxNeqxUUxaAYTz
tK90abOqcjXY7PSI1r6ywj5dEQH8RNAVcPGiN+5A+N9ujhhw1XiehtiLVhINnDWT40oB/gKy9ooP
P22L0+GQFSaNwglhUv98SL+jy2NCFV6sc7v2KoypBrNRV11f+5PKJK+IL6mNN4oXWTBufpNE9L1O
KrjtlE2MHIrlxWXCZ06Ngs2G0ilIv2IBvxabUD+yNVXTBQ7kijEpQ+YFl/K2ypdta38Qb9vCgRp8
2G59b7XLhU5sNwKbLtNXf15uctUcD5kadtWbLeSBBI6h5bjvU9zpAKgkpLhDZ3yDAEAijcdHhxI2
+gSSNDac/Ifspy6b2MrJ2wS6FjyT0j9SXLivI+sGBZH0QimTAG8+i4VGBAbWx0FxNnioL3WyNc3F
hJnC7ktZRg8R5wBmiPucPuW14w6ryJDmu/Qw9XMNthaoY7YePBm3MGfoSJ+8i8NcV0N8SOc16/29
CN2h0IbWZnOjuQlg9VVMuPRoeXslXw/hDMxPVLfL2Myh0qRt5ttwf0/n/cCpUpMphX3JY4et0Rsw
OQxOeG0sDLaMtEgmzVj1vV4rzkEjqhnzad1S9Suk9zRr+UFxwNTr5TQSuBOyz38NN/6DKAq87GTY
tBFvZ7tVvWb93Yu2HY6JWoF/SvxIuMoDF+nf508KNzDgQ6F9jH7i2LAxS9QUNFekyyP40LwHL4PF
pygFQ3X1DUmHaatnMvjvyedxWRENbhh/gDLsnskxHdS2/AoED+FyDs1RMT4HE4z/NgVNOBRA/XIF
LZft/zMRHyi5ww3W0MYWUgZ0c9f6HNbt5a5Sxx7YBd3h1WoiWW6auiG7XgGvWrx2U9JLQ8FmAVly
klNbfmepE0S0c2dbePBu1DSpaBoyHE1apQnBZUuI6umuy/Tq57vSQKzFKtTeXLep1QSqq8d8B/R6
o6XUbk+8EHcLCAw4bceycPG6Wc7/Gnp9OhIYkcN2IhciFCfU0RJ4HmmPuNkuCPaG9O1nQSDPf3Kh
BW/bIqMDrBRu05wCuOMNTc7afCUh4SnwULXN+zBLtcw2YUedvRJY5Yd1rlbbnnQQVp0EZXxTLOpL
QKyfQrmxH3DH1LNV+RR+ZbTaS9SqiPqb1JKVzkL+weASDAqNT1Nk6RPfH1IZidojffWgfUFk0R3y
GYEJT547t8f8T7rHtSwLv2ghhxyHdY5zKsAtEPl71jj5RFg/wABIK8kVIBCmo0B4jNIJ5SaqRs1l
9m9/+F4YA6cRdvmbdwAp7fL8JsW9rddCnryXPZo1gdXfEcN8IWsiVKEtcTb8iI7V2aZkf/3izn/a
UR5rC6KYnv+i1ktpExSFx8vtSYET45tu+KQqSvybZJGCMjeCVwFJ21hoqwNUbYokRmopz9HEM8FI
6rpv/b1BaBS5u9rCt13Q9GeluA9AOydu9mMAYLI9HPUOFofO/FGUw4KKA2FKOa4hP9T69r21A1qh
G5uOexoOGBrPmyJpEdSfNbk9NFps8RHKe6fBvhkGkhCpt/mvSDHbrMEDKDJAzw3By5InFLwx2reL
zKSx3H8Gwwq03OxjpqLjzlD2WrFYvRIFKG7NS6tUc69f3P9OaPwOi7EC9NIR77Lr7ZVyfqrxpGKO
TteBNn+Z0NTtTx3lRkddmWOGgcsf6+T2qkZVYLvC4anYohQ52O6vPGNyg2u5uzDl7asTJyUs17q8
EWyLJnzTX41RyWc3DO7oji5R8zrIUXF1a5Qzf71QGa2ZyRvCsxJa79HPGG/DRjUOueeXVTSJUCDa
zpGW0RylvX6FhsHC+Z9wr4EIzJwoQQJ6hQXvqt1jUPdd2xB2x0u8O7XHtvmXvq42Wk60Oi/5kNTs
sg1xKWIujNMQXn7GlMCyoPxSLlPEUHFxckkVEQxn2B9V89lunickAq7kWget38AywB3IQY/z7qn7
cAtQ3auW5mW+SuYkc9LLVApq897S0Rk8BukBz17TcSsuTQXl/6o/qkzSE0N1iqCAAdPvhvDK4OOl
mXK3M7podeAMiaC9lWSxPxEbaGBuEyAq2bajEaYxSk4Iz8zuFg9nE0CNynP5tcFSekEx+a07kkrl
Mqz72ouuUaDmsDmUbb0mgqWzoN9cKIMyt8v+nLsOUMYxEAWqnapmYNLuXy3J9KfTRqEIy+dl/UmD
oBvK7qRbZ1FWhxfl9vlQJWAn2T9uTcrc/s2u2KKILFwspE2HIWOyEj7e7rnSF4URXINOcS9T1900
DRTK6hjsME/9kL6VyEiNZ05EuAs45AcK6YfEwp22ogo5mqSiSI57lazE92rAqGMRq/FSY2wx7jHR
CY/ABYXZ18KhaOYqLy2rC1Oz32q6bKaVW+WWCdF0nhGiQsojrBO629h8AOaJvSL+RcWAoXNGVBMd
SWwYwMZCFlfz4hmUXXXUn0DfK9NCxf7K12XMF5iGfHs5pMqgRbHauz/VrwCkLW/O/FCZlxujVDae
5yPhNG8maP7EZIID5lSh5TP4zuWi+L42ZJeSmZtEIl9/hn2jIt25OrAiLe6hMN39y9CB90SnkWtY
jJnJE9nL3dFRC8ZD2FW0f2VknkeWUGKx/XH5UQ+y8sxImoULtZexByWLtnQlH3CTOpKR2sUBy0eB
BWshbXaEUA2YA8A3s4qF3jd9d3l1nksvuir4MjhROO9qD/8oR3Omi5LrIFIG+B9I2Wv45VFUEq4h
kSUHkHULB76l5o/2Qbxyr9WMxpPmHDiJOP8gdHRV6z6Of2YdyLRu8HXIYllqX5hGTRwYOL1lWMs6
ZlO4Jvm5Qt6u1zJL2m+7+F02OvOBWNdH1Raf7WSPT+TmZCpb5L3maJGVxhNEIL/iTjkfjQhg2Q4T
ow6JVZwGa/meORfZyZyk5Z73/X951aQ4pfwSxHW1OOtIICjrK+kyVxK+CSK2tWegMtGRi5NVrsaN
7eLlPWIOwfTuL/4box+hQWHn8b3XThf315aOLJ0fK4Ki02HW/Q5Y6g5OH9tzuS/FgrF8ihJ5QlMs
Sp9Osl2g2+fuHdkXIODemMEM4KL0gjSEnPB6RKhJTeJJ6OnxMBdmnYhN58eNPEVLuV3di38OMMdS
V60Ez5ZOcbKCp2m6bfRcQBrE3Ku8crUyBL/1gZpriWW2QUKngESum4bgPO8PvE8Fs4WOROvxsCwM
vN91j4VE4qbYshpPsTbc4I3rBLgLCPjxbgVSP7hG3WcHI8PwW5HEtdH5sH+4NgL3+BM2nj/marFb
crz59zcZQIHz6j8Y81gkTxG/S+drvbb/py8j3qawZpc55NsoAV07m4TSX3gcyblZiLN6gT9FxAWi
8v3YxSdnC0tJs5EYNJ/4E7rGbwn6BtxP+4O0Yw+stqHl/DALaFDaQ7Mez1OCSjtEzy5aMP4l2s16
SB1yQqULAyVdtKhCYeALMh9GLMfKmPvNjzXRIblhkHdt3CQYrSgveCFfyYzcjUH68ymjeSzZgti/
ZlNYUfqy7kXSw7hdizA3IN157uj0RusxxGk3UQKPgWufdiEUxJFOJQZcYaD8PegxvjNkm+6HV7af
Hp7+xOGJZzkrXqIsONscu0/awZaEtP3SrUWfQUaqXD4JruAGw1tSTwUVaSXxgCdhmxO89TWxlF4i
F6RoWb/rkiAoHwp4leuT2Nc1xsHZaC72giAAZ/7aygPEnGRrEMbEBXNTg5k0pV2OOFRInWdY4OuF
jD2w8TPP6fpf+uVrEOry2x1sSlkCa/j/kzp9/LarhfjcJz9gfCB7Rmun00uKcQixgbcvws99oZj3
ukqOH5Odlcp+Oi2RXuudLGSS2oPuxekcMQeNegpVEUW0o2mlUPXBu21m6qfhha9yXBluFzGc8s98
+xttvgv1lo8yhbPvVIb5wlRpWiGlCbkIGaFfnRJ5DWSpA26BPCDr1qxpKsR8QJF5o35Crc60URrn
OBnqQCLetBQYfwiNodHXUy+l1mpW99Q5sGqrrW8pI/dt5cBBpF4EKUu3yf9sodp/cWEMSf0KIdgR
L8h06jnHTsI/e2rjnVqlMNpTNQ5M1iJGpFyaPYsDP8n0gv595ya2osjZDXlSobXwd1gkOB7bGBJb
QpPDCtS5eV9Ln6mqoLZJ9a6RK8uDLKVLK/pnbyAX2K+tUkptymWz6o6WxHLK60CB45vWmyJHdkSC
T25cpyzpd+x5cyfcRNNcX1zHyJwnt3YEt48Tyn/qKbtjRH8lu9Ih9IUNw2tvx0Zj11A8YzotZszc
0/zxsM+KpSG+edMwTTOCXM+m2rB3+e7dTwYlY/HF7qfCanaICSl59RswbWOOmpEO6TmycSt6gJxI
Ak7fVabZVMq/3kXfmMIErjmwsFYWDomGc/AvIy1zTU316TuTLUQx/iOcbzq4PW3f8psa9UDYZI/P
4/afFVpHexVpxaQvIwJX+LhFTSzH6lLtykNJHLfcgSF2Cf8UA60C4793OV22ugI0dEIex9BOy+sc
WR24gVZPzvavgOojCW12Edzt0jsqhdbxtmw+xhndC5qu43EwR0oQeXlV/WW1jWpVRRsEWOrhFAKD
jud2ZqVdfcW9OcMFlXDBHxmJggOH+g7pfkay8s0yZwjHSZnzpVvgPII5qamVRCR3UhGv5D6QVy3o
SAFVj7lIAdZqU2i7abu0mE6BDEV5UL74eA/oQWfWYeiwrm7JwCkrrPfvE2x7u8EQHD9wv0TT5pxY
iU07AGfw61pzJMbxkyUwnlntvUiNae8xp0/5O4jeoS+88GNc973rTzAeRiwLXuCAfiDhwWlGl6Mn
dpwOidBUKKMSx0xfiH/UG0NUceVYHmsdkHzHTnnvfdns2FEKufknQp7b455B4gI+ULNE1Z3DnjOH
HAc7R70WaDdi8nvPMf1G1Rmj24u1niqRY+scJIZkOAka8BpFhsQBTBMb7guLA+VFLF4tw8IyyyOw
hnWTBOEtwR0+mU484gJRxDzX6IgUU7fTFviKe4n5WFA42qpbBAGF5ytn2XVKSXLpDgeyc2xscZmd
x1VrmmdwquUp2mqrBXhLQ99PCU6RDR2f6Nu97WzqVX78BB7LccKqEfJ88cEG7SoNsKwaOFbJL3n/
4WpnmiqBQ+9KdWYVoa1EmltIH+2BFeVpCeuoSThICGnNWOc3zF1W75bOjpdZ/ewYI6ZvYEZJrLIj
i7lOCUSuXhQy3ooHhY8AeOX1wgVWD19g3OV1Lk6w9+R5Oadqeuzncn/Vn8zcfxMdsO3xNfx5waDq
/XCi8wed4xwBDIBjPYGeTUP58QWxUC9XzYZcKLCraIZ+G6+wvrveEaHWIGUjPDyCBQgYMEcj0NmU
/zlmdIVlrCQkLd4huceE0mfeiNPJGf2kw9s4ebWJoyT5OY8MOAJuvMD++8ylbVcNCLj62C70GuKZ
fz6OsCYbHIua2WYk+XwKxBdfcCKc7IUEquLwlLqdEMu4z5iRk/1OBivoUcylAqrEJKqUT2u9zfAc
9EHLHYCnSJigFXphvbJK0TgIcmXxkI4N1YpHYtRQ0zmtofGgxlzcGjuIku2vPPlZAtGLlrwhRsnL
DSnAfzfkbea2JG+NwWrjrqHPlzEAMfneOKVsHPfMPjmkLhLFjwsFQr1CEUqf41zQPuz2R9gPliwm
95IJqnppvJNNQy6zom4b/v4znTrl1FDU8UU9Koo0A7lCJ1M8HnZcsoJGNQiBVRsEMWuuKaQybk+c
nvQOWJtya0nWiWw0pYsZiKAHCadfGt1bonZzc0QUkpXn9flMrI7vLqsgtSNCoTBX0rAc+EjV9Lan
PV8FXy5oiv3PJrBSsIBsBL3FHgJ8J+Q0Lws/Z7azcBELgNaSi28ntoU3CCPzTsRqPIKz4EWSh9rd
FUjjX4qIQXbUTjax8cKub1A4R1ug3yHJ5FquTVecMW3AweW1EFcv6TW2ZPgI2gasWXtm18/FiuDm
6d2l0/yPVKT8SGTqNNJwGOXKa3/R8kFFH4wSy4l6A5Uqc3LpOllDfgRVHXlHxG3fvViibiWww88w
DpIIeA4vv/4jA8mZmKLN19NIF9PUOqj8mqKLnO4fYp2CdlbloL3P6TEAFtBDRS/PIfRm3fkZTgsF
7S+GxWVB+2EtF4rHfL2H9ub3LZ3a1CPlqbwnFNCo1EjBjS7Zx/ccF1N1qjLugjZE0kGyDBIGbj3K
H2bCKjfQYgMHObuzP55l8BG1vuyUEImB2fhIaJfPX3EXjtJj61Jpv5wggu1hlmi7n8W8/6AvmcaF
HgHafFX10YQtP2JTmxFBD2zZ6LfYmWMEtZe0b3PbHIsV0CKgUjfZA34CoxkvUi4DLdRfoGQ/azaI
gk0fLwMY67UOKxWJ6l0SFcbQHNdsCsH2Y6vc89iM8zbDJfsJmcvUBYry9/SzTJdwQkyy6W2roUYS
a019Cu524HJgeTjV9Jga5nmkEnsJeD2GGjI/UKRdGunTWqWvj0aBdWex/RqfL5fQOgDLz5jgClyE
/FI8zuoSVGMVdlD7OkeBaqn2MFU5ii4LO7kAgdODEM+vHLcQvrQnIr5Rr3q/Nu2ONxrm3qkB2ObB
bTQXaI9XP+UnbeEsGoGBOzhKf7hzcR7ZCMgicW7dHGHkv4YIXCKst4sutvvaRFaE6IIf75hgaOag
UpnLGRKUhUHD3NzEbdMpoCFGCpjB19ajNuPKOcGe0B5pUoHh7Babace88Li/su3AJVIKRSnj528W
VOz1XnERoWzzH0ZvZlk/a/3ZznnbXEj7H7Q8+w54EjehS3oSWK33Omuiq5Zk4njIc9wtlUWjD/2x
TnQVGke+EZnaTlVUX4XyYUXME6SMPEFqXnY8WdNp7OCjTOuV97XM46qzoEtVTD2io1b7VUgIRfDw
izSadI4Gl7S4OhNA712z6y7HX4kdUJSdgTbvakqn8OwFBRQd34W9G2GAfyUOATrAU4aU13fM/3T1
x+C2ijU5wfXL31fX4ZOPm2AWAED7Nd///KBLwIrdmqZHA6UFml0abVtlFnF6YwhUQYGaR/8bAmhi
WMy6v57D7ooVrHlXMbnkHmz6/+4Zqnb/IJqgFNjBPk0UkkZzDX+ye+ARGma2iXIXwDBYCSzH9V+1
EUjoYRxZ10YlrIG6/HwrasCa2p8LOqCb1nn1ZvJ5r6/Zj8YsoE2FRSqfuAPknZLA8A2h9c2vxErN
YcX1qx7HFhc9FB7JuMkl+K6MNgtGsOU8apql85C3i6Osax5QVQAqZRg/0EM1tvqZjG54HmFS1AF7
K7gFslPyd3QGGUBijpOd2E4OySMl2Eynry9MbhbFOcDl7OTTaO/zZtJm5cqItLfxuMLL1FsBywMK
wE2fDY9WvrcWpVO8OpGlgIGejGS1ttPJVaPXxUrUIeZ+XItosbLnZFSk4mAsKsaIchvO6z6XrxmY
de7XhhnrFX2O3jHFg2p+UQnST5Dc18Aow39kTVxnOtvs3/1SOhd2DSM0hbI0ty+q37S5ZuEl3tKn
f2NEJFW8aZuuGwtoO0033giszBKOdL9QvXBFJXcMUItc4dldeRP7nqEE/NTl+q5UKReT/eQ/mxt9
Cjw4VzTiMs4Pawf1tnQGKQMuxbVKK+7cRglLFDyDbP64b2pYDEhIgXKpOP7fa/+h5rUlmk+kXloA
kxaA+P8Mu3bBua+2OMjrTd5xiXjP86DtO8IV14hfuagbDLhhsmkLPHDv/LvTHuE6y/wzwjs/Kube
WR7IDq4o6NhCBFnEp/LTbIZuKxoQbnJko/bwDo29dp1NZLpPoE7C/zWcQI/ZMY/0a+eSc7LJtc/A
37L67QXhRBGxz/2Pw/1syopiksGeHcrdREtpuxmYGAfXCibsO6JHuRSkpMDscaZ0q2qMrdMzJNgA
kbAzGVaDRLZNco30mtrKgnwJOS40FULVNh3pRcT4xauVCLd4z4CgRLYOGauraV/XtqVfAl7V5NHs
ngI1EdvTDgiRGoHlxx8XZp1Q+YRq0J0JQLWA4AzTqIcvHALCIMijT9Pl77AGdSUaBGFJBlndKySX
KESOW+oyLQ9s6GHjFOXZMwyHbNW+IwpK7ss/l/nF00PwBVohzDMe6XMouML4fY0AWQoZmIfHDOdY
uotMe/WLnr0oU6RwqeDhEpf2Gu4MXrp27HePfoBad+/lvTr0fWSYOKLXb9ICWRFkgDS+vphQGUw+
Y6H1Y1olQcGbvsaHPYhis9Q0f5GtJ8c2Gdm99bCvRDSoyQgZ/VNHcbtMORuFt1d6qoqMPuvOmPXR
C8OAFGxBYgn+HiB+hXtIe/DKYxsNk3ddbyBSX/DVrWx8O18ybrd9nJTPhZDuVqpx1S2kw8OO945l
Zmoo7TgXztUPY1/d/ENCfIOe3XLWeQYNuWtP4aQfGIKm2auPuKG8+hmvlv62iLxmpjn2Fr86Nacj
ah9gvaktX6kQr0XQoEADYjpr+RDlGKv2lXamb27xF/qo90eprCOqWZyqmYRH1w8HiijUMuJU9hvi
fkvFVA632YTapT5UXvcU3hTzuh7LeyJFQ3i/pN8pudpOio/qMj5rz/7Ruuz/juV62W/pHZLfnp1u
E3CTn+CeZiK4jc/KOmioJDTcrdkolu5+Z1aEDaxhBi4C8H5X7OqRHglGWmEygL0+wzEqa596Qmk9
AcCWSYsCUfgESCcwLkZZlAE3qXMPciuqayEgrkRBpr4UeORU14fmLMM7JtrMuCKaV2hkwhGI5AmO
FPKPm+uFNnOzcUIizQZ4AWDFog0Fx0tj5rKzphhv/q3cdGj5G/rMK7MYy0xbpmLlPHib+ILzEHvj
Bj6LTMLXuGDXPRmDRNru2okkrt3kpu0zW4zJ7g8v3u1mhm2nAo5QH9MV3BxNNDEO8XT+kkkr3Acd
y4k2XYOOsYJbgAVdSrITIDWlYvFama8tyerPJeYzGc9xrsUCwKjH98K4UYLpPxcJIl5Mm/7EgPva
cSkW70jSJUR/tFAdm6yzxhqMG6Sx4FpSjnixCerlR/sm0M2WhfcTsLrQEbDYRGiaY7Dd6V96GV9N
7eOBD2sn7dMPY6k4hZu4a0DIJEhei5S0VXHkBgd5+YBNmh4t4OdbigT3wBoyeKPH0SiIJ8w8FTON
ia7DN1dwHCdmhfe9tweHTIBYdzq+WbZ2SCT+lrEFF/87/PN8ZiWTnF3xino7b5HcWnf2+7O7xIwo
36DEP40N4zn0L4l1jWe87hP1Q88MBLZ0psI33r1mzBR3G5evKDx6pr2BnhF9f21GX1E56hrJC1t4
jIrJW263YGe03Pa5h2gjGDM2ltFHvvWKwaGzRBIuDr0Pfcd0l+SCg1HGNwKHHPRlNmBu5vN8WSYb
mOjqCG6WwdawVAYR8P6YpATpfFn+AhimboZM+G4oGY34Exdi2tj246+gstAWVa6MwaVHHVndgAbx
uCYoZC+sQiBgfrOliJFy5GUprXlwJ5/ttW71pJ4XytGoNZDbwTIGvYjE/0dTKmgosl73O87GAO8t
hV8yOGEcfqCz5QruaeP0LIZy9i7NtReiwhuI/PWHdn176OS2FVA9OoYRD1kqOABAvreoVPb9wf3P
Q9fxBOZfIqDr+7pq/8sJGvMvWRjzx16AoHqE05LuRNCX803GlXmssGEoKEJIcVG1XaCvRKvXHEzb
5jaRkci21VrlkbjYRhRt8n9EyXIS91/Ic9ExcUM3ueVmq1mf5BGv2TW+HCg/WgXk69MmoWSKgEQ9
+00ox5agrarnd9lWoaC2fFUQ2QqVRNxoX6gyWn1B1k3ufgah7HqbjC2vQouE+Y1SKivwtQNneq9q
op1hP7jcuFZMeGbJstm1/7HOuQMajYgXNlIMZYI7nFVHs7BhqrOV8RQzGxvOqM+vQjJOWRg9EkaQ
bGpdSMipM9XIL1bfPjx6XWgxyxqrI98yVBVZP3tHwDP9wtpAF/+c7ahxa97EejcFGno1JfNnquVG
ItArZ2smerUIvrde5FoZBMi9GewUJOBc/iqBmpfBnTUlq8mIw2nhOz+YVAg4YNajpxtlyMfhB/6T
PndrT1a3NP4pyucXFAl69y8LbqA0z06NM+NXGce4InCpWCdsnGjHI8QqR5IqlBIm+38ZDKWvcAMq
AXrRMrQO/H2bAnZ433ISyocCX4c6BDc2UR2x/XyAwFQGi7ZebP0Id3ezYrpaKPHC5DwfJ/9R437e
Mi8g8Np3aHTZEeWglxJYLFwk0OJqoWAVGvvPNYAQ7HJatECwH5hsn94A4dAte2x7Xez1YYrjJck6
yJFFQZCPJNBRRO+m2+VFiunoNkexLJKjsqrKJl2/zkhEq6Tzo32hAVP4DcXXOk7jA3IvBSsIa1ck
rVZGlZ/zbZcsL6CiUq3TGsIs1LECWGxlx1gaNF6A6bCsUutysDjEROPvi7YnWqqs7ybWhFdqGUXl
67Si6AVirVuZRUwLZRT7C+LH+5qekoTIYX1mGJQiv4WbZbjay24fKmO0KTwCD25VCSLAOXNrTpvW
6dVNEBin9sTysm8FXFhgwq8pS0spWYMpRGOeXtadZlx8YDvd1kch5ZPRDkFhD35vlXt09WmFnKth
rLOLsvOBSKfZd9/Di2eTD0PcZEuEQHyz3a3/4rlggpfQn+TzMbcjkEeGeZ97pJ5LrsC1fWOXyLOy
nExfLu0ipiddJ2sLGOu3o4kzkOyGlA3zDnqG3Cg+fiNHT0am8db1sZIhmz6HhZzlBSiuCU2+NRNH
FF2JmQK2dA07AklXon/FQQx16t1AtyyOhZa5duKE0fBTe807FqTrjnRFY0UdjaC8kL3qIK7Z+zhP
xE9Y/gjbPVXMViYe2ZkEGsyrk4OcDi5OMbkLd9ygE4NDqRObkjh2urStL5LIwG0iQdAVQ5u4uxkB
wblVs0wdTX2F5AaynBTYiqHn7Pi4+5jFQ5v3s8uc9Pjw40rorQW/PWGMoZKDmJ5IEQNh4FxA1seE
E0DSmgBEPbNnycFjPscD+1nD+3DwA19KgPF2fn8rmD2EMsA2K/OZ+zz5VW/vg4NDtRLRvAsNqHsh
cIHfQHDyUWXO2SUfA19O8OJdayhBYNn4dk45opzpTDSqtPoDZPETz9+lylEUHpyUsQqkuhO/9adn
Wara2k6Se8PJnHn4InQaajN6FGfwf3Il8/N4pEzfr//MXvi2Y0bvEIqnK9ZLZznj2iha/zN9usnB
ckQR4I/1JFcZdBaqXeBQen41T6IiL8OqCPSVmsBPflZiul72evYAMQGd7Hs9LvjorAkAsPzCXs60
tsGTRb0w8yS2E4ONiQaR9yrkCFly9x2frMqwkaE5i9NK4SNHq1noCOa4dAykXc+iIQTf2YnTcyu1
XrnA4KHKLeED9LZXxjpU1XFGTMkuoGdoQNHw0lvURqJIoip8rAGzGBg6v87FwS9BpIgEXtXmgTcA
sPo1DJPGAkWN3PJSQDX2pp27XXMz1NTC7LemErBsPCi6zcdbZSxWBqGSN02QOBzjboRPFFlAcEX7
DsKtF59+Vw/D+yTY1Skrm3zya0WDuBPFpCff3x3q/pG33LBJwlKVHlxOMo6ks36lnyDgtfFcHr8j
9SoYP+L1fZkOAUP2yM9byeiNB52OufiDRplOwTduCb8iB7ndAw/086y2BVPCRxAKtrZbN/GNyt/X
+0kGkd8wcaHx1IZZtYDfo/RziAdaC0FeDMVGr1v9cQPCQdQWK2CVd3qQPMRtkH/z5FMntmGXaESU
alb59rsVjbK+FolFIdwnTi48/WD84lwi5TEDX/oswJtjLVd/oxP+Q88RrratpMfulJw11Yl/duEb
o3ahOlhUh3tdc0thhjeFQi7mkgqWJUrN5muSY7+M4dyVfmcJsAPSaier4oMF/9TEyFXFNUS2pNY3
kDgSNzrBct1ulVitvQfbaZzjk98qOXn/bYtCK0laoE0M3YS80RGsKuay+wfHjTu2Jo+1nmyGxvko
ltGleIFZRareQXpd6CaanY/GdnIyooiQg2DW7RyC7HxHAbIqikCruZWIFMYt0/ZzIzrJlmVt3zdV
MWezBqRUin4YbfQ+ubmNAn13oJvuAaMcyo99ZYkMzNrVa4juTaGghqNwaF7ErRx2wv6CNSH34i7W
G0O6sREtnp/2RZEBC7se3qrxhVVFOPNxGCjI7QhQy2kPgJLu8rQEP1/0xroOCDDEyOs8goaZPrt2
0Bm047RM60gwnwYlYnaiSwa9peto2anW/8lX8qP4yoEEtuGZuE3m712+B9sZxjo6N2MqDGGSBsKg
TL1UwVuCixsv/JSCH4J9iSs1s5FfWUiH60UrCXGUPcv8r6YNCKHXzy/HuaM0+mN6ZPXU++XYiZkE
6n0q1MK62x4vbei+Oz/dkqxA8B7ANrj4nfjMu520oaa4o+gRcqlslGUVLVtrexKUxC93g16Xiu1I
PbKr74m7nUYh4PFGMiCy/rN/faZvPzxlZ7iXFZPTkX+g2yz3J/3/qhXNtHD+knEZqbR0t4O0HuZy
Pr3pM/DZCGTTo+0qMFbxYljqb0VosJMhqDcsw4k+ehdykYkNVORaz4S+6S+CpVtE+BZOQvygQGmG
VPHxe9Qti01SeV/JU7agNui4C+aUdKynh+L2Ium+hu7tsgNQCli+UDJrZ7To2zY6aCrzapzRpbhp
cn883dNcKdiT6SHaDjbywoSDX3ViMEIpzbV72ZCsJWc+Az1Rjkt2f8jh+erN+PCmioLuVyK7hlUK
wq2C65nvLXVnxWQfrFRu/GCH0MQx642UOQYL/w3pmIInStx1aOik7dD+yccOTxBjmL+I90fuN9/b
DCNxHnKzwFeVR9a7VlEcNG1j6KwiOLmJEfLY+Z5krYYDrLtHaZWktXqAkkkVHyn+vS4tq/b6xPXS
dl4X92VxTLCCyfQfrdeKIN7FtF5TC2lS0XKR6BFgYzk5PCKsZVCFsLSCF3n7+7Bfs803tOLxvjYz
0xWDtvEczF9CcgFyBcSbfiAfmYnZQjsXBsy/woiB1EKvO03yW4V4RCNmfIyOqdUb5KAM0ssTtD2B
bRCSRFXA2Fx9YxkKcIqWwOxUdLjaw7KkD+nz5iN7r30c4iJ9aY/I0+3l4hmsb+4XypDA0pXui9G1
UKIwWxeekfJIvpPbhehWAwF/Vdw6DKvSbEK52VvtBOE+JskRBV65/584+GHhNGO7hnrSW5AnC8ic
fULCnKHjIax+nM83KdJ3hpiywawjkKc7n9AYn9v6fFUoeIdfseJLrGUx0Rf0NFHQpHp48TZlb3NT
Ss8XiexRIE0I5j5iQKB0f489Z2/gie4O09nh4AObN6IS+8mAr9KHU3bcRZe5fYLiIgLz0mw1YpMd
nDFlKamcQezGUFYb1wcVqz0svCmPXGbwxndEUJGWPwS46tCW3iuhYDnwS33dUfkLEDSFgrVcif6T
5UknbCetBqpEIbtfPGUIj9RU55ZnS8Kfc7HjtGjkiLzcwsz98iymA6ndNIfYCEKxM9MlBaoKy7Sz
1qa2DmXvvEVwFlZtM7vgrC5AYf1lxOlOy6kqY2Rls6BhDW+vkQefEKmmNg2xgt72QDcLLhBtG5rd
M/2x5FfOjvvFKfLXcNO2t5cldhccXT8tj13nRnXeCJ5Z2GNLnJJ19IkAwFvZbXAubSWnKsdJuPc6
6X0qbI71GwLqWfjfVvqlTSL8zIwSjS2jxTV0fhMXac912rKp9kUP2bMP33ntzarF/ZITaTmL6ZMx
Nho7/f7YNnBlD4vflUUL84kw339T4s8Xk5mQSEjcK7vDn878LmHbkbLkDYchipBdferQqWEO0/u2
4zlWYSYi/U+AUPt8Gp5ng3Ae5pAQJPIOPX0KsKcnp8zgKPf5IGbniPc9t6JfqGjkrrz1icuwl0K8
M0HXjaQvPB9V0FVuhFcWysc7sUJ5LhmO/O5jYWRliafKWeaAL66xrQPrTmxBz7oVt5UILpD/128+
7GayFAr0RtaraC7Wj6JL5SYIWy1x8uf+s9mzhm0auQ1dGiXyjPfUxxEtyggwxIbXjLgSLsGdfz+7
AWwTbXKGiVg8eELRd3AD5NNMLQ9A6ytSGp9PvseBbBVCnITLrJVxWLrNENl34bEklMc3AYmHuXWB
GJw+08JXcb3zCU/QrNOWIK9Es7Slync5OqJ63ODkdt1p4aLrn4cHp3FUPs/YocisFOMEs3Cbg6Tz
gRPdUH0P+bmIM1RAfFVcbG8ZVoIt9els/O3LVdoANVNDr4vzj1G5NaZ1MEj1iKqJbGREgLjBr5wq
m7yxMGYZYsnBYS+mVs+Rb+ZFCK6Y6N/5pBXWYgG7tMNQh8pHfpJepyvc7WZgydOrJjwgzUp99Fxe
F3ADinIfCtfDjK+16so50Nvoj9BIK/K7xhEBrHhiKIH7Q3m2RurgUWbP/pK8+JEu7i2gTcQ8uqqB
jGNPSUHrgUGnGVLZYLvxrVmDWuOEGwxpjz/4xdjTOyRsly3ruEATRjyKit9uojETOmTS9Zm784Bq
ju9RGxAXuzflMuV9B8UF0IXTRhGt/RZ8WQajbXy+kOFThoGNhYDD97NnPav9ggYg24p3zYuvlecB
0Lgqs2paQ20qArEZCVk33hFluur5VL6B1TE6Q98qTSoNMXyk7oXIAK4usuJ+h0xCPJQBd3uAI4AH
0e4HwBc2zsUYmhX/2QV766l3f9XCm4Ebhja0jdf+2yyA/bbH+JxNstsOlN0tMwUd8y61FSUtSHEu
vRHK6aR8xTZMGgurltLj4Et03pX982eaEcTQ8CWfXwX9rNmOO2xDEhBql6MVH6TxaOJ5r6YhtXXU
9b+5iXj5kfoaedeTiFBn135NMt9JR9YRy+HohK2neFzR6WIw2eSwCP4NO7UPrK5hwl4JvAeoG6yE
LI+LbtNDBGeZ67WNraf1ojMJimhqfPiiB8ZUrGfQbCo26SCSHSNcM4NE9uNr01bq7VFnk9ceGk3U
XViUGiNBj/E/8hMRvnZPTKU/CVwDbqngE7ve7hD21HlRPDZwtP/dQSnPuFaqW1TwGsExWGmXRIcK
f+cRvFP3xckvYnc13hsdTs3py34+f0qoHWDpdwA9B79ZZUFhVqtwM6BfIRb/tU7J7JDVVXga7/la
aDgbffJSijuJhXmWxEn1S14hnrSJDBm8F3h29E9DP+t24v8+pHidX3XFkSpImvmTuEMVuE652SAu
nYe/xH/dki63jY94EW/8Jexz+FQWai7Q5FDfpJjZ3UhhjgBP0dSAgukwECv91Nz3pEeNU9L3irYB
rQUkAkzhC4rk31x7r3f+jJf3sG5S5M3DXpNC7VsTmRvLJb/2CG6LG+aYCOWKXnfNPQptLNJpo45+
BWI1BdTjhA/gV9afE4hh9VpkFl++1o1SjmwCwaGbVh2PPA/mMcmiYXzcpu3ZeMjFrkhX5qLGi+NU
qrimbWa6E64iZKgPGF200rHyaraL9GItuqTy8aMzxGNBWkTk6TyvCyo+E7FTzjUWujJ8YQq+Ct+q
DM33JEUZl5sCQm6pwWpFER4xtjsmHKz4WN1cnfDeWaWDlwMLDWMzgxkKy06kA2nh1YCP0IfigBWM
tk5iB1v9aX4ocnYvwO7xhitXShhWQuO5HKB94q/4RqOImhWoC76qvWkytuZf2wyFWdtx36ZPuAGK
wJ35B8q5gacAKSKnGeWT8ukXdyR/hd/6ZNxkWUsQl2rTOPe5guK8Pvw8AMdzJHQK2yP00o3fWZET
JzVFIjMMQlcOkYhCQM/hfo+4Xu5zWebkw1HrxOFG2KoTykwtrWJQXJ2CBr+QaGgk2Ljx9ndeZpMO
8RzcFRgBYPtFNLvUi944oAmNFKsQOKaLaiv/wdeEdyuLFUGxTMI+KoU74q/sZ2mh2ih7vfst4BD2
ufkbiwJ1uDhNdyVqAgSEGFQQlw8ertQ83EuaFkiTUu9jeJg4kUU3rbGWh7tvTcwzL2tctnjZma7x
dGxa5XfAqWBYzDfDfQQEX1qvl56eRRCtfrhNSGnphvSBEAIhHKE7nryk8Y1yI8oCmG0vDMPeZwM/
L55+AtJC2BILZiOalON1hOVwhNo4E3DyxXk4GoAn0DOmRtd/tVfwr6LXaeA6F9+HDHFCKryQejnc
NxOBRkKk3KqIvyK0axvTyO0Abo2yvDboL3F2NyMZBcxskrDquQ7t8B827RGoOhXKQReGvzHWgAx3
j2dgHyl9oOAskr7Qj21GEHlNNfBwb6KYY8rRBESDfDSTfvbI3Lib+DvzEcNRNSRbNfUHoEdbjQSL
W+QYL1PFDjp1t2p2iJUpV+kMr28B/Mq4csxSFNMNa4Y9Xyj9UYrz3xXZxcTMs2mjs5vCykpgHzr2
O31TMJzNDaYQtyUK2gi/J/hUEzRGSySLWzZ39x6R4j9q7FxiE9niAXkwuY6IJzEHHkWpezauy3co
IhkOHwM+WH96A4vWszYc6P8waVTd+SwqmUQJ4AlMOBGNoNSHe1Y2dfF5Zyven096YhcjaLjKcp2L
FI5IihUgtS8mylgW9TuWJtS/gY9652+PgdXn9IvL4Tivi2pX4ffOzwZeVOvX+CTiInAIO1feYBiR
kRcNnkRgLn7/8lbiUg1CZrfvQRvU75ZHo03z2N+tGoiOMP0RwOwCaL0tYM7GlZKMepQmmAFzcKZX
jPP25rleNkZrGJq/F33oh0Zaz3+mz6Ii3HuqQ84RgHbqqvmC5ksA832hS6SqjF+4+8veCHEudywj
Bp3F44x8J70jYVFU93tt5HtExQ/cAdIGj51abIaQIjimmpulSw39fTocwT3zADsAAxDDRIb5TvEf
3oNPvvVkJMnB56vOtEGrmd3iYHEUCKo0EvFpUlt50x9VcWXWf102O0AGmxCFSpetMAMuuqoIpHeI
cxusInEHt89jXUGxXYfoIRpPwBs+eRARc5NdfwXSAGVYp0pMZEbMAejNfSSxeK6GQBbLpO+sHDxh
hhiSnD8VZKCN02L7TXeyFOffgOkPAl88uxPvo2dMggJobOsFO/8OO1hcORo4H7QcNZq67PDL1bnT
/mKBetFwsLv9qO0DGLdeyDLKWj1BPztapatLYj6ofldpgUXAJciAcagjNzWVAqB3wGxdKQA0kJy0
zyuevqQOdq5sISk5nrs3LLlsQU13QzrNkTAhR2gtdISgZtELUgUkIckaX5Ve6wejO92zw4BrJkOb
aYMOEmpiL+BljHdBuGSta7VbIc36X6naMRbT5em9eABb4BQsWGS53MNuCiWvmhsBKXoUQKGaCSJ8
wNoygEq/5mYgVnC9SGxtbiQpJRLCfiK37Uz9XSEX4tWjMRZMo25RHWVCsWz5bqxgYWeD+BrEcZzc
a3oUEzIVZq4ltOn7F8a8QPdH7/LIR1tuwnvF071dnjJwiO75XGeuJ9nW/Zdl8GWFNgxHVtHjMVYj
LMFknrAyS+YKIVOsjnyDQ7oUZYycQFtyvZNCP6zY24p6EAfjzHL5H70iuupvjOhEB+O2tCFXyTFz
iJHSh7IgbDKV3Ja5ZEeNZJUHB241QuAaBmlStuDXPBOiKbzZf2hX2DzWfbtkNAtKRS5VWns+2D4s
X1bj1UcfM8K+LU6q1xoINmgBjGb6ucGlWzjHf/p6iCInDIDMHjd8XuPq2dBwTatOGbPPjRqodJDR
7DLGSfDEJaj2kMimw6UGHOLbzocJ1encM+Gwu1R8Wul0hSdb7HmKBQDwHqi2fTrGPJPhjnPf4uNa
JGtneGPdDjVDxoXWOVnB3VdQrwhg3KXcYV4lLtX1LZDTgtkhxxpgQ1BEdtZ9rDe5hUgSMo0m/Z9m
eOi3g3gV1naDjAVKkc/eiUw7daRrgYyRJj+yFnVRdWdS9e9xanyWPJD/t8tFjdZ2ZrL/aCHODDpl
UhoUvRGflQjIwfeVEFYBhkieh683XmIMce3reFeA8kn+oeOVbJhax6Hgvtw4n3YHTqhELtEBJenN
XemDpEgodrLKrycnPMpGC+dTBqOB0rhiHKASFyO2M1Z04J0SWyRIflD/PfiVC4+T+kUdby4bdRGr
s6UMQ8tsUzNVANTkXrubU7JIuVUExpBH7JGLzx1Y6R2XzgmEBqORrDxIsxl+W8lEJ9DSh9GYYxM6
ys6t3CJwyH1HOtcttm2UEi2xSoAcQKUirtQEJUKEOIrWLZb/vkxpF6z4MAGT0Kj8mnWVBej58R9Y
6cwFmcAZ/naMbavqKpvgFMQy960pAZT/q9SjCHViyeJ67N2R5j8TnqSzn2QPIN2Ihdil89Ch7cRY
PnZ+zjtDDFyHR9d62z/NGvGp+w9j9Hx7s8YdFvjQ3KZq90EXIXiyoldkQycBpksh9ixUl76mxsEH
qp89fCNebqBj2Kp2w2NrDdjZvvjBG4ob4KTBb7XwVSoZHMQbKzQCRs+C8WslFrmC38ok3O7KVrTe
N1jcIsvZSKfjY1OyFmsttfFttmPT4gmZEvZQGE2aXLbwK7e4PFXJp6NN22PBaESuHH5X87GbhDKi
8bAA/hBH7fezGckiMmlftpiubzBH3CY7N0471uOS28gQ+y7hsRiUutYaBxNYDk93bRIkG80G1f/l
3CYm6IKFXVQfsbbbE/iR/kr17P6x8vH3n+4oR6h2h6jkZXqESjgroeFB2iNCqCXyMViNFZ5Rthbk
4zkntngA8x2dXewzfH2vLUts6e5ep/jLE7Ph8OVeIJmaMHsaOakK8AvbysLGGi9oSCsnNj9z0nj/
Oz/bMWzjndqDO9j/QRtxdXZaWZjkTczJ2owYBXunppTMmmNZ7UMY2B4KcMGsJGe8kt+1IHxXgzUB
EdYO1AQsUgAx02UXNIbtBXRJr3GXPSjH+1uENvLrjIoZn8OCIY17UXIpL8/qVf75tJPLg7yakV2O
3nEfUkGTI1sE2lCZY82IkpvEpgQZ7jb4Iu/1tWo6EEn2Q1YZDzPqC3b1QliYBUbSWRslHmVv8KUr
XVJITRO75wcMqL9yCmh75PNFo9gcXTw07YWYMCbvWaf17GyAduIN9bSq5hDNNHpAed3K977xeA0m
O0eBQcPHKRRhdUJZDXTDdXO6b7F1cPSTHOeIz/5NiYT2khAXuII66GWonb8QQSuhiwtbBE0P4X/j
Kl6s2QFe4JX2j9pAl5IA/1uzjf1FLpg0kw2oyB5LjE24S8tvvSj8gqyHi/6fLFGudxuUk4QAmHRf
u2RzrANC33obxtya7deVNfdHenUPMULCkJiHru93rxSVreQe1uwUp1ZsazgjS/aaXPgwexDbsYyi
gml6BboRlVZ/123vK+Kaihjnimgn3NrgmG9Oz0iRbUWlGKjy5U1eEZ4ilA6ddCliOKRhYpEm3epY
fnQxVk36TJHGWDfogiZWprMGNHHeT2fKNGv0+7/fFJ9EGgeVOMJpS0UE4X1oYRKliDzq/J69fPTh
wEvU+2s2oaQ8sNzEyvVVJEb71jH4V3d7Se+qVRCUzEOlvo2o+GTB9wcIT1nFJRrnfKQipq3Zal2U
vUKyzJQ5xUlRcC65YD70OgoH5XtuttkihKHfgoReBrelPltVa7weDFlj6Dq1y6Ke4hSl+uQzAJLB
T47kp+zjnz++S0YOhjryTb7Cj+2Ntzx9xN9Fp/4/Ktb09HiprfqJoGsIkIkhbK7HHGD/Z+yHhjVY
v3tPxiB3Ftzvb0XkcwBrqYFjy//wybLEkQBRmFehLdUVIC6+h8rmUw2tOX2m3eCSVT/oCo9OUnIa
JTKXQK0h7RvWXMMI6XY8jHnL3Z4HIb6sTriaF5eHzoZnoX540DrpDLUeW1PCNIqmTQwCP+AP/mmW
iP1erqXWdcA5joAeuOez037kMcd3eCGG76yI2LUU1V/VnycW8mNDRURsku9E7dB6H5G5Ns3IgrVq
2zqeNbo56U0PrJ0ISwXTIGmYkpBVNQ+BeBq40OY8wW/G3u7NyWwQq5SfBgzcG1bxm1dh9sqjslqq
C18UiAC4jsyqlEWWvOkzy02oYdplNeFqnl701o00SahxK6iGx12BV5Yr81W/L4Tvy6MNaJ1DAYZr
gcdean7XGZ87H5DRemrpBd8XUgUM9Sltyrz3zQBSzcx1KomudhrX/oVJenqUcr4TcFlRx4fxfyQP
nFj0n9bh6sWzPEIgTYT/hVrB1zKAirRlAh76UPHXwosRAh3KB3u1mvH0ADh7uBQleKmdKd+57Oeg
a1XiMqPjxsmmiRlIzJhCWWKgSUs4lKPSlZr7rscH/o4Zn8FFzUTnB8FvlFtQ15xxmp2tKhCsh87B
kM3u6MnAOsTYFxoVukgkYZg4nYghzwMMPfRysvdPpEe7qiO5aq7JGAk/tAVMtkId/ggnCaAGKifI
JI6GRdywKPCQGyf1oIU8AK5dFLMB8w7jjoQAP5o9JxicnsVxCl9Z+X8Kk2gn2DhMExjqF2FVWCMx
6kp2CneFuD3R/f6lL4cnTXvr7jf7WViBU6K1IlJnkD+U5CH0RQinJv67MwEIzd81/ybF1NKLr3Zi
MGYhTQy6CUS2//d6v6HWiyFfX6xSEll92A+iGUDsTc/zkHzoyI+ZwwowPVjsy8iIQqJyGhC4Yogm
9gRvwkCYhHRzNRpwD13GMh4ZnQ2zN+qrxRv6+kYj5aW4gTkj+uBoQYyud0ydWBdk0KhLwN857+8A
j3EAKaE/yyO2ODocIG/QG8qnilJzVXY9SqDCTA6S6VjXGd58cwiGXqIINS8dxrInKwoHwuct3vOf
cO23gHO6mUfqTlBU9fmMlB6i6JGAcztosXGkhH8K8lhXoW7AKzAwjNMhwrqmS4ms02T/2ZsJ/BdY
Ie2jFAqArgStq+S7ibkHDlUOSbTwqCxpU+/2cbzDfCqUZyIA/whRiJqswBNlmFfEv79r5AZC/Zsd
eW7tJoxuTElAwiNq7xKKudWDIYG7s0+aN9W6cf+Fj5Z2jAUU/tw/YPbWFui6kSk+6mpgytvyyz8U
Tn7BazNUBvCCYBjiLISQHuTa33OnnbuwmhB1Dbfr/ABYwBmsT0Nzfzu8lNYoDPgd5zaI9ElpqHCs
i42UArnzfl/zxxqFA6cMlFyRiTFON3MVi6AlfnDod1wgkXEUEGoAxuXetnaNu+uSw7lMqBmu9vFf
SiY6pupMMqyptpMB/GrsNr85cblsMKMDhPtjU4JXmPGW8ZXXQQJF3tu89rKtST3y1Z2lDwsxUwaS
+vbNodh/eR8B0VodZLKPwL/zGYw9naLPgT6NEaK9/fZ0vYFB0C6PHKe9huB20hW2TDBJVSuqjJTp
nKQvGBgABmvfy5T+zVfxEELfFpuPM81nZceMuaVGLHYqoQnGCsPWqbPdo+KtwygX7ntlwXA03+cc
kUl6hEJdzEdG6e8HZB2g+AuUANScpVNUbRmaHslj68k8+/THL2Hb8FjQW8wf1b/Y558NRZapDwcw
hvUBnSX632v1Ww01VYk712nW+vMhl/AKGYypayy/NFTJv6PdgYom8tqLATUDIU90ux7DCimTn3FS
KxcTY2sJguHRBOZm7c1DV18qV8VL9Unqkm/pMRtXNmGoijV1wMGlSe6yvOk57OJF7olE6wjskMas
RrKzM/y8Oyqnw1Ja6suapCx/Pywa2qMZZqCJxMkSw+URNuRXd4WCgLvgBvl6APMmQRpyfeA8BklN
V4xDOkGVTJU+YI0Vve8JOq0JZ4TgvoRv786QCiauLwVo/oeO2mOZ3dGO9A6qi+Z9fCe5ZLbOp+c7
vg0jMtr32J+KBIr1gA/cZSmgX1MXZ8m4phLgvVGwPssoKev5L9/hTmomrTevV/fxnnUndK7uxKZH
jdf5mrmVcjhPuANc+1rijPPKyGjGA7g5lLPy3tWwPMkfqH5U2bycy2wSSuhRuX6CdFx7DSN5zepW
c7zKz7vr6GVgkj2Gun7cGQCBavLmhLPOkQ7QZAKgZTJNNNx6QfIAJKRw+yp2B7LwkSnF8oPv8OAi
XlYIAQWxh4gCcmvJuaCwA474KzWLuGtu5+VuzrvzMBR7xLSNUcL1wSMwdRHEUArwwB+xrgCtjsYw
nwK6Wcyri+wJs3Tw8craN9JgmzFUZfUeywoRtn3cArYtUYcKj+qWcYoEnd0pVVKMmrkmEs0su+9K
YecJiyPJAA2aXUT3SS8Hx8DQUOjH67b7LLsOIvPFpLDKYBwXiSJZhK4cvGyrjSDTi9GGzLQy8irf
dfa6gl7xbiP5qN5fRgHLYIUBKoWIM95NEz4ioLINAruGCJoNBbdAypdI/qZgVWpdNcEiCXJxgZau
gNknUgLWjmM2ZC5OEedvITvb5CW0haZa4UmHEGCJdHDHg0sgZrrRhQfNux3InJSutamS+X0+ubHW
zT9lp4UpJK52/JQW0UYevDnh8TBqzxaj4rzph+ZQkzmxCStu4ySqTNN3qNZlBSZjxp7N2boHvd3S
vvkQpqvbEThTBTL0lx49nXGoemo822QtWV1tJs16gSNOALcXQWcwncw/RS6AryYnbvaTwosKGjhN
6lm0SDHMaoNDee/o4fxJfyBR4jfZco7wIfkIo1qIw48JRYY4MzI52qZYVROBDXMTcqDaCwjMyRny
c9eZTclxSTthSGamwn2n9i0I66wNBnIV/lloQqRh2y07b5nVsjkxSuMY6QEca5QSiDnYNqGyrdHM
eWG7Hn9IoYOK6FKgNncFSSlDndfzI0/WsJcfMkpZW5QMaswlwk5NxOr83FLq81bI2VQw6Kc6s6YA
D/PNj5KjUpVgdzNvouW2JKUzi4Vs0QZxFeS2XYvVdZhc62plvJ2rdfeA3Rxn6s0sYVjUmyNHvOUu
gjNmMnY46lV2BwWR4V/vwCvPXeEl9ZZkQwzPegu1AEAWCyNSMNvLMWGPSgQ5ReWIlvDdCMOKj/C/
VuV6Z1c8T2nLyXapgn3Vx808V1+eT0dQnS6fWHsmd1YtDSdKi8RO0qUeLEsVA5fix739IcSoW78p
EUNSp2S299Fl8rwdno3QWVFw8n/gQEHxaUEt+0lruMvOJ2beXSKrAwwSw1ZFemVyVl9+QX/Ct02B
rGmGvQ72OFjSX2pbTGqbdo8tnAmSW4gyUHMhU7YoGh0XClgPH2gFf9xcjhy2/VtuKwnR8O+3IvlJ
KmgbdypH02kBpnhck9D0sazmNPliz9X3gamxw+ddUKYiHgKnuQuyJkrT+Gi+l6Mo0yyerSMRhO36
AkAbAwRnOn+Vf692+IuZq2x2Y/l6BDtYFwT4h9lAxUqBkA2ARAWhR7h3wXM3XHwHA8XNyAMdpSFa
g5Up1lO+SEqDO68g5htf9EHynoY6RDlQYVoaR4xvkxHWo8kPJ4kpBZSUxKo3D6nckAok2K1fpSqK
LfbSKYhTS+lOqCVGVumEuaYSBFgCmcACVpNniBQThrqHcrrf3NMXqQJ6wk5k83MEf355dr9s+/+4
kMUbvwlOX+YZMX1DOIf0MYjIHzy+QtYt3o37R+cJsaue7fXy+w7LrQe3L/dsp053J16MiL0BL/ma
wtN1v0jjHA+iWA/Xh0o38V9HfScupeeWEeeQ4yGiz63fb89LyQC50L5QgKeM3M02klg/vFtlAlrQ
u73CBmS4pDGfdneGEryyQpi8yMyxqIeZ5kbQe8MaT/ltotWFhQSwKnLWkWAqtjvilXIVzKK1HdL1
rntzliaPNZe6NmE9zgsf18yFYXSPpcXQgel2v+OmW/2t2IB4nQGyORhGfy7yLp9xbYbjPfciIPcU
cMhgAC+iFQ6Mq5lBwIhxZRrTIrqq3jRcHj3kTeejc36dYzUb7hZyNUFXryoU0fTIgAK0FwBZSED/
N9QVpjklhLqsCNBIz6y7EKPFn9TSUaubffNRqMvVEED/PsLex9M6dwWk3V5Dj7iYO+iUL6Z34fkz
cKh84n28AA6wjbPMsvEJyYSe1rO3CGLOipoSpa2BeyzeZyEEFBCnVeoj71o6xlnuLVTN27fqTKNx
8TYIo/JGSo2cRQUvnoUXRBmygRplqutsk3Qvl5iHFAejmC34G0a/R3uiQp4Hqc1wa245yUcB/iKC
gjCR0d+j0P/g4XBMNB/RkksvpmCerB0cFve2FQliz2TkruH68BtNO1Stk2Ji/1tGu97dyVk43I6U
pXV3XEm4Wva9e0qTPMwIHwpTaY0aQFF5rPn0gv4QmiWqn0MdHp/KdPVjSMI/b26VJShvKJEJafKN
6NbU8lqizbMwyxGLkO1jJHXQ6pDsyUrwKdBeiXyFgTuNFJwjxxB66XzSq6Lgif3vGj0ZsCQuaz8Y
PD2Dn+pNygSMVpYOxS69GXKdf8kOq6H7d1YWHpjqZdErLgWejDa9ZmmPxCe/uXfIEBNMtcv/5M4k
7zJisTZ0Hz4oVqC4GgSp3+mW0onTIpoD8phbEe2yAY/d31KM5toZsY4YcLn00n5SZqb9c8NATebG
91c5Hg0ckAqj2jJtLFIZs+fIF5XsyCSona0qkARVyM/G4WgXDwt4ZQEgzLLFjVmGfmFEzrGn+P3+
jgBpbDjMoVy3A/hpnaPvXqvnMRtZOK9qM0MZB3zsOuc4Ruj8x6BTHxeUbti5jEu2kdXq86T6yCNB
rHdkTuRAJYwJXYzAV+Euiw1jvK0OSDwvB7cePOh+cRLX17rhf3c2Z+TcKG3AWu6E6uAx5tylHij6
L3KOlsYapUhnTCE0VNoiKQm3ajDVzzEdWT+POuO3PMxNOvujpo5MEs3c2R15wMlmM7waY/G0kedc
GMJugWgiFfJ2bxP06oB55BDAa5ucZkv5QyOmIdGA9ZCi8fvK0WlitfZ6psgNOuOyXbDIV/4bE0fJ
hu0AdiOz7Zp0EPmWmMQ0eG+fgnJTqJX8PVxfLcD9agzusJPlKu9WS+f39MNngPmnL6Zu2aQsl0dH
4N7hjbidd1VBQD/SOVlg/bm5kBjpErapxQFmub/5LMLQsGv4/mCte0ys3sgAlNGHtv+CvaiIQ/Oj
Lna2+CnpRfnz8R6k09g47fNO+IpzJeyH0hNZKChEvr1gW2thyHzZGvJ5MSfqvGAszfAw9unVYIJW
eGKt9CwO7xWVResC347bmCmeC3jdJe78gQkz5SHyNhbTNlgCBGvVz+gxf9YQr8GsDNc26uzAOHXh
kI113sGyNMSj/+orIfhz69h716TLgqjC21vNBIT7GvRw2lKM9nJ9JT+EbvOyw3PNBNo5LYiBkDj1
QakA1UauyI+HHeaFbUjIzMfOKCdn7kJCt/UWx5Cwokyp3HlLg1YA0HAUV9UaQ7H9lnEhU+39w/XA
r2N7C26jrsBSmE4DgX/rHTc4Ged5w4jlGPvFe6w0JvqR2JTDgQkHkeq3P+vfNrguliSH+Du1w2cA
6Xt22dOvak5BnWFtfi85c2lO4Y7inFHwEg0hXdHpPzAGt7PRLOwnQUJOJA82BmlUNGaV5Wos2B9l
l7sYnQ7RyOfFZnE4S2M/gMYzFuOHQ96pCm808PZ7EdDq6fTYhemBTmZC0GN0UlZpLcjS5Y/+gx8b
EFu9d+8DmsF1ZBiNYsUiOgjJpjwn9IdKbYCf6FFumMNmBxWxj3mSBzNjm20RgltQCibuEj+XJYLO
7zGYGOwciLhHPmtyibU6juGgxzSo5qVMMrhGnKgACn73NBKMT+mJpUSvzTxjY3mhz0lbReiymarY
LB++B+LEuux6GFOooBAqu1hBumC+DjRZt8FR4GegZFFM2hspDoxdB4w9C/uQgEpfXPyoPG7CL/IB
Lwcr3K5qXtLJpxrejpcx1lRrUmWMcxJCS2LySXb7XUXbxBV5m+JHjx4hHk/efydfjxG5qeKJek5v
9AOZwEPbnYOfxBu73k5CQY8jiFGcZ9eQcfoaNmGi9PxMjtFp9Mx6edf0eBh+XxZ16IhvThmHdSLZ
cYNPIQQVDLAUpAtivl7kEYbNxPsSJ0XhcVEnqHezoe8OcDCeb4yjKudqCY44i38vGN4gnwLoCdzf
LBIv92tn7liKvxsv0TzzeLErz1MNun2PTb7FFYRPD02CLGnXRee6+jtyKZQIWdsbdrierMTFYlsv
kxi417s0FyoctnutuGJifBPtbZn4G19NKV0fhautGCU5MM2nPnyUpwIHM91ogeEhsvmd9Zk7hGfE
xark9RCEtiD+uZVL8ANxON0liEvzVELrKqr4N1Bkkz3mzu9T5miT819TLVC/a2mr/W6f85P8/cf6
yZrQa60FVu6qP+nV7t1lqx2UdEgOyqTGL+inqpB94lrd/fZYYoN3BEdFo0SlY9VcpeLiqLxd90Jl
EYJbxtffjCryNsUGEIgDa7FqGva8XIs3UQzlifiIHt/kifCrvPf1FGFBnNmaTtEqhC3sVJiuSpmQ
gL8kEowOrUoEWmxwdu75OfmmGih33jOwmWBVvwYG2COjueFD8G4Kuouo90jQ7019sF7mSVbfxghs
laLb6X/gAOwKHhgwPvJtoSv3Q5wi8dJM40HffeDVqkedG+3Ua16EEOJeO+TvsROHXTyMET1Vm65L
CwynjTXIxg61Nx1on3bHt+1VmXJXZvhs9Sx51xvXUJHDTY/tZMPhzA2EXB7/RW+6KcHlIMISuQhU
f/tLeYUGFIlm+03HqxBxd5r+rme5Lg6k+NZxTqcfw91gUcMYwFOOdIx5JLv69LMZ2hNk4IZ9NSzB
4MAW+bpHMAFpRgz9rT0B+9NaOPYte0MEECMhrRrioB6GlENrcaXnCPvSvRKoy2my7aJjDv2MHNhe
l5ova0zcdTviVNL7j1WnD3+m7ETlC06t2+GthuW2EgbTQsIv+tr52IgCdiHtlxM3DyTacqEEim0f
b9+f4e9RMS8EBvtwcBA4qZ7np8UTpviH5mC/VfP4z53Dp2TknOk26bSKzbGaVIUXXVkvfBUHYRbF
Dboej1XtGTiRstcRcH2rLLwnU3HfxOFoW8KSOgZTMH7k4w8VBX8hottsmCFdkQu49eZS5IPhwDaL
YNCllDijZEd2EbwWlnFl4UQxUznE1KhlszDFdhSXSz5WZN3SRIibD+EjwFG6pv4z4nbPp/2M0/hr
E8naLfEasU5yASGhoWJWtij3tADvnTbqNDwDz2/5ROQKgq6V9vfmNtuqEL6txVdJxiDYdy7K0E81
o42RWyJ1OgYNEIKDhWXr7yu+I3mEPrn5k8OkyhxAdWw6ffQtolXzPjGpsqnnB+klVN454plccts5
/JLzgVpfz3hmYsdhdm2X6QyzXtqEgaGiSca7PVRJetkIW9xPvBX2ziJmEiw7f33gPHJI14gHiN3L
vlTjYQxTQWoA7Ecsbfq0x2aWyxrDCuJHCG6i6q3YRpjkdgfMG+ghNQIaBlRQc5HZ+VHvNk8YFZVD
7DgJ2zg0UlTFq7ajqYY49kKxpDKzMdaBZRFCNZxHdtHN9cjzXiKRGu9Jn2I7hc/YjlcswqzGDXAY
OWX2M26WgHOLNWUbuTJqjnLWqVpwfWd0PZn4/GPcv0czHR6gkfAAl4YXxltioyumqJhSwnq7UTnd
0jUh2wBsWnIDEMmsLvsrmx57s+XW/kB3Fik+tNxMZFxEZV2j4glsxGnP9ioXHwc4mXtcj9uLAWHM
3BtXIAW+Cjz31UcQIIyX0QzOWj2QI0tRDfW6R9Y51tm+W0Yj/sdKDXwpHnlzdgpcDKgHos4l7cyr
NLD+e+Rzp2vqN7pkSFB790R5Z1mirOKueQmuqElE9oJxxVsdwmjL8cmOBsM7y3HQOa/ZBMoGoz+/
TGbb2WISwlmTcO8iyeCPkofXc9wGMMYF0jF6LiCWvHJE9emekN5G8cNXkYOkVYj9VWla/5pzWSYW
a9wr3bQOIlDMJCGskQtgJMR8GCEXeF+RLm87tlo7OFDpW6y0CSRcBmSQrdvkEKE7245wbI4R0/tB
kTSbUZmS78epz5CPV0DH6/j92QFNrmw+j8VDxiOVhnnZZ3zvtzaZg6ci1inJY2/aUFNNlo5g9POB
nD5R2x55rAlJ9Mkv2J32dRr8vAg6RTw/1iJk01jR6m3X9/dyh2ANXbO7eYpGbgOpsOu1dpcjg/Q1
nTpDWT0uF7cGjV0roSVr28DwbIFKpMItBEytY/AaGfFZRu6+XQRqPOPn9mQVEpy5h3R5SnYCq7FW
Zi837Rc5C29naxtSZiPCyvVrfyTx1jRKoubu8ycHI+Sw01RZXwMn1pRzebaKJ22ULwxA1jX/8ulK
5x6CbQh6OqBkrHuvA6FbCUPGMKrd9mYsJaWvmmQ9qtRQt7UgoBxUYSFvniUIBVjGw/LUowPzraoy
mKMZbELcqp1M85TMQwET9B3kAGwZ1iVaOfU95J0NU7Eseg19yZG1Xl8GutieGVvzh38CREbTEofK
lOJ/Fo0UrCe5XXB2M0EdHOdlKnt7Z/GqIoqesStwwK+zzoCJJVnqsbVy/b6Tvj/rKq/PNaNE1kAt
HLRHYajXV0Y701GDJoZ7CPn4jpNgCykGfJHJmPKGyqBQUHoAxTESdENBLOv/qi86SZThz7/+Zocn
0lLp0D6OHBU3aI4q5llMCXk+QnMzdbd1N8ZQNvERjfHKb3g8/vr/K4ax/CvdyzWBYKFYDIfhkebf
IiDYqkbAvT1XhjKN/d/LI4LLXFK93XJCfoQ67lwp9YOcXWUxEGJVNF+Tx+XnJB7SzAW1E0bsr6hp
XzfBrjw9bmgUw/iEfRXYMEWad/Zb5Jo2ZVadvoO3NChCZZr0NkGwUW2DWLAi2X8g2y4L8p98wi3y
vNTPQTApOWVB0I+L54GaOWr9WzeifReJApb2xmLE+/qO8I9qMkG5ph9oHhj/5RGJU6DGwn2yHD6k
B65c5/x78YO8LK0+efCh6EdScoXEKtrKLrVwpgw75MpJcpVgHhkI4zGwPvyfSlNr6C2kTHpF5pwh
mwWD3szjwF7/URuaCFrW48XGEaiIPEruNvvZDu1Z9k3OghAbNT2bpD6U4/jpO81h7SXqUVqfqalR
pVUp9JuPzK17su2fVex7uXuGZGX/Jx6S8trrRbYaMJBI0+gj5d2J200x3u0Ss1SjUFN98pfQRuYf
KS1Or8xlroi5vnP27R3Jt69LR8qUBt10+0p+la0A03lGwB4IPm/YZbleoyjbsAvk4wqsT6l0cNCY
QaHUEDcrDEzg75MznA22qF/kbDXzlafr6vzJ0qcrxW3aUzCgHvR7S4LQKotjKFmFBldx2rgwAkbZ
YKQ6O96n3D/OyuhqWUytSlGZe4R+5Jo7xr+R+RHxu8F4XePuAeyV51tzbv65rNkohoOML6Rd8iae
uc4vpz6RJndadjC656864eZcVD2kPIGGvphhAC+q/tmPiI03N1dXQTM5edjVFf1Xsx/xPcC2KRpO
qjDpRVDyZ3GngvJnvsSnAU85kuL93sG+1fdSp/Mf9GMumeYOQyZE26DP2WtQ6bvdz3ffKQVjh1f3
Mk7I44GTwcCo7sGFV6lNF23dQtrpXxVUoSZt0jlLzXIywEpSG4etw0g/6tRq73oS3A3cn5ah4JV0
L0j6WSK1rU4rEKK7L7yVNgvoGQXDemf94Z909gb+YrNos8s9Bx0oOOACrXy5U+4KD4nSjbk8Gh4H
VBSgCa6cEdk08z2KPsW6MAJAtKo/SymGSar8IGZBAqEBcPcU1eYNK29DjCkqUsT7qAdgzclR2GTs
o8QCQqYKW7K5GyESL2prDs0lRTrnDCHgGaiJ45oLfCcrWlVMw6sVlaVzCTfNUZ7Gd3qdT099NxRg
tWxRomkXayJWyKE/C8sNUxcxD4F4mjVIXdbCaTAlK5W6stFQ5pqgDfb10sI/rhqIfmR5I1sqD1jS
xqyYA/bfG5hZpteGq6KQnQhiypC+cH/fJ7O+xExwok8LTHSBQBeBx8X/2NrfX0NXPoYjcXRlfZ0z
XRRNe0FjXN+Rw2nmR+qrgFXm9D1ELV5dOpjI2NImDErTHf/5qgXXX2h3IfVpX3wZmNCvLDbOmccT
uheU1GbnOq/dq+x05aGih56ONCFEWhAU2s355UzY+ZlsEkXWbOlhnIw203FIk5BFUamiZ17jspGQ
whm0TNuFzfV9MfCGRrQDudoqESAjqLA+ac6C/yc+n5cyzNfdxq9btLAfPKHnR9k331Z5V3VLESQM
ZRsdqjtdahXqKXeGyoocrKvPqVzSU7Qo81dj31j7+T4cMPFYXDzNKUJWw/QTSV7ccHBdnLTePh31
3LTaqFPcWOwWELgf6K/5GiUJCGMwBkLz/5i3t4I5kwZeg6OlTp5nzjfhc/BRwgOsYdflRN6Wjdox
8bo3pGldS4wprq1T6eJBpa2rcTZwjgXLN1MQj7VvfGCV9Ml7ldKd3Btp3Usxk9h6mfUSj/iYoXUw
2YvhyzP27DM6v35tLlUQGBKpSOmeDYMOTM+xVqOdB7vyI/VpcsnlppBJqWiKhsmNiw1PczKt2qQ6
5OcTYrFNPpWu3qGYUnYl0BIBl2UJWylC1JkzDMYmO4wisrPkNcHC4P72qKd5OWSQ1lKW+QlIa13F
7QBqfp0AzBZeNgGdxi8Vhqd8Z4zH0D8wCzUtS5lCxrMLx3BfoJI6ncwqY9rHG3KIsOZY8yk07MVI
oz1hIb0I+7LjyBaKzkUdG0zCfkVxKU/ZnhbgpiYS762m3UfhcVkmEjs78CY369P1NQX5jPgvCCZm
o1plk9rIobQogzal5LXus/Zy7zItBl5+zAq5MsLh6ri+Du9mo9M3G/xRpU3SQT4+vocU9ybwqujV
+aMTsLc76QTGjrn3RQflniQBDlc4ugvW3tvp61de3fpy3ibEydLdUCpqF/xnm+BN/+aO0VWcMCzN
WZlh0RvCA6YYeMfdYDmwR12+0RZAF526BKHGDlN+cf5S0NdrCRvAnWbqep9qcVDnKphYm0rJXIT2
U2mwX1VspEH9swSFs/timni/gxR96bU8Tin3Yq7ibaxs6lq8TwKXsEdTUkItHgPUaMlHUoC3P1NI
GSy/It1HFb8dlj8BdtDixN0SH/Rw32XaLDCH5DgCFTsRQIbXK2PY3W8kjMleXqQ49sEQNFG7Vmn4
2Ow9Zeh37pbpaqTsVESXIc3LTPlbgCpiKD2EBHQkj+L+BoOrDO+LbU4zrmAJCvZwiaT4q4GyA/R1
Ut2+UpYkxw9xfji9XNKuBbYSbtfdGf99SEE0oh03Ot+lyBY1LpaGrkAULbSVTsbkkcLtyATc8kbk
bpywHCrTT8cgTwcoIxktt7lJtDP7NHkrCx+1hQuF8l6Oy+kMuhVHN4azkBt6RwybsqV85bNMUiHh
55RLN50uAklh19u4JglK24/A5pdrie6s7ME6xAOBYijQqmUWL/XE/6Hm1Ba3SyPyM+U9ikSU39N0
5DWPI6qsYOEKMSTKl5ytUKgE0509Tjb+avE+QhZwQSfymSi9NzJZBjzawvsltkk55CwlkahsjC+N
AOQfXIoXbr1c0PHU8i/9eFK+k6u/hakPaJz2UkoMTt43CotClxHNiIXRuvhzk3lxfqrPZxuLesQE
esnSaomGRz+PgKCyxgB9TDZqy5TnLPAzuPeIXpGiyywU5fPX9SY41xuRM/VGmgogYTxeAxYh1cub
KC202dsGRI9/N41Q7H62JOBJxs9yUdtxQes79LTbn5GVEwnHyLfwCzEsnr9irPNj3mUFkSP5a73X
enV6Fuyu+E8XlOpLsgf+3hVPy8mvFDK/Glaa3LAPYAZVXabKosj49nxC/Clt9JDT8sv7vFMdsh2P
b5HJ1Y/vGtNCFrPjTmSYVgXVxHsVD6K3GcFQip3PtM4Bv112vbWJZOLwADvf3ZYGZOOklssi5j+d
14H1CVxZ//SjZ4saOLTO2XUF0rCciuOnR013BDvzw62U2wbkCfEELs9gZ8+ixTU1gHCVbTXM0GjU
iGmlJZ/Y9IeN4G1QvGymP1ebdCC5qQDKgKIFF9KxcupcqObwF8BrXt85+UaXGw5/0vANSbqmbCoh
M185LRDqjBSfPVA/yvncM/CG6eatMaWTW8CaludOirMJNWge3DFxDAMCAguYRkhrxjncimIP4CnY
occxSocQw/RXSOeqpYLEl7nm6Z7I4sBNqZaj94KuGd25eDJb5cwXprGZtggDgfxtKrik8kYwavGQ
xsxALGbC3vXA2/+U4ahlqEzDOT0P8ifIZ9+XMzx2rhVMjnucCHi8Yxde0gXq1yHSlaWzsX+RIo+a
EO/EIX6IeKzZCZLcVvlesaXrQcEc9kVQK/xELl50wj7mYZy99gEye8qeZ5CxfmBODsuC0sttgZRk
17Ok4/CI/L4GI5dLvaVq4lRxR/b30QJeeWOjzCPFC8uttHf7TKoJpBT/ZxzbaHFoqHkPoEnPGVPk
Ji8W/4dab7/WIwyh+kAQYotyrCYQ4sXSH6IEf9g0t8Ch+fWGbzJXUTbo0F+0XtVXUaQFxsOHk9Q0
EkSGWnsF1z7AC7GC1pAlGtAEN3mykInSKmTYPm1O5P1ZPBTYzkhSUu+6XMG3gwnloUDKdiBExsgV
n36WoqR7z5X8Z3CvKGy4critfHGj2w2gbh5YDTQgPhHCAkB6ozpPKffLqXntIFHKzv0/wbYNUGmz
M3LhvAoRvfpZpbCYxy7WdPYtB2sWGaDtrfgTkws/F44ar1JTSgBZsKOh7CPScUE+dh8xG/cIxZSu
Ru843RaYN+W0K33sU+LnMyTqemdbS3s5uQn8LA6VhLPqnuCPYu/U8PWnNhr1keiZ+FDwPwDJQXNi
dgGYU4wIOwqavx+dCtRCxapTyf943PZnCZha0pAfbL9G0YYSbqx6g+x15BdmbmrfntJpHF2d2XEI
s6VuznxgY+1fed3hP4/N7aHMk8x7UcuWEJ4ljoONVQ+PPT/xZpZ9ZF4ipP9WRz2uHiUvptOy/RNk
gCjurex3se7RE4+KAeNazMXsA/YuVzPBa65KgKhVU03bt5O3vBTxqdCygHZJtIicJZujuZKmtuT6
gRVnqXF8kTUUXCjVKywJegntjp45FnzI51Z9fHLOzLOJC+X/99MUcYN3miD58xCcIoZKGTi7VO3s
dW/rjXN6Na2FG7EhLK7pFX6gKujpzCKUTt13Wy0WGIFRE1DUJ+erwIpm6sLC2/F6cvfXXHirUP8G
TBbEZdvVRtF8PbrEndMw8DpLKDw065MOsKAZD2XGovjG2uyymS/n6DecyGY4PAC2pxpnete9wFyh
sKRcDj4Fa3tKhcEg2xeX5+XKchr07PRgFxpfStlcQckxnWzuR4r1otKexe58A4VZHNeZSihQj6c0
AzBiBmO+pboapikswdRrS41kQAElL2bExiTxpbus5Zf0SAENL5oNIUN8Ya8sYQhr5oVa3WT7em8N
hrfLb3VTowmZK2/jqpIJ8o0/ht70KqGffnVvxCPIIpV2YUIElE64E7wvmbDEAbUF2B4nCtnisDor
e7ynEiwBMjkeAmsTDPXwO7J1W4lzvyhgq/GEvOfoWo7TL50z6Ny2loyrCtTgTPWj68v3EpoTcREV
fZjyhZ+SPHBrz+PmhdfZG14yXKoiH3KB6yyA1rc0xSYwydQ9va3G79b4ZpXhnc8Bn1kezAUA3+nv
/FxpcwjxDrVvSIVCOkT+v4RbTZ1bEk9sPC6Jzf+WIvus8Rc9IjF5m5euUKSdAeWgOJIlzp42VDly
tXx4PaWz1chniFxoFFEuRA8rzfeQff6ZobbgfyHjgFxa+cP0IXg4WVtO/1Knj4ODHZZj575B3Y6Z
hZw41rnmBmiYrBzSqOS95Mjh9UI2lVNCcmfVmFkmVQ319XLg8jhiUTXRSp3ju2q8eN1zhKLjJ5kw
kBXNsGZRezss97P5yaGki5yynZhxxpEhfZOXWrSxExvg1/Ec3B4WC4HmzxNiqdp3fpY1AuyNLfdR
8gzLZJltkPMyx4fS515wXVSZoVKVvS+5R4fEojxeF+6Cmrq+V3Uog9L8MZmaw6/8akH/Wis04RF2
qHMwYvBvpYQGXFWpxV9HDPzqzZ6uwkKlPKTf96ltdgscqlOzslgW3jQrN5wgpv9qaubpQlLd08wX
ioCQR5MG9wFR1hutcMliUFRyiwJ8B6ed2bSyrtJZsprdSQRmd90fCExCCSnyCmBApIdwX/ET/EMI
nkfuJrd6P45+Y+cID1NldWVd0KtCLcV+razwhl5JgpZ1cXFjlERzUjYDZ55LYQhMGcHXo20zGdZU
VyW4BE+oHiuDn0CcVxdUoDF1/KsVErNfOsjeblER0mAHQBXL7E3psEkKbj/PGjFLqjQldy66pGPm
O5iFngaqIz/w14Yvm6bigw3izol0jDME+zqyTjXQyYAMJGZPvbYnCHFc8e3KtsDyj2b+HTYTrRzB
rSGUUDCI4zcCI0hUsoiLmRzZnXNMz5sNrwBq1dGO2EUi7tb2VTlmRmZEVbsUGwm2KufMVWuPVual
J/8bo5Cktd3M8HC8nS0/dBSke94wiXLcCH47TxaKwwIqDRCBjA9/oCXDHUimShLnTZQHiaHC6nV9
I9T6XWuIzx+VZL8QW0U1GQeQI+b7skzQBeIc+M3wsrfp0RHjpYxgpvd++KOJmfSfoBG72NM+HjWw
lOSzYwOC3XQkXFc/8RxJK2/mRMWzOyiRjasswo7lX9ys4piZaisOgOp5pjKuB18KZgMb1+QF+QpA
J/ScbbeyGXHqkFpC5TRzEemVCq+MqWc4vu9kAqwlsh5BdHsrnNIH02B9+s7z8qN1TomnjuEN5Kv+
3lGfD6UTntg0jD0VZTP/HI2GZPJBYWVotwpoxevjkQKhzbp8YU+B652jHI2adCE7CAq4CcbN0fX1
Xj5yyW00thfwJ1LlIKPdszjzDkzNn7Vm0veoJuqG7lGUJ0b9r/XOpt2z8RJ6mUDzohW3daC2qhio
SyKFJ02dIk5ZJf/dXxdsLts0VQcmAhH5KLw+OQsZI82VZA3mUOVS0l7G0YOFjatN0V6TzJPi6Tv+
a8tPrVoDjg6uOm+P7fhxjB+NtSWSBJcaVdjg8PmKLnkJOfSnp90Q3izYCsloks9/4MFHQzexSgyS
goOdV0gGKRz8ANYPcbsp4ubKscD/Hra7awcPa9iVjHqMr874aSoL9o+gSwIJfT9OhhudeBdMyn6d
1ofUsy+9Iw+hZwg45w/kyWtq+mIj1PFC7FJvFls18JwtWNNORv0yZh2INJerufRyBiRHFslQV4VY
g4b3PjFfvAdml/PTQIQO5/4ZYGqP0ph3h7voXrCB24eiamSy3b/SuNbOVGePAaUXAwR2q/W1mli5
hJQWFj/im8hAs4OAUURdIgEnNa0LewV5F5KQTIeR41FH1LmGG7dXQ2PJU8a94GPO2nGOYOkohuIK
4ZhHquFmTZWNj3s75/jejZkdCbRvI5Xf0GmLx2TuQXh+HLD0Cb85SvEf2NzeqiENha4Gx5qqrRe1
t8ejEQRJ8bgxnfsAJF2dzOaUQGPeJBqfl7+TPhhhj4KlnLMZt+ELpgWUP3A3YWK+w1AeNPB/r0yD
VOA60NUyo2kBOM0ZnykZyK91Y4tMZks8A9RJ6LrzQAurVRSuNd6Du58ReU3RTHrRhD5zdgIyj0BL
bqAUNsqE42d2o5wKqwSJ2Z7t9cCiC2FOl82zJezlIRYZhnjaVKBV/gCH5Q5SzPHcqJzf+xqWioiL
32pbTJ8ut7dp4Jo9yOs28KermDhfFSzZ+mwMywOSJXoBleyNDhykMVp5xU7t4WnTDykyvtEgpY1G
Id3ZrO1/Xtsty/0YyeBTenU7h66PYZMepsgfyJ1LciQupfdQo13i5shu/5yXBgvD9m7QhMWHOGZX
i3ayz78JrTtuVdSpgi3NgOrIfhk0k3FgLbFPbvLbgYwj3Lo=
`protect end_protected

