

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HpfjZK6WG7sYhkvMgAngy3z+9zzwD77820wau9oTTb6dakSkVNELcmI1vCDbEcS/48D2LFxL/qT8
BNFOIZ2d3w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VPnG2AZhAX4ivH+F+USmM4TuIe2lYrNUq3Xx5puxPaV5guza4OeVGJP6pYRxsBYzj3S4OGH7b6n8
K0l2LCX8eil1TGx7VbJh+Wd7uUD2r86y3rluWkRdWUlHXjFOxoCZGO3zP09eR4IRsG+JxbSDSiqj
FoMAGfR2zks5CEu7dtk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1IQ6dlJ53C6R12Hzl/XoBaoEA3n6gOO0fxU9jZJvCev68EW7XPnj0pNHAKpShucryAUuc2FQgbE
BwIwQ+0yjh3dOW/yrG6sHXOI8NvAIzuE1LMkRT00JCNCjyt9JL0PrhVhWC3cY50b1mAkSZBVfMWL
G4c5aMtB6wF50NpvOm20Ptquu8OAMlN0E+mHAN8qvWTR+CwIDUV/kvH/83yRaRonCOBULUP7XzwI
uAjFnciSf/F9eC2blbPxLHlWXLQDQaZnUw7NGNc2Ufyh7lsh0GoZzefU/JIhthv3ktn09r568XNe
kk/w7iRo/w4FLMicA3dbzrMyZkiVt8z4I74KAw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
x5ctSMYno/7jD9HwXtHguBvqXjqGDToxuRubQZySJLeTm3iuHlQTdlRRlvw3jNvFx8WWN4nEmWap
sLwuJFUESklgDZc8wPsu9plvibxKvIUprit+FQWsTY564IYlM9a003tG4rrtM7zZ9yfolbWe2MY7
qJFpoVf6XAxMMDrPtP0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JhbANRgOr9SOBKZDRGJGrZPWNKSEG3awknWUR+2QiYueCqJ0p8+Oq42E9W+XtOMQqS7h6dt4lJzf
s2rJvfuxWWYMk0rVRoGeqNzUfiVHbjHTaPdjhGKzIm4Kgu/QJ5ooRwBflBurdW1+74PtPtKpfjcs
79ijwPcRU18IbRTlWf2wzAlLDLkDUewye6if9pFfqGP8EVIxQIb2A7LmwWnM+VpfHc6KRQhcdZbj
LsxdBzKwdjN9Cdt40472gpQEnBtaoqRMW+4LW5rSmhm7vTXSum0cU3Afl+AWq9hUcVWPcrWeYdm+
aNrNDk+A5wRHt64iDTF82GsVuvkYpCi38y+ffQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12144)
`protect data_block
VbYVE3NXG2i8gRTZIzIYw6DiPUDovJOMs9jTilufP1x/wliCoFjasnv7cA9e1zhlBSFUEDuABEw2
3vfSumfhjJYmddHaX+R2atVW1CGfv220aymmWvW9LgHg3x+ScfXn9D0xuB0SX/Kt4ukqzoReuMmz
xrV8TBaaaQYmckc0IM1hHyirK0zBPSrmPleZQq7AJ229JeHdsbhWeZaJ3uKywMLWeQayysAxNtU6
83za7G7P5cH9YkguMdC6JGZ77wEC9zoMbS5D66R6nnaY11vjFcD2z3FAB+ORZZhhYEZhD/NGQ4k5
Jz8Hd6cO7AVAC55BDMYn47NjWKkRvMnIlIr4gRgWS9PwID9NynkJaF1V7KBT23L+Mn3YYibw/scB
dbPgOF+VJgnwunRVevoX9gFPgqjltFgMpeRlGMgy4+627C9Qk3CYLgmgG/iBgcyAqvW23AFSBz7x
AI3rliUW8A87zpeiv0poql1bg65KOoDKlfSDRhDmXKoHgXXg2dKzUDWoIIrFb53npiACuvd/YL/N
vqPaQUuzDZSyl8S7iumMDbpSxyIKIem8QK8LUDivVT69FjJU/hw7mtTAJ/bib8Wum1RpmRAXIodT
X0u9fYnOXZuSDYiUbs8qBdz7SK21xUas/ltcdV9Er5MhsSVWpYMMasgPdPiIKV6NtMymQo4FsHEH
nHyft2/Ceeulgof7BMiyI0Nktm0rdn+A3n2muw4JDdlXzHBODXEV5da4FUNd9ZGKDu4+kC4BfnFv
xxP4tZAZiPY+p2+P8MzigWaqGGWDvVjbRDrli/cHYEnbUKewwSGopll7pWcEtYuZzCAPEPEQkv4s
oAZp68Zzv/FEe6A7zUWvZ7r+aC6RnIK2mm94vVMC8IPdx2eRB7czicuXcteXTZWuct4po0Eqishy
yDWeiAK33ZsU3Y7k1laaqtYaIBb2ga5giUkLFt+nxiAOfg0GlTYrgt+uWDfI5G74wl7k0yW3jUXE
kxDEoGOy23ih4lOJnF+CDLR0EXDGPh55FJe3avKE2GY1WZd3G7c1TPfvtvE9eBH3sBBfrXtfZGpA
1EUNzBcJqhi9g/4J1Tz2PeAiZMcQEH2h1MNaEqaNv7Y8lT7WIPpjNTS809t7qvMhc5TClFLu/jX6
a6WQ9JV8W4Eta7XtA/dxu70VW3+WcFrxWDRLxupL3DoNT15ymSmJr0o18l9wKwuL26DNLnfHuv5J
mlq3QLizqdEgY0tfrEInY6bpxW7hXHuti9MI6/B9eZTze/wDZcwnHOHPyS4SCNaLV9TbJI0+YJIQ
s1jLAa153BRtc3A+CvXO07qEq86G2imIbcQgmfXzzJ60DLrBzewrjFO0Q6YB1iXl6cRbmKhlQcYE
BMnVGkFAntdWhCD3121eAJHgS3xASa7ltpcqLfyJzQOu0g6IoHeQOyHhVQ2VwlHigYQqP+W+G0ZL
iW8lcZ/rkXZ+AR6tNM1QwzFW0p+yYbXpj5XRdFkT+fzF0XAc0d36C648ugSY8gtF9XEYSzWuztBq
5EQXM/Sn1CFaiM7Vb/aMtZ84HNsNDhcxHn2tJZugsc/6SNYjSLo3Ol0kthN3dbQyw7lIsMRVafDO
LjuvhK9CTBU+RaOVwiDGrtuhG8T4y/G884MJCqyCRPJ39+K3H0DY4hKDioAJnwlfmfQZHleyZ2Ij
2JfZWGH6snIAusg4QwacrhcJFaaK1+HFafTRbQGcuZP2d6LOrEMr1ftlPkcpujOR0nT1SrvvwRUT
Uc9I1usYXWhuyFb2n4HKTyV7uOTKCv0LlJu2Z0N7OnaOUDh/5Kc9QcPPbIpAJiey0cO3m8aHrcvx
Y5HurynQaVXPKCjSdJUeymeYGBXGP3NCrNoshLSiBQfdMcs9//C0atX69+vqW7NN6q6uNwO/UOA8
GpWfoO+bheIdbC5PfQ6JcakuxKLZXGHcGObEIMEBLdr3V6RDAHI2IXWE1L9MA+PfGbxIy/ZDaC7j
/898kALrjwO9w3seAxXqWU0MqHMCZvNy3uME7l2g+LuRSNx/EG6e/zfn66edHDpEx0Vv0UtVyLa7
zJN/8Q9nHpIDLtVhQ9OKdDlUdZAreAKWXayUpawspJFLTpIXLhIfBUJXAuL4pTeRNubd0E9YQpb3
pulwNl7nhst/8rAJBfeTnVy3d4eTzOStxS/3Lns+LAK7J8t1Yo1coDsqwdCubBLa8rntQ3OEBZML
h8orB524RwxPl76s66dtqTahGVO0aZSfzPGlA0dyDKEIO2GexaMXAXh5NA1TItmBHXdMczJVFRod
5Ul/Y0ZOE4Il1cWLT6Je+X9AN/9CDdYRqNXbCCCb1fkmLlrPrJY4xEZB71ECNk6kcQCh2+Wak93A
lo1oR+iM3iqmJsLX5F/5sBsU4wTz/77YJgAtrRB7OvRS4OkJ07p4b+mN08rLsL3QvDibkg4HaU0L
DSlx+YNY4Rk3e1nGNLVDmnfyGPWCxqV2ze+th+7lifAsOV245o+q8JNJScDrPYJz+8BtoJ/IC7Zd
oRHdrRdsvfx3r31aL8IcU/9qg+gaYVK6GYumhdpVMGv5kiREzMIt+mpjH5rs7idJRmM2mMIYMqQk
0nil/DpSbXAN+LDUh7UG+fNTv4aTb/h155P/pSQl0v0yfq6k5+76+jAvOhuD8LWpSvwLUwSS25e8
raJt4JH25gIJZnVJYoIPmF2o3bk+blrCulr/Seox3KCKcsh38UnIR5eD5eVAhTMneeEJDc7nyHmM
4m32ntLYl42xX+7+4r9Abxmg6VKZKR+R7VlYXIzOkLtnshrMvMqTLDKoolaIA9RV6c/PggyeDCcr
BnXvN9bOl7BpAo9d53CSgpfPBa6lumXb0m4XHnBj84JepTRcNrR0IZakuOFTyf8WI8b03uIe6Hu6
p5ruoroiu5PXou/QylZMJPDZkXDWZxMWpFYZyGWdbUBeLqqsiUTDY/s2vjDclTnfRmtJ42FdayOK
kl/8SHet/aNvM1uCdMxCL98fT5inYiDnYnEvvD+xA8acFCj1pYClbEY7Z7rhF2gWRl/oxsrD0BQr
I12l2mbxrgPszu3DU991MXzwqEjoHdg6W2s/YZbQmEtvJpAfP1C6FXjchcv4GKSx/C/CGWdtI0u4
TBnmlblSmfvKyxwCVx//A+CEZ8J52fe8kaf+IaqEmk+9qaHDCjRP49Mev9OrKsPYcJo0mtdCIhb8
t+vD5ceL5P0hgCtd3FTKkfISzjYWDY72IN8rm4AVizP98BeMg5EhlSam1puMbOhX3cXIGj+8NNIJ
WhydDKnERAH/dnXf4FhNOo8x57hICSIbUK/brrDiMK7DRCNUaOIOrg7wp7ukgtLAuW3DqpCrkVYE
Nig4AbadWGbQR3hkLyFsgEk443l9/j6vdt4hmJykQjVVPNYbsew+TKe02AUUycOGhh6ILEtk/ZJU
UadMf8qMrGMKGXVf+3sS9ojRfUcqOZXXIAvm0/HBQHOn67QxFdC/6FCJNmOk7PoCMTNnzWzJELhO
jgTh6h8mXDUwKHosrGZuoK0ExfE9MVdO+n5YI89yjfNC26G8rpE/pLBYDWlrc8CwGmsoE0Hav9Jb
FHqj5h1zf7bWbDjDlGfea4uVOaedpak6pARYqzLdtKnlCRW83qiDPOTvJRRGcZyrEiCC2aah/jOi
/I/XDxBgcdkYHgWhipvEowykWZIISPykXRvk/oVqrZrh4BGIE2AdSjFvbD90l/+3rWBe4g3KrLpT
Qcb2CVjWCbydmJ4sm4u/0+gVK2SU843XueIwTMif9H+bv43CrJVx5qm4Tgzvc1yqYNoUAeNXvWQ5
0lJLVhgzwXhZKowYIpyMKaoKVHu5vIm5zDC4SyldpCvm8doCLKrxr0HZSRD+4jySa9sv0HYUkTfm
I2+g+ZugSKAj6wNqv+ec/POCTBxlbkkA7XDqqNB39yJ8KhsvUn4yMU53ZEEvsK0isVl6KAd25A6q
XFbPfjclZLtObj1FUIkmwHtURTT9CgsEfC6ANIccWb5+txZVANgnZDprzPtbhSMDqAFk49WG6vu0
3ZhbP5k0i8KuOHYHbmPB9g7mJnxWYrqyed/jAygnMFw9s7mhUR/O1vjYrufjyIN+Rxre+leBv21z
L964vY1j2NCy+5LEKXzuF86hru3rL90vMqyxpg+Z12JSS/KzmD3wPOEB95VZsEKBO0qYDUdfflJV
9NtBw7sJJ8N1tbDkRKVIQqtuZPRT89I6oY+eF+AzyEYHC4xyZigDW0EPcvBu4fwssRw38IAe36Tj
M/sYhoQudALCrugfuL4T4CPu3spzULHs8PxsNbeYa6k1AMNcdKhrACBzJcfYMfInmHZAG5Aq5Tgg
FIMGuIDB0Oh+yo3/55W6PnnGj9MoWlBCDyue5AXTq4OEjTWzFoHGw9xQZpaXWJrFzkXWNH5xfSEt
PR3UH+0oT/Ge1rQ/4AMyWCCHIjrOj3H2KUHmKEkIuubvyC6QxC6NjvpowKg87Dh4Ib6XODNGd4p7
UX4Jt6+lvWwoDGB0vxjBwl1qfEE4qnq93BW5UK+xSpT3/rIcFkIQ3JPVlc0CX9gx52q8ZLUjWemw
8GRhRxtDLMlgkO5CXr5lV5geWPIBfErGRszEMsA+fhoA7Ez4WV1sHD6Es99AwDJc/QZJcSWMVIkU
KUojXR5yfqgaJ9Is2+2GRHwZnwxjyLUQO1CcBMFwbQLgX1bcYZuwNt5MChFxKnUvMTiW88py/M2n
dsYk0y9QHFMVH7ioL0unUpGsp1cgWmceYl4bHepnpHxbPMoQSc5yYpkcy6oA9GixVht4erT6935F
tuD/TrnQVgXvzLrB9vXMYTON9YSJ0KUeEyrJub1UpDDewB/4TYrnHGOuYlY3QQHmxy7FZhjl4uVq
X0HXnH1NR4ptrU24qp/eO37ucWq6GI/Vx/MRmINHG9Fyb5i2kJGMRNAaf1VThEXIWpcJxOdmfmWl
dU6EuWTrJmfMb33ORSXfRq5EENTyKbkijHAOLAgRn8AytRDXCyAXYqAwa5ugszI3cU9flqH0HvU3
AQnnVfPaOz95soj+MhCttjEKTFPex9ONSlRJ8DNDWfeKlLiAjWefF2zUPYpGU2xzSq1aiMmfEgKU
94QeCAvwN/pJG9Yzmj49dN2tZQ3yDBFT6YY0dcZfe9nJxh4s8Ry3FoKKN/y6tuwVKy58HXGZ5tlE
3D3/hvlEoQGJNwEye+DgJDDyW7NpSUrgoBgWdf3xI7aI5JIfUpyITkaIrAjYLqUBTmmRSijZexRT
a0Pg0jlWf4FCfqz6whUJYFpWkdROhaXB1DDcwEwx3uGVWBdA/RQPXR4zS1mU8Kh/y63UNI3F4Xse
Hb7rltZnBBuPtgBgcufuAWEFr24j/GNk6mdz9tJ8O9UnUtr4FWAJ0DEFHPjHRxFXiFpi6xjO9/LJ
Ff2iH8NEz+CJtP5cI+kn+L4dglFEkjDAIsf4jlWUsHLZ2WVe2/bgZnnwFNOnHa1kH9FmlYrvAFxm
g/KiUKqRqRoDlfqTFe3dJoKT7BLDZBqd0lYvBZT1Y4h2HDrT1CrD0/xKa7+bD0mwivcndfK9ioYh
7DksaqrGQ1BdF5JIpCSFu8xJlzvcwRkyueidXhW7ZtWqotMOnSA9JgnpvpzhZDKIgvC01SVXppzz
fadTnZ6ibu6fiNc1bKoB9grrFy7Bb3IddtH2DpHfnyXzxpyB7c7aBKeVialsNLdDSnFms2dzz55D
eYw135EBJaFxKqO3ycTj0zHBDez2Uw7iUjdHnTnoRsozYX2ZRjgwViBShkKETERf2MeSTWGFX2bF
CN2JKADIsDL4Dq6JBJ+jFRYmOTBAl9HjJ42DrmqscjPIPK7P2Icrzp92fJg9QPwsWe2UsexgjWk1
nKtfnOu79NoL5hI9k4tfEI+3QFSNpFqYtuw4jj8mKgdR5cVG7ia+ljKLhU0CD7U7w1PzTRkdJBqd
Xp11ka0qvU+txoz8zwhS4LaOCu77pc/WkAhxu1HYZIiq8RgNDgXpfkFUMOdo2+WFnYxcoQegBUDr
c3IhSWf8xlEOrRaPV8kYPNMh74ENLUgbmPEsGLglTArutavYDQKthzvVqmnV8O1JCxxNvWHVPJoR
bRK2mvZtOYXETVJvvQdJIAF27Cy1Hfu1k5YpRSpNgONLaYwMK45fhYwCQXNDWAEtqcMvCshV94HN
AzzuvzoTkeIBY2XdpQX6PpO7DO+DjweGCzlnkpIfwLZQQdn7GnEF7/9qdd2RK8JSCduJI2uSYjkj
5LTSiYKf6cJ3JTgQ0AmKIHSwaGhPFZE6paiubyetS26Sbg587Ta9XDARRyoVZojt5rsAGbnvrEt+
4FmteYgYOcA2hqIGyr0C1/DRQ2YaPIXnQ4/TuAPSgCuLlQolO3Cgab64KiYCHZarhyIZGYDL4EqS
ItxpqhEIGfR+gVjlTCU46MDqk5YvRmb+XQY5G3Ywe0bdZR5hGMZh2vlHpOeVJjOKLRMdH3FnFh6H
Teo9V8nVblwfnWgW+NNYOy/Vw2X20JedWxWZgxR0wgQnzedCGNwAlxX7rBvmwx4IhJo7NFp8BeMr
XSP1DfH5AXBXepn5HMbsHFEjKC4g0Pl1/X/u2AJKa/1BgIq0OMQ+89fqhZUDMdAh4RZPmgvqWVM5
wMkY9b95Cl4YJRp65ZIsOI0gRoUCaoMzBFSautpd6AhaKhZDizlsC525fArgy4MMMlLuCufv/wxg
q5VOjfMtLolRgAaYUmD95zN4aCpHZTIYZSynhlsUCV1utgY1cxeghvX2nC0Wkfs4m7YCKO083R6I
qjfpO/bKnyxKYG3LeF11L7a6iZGE3fVmX2zTdICt94OP0BwKpBcQ10jPAGNzdLPXUB/ndAiVVMbt
8L/6IRZEFmmRw+oaXlQOhpSsIp42oVZcxtje2/SFOS5PF/I1hzuFB79bhcpqU9UwqyQ0M46rBIdf
dPUXTZliQ6pOJL2Gcnaor5Y9ggBTgUawOa/puY8d6Y06DzkDvboP1VJ/sxaxM61mVa4PkKClcOB4
45jU208xv5guc0cGs3l43PNErqtgcEGoyqGuks/4NqGZLPL6c63Tk9wN7skcwvb4evkC5bOCiMGA
5RsH/t7zAy9e8YUmyZN/DcWaQ0PrAb48DpFDOpUmy8Nt3hbjVCpAW9mJ3KwBGgU6iUwSAArJJdfw
MfaLXwH/Nz/dut8Pqck9AEs4l17lAfyGbIrQ8gD/44gW5UM3Q5mdp/WZ4HURUSfRk9uikVChh589
suBpoZE8bw0qHD9L83JVEGGgJfAu1UfGyzCdHxZIpQZcSUN943tLfPguL3k0kDqnvPg3kBmStxYQ
5BSdtS+QyJ/Ns4Q1DaqT4vxXu/otv1e8ZdczXe5r+7UTdxxWWiPNB9cPETIQAG+m4Oy7KwRRoeds
mllcEDsmILahhI7+eOEtUYuZldGq4aGtBl3O5oOwyJzoIP5+W2YjFYR1Gd19+KbuJLzVidfCgYqn
xNI6a/hixR2tkavnP7S2oj+TFqsaZ/R8NV9KBpFFr4kR9AsA9Bulnw+OZYL07WWk9S/nADxy8Bp2
L/wqyvD5dOhijWDtjBq9kQSlr5d0KtL/2OQUonMXqsSnfSFHOma8bGfZ+qogGRfiswomDdaNRN3Q
g2gMBGgDsDrKaRT5aJ8Cav6Kc8YhvZsYtW4gAZUg/mJrpWOrkbtaIFOZcCeQ1g5yExTkSj0YAbBL
abUcnKqnZss9/kBgjl7MNAPNOJFJtWDePtwvAyIFcCudnaC26oxoHcU+slMo4PA3I46vpQl3N8w6
sZWkm6qPZFLODyjGyBcMeLJ0BP8akHUsVn1b+9LmKicGIZ57l4DyrnJdocGezBlSJWKb67iG6Gjx
rz2ElqMGj4ggKFEG4OaNs8k7i9SOGdmQLUU1PkMdjVDxNIvW0hHep8s8jyjQW865hV8a63wofmUb
A7EAtHYjdpOeo22mSMjcL1XqbfiiJBq8ofXgbxOirEN22a30Mgn5N09GVRcc14WxagmSfCj5utYS
TA03N8mfoVc6oGG+KlcVv9eWSvcKb2GhZLQuBeyxgcHHkoPAnm7b/pWvLg6wqeLI5rMAFGaqQVsU
glVUobS/ck88lYif4Oh7J8pjayRGo1hmkoP8vDZqfXo1xIAqKfj+Q60dlpyzWzGcpgGHZZhr2XeN
c45qvzpwXFoGy6dvsyrU0IO1rMc/EHPlSMWlssdrVyIUr6nAjD+ZiDOzxoGNcuwQBKJ7tC6MyYz1
dB1vaVSSdTqyyKMIa4rewOQH+vt2AedNPttc4EqThQTseH72p+A9J2YkmQCymGg7zm68hwza4788
NWAUI30Cc+urNOY9ANndXhWMnzgWHpwOtrOcIpyqeFG3NXraEjIRJohHYy/KSa401aHVAvep8w7Q
tYENjrzFBOp0iEEe2O6LuNr2hgflYLYnuERaxGOC+5hoqXnccpCe6w17Z3hKdEEboyn5F8r0ujb3
I/gXpyL8bLZngG47NS8mpyi+DODxOvhjLuQOn4G4Jap75LMwbWADzILG6SEb0bk5gW5qMw1pDARA
rZpua17n6yvYBeVJLFPP6aSTU+SUR8jVWFf1Zg6yKOdzMP2fdmBPLQMrbOpqwYV5e0wUjgxsMGSt
iVfXwJroWVs5C+Bup3+pmddJ+AyJXv/P4iAQ4RbFeX1XrESBAJl+fJk11iyeS6Y9JyzhNDOSOUv5
tmpaaFna8TN7CFoRR8JxbnvV0cB2batvFIG5O4ukUvaJJtHdpQnoF7Avjg261CdTtPNXdJRxpw9s
q6Labb90cC4A7NNlMpF7WV2ZwnWyJAHPWlYeqU4jWOifdk8D0xocj+J5I78UUrpocB4cY2uKtzTm
pwcPlevI/liqmmzDdzdDjhO7AiSWAb01iGaW1ItrGOW5tz4yw1ThBKqZWINCBZXgXqpFZIFgZSw2
tciDf+UDFV2ZO3oOCPd310o5UUXhd5NEoePUyrrgFGuueJZ6VF0eEydaaeRwInbtugHE5BfwVik6
UhoT6tOLJp7KplEBdSqaNTG98Hmbcb8xEYfzb/lgQYZb8BYEsqxP3VxzyKCX2wu7GZICPOjWStzG
reFF3gVnCJgwb3baVWqS14L6u7Hd8KEGZ+DNvNM0ryRzqN6D+DSMklZ9y40o9AlnWiwPUe8ljq3w
OiqnQRvP4bcZUoIySEBHiRqcZJ6ZLJp1JERB19nFZHkstTEebN44Fs8T96nuooifHomDvXaZX0oc
pWUKiPbsx6fUEV5Fc+owZKuS9ferPzjNj9I9bcxmq5AjylfuAbA39XBC1qVpveNune3JZvrdIbse
A/5xIBtAOeAioB4tKgdHy0KkJQzWqG/RN6KaOuWKfBUTugvwQtdCBMb4SirNa8Yo7V8ezCy3RfVz
YibtusPTYfyxmuI7YupkXywdssywIzOkt5Ax4HgroLcpKq7UAG3/G3h91DCDzB1obd8DT0pklu1g
yqgRtqe4wAD7d7tWp8druH97E/DrfGIe4DVzlhtk0s3RqH5NDeD1XwT3jf0+L4GqUCjp8RtaZcR/
+7OV/xS0z2ttv7BvBRrk9l+pAcJkjnibZRzw3PWwcDVjzDKwMv+MUcpjsZC8LVjhcBc9DD8KHSj0
mAWN92CL2xlEjUWbs1CiHCJFlM3JaF2/CDd/JvtOWDHIO4ZscEugjF0Bl3yoieZErE4UTfnJWVzZ
tKhrwYb3Lv+oBAMRSi7mOS3iyFfvkccogVBpGZ+z1OnMV0091YZdc+m+G5q66BF6EOF/8fNXlWUs
XhykSty/MeLXs2JQgL5hPTYUNXsAyjRgVYRAjj4nItiiM6I8vaYEaMYaSNoYcz23+tUhdmBX/t3O
liAIHsKRfJIvFw6Th+qKoHcrVxzZ/G3DhiGELlMX1sr689UaTfyfds/AuSizO7XK76SOx1UHuywz
xVzC7OEp9ipTt2/3mzab0VvhJz9uk1P0oDY0waZATyIFuh/uYIY18uoLur312k30iERB9EgkiQ/V
iRQ9itGlf7BHKFBjlcXubsy0vXMzJkAmWkJ5YIuBWe7r8wUpdsySlT9OeO2W03NsycaWplNBzhzq
52QZfrNwoaQHlJh8FDm8z0eWin/8nNg9D+O2ZKM7dSYzZSr1AwmlwT3w4nA5lDV5RzRh5V5PM/Bo
vDqjEV8IKTu/q83qIQkrHxrQ25QErdjaQkjIhdx62xkRoptE9hLVq697Zovx0v7+9wQ/SIDgMqMf
B+W8GqP8yXMRr+wxy3OZpEiJlbQNa3Ts4xGT8OMPFhwXgIcSuAIJqIIqQkKW0V5SzmaT5wwcVBmd
U8rjcZ17xbxjBd+i5oD2jdASViYLUqXvBCn1fwoKjXt0By/ner6J+u+MfuYpSa2pg3a3fZM2ivQm
E0nXUToXR95w22yxTymWINulCTsm9JeDOcPsy2wQ4ZMsozWXkXNhlzWHTmnF/cG8+yf7qSsACOcj
ZXO6mkzkXfKDI4BxNPq7rvpkLzWsoafgyiTd6ZnPP5z1pxE3YS6yLVNwy5enWg61EwVbRGbk3Nw8
j27xKGexs59wkNEqNgJhuEbeXuov/Jw3IN0H6YKw63khCDAPWwqEVRfPwePWGtGeU4cBYYLKDN/o
oC04gbcE4kHBX3YcQa4Xg+d3CXYAFnvZXUS+p6KufAoV23UqNnR9CohRkFx+G1C5Kv22dpn4PRRM
kCA+1U2L5gTvNMEftfEPEPqggJzUMkmj0D8N9ZcSdNCmNAlI9migVOPUg3TnKCmV2IJM75FHxMEp
l7XxKYsJmmQPdE1klF/+WCZx0ugz+PBT73sdl7cNf0oyDDto+GSOMmSGH1UZQZl6Bw+vpfXDFc6N
35/mLW2vnNh9h06sBJdVokDp2yUXRHGKxEGxOdHi+hg2KDHPy5N71vf/bk2sKCCP2vQDRWn4MuLK
OwebZ1/+rwDvRb80IWlt8ttqwDBZKXnH+k2D1g5rWNDJeLNm4XpLEYYevg0gEKznhk6FKhk0ovoz
9VHq+qCk2hY9RsLSaslGn5KLy2kFz3a/vj/6eV2IUBG2OuctxkLTw6+dWBIrxJuyPgtEagO5HddB
ZdTaYqE8Jn9zQJnyfAHEWLtkTF78yY658qCQKWAtPNHlzYVw8fE1XczgizjeDvK0e63kS2nHLPei
uk1z3s0pIKpg3SN/lXaNG26IifsGyymjR76leWVcxUElVxWzbzP64WOtAFh4xdaY0m5iIeaNHUHz
11lmJyyPLiT283LV/fg2bhyRC6mZPhHb4IlyY7aajjMzs4isn3p8yRAJmpcPVq0WADks7UA15x7D
PMcTXj62lER3LZv9pH+NXHJl3Pp8KVR+UNgLv3SthY2+tdSknRDt6tHkXiTYtT/RySKoWA8LuNm5
/CqbmXkNxkJ78UQRvw0yrnkg/+x+vAN0VVY4/j+Mz9FFY2e4zypQ+D6mrK/sy4HFvYmrQJh8uLsX
Fc7GPNvPtSayCaEg//AFfsf62y0mJXa3x6VsWc/A0gLTm48HD3ckb/5ZILx/TPULCi2qB1LtrDYp
KFNZ7QEkKn/ErAOYZu5JxxBejov9oxM1XNETikyHHCwv+EahO0yAf6Irym0hxGUKk9tooIImI415
UZdcr4wGFE3eiyDJpa8PZ7AylZTwZN8W0VL4k+m0AEFck2pu0SQN/LIY+Mum03QJMPQzSiHGfVnJ
aTE/hA+8mYhEjJki72iQvqpdypJXLteCywWua9nUdoNn58H6IgSe+3BPCy6CoAK3QV4IfPygVWRg
fwagK9g68k3g/UGo4h0RdiaDH4/NEIBXKamAEqxJGf/LEzz6Hi7vArE/7BDuI68HzkckfETMFnT9
aNBS6TtIQJg4NRR5l9aV91zlb4wPU4khQ0MsSG6Xe/pIKmQ02XtIe1M30raaeo9bAKl6QTtGfoML
mTtntp+LkdmM7Msd/4hoMPh0n7mNc1Dvb173Mbe8NbdqNG2yWYs7AKq9nIrYEiutfOZ6G1v4Fz1K
nmOITzCJjCPZ4PkEORL8qHoVjTj+VD7qlGOgcXY7+/QJP2BmFFJ2p55z3wU3+gML/N8VdGeLXnPI
xEj4NJ+gWbaM4cli7N5eGUyhV3px0TLiN58eqf1huHIRHFvxq4hr8UT1CUKkYXxY2vlNJArwPzoV
iFfV0EGHJZp1y0X9O00UxnGH4gadfR52sh6I+QaU2ucawIsFOA4QbJrmrmUgioBEeRTU2lnJi8M9
1qfIHMV+xP2F97nCKquDf1k8/+0NhlSg7c5fQsP76g4+vs1ApDPxvMKgDK4J+sRZjjR6M0CQSU5k
rSJSfUHsRKgUAt/yZwrTmyQmo8ppPJCWEfD0fGDokD7zrEzYclnz6dm6Ge1sF3ocIlJM/MEUvDsA
FTOhzpH/BwvIy1Yeb1VCORJTY+sEtXikoVoU5pA4pQLZl831zLHXVR7Qfn8nxiIOWaJbGEVuTf9F
dEpW6tOxzrdakU+dNYTk+TtR9T34KkoLt2HbFRh1waTtZpgaStsx4NOH8lN0Xh02ALGYpQ3KJu0x
1KuClctVL5iNK00lLKv374lugAJsfxSCOkgEf9wZUDCTUE2eXlY6LJLmCEUBq86P1Gd9l0rGltv4
kaxV3BblrGCUlanlcyCyVRhfwc0wc1G1i3nvTxKPlWPgOZ3oCWnaY3Toi1tOCDOcP0RwqEfrT4yT
W5C5nHROzITqcc2UrAgf0sjcYzqrKR+UARmwUOSAtbjUKt8eD52j2QCN4RQ8NxzJWBS8+g2NJXHC
kXnfjJF2aVupH+uRvIulN+LhNRrWqNyJHlgbDc5vK3t3I8z8c6AfYoUda6J5+FOTgQMKSbo7d/Ve
waQlSXE8Nhw2VGVGJI4eYkUokmVJrR3kQW8+o7R8K2sklPpIU3VuMarZQXfVmrhuiema4sT3ovkv
9WAZ19H5a6uTzn70EFLBlF3ahSjtS6CXVcjPElbp0BC5tVoTc79lD2ok3nb+QK4RY5DDvxliJnRm
oOi8ogbwz0QzJRGpKl0T/sXseEqs0SV6r2u8V52eXQVrrLcki0Ra7AnMrAQiR2QLDhMJ9ICAp009
XsUeZ+q+Mb7bDAnPHLduZ/hTf+dGznOuqeEJFKQdU61D98T/r8xyz3ABZpieMlW6zv7+XIHdEiur
BkYEFFhszihIqhGV30cnYkgzdKI9TY/zmp+OxWIWuCcpLujypFOdFd3FSchO1G326caGeIPzpK/W
93xtZIuAkt2Xy4EcO6KFbSFtNWyD7L0x6bulmNryKr0lyn2PIAIzlJMCaIubyxp37oQTjgXJ4VkU
g3hF2EAj3Pa49LH1/VHb1/cSdqLXURrxvII1+LMDQgAK8/NydAK3Vx6GIrLMt459aNdjueVNz0RN
85pTnEulUn9C0i/M6M6L6MTKB6G8q5Pi2VB1QyjtSWcUrqsm++jfbjc2NltC9hWC/XY05o1gM2fp
3NJTM6XOCLSQuEFJ04VSPC3gOXNBmm7/yAi04NssnoQT7rp1RHGKnv+d1GQsGcLZWYg45IsUmkQh
k1ZGdcN89n9LRsWyud5xgz3Pgdi1SewCBiC3C/ZURKGhIOcep+ClVV+3gM+6NjrsGsWTM5OfroN8
t+dz5r0YveFHOMeBPx0V3RwdrrASuOy0awb23D/DGaVhf163lesag8aOZo4qRjzDvZoyV8174436
qUV/y0pIALI4PwGuoMNEd8Sj9PAxARNXYiSEHeNABSKPYINNBCU3f6YZxlQQLBsUAlt7KXT9Y4kc
5enZp4b0DRMgR6yE70yV9GkJ4XTqM+IJdX270M5KpQ79/Y0l48eXNsf1jZspEaKVv0hPWuX5pdJ8
x/Yjb1NTU3R4Ou2QpNB5FnNUxopCWP6Lp/Cesx43psRs5elmjvPPkcVlKLegbYkzfpkToDnjsC/4
koDc3apGpRnMbP2dK6XJyov3niL9I+1VFcHGsoUpbgWYIgqYlnv6gxJtLnmCp4w+GbGr2RjPBBpY
OwJ+49LlCXRhzOUCLSlc0Fg1x+Fu16r158aExzKbH73GYmZg9OUvCV0vk95VoY08YrSy+IZqcGdJ
khQ4eNcMmqTTKcTla1iDZ/0qgEWKUHBDdtNNSNsfL0+8D6R2VyNle+yz/ux0ovY+RSfcE7afB2aZ
C8jfp68FDe4UMKcSnuzbmaapJvtDdXAKphcma1/50p02PHn18DbcH4bRsf/uOZbzG//pQHM5X0PJ
BxnKHYbKKtohum4cJTf4JXcFtqMryBlw1eLfIJD7BID/qYZoErBfzLWqGPsAblCzD9wzrm2TO5Eh
lQNukMv35T2qYiO/RXO+TOaw1rVkvufUJmBXHQIBsMIeaRTqnr0LrTQju/IFeg/qs9085jlKRIov
DRX6wJb0rLQVdajDqHkQ+kPs1FfQc61nU8szzGLJrJOR0N+nBk9GqHbnv2qBQqhlZ+7rHDwzd94o
/7XKop7N1LCqJISiszzgw5GqvEIlr/3ZZl41m1DgWYHdgd2EHLA/j4lc80TB5MAetcO9sFq2j8oj
5Bxfos8G1nyZsgWDYIeAmYEujlwp8C1V6nLiBtAvdK9vRDtJxmy5D72eFqSiGc0Dsj0OoKfbMqGu
qU+umzcj26iyKQh5VrVf+uftsKwc41LOCCMZD00zrbo5WdlhVgFV8NnBX7dCJEuV+lJXg5mKbNGO
cBhrXa8ptJUKtXGQ5uvv9g0YI+WGqwXYDod8Ekt5QIqhpmGLKWhpAwcVud2xalTj9O7JMEHmRyr2
x2VpyaNUd1cBN09tqezKjHaEu9ZpnDHlTcVUY9oGSeviDTPZgiSeurOxWbnRHit8M7u73gGJge4B
xscMpU/zwGMfVjmDqbQI8YZUyZzRIw2wWvkqkmHWgR4SCrbS6t8kauhbVBTNwmJjxenugec+4TCl
1aV5jkKOnhIWfEI37LdVHbbEPoAztqzvKmIJrxv8KGbnCHhB/w/lrfi6b36TwuRqROqeB3trOlzN
znNJSHEs3KzEYy7V8aYIEdbpebo9p9fYPWgNqA6ZhAHDIT9Ma71BG2XhDP2WPNZJMQK8NhISORTo
TRc7mKCnWE8Jzmy4whQxFpgDgL22bGAh4NiyA7dzNdNsnOSOow5gPOT7iyHcWTzazvJecfYGtQ11
B6C1caIEE+VgdCmECKHDXDiLsNts1t/7r6+DYDthV2SHNzbFhgULRcic6ur3QsR9QCzTXwYROCxn
5Lz4dTARsNRJ1X0TQ22hp0JD4cZ/H6WQdrMkN8kR6UO2e4m7Gbw2pC6zvAi0EV4/OFmMlu0lvviQ
SfSnYClhtXJ7nvV9WZaU6Ma5uIeiN+Td/mmzNxtUr/IA7AZedYhaNKPpOb7qF5T1bgPG3NQYhHsH
teukmO60/7Y5SWv2H5L7T2zv3OlHlUgm0j8IE+NyfnDDL4WkstdgcILkaDs14C52a5YB2FfKDrn7
Q94EkqiCj3ORu5IH53Kk/GCDE7KTkp61NZO/SlpwjS2Ee3pnaIAawvBChXNUWzAdIo29VPkjUTDi
0sPoVuG/PzgxpT3fZVfJ6INKg5cuedmZtEnYpJ1wzAw5MowqQajaF10cTqhImPQFspKmbqfvt4Wi
1gZi47w4XaYmLJj3jrMwz+iol5Aif59l4M99u+6jBy5X4Xp8kK0ZoKw3N4VUaxIdU6GYru9a8KiI
pKmrKg7q/X+tNALtoJBPf6J5SAmzTjgt9hU1WdY6/m+lKa3WzX3dgKFPfG01p3UDt/5ySwyGkXQm
qbSUS+S1wPoHe0ZpfJx1noFQl2GWzkR6e/4kHjJbSCGdZI7/OaRzh3NDLedAyqDBO23myrc9OVL2
yxlJlGTAgWEeVEUpFp79TyhF/qV0+ZPt4kG2Be3wJggN9vksbFGWl7g+p4Ph8HW57CeiUwAs8QVc
C657jrKDYad9AaBrBbatBh6cIF05IgLimi92SVAKvPh5keQpvaI8U7ta5Gt1wpUhW0xffOjxBuCF
SDKU/s0VgZp2QVxCEQ1x65lvSQXvIZi/wvyEeVzNgic/3d3uMdU871DsavCDYdNi+BcOGc1f/l23
VStPqGcwz+VpXkx26eZVUJwBDDEjHiQ1jbemx8wvQoMCy99LKlubPjUFzrDG9ZdavrOl6lRiD1mz
LT++5TY6Zn8CnBTaM2MbQTuklchHhBq6UJ+4OHlwXlUWI7c+hS7Uicwf9qPr+n7n9viRRLOGrSLh
VMNfVQVMujwuiIAH12QcoGU76iyNRZvqlC2Q1YqIH24NFUexCQ4Hc7j2oxW5KWmQe5mxzlwNRcr1
t0yy
`protect end_protected

