

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qYvaWTl2dVn1UYauUm5HneGLdmTNfKYL2CALcG7YBWzuKWoXlk0Id+l1oLffyjtPstUkcnB5XMcQ
6NZs7JK9Og==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYtaB7bKNbwxVddRWt78CWZ0keZknIQG6IQKSIZ5COH+hNdpgy+tCPVsEHq4IVZzTG1P1o7hP4Vk
F8E4xV3B+P4d4XumR2TMQt1O3p//18K5GFLVc+tXegTNm7nDlHWB2EseJW3Comce24tPY9JdBxY3
PqZ0pdNcJu1q3elLkyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dcPEPRyvFmW4PpA4iDmUUiTH0W6w8Tp3x24VnlLzTcuDsG/S9IG3GcyE78eNrT/x0pAgwHhrMrSY
yZo9WE5CUIc2230lFJdjwqsu1GfylgdJvImjNnSRTPzlw78/vxcWd8GQIKrHyFhACpS0FlCWX80u
ir6wyey6yythPFMR7YL9alngEab5jqlcDLLq05xFb5xa60ZtUm6H8H/kSZM2WCTQ/2EYo9aRaoyP
YNJgznw4M4JlCmjNGCsEEMbnrUH5XC2MOkUpPSJ6HpAPhZTjHtmrQy0MjGpBzDrrGJZmxlIzL7x1
7fFFHCW51Ue16QvPlxZlJr0kCC3nTtDv9f7xsw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zhiiGh6iqBtYa8uvzkWpAts7vZ/x1/EV8yeLKnAXP52susoGuPOfmWMYojIG7BJlvNdJsqMcu4aO
YgpCERsfm5E2WNcFxUppU1uIOa+cnCBSZ6N5aebRGghJrQL1tUzWpRnQ2slMJ8Q+gRbsoc3N0qtc
A+A1dAH+z+hdTGoZBRY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lbE1QAVb48OwhlUCQuKav8khO5ghQAvoWa4EGI1wknY/PAoHSz/mN+mHHLZytFcumXquM7gAj5vW
FkPYXzAy7xSUZBC0WEUc0yo4Xa33jDRDxY7cxGlzHmyb1RsXl0duhVMcX5rDmM/+KiXLbAmtS7n6
pXv5Z5tj4x3AoNn90rxrYgdqN+pxQ1GZhPZPFZggV3JHWj2LJUr0U/7aGlgZSQCcdWV2V8ktlt4l
b9BA5BfHfgn1UuvjTl44uqXII+j7cWg72Zy7D/yYZ92M5Y7nPBoBrEiv0PrxnHLMrIv8+jN76TPm
TMiyhLNg8NAb1xNexvBsDmGJWQnxf5cukp8uDw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`protect data_block
L25tFnUSScn+NSNZEWHyUx62X7iOgl4pPW6qXX/RlCYGyI5zj1JePkzoNWyhbhCLx6mrDlDSv24i
WG89UVVJhyQzRGU9y9GZJPu9YHXfp+ojQTEbSnNoarZ5UV06bB1DHH4Xymnxh2BERmPAwxdPXNmS
kW/S6o/9TktZEOsVx7TK5gxRVoBKnTfRHSK2g5mkdhHZ2XefeEVaOlJUJDoWKXCNUurJTFM26Cj/
/8ebfiRJBJ7+N12xrSUzrtRM8XyDja6yWqNMlna3MvPiEDQyCgjTiZjy4mNcn39w9h4EWbL+lH6e
YPHORhpBJRgg48hrsldPsP76DLovj70vyWUdj2ibX8bJj5PyyAZDs/e6juGyRP1RbixfyPH9PtSc
kX6+ZzohPi3cCWHo5dBw4eB7X/Yv/8goRoLwMdxirNb/FgeTHW1CPwS/whBla7YmnKWBJhYh0LkB
qCg22nqSVraCnA0YXwG6mVc2QW1zFlhrKZ+fJEThfgc+7gw0RnaRVAb3HWqQdFZnCHy/2DErat4P
Eb8RZQOKkfuCc7em2veH7VoqRpePteHC3FYCvaUNajig1P2VSRqa9neQwl0NN0myLphk+31KOCHz
i3eKYbqmgxO9uOYty6rvfc6MgVyl0ZZ/cOJ3S315fkvWbXyttxnErLC4hU5LL9xrAp4t/Y7sXVLy
t1pDCcoaweKA4SanFJHXEl3ZTGPoiW4mBPMlt5QyrdqAUVaoNdC2HyWAMgIOYgpT7Z9ruc4jxTUj
KillS9rw6hTEtCd4lX2yA0reLGyxt2vU+nM+qxkmhCWRiIf2Zv7rFjdygCeD4kN75IwioxBXHjty
UVJfttFQd1/Q+o0zVldLcciymHxOW8RNtgvJPgYxVjtJKnXvdOwy+8pDJdKB4w6Eu+65uDqYJ7D+
2NhSqeHmmGdL1Il/IElMm3XujV/isTvn7/CgHkCUTdoMYm8yD1DDakGAtTDkHmvajGxceXtqbUof
axr2vUC7H4WtopmHzZMpzzrTpLoPR/ttUGBTtUWIL1ltfGNYUxQqbGGMyVozQ5PPTuEPmqBIG22q
X+Hiqpd/u22TigRfYMXhLYkWQmbGuu1Wgh9SuT3bBGRx0az2DhYQj5gg0Hk84PnnIeeCuFUSWP3J
88D9YpJNm/EzexBr9zmQz4dsU90JYmLNtXf9/InRzWc4Mwqrk3TTVo0OaeWEKwTQWA2zu4xQQmyE
wO6P2HoLBdR5PB08XePaD3U6atbkIwj61xx+a2IQWy6Cd0LCosuyO1LA1uoZgKGYbrQoWRjAfvUb
AN2m2v+DIYvgoYY0Kj+/xZuow7WaA2hu/nFVzsIZlVOl59af5Tbu3YlAGbQH4I0sg5YFJqgKk4bq
U8izz//aIYdthM2MMJJv3j/wX2/W1LG2+3T1NUbJSPzav9BK7Jmi/Zu26kmd+WCTRPICouB/+Q0A
ApQfAC2yvfQjfV5z7rrnX8xWaxzk2IDP0mR8u75M3a/jmKOeW3DjEvwyyypzhsiBaXunOep9vaCL
mPhC4biaOqqeue6rFUvmzrPEhgfrUoyzTq6S9Un578eT0doRE/fURTb1GCsYpI1aETdS8BDFWNxp
/uSXSxCiJp5M9KETWpeA7XgkoKebFC6ZtB2MnOreZ+RKhxATakV6+wG+j0DBB3Fi/ZuHg5gYcGIi
e6yLuybXdqTK0xX/VfasMA5Ax/pEQ9Sus5vWFzogRMDnHYd8ht0HGT2I5dPGREv2ekZIy7OkqpzB
xe6Md8IlEDc4ZYptOn3UPbhRzcbWpcWbyjkmPYcrztY0aeBmNyBzRpAIGmFfRp22JHIkRPZSdUQ1
zmXTNqxBxNc+ZnrBKftpNV8LotRLU/XLmeY8BnIgNC6psgIiWQRFY4hAM7F8uJ/HLwRANuYOwysn
+/iYZJ69TQwjahHvDAeho/OrOIoKGD0d2gFA30vRtTbrK7IX/jp9KFO7gTKlbwxnFgY0xI6N92Hh
xiF0Lx0mTErvCxj/bgsr+GI3lExP/nUXUZKDyzSqdfDvewM5oPQwzgcK4Y6Py3kOZn1u0BV5+bwt
j/OcVntSDiGtY96uqBkJbDfzhEYojJ41TL9FX+Q1Eq2HZVbZpyQAECQAd28o99fAyT/K9WXLJgiO
TOnLnvE1FvN6Kr9mFFIBk7yA/eny+MBlnKLNfjqsIF5pA4Y//YzdowA8hCW4cHGfb5Y2h0Jdzi8X
R3DDwMhZ0889vs5b1NP9GUWHGPZc02cEvfLcrjkb21brlvs/5IdCJpL6iATgZLTtMx9vsujli4TI
1qbUaCC9dKhrBHvthE9YR/U+1iILQDO2q6gjRnVVHjLyoZxqNiU/xZmg9ja2UtekR7+nvFolYeEa
u6h/lF6UhDoKPiX2tTg6enEMb/9bJK5/64zZZgnQXyMVyBhoVAHSCb3utemvGlF8CEA+rDSwRo4c
uDmBg1y9kpnpKuEDsAa/y3UtANBHcUT+FN4MA4Pdmji2k+Bv1ayhTzrr0alDObTw1T45q2iyOJvc
ToSd6fAkSfED/6PLLephDikWn/eKMduExsN5tjutYYqNx8Y3FfwQItvZpL4YPfdWQJN23NJZ7oW9
2+izNuXZ8BCp7FCmzQdQ7x41Ry1rEVFUXx8XXc36eqx3iwjmGyZE5KlmeZFpOLzNTazFC39pzmA8
K7YSuT//Foem722mtIKynrDN12hLTDUKJxJy0McJ/lwz/G6lA+klLfhc/mcAj4G6iO2IVt5L6bpg
6nVSvDzkXvJOVMPvhugdj1wJJniPXJ8GuYEP7YU8Xr7x9QZA5xTkrh7qmDpMsEooRZFIz41Ax5dN
/JcbFROJK2uIjgmFR6uxU64uqGc8HqisNFE62hurAylHckA/TDoAj7PyjtMh5iUD1OAS+b+raoEd
oEI2OSYi3y3dfLD/Qt+0n/O2aCN31pAJwGqrtU0t4wS+YOG/0nZEK5MYja6a1IBVxWa4tAwg9S/L
tOzS7C1FVI/gmw0PYwmq4fpzEexm8A/DNOYy2AcKSYjqm4sgWUIT15NVeLlg5qoyFG2xl/ClakOR
uZjgR8e9UjkHK6zn4xfGLbBxY/t4j4Z7jQ4pfyHtf6IC1BrKw1rgMSi9C2b5/91DYjwBJYUVYazE
fVMyrn+Ycgmt4xi2w2RylAnN3sxJcA/dn6BEW2TKu+3p34yWyuWlP3A2OOyaVSQ2iNJ+EfUVCwwN
ie5JWJlunrt6DfU7lea4kfPyMzzXdBEoea8i9N4JuS0QXbwoDAO9Wp+WGUCXpvx3nqnkWHjhLsQE
Wp4Db5Qj9l3Ma/RnpAu1HYziC4yorLUfSHtquMUFO0TLsW3nnuSBqbAVOHBG09ED0CNesBH+6jQ6
FbVQLrAwbmb4sFfV4VyGyoS/6rsExl1apr7Pd2TKEJ1pGabRLaCF+dBkQKTCNI1Z+hy03/VD56e5
IOvhHw3PhUKLMkzB5fPFI5rIUk68nBhNtkoFNOmj2nVfg6tB+gQG8H5iD2VlyjFpEumKyVt7ZFY0
CHiWZZoL7CihlFpN8BRqvQoERt8w6IwXy8fBkagEVTI/nAuL4orGTBIDXL5eN0Yb9ZRA8Il/hjH7
NkS0gcrBSga+7DCWw8D8VF9yHyibMxkkqrnSPLyIOaKYUMRH/Yaey+nwzfPTc2QETgBAVQoo+b77
iskb2tPY8Br5zOyrYbZnz0EsSQBHq4j5b5t9abwmDmN9Gd8tcUV5nbe4UcUc69iCfX/sFbb4+59q
rR8Ilqe7atnZhXpufFxDiUZDTuUOFCkJ8UjLhsbmk9ArwlWDzjKagelemq+REx9EahrAlAv+yBqR
sGn7waNNXlzJAkooTfuezx7glURC6niAMAN2AVg7g2uTV8WNMbGkice/of0uFylV14BRJqcGTFXr
A7W+L5rrKnbWbK+ke6tv0GmFjRqlvnAk65eltUxXcYB+HsD49tXGAKzx5voaYWoloImxpJXVdMpe
9tYMqTT+VTBaCRlfmF3JZ7nxyaAuvjznO/Urv3GT6iWhkOCMvb20VsKPrWw4yLP3sSvgyaS7ciec
WQVQKxueHAPuhi6MOIEtLzADzQ0xxNV7WOrG9jVXE4rA/7JM2QcrU2AWDFvZlJUUM5d+hWdzQpq8
aH5cJKoDza5I5wo2zkxLICQHqFQ07MryQkm+H9xCIqNeGnC9e9BOSZ4tSG7Iz+3X7jP0EW22oUHO
0PStLmZ0ezvZwKiZ8pzwIQKwHYQ7fDkC2gBTo/uHcYPwuf4qWyrc60GkU0YEotK2ejlhrX4ThPLl
QrjMab63QjYc9CshLkvxu1muMINPx9wLhNw+Y2lAYP1wfUPoGC7zbqr9zAgZXx/Bpx3HG6pSMiuj
Dw+/Rl740+9Uqor/5y6n7LGEBeC+BvmAlBcGH7qIgsdqHmnx93IWqi3YtFVJAUCEoOU2lISZ0sYK
vurObCl0khJmRkhPKJ/42L5FbrPb9hDIv/i1+HL1paUsi4eckEwM8xcmTxmEnOBjfw6ZSj/4kXPV
aF4XvxD3UaUboX3PU89uXhExeYEvHjMQfFuFCGtAhuMwk40oMGJ2gHy4aUvqiZFcxLmG3MFl3I3E
hCmidv0KyndiRzo5xmHsR9ra6XZ6wk796AJlv9vGxnPu8lznxZySFPet3fuP8t+DihJ+H9TQQ1In
Xgy8XI/00ZsqsLHBKyF9cJviKnPjNrcfFYGRVuBH6DyFPTkFsLVMSKXIhuPhNgJcz8TfVbyN0ztx
HBLosZ/CWgY+8Y/Ds1795Jcph992jBo0qjtQrSksL2p8eQDs6cOQhApY8Eq93JCUpoZ1+AdWT/iV
toxfy1g/83hRsX71BunSDqa+T4hlvnTyiUNqOQOHDCEke8PYE5elDlDbpazyeBkZuj+f0XZdub65
AN3KnTInx9AXdBCTc+LrD1Ba+dLQbxOINr8zfdYCscseOYrCLUgP29wrwTpaxIOffZT0PMXkX0mr
H4mocnT3ncCc9UVi+SIWgKCRaGfuy5GBuuj5zvCIr9cpZePbn0XWqKo/X0+nkj5i9+3oKUnw2WVC
XrpbDNFNuGaiSon9F/yr1Oho8q4B4k81RYbMnqOjBbMeQfVPaNHhj2KO/QhGi73bCKfQm+OEpB9m
Qg+xB0b/XExKII5M4AQ2bTBPM6uT8fytgJQG8aBKSyd752CYGYAmL0NkBl1cjEVuCpr7w4Jpyep2
uYWH+N6GhJTeHy5L2gJBVv5WuliYoIk2no4d216kJtwedJtcxJ/CTS0poh60AmmAySjXSUibbJoW
DOG/aVAAWv0PY2pqba0CgS8MIE7p05teIhARBGQYaFcF5v1hRNjkWPmdVqOy+iTC1EOrJ7/nouzA
e1+zBMN9BhrM5HRwmfC89gqQQNcqAyvgvuGVqnSstDzZCfKLIuVww4+PK6kc0ilppcNGUhcGs6cM
XtyHFr4QxLQpyZnZApXLmjP5K+KiEFx82UKPVcpolAr/ZarpgPnrjymnsRJGJHsdfXmfqsjtzxoF
zgWApEqEaPqns+XZdf/K8TaGyjlraz/6DjEnV5T25h4eGb4uWyeqicj2gEcLuNPXduvTjJuGdtJI
7q7rM3BU+6RG9UWigrrxGm4vUK9gW+qKtGPlkcBwh0pD+WLsYGoMLwWbk3o3f6AVsJKY5cQGVWsp
I+cPfJrnwwgfdDtbvjZ2v1TwxvaUAnRoQr+uaPoNhZoZM4QjF82KrY4txsyy4F6/zCnFyyPdsxDm
nfOCVvRhaa8pAbC7HwK3qqr7byEOrak2n76CTpoc4jVdXmHUdxUDQ43nr9cn71TYNeiIwjK4iMa/
4rEvVgbRmVB4+y4YxJcnLRDqTrQigdXwNtxmnbliRRawDvG6JTiDUUbwZFPiqYIGtjTW+y1IPxiX
FpwYNCeE/J2kdBX1x14E8zTAojkWaIgYd2mv+DLfU2bNKMZoVb/uZ0rgQeBLIiqEu+Fctk5MF0y+
SjzKuCUSAf1BJuEuXOq7F9YtfLFlOvlHBmPi84Bzhiy/p7DlOdpcUeklFmVx7epuGLy5gBjCs6Xj
ls31YXJcABJiXXsMnV3aHiA81Af1KOCBcVNor7RFXlIpzG0xaXLCRFQK2XPQLt5H4s5mgzCYq+m5
YC5OBU8CpI6ACIJO7ADHsWuFXYNIw5X8AlPqxKhDDtupOtkctM0XfG0s4U5wL/8GCiLBP5mSG1NC
B84ElJiNG/6H4Ps/Ev0S/FGWoWlM4AXY+RayWvp2ocMmhMPUd5XdmTmpX202SFVCG9yItXKXtKR4
A93IC3Or+ObzRuETDhVPi5ddtnlTl2K5i5Y7djVXpnkn6fhwXmuk0Q6OCAj8RHqmgNViVNc3+18Z
Xo5yh1QQNCVC9dTcUowJuPqCX945SOZduxmA+Iwfzyu9dwAijR18Y49k0AOLdpZ+q/2xYPr1LGJ1
7r0FqOVq/84oyf5HU13TfnqVTtkOe9x2DF9FqDc4ELvKj+OHFwBbE2G+x8703SV2XW/zRabmVxCS
FJ0hzW/JgjlOkwBkyb0tv9zkidHPox5ebxx5DslXXmh2miPQza44sL2PucldGSeRY/1+8h5Y7r1q
fZVw3wvHKpHneG6xS0mbWBwZGjaUO3sRFhzPxzkr0rLb+zMpAlh3DT4ufPoLu7hVKpEgEfl6OhR6
3KPbkmiyouttvd1EcWvlJ01aLmYFyGy49Kqk/LF5PWGk+YObqNy2dFcyL1ay4Yc8Pm/QIlhkaPt7
D8K8D7xPYEtQ75MFvFl36J6pbogNcAVn4H9Kd9+ROuIdK56jyerT3VnS12sypBK1HjX+U/nqzoyn
mD6Yn4j1P9hZ3iDKY399n2ZUgDuVOgyVtsknFbVJGkkjfwrIjoF1PxCFXQ7K9ByrZqtox+rohItV
7lBuiVCxpV+z3630ZmIE1HVbpe0LlaPpqY5sDC32YHPot2WghyZpAYlWP2DEBFAI8tSM+pZIjdSF
jQ8ksnjiboNkZXUTAtOfZp0U6eAyFfIYAjEQcOKgcaXarhcMs7xSw3NGczDgs0pH8Wyzp+N6tbuM
uJxq13eyThzdqMv6+L3rQXWosUZiZritoph3vlv1C99QEOGua0yMKUx86fJwuzyiZ5l2+r9vSB2X
o1vsD+v2K20R2RG9lBCSnrOC2AVYrNVil3B8GDeBLgB/z++ahKxuIWBQZJyNEEEjBtnRgchTzgXv
RLHxYrZf9cNjzXoeraJF/jUZW6CjbTTP8Jj7QHzh/8XaY5LRZw0RUzWtaIyrmIBR13XtkB0Frr5a
BWdyPeSofXnDcAD/vDfOwy+Lq0vAXZCJ9xtwoMxghxqTTz2vcCKXBVbqTsvtGITKnjmBWGMWLUkB
qQervkdwxKbuz5QOS92UPF3FSb8w6J1ScvNKm6lt0aU8suOmXRMAJVfffsU0aArq/lOkARmLRGXG
EyENL63CrSpElGkW7oZQxlK1LH6Qb1TbF+JVv/mHpmla69AglLlyf5kPlvV7iVJiJ5HyztOLmEPx
IrnVm6SdlqyD3vDU7qXZL60KGSlbEk0ApKJIbY4oKtp6ReX5tXx1VvXMsbEldIKMx7pjD/IWKPci
dDiuwoYaMc0D31bHRs+YLuB9WO3QD2XhtrNOnL3OV3mTTCB8+n3LJJTsKNrazN6S7iSM+qkEDnoh
io0lMxAR6BE49AKgYKSuvYzxuzw4ZSG22Gn8gP/uEcmdLmbOZR21pnKUqORMm2rlJdNJorE7YGnS
IzVgqL3e8KMoEK7Y4UQtLCmbWRd1bBgwvltU8XAxNVo21C5W9AuGEuHuo8QqUNQDQ2cwz9kwIq06
mipW3ISbIy5YL1BdFop8VEbBH+/HdqRpv1fsu2HqK7tgxEx85gYrJr7yFugVuP/SCtdvPVxHzAia
kR3zWLq2YphMnhyd8FAG8pbyUhEwEwm25QQaR0Jc0Yril79PBOR6SCOGGmWxvjBGqSfU4m3sf+lR
oOcBgaR1WXciUXehYaXI30S4E8IfplcxKK5xO1B2z/xT0vWiWdiifLGqo4ltjXLAngOwM079FwcO
jGwCGCSqQaM/Acn5CN1avkcYkM5YUinEHEf+wHQQLkUOfNGVjXrgChff03CG/SMjI695Y/WPqe1+
YesaMtWXg1fnYaR+dNm0BJye4M9aMJMhh6wy/f7hUflzbX3jwX/wWhMRrWkaAfK+nZROobXsEKix
RudETR47i40bdu5AN3NONnhFeNrKjVoVu/4RMmij5TX5dil9nNoYEasNgCTgkdTnnqShSsz5tnIB
uJ6E7BXyO7VUKvKYJu7GdabHbtZjRXbygD7FEuceHgtAJWLxVl9KTq4nvZ7LyluR2fKMq5AVsv9S
aEnJEPXGqMBP817KszBdP0d/MgpPAYTLEzcoU+Zp1J4x0KcNbUuuhgfh6tTOCBTIhtlm2i5Y/IUs
tm+Yc0GTnJ8RUVsdkSCyBU2af7vu3v5Z29lyjAdmg5e9Yl6t3F0qjh6jNLsipRfisOVYGGA98bFB
TgmLb05k++pgOgpuONYc2o+UeGggVpW659kHnJyyncK5aincUJjMT2kV2DqjSZogJMYt5HupnCb+
q8HOG9ccYkohOZCUkSn6PKwJ8fx7Qt6FyRxRDR01SdAMa8Bfc+FCRzq4xVtmUsCA3AwEB1HMTG1A
ROU7d9SpKte2NDFsk47LvlFhsEYOcpBSyZ1hZoa6yDyiHbvLKBws1v6e5oZAbuG3liYjmpEU1ZOu
R28CgS37vYEPZAkBYlf7WA8t3lMXR3ZG3rZ+b6D2pCfUEPy+EbVF32rxhnSieARN4EwvUcZwzqbG
X7G7YimOeGEA7pKIJyELfsV4WgA/TotPXxrHPf0yjVCwKfJNUi1wzIIi4qapVdftt5/yhCQY8jiN
+9XGTC5rgHKq+UpxkYlqILRzedUWhCAA/ADsq4ftQovX3WV7Ako0IN5GcdnnMQD7RKT1HOWm6+LO
YX/2E+zdt9YF6sa/BEckBLxqhmoWuWdZ1FL9IWkDhRULfMFjUpFmvcPPGOm/2M1MPj8pJ1JJnL+N
Qk+3gHvZMQyzrRV1rWACQMVppO0Dj07GlvlQPM8hTlNFQjGtSd+Cyu+cYpvOXMZXp65bowL9fX+d
4jbD5nts9s/RnSADfd/gs5p/oppbNKNXgbOEoc9Lu9o4yG7SJUfecrBN4lKnOhahmm8QKNyu4uSt
6QDn+muhdNUpOLbZAhpyCJ4aQxhlT0XdIq3upUfU5H4UBbH/4jLQP2nNPfJCKzsgF0qUXs6THvN7
BM/MC8See6C9QUmjiQAEYge2h94Ew5Hybx7uW7t6sJSUpBOBGiw9sc0q9Qveg70FTMlCsCmj4zJt
+Abh3ROhdtNomhPELZzJyWKz+QrDqtcFcOSeAgIJ3EMhiABiIqevjqQDKHUqN3R+tz3dwRnXiGHu
spg0ca3X0hrU7Ho9H9uERk9l1f2FsCfECG5RFOHOMdOqJRu+LFyYKAzDzocm0gB2lo5wuRP5TU3c
SSDa6oppMg+Nv28zC2WRqzQDZxvBgiFaR3MnoqbaJtZ8ZRQaUanRPvdmlaEm+xcSNQygfIu/Tb6D
RUivXHmuo1jw81jj9XCHyGwpzw7XbwCodPIGOYYqjGJwfbRfL5Rjyp36CjauxOmj59RcdwiLXCge
AdyQHefSqFqhhBeEbOqWkMMtfeZQS5ER1zrx4RoR1YQHzujnswvgxbtm8XHm0fQAcRWycGqSUmth
K0A6HLK4xNeHcn7Gc/X/Od5uLopVr1yMWsT3XT8OxfdvJMrlJUavkITRUPOlPRQ268nTartBVk0p
jv482BGL8YXbLkhgvctj46LmtVqo8okYKsJL9F6FQO0w5mPvJwOtlf0LTWJRMgE2HvyliPCge21Y
teKCPQ2lQra/tFJKqJ5ntxbQwWzW7LYpccsNqodEENpdy+zVH4GbBsODUZimGgV9tdxRMCMOP6n3
DUHznwPXCwQLLwxMx7JJqGPKbyk5taYlvkQHYkpro0SvkOT+SXsNfaQXs2NF150isVxC8Nz6QE67
lbNE7XGrzUP1Ya20jxWovXCs8jmV//mmN3y2XJisZ5clnEqExRaCJ8av5dxjiYctCUccKTKJ4rpx
PCLXWV/10fEyrsTggzLureCCtEQ3A3tySYMmM2C+BBhe/y/T/y9WAEqtGfl+1x8N90u7LTr1Ri2s
/AVRD9fm3yS0wsHfpzJDHGFqk0d94tPE8pRIFD6QvlUCczLNyxtAKs1vT89o/FiQFhCrtQQKSrXa
RvkNIwsF7q7u5f0kMlTnbIDforYyv753usjL1WhLfWGnoY5+hc1u45vUktUtdPZXFf2IYq/39tpt
nvFOYDETiSQoMe0tXnqhzmWxxPHzQ3C91Sf1GlpyU0xQ6HooEdOkLea1+jGHtiRVlfI7cG54tPXS
dyWv2UtC0xSo+biwBnyIw4VQ/UK8fz9CgD0bgoeoExjDYPf90QwLnFaI5Rrh28xieXCdOTzkVhhR
T4V/C1a5Py2tbGEATrKYT/mggwSZcfQiS32EeKvOFPGZD1VEX3a42WCJC2TJhPVKr/ou+Hymi8Jc
xf7tYies4vamacCcet9oQA3cVvhdT6cT7W4I7wscBkcjEBNzihgUtJWhZy34sxO6WInJRhREXQNJ
o8ZjRGTd45oEocCrSuIm+gmAtr8NVa/5jeQo/1tBXSYqb0cHTHvpvHUPuO/PWE7aNGWnhY/NfmNT
uZMF0gts8n3eOSRGf0tNT9N2BmBv9sDiW5isOAal1MDgzU5clsgcsX8xoPw6pN/vST+6vfCRcmwf
IMM5H7043dGRNN7mXrya8C8Yoif4BGy4qtxGlOsWnhg5hTWiQY+6Pxf8SG50MGPtpfShzSrBV0S7
w+3rfzMMEY47IpCu+IsjL4Hux6lCHKoLRtqJ6y6meyHatX+whPKdiwOEVt0UZnOuv27hLXgZN3Su
CshFSPlJy9SDSpjZsT83QuSaPg5/kPhwQZZXxW583NPjXdwl3caT+MHQbzN27sH6qKrHY5v7xxkH
mVuAMhBX1HCIXFc8IjAPAIC70dozuaThXyRkLFWZ3oeX5UodY3VcMAKFP6srTBEplLtYNEnMCTNj
jrHa1s93RB89Q5yJjc8ecYM9BEvM9jiZPWKl9VWrv89b0B1mQhLnQZjbi4A+f3yTIhendW1Xwkox
imwU3tDkExg0fI60BvJCmksl8+BCrAom+bC5cSch0agEFR7inn/Ue5BCa2WG0EoCuYOfI5mosRwv
QA7G+/Onf5pW2QnUDL8SK44eHbwBQvDH0Su2HiwFHXsxGl4zpT8FeaX5m7XOObGiHExtpiPsYzjL
WatixUWZnT2XPG0x+OSMa0pY4U82kXUp7j8Nz8J3C7UBm4NNKwTkMFD06kRYOgOLbRU5fQJmMWrn
xTgiAbOdapWEEmAiQPIIJV5L4yT09L+NakdSLyjlRf06aj1qHpJ7G64KDUtoqcWh7JzM92CrJ0F5
HAquu5f0XaeOlm2Gx9dVY3M8wK32+YeqffzbxIFqVktYAdZKpabB8x+/eB+4ksWjrKi8jkE8kDNo
iMgtiIHMe5i9R+b+l73g2Wf8uq9l5V3ssy/kTGkNzjpPv3NkvZ8YttpSqre5J6Vkn8KKwb+w712y
T5UIUfqOOTRTv7xSlF9sxikuqj8cZpY56iVDlBpyVDiDNJi6lBGrPYmUHTvWIcRNrX1sX+4lSZq/
szMwpyHeIi7uiHPGxlixfQlQK7BalcsKKYtZiTjsabhbS/dM4i1eRKveOmQ/yDdGN0N0/hTFMYCl
uW7I3UN2Q74YHsFYWE3ssApD6JOQaFPkkw4KYT2DsqeMOjdunhpKoSpgmcqf/NyRoYaec1bBzqGo
kFbthEUDMABaiAx8qjVqR/73OYrojdkdI7jU49n5EEg7oYWVRSv2nrbxyz7egc9zvJIrIV+mdy3n
zNFgDAHQBVJXBshxNlCIF9o8qp67pMrC1I/gsU5g8mufz0JX/hJXAgvPibAgUr4ThtlkzBJyqcth
ZZ5T8w8bl/NzYOabyr7aCw73MdUpa74bmv2WIjelaCgbhh2JsBfPcUZA7MkfWMcRD+wqOjV0F969
84UsxmW3fuurGIwMn6Ccohk9BPNQZt9MzQT3UONXDtxQnd1UqM5Ovhyxh/f/sybthEC91aeS0IDo
71kWE6IF7VB9HePn4DctDVO0s69YMuAdgLroUHMsAxuIZcCbUulRyE++f0Y13H5Wu0DFlYAawj96
WXIzFnS/GO0coKvsItPBmld6mGbTyAFjsUtagQWTiB9JpClL92H6wHbONrOFbBFVeTfbMq/r/Wso
aYh2PDuNBToADXBCZbDFAzCN8uqt4Yz9KXN63EAZEUl/arA14zVQZU5P0RhgHzXHPzSIwT7o+IZP
5xWhLALi3TALRwad+wiInVjQ0zWCdlbx76RQuq5zY6LkbvOk+jTG7CjRQ8UdzNpqXkWoQxAeJIqR
uOwdm9SnCD7UOCZ3AsVpU0DCRtS8TLG5Yh3UfMrN3jiCMEm0Tr4A6APGAXIASFmc08oMeHI1iDkS
IYLoiah+BnjxRmpEi1n73RaG0oqICp5+Um1taVcTR+AFtjLqIQiEE0hG13vLs+KwWleJYDYl5frA
xnUSgbvyMNH6rKZS3EPiKOHtZ9ayZBIJaYjkuoAx1qofwt4jWPXk78PSJkNK09ntlziXiQt2FnQO
Bo7bLdveyu+l+6NbbB6CaLSDJ170mD9zQ85gTfUEGtQKoQgCCE62Fbw5WBlpTUQmC76ZtyCOkSse
lLgOygRLDF24uW4XebMWwFhRTPwjTSipWuaKIAX7N+zS4TwL8hfFQ4/BrzwI//GCS3vFXPc436JA
Fji0IuRl6ip6uSC/dMDWkbpE1daQJLs4VV3gUCAgTWJW5G2eqA2pNx8wNHSIoxVQaHd2WpbmgBCd
LQF+QQb0iFiuy4UoVllLXD1zvSgahsnC1rM8+ou3wqwZZ1XQ7iRGrLUEprG+ZtTLlEznXRyo0DvM
5+cv9CcMxQcjU96FC5Xk7wTsc3aJjJMivn3kk/RpZgO34gfh49ZE9UNn/UKPF0TsQ/Nz16Z7nBBd
shjVWprLNKG32WN+/8RARR9Iyx8P6bG6qvjxTk4VzOmeqAivI67DUsiznxqQw1DSEc4v8sdAoDXs
r4VShXTJL3Kz3Nw+5lpu4MBFCsdg/MYwtS9W5w3+mh9BFPWJ9VLoTP3ouxh4odaHLrZyoH/vEnDg
nA7WvkhcC8ejc1/yk9MOAEcCyczlznP7gLaEipCyeF5ViBA7RlfcBYasfjzD9cYANfcNrW55Cs3N
bTb4SYe6qnRC8nA2fCS0qsnztcw+LADp5Buf7SS8xyTcn8YFbyVCqXMUn8HAjylpkDW20pWNgx4z
eSTO4otXo5mK4KMdvUM90nX4Wdo0hkf4r/pR9iRiNV0roV5oR1E3vTPxAQg7evdGwY+tHTlC7JMC
A50usO25rsCV1njBu1MAABTZ6rHVLjL9DsM265h9OT7usEbJwlxcCZE728yhlhnmjZHdERZhoJ3s
rN4wRL3+0eX54tzf97mfUWi72ZzF1wxwYlH7yBmsL26RcKIdNZokg0D7Ud1hQcNdgsrbUbazdq0I
ZchBYk26UHxOFmI1oVV57i5IsK4pKdc6CObcKA8SKFYka/p3UoPW9ni17PcAZVlzU0LZnZ/U0etQ
Lqw2wdTLfiL+SgeUsMzRqXwGEqVLijz8CwujKIZ1IV1y02kgoSsyMn0LV+IpnKITzLFnoAZceFMS
zMOlNug6RlYuB5RL8LFu6OOjxHMmGAgol+S6EE02QWH4hkHvaydySHfGPO8BBYMIW0dJDBXr8BWq
spBad60Z3Q4jyraWZ9ZfR6rk2/VPvSMRujb/BANsAbcq/RDxl2vrMcQ9L6T3uGjpznBustyHsTFk
yqOBed7vxwKs7zbO4XL2mrk+WWJFFzH6zmZitYLbZ6/1Vw5CA9K1kzcMwwhCfVIpZprgnGmjgKN1
zF+IBO8TMuksGder/WW+VFsQTZehSjxtcR7UrBOUctcO/5lNxPn9kc/YlWi2AmSFBJKDmjvZVN60
T8xVwv+7v2+4Hg3LUJEGGf4h5HNsrR0LBVZaFyVLQFREkXAvbKz9gNtK8wWyE8SQzkN0rkrTN4Ex
IUeTogBQx/GMCNm1TzoiHnQmJ9h9g0Y2+O11YsD6wmL26LaTCk2EkHF//YF6R5yjWIYzgmdnA772
BBT1QFXEXErUPXoEjYLydAhaHgErz0SotHOccUlOoFyCVQlVv3c27viWWK8SjZ6spw0Kyf64Y8YE
w8hsVyTe1scOXpV+sQok9uO55GQxBDRH+xj72jo7omoNXN+1EozgHhzP9D1s+GGmT/QauU/UjO3A
9wcQpTii40Q680X/MKRdEaI24UgoICyxIZvFOI/K6Fpf6XTkVVf/nsw4mBE3/DwxTeSWfG9rnCid
EEoF2/rTIXdgDCtDAtjNU5HfXY8CfKdkktcMWKl4iSW61ay3mWsKz5/Jg/MD4F8QcQCDjyWB10eQ
quTtJokZaYqSIvp2nWhqv9ENSHbuZeIlvXl1ByJqKLBZMwdJfrfOsmJXUxD8CoMglZqmarQObdCe
8PFEZfOA3F5UfgTmAlj/+5T5YhETbSYCaRv2hpJJznXbqH8vBAHNPqNLmQLww0LCZnMDbhq4iYtZ
5JoqudrqmgXGWe/P71Bn3PFLc8vpiANMc6iT6jQUIsVvZ8O5o2XU2fgPDY+D9jph1TKUKatciiyK
JCD5+WhQ/H6viSJJlkpKaw7Cea1j/prYxFJEAcqz7M8KJMhWy6KWzBoDSml6S39awTGUZySR0rSS
LY+ryg/wmw/uEVqqYizQ5IZ/b9wPak2dJrzEa4L4xFcHnhB/OYfrL66rHR/Qpv9v6msw3p9Jzudh
yQWeZHufCQa+hxCOK1DHYzRSyh8UMM28cmb1EqrMsZQuexG/9Yz2ueZfc0MgE3cdkNIYdvUokZ/Z
wGWhOmiIhIUGIOU9XZJgMCn/upRCXFkjLtS1FeTI/xZzIEOqA0hS3aA/j5KXTvRnJ4zgtLYyW6Za
g+c0Rb2ft8PwoYe8LYlx9h2TgUJj7FV0bWn6a5Axsv9uOoDrJJdBv0Yd5imEmoVqdlhk5wOHhYyH
s00/gc2xR9hUPHON1D0Oi/yS/ZPXdNmkrDKQzr15/969bRB0OgCefjZPiRSylypGp3PD5Kfyhu4t
rTdgQ1jpH4PUsyGYHF81XP7Yr8tSXwU2hen+KfY/scrJQPja268ERKpZVLqOKcTvqRzSNUECdLGr
6wOqT76jbzVDCqFe3mTJ4sS1VTQrkJXpOYRjpyty4a6thrRBMh+kaUdcaMmx4ukYet7BzUhw98iL
y0M0puOqNkVqGbxS/GmmYv97L9ao/W4J6H0C74bHL0A6jXMkyEOuZbpLZgJHFkAQtLLTdK2Cgdmf
okEsOJTkx5JuGp7l1gi5O/sLmYdBQGM2wpmvdRDR7T13o8OBjn74lI7oAi/8IgaC4pMSh2lPiGCn
OiOh3cyUMG6xfHYl/0GyQLN3PO9gq4Jtg9LSI/4h+BbjHENaMXQeqM6UGdcIMKr2pbLNYPGCp+So
/PPB13ya+bv/SFaqqIh8iV7rRWkhxpFfqU9+Y79tR/DsqQ7UP0kzpX8Erug5rj4NAXCyhhMXw4Xy
ZtsdK+oSMUJTvwkXSa2/x+okYAWyrr36gRU+8zlapRpj7p1zma6blwYZolmyjL67CAmmWVLXQG+v
yjEt/3h7YxXbUYPYdvYyYLjJvZhrIQnTDwlRQ9vnlskzdXYWugBoXkbieUtniL/xSsmwG4COntPL
Ts1s03DAly6EY/2KSKxF7ZLKwKHE462FNG4DAOdzTUCZ52HgJMZI6BLNNfhWYWMGuPdoCUx6U2XP
Lfh+fSxpvjvzpsf6D2KR0vg8xaHl06vpc+8LdZBfavX2Myvo5pywJzU9QuOgKAJrps3+y/C/aogL
IwbDFpkUkwE97Gtu0c1vSQRP1SV+YjabluSWICAQ2s957xf2nX6Z3Ict96ApU8aEvmoj8/mcehae
UcrBzKQsRldm5Vjg8a9KU4irbPAi0YEoCiAU5JNK7cQ5In8Z7dh+8aIm9CofkNWIbRO1TcMk+UMl
ZCFzp481BMxiVZSnh00nzh4Y1+BDAFJQEGQGgf46adnK5b1TMQuFqAqXPnv2wBcuKplLYGI7XH8Y
ginhmKB6S+zlTpNA164W++pkOR4qbioDCIj+a7sDdMfDsE7uKTYyS1f4DLXbOijQG3fNy/MZdqLy
po4QQj13RLwnD6P5A46xBvVYVSuIOI2KE/Wrlm9tBlnXzguyvVKnp2MxH3pX6lNtpEEEGUoRti3+
SgFwRSoBnvnYGAcf/f8cnRoB1yZ9SMfSUOtPGjjzmAPhNRD7bBkJbRPwW2c61+wfSmEGnVeh6qJm
UfHy4PKVTT6MNgUrdrfUAGdWkbFpKTnROjpYJY88GyhYal8lSmzQlFWp0hOLgNXiHi7TQQ9d88DS
cdSslc3ZE02zxSaCbKheWq0s7CEzkpEBil9rWvqqWIE5fQiQF5O8dNbY1pD5l72V2RZ0AYeMRL7x
T3IssvmdxigJnBIBGYeQLdK3Cr+uua2qCfY0UzGrU/XoXIEc9KhIUFobfoEm3yLgSxb+4fRa3HP3
PD8/F/T8GldSQlcxo9ZKE9n0kmTGFTGVIlVitTBXqX63Kxu/jq0ou8O/IMNFnsAzB5KY56g66dS3
eBB8AWR/ZJF2TUHzjRAb6O47iZihdI1mYBugsh9uKNL17huBTRIN2hDrQpOxH2IGz/NSAISMCny2
2rbfxUFoUzgDCWlWv6dt4AwPcR/m0foiBJRK4e8iaPW9xw30PNdARLmK4/XuALO9WX3ViPnLg1WF
62KYnt5No3zEXISJvDO/f5jlxj0Qwa5C0/mFAbLXxcI3Mgno0ULOwhvubhtoHi+D8giRFObOnjiW
AmFu3H4zss606b4k40jE7MMStaF797iEaGJmp9H31FOIOCmLbvn9mVUe77WZIfaXPWUyl35VAL3q
e+yr4Ra5x3jGiT8Bc7bCz1NKSlq6Fv1ca2PyuHp8+VqUlVedGZx740PNZdlX8vIXQ8vY+PZJeO89
B5vFkPaYmDStDrJctgrfcoBSwdouwFgbO4ALzGBbRhM3bG9x3lb28gYKn2jKh4YuhN0ZedOdoanB
kgJLH944UKlVjudgaDXfmXqdvXkmWMWUTLVaZf2/oYx4saDGs3PJ2OPZCI8VgqtHhoWFYBV+s7J4
B2Wb171Bt9P6JCPnjZ9oGXLzOdmm/FV8cDAtO0nLCvcWUwYWUtTk1hNF5vwuSry4C6+oFFsbkLUN
yCCbBmoxHWn0W3AKc1vezSABNy7kbuvRhnNupqe5mIBBY0/qV3z43D8PuqPUcHyeywvBj7RhdaB9
jqHHsjJXxtEuCPB39MF0dQZkih9SmHD22e5KF6zwPfHkjtM3F9+PUgBsirSRUTMQYmhkPrBWwJxp
NHuM6c5Brpl2ixn77Y0rH0U+zb9NunYLRuzakDF+GXWhZT/P3YGltpfRBfgbDlkwThbKu+MGqlhl
FiyEP2rZ9JoWpjjJU/VYol5Pj1aBnlOrTUUQlH3FJE5gfOy/vn7hg2DwYlWQTNldkUQzh9nvb2aM
9KPLYB5TPZY1Vdyuq7yU0v3ZyT3RI8AQSWnCds/Y4ekC9P5kY7wRh1kTbMuBnVFJ0zlSPP2htgf2
+/pQvfa92csWPtaqielAZrPGFKUjCtHrDAbXB1aq6mCEn9rw/PKg7gR6RWyS84Y/WhqEPoc2YNue
xSZASM05gSPt1gUxBbcP7AiDrL2UgyjIFHQhEHBBZqUH+Ga4pGjMd/5IOsK3NjLNulkAN5F1rRZk
oiOLAkR/54FAhzQC9HBZYLdwxdwvL4xJiqeCuDO38/R+a+5fCOvN1FIJjbG9CVFkZnZB5JNVnL2m
fcs3KMP55ugYcxe0OhQrueAg4B84URAY5u3JV2r4UGug/wja6F2ZknYNIzqlVUoiSTidudWY20Ya
QzeDFnbE2/8BM6+u47UY4OXfBSlaEQaZCjnD+olfiKFtBcJhrNM6R8Bf1bFLirmhFNzzqHUrNKBw
vYZG9M4mHcSwJn9nZyPDahUeCOlrO7FjpRceDRfF7485V9UJQJH1DbhI1d1dCyvlGvtAvi44DmDd
qyPzpv+wZDlu07jNr0XhvT72usnY+f64GyvCo7WuPE09iYx03qKGUeULhjR+CAKb4vcBPxteLMRI
Defh/VscnzSN0uhGCDL5oW07GVmxbGPDjCkt/0sVubwlsmxa6RtzEJygcY0d4BBOtzQAwduGdQLx
0NUSNwWxotAxWY/6CT5URFCrVPqiVC8ADloGwiwJyRmc6aFtzk9nlV89FUcWiDj1+n/AejKhKt4D
6T3gG3y0p0ascLEYXmk5QmOui4mt96AyGajuBIOpJLooW1nB1VFbzw+7iHNZjTJv0p4TTtka6wnw
cMOzi2uUwOvXKqhae/gbGufsYvzliCvZmJqGOcdpih2u4jDHNAmkwNKCabPAYplMtLx5ksPPC9iJ
PdM7OXoPdzWWT1kW0JBhMPC+gBTqGoSLsN+pB57H6xvsIA77olb8RyWgoRs1Q0mgrqCWDtd2MWVj
+S6QWyg1Yeq36bHSior3tV6tu+wTIPxoY1dyZpClfaGpBR8VhuyRCKEMEnh88oRrMk+DfIQGg+HD
in8Pmmdm6/47HFKNQF/fi7jecg5Pu5o8htbgNEqeN9oFSWhmdsujrAMBtpxtji4BQAMV3cClD+0m
aWUhwKk06skp+nleCndLLDxhCZjNN5qjtrjIMV0+y84cx8gIZEupbGuxv63Ln7EU3tUMCV7heZRb
9i6C3cyGzQjHhtuemmDAV2L0YaSKM/QDMuALdMssa4sLZyFfY72HVxBYZBueh0QinCLYa/ZJYZak
gr5SUGwntpI/o0wTaXsBiZerjbpb9/Q5KDz0hTmG6RgmI4IhoUlxNrkhcox/VvnZDExQ4uigyV7L
5qgkkcneZ4sFhzWPY2wBSdfnrmvLCekgADpPz4L+MyXrNhkrNrT+Afq22TjR/T6QJ7Ea4pan+zej
siZudBWr7f2305PjS4d5LwtuC80sKhw5ICNE9XqigxP/SSmSTyp6S4p+Q5J7hX469mF+WAl1q7tf
Kij2QYObfunupTDOwu9oo5RmjJ8FGKpJUOrOnYD/iEwYb8zUiMEoX0+OXB++ZMO31MaaD/sp8nLq
V+1M2hU+4w+1/imGoGpR0jMAU5pggX/Ubg/Y9gXHqqFxEsF46eeydy3L+el3c2AiZ3lRYYWPHrVu
SddNfUmlzQy9S1LDQ7YDhq/MpIJst0uhWeKBTO2gXc1m06aoWQOqb6ySPb9ML90xHW6OCxdmYmah
Vz26pvmwLbNL/S6DDYuC9/i4X4zugIaAgrwzpKxP248QMPBQpdlOWKcK6sp70y4y57R/YnzxQjON
xJJEsJgqMzPfQhAWAOtsIbX7Yw98RppztACp9pfJvb+yA8Uwwnd61jWk+tKKq6mKbDBplSquSWBH
vDD3DKCd0iD+dM6f6rWSfstOJRGRssOODYC2YgtpYvPt8HTiHM72MB5zpo1cVTLulzIBzBLWNauZ
ct07sbuZ77cX4x1+95I+ZBH8mfNTKhkqaDg1LWfPlRq/iui3A3+ubFkRzpJ+IJC2MII9AosOyTFo
37uIyUfndpXmi6H3TVTKSTDfvkrSx7wsO14zvozWTKfMwG8AMwRr+AwuXch03uaLnILqwQS8OrkF
I9JbRvhdS15g0eOJEUkB2tU59n50y/+De4aTZIwsAktHoVM2zPhazmMaf5sn5EcVnxv6RgqPe6HU
qtG6eXQw4n9/dOnPQs+arWCX6DEvfSHUGt6l4sc7d9pclzz3SB+b3Tzw3PaI9wdk/G7K6Ve3zz7L
LWIHIY/sltu6LF8ghXhjobIWui6vjPbiZZvZoa7N1brl+rjykMmtb3Rl/FfgcS71IwTQ78i/bQHh
hie1b0UmzxxY2CtSkpc1u66+66LuC9XecSXUtHfmPkOesl60bZcO6brY7j3aVOJf7ObjIuzg6lpA
E4x0YH4ht1dsL0rEHtCoH2Ej2bTOJQk/J5pmcOhDEJGuK4wOCeopSmpixapHHT6y4+Qvvyut8bR9
Wb9SG+qRFYiKPLMnYRoDR+Xyy5gxL7DRJ4Af+wITFaSOWTwN4YlnzH6xhopv0K/rG1GWKvZTxIoV
fB9qma6Iv++HOn/Lfkdo6dlOB6/rjqZuOTzhRI1VMsSSPS0imY/ImI+C45WxsKqTUj1nStDwK5bp
T2SMVRhF6XsEMgl2MLqrV4/JELWXcwfb4wNMG8vD1pUjNXeVs7HorxK3miIpS9X5p3VADjbQfL3h
kZEDoMbxAsy23lKpS4JokQ1PGxUvN5aN93pH73cvjE1xChNY7AAth4pSsTiPGUao43n+r54SuUFH
OaRCItB0TwD1BVtzbLpF/oKcy7VIM7r1XswsIL8r9uxcEXko9iAU3wcyMGDNMzJWr2ohF3dDpX+c
KXGjnwUydFzZclf5I9BhNuKGJ6rkUD/jygziGRypQ0zRgAIGJBAVmXmRM5KEwQleZYq2ozk/gmTg
sOLXjvyCRty5f+JxoBcfijUTB3cBImDv0KaoSBqlG8VjGdyXz1fQ+UaBqy/R2z8LOqnTm5jrp23q
KXoA9iehlMYmNa/CO9URxkaq6gndz7MXUtFeEvLQ5lRPKLm6FNGIuZf7HRtXZBGqGb15LMRzRein
Zx3iaMw2qutkoEp+zaou67zXD4cbDqU4T5Yelhgg8cbpPw31P8nNZmkHTmF/O3KHY40vRQiSbSMe
VZ2uPzrltwfrBW294pP6NQ77qc88SclPs4Xy1314XcuC0xJYsdWoYPzB+cQSMrjZUHESsUTiAF0m
3lHDMlYQDSGlMP/0fItvBDhK61KMoKrp8y+9IAweJx/PE94ZuUyM9qHAfBYhqyIEizp/AtMYXGe3
EeMNIiafvO8OE+wTkCc0QIjTXn/dvVpJfS8J9DDUK/VCHbXI9ePemT5dBfhUVVaoZMOzwxVKs6Mu
5TJA7OgiAy1KlfH8a0odSn3Jb2MLo7iDHuooAn9rAOBP57UcyW545l/yL6rWoHTbKHwmczzwnXhQ
xrB2qYc9mIcoZpPL7ZHpRsLITVaKN+eBeCfNmiCF3QzNbmVbc6kssvTRxbBNQ+nB/ZBxs1yZzH9L
qSZ3TruRRHdYyvOZgorQc22dzvlnx9f6VnEEiw33K9vYo3MK5gFo7DgiTOdky/JtWROIXJAL5uih
+ChdQfUWgPWxpT6OqvCk6YllmJwnbkGHjIAlv1GVtfCnEP6EVo9oCSAeKxpKcX7iYfFWRYtrZMNh
afSibgvOU2DNZF1BH1fYwoVOD3WGUFu7bzB5GjSIpZArBmisd/kL9TZCwjhtbZ7CsB+jtmwg68FY
ASRNR+gGkHL8tSqPnuM+8rpVkOgmmwUGdVmYdwMllULlpuNcfdTavQGgj7tJ+1qnFUpTA0pGZDCp
eSHVeRu0D9OZk54yhf36FQNTKbIfmvr2+PqGxcxr8BxVXO7eTLCEljbvqVQjewbc/h6CQw4j2ti1
tPV4SPMcce+mC9ASLFgdnNGHgc2yjYW4dtZpPH+Chye7oh9Ul3yjRphme6UKSisWX9BsxoA7mm2n
hK93aWPYuimdABccbTDEEwLZBSLxWiKVmL1uCp0izXvtuktfolhKyFrk3zLwGOnRlkR/7tRED7Sp
iENcpdqp+dsbX7dhVJ8t6yIA5KF/VLwO1rVAK/WhZv0+p626RNhGWIN1Yp4byCp+uylNZCmyTjts
yJyP+3lM/SanecN0LMP+yXLXo7NRn0pesL4VAAhn55BUfpU5b7LcZM5N+bdXUCvqvY7BvBwYO3iz
1FOeIAFksKvOYh3dYVfuSSIcZv19LGNOP7fedaWQ6TwB/k67Q3DYPkZbSrs4Sng9boN3iSzciaW3
KQX4MT4rO/kglwjEF+dbXYo6SuTMuIpih92wJVGsOM8rRFsXcz/p+dS4YbtVv2Jnss+QXTPdKXuq
MnEdvT+aN8gjNsKlwJv8GDPR7jrO9rIDcRXpWNbmiCPLzLaBlnpB66KEhIUtI3a9TGc0A+/z2/Od
QIb2UrBdVxZtZlXvoNxozCRe+qvpRhKX+n1v2oCAvvRPOc4mj4FKnpFSwwjVhtmFwZ+/5Bd6xzE6
L9TDy963WpUacUBniQFXIeaPUp3g0jfkWQfr3u2XdwuB6zeVHuDMQM4K/vP8fC/Fbk4ESBHB9opF
0Bp9EVrjTS0aa9uW586kvsL70ipo9u3FpUibg8Vxh9lMynw0g+weRxdecjUKu5BHOpOdUWms7Wm6
bTP/fX+slnPbKHiRh2BXSvD5CeLEACQzvL9o0JySNRTaqIHzsIoWvdq+ax8H6FVnft7RG4CRMNZd
k1EjPP+BD1XLXksOs+lwAFXEd+cvQE3g1Ohqx7BYA7gW56D5wioY/5UXr8i5TNCefVM7dkx8mmg0
0pCera0g6XVcdgqHsNHXVFwFabYPI1wiatkccNI8OeLaxFG/CMvtxwOV7LrxtO0XeBAc+UMKmaLO
cD2uRFTSWSgkkpo9TAPPLV/iY6/EuZWvs8VJKfImNpqz5ei7UsCNz+EI1gxweyVv2l5/JY0N/D1r
+MWA3iyWO5SCHQ/tV3CQIPvKtUxnCvXaQ0S3cu5l5yyL9/BXoany6LAGrdxkYafPFlccLYadXgnp
LD3fw2gJhFup8NaX3X2pyLvTFyb+4iK2/vqUgYXGTufIretPKqCx+l5SMCCKmU/KeOZ/rpGGCYNW
8vP62OQYuLzMuy2xmH/MM8vWXy2WcVJv+DTn4oT33wFICwRPI0H41whrRmxXlBk7nWS9TZ5daTS6
0IQXCdLP2ZMO8yZAtS10i6IjgkA7BcxUMvP/eP7SNwNtAmp0aV8GUf2xxepGrrxNSNDfAIanmmWU
uRhMYmdUsf2TvRDiqrq6wBe/+G7VcrJ1Qu2r2NrElkEBPCcVk27Iq3QyNH7/SVT0fbs7DMYc+dSZ
Oev9XGhXnMjSnbm5z4h4rOScLiLxRAVVLlNJCrYfRf+vDU4VTTb+vSe+aqhUrhtmy7ORgfG7u/HF
sFlQpNC2nHKlmg+KLZm3ckukekrivPMrtRSN37hPzTVJ+8lGQcyu9phJdhiGofhH88IAdxCFD9ze
xDWTC7J73600jdcALVCCrTCt1wIg9OGNJFtslP0j2x/su/jXJIJk7Uxu9w89kpoDCoPZTLNby0WP
bl6pnTfZfvFAHHuq1UTcjFnICwtTHUvHfQ6KoQdxzuvCfVr5ctcZjjYQvzKU4Jq6J3DMlC/LvWAg
iW0NltolEdt+fa38blyLuqKlNIHenngs62K5RXKI61tkkFSDFV9z8lO/nrGiPEVPRhkUXajYSpqs
OcAzftyIltYpPlC9ualXAKqgD/blj4WtC/v0nULxros+MaErsZA6zjuPjLLNiONEwyvFLE1eWtIs
bzFwS0SuYVXTVFD4rMJ05zAssMkbfLqGmORcW02gJKeQc+gtnUkAqX4iINXkuMWnmjW0NOrPyCmk
f1Y4BdB4nmbU5vzdfa1KVkXgOGAsMV5F2EigVK9/amitkROGU8AuDV6kKDjrefBq7NF9uYqHISkJ
JMlGgXHV0cmpH54xCmaQs0Vi2wsSu5A9rcv9//8CGoKM97dIlh4byG0OTwyjFJr3ft/t7UlK4dVR
s+dx3cKexkm+4yq8ffuyUCHJ4SGe4N9FFICJT3pl9Vd8lLOFjk7B5ubbyfLRppePc2iFJhAtXbtD
w60iMORHQVXCxubKEWnwiWIls7aqaSHWQkasB+YdR/xzRNYRWSLia9DxN08NpBSowJVAe9ppym+s
vKa093/ULENEatxWeQl8l4hLCcNqeLdEpSUdj7aBsfOu9Pq8FzPqIdeGHR8NOCPrQnzVWvejfmOu
iK3iceV1AftWweADNYsh3Gc3XxM+nKYpzpekQ2iDKMRdOFJjsNux1HiQl7m0mmzcerZihbf5KSbC
pOdKPQFafgHibjOnf8W/bpTyhiGyE0IfHhoMXDdgImEtI9cqVnjZuv35Rh2yM70nO5YBm+sMrDj6
3OpK++/4Bt4aXcmI5QXElzFxX3qaVH2N452uVf/W/lQFq9jnJMA03RmMACRTb9YE382W8ky6VGsq
hXg+PxEkXh9lpbKe3HZb8bzMDMLuti/EEfZYbgZxFTcczP2qM30Z6AkIC3wEniflm4DxJLkaZOqV
rBQM0a3BTevh29xm/brXk/mUA8xnE9B+HvIC7H3Vt8CvWGOFOGlbHpZ1C05zLqKJWd+pB27w9/2g
Xi5LxeJQPzAtds675+hu/uPDnVhdgQ/A/l/MA/M10qEZWrE1TjA1vtHUJHz4sSseCYTUf4mXg+9r
g9QFkACrA+axAxBiLZR2HZIxEaa8iZKDbXfLrFAwkFNj7Y/jiA0ccpwWe4NumG6AUDexWT8SXRYt
mYvkhANzWXXen3rIxldDzIRPwykP7GRga7LT7wjUA1vWG8d0AwWvXBXsq/uu4iF4Zdfcmm6Z5ZS+
AsbopZybLBzg9TvZjQ67AAeBzDp+7tiqM5aAkXrrnT/ARSHgMmBzrXGVjeHa/B0RkxepwK7AxdEs
hE8KCGT8LKu2ainOAoMYbQCBEvCRhKgeb+7kEVUcASDHzN5YMJcwlnhnwgQOUQvegKG1Je8XncdN
DIjN+xMZQZZow6SCJQiWLYUZajgm3T/pRewLu+Ut9L2yd7ByafJIJsLeBML6DoZKhjHv7FziT2Gq
plBWUQw23X05b1PmKGVOzXNuw2E4ld3R6hvxGDcjPe/YFehTvPw0ygEDBc14vW7ljTpW3NmH4TVF
7Ee6aOpKfK3OwbuHNJ35mvS1BAXTKo9uaoLVLLEYefGPPuJl0vNhy+ecp2hfKrBuaKh9yxY3OmTT
IOYj6PwYRDjB1GS6/iY6Pt5+1z0AwNT2eyeBYGeSPWPBSX4600/3MZw8T3TXEVnU2UQ/ys/UEImi
CKwT/87rgmhZiFQhnGQJgVRqSPGY+iiIWAIifqgEV4aYWBnr6nXcLJd6SiS3VnoRmTPxZ4ZqFYuZ
4dMFRosiRJfclAMtxJiSMVNxqc/UBR0yP/LK3bLp3X1s0R81YEY6t1LlnquIt+j30V6t2z4OLe9+
dLoXIqmo0n4e7TT4dszpxC/Y6hW5HWuSgNdrXsATqL4qjlhHDnSeVoMpB/Z+6mocjd/58AAdq0q1
TfZHNGHnsK40+8nngSyQGRZXu6X6oBcoOj5wlwMMB3Nlfqk6gfHiri4Yw1lCmrj4UmYIvmdzV9QZ
RTOi1hdm45G+eqK7TnSrIhuTRkXi9yuxNz0+PNDjOBYnui4Y/peJHucBXUptEZKaLHj2xHiLuOIP
9/JNPS6o1ts9G7DL/+IYW3dQSxZJHCcGSGDYGOmexWBcSMF1GH4nAIde2zswyVeMXDOC7bTfMLUd
lj3csT1QgxfOkZb59MmDNXcNDnYq1LpoHZyrlo/lJCPcd08p3090hVdIvZwMdft442JEsnXA9vCk
klYhAP3+lEehx+KN5H+6VJjXOHE2AcqqRv2qYRwGcvhhFB2/5cXw78ilSC41kfDKuGgMd/JN6xuZ
e5ajY/6DSkF3ygxIyc0UkS0LOf6zheXTIQB1XIJNm5EPKbc6ZUOIJpDFvzVcE/h8Szw6TxYxxDv0
8eOD2VvDNLS1cJrKOtjF6lypoJaGx6xo0WsinhlPDa4z+sxdXRcvzxARLAZzSTHf7w04BMLBqTEA
gTtb6gPpWgVhwwMkynavlBRd22u4sHV25xdJP3ydUXQowCCFTvohCge97k0pk5j0P3yliaorL62/
dFF07LjUgVs4S2E3h8zAzJhpj2xCfTqH9zz1WvdjWjPJBhirlubN67VlFHGXV6RwRxU/6heGQf4T
UAFOd47qj8vbW/8UPREfEbmbyRfKbxkhgUkRcOXgGAvtUewvEcEgPv9lOM1gljv2sjYdQwEHT+8P
rDHcQ0aHXAtlMTO8GarEsP7rbqqndezdG0q8F73InoZiSbSgjHt5e/UtA6F3FWIkL2bRwjGoyQ4t
CYUzuYDwkCNN1l064DG3mcRMWzqD6LZ1j7NLLIhZmTm/+z//r9RKcEqXUDZ7LYgZmdzgFCBQPxYW
qnjgnLqUS03gsNeaUyjoMED8NuWrq6O8z7IFZG98qQ4JVFpcuWAR2AD1un4ZG6vMDzXtihBy/Rb3
mSlNV2/ShwXKDFfTaCTYLHapdYH3Tdbco4lmxMLsj7OZBPJ03OEWQJi7VwDCAjDoYfujAkwEKUtL
5i8K3o5BLTkN2cnN4SUwd2xTQYkjJsCJWwSyv2ZxIyMjJgkz77CTUdRyTUHoITpl1t0ulFRxq/2p
cnW1gOPua5pIo2yXH+A2v1Vcp60cdZ6wkSzyERwaqghQa17nWVrIZuu/w8oW97NlKhHMmTmXooTs
LaKLebU2kZy8/45NOiyoM22p7lgdtkzvRi6I78bpis/TWm669hD5zjg4al5OSzJ4OhgUPN4T8A2X
KEVeLSCek+p3zgzaD6zEGhQT018bbVR4RbDpZ2m7BUquleo/aMp0qye6cGTmgeAY605iQXhEjRWJ
41IK78OnHyEfSsyl/mIg6piRJcbHdfBDc4y3dpOxlSQ55XJMdvsl9ji0Obokpb2EoxeBpJ4aWPoM
8gMEAVkXBGlw7xhK1TPCWqQOM277cprnqiPQjg38FT8pLMjLXZDjqlyOehLG6plEG9nqg67OlHLy
FYUfDyKqfNOkxNMi9iaEvZkUxLo1zT9xq4FHj8BbIbfHT32ymr1qmhBDjIJcSOIImvOjdn0hLVW9
fd5qeHSNi2Rqt9SF9W82cbnM0AecVG/bUL+lgHDdQQHFZpbgOYUbeFXz1eyD4N3cwyKECgspikXb
tEN1L9vTv4gvUqGoMiM4XdIKObg9lsPe6RcANedgZpw0AbPxFlRiMMCzvkNi91SnKiYNANoWBj0J
/gk0ZLwoSyHrbEPapPuU3/K2grAWGHQcjbjA4+YM7hcXy864R1AZvTYuyyuz7euwe6x5m+TjpWyr
wRfbh7yKw1+Ja5G98SHGVFGOEXOMyNXyPeTS+8Y/YFONNMTG5MDaKTSJTniDkrMJ3cUZQdOphjwV
7LCpDBHFbUebmrLFVwMJ+4uvAlRh1LR2Y5h8HdLU/Ly69TVmLD+ZQp2HsR/efnDP4eRZ6UrExaxe
Mt+GpXg+G/aRbPPsZPGL+dUdoFhHUu0e9I581XkME/stDfLDzcThzpmeE6lnQdgd81FOtExLHHHb
UThmGtqwYHHjob0v031tNJR8t7ti2I/do41JyIg8quGO5kngVDqkWfhSp0819oTQ/TffDT9fjkaQ
0ahMi2RPmAUQrBTIKk50eTMeNDK9B3qMB3jD7Tv0lZ25c3ZGmOjUwZPDENJ++I9hMjw3/Z4hUR2t
DyOYJPjGfNZ/qDnLwSe+YvVozmgrOHl62tBMgYHCXyNDElPhTl2Ng9Ewz1PauiybsEYU0R7fKOxM
mz4+A2Yh/h4VXP2jsPMZZlaEu3S3tdrWRPZa7XckY6T1zBgID5/vM4IaNca9xNNNpmJNVZB+2tD0
eOfJtQbi39Bmbb9IgCpB2jhxozoHzC16jMW1K4zt9tBAtYqTab9waks/n+E6qFV7QIt7ISYFIb6P
rmLr/AIWTEC08LZcpn3D4OdKcsDy+8ZZFBFVFftIHQcWuzdclTpDJb3xkU0K4pkKwsSVRh6Gkf9q
VbLMTeBLAGzQ0JFo+TyeWrA2MMjmhDKabzW51Nz2CgSUTfMYg48GrA7NTUPpA/Jn+vIcF01PMfYO
yXVInFX1zY0htEWaEE7jfADwr6tU4tkkx0cbkN5l/NJ6Hmk+dMeHIX41oA5Yw3AP64xd+rVwUXI2
Z4B4w21RLsYmORwN4KO2AAf+e780yS5wb1rVXkYkEnLVQPsrUMvtk76HZx+FBPOn/dZBfNt/rYkp
Zbg2R1KEQhYmzqVGu5WnmwCEQ6BgoawEHgwJ/wq9MDmiR4jkpuPFpgaCujkZXaTPHqI5+w4u7WLU
y2dyKnd+n7YPsYXLo/89TTP9dMCbzbmGnMvArFROGps7iPalNxQzpd1mFLk4rQncyPbkCTPhOfqk
2MI+TzbzNtdJm+wxIBuvODWEqrc5Jlw67bY7u92BGDugNLu37WUvUCNNoSODPQIn7L8ZoNIssUli
CzCU7nVWl9wj9NvGXVdeTA48CL+xI6W/Y9I/wcmqxZx7u6tedlM2nVz1a/eDBGWrVYIf84FXgFq7
TCgreNDQ3TPL+f97cJgxHpc0q8eG1DMMUTfRnxGCg2PgIIF4i2al03EbfOu/iaPOhYsqHsKxFcOm
g2WIx18VolVVXZON9GVVcvDBs3lxVeKXNz90ZrGK52vOYUZxJkJVzJEFGFCO+cO4rMf28KZhMVtL
p2kuLBR2dA/elErjztbKoGs7AztQTBDiggthXCDWh8PMhlSH9V2AeZDwLS081qPMXou0PvKYAOKh
675AJQp0wJfwrDRhSlBVp389DrGfsKuaq4kd7xMARLqdGPCj8jEKw4kCVUNQjVyySNh+5IZw/9O8
YKhC/XSg4HeoQWAALQ8PP3XCRrp6SK9O+n6DikCgYF4Dv185HVepdxVTEvWpPYasKYAkGwBdq3qy
pW53FCW4BnIIxRNrGLdkUYpy+sg4Z8uFiERCvPkm0P5dsoacuRyEoiH8YjmGDqVeqi4IPxJ8wm4V
2P2x35N/qCCox4ACwTeKgCCLpPDPEV6OHMsIjQq00FQumWZiv0u1e+dXfK6jx7cnoQqGdziQV+HG
FLC6KRdmTjO6Y0rhUdkZn4EEOA3cJOE+kLewxvoHN2cOGmDKimMtEL7904GbUhsus+2uZuCJOGbq
dIU3xFemfwpD4FyUxl4YBs7E7VrDAb8kWWGaVI6w9jjuZINqqB3g0On8LgBVKUul9awLN96Qz7CZ
pjLmPC4ODV8C29B2frvW+ISOTaPMEY65LLQzwDnnuKjdJ3wAq6/l3721KTnOqg+Gonjn5NdUSRG8
rWUZw0iMRUsSQAENzNZSHjXkd3KruwvcgntFrVu+SUOairJnWP9mgZakhfwSaz7ExW2mio6NY2XM
th+VLgjCnXPX5tzkBFcI8ox9GiLhNDTaGNuictTr7/wMwsDwoRR0g5hPhyFGfF+anY9huxTtC9Js
YR3b5CvUGvUfFYkk6qJ77bjygD+XCh7eEeLt1OOHPzz1w7LgQMWUbCCrvcg0C9NSOBL+L6KiI7nG
ph3zMq0Ywc1SnTZ21/xLemSiJHeL3mBH0TsjJ/18EedaPpraOCsEnpjsoTfSJ2unIyrQrAPtO/tm
NAPG78G9ZEJVaBBo+HEopG6MeZqyazSw9VdJ5hUIoFp3JrCuxUwYh+s3nPNyWYwzc0qCmvgei8PV
0ZeVKdD2patuPrsPgExZMlV7L4MF0mEX2mK3qL7SpUVZkaOaBpceFytzdBAnASTlPBdkQj5DYxRN
XJRrl4p+ZBtohdfGWLWrlrrlzjecTWn+glMYua5mPRVMJwsq5VbMTlCqe+YpsefxJJZn5n82XHyk
JqVCfjhGGy3ZGMUuVO88vzIqLTN2b2/jvMZ28uSSBd1mHTWV6soNQI9iCsNFXHDpzU6yOTt57AfT
jsqSLF/B+ZG54AqhQUM9kpBuTk2CwWBspqxhokS0LsyWc2WhfopnU2WWa95uivrzPMvmTv+2EEm1
vdyd35NgI6z/EFw5HRr1WH3Ayve0EVS8iCYaToWd0//3K/CqXjPK0p3FsuARl9WViLNpQH0IWXQT
X+39Bu22kXxVEM8vwBhj/MnN+BrXJZr1CXytmiE27AidqZqrT1DTRrwEimIQfdij8oiS9k4x+I9v
I55pyItbWDP314ngNWEpQdZa8pijq/m0q0PaciMaZaMynxsNeVfhjoVDF0c/A4uWBIccjicyVG8I
ahrByjYTNcp1pV4npsy6SxLpAs5G/GkXNgeErtA3WFIJazKtYSMr2oHkTqexwDwm6SzYvouXX80A
QvH2ICOyfyOO8xe53L4ch+Fg2DMoNwVt/cEhhDkONW0nvt0hxxb1gj8T7JgnD8g14onKG5fRSAis
NSSbF3ZChdpxroNDJcVyzypuxyjgTrieTGQ+UTCzfKALwi2pAE/YNyOGDGtDEOvBF/qU38T8wbsF
DWqkSv3qeoVpPTzYynOFHq6vE85qp5sBjUMrf4nE3W8JBvOCRZLTtV6ZgpzQUELel7WSxxqTrF20
8Mud66s8gELXciyirdjiu8OpDfP+rDskCjOKuMcF6+kyFFcu1NJQonvlsNJNsEQmil62SgFay7cD
nbb4iUtAMs7JDB8a0bV0iTMByPknY8LvfOlcAa/pXQ2p+6xhmwEgQkKZwVxYUz9gUZfEi3PQ0Ub4
nrp4ZJ4MDkAKZOnaQV8UYENyLzm7kNgfKOnrBSo8Hf6b+lO0W2sp0aQvcAgO2LBXDfLoh60b4FO3
KLSUZBCsbNXnTFk9c1f2RR587W/aIyx4N46HktUmhdaK6ZWcfQIdDMk/mc+7wiEayzSJ9mECjArz
TpXUVy8yMW6R8h68IMdV0l28YzKRUE780jltNdGrE4AmF35ud86nQ2Mje675eJQIUUkV5xbfzHaP
Gbpqu3MBXDu1SrA9kzIpok+JmwO8u3B0McJvH68ycc83Ls6gRIQcoD9anivVUqkFtrpFiLQMO2Jl
c9NwU4CP90IU3IH9EKUMw43PCJmkCUBCy/tW6mA9DAc5NX52hevSaHbkPF90n1oY9q26raiu2ble
SxKss30D61bZ/PvBgLm0xEkqXmZjz0FamzAsWCUH4g6V+eRZ/gVG2GfqrabcXg2kRkJcVJYbo6wP
iGDUyoZKZRXze4xs1NXdU/rA8zJb/oUeNqOfjrcPlqu4TNCZigY+Ksz296UxSD8eRwmdk6ncZHGd
kQvGA6Vfrzy6VZwW6lRncqL6muUCArnormRZRaNVF81RjQRSuaO5BpwAYxRMvHoKr2MVKiPNPygP
GFBPcjCV3eNdWQYXdn1Lswy2ujK3ueMcd6nSUMqVc/iHPe5MqXbLOA8o8bdGZenrSblcgH/JF7rv
Cgs/emtBEn8drdOQ/RNu4VDIkQuuXKlnVCMPkSTU269ZDFZOmNbS2XNaTPpUJ/V5U21v8noiLGK3
lKMSyhHAvnmYw+iZO6RZRWHM9aak7i49m58+w732vC6fgFWt6Tyis2XDtUEIA17Ci6awn/lHn83R
vRCi3eklomCqMf5gpk8gMRI2V7D9EQsuqr9wIcOzp4jy1ZBGNo+z1QRdsBOy5khEzrncp4531X9n
YGcdBG+huLB0bE+oYRiSBrMYGJYiK69p6pRa+ok3r+yhAF2rNMmyAV3UorRPE9l/KtwAzVrPwmsV
eYcbzYMdoP8v4WG/YMDPqYQJe5lR95gWl67uOvb538e/u8Ln+wFBj59q35WgcNieonqTHlIWXY0x
qpAP9TXG98y4cQQpf/bajHtyzRtXIH27b/BOGCXp0u1jnROqo/Cf+4k0bPX93SXJszP6rbtf+1ox
HzdU9bxAJv1fsNhlsLDNCp8nTT1DBpy1lmCnEpGhJ/ksHtTK+MjPtlZADqa11k7ouCbmu6AIJDmc
bpF36HK3wimQI2aZqB22bsredJoa23KQYpdeGQNAr0oMcCS/RgaShNOvYuzfmUUjGHNGCx1unkkO
N/evTG22FcMQH0BArApRC4fHftdKfb16noRQT+xmcnV8YxH/8B9v++9djKfUMPfpEy7Kf3B2xD5A
wnYbe0nljIcUB5SfKhEw7uEoaJvrCY6e8FRDJmvm2STSlHBOKM6lAgLZBkA6LJUS3bLG/3bu2oVP
tcVnP3iywLg7agD7yo2uROFA+xZGd+f9JyMXZK2Ul/X8gyqsunHKPqgMZpDcbo6+C+ALsevz6eTO
dDnAYRtV7TPgVnCBREHC6bat0aBWAEou0E9NCR3q+u2Sv/67GLHx9eNhFt7Z0cB2lFGTH/0OPW9k
UyrryqS7RuSkRopGrMr0O45sSNMNlns3eEOoCDNi8GYrioAEbI+Mx4UEOQQ/OL0tMv/EIPOMP9Mv
rbZzRhctkkgaMQWKD3u5mQbvBXfKhZw9+b/l8x3r88kC6M1XZQ4jwrJp70nXlBowV9hvpxG4wxQS
RduSJJxBg8PYzk3vhI/dyidEuzEUhy8Ctb3+du5dCdDKsE0F68RBnHuiwDOlTxi1FVVR4IPkOB5o
Jb79POzVWt8NJryEtNm9Tt2JQd7FuG3rbkfmmhS5+Bd5wKJq02JexBlUKl778MSxu2L+kDCQHG5a
B9Xi3J1e7n06UhHGSZIytpnhHmOLr13cBI0lCLrmmyPhSt4WTRG43aAcRqFn2twik/TxSIdSO/wx
FsU4u+W0V4ZvEjhEZS+1MqyIUFJKF0ZLcpnxwhvWUAvjO0rzZvJwrBIFMSCmmXUWz/d6k1oq4oIt
OCMw/iQW2zhU07L1kaCihCrRZNpFTi+DLT1nYtUWc0BAugQVBtiRyoKlyNzZmzyzMiwRNaNSCosY
b8ClCGvk0ZYPAnC98htIVzcHu6HRcvsH4cSGLB5QPCie1JwFjStcY55Z11/WS3929LxJ5Pg/MPkj
iiayLUz1NxMmJixhqWLUlzFED27GJDL9w+/R7nxYyEAsr3L1mxle44B/h+a/RMPmguS5sbrT0ilI
4VRLf62hhpEZjMKNVg8HIPlcybDv+k53dYKKrQ5NFVJgJZXFh7ENhz+rZqIFqEv2v2t6kbg3oW1k
r8x796hNt/i2uLbeOLO69UO1ByeEi8oyWyoMFW8Z2egldAv513RttfC/nMADBvi+1AwsAa6hKT4b
Ci+i6EZZJtMKCO4xg6f2P+0zn8FnudNUYo9IshbKRL7WdOW2u2yJ5ReVZ9LBf5G1Ncv2K19peMEo
r5COaqZmh41oRH68xqXcA1G+p0mUYJkQ2r6NBSqLuJQLHCnscoTE/VqfaEfPDzMSHiUUDe3PBsKM
qcpExhJIMGKDtDm6IBSkL2V74jQ1oYPjReRzMHSORZ/pG/M6PHXdz3O4CEfDF96fVFK8zvW51iro
s0IDj8349DJqyYoIPRgZMsCzJJ7h0TdCGnel7IpVwLSpXIkNPvdBfl/TjU4Jk0ExbkqdGhMiWKXt
fl2c2m3ryxSd2P/Xgg7mOo/E9141b3oTvW/si6rplid5kQXsLKtg6Q6wvSfeIjna3OpVEIp/gEHo
QeteqSO3mPzQfHo5KikaB+v9KbWY9Wb/Dq8FYDl2BKt8GdyMvlX2Jg8/ipdYGofFV7G0DTmOTSKD
S1jcr9fYZPYh+1jeTwLDvbjWMKOGjNpagxvMtbyj6Wf/sPCLGmAeIvsQNoTdWT4TJJSs97e+K955
qYT9eJI+SuaRFuCrJwyp5esZwLw26dS/LlCYQ18D2ocFLvct3hbSTErLJnW1Ug4cOmlQEEpA6upm
JdgaBQHIKFLbrWMyA9o2BeEUWt3b6YGPjoe6WBlGQkm4KsibrxImYaLdFny4x5fueCygb6BTkFB3
pXeE7Yk/l/YIzSDr3kjgfzQBlEaXUJYZJqtuHHvOdKZqpR39TsU5Yzc4sPvGkW5Lse7a3ndsbiA6
cwcXWgq930DzvryRTskQZQTffeYb+zmWs/fhD+uZx7zhRHo8NzS5sNLWd4EP26POUMf2511J97I1
yIgkHT39v6JDUSlTDT3yNQDJY/ze1MIJ1LvYbqxUQfUsyEFrfzFm7746YjtjnNVU9ZOa0mz4HAjQ
6OcAQPFF6SlN1numZkISCRxVIUcHYjCBStA8RAGz2PfDD3VyrfD+qG6wBhOaAoUnv20MdZcPrj0+
mZclitse+X8yD3i38/TqqQp7GL5jDLLLlWjtlQT+8XlpCbrHMkInKtZqC1Th5Dt2/gpvG5TLTP8s
RQrwHQ/9zlWAa8a/o0wtJv7jeIbif+q1MzIRlRRpV7j5puQ2bUI1gpTyrZznMymjUpacLqHND/lV
cdV5r7Q0IGmy3rGdMup52H6NMYHYBEpwaBqQTzgOp1/g6EOVJrqAiS/THN7nsBuIWB4FnCDaKnVC
75uON9FRIpDAaAZRwRgRufqlUGqVKA6wP7yuLvMVgvYnIBQn8VFuJePVgEgyITquTVEITRUTGidt
10bwkldcf26LaGwxCz5dqpo2hKpKEiMuCEbnJWdE5N4B0LzYahU62naK7qD/4GAQQy9f9E363Bu7
ibop41pEZf87aSGp0a0he6kRdNhbMNU0qrrWv0bNCwR9JVI1LJ0bU1qzhiUUya3wm8yqmrun8P2o
6v3VQmvje8ksAF2E2mROvVFPhifzGaSSt1cmSULtEw9wDGUbo55vJaokDd8W7ZuiG4dYjqjRsS5h
sQLgBrCVf2xq+v7hEXh4r+o/QjnS+yOXGhBnoqw1W1IGqrSX2P2ywBbCGAg9RbxBknlQ1ndRP+7b
iK57vpjpQ0aAD9/CbUkmbEJ49VnsAV7sREaLR9uWNDUNAwK5ZSQ5I1aXLd0fydiOShsKL5EPg8Wl
1ePBWPDsdHuFYDupfgdQJxOiaBxT6NVFbnHNfpmmANBdAz/XZZEFBy+btQ9DZpfFUS/XMtOf0M8x
PtIdcZNCRZJJhryh44YxMX1bO9OXGV1vK06Bmx1sZTx2ykUE1bILojRhV8MUbvAdky+lgXJd0qT9
bW1hb+LDwMQU0VC8Uj9fRssTjp0Oi6f75lx1Lz36Z4XutaNaF/IcBfsLPWvjFRJ+ndY+kng57QB7
5+uCe7Y1Mw9/QajMA/R9VJ6WUDyYMR9/g4QHvLjglrOa8IIV2hq4IGh5IjOLodzHCj7rLe6gBmyG
CnN0pub9Ab6ZDp3xDUnk3kDw3CcbVU4ax1pra3l6Max/me2zaP9DJK65tbYXqPXud5M5MMovYATs
r6GlmbTS59n3sOm/WW4P5hIYyw9wR/inT6Uw2+z+FSjFD0RtdnlUoT5chHVwJVJHjtfzUHSeB5nH
wmOhnnj6ztX00kdpoPAkuP3mSop+Q8VVEw0t6uykz3pKOT4kRpcTKDpuLvJG9Vkzqlj56SfPMylZ
HLy3rORk1XW6FEmVTL1zWop0SVb2lhKCal7CmSiRXldsONozpaYFuWUsjfWS50Qbv9rDhkBCOV9p
TfhMU7VKfR2V6aDrbVz/43m05AnVP2jZbsUTniojbM++aL6o7ufNIvUWwBJKEoSmIpkebUMjFpAt
knUCHbboKQvNOnWJtTclGV/g4CjTwI9hI77/trkTbVXHefcxuA+2K2+eKfzkNcalIEPdXmRF7hj/
v8Vlg4hRpWjXtfFEW+bsfjFXHFPBaX8tMiEDz8V9KYrAPB+jHnCfx1TKFpIgA8APEGaSR+b8jGxI
RIQq+v9vTIKSsQeR/Mgwf4z5CSeuky9QFEwQunImhzmB5Hw8oryzm/t02sRPdOELK6a3eAJ+j1gL
PIts8X4Dj8O2RdyUCqqwqNgItCLM4ONANOOcG00THF4ut7hHmzd9UHj4p9njEBc3RGM9xSBlcPyJ
BvA8w7n8NUV6k9+M09nJ/7AxqjEidStxFxr7EZH02Y1vd22uIWWK899fHwTjI9jtQVbx6tAojSHy
m8XKIm/NVM/QZbR2SGEGlbMa43ng+/L2s7QGS8Gr/ur0e8buPMH8MwtLpHwIMZ2W+WpTRM1jPcDs
TROhYQ70FnC0V8t+IRaPocR8f/OSawOfF9Bit3uDcu3WZfnFGrv5qvYwntGteBLY7R3zc/sBxhsF
R+QFSw0QuPBvo3Xt0QBGcbWuOv0EmskaNLqHHDPZlAfOoz/ZtAjB9tnTMINr8IKwXqLufNwHgrz6
QJZswHVFlaf1lLjSK8Ot9KSWvEaY7n5LCzhFolaS5KWbrOdtQINF0i9DHlJ32R44DO6i2QbYSrFD
jwQrr0CxywGp60M0Dmg6OZbKWjarN1EGl+KXwQzNSDg0pEHyqU74k6L8mDIDiM24bgFVU78Efqut
W/D92EHj0qGA48ZCm6EpAWb8wIUI9PSkJHWqIdSc0JPxs4UQOOn3J4yGx2RK+03nuJeLwDk+E4Dw
K+Zs7sWNu1qR3NXyrYnekaMCbZYk6bLmRmb8snKRPdRTK53bcbY3WrugHKfeVc+VcfxYZV0ANl+E
DOKrnYHeUmoBb6ATe9HdgUCgdZAIU3XIkzHUeB5nDT+hBdpCpLDxzukPn9m2FgdrVOSh0WPfQOM4
w88FRXulTGO27oquDa1gEcAZeEANq3cKDLEyOcfnZSQ2qLUR4UjoTiD3sWPS4olFxwTXGa9U9cRi
VlIIC+2A916THqUN8FXFueknsNz3YCyHV7ebNaa0HIvTbrCnZOoBgsVsFzoZr8ZIedRPDpiZN5Oe
5uUSZHXQ/l3kydG4R2F8Zmhgk7XbLknC/MJOqBmDIp6vdHiQsXPPtu7gmz/MJ0IYeOIYSS6YMyZt
MagAaeh5k5Or9jMG4H3yvbWvasuz7m8zcrmyUtLwQaMa9cv0dOR1gmuyX7OVR1iHTGUbpopMH2S6
JwMFGQXHwTGbQ+fV+1aAc5ocyqllSIjJtZwyAMJr1jwwTKnLdCaAl7advydAY+IC4+3F3HgGZrZr
jvqoqcD35AI3AR+pmNwRzQQXWAyod+6ePxUkmseOiNOAdo5YICqDhGGubJbHjXjgaW/HB2TvhYyU
Ced61jk8tTr3T/J0LR9o6xRfoq5B80wjVRMu2ig+r+ffJHbE2LxMBoqg9zgnt5H/njNo/Vt+43Z0
0/828/oW/njdoqcPYa4cXOxq5HQG2QkDBs21qLfIjbz3nvD1IC7zzerOWfYTk247sVRI0L8rlE1N
YFJqFwkJdrAW1jUS+I+gyM4/G7UxAc+lJF3nL+KfxGM7KPuelLFk0oyt8rOG73OeUHDfT0lVCIIY
0tKBG5hFBUxEYcSJNI3h0O3u/svastaFqn18tpe1yH6PlR78AGcELs2lVI02KIgixqXG3w5t5nLw
obwkbGuqNGrIWWenbvxVReKQILqY0GHg/fh7r+osZZN0dQbgbZjaLHhzb74QfP7H6MkTAO5E8FtN
7t5nuo9IODLCAjAf2jO9j528+KrrmbCHA8rV5Mqlh+ZnFmLKpBQIEiiTEAqWzOYdXyqbD+qoh43a
KwZ+2UJXjGFWn1PnQKJdTQMRINE+NK3m/cCEUmdbfE22rEEkahybU4bS3BBVYsFlhSkT1/zEHBMN
sI8WEJ2amNdVgqYULXRigD4GY3KDzGihV+4aF6at4ht+JCPiHPOSdr+J/29v95gAvJ7+OMYmhixw
giKhnrVsx9itqPa23EwnJ0OhIHTOyp/ASEwRgjUjpu5lF8GcGYgqR+DdlSVwY5GD3gyxJlWW8aQc
EkMV3WTi2YNABwVAQeuKllkrbB8GeGwIQ9MOSMbWMTe2MvuGHYlu8TGkS8nD5f1CdQ3+jb1AW7BC
UlQH4IShMI2AycnNMOjqZ/+mp1oZc+ZNr+YEqxfGcyvxDKJpA2Wl5UqownXqzBJLrbWZzPkhydm6
AE6MOwSKmRCto16UBzJ6vXXDXa26woux+Y1geoN3qFXHLGCYaopXsEH6izNN8+ZvndI0bZHi4TE4
HM5sC/nIhhqhlaN9/Ozs/5+F+QK+k5HB07OFsyZ7LWGfKXE6GzQTKXvWefTjNKZ/Rg/WSockaekt
qRVhLtlpJoRXftNCXsTu51zxrMVWnMzEK/UQ85YHT3fEvWoakw7eV6FG9+t4zmcLQt/VJl3of7uP
sH0mruBfhLD7IRmECVGos0CcQh67X2mWO4FqqJDUpOJzOFkhqM+MB66ymY9WxlAYyjrHQs6VQi74
J/t1zzhC5QuCBr40GQBaRIpvUZ5xMOXyJWNyaa2P4MGBfRjtBGFYu6YEQ1TC+TWtl2DwnVIdEhJD
FzgQYhqK8h7q4MhZftIug1BYjY6/6pYFmaBDFEptCxRBOBx74WZ1JSBfCSpAb31B+SOB6oT1+W+u
rcLC/OR1gocWHsntgZ1BYwDoNe6obWQ6/w7ugbJc73O/+2LkU/s1xtX51VVs3LJpdW5J10RAB7Mo
PEAixmK8G9Y83BUl+b6NG96BjnSLrWaq/4vmacaZjbqec4mYetOL+OmRTXCv/Zy89L1Z2dwg9r/a
hBHJUoTCSU2O3cCV4Np74FBkqmBbz8pPR4KjITUH+RQTFrihpqF6amK9o+pV/B1zbJKiGqaO/d1m
DaG4TSwTNNngVPHqL87xUJ2I9T6hI16qrUE9Wi85vUeoSySu4aEVXksnTUkai8ehxFBAyeRbRnug
nBjLS9dphheWfnm18K9/NvZHbZNzGe3G/6fOb3v4VApp9xGLYNdi1WDwhPynzN3NiHqihZOGCHIW
QevndhnMPuLPcp1hxUgj1dzizoLGf581/b9rLtmzKZbyLw9/wZB63+XemYomjrzN/dxYhDoGikqh
WQA1AMjG7SUkUoMJsup1IhILSwV4ox6pi2aTpNzkxgSrBF2uR7Jrcj/vUBvVhb3tWGeAf83IZkPh
XYelSspnDSepeDsNSMTMPJKyI/hybvirSrRls1jvoE8DSwRbi+ckCl31Q1NFqKLP65tCtYsZ293y
Wjjr3roUg/Qi03NHUfdXdI4WV+MF+uIAcikil4HmuZjG1EEfCl4loREIXBdBxBFhBCuEep6vAhPL
cG5RkSeIrDK76B05ho8PQlNsDTBpg8Z2tGSU9YWw02dPe0f29jcSkOlTU6TKsI7H4K5ZXUTMKTdj
6EtoJLgcyHTjTao0E/5eO6Xldy+51Jpq2vRe8qwod0JO1yZYwVLzQDZIiygkvOC50ad2h87F/fj3
yVci0bU+bEhBsJUXUoGzAQGg8IHM/v0yejDQY62e0owoyLP77UwsQY96CP3ZhWCWLnnyrvfLICG8
k7AWwHfmiWILet0mDJ6KxfTY0aN6Aqu1ZObd+C7igwEvy+kCkrUv8Q2WlPS1LIEcQ2Ghd+0Kglul
KjOLRzsslpWY2ZDXpL1gOPNrn6s9FkDxWe5gNjOxx+HEVCUAsjgvqhZoly7xbmPsINKyhbLX47TK
ehuDtkIvfTGvD1CdYncUC84Gcw3fC9chn81Ph61WGmV9KdyLmQPBq7p6en1+g3SoYa+nixbTRXv1
g1vfsQiPSz1Q6/QLKqthCbD5G/78wNvKheTzHkFKC44p+cyGIhMxkb1hrm03Yfue8nnC3TN6+zS3
sjePKYToC3NlQOxdbQ5m3ClyCYVb1aZmtb2GtZrSeklPLH1qkZz18Tnn1GfiP0gTgmsScj8V5Qgf
wr50Hhsks3Qe2a17S3A8htHnKB1lePI0t9AFrdkd856GjAdCWHKsmH85hxILy0JRrCnXuaaAhV01
lgKfxbmYSKwanz00C5pU/nIkxq05uu6KJh+M2EeVUK1VwyKmHU4ae+QbK5siBV1UN15NirpJsl8F
RnJpKpcdNY62aAoNd2DLWalttSTw2/rEqE6xjGiunwhatCJYasWjOiaUBlUeE2pZZVSPOx5Ze9yG
uwGGz1ZiOYTQEDDQ7WnZ8P7djO05m3+764YQThPHxJIXL6+6SqD1jQbsIV+qlelf2eZ3nY0yc+35
r74gOZav7HmqC4eYRpnJ8/HzeOCoBwzrE4UrcAbtf5n1ouxorkwr7gEluHntxsNDBhb083sPjEI2
M7LIZidaGbF9mxsGKhI0NhnL90kX011MBTW9hRXulc7CxpNEY41BabOAz6aXZ/EQyBOqwZwtaekf
z9EzHrnrwyF6m+GTa3PLHvo8IH+d0Nwo1WUMw4uZrunZ0+cAbsnhrrXz+9HPYZBbXYkUOk4dZ2rW
qfV+t3llH0HTYNgL1eS23+quC8rX9I1zp4fOI0+gNfjv7aQ0y9xy4ZSz/30T+H1BuuBToi+5kSp1
MnwfhDAynQQJ4OKH7qgTrin+qQTbjBYu9OcP3vH9AB6C31yiLo8IjKiGv54aemK5YDW/J6MpWgd/
wq6q/Ys+BZzcukim3fmU013xURLtpymH0u730Hk6o7oKCuHfSPVltPJW+MNx/+t9Mmjr7Xpmhg4g
lOxG8F597YNuHJm7bjlLR10iuVYGUTKugVlBZ3MYFI0Gsuk9KUb65ebFrOH8iA+efcWbrHlIxgl7
suKe7BYutW2b0jIr3sLch1XCA3egLUMcHO+/IUv6X/r/qKW6KtNT02OvNnMntMlKEi7/DE4DCc/8
8Dp2vt4RrHr8Iot4RnFiVGSDKjIA78d8d6gSAnHrGgoQNMlvS2i9W78cg8QrKvlybcKpa+yjBUch
41WZ5MORcjrSV3x4EhiWAkIoTyio9rFjOqmE/aVvsODTz+e1Xi0PnofruuCx7ZaQo0P5lbv+4nI/
1BcM1RJ/I3vPhPoeHODYncLmIvrCmzhCzLt94IIIUdVPpVhgQiWQqN6p6D9UPc3KvMM4WhmdDrBu
v6qLGVdrNBRUwS31n7cUuOtmCNjV6f8tTijL9SB4sjZ10untYkIlTm7HKPSSw8ixwR5EGiOSuG5n
Am1+RF9cluJ0CYy5/+HuncfDQm2ZZi3ls2drQRURI7BKLRKiHFGSMLEro3HkVOLRQ9JE+qhgjWmQ
4HYGdLWJ+KSkFvyeWEeHbTZOMWyx0DvLuQHlJct6o+IOct/qPGXwuCrc3pWG9yXM8FxJJBI5LFrV
He0EpefaWDzegKDTbTkrWoy7suc/mT5lzX2nkLDTWK036orCtq4xUqLdVXtSy2/ZLMn9MgCaOve5
5KXEDKaJYB+ubxICnhBYsyk2+VE4ZaXk76yekz4XhiFJNqUZk6zvSjs/S3mxSoiGJAWJzIQTlN1f
uP27FoD2kUJV3pb3371bxd3aJ6QMhwEynL9xGc2SSJXZiK1d6DYtNlB3qxmUDcGsXzUHOjLhlcrj
Auo3p6m6JLfqH7iQWZDZEhx2QvbTPqpAxJs40eC8mHIe6Kc9uDxl+wQv9cKNBNoOqckti5qofWdD
bQTX0FW9C3jiW6Pwqj8uR+3HAVz7P7c5T8NOlZFFRxa8HyNXS73UCTWqECTnTV3nThoaP47HIMo4
Ino1RHTfXkus584LFYLi0oMjCmzm/t82SgPd1wu1y7LCL+RkPXxQd4XZ71mLBIKHLorJPNW0Tpuc
EkzhmNFF5eriMvtJPt0NizuByN8yV1r5WYJMhX/UurTIb00cZFo3Z4MvF2KIn7XG7vtrUgupgC9H
aQy024vwPWjd0dhXne69Yv+uumMpTsaE3nYiIU7n96I+8QmiGGkIndSPLn1GfhReGZmEtPGihFg2
Jaya3CKvnS3oa+V0eKTmQGCe6mfQdEcAuY1/xRY43GqFuEAaWAZjg7rVglrSJnPKzvVs8Od+VhJO
1HeVs33Vxf+f6OzBlFoMENH3NKfeG0CV0memL9if+ZN4w/OqY8IW7Tg8OVAWa/MKHU7EBt33Hyf4
w3ap/5eQNNURbBJiSv4uPVsK6bZ43p6TN+tTy+u2sP2W/gs8GD6osWSQvOoIONnwusx9QJOsBWqw
ldmBJYTr/RsYsLuQMOh2DZSjpsazs0zW1nYqYJ7aDXp4R3F9pymrqP8dF/CtHP9ie4y01Ekie6qZ
8G4lK/WwjRF+8DC/Zi1i70S8bo3fLK2u16sU5K60vzaxA4rFVKBIJOQtzbZrsPBwgO41hwUCZ5RF
VfwRaYdLERLvDjZESZgmI8dJ2/cphYUrJ17OaQIKkfzNyvmvItKKaQoTXuez6rInr10azosrTZdQ
GNHtcM8/9gS9jBkeDV2vONuQCiWh1oHSRWtreMyNJd/WEAnjNRZTlSyIk2btm9A7nQyQ9rrgMsUi
R8Bd3Lj28/qN9/4M6+ygfa8E4VJTHmk243BwJbeX4RvjRbrzvSMj64wASnaBoJJXrskYgAkW5rA3
ntMei8nUrp0i1bX5rVGq5emJ27Lf9MoLGbPPfbHEpK9GxfyCrELn4Me5ZnD+gTRkhVlPX2wsJGQ2
45nYEtHSeikY3jb3H13XfYQT88EZYhwTc8J2o6aN2rgkBaOrUPk6vjTGMJq14iOhenyjKzdSOwoY
mIZurlF/rpAz6WGSIEEyjpBCpTrvH5WziyX68YtalGj6ajVey2qPGPlYBl0JQMTdb64mEkDdJbqb
T+MQKDpFQs7Ocn8VYAtfWhiMd6C1HQ81fJyhrTD+FHm0ZiwbsKHMIlJB8MJ528u/JaiOob2q7tPG
VnwZ48VJP75gdF4CWkIKEEdLyzJdrOzRlAdxh5ntsmBdi8bd1Equm0obzZtRy2DZEndj1ATsijhP
dRsYvcF12AOZk4z3sod2fNqFuVmbPGIgOctNf2WKUoewB622tAfkJTpqmK9dbdqeIyFwfA4uxmeW
OYi8e4bm/LGHl9Yyfx5ZqiSU4nHLdVGJBvu/rVdQoMGzd7uTw7ez2jn+G/B32dYDhY66apAF3XwY
nnu473RHz+S+nGqLIc4RDXiDeI75czDrlzPjXtzVG6t/ayDYBVJkZUUri5zy5cIDHbFgqq1pcGjl
ayGltV8iePc4lUazq+QrAcuPSA5C6XarWmHe7P88hEc6HQkg9Zhf7w+/HwZwfXCWDa4tnPHGjZzF
K+ZT4nkDwmDSV9cXOjyCDvVQSDB0/5/bTHP1KhBlHTClEjIPF6aczsgeREWgfvitBLSs6E11tAUX
pBXUwmXI2o+1mPor5RAhQpJRDFAKC/yuOuMFuh0/dyQHIsvZSHNYN9NeK3R29lcFi/y7AYbJ5Xx1
rTr6ZJVIsogJThKeltccG56Icabnr5wUTMHVmNbSNBMizoH32LNT2p36wuSuH+yERIdH0P2qhb4R
WBI+b4HMXBqYF/q+fVsd8XItmJQLGuGwUJKnip7cpciY6M4707q8GVaBLueZMvpKX8RIUy6ivwpo
QPlXBE4yt5sctKJZJU+yFiigo/NUMnbpoqAKN3D6GXiGZy1AYUgB3VFbmVF2x7PrZw3jGIow4hTc
GLfELdEWCnLBA3zdBrP7CUec6uORRoqLIl8LMwyaRJZV3gzRSvSBPiruPZ3yb7x9sbn6Ji2o1Lec
MpZuCVSwWfgkJa+M3EVsn5T0W7VARNiBIxq4uz70gUe/i1SRm5ZtNJbjtiWNDmiT73INungsKKcM
GB/alUCaY0be3852peBZ6GJPAgG8aihrYiE3ukplr/kArY1H8aGsRTOwYb5veqpZRnm/4BzwRzdE
vXuwL7yUvNYg6qa9Glq7lHjvyYrECLSs3jo2cx7B6Cin+f+80+ZJEej4fTv1nOCaMkxBdA33xXZH
4YuizdR1anXHA2/YSWQdp/2sD1RQTY3zT4geojWkXSLZb6KHU12l8Q/uKTkxiMd0nPPZmrBfbpTX
x0rlLgZbRbH/vCn9vFUsfFCYek3cknzclhgR5il0869hu7kpSDzjjddSf4YjHLWvGZ2oH1/77Z83
1XzJ89xwWQwaTix52Pdl3gImG3JV95keKbJXwVry2EmTqxe7s8SH9r/shIsBfnqh6Nz/i0DEbHH8
G1pcmyTAOvZDDicZy7eI4thnChtkhrEMYvxjXTCBE03vuM9tG8l4QRWLsQMBnSq2eEN8KqWMBoW5
Au3HnLiTjWlEPgAOwqCnteaxW4Tlp7VIbpmbEn/hI2rlNmJ/NigI+/091IbrwBXs3EUdCElHxs66
4Mg872duTBh8FRHcCIyMzk2jUFfENe7kjyeo6tXO4z3dzozJTAGLy7UdbFIvK9CPWe58AqKZoTFK
n5t96dLYjJBCHbxd7m0FgO3hd4NR/kRT5iP+11u5cO0MyNTkTU/hFjQsR9wbz4zm/fI1gSTX+xK2
xxtpVUWdfB7jx/8IX3gqLy2VLGFw+ds530Yjo/hPnzSVaZ0NvyDUDWGrT+Exxnc1u8oRkRtQCDx1
DPil/qBgImmEXtDucmC1RtBYQnb4q97zqMi/jxnmQ0zPZPfnStQfjz1VNVv8eShzfYsudNUcvwRF
Eun+BLQmhpz+1upfm0nS2iWl9FyLo6UzSuSZxakc+JMw3LHntzWeC5P+krPH/njD3JfD8pSPndE+
jFQV42F54TPSB/HTuPkEpda8rVbygMeuXWs+lN7fwI3Cgx5KEJzO6UZ98GzeRnI1eUrg0j9bb7Sz
z+MOmTlwaTWzn6gXPY4lYgPxeMdQUAFhSXVSGhKyWaSSxIO7UG1Jc4ejRmPbMVVTMnK5vpC01O+q
rJWKCty3TuA2jhnuFOQq1CMQdRedVY+dsXVhG4rPfSv9KbWSrG6cinuF4Z43iEzgjZOfq4iOiSn0
jVBEQ609HW7aS2WsngB3FlZ4+B6OiqAABHms4Fwipcr0Ke+Bq9aLJra3XH/w3xqVqV4GegKFwGwG
84nXsg4tcYlF8rFM6ap2I7QGtotHrj7iwRa4wVfiT5cOORDU68be7RdXXw6MntmnXMR8oE8HoLYT
96GAAdN85u4n0jbj5dIIaQTU/b3ZZOcUVJHce0RiWNM8n0xHwp1OMtJisxiBGPHZcWPU1t/tNjGV
TvEwiDSEx/5kM4IB/yFUmfsxj8wLxfH8PTR/lOFBK+nsREnohSu6RDzezkuxABkxYKVjBq8Mln7L
C0yX8Lg3oe9SmfaL1cmvS15soDtYStP+84z4Irg2dSxkfxei/qe+d9B6YM6sIj//FAiG3gAz3Sxp
hUJZ/GL/Dbf7xgSed0dX4zrJ+xUJ0J9rTIuLsU1OGGb2+JWm9M5DcKwvznch+ARBoQU9KUwjjkdM
OKAMsMFbY5AiSIH/NTNqrQKu8iQ1UeCDsG3Rvsi7n7LeDM/4qKAxo858aFKUn5HKvxRkw1Msxth/
9OorUsqU0wVAx7r4LYJM2BCL5k84PFjpjuLAdgabOzUzcMRSFCFgHOHO832p3mxlzvecaRGwJl01
HxYMpa9zXcLihjP6i0CR8/rC+fXSfqFuEs+2NKPGdRqmABSHvByJEOVFgtptsag6a9PfLfXDXyu/
ebX1np5bNXs5KGIjkbB8kaTRKLnQ717BDQNXZRF20cbDiX9pFntjPRNxcRIyGXc2vnz8TJJVU8ru
t7vOoqIE5QOF/aQPWYcrzZiZ5YxudIsRJRnAfGbYfaEnr/riezXLiUmH0wUtIgPuEZEj9azNPPwJ
J3x8+N86D/d01QtXbnQ4ljo6Mcbog5Ycf9B6N13H/b69Au/GLM/VTt/+ZcEtnxubTLadRPPThsVP
OeZCF7LXU6em0iz3XPH5xMX4yuuJqHA8gfDVI2mqJQUpG/afEsKBOQ+3jYQRaa6OZEwhDZk1kbNZ
ErPBlQIC/AoHocTgQ8TIeoNzmNYZH7Rs11EpWqRwqj0LLoFIsMqtEFxX8t5m4Hrb1MUaTPlBzqa+
/18ZbldF59u4Gx/9/yOL8rv7bFbjNSltC68B5Qy5Pwn/KaCKHFK24/RVvIDs5nqW4RVvqJVe80P8
xg8BOuoWE3FqT6d20TQURNogqJB9Zt8X1mnfCzcy4Ca5HE4nnbP+0HbZleyDm+K1TknpaPiL5fHK
dT0z7QhIWOFTwqtZLpXM5zK6y4YuSgJUYw8CnizLBtLDM/efRnlOwZhCWVGGFYS7DjUrwGfFn1Hn
mjyfJlawuWW6Q0CooRPjTD7lQzlXGHTfM/Xh/3Op5oOcEabzqfFTyDyiisRIG5dnENOkH8QROPT/
N5JTaT3xTKoZUpvuek0qcJYtFdiZS1AVwGKY8Aq6i5F0JpqavkPSmBEPNqiDY9CrTHwsQEAbVhms
i29hCqTmqmILibs9DkdnLeKRhb59x7UlevEv93W5q8V7t+hLMLB9hNZOe+03p+wojUsezp4C6Hjp
S2PWNVoAxsPWJHf/QbP5eW9ljaSzzIjpp0XzBWQy0UI7sXcS6063aRmJ2N+8amcc78i0vizwtnwf
PCLkyu+e5Cp+NYjmzj4ViOqTVWPd44Ga5G3CKCF1gPtWfijXThIFFmgF7U0oDhjsSrXojnFmXVGL
6YJ6od1s6lsyUsf1rHxauODtSr6q7Vq+1MDx2Bj3CXi7oDevDBJMb2UcQ6VRjQESj8YaKVruN3n8
W7XY9X8h4zvgZBX0/5Ki67z7lAblJ3OPcoBNUfROHwor6YSdxkbTx3ROml6yNAXeyJgJZf7mZP/+
x1q/TGddU5Qi78YD3boayfrU9hxbLrVlHBAnV8giKZBzFt8SfTO/H4Jlxfna1SdrMJXU03oqHywr
6dUfTG5IrQvB76kNn5PmufpLnGBPY0o6G1cjueTmQhCQImggR5dBjSXMY036XRI0da+YX/kGqrVV
BMneUTkdZ7HFgGJw8Pyd6vbcBLQpByr1wWpPZta8YjiN2RlyAJ/fnofArlUXZlgEKU3WM/FR/5gY
zBIYd0LmL621+/3Va48oh1+mIWO8JXgbOF14nwUDcztGeAOw90dMnz+bKo7OsfmOYSRc11mnECPX
gc8jtcoG14smjkFXoaUUNLo4zdXYif+1HUGLNh2Ka4rGg+bxTJ6KZ3iR6EfjTizj3yQsgJHdzXIl
lNSib7ucpK8B7mlzH2oCCfWyrLFUg3VmW6i672EJPJXV4IlcMfQ45UusntPfULyOGrZQUiSSH5V9
BrYOqjdxIsSEkotRSKv6HnG6IAqS7KqwC5wmFplLukPt/rsleEJb/VX0C1TivI8n0GcsqR5c3opT
YEXNgJaVt+huTfNln52rNCuuexZvCfR1ECOCOaL2SNk8OTCz25pDqw5y0PlThGW3DN1RvKzo72Jy
YrEp7xaolzXJDhPdIR6MIGjyqTRfOpOq7rryZRRVVH+DWvSKj71AI9GSsgeDCHjgffn2qGKWBcTj
s67fnmpRnX8eoU4qeyTzmipX+BvXQz1uZEMrbSa5qVuPfuIp328FZzoykGlkgGgQwyKuOn8cesAV
eHm29CARWL31fdc/kp34h2mkfmWZyT0Jnl+JEhU+jxX6ib02njYm709DjYbOV3s7ssg89H8Y+CjE
QYG9fIPxJdt+Ht2MKtUgWDoTImbDPu4Y+7/+4LKmy6MV5Jc+flNKTMqMp7fiFmL7eYY58vUuJ7sJ
bGKw2pra6ioSpTAJbtjW5GwhMAZ86ypTasUqrsUrOF8pk4D8Z7ZIr0d/8Y7tZ58+CbdE92Rgj+D/
C3Kb1GHRBxf6meKO8gg6PTTkhxKQ5c/UKy8ObEtIgGrvfhqHe8ffANWA74SW8Esxs+8kJY6IT80M
WZ4qfWHdWXX79UooK/NcyczBR52i0TT//1+UySWUW8C4l/puREk3XxQbnCafGz0OCEorhqWsejZK
/KKLG8GYIVDBugnUyh+cYSbzmjegmiZSdjPiEpZcXGIsvwcVqWw48mzeXM8wUJ3KYFHeJ6H4Xsgt
+J+ex3jCE61PR+ih0iY26LAEd2SoEaHa6bkoZqI6dEjXSQFXukEpNfSbtFADUo5e3ScV6A1hHlpo
rB/yC0/qqxvTMoCML+mfYQiZW2YadKBqEJW4ZUHNam/G+MiRfCzjT10BjHgoW8mXk9CcZAzRtPsD
LGXz/mjd3oVdJryrb+KXTK3gzfiT7tyxDJGqWyEY/Iydj/+tWtbtk4V1ftrQMiB/OrsOdrXZ8ByL
vCN/2JGHwDjfOJoDnEcAJhXq4noTihNDGQzv5EVfYUuAuQpFzHrqeFZQZB6lvBfAHkMXoH4F9FTV
4VR4jbMrV3Acdk81562t7+yjDzvnQlUzhLSyzraQdNnquOW3658Mwoldt/tIWlGfa6MQzBaEANtK
vZRINL1tK2qn8A5umyCUiNrPtWyqmvMQIc7jHPnuERmXbRN8AN2MdFQXDczWaBdgeDE+HH6rhhyu
+4Y2PX2ZD2R86qIO6KFxdV72OlDTS/9G/LxYOQt7T1T/oF4bXTjsbGKQI74usshcYtyk1xJZGoAk
XcEyySQmfbu7LnHbR0uQjDJjtVBMVNez02OJtRNrVbV40+bfI6nMd0QwfwePpqFzx52qMwZJkenW
XOLTLbDFimKInHFFeekgjnX1Co4aXFaxtWfw67693oBrMPNs/F/joM+0clxVyE93MjqDu4kewX9u
17LpM7dzaATEuPVkojMPL0uMuAro84QTmtcY3x880veRbPsF2elYKVzfTfv0iJBpg67jozl7va7f
pWdmhmWKxf+Xs/Z1cIHx4sM4C4c05GgZ5RjtAXt80NtIIFKb2TA1sP6p/WrHSw8SOiPE4DNmUOf0
VXFtbPkBv+yFZf1MQjXS2kUbeoLjcw+vp4Ce3TF12hDsjV5ZixVsH7Rppjdp5ZMT3ny7tjfvA4Yh
a7LPmLxO8WQWJL5zHLWbpO3TvFyzwjfUTkp4WARxWoC822x/WktZ+zGlVgbKL2kJnZqe7HWj8PwQ
KYPF3yxmzody2QVjRvtTGxIsYamzN6SiVpIhDFQrRxEWVUk9wTQB7iqUuxABPjxH1hWRuxyjxcga
EkMYA0mxCmeq48uElawhSJ6ukaTyIEKMJmcMgqUPZm3lYpvqXkRpSKZPLHFieYzGPBxvPOcVTgJc
d7KNmKQ6/Epqnlzt0U5povSz2tUbi07FWNDXdr8R/iA1M7h1UDNOV/K4hlCkSTvb8P1Ww4v7KTnR
f/jziDHvKxlPEfPJzUfCre/3hAddr6x/Ac76C5bGgYlB1Jstrb4hk1A5AoGlk26H353roqBR4Eyw
sUuOk2ENCMokDZLvn5J0HG8jV/QtusqVOUu91Zp6HFzf1u093E3f//DU06/0CtDgMcTreYpAdaAS
YxSQnNpANGyK53uiK/60Qb/JN7ILM2gxPXUl0nat11vPyaNwEvLEvAQspYxqdPMRR+t+2RMApuD0
1Y1ketPl9ja2b4WQ1aq8AWTmf8RBL525rFOs8+g4aiLK+kjpE+e9eAoezy97WqhUuej70alKepEw
yuJWJzIWBclLDcUI5+7SACF1A8JzydDaWPZpiGrTICJW9ruMvar1xo2NDzkD3YeJK66h2qZCyhrQ
CSI4ZoVrT/PPjahaWPShzycDHry386yvtXWSK7yvIuaA5lo0z6YQ6aULwwDWycDk/PtOVRLB772p
ARDRMyxhounA4h3FsYD+3jWsNwhdIaqAVG3ar/p6i7nyNqXUhGmkuPrlQz7/7Rxyoho2iwWM+5wg
OnMjF4EG+OW1ZRdlkv/1Urh7mjJxr1bLwZD7NoobQLnsKvw3vLxiy6XnQVpcly+4I6NqQjpi0vQ5
GkKlFUVbC1G6YoBBT4rHYxfSlKKf48J5Vdfqdy5ywyg/pozr0cE2JHjrayXao0AKsX6fWHucQoJ0
41rTtxZesVL7ET9pW4vJ/x3T0ijw0wYPIHsBWW/bDLBuPf8Ol80cpG3zsJAqCzR3Qbng539XmILe
MFkOPPgDvmZizr9/OGs2Ek1a7tVXgkMGm1d0z5UvQ+BqHgTBOJgnYIJxLZ/KPWBCaWTswufQt7d1
/5pvViab/ZgW/S8yM44l6PDwX3o2fIlo3IVo526zlgDRXhX/tXFHUaiYP54usl21P43zuO3X2K0p
hPCvEsV615DvI/uO6GpcHMynUTdsyXmCEbCTO9JCeQMaABpOMdN4YlyUNqxpxiCkoTPAcP/Dcpza
0eZB8mw7jyxdBOj8BP2i+u7+aRfLk1h4mPGuksmcutNN0AFdMdfpSREQOQol328KQobPyN0NrkvS
o/BvaYfjMQoXoqtb9DXoMw/HfgZRcvEO0YjLM6no7HXzSwMS/AUbQdDSO05DspZC38zG0DWbDo5y
faeRhroCx6zX4avGn/39POUtW/bTM5btSS7HIKGH+l9374Hr3HBkHkbqRGZCvE+C7bk8wmsR4hRP
ZOc4supowWGDnmBzp9iqpSHxXtFejmumJR68hmxGrDbxTThZilM84JB+L8gZFNWw4MB/GEjWHG40
w85UIMeoxl9pe9EVg+L5gnnYxaj9SkXc3vyfQvztgY3LCZiv1u6c/fyK642eNfl6rr7rzGJ06ofU
/P0hzni++OYhMOAV6le8ukaP2By0y7dmNMqkYZBBDV6ThemvSygRhn8BPwmRjUxG+f9B+fhjoqBf
2thYy83nxefqxs8Q3QApnK0s3ZKHh6RdmZL38Y/7a/8O4+PjzdZUJSrHa9UahPs2z04kSdIYLl7N
beVYwQypxALnVnqD6sepKotkAoWKwWvpUcAvuDjTo0bJAKY7I8TzBRdM2b9SLV+pIkoZENMAgPuN
f+FuD9yhLR5qVZ4FWuSBdN4GDaSkvVicMsFuRHtFrx8/9Tbpbcy/Xwkrqv3UT3G+2hDbWqNE4+3J
mNrUQf+VBuzCK/VWwNbLLSUsI0DUqUycdeJ5vC6hwA1Rpz2QHaE2sqnJOSHic8Bfk2c2YASEhTqZ
pRPyrrYGeJM2UZoJj49v1apojLa22aCCuXOck3rE+Rsh52SmbOZDk6UwwsQwsWC1ROlIXykUJAyq
sg6B/OdzaOyk8XwwcaOGLvn105JfGhvjB7z8Ff2lTEUctdRJZeRu4PekhfMCky8qCwhdDAHjB1By
YB0nntCea3gd2ifJA4pJy2iLc+ZfRu1UV6L4tKSU+ojsHObI0qxrrDcP1hlYTzn+hMLbzwtGUc4E
frAgF5gdLxbnYmPtMylEiCBgpXaxV3BkDdtyXDx1kDF4iBPJMqvRLI7GhtMYe1SrtqFotaBkRB7A
KX/op6jJzIMREiActAcaM4YAG5TuavWT7SsIaUnUc26jIXRXUbBPexK63eWA3eHKWiSUQmdB99ji
Yicwp79DPLuUeE3X3ilkww6Ujx1f1KbzCxwn8+F72POBs9qXuJ2uR0uT4/aqw74fvycll338WB5a
Gsg767VCWpP0WmoxgFyKi/V8lOlKd8JC6a/ppHotfvaM6SFMirbvTkPKR8rjU8FxVejeu94UXGnw
+c6Qqe3sJZZfTjecYKN2LWwjKDNhM8OXeCycQ5FnKTLsW8AuMrVmeUu9Q6N348Xlslw3My5ELy7+
XNCPD0GZ5/aZeepEtjaFzkyg7Cax7uahxPyigFEUa45ENi7k0tsgicbmctSQxnOO+YVZ0mmBZRU6
cW27d5KoVvlbHSzjd1/IrJl9ba+TgsLsiYkfNXlkL7kz77XBIidEwwqa6vmBrVVubYgcKhYS1/aa
Fc9aXmTlf1arycgwrvta1bsKkuOKR82R6tZbRka5m/s8kb/qN217Skgh7ys7nsN/+OttoKm1OiQg
jC009qHBoFeUPAU8WUBD+eJH1zYnc3mvUfO5UAA8B6T0cjdZqElqq9eueTzyU2OAKxOHqfYyUzqH
LzmqrKye8fwIzwA1quyJeBYpK60ITNeD3dmPy7tXttyb4YVKfajMm7NjFzRleBg3bhpEtelRRH7a
+Kev1E+z9G3bHr4z95tD6zeCstMmXwQz4Bi7AiGF2SKH2/Clg2POa8iJoiHINfVpz4ban2yn8RPe
sAMYBL6dAn7ADUSjESFWHseCFj/yJZbam/9zvKhudwLiiFqb2m8rLqVlhjnpKzbQdf5hSQ7G+s5e
3m8GiVO+GjGtn5Ph7HvtxTwdFLH/OyZpViBtAd+ez1NrKUdu0pqLr2Cu4ceyzqmjE0Td7uddG+MA
G9a9c7Lh+jJyiR4mmbhN1xv3zusJ9871+NImvdebUq2dTzz6ZrkPWC6buuOMrFjg3J82j1wN9a2l
iMhWAEmg/UlB7TvE2AWRlxpJO/U9mBui34Og1lVX0Arvk0jhB2iLEaIyUOhv8oJFuuz2p6Oh5PtB
qXmPtF3KHZbAGSZ9EDzLm4q8KhuqSa9Tz5xiLi7AiZqeQACX4xCBWPeGR5Q4gs0wjv3Bze83IAyv
tjSJlrD+w1zzi0f+S7vUe0qzuJl0r/0kaGhDKdEY0+po3NHDI0jjvWnuEjm1G2UKOMvZjwqg2iMh
vgfP4XT+s0MdVBZ07/yiKrnDZqzynDj64AZYOlLXoiKin7n2xmH/sTlmo5CxRghtGtzV+5Ra4n5T
c6Tea8xJrKoahP8pc4T9JjUzv7KIs124Ql0gRvGxSZg8as3jis0p4B/LBPCmfeBe5S/qNzW9Uj+e
UmAnodrVhTJo/Q2OgelueFGc5NhT2lVe3cM5f/SWU2FX6hxInhLOI7O0nOyvUe+P4EjlcgkYG+5H
x1sSlvvjQYdqywaMk0CKUTe4ta27dZKQNIJk1TftAO0nMGRUEsaOE/3TlLx7FVxvpa4OgcGkOnmt
bYw8C1vXfbjdQgP5dnl6cmgM+L3krrr+xZm8vYxVLW+nk5G1MgRY3P9Q8TkR2gHQYTiyLHzuIBJh
5ieDjF0K7Z7s0DF4FRodbwYrZ9pbNaIjWjhujbznF5QnBFgM7TrOybNm0Kkcz3s8z+cEZPnq/CBH
kCRAagYwqliGnJEfk9PWw6tiOctEThI7WQ17u4tk1DS47hbF5Htm8/rYTSo4CFFXR4lehR6RsYxR
rA/Zju4nqEBHjy3HGw9ixYYdYQEPzelKs90c5TIVezbuJLcWl1PwQLkEAwDWr/MVh2ABa8wnSFuF
r5nPwSa5u9EUztx3lEOALcWzXDqpW5eMN3s6IQnGISZnG3oISKY3Z/bIGQ8h4LhjRpu0cLajrS7d
xqba8MwGDAoxduz1QjaPpgp1ps4eFuAUTSadN1HfkkYe+9nZ/g8LLCrF9rwKji414e0xz2Z/Nchl
voYGE5PEMoI2dxF0BueUnbYBstFs0Y1EgKD1OLfmLUcBLQ4qJc1fVvrLvm10QpT5OtQCBCfSPEYx
MGKUSBdhN0h7ngHwHC0cvVelxRlWBDJUEy78bxWpXxUfH7pTfi/BjGM7imXMyarfXMmC4eLhuIR0
5QMguPZRja4WfEAdFYDy8sBqU3mTkvDQuoKFB3VZ48Zqba8NrwGScqdnstxBpdnd3jya0DUOMoQT
+hs300b/UOGOd8cO+yHnRd+C9GuzZEFu2ES75gMkEodwzFmJeb/TsfemS9NbuYiAjvMX9Gq5V9tW
4sbToeJ6gWpb8+/GuE/XNrPkhhUfr6KjWkmlbvSEtAigCDfzUqzEpdFVinPLNHr0uAg4XNbbGd0X
F0oY+jHVucEXCBhAr2TkJad/DDRIjjAEk8cR3uKEORHEn2N5XHtOiMa5OBBx9NlE9Z9Tacb+EPwZ
k3O0KLvrRNQMfRFlILw5xS5NMPEf/w17XcvvPIqmDbL9jnZMKx39W7dcGbIcddCSsCxbeeGyIZhg
JpS3XR6JUCMaYWremdkWLc4uhwaFq4gxPz46MYsNEoHy2cAE4FjN6Lhqrn4jaJLbbyuqxJ8+OuH2
VxLk05ZBpgAj3AwEZkGItW0LgYQLi6dllQrPYR10w6UrZsB9MhoHNLDL/9LabFvuNNPrbE6OXWDb
UxE6kzzZMlC66Qptu7qQwXX7mpo/P+ZvSIbAWA+3x+INbsGICoNs/axak52I7+nyJSkzvFFuGpGr
PfjdWJCTO22vbINXOaskSUi3VhpXnn5l6tSaRlsH7EC/9fi0b9cUXXHl30DlGlYrI77i1pcDqt9o
wq8aHexOAA205k1XDmObBCoC7XLDhGkCSB+ojzy1+Z/md/uoD7tTr2DZBWIRZ+5E/Suvvk29kv8O
mZ9NwDv7EkNA0SjJZbQrdI0C503goYA51CngTXpLjZuHK2wVehx9CaXK8SI7ul++nrxsntQrZR6w
pLY521x3r9lOMsAhys+8q+sOOtDHNRo2tmVOAWHwRTG4iWEyZzZJZVvM7j+n3/9yfBhRoFrIBTcJ
QfpHNVRZZVJbCFQCDRVsxibw2gQyjH2/4f9RlmqzvWP7zzpdZgOhSAjEWz/+jrspU/C6zhBMVuiq
5EeRPvwWkuw1twnWApm8GHoaz5OXTiatyAWyovrjg0z7oYWl+7DgNV7C7BMOwAvq7k3gJlFqnLEM
fg0Yk0Oc/jBD2VzFJUEz6rp5MDjA9p3tePzGLFDEl9Ns1eaUcqjIQpQIU3KsSXLBYJGIxMbAsd7v
sTy8e7Ob4kCRbzo+38KHA5Ben4ET06dBVgHsBSPZg89vfYY0Oeh9pdoUjMKoJoVbrXIKQA9lyc/5
IIylAlQkPgED1Mtos6OrNd9ZRN+SjgKrqbvuintUSJDvBkpUL4a/w2X3MKDWNdLBFnK3hfznbh8p
dCoH0+pLoqOYkdwO3eabbr5GkDYDZPL5iVP9JDBB+NZDVHGP4a22M96I4gHjtA2YJU5QpREfX4PT
PDA7v1m7X5RaDXNBrY3kXAvDQ0V0bPrI1PFcrmcto43U0YXUfbCLEQ7A+dGCtwPrjPMhyqog5Olv
pV9ksg15BYMf10HY9sosrz2665j9Hs1gqBneHm/VcWjBlQgI/mV9U/7h8qxLViuq11f4zDl3ovO9
4sMYyyMS+eQ/OQFHZraJm+/7kxM4whz2Lv/PlDlXhl592LIU3rl4ejT0Q8/QZVHzq+MmXvjBLXIB
rLx0puoRHaHFMm7O+Lx/QcBM0H0MxqAWp1uRAWIPv8UOgrEtXvR9auo6rKB1m8uGqsQpgf0eGVjz
JJArCEV/xU7Ekk6w55UpU1esx0wyNVzkxAoAMHzywksb0ebUrf3gmXYHAT/dV5hARufHFKey7xv9
5ZChlWoedrg2Mi4akKvOQ2ZEDewkbyFXprOkucydxAp1Svyipe9pTpbXyK8ikDwj2NILkqInx2Kl
kePJPyQ47jFRGXE1LgBfVjtmAsy/5VEI4YJyxrYWsDrU5oGGtkZyGRlSpSTly9765uyVBRSlSei4
l938EqYRRwz0kw5QkhcPs8SPqtTXluucL3u23FByS3dV/vkc/ZYczZyYaiM0p9jKD53MNHSj3x08
tnjJ5ahxL1dSTDcL1l05n89DZIdwjBZM1l0od9+1Pfe8mK7Kqwxce2zerSuZRjh5XDx+Y6M1rP+Q
9GISNZ7VGZlWUS7nmY5Wkl0ATctDN4hzEuHHZqqxv4pbCgTEWVDo7yfNqwQofiuLR3EeVUC7VUOI
jU5h0ucezVxs/MEevpJnIkPRAl6WSL3W/752VHtTpaNZH7ESB7jaHVUkh2f0jRfR/cN7gf9kc+/i
PB6xBwq4e7/driJ7uvLadDOIyYa4/nGnhR/tUjyF+Yg1v7MVAdLHza81/u096vfEtR4hUq0+mfmh
LohbYyLx/9hHXzG/7iyMh5QqTfhAa/iTMwxfk9Y/dr7LrTPB9q/cWcrlp3jeu+zWUC+iC7fdYJy1
/lOvJKyaZ6HT8YDHmNz60XPe+6jhKQDbSviCHIz8A+z0oJ3JJcTtzx9+2BIPMw9xCNakewslH32Q
uiMc1GvxYv3RgSYWcPKbKYG1Ym2R2nndfNqQODXZ7MnEGnqX/6eHMEauW0THxEKHb6QA/v0T3BJy
Z7GkV6zuMhqOCt73ecZnwTwAt4nijEHCLXR5vWwEnrspfetkFvFk4ABOWAmMczDz8GA06bqS+/1X
8I5cz458t6r4jGwHSieipbDyS7YohGaKBeizVNJGK3CQ/08A7hhY9usfE4ermGDC/3JGZb5FoU+l
vJjg82JCcI2wNB+vi9huoGNl+Q/KAuXIpcAPKbsvTXsJ/2uOWD/R7yLObX+b/n9QhKiqxWxWrrXu
IYzsuV3bdHRYGrrOuSOZVb3xZf6JP1IuCxjaf3Rs60SduX41LzmoB8+4YTFOCS/WYCdn5GyR3QMA
uzGqFNgUmzWpN+2xl/mBxdKg/t71WYryVwc1oGt32hj+YNdTDzI5xVBKVUgw2/AEeFJZ5pF3S6al
kDPnNgb2Vp/rv0GPxFbTSmjcw7cmA3NWiVqEKMsazapDFePVZAvKeCOuPUO138ZYi87CgufR+EPL
SMN5a7XbxzISAe/pydS01OYckd4W5uvVMW8QjHlFMF8CP409ZEqVfFPdBMcuuExnX7yHpKQ1u6hD
j8J6xzCriZrLPFgxoxi+GXkjwbMyq1m4adBxTK2LhUnVnK6VB/vQNC9LZXu0eUIOBhnCOF3B/qgq
fFND+pvAYWtcY8lBD5MVkHrAEJFIlx1tM7vqneZ6lvpcHnGBKhxfxQI3rSZB74ArfuoAxkrf7idV
/+N2MY+7NKj5tgc6cCQ++MX/BmcQbBTxNN4Bv6X6055JztL2mMx+JgNg6haoqeHp8jKmKqYpNQFh
I4iwnFeHkk42k4VL1vKgQ28z7W0AFALQgQxCUREZ3oPR6OYuk3LSBAwJ4eIaoi3GUvdZCX70qydU
Ex/2nNWsrLHgGYzqWB+I1NFggEh4fI7krN25Hpk/r8MkQz5Dw09Mz8/cubCWJUEASC/8r1UnW8hI
9Np3YlL+/o7QcbW3PeNOgvarsOJ4Aq+YaapDcSUVlI0MJdfDttILbWtTsTDgzE5FPtvqfEdZWCo8
G7cNJGL2nXkq9kCeRZp6I46BLD8oo2GBOFc5jECNH0JZhyFLXGgTG1ehtQHt2x4d7D1HJaCr6Nq4
s1j0Vp6qG2fYn9iPNzA4gpJ9bZEzsAw3lXCWESAg6fHknnGx0coT/9OPYH7wVBQXNfSFokr3VsSZ
CSmP+ERR/4gbw+6m+Wd2N+ZVlDvlfnir+bX7VnAZYZwLodP6biwWe6MTDEtkPH+v1/ch5lR/REJz
P2u8MNqgwz3uuohLCQpCoNkiQxVR8j4o1gzX55hCgb0QSc9u1IhoGO4HNJTzfMP0xeUaf3XYCF8z
n7YRAIqa8PzLf+DE0ai8yDuCEofLZczMKFkzPoJeJqy+8XkuMF78T1HJ4Nzr5lvsk45iv4g2kAar
Yf+8QV/mhYtpSjefjYsxo7jMtgQlsGESZDe8k4qsH6KnspFRrWDCl6nvLYQKcmYwltsCuAB9RBxg
/+GBzhKd/jqhL2tjc0GpxMgYXWFszbX00NkxbS18R++tBjTPFjj9yEsvrvegf7BSBQy/We/55R7k
NlhbycnYzNGKq5E4XoTJEhqr7KNbsDlIWFaRfhJeID+OBpRIVl/w/VGdVd93lvUKE6QdyERaXKuz
U0E2iokbRdv6Q3mBTCFXB0KQalbR/DOdXTIx9QRxuzOOcB0PC6/OAnRObbFFtStUAMF+aeDQ9whg
Z1abp5zb7alAa1sfYfWEkw+fjZsNYG9u2bdtiXq52oBB0gmqncPfjFWB5cgkmxB0yvX+C5PJkg6L
RAUn6AclNxOObpTDDl2J/vmo6mTIL+5GCc7tg024OQZgOo/AOmVoFHzeROf6iW90S10wive1FZb1
UOHtBLgR0JUOwYpO3VOppJ+LK1Sp3wsRSlDbnaLo3utCxu1YaeoeTQCY4DeaMTv/WvWRTWuBI83W
RIKuTu4LY6EEScmTWFUEZoR7IJ+R+S59UxZTAGjURBfSNYTYOKsVszvuRHvonk5fun69ghrlotTm
PbwCXdVRL3Fio9GS1oQtt/A/GSwByv3r31m+41/E5LmjLb6KzA2iCv7G6bTo/pzuxFhMeh92CR/A
DEemZ4KkAq5yS4jh4h3sFnPro94cBT7RcAoq1YPwAaae6QLYelWmYA6yS/1tuWiNRyRJ0C/lDh+O
fTkl0d7Y/MoSWU0Pk+utF3z4KJqh3xPBV7Z2TpRVXqkGRA8z4EvOzkUcixNK1JW6DFWGog14OyRD
Tssxv4AJUgyokwsUzmL/yTjREl0tO4dlQV27XjxYrBfrmNT4YDeUZgho/TsdF5Q+ZwlrLv3U9jDp
BVpiFTDIQdkCPVljrQLt9kPLm+hWbXcU3/MRxBYrDqtlCRLoWLwkrOkTWg72Z7cgszaGLZrlhiwr
TdTSVmuQHHpyZwd2plXJ+RiLtASalDXxCDcxvQSOezhu/N69YX6w81suQJbgNFFOKKZ4O5juBZCa
lCiQfOI/si31R7lNN1yH94t5D2R3bo3StWU44FMJEdeNgx/Poc5NV1xZ9FkeqTe+iFzru3pqik6w
64FrHOWPevDzWOFQGtCSN/BgA4CZHGv93c8FTfTIA96eTencRrbdekLSc+4oQY9kxx9sl2vjIQnJ
oqiDjJ2aCwCv5MgSVzt461njevXgT8c3jJuT6a0RBsgv5Afvkge4183rGj/G4xUrzh8/z6nTd2GK
CZ4YOoSfZ8QDBR7EDPn1iJr7pBiSHiYlM/PWAT/srdmaopMiqmF/PDWi8xdnW0ELviZeK1FQmbas
x9OdFA3HXLJAKkTAHV5EBW9OOgoC9emZdih6NDgpCX81pV52Ewul0wctPKG85dfi2P3QqY1G76k+
ZMlKuj/2RM9A+/PZ4Sx7VifaBCG1Uwg0g+jeev9ikfnYnRmYRWZpk2cVmWSWf5DLy2iNxNaTh35g
thR/10jKG2fn4XRa93t/V6zwzpI2Qd/i+TRqxyLQeK0Nxt9nPtwVxC6iVEbf0t9uWPqifVmRBc4n
vSGlFhGUdZlV0gBCZ+41rIleAh4ATIYrjkAOOxWIdvClcz4gHtI+7A/CjCVe4ICF7EcfvuCnU9Q/
oSd4AnRrBgLgzBL0/HVVcEAvA4zFF76YEJqhbt3qFNr+X14BHXZoQ9axoaDIpuR8BTYqc0hMF00a
xW6vVn0tNxYhq6v/zC1H0yDJqWHTFqFr2HG4OuBpcAdNeTvEbYzPBknehapSMd4P2RLv2l9OhwlN
X/Z8+Rk6J90qIBChl285wTg3F9e91mCIK8MG316c8z3D9vwE+rmHgGoTYTuuEzdQC+QDFCE5+Mrh
6uQOPt+KjvfFkEKoV8c90GPe/DRypYb5/lVlgmJdHOO1hzNoZ1YInFSnQXX9TC8cSqCobkTixPp6
ph0LQDkqSj/F105DhHSWzyJ/79ARkmHKHZLAw7zm2yR62azFkSkuy6Dc2hrat1O3cAT25wdt0wrE
mPbw/N2u5b9jj+PGnnTihhtdRpn4x8N+uKtY/5yOFqrPmCpx/H73iwSHNpVM5USdhB0iqYEJ+Xb3
XPRdLoqZVRp0BaJfTTJBbtdTIofejMM//BSlvnttpH4KjO8/naXdwyV4JCyZR1QcTukQU6VSpFT7
dkiLOLV88rd7Prfz1LdoThhvwAIIovp7LRS/+mpwGTXuwsc+U6IIPTG7BBbiibkzDMI98werOxMp
jO4IHrWVmopIQAvpwiTnPoBCt5q+0wWylyh8rqJml6WupLvBy3ceAPfftJEjA5bMsofQLGvhdeay
B+uAoZlSYryTYQ9d8VGHswDL20OmgruGNw633wXrBj2gpKSNWftZ7vjeNvkrJriMe6rCkuHLLZ++
/OcDDkxiODzZvBP33Dx3IIBj7fDx10XRPdL7s/Tjd23Pib7xnTfG7FxYq7jO5zLLBERXxX0ZG63+
SOy7hpiG+5Xfn5mRga/TKDTRvSeBsy6vMjlCyUL+/4NNkftKWF5PbcbBWAmHTCWVytKKGV9RpfYq
oZaeM8ntdWHxCD/ixe6O9p3iF70wM/WCsoPt029p0mEUVWduDOiP4p27/ohiEiXpRIOhDNYUoGZ1
gEN3QzFjqxhWGA6qSedkgYPyrfAKQiTOXLra7GarVbXodTkJJ6yGoIWniDAtFSjbjaVoE4mKBx0C
wQLcCMoB+X4qWrIpmSgatxUEl6lNRtnhAHeHgbPn6xlFKT4TuMdG/cVXTk9qa7tLVBF1tdCMFuTs
YbC69BZBMvvZ1hk3J/ylTAFPqh9tLek8FwcZCtRfS/HdSXWo05qkihA6VyTRkQA8UG9j25oHhBpy
kSBw+R7lmuSuCn34BCfmJZeeM4mZH4Iuc1VmDNhqwStrpR72+vfscPsXNkKymjUcBXre/4xtlLcL
St7vULIXnMB0ywIxU4XNl5GFmUEWhFfM0cwmO7D/VRpgsjwgBblWafcCnOrBZ8KFMGseaz+vIrk6
AOT0ltbWA7fSQu/wJ/Lw6BL7GJ7FkBNaVbYxD4u22PiMcNLbgXO9AnKLWNd5uP611CdYUqVIAZWI
6egCyzluzXq+vBHwz6TxKih9A6iGmtbaQW4MDzyiUimejIszQqWTikTwXWCHxPtcwGCmSCDbtG5i
7XX2xf+e1SBnnltZ3OdcvPqA2MpefOsP73s+h7USa22dor8iXAavBY0X7TvK/zTLeJ9JNZ6fAUA9
6Eyl0VAp5KpzFwcg68499fh2HvfRTyLAeRbY3HOdR+258YzjUNoi2yMdhGvjujj9GPGrK8IBxkCH
XOHkJJ5BSp+njdOkQXT14bft0CB7v8e9LMrc4yh+YQB6BuEs2Ac7HUI6k18GPqQ/VWnPAqatMn6J
AZaKUcIRXMrV6OAOngfIEW/5juyP8XhZwbF5gQFBBaPwRJbKUrgy9uxp+41BiElb1/ZlNkC/BdSs
SevyVFv5brwYAHtZOutysNVmrcORBsmaJ1k5sCjj34N82wU34u5GglLyUO7B/zMtMA8G67omg+Fk
uu63jmBkPWIM7+jSsuAFc3KzPdUqWTofE/9zuC8c+LwIzgU3aRaQv0Lc14Mhz6tpbNwtbp2FMBAK
rmz/eIeE/l6hi5BDByjD9mLtqyTSh2mt+ObWSVTReF7HW92xH/b1L+nDvEv46ufZqp+C0ZsmSuzx
neUciJaNLJHZ5D34nlyMGaUacNVC5WvqP1W39uu7bGiFgnv2HCRGy9BKnPVM0+LfQoaKCbzrd4dN
tVYjJS6XFbyDmFB6kkWBUS72rzJu+zlhWxEsI2OzhQYRMEIWAvoQw37urrw51Xih9fii/NemP3MJ
1O+SwKZhPW+36Fq36G3If1jrDlCRAoq8embyJvrXESQnm512mp3Z7Y7aXRmKx7qTm1YI4YTkUAn6
Qz+WnpUAVzfXzfL/cxpAvMnp5fVWaQKQZTgXp+KDaoxgsOBfoKFvvAtiDU8zZ8Y6ojEGPss2v6Is
N2oEaob1nR9V0aOnwuUl+YhEVxqnShtmpGm8bJHI548ql0IwIB1etOYmI+vK+GNJIypF8e48H5to
+N6jMlCzJPR9dai3I47/0spaFHEvxKrk+RZzyDXzdcLjgwKIVM89896enmmEirH5IQnL4p+pGjZK
/huE4iK2kHKFGWPYlXfYbpmDOLG20nYFgPd3X2ayHRpU7QpsfeDTMrvnK/oEPKz3q89TQKFKukCw
Yqj+efPNvL8UsWJ64R6rHc+KnKfkiG0X6Qu+o0sUQo5r+ncIvaYA+6jlMTmETChdShZ7YHgmkyl9
ZRw4INUk+mus/fC2A3pCW9re8/+A9GvIDGYDKHYSDXdcVnd0yR6zQPpexrtI9McIT1fJ4At3+BKJ
6mdwZL4ioypO51wrhm8DrBn4hxlyMYZ/BviAT7CMjpgc0YsQ9MLzs5TTEk0IVmmqnL5WXQDS0/62
IkIasqbQ1P5Rk1N3iGZP717QzeYUYr/7CzywmgfgUQ8Q9AyjTJXrezJ7S+auU/e0vkqAvC+vSGNX
zgd9vUm3IXKhmOER7CZMEwGu50Pi36HIn0n4nAQq7DGx0MXAG6isU9tfNGBYDokDt1IOUFAXegFc
91sy/K3v0TBQw+KktsqxCIUiaEgiqacbbJnYExCeZI5FHH5zGgU+3EcJrPTyYqiSVed06c8vHaol
Yf3YBkKzQpyeEZ37zoDD74J3b7Z5Dvj+7MRCPWBdvnMtMF0PPRbTog2JfAiJIR/GI6YgOm4tAJpL
ZA429hudyjDPh0t4sdTXcPLn88Tz11cQzQEUbsCg61VCNvbk7GxchIPiG+Kh9/RfrxOLfSuft5zJ
DuWsajD3nOAY3xbjGKabMUqt3Ad1WZNhNc3mgfHScNDvZBAjUzCOunwPLicUVNRvwLx4BtBmeAa+
/0D9vQtpJvg89C2GylySiPRuenkFu1Th7hiROnzfatwbKfz0mbXFx87CGvF9F9AMs96hxo2Gr2mY
A7gXlKROrdeQviS4SeDouAjNj91I28SvOIAWVj+xckl8K/uUk/z4PJv8QuZCxUgJ3VkiXKFigbK+
pevyV9qrw++23EqIkE0AV4rYppR4JLuFHO5IB4y4Yp2ryJENdU4euUFMjpb5KBSvDbI6hcMZprnD
u0mVyvxvOYFhUmvcFCRb/VRMglM4HQSTJn3zhMb/+Jr4JXe4aDmAKsNSNznCvr6SEqhwTMctxYvw
rSQ7WlFm31eXv0Id8Q547yRscgl1Yv5tchNoBJsj49rn+8z6f9+Ex+qn/MKnETSFmeoSDxW5KgVn
MSg04Vg+MITcRc/a1Lhf8NcE+STC2CNhhn9jHTx1eZQvUoA3F2E5AyuMKMSIn1KX/2u5F1B3F1C1
pJubf4sIE7pUB7pNw87KhLUmUr+siRpsL1v4QaWWiEeSaL4DcmvQECjDWUUS+ikVdaicGVZIqU63
fp3KUAeP1up+lgzDxQy8IetHMCFmzOjUunoM7lZtYqWZHnW0HV8/7PlGNLjJX07DZyTGtji5Xqtj
WMWSA/yEzr9tZCXDwbBiY9yRi8h1rcA2qgEsFuj6EAOXwn4ifB3fn1EbMSH+Y2Eqo3DU415VqfqZ
UqHghZz9UhHo3OpTKHpxFLt7Nx5B9MhbUR/UHJKjLJenmXgsx1UCYGQa5hKiILfdDRlbWlQsQKia
37aSrQDaPCeDfNi5t68BgTnbpDolPN/RMR2HR15d2Hjb71EPjNgbwEKS2Jcibn4XjVwoYIqpe9ND
zCPpDBPvm3FaveRlw9Xliy33TiGcpQwcOPBCXjfWt4J1myCu5tqprftFOc9Eqj+uHc3BaT9gUtzl
sVgQOqQ8k2UIxTvAk6vPGwNWKzJPe6XThPAtNahqfNWBsKXceaDmGaxejJVLrh7HMKN4Fr/uVurn
LtFwpPUXuyx6+YjLhM4lQhyrpQsWie16Iw4SEdRjeShLqvIEjgp8k6q6xQMBzT91sgX/JzeBt4fJ
IpsuEcjfnZfWaRqyZJWTNOPEzGOMnXpGkZBZpEA7kkraSff7o8UDeSk80se1s5yySuNvPcGNFrvC
WHwVXUofwea/lafbxML49zPdkly54JzNBoUJfszCKGB45r8dy/m5AbCLw+XVQOa8R4qW+SoXngSc
hAvFOnoV6UKjFwq1LCsdrUxJ2AIRZgsUQ18W/ADRd7Wv5/DdyxqhR/SG870mNOLRdDj88XhkexWi
7i7ZGOO9naASN0rfVjKw0C3fWHgnWQ8p94kkigRciXyOSRBPo3TK29HY8xQNaznyXchXkxxFEcVa
vu8G8O+MmLVUUmFoL+8gQiQPMW1bUW4yfIRbWPf2ZDiK2U17e0mJnVQlW5WApDxlkM1QphgsIMMG
96TEAm7AL+JpIQqJGCPWkXgjzv1V33rsgyLt3RkQkPMlDh+GwIVkK54hb+UOk02vGmDHbUX1H5CK
z5X+7ZklSwHV4V/GBL+e5SRM+ufSXFXhab7zrSJmVdLqYjj7GJv6zjZ3xIVY0R0ZohWI6xUVCWfd
gW1bXlfOmvr7eN1hg7ASj2i0HOJ8yONf1mgCXGmZkOgG1Vqo7nqfPa7RPv2cEIigvc5X0vVNDd37
mhq/wFVCrtG51UeLuK0T+7pKq0cGj/ZTtlIa9uqdlgo507PIkRxTUFkhWChpg4U9y7XacRWUSapm
lnIg4rUWSuhi5UFHS7Wby0OAKIzQR7Pi6ralCkGZHE0GarXsNXxkS3NIMmEkjY26Lk0jmDq2Rx1/
kT4j9S2OJ+bS7SVmDuIpipq8GorvuGGUExJmoXf3fJHcelvV/rKbbAtFzh/zkYtvRHj0sS/2kZdd
kqIZ2zTKoYYnF3rn8wDk/JmCQ4fw7GYmba9+gKqVgNQMx8nCzXkTwWyCcq01OpyfBHe5OiGtmNoj
rgAR0nOXnfC0RZKlIg/dP+eQbRLLZ4JwhTGyo4qrra/zUUqr0fC3px1dQKtts2kUJmgQtP8/hsHp
3cjw6Lv4N8Hyllt316c7uQN4Vk6bsxEBPKARoj6ifepgjidZPQsTIX1eFFEin1t5cuXEyQZfKUtL
/1ja3O631jU1mMJNyhAeFCzAbPCyI7XfRXxgXuCXKBhT24hEEzqjvZHV20wq0zLFytX6ipHtCHdO
xMreHbmUman4q9DmoDsNoHjuWtEY/wNIp16/R4/71/WMjbdlw8EBl9aG2Ho4Y9fxB7C5dky3JQSk
sGS62KuSa4HRjnjHpWGJy6zVHcYhV7LEbn9ZQtayaw7vKoqMJrdjugodVF5uBR6kB4aLTRPh38nf
iyOK06eyXxkodbBTnNr2B3ze0W2zuAncco4+dvuFUlviJ5Uy3MhAP4VZSQ1uY+nAkz7PxzoonwQh
pkgs3EEvSEPMbA4D5uzHZc5KwjvqTS11efLW1SuSWp7ym/EvxtWi/CW4VBl9Sg7R7u1MQQxjQ0OE
i53D+QW0Bic8S5/7Itm8pvGnJa32TpESgHQuq17IuyRpqbuCn1q1b78cSZMcxSW6Y5rH4frgo4mn
6dIrNfv2C+8+LezN2JzfaLSL8oJzeX+vVGCznlmwU1Zd6bmqnBCiLQmFeMX8tV/zNh5o8vCheXBz
7L2RAzWcapMgakLVODPp3g9XLbcEa1bZ0kCBie4kBuzM+27mIIfJQbVZdkT9B+ch71AdqlIOyBdG
YMDuleLGxYumsPJYU81gZVNHVHrcsJHBlulUncBNGcTbPfSkLicUHnCM0pIwiihr9iDFXGmaharT
WrKe7K9p0ZDSunQwJZt8KDa1y4CdULhANGyR1agHcGakV3A+sixCFucvjNeSo03XjsAIm9I16WVE
lH14FPH1YNfBy8M9En5tTWXd0w5kZqB8CJOKX7Pm6jmcp7mRc1dvYNsJ2WdlBAYhtLr5fdcPDTBY
Gq+UJsz/FQzqNhrmp7x1IDrmd9wDmmjr46WwL3l7iZ4OGm1zCTv+S/nYoCUm9Qxd06fOcveX3w8u
a2IvLoYBIebVdaiV6ZxTFVpdaDKJGqxsSA8dMcDjGAy6UqSQO+OZqlmQbNryV1G0FBhOwzE1AgHQ
TnbNHIz71sUe+oxPJ6W0EpwzfA61lTXjcv9ugELSs+GSHtrnQk3+eyuVePX1WkAzhzs1ze5pPNrt
U+q/04nNjNRPBklSJE4AGGIBrZeBH9t2dBS7q+A1mriaZVAuJM1fW7S5GR5n/LzDjlJImS0CpNnI
o1KfWHMCI51q74wzzGCgmRe2nGaeItgLsW9z/+PBy1ps+KEPnGXeOwWU9DqvUit4FWVyh2/QZuJG
Mb4qcvn2zigVB52o6eH9HWaSTp8UztlLbgeFUzsVX5fIP/DsnljRmFFC/hEjHHWDzt5PASyXBzAZ
CL4yJSfKiimiXjGgzfPTVmJX9OHrSqHO4KP1rCNIIIxQy+UXRcLWuODVZEiQdbf4ajYscLr97X9e
Jjp1I218PLb3Z2cffWlq7AbMSQFjJV93WQcoyXfKcc93npkXekYTfg/148JWwTdfilUYeIKrmHps
FKrYgImdhKO0kdUiBYR10CpfijTjwMOHXzO0ENtcuGSFKt/F2ANeEFd3FlpaKIuopqzArbQ4QZsx
qCeqQpxDKId13Tp6xNuxo7fc3wXOb8Se4rVFKlOe+D4zKAiOKyBXS1jFMLe6r4h5P5lHYzVSDq9e
zrl0kdLWLSBgzWD/Tu7o3w8Yoe9dK/beZot41uLT2dIRuhxK+NzGsUpKYOWk6lXsvyig/6wtEWli
2ARIMD67OjifN5gtv0s8FBrXdyOTWDTKend+daqYz38SrxyRalUFwYSZSLT9xX5ZNwaTFpwIDiyV
EvUQHMC1qOPXumPcEv00ZigVrno6nGKmOV2lGwbBQJTCgFTpPZZ6/NxhMtUfZlcR/edIEn/KaIMI
869sGHSkymE3w9Uh3R3xMzp5hAUgF/1WbcXCRfGjQA2EwRL9FAuLDGbpQSFFiCqZfNBUtPQieKnh
cnZXom3NP2vKKPaO2zKPFx/heTPH9yVVHU6vy68JE+YuUUscOOotZGUNZNPhlzptcsn118MJgCdW
N3jBb6zLPhW+NSiGOLfdo9t9MOPsUbgJmpiTiNmXGYgiRWcSv21w3FkfjW5GZL7Zt7K2fhGeAY4+
YMMVMCxF5IUEtpNB17cZayZEk0pazWPq4EAFOT03y2OHuN7HQZ7z9HXoDhoSCDenTB/KYY9mMCUH
9NfdBsg+bBQTDIWP3pfdlbKvMrwY66/plrQCZ3o6A5WXeU5QeaBG8HNEZ/PhHY59N0gSnUSCzunH
xONDvYLrIplt0bRhl5xt6kxZOSQqKsYP1THiFKD1W2G7V09HCLKrQDUKmvTtFJSodOXAB38g2TFb
yodQsG2WaFX/oeaV8FxylNPRy7Km4si+be/FNYx1BKXTUlNxjPke2xWyjIvyl3/STEf5E/g9j5f1
ByxstG/Xu9lWZ9UTRmEHLr4mGjjiNkEH0r4tR9jxk2YeqPBt94OIjRY9LSNk3x0UPjDw6oU3YDWT
PBDePAjPRcVf5C36cjBD7ofdwlViKHqZV86NVjIcJxXQbw+y90fuoQPI/LT0yMHylls5x06Q7kcc
rLgDaPaxBbNHDdv5ROmlR/zoHu1SfiWNy5E88QtgS/vXOtT+pZuLNr825O6W/msXO+AlYV0tYvbQ
dMv15ECAhBSvNS+lxPOIYWMJsuHkkMpwJ0eFXFhV4SqWpqUbmcJldHZxs3IVeiuIjFQ9AGSKgJ8B
x5bJccjyFE5uwwV7+02gIVck9pHTmR2tRBcbkRuyWDCRvxKLwh8go2RbYJN7dPx5esQhxmdIQrdJ
gb6DO2B/1q4gfcN9TV/5PArosvQztVX/0HFKtLYK55tgRDaA5oaw4xfPAYpjZltxmaPfds+IGTgL
IjR1add9R/3Tk3uitedCQO8OL22VQVRze0vaC/2uFBPyz4g8kSSjXgC4/RskR5ZD5zN+bqTu4VY9
+yLpzHMPDVB+2jYJ8CKB+Ym7/c7RYfwczxa2NqeUdXBIEU6qBfYNtdWzgRoPkAzS+OKxRtc5zwHE
L35z06Fz8NJzKqeWD/TD+JaeDomRQIufYd8A8NMBdtZmjunMLKaV42Zpuf5s5YMyFhKr88yxTomL
XebsvfVQONso9rwoZuZ1M415fRIvuBFd3TM//d6PbftET5tlp9k9dFhWwLOQE1fRCFtjpTyflVf7
qShjNBH+Qfa32wYROgZIGuMfjbTx3qZ+Uw+USpRAmAWzK9u5LRRc0JKMMXxlLv18uhvuD/O2KZBt
qPQwex+HceVg+NprsNIaMlulewuEeergHOdpRqglbNetQjw7UUQQrOybFC6gTUp+TfLWn2sf+cQC
M/Mk2sYXE6K//lFuLdQduUq2txsJv96WW9g4czPds+vNXoPUO0ifiXPfgVEfTdFommMt6TMAvctX
S7Xv4FtpfwscR5yIT7sayaTrp3aB/ezmFMFnMIXimXgSgKgHi9oUc7hHLN9AyCXR2i7HtQgWfhDa
WBxlnrnU08vJldPVgq1UFd/i8988XZ0NaNmWt8E6WRG0j/TAM+rbLG4Hfd6DM5lEzdlsYlbtSPV+
mBvuGQ8HyrT6hO52lZZNMxp5OYCFHCyMgn+S+JdnhoSO6kozmxbb8R+w2Nq7eZpk4ZJBH6GD5L9w
aOnBT1l2otnTN37UYRBTAiDUGu5lxuuJRsWZAKyVcu/UuFp4BU4Iqb6P8DzuZaz7P4ZETl1HebH5
iSmLNrNoxM0nJsWHxhCXII+XZ9yLOBTr43szSJDFi3mZxgIgui3lnOHQcm0CpV1jn+m3K56Q92tp
QJ1I069U+yetrvviGa3dOCQKOikMv9yUvea3TAQ6IOat30xFQFRlH5n1a6mEtjBHDljTFLTzcC2U
bUmXWCgp9gLN0l+9lrVIiSkfRLs9RhNfxUgb864odES0veCWGV+JatHapmaWUTv8lVRL1y9k//iD
kVU5eITgY30cDc9ywqwLr3nxQ2oEvz+Ocv4mEeseobFCjNNayXvZvf4Zl2Z0S/RNnXgvF9rscO+U
wj7GT7w6vl8MjjhBt1aDKAGOVmdLxL231pn+Tt/W6vn4BLjIr/xVVSkraa4hy2nnUwjk58R5F3LG
2IptUw0rGzsFm13/mOCInptXvtMsa0QaPdsTaZuu2oaN/K3/GU0at/iPe2OyH9Dkq3egu5sSzLPw
HeWXPuqgHKmqsfc6xxl6a2D6bqgfzsDCEApXBYjiQ+jSDnKbbtH+ALL3c7SwRb46tqgpuxyVlktm
WYSCQKRwZZFKKgLjcBhv91vXORh5QH2SyG04Kznr3/S0i6LSMkVOK3jmP+5ys1D59+BiKQAHpPlm
oHkkgex5DiMcsPAjYZiAAxaiDOOcVKGxHzx5Lf7Lk7zBAtnTnioCg5ZGLxAyPrcpOP7CbTOTvfDE
nfuCw4/d4PnKhXHZAz2AZfhJutvqWW3JgzSQnoDvOQnabknWrVxzqAeC2sr2extCiXefe1TUwZMH
r3yFSgPIAVtew5+ms0kEgOIS278A/a8VRLR8mxGft6My4SZ/RsbPJNhRAi9YpLZGeuvw9koHtZTi
jIJ9qtYdRj3nTLvqg/HxovExjK614XUCy4FZwTGD4nr3vtgYFNx80w5f/TTE/z69XCfRy9ZWM77U
q2p1H6sgSf8GND3Nrf2fM0WmNGPq+VRUqZEC7K9s28Om8M+9yC694l9rqe3DtQQjEf1ZiX7uDlo8
Onvc/2LY2G7sJaAMj3LMU+hOzM6i2DPbt9yYvrnokp92v5nL1HoB1f1vwp/k/ChcBDi+QeRYwaEI
llNHXdQhS5ELTxmmZzTOx7AlAI4XFR1IkKRAKQaQXAcEdKZkBxv9vb7D5PdY7AreHymdge+TlRlb
+0RTwkMV6RDjfTRiM10ZnRdOIDTYahyys/TmlvUpNbc9FVUuqSH2DlKWpmMFMeBueNsEFgcP7tAT
ci8r+7ReIxPJmonlKSWv8oqinw3x0GXLvuqsogLwBikMDTlpVXUYSVkDb6PrL/ZhsOtevyoQPGMB
JDMrZZbjU8MDUkqboj7hNAs+T/1yfBcC7YOXe/RHypc3nyE+WvQMTnuUZ/+c/7xv9hiLmFJGgTwU
uVBbMV7RG0le1POdfl63ODTlYfC/g8mLKth6yJTcRoJ86Lr7D1FU2COmguv0PUfEedP0fRUUqMO7
c7SDJy8+1S1i5Y6Ig5A5oGh46vN1MpA7OQTlgXyGSbwgTf3cpSroyXA2I/onz+59F8GlN8XgO8Sc
jPRdJaSxPlI3v8LDMYtm7GTBNMfAb1k4Ad/GnEh5e9IfykFlYfcLJ/ET3WUs4hauyE2p4qp629Vn
3mrZ2RicLRNi3JO9x2FX6mFt/Cr+BSkMnjml9bYJGMomG92CVNi1NyhONInEYshsXjjSsifW2/IZ
39a0ZD+aGZX3U/JNB7/znEk43MyM5z+Sepczds1MiITMGYAwduksewQJA0bbYJFHY8hUayJvRl7g
NOesfvhahavKmwLFyYboIIbnhD5lklF/zT5dofr/07kCF00lJeZugojFvWxH+eojXW1RzXZUdTKa
S80vAcPL2zrEs7gajUlDE83mZbcp+M49ghtnZY9yJaeAAz0FktTCEdfKkhKmtz+SJgE3R1PJdyYF
tNMxsWRJr0JaZqXk0qaDbefu4vcGPzvK4IcGnY2rxa8u/wUxAlGK9xf+O21v6Aq+2EcUMfGWKbeA
XVCaAI5uWzBNqn4qI+A13795FYdET0bMmDBHUcdgurUlmODAPeWA4DB4w09D2CwWNjCl0Hu//fye
mvL9OVl+wHKS90GEtXJKcQw5SAB/XOe3plRRE3J8en3HxImKJFGDzDAM0KFAi+QjxHdaxjNV0lVu
SeMYXXz5+DVAWMIuyfyGTHfRKP0yKY5LQ+dikFc7STXDvquhkBHRWYEhd2s335V5UrAAegI5Q0jJ
3YHu4s/7R/jh/3WuBJrsluCoRqJZHbfPhaY63oX9a2OnzSk2a4M04GfYMPgPrN/pb2X0ZjUYDTGj
zJidTPBCxKVul+/nQ5Ci8XIdD8QwcIAYjE0GV2WI71nX6y1jaNNHB6+M9DJog+Iu3npraa1FEuQc
arXsDBkcAlymnC/HHkR8a4gBwD4zdQCpwM1J7FpmPDNEAYO8V66bwUi7eDGduaeJsM36P/poMaSM
sdbdf3ByMXKDFtUJ20kHX5GtwAY2W+A7SxDTgE+qB9xNtkT32K6kpFyi00w2req69D7qHunkMcw5
zn7A5SO3ylLzyd3WPFdT93DuX4nPNe6gDTRGDNKj1LtQMNyg96IqbB/iSuU089vfNduxU1VmmBCd
rXqUNuU0hW/my6MwUTo3+x4cizBc6MmDMEpeULBr8LIZdRakZYVUjUTPtvvQvFrm4cKXjamr9U5W
q4DRchdUrudUe7ErkYM57ya0D8jLO8+56MdX9h6l8q5eRfE0Awcy82m1jRzyrXowR8XkJt+azAOK
X/3dqvE3ZLTKR9lx5MnXBJx/ACtKWpK0xcEHynWbAqibY/sOexPWG3RJ4edzx1KIvp/RxtcJ5gv6
7AYEnNb4OWgrHEDNg/MoT+iG8j9scI0QUNfxteGR+aWuH1J1e0cI+xPYg+zCphyuEZ78ebiXaNWQ
q7EFo7qIISf4boSN06ClTktmuTmkUhlqxum8zfmW5+ivwfJenHm0I+ZdJhJvnclMGtEDnyHqyDZs
sJyMwqqmEqAuJ0HHJwjGDvdNWbd/mRwZVMiZ/Ra9gDYqOBUmhs8CiKMQ1CqqkVZtL7lOGJVqPq95
V3e8HSmqEotclwGBHxvWCjok4Khgjvw/014WervqjIS6fTBRnETWDylUmvVZRdoaN+Z4qKDPNEMb
ETLpzY3sa1pvfHuRBnKVHX+NgQWix0HCtQSpTs+wzAV5Nbz3lC9+ViBtqUzdHfb4dF0XHJoOr6Jr
ir5Dc6cg0o+auy0/i+fnkVCbVUGEg5LaxQSUSVIKT11513YRhXZa/p0N/sasgFkiVq862bmcFYMq
7/VZKgowvEptYaw3s90JQFJlKjkjCU/LowmQ0HS0lPUKTU6fCWgjgBMe7rI5pIKhaLT2/Pl1gbfs
nNsw7aucLnnw8MSRTPiSMMJCm6N343a3cYbI8CC783xlrPl/bziIXBI9DeSi9w8456UTqCxBNpWe
eJRWm1nf4jGn0NEUMeKxC001qj7c/P7U34gvi+lgRpgnm6yYjBacb4WSUDDBtLL/GZ7+ljuArJY0
jp3ALd8SIVx3taRlBNQYmfTmoPWS6QovdML+Rxu3XMQ6vgmdZ7qU4XNW883mJCcucx+NOp+6it/P
m97syYxS3GeeqEvZnrYYKsFsPE1CP1gYeI13JEi3s+wv27HF/YvyIWWLOqJfg70UJ1kabp6+louQ
sDw+Tz3POOEYFG74rBfisQ45lGmL5+NNHeqyinrHS33vZSxJV+nretNoixc3LV+mn0Cv5jfpjJ08
YluwCIaKqjk7qsyL89iZ6UC1Q/mXNcsy9FQJWh7ymC+1RhWc15YstJq8OOpTInMSRViyyOZXoABT
zBn/Al4+MNSX7den00vWEN049C2FgDSV6YW4m0/81g+nFWPFklA49+6YNNvktdDio+TJVYmbFyrC
QPsMsvaNduBDw4c+96xc/dPmcxslqMoq9Msb6+JPRCL9XW/jZ6oVomXOLhhn5tQdue34C/24BTqK
X6U6+hNeApu5idOw5lk8WJw4qN9/Tu9diK6gKxAgsJTdUivaMI7NdXlHHCSfsXRx6GHLpono5d5f
o2NtTMdnqAk6C0R+VIxFx8nw4gr7116mRHSO16vS87zlCVwv5xWmcltHMFIEhCK+KXB6VluF8gKp
f1d2U1iTwjp6JHiDltfNEvmOIKaVDkLy7PPXlRA11UKnt7cUqbbHgdL4SzfzkikUle5HfxB0l7xo
khmKa4izY1tXYRLrZaZzXcJT9otsZ3j72WyQ1R8hHb89qO9oW35XjJ8GvmZn5/0UbFhkLIGGOldo
pJ2iaClkb3Xo7L3/Dr0fAtX7ly2EchVwoKXBV9NfyMYLb75iaZMcVdI9lx4p/RTtN6+kUdrS4lJp
Hn/GzHIrVzfhdzA9gES9bu/v0vv+h0++If1qx10yMgT2WqPN86NKOft1nTaoeP52u5odQ57MPqE9
8La3KOUmOocNNfrD7meYPja6/a1OCHT04Vmv7uavEoyqKlvO9yEsOr6UpuCbwj4ssGOf6W9iV16d
ZW4TXiH/BaNFhYEggJwEPbaoet06r9Bm/Rm41DOpSHOTqSvG1tPKJ8M0/cWnnqjx4CPqFhQqEHpf
1vpzeEtZIw3759DlwbFXgYN+c0JBSizPPTFiJgkv32Gifj384SLY3lMdma4lCow2jx/ePujhLUxK
5AFtcWgrQQ8b6/qQlyFIZ233fh1wEj/YN2lijKR87tSwR53uEjXHBgPMp0weV1PSJZCVfla5ABEF
g6JM3+bLFmmqnkWzLeGvTdi2xHlGTRPuR6QpBotfWrhSlZH35hXasePCLcHZZ43bW66gSSb8AdFL
sDk6NWySqU/DOXBP0JhBFnWzNG7sR2V9aNUOb+heWi2/CCahdspBof/bcv9GOXouW5CGHD4ko/yr
IeROhEd8KAFxqrT3qN5b4gGNNjUwGS/dX7wPnO2+lqSM677ZjHpTQnXwzURRGJpfJ8Fhj9a/AgRz
ivP0lhLW8Rv/iBDoJE7SVlk6NOzhcmINw24NLQPuASbG2K9TgwSqrOVliKNMD0MiqeXSYVcr466j
J5T5q+9vfFTJFdIuiXl0IIZeeNzuJuZzE0QpN8rPREslRTxBmeIx9ZP4y6jX//02cMdVRS+cYdew
h2GjHGfPcaxFKHj7tts9oxYdfTI+cXNUyWfXLYdPT/9xEaJHMVyd6AVABKKcy9HKO/Z0SW6N4X/d
QHil4Pol+HDJnP9rPXMXvdxK5Si2XtuVbADB5XCjiCsUaVQZbQffs7jI0NE4NKeRvAEhFROhBtmu
2pkeWFopd/Cll9n0fhvmxQTWDmU0j7GRYZBT9plbIy2vCvtZhnnUSASHPHAZp70Xxg0wgW2XFFV4
km4Pu4nW+C2dAqJ/BRqwlYHdPQjMPPzLX8ICXk1kL7kK+TyKJElJ2V63Beg4clrsYP/avkiPWbuL
ZB/d5orZNqQdnJMOO63ZBodMQBcqGuv6Gz2CbEmQCkfo0prNQc5ymSf/YRQmj+cLRcF/RzGkobXM
NwLpvCFy2S7iC62zr6Uk7AB0WSw5+bAyQh77sY1+3UaMTQiktbq2fHCbUbftszBpzoNNtcudZYc7
u8cLtLocjTaQQWFNbGzKaX3qvQBtYOc/wnFElFVj3TKmuU1Zr+yauaPttyTa+A/qhjgdAV9USvds
6U7QfyTsHQH1dZ6IJsohWDV9Zgex2d2Q5w5EZDkkI1GUBGFa6TmAFHG2e7nIkkoDRyZwZKWASPhH
1hnk3ZO8v3LrSUVM2Hh2a66m2jPtXN4hlRT1ZszuQMunGLSg/9fHa4WPOnZrbDIaZDcD5JqmxGR9
VJBPRK/wpejXJ9D35gzKHmI92jZave7wcRmUvd3zjO7zp5nSr455mN3exuNH1IVfpQDVMRdTYBFb
pODkYAh1kjZTe8utv4cwNR4Wxl5CBMm6RVFHfpMHd53OpqjhciDcU5XLrQ/qXY956nATeL1dRHGl
/i/VN4NYqP/MdTmuGuyW6HcqWhzISsFrS+1YaSRNVFbrUQ0EDmAtV7r9UEKbQa5X0lJADc99gC2v
q3bpDkCJU3m8UYBVggM6ijEuRMKx4tz75vuxKk/lwkcsQPqddE7SeaXLoNHdHwI4+z8DT61h3M/5
e6HFKlniBV/rPDSjdWVTqmmL0m7QeSLbF+SG1a2kEKonCnLRS1kL+vRYsWXlp9E3/0H/8XF/GXiR
D3lO9aA3q1XLOs9TfccFJr2Lzv7QrqO6f9lTDeKUjXbgRwaTCAhZ8DkeQBq5o/HEfsdN3dHWi/5W
fm1uwbadGKVoTHosuzD8QQh7cgJeLJNKZfOGI4eLKfkX8oYJp6BGXeoQR3YVMxgaCvSw9uEFeRQc
PhkrPw6+8czRa2es+IyVgZHTLjGD7yUKW2OQIBPFX183XWXIdOaQcdIlPlLidHJRpeOzqHQJy5Z+
IgNKxcUKvPHAG64900+B8KWs2bBn9tchY5iVhvP6DEf6Va2Jk92WAsEPNIKxvatKUhZkmjeNb/Pb
9cI4B9PiObxWWfiTaIzQi6QWiSv+IaRRUCI4rlkB21IdIR887VvOuHhyvBWKAJ2FjHMQJkTghRZA
LItE0Q6RRBm25RD1A9CgB0PNW0Xd4c7QBoPxDrkko1t/EGekJXontE1bWik012mlybFU7jlH+om3
PS9tM8YKlb3Zfum0WQKlxfdTs4GvsrVpqPL/fotx+K0pgZNWj3x7sm7IRz+za2PLyNJhTm8xzF6J
Tw3Z1Teuap4iXbpZFyC7O5nbyucHx67HmHTshHq2Wj+WweKgldgpm4NnBi70PFZtbK0PMdM4wKXp
WZxeCTraWr1xDpGGGqjlhc6pSfir2KAMcfeA1VvZ08/D0+Pg0ydDJyLKeKWMLfaiI2y7sF88258c
ib3sNGxVS2BIsYfaT9R/KwAJmaYwbTYAB0Wzo18bULiIxRx+GQ125VlbXtfgCeuo9dQrx0WJkG7b
qkHoYh6cRox8k0MMtzPit+CJmvTjr6v72RHuJExAV9hBftbCFMXbOUc03+Te+5R+kPdrve5cvI2i
zBbBSIW92hVrJG7M4M6mVEb1anbyc8iwi+7r5GreZumlhj5QCkIbwBNtRTcqjxmrw3MFLNOQ9x2Q
93l80Xycvuxhv5z8oCA/SpbMqGo8mGv9SOsmFZw4iZ0lKZS9AC7cTZfixzL0w/xzfYUFJlUpjEmy
1KNd4xFUnYRtMWhW7dbTQKJ+EuVSMEgTmYX/yDl1MbozT80SUJEVlalumxdry9MTjCIYW5oHZtEh
WqiMYF35lIBi97p4TBpJPThvi2vJZt4fZvs0wAiu8X85UZ0atWSYWJnN5S561GCsmcOAFE0o1QJH
wFV+CRbo5fFeOZ0KhZftGeZ/CD8QoTWEpiVnSEdTu42veRM/CmRTyCg/kob4RMTNstZBSFajnEop
MgedmoMDkkWmca5BirKu/NiNDctzxLtcW+mJaT9/C4ohg8PjLt0ncz2mhBXnuYoyfpuTDBYeZpE9
n+Vxi3qI45XhItKA7KsPRoCyJLZZOBaBYJ5LHH7NrhUQxCg8q4NAiImtCgiMmHObDS5yV8udHVz3
63GB5CeMXiZLUIxT6POeJ3sOHT+lFEdCFPW0dv1DLySdzAodqDxJER4XRC4AJJ58v49AknRU44+2
uHWKFyZEYij7D1NTkQKkc1zMB18gagUwTlBaGJQh+Erv/P8O8CRQW8C8SMaiBGdN4ErTAecVp0i4
wiakE0fRXc7jr6B7pzMdkX2b+O29qADezewEViken0R/r9Ck3ZAVtyl6dS+k9r4hx3qy/RpgU9oe
8TUYwMnPa7+OnMyXk/GGmljN+X0b/o2l17p26mxRmJ2aWSXsNpJBLCiiQGfrOAmcouIYueUFT257
LOslLOYUckGCPIikvK1NH6Q84Td9Nyh6JdcTLZyXTdPP20Hm+C482YnZZcktU9caPnLzXIApX602
wiLleqnS97M6Egq2b3anW7BzyqyxrG2fJOj5qa3PnsWMETcmtXEIKdhcYudCQl7TD+yYzSuvMmqa
FjGlsUkmF6NB3s8s/a6chwLYvvopJ8v1EJxQJfQn30lDx0glkTxO/IZMZJ97frapYwG0IXiK8cxk
2Ob82seNHPlP0d2Ggjl/HAAA8Y4pdbuWZT4iHulA2PdbvwuwByqkbOM+lLdIX1Oo89OcAZ6IBww/
UT8yuxUZIrKn/HVBwF97acDv5ccsbC3k034zP7rI4g7aCcV7XZgLWVOHq7skTiqiRdjE8KoxEAjv
Q7f7mKZH/72OWx10p07vHHkpEieKZN/gQc2erCtE2BqDVSMQCgM9iXSVDdgMI5E1y/ac9mdACKHc
FclXc9PewqfzwRHidbsxVxt4c0tfyIJ3v9xksFQxX3pxRRNzXk+PNnYp9LyllLmFfYZGVduMUef4
Ow4fRD+Pg/AjjiY7+WrHZXNeCZB1wawjynMK/05Be6Y4rMAk/CYGq6avfmD787kMiuPe6lt4r3JC
lUSFyp27fVCorEt2ztJvDwkeHl5a8TCqpTff5SoEEIgaJ7M5Mcq5lnDDkH5AN97Mf5qZG/0mq+bb
BsLCfSXzQ86cOTK7A5MXkR/iUHQuINFASbTdNDWEmIFFYxv2E4kXJpdEmf4v46Dlg6T68JzYJbXB
9JROfBLGfroedq0L12Wnxuq3NbjQeSSaedqN0WyrVD10BCiLu+3QMiBBzj1VT6C1xf1OL44XTR5n
4EzFo8jHboydMq1e/gHHqTNlgWX3n2zlKrJnwweQUeuBccK734veZEKfm1vvBt0lwdp8tRKXtmdT
L46jlQDcGP3vs9fuBg5LDakGx3m1iBbwmCG1Djx7NJ+WMxtjFjSTK0kT1QdFm0TSCiYWOQoiAdM0
q8Dek0RW0O6dkpnKRZXf7v8WIAlX3bV3JKlj0DA+GXXR1hzW0IYD9fumQ/dGmb2+JQ7iZZApGUwf
7hZKfSBwRPdcZwMd2Q0NdN6NQv5ZeGMaDgzV53iLAMtLXMp8wjiiR1/6H6edPSYhIivkb45Sp3B5
Y7ibubDpp/ykrr4uEV9dlo2il1HVqVQ42fEJPhyYJvYvyp2JQeEOgjPxuhOj8LDKQduN7RWjRRwK
9PlZ3SCdk9SCXVRHkF6ulgc28PaIh7n/2qJaWIq45FTv2p1VUKZf/picMZytYKyjjuNfJp6ApZQx
1+ek1T+XzlPWN81W7fYJJA9377SMgeIKwL89ebYISaAuPC63NwM75L5cNwW1ZvxtGgmAeKJ2Ih7k
4EEUDYU5zo3kv/oAwAer2raVPmdh7sdEkV751ZzZLjKGv2g8j5JzaSemFwRQNkPFa8P/2ybgtv/s
7bCjsYny96KQ/Pj6oDwACjDx70p+8geWLUPcZ95nFBLrb1vaECMlPeU+iBX9+zopyqXNsZx6YvZd
1OJFgpjl/gQlEoFbC3Im3j7SUH7vhla+KHYcDCuJ7mKKh8g+QF69dPn85I2JeSKHLOobxhIa8cx1
+7H1bQCF0KQTE3RB4U4JU6PhBNXV6IF10n3T9z5RK6lISfYZq/crusI2QCOnLyUWYq4P6PLBvFDI
oixRVivWoWGAgASr3zcd9ge4C9Q7608iD/tqcmohXgO9aRCuLIz+N+8FtXQ9DticlYRa73CABL25
TWckA1PkGPAP+nQcVUaYJr6c9BcywwXVUSCeqxy4KBYAXC9nd0GaO9kgqdnD9y/DbAHvwpGgtFtP
V6x5JWOnaar3cS+rFmeSYm2CdGl4qxTS3p/dM8D89VCMBACZzu3fA3aXLh+fz0U48nMdhQqLWYG2
oJnxLdpwo7ZNkq31azumrnUwQbd3eWITTQw85xi1HRRtbLIa2BhWlRS29Izt3nw0tfqgxlnj6a/K
RlvA+XWJ8hsB1LFyvdYOzHfW5839gbZKAPP1GBy7rhG48vi8msL5RleJLIc+zGvEuN5U9j5fe9WZ
H51msdnQph91jOxblnUbwWV9shZlWeWBtKHNHD2YOv640r55mqDbcVXu7/e0sIKGuP3y5B5xoXc3
dIioxJLDP0DNlEeQ9s0cQVJk8mPyZwdZCJfFasgqPiwVehkd+yHifbt8+kRKAkIT3O69gfxsMtAP
q8bAzBPCKdw9TswfG+AfZb7N9mxYM785F4lHi5a6Ih4C/5dkNlI8wMoJJw0dNp5CMPBPhP7L07sN
N2B2bSyy92jTMAtAh/Q5d/E+aMRt62t6TcJC9+pUDJmdvSkfaWVijX1uWxF50r2hmllYFEQ1YVlv
d/SC0CvkzoOXlG2QLGfouZq2vQ/FlHKUz6LxlBx6dnliWFvBLj30ATFkI7d7RK2HsQLt7EwQCjJG
vJnj1GTXW49Els1bWq2XNOWj/nwuQEsGzsauBkNBgygUWD5h2HLPfE3y7eEqBVEGcC3RsOjIVLQD
bJlqTviYI3TiWBd/VzBOhaJLJpFOEL/olhckAPkAMQ2kLqf+IRzamCiZ/7nL7RkkVP3Xst3EGAy7
AOKMkx7A6982C0eCkoHWykVa3q2636eQHWgwbpLWnnOtItBcljfguY+NAuy+6KHs+b30i1Up1NMG
cZgKZ+BU2IoAUXJM1djA+68TBQ1BSv0Kw8huKeaHpaEjB9Ro708ahmxbrfg0mnFJ6GPjL+tmCfgU
fES7gaNjZZ/9BTc1O661XeCpertWj9/9c1kbRBJ9e4CnN7Hu+wS6exxH98ehM40NJ2Pn7PiE1PQx
mnDefK90zeWD+L/p/jiQ3DDtcTUi01bBN/+X+/LwSbJtBV9q1d+WItGZ7bxwNEM5hagqEcpAH4fm
MYP2w+SE2Qdu+SUzWzqDFTwPDzzIM7p6y6RrZEZxDDe0cosQeHYm4mVyt9uIu8E5o91bhQfv9Amw
C5oAiqfdfG56C1bKOBluvWJlS80HG4DJ6lVAgDmV0tXR3Fcl1m7/CQWdzhQCkgwB53gwvwBsOdQ2
vRq+IyEWWQlAAvpBUmL2/Mp6o9mPJWmYS25Vw6zdS93mKVIZ+/IiRkeq8v+Wi2QDEnckpBySKk6I
Y2lXUUQOpRWgKjl0NJ4pm8NH1wIyng9ycVNoFxmvQIVPfLvG81aYq7Jf9HrmFrjireHLz9bQxQRJ
OjEFTC2UiH+WXmUoCmSDjYGH8bO8QGbzbcAWRDZFrj4QMW/LGK9ld+iOCx9D+cmZgbI7uK9hQcsC
fHnxuYYUMOLL+ByMKpeTzMWfVrj5y4mtEStdhPIRM1vCGfyv0cZmVYrcGeuRvGjPr/I6RMP6PTTG
CI6bUq7LvNPPkkxvrvGjj7ZceN+J/2lX8PP2PKAM9d6nKjcTlV9ySMjP/tZQX3/EsfBzVMBJkTTE
ZlufkOQa0yB4lQZOUoo4FXo7gdLt5Amuim+xjZn24b0DiW/DlSwgi5oPzwhWjRy5Z3dLXAGh44iE
ViyXPn5vyfjNte7sVxzDRUZjjeMofqa1evATAOzujHcZV7i9Mc52UYsgRudZOrfJV2o+jkXHbAtp
y1VkcIiM22fJ1PnZhaSyyUugLdXQfJiRsvGFA/qFu8AlE7mMpnJZtr36TOYW32thH6JvVATGl9op
xMurEUl7zNifHu5K8x2t0qI8enal/jFLqvmNA7yLCY/UwoCrD1l8T5saiG/Oxm+rIEkeV9aGCZD6
rpDCnkcqEfLB7m90q66TEFsNGsu2M1WeiahH3Sxl/Ri7bDZjv5F8vGgiaoPlMz6UpfjcroKfAUVd
o0uHh9AFgBRMlWO4431tXCFkTwhptHSU2VA9NRm/Eh8gTCbRE+6WK/9n3MgQM+OSDRfXcC2ePAz4
/dMQ+47DeoTT0YfmQSOkaVw6Bje96h/iIixJKs5P8ztb95j/PLXdVbd2IydGfgaJ6rxxYGQvRuE3
cpn2isSgAqqP0EKsBrTYa1oAN1ycnHRvT/wKhfUrjCJG55Mm5VMYInGdvVfVkOCbX48X3McyBBIi
N214RHRnv9crXiwbswmZS0qaiaAuIkmfhvZN44fp88wX2E9a+142m8mJhzFRx9BCiDyHQfh/zXjY
lRX1sXaRwzx74wQcVptN8yw2cLkHdCKpCoQoqFLScXPGvqKnS8Y5cFeeWR13jvht9vyMAnJefNRX
PAf6tHTHbjQtYBGfozEIJLoeAujg1bJNU9Dk+aWGtaIkjsKC2/SudsEdiU2qFV8e9rF87qSBsJVh
cWKlx3WemNU5B1TCM9VHfWRzby5Emja1GrqnmbLg7e4WgJ0p9B0laApMWsBJdW/nuIddZnHLn66D
k2i2C0xoeF5r8TAxY92oY/1Ra4hxShtl7HVYI7/zpre99/NlUcAZz7qBPcfmVarDzHPy/GFIOeli
qrttdfSq8ZFDHizZZRTtFp7BcHU/5aEpOFutL58xTn6P/v6bemrNKikSw2lrjY/9KxzLxvMtEHpU
cQQvHwBDvq5lZQ/at7Ensomhp3fsgSKauHilECWnKNcZZDYq/VRf7dcD8SjC7EPdcDdVMHoPJPHE
NoSFPXsZMCfEDlyQ/rTZ/OLUierE9bZV7hagAXTz6Kv8wXTYGELzDJiDvq7ZVZtabHSbEpAJLYKj
x4lLPBU1Ip2jVrN/83oVLzgchrjrnLIV0/Ah969h00JkA+rXR6Gbku6CuOcMiRQhtqGhfpjs2LIZ
ChBm/kbNnC4ZsgIw2UsRtwU2gRyvKTnZQFwzTnLBaK+oszaQY7sfcexL51UZF/ZXEsAkvJGUWn6i
e9RC05lTJX9H5dcvh9V05cI4W9uESF77YNdzBI3ETeZHMLhyi6wF0sbQc/xMFnYqHmcwXhP1HI0B
ZekZZDYkHOvjoGS/PNn25bASNQLbSEvaZRXFkpA03VoZRbzJAeFDyA5gZTBeH/jF6T2u7NAb7LSd
CNByhsF1wod6ecTb/f6fZqRCPRme20hOarVENGW3TiaaXnjo7FZRgH9uY4r+fNpEBGMLNdEuDCTB
3gInFjOOGbTxtYvLEIKQaiNNeCwSllKKQRhLVnNtzNPjQPBAulCEHGeXlxJAyCrn34gy3fAonngN
gPG01robRSLTYH5JAKiWyyP4OPBLYvyEfgyt2tOgqVAcNCCMhDtz+7lSYnbn9pUtTgmxcb7S2hbX
gjduDb79BsFmzyKZZv1cIRuL69mcRtTrB7SjPenKACK0B3BzQt96bNrXyHZJWXzLT7Uj49aXRmlr
X34m4CSXlC0WDdhrSIt1R4cPzW+37B69VffwMqBrrBi3zhtgQyzTzEmNmtgoBc0bukXtDux4J53R
X1tHGr/DI+WmahbSP4XkA0nk0Bz/sMC6lDHbu30Wg2yXGCmupuSCZiOncOD/7APdd0mh90yJpeF/
zKg+8Xpx4QeI21e0JeGgv57LRcXOr3LfnBk6e3jPT6nrWi7dfx01OGiE39u00ZUPoQpSKefGHkkz
sxKQ3bIbM7+HYTnEiLXzxCweRUFXPTVjNu6TTdMkJpsuM1VrElPnPVHvjX40xSgaEtXtxxsQWKPo
LyLLyIw=
`protect end_protected

