

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZF7Gp+JQYN4x6Hvjz/p/glt8+Yhfw+y+NSJwSgFAT75FGfBEoCi9gxGC1aPKEYH1nKSH9HDVBmjN
jVYDQh69UA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bCrwACZO6VlyUjDp7F6NflPANkTfGVm4hgH/4AFvgK6LtR4U73r1HOWXfaKa3y3uaefm3opyWNhK
nV2TI2PpMLr9LswzFSOsgRzHCqR+XBS+8LwZ+lBVN3PhbED4ykAJBbHjWQapS4mEVXs8Bors5GDK
A5lW6VBcepABjdMHcOc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sWMXC7ertaTFiCso7MQnbVyuVSvzDQRw1zbA8jCBUoJcGFv+Da5uM/ZInIx2vKnorpctjF+RfQ/I
vLvHJ4hFA7ai3KLDBa+osiqXeR3vvyAO0dNGGmO7GQ1dYRUzzSKKrGTJhKWqDfnAsYaLroy6U3UI
uNSRIQtxv1ciGPzcMfrykPy27NH2CEGiCobfxP5HXDyrOVBqWAZuLaPzQRv0D8Ie2O70SiCDKawR
vbedGBup6qqgOpbOuoCX/zcbW+qJ2FxQY5Zrju+0WyLSf0XnZd4src68n6rXZlziL4eo4Q6lUGQv
gUEyqpp9Wiyw0QLmYTxtAKnwwMsfY/jCo5ZFSQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d4cZTzaonF13oHTIDZgb2oXxuKQXQmTrHOYXqYqbAU6BYAx+7y9fxq+NNlLqPYeukSU316ZJ2R63
uH6wrMfXFW1V94ov6Pl2EeLSPre3P4xtwdLCKbJrudZD4i07Cl6ICwNSN//h6MJD/kwUIU4k7zeP
ni9WJs+GmLVsVx0bOck=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W5Ic6b6KWpsR2htHXte3+6CjlmHZcuEa6WOajuu7k286E/JIlKxSU0tNrXH7rL8k7QTBc55tiAC2
sT6Jtn2FOqn9b4N96SwTUIbdNrh5Ew/7EjwCsd26VOwpEgD86kAwm7rEEtRCtStJR4p0yrbCQjf+
9+YuvQ3Ab1Y5fgtY5ijqZPgs+knlZZFAxm+NI7o8f97lEMTpHDonVgfj/KtK8xhV46JSrDB2FPhp
PMezRFDPcrnrGio0JnUe1oPbSneaSJZPAFIoGiaaxfjjDJIOa0DMtbVjecaL42P3+sAmOk0R5Mfk
8MlmwedAmXWwr0D9NdqrNJ68Zt9aVa7CXXiS/Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7632)
`protect data_block
Ec/bOertbDn731xvlelQPeSphY2LEkq/GEKfRNFjvuazoWnGbypvDWYXnI3d3IMD2DCEp2vKW2js
qcb031ouwTiKJYr77fRey/i3tWWLUo6mSmuhWO5MEviYhQku61MbneSG6vHXx8FQ36Y9HugZN5XU
gn1C0Ys11Xqh5pUeH9wRu2KjVxwCOXCzy33zx9qxW4+vljCiqfDoKvcukSTg7M5lCTCru+9/f93V
EvYgoVa9AIO/TRkZg2fvjtQHc+cFPasjwM4tGaBSN93d3UMy/y+cIt8ZC6PCGuTvTL5oLlkSgqct
4TZ/YEyGHK31WY8RcrLJE6xFYy/si8EJhO6Vg5b40dHajXoMTiu2PzQ9lay47d/1xZ/+eGi2Cxn+
a7b73EUPKjx0mVsGg/DAsK0XCsX3cZQ2kaVTBPzhjDUzduX0p4w9f0jDg2WpR6mggnNVMrS38AnY
Dn7w9XaMJhoPay9m8ILmZi4vqOdfE2i+lGmXrvD9XbCZthqi8qxUKnaRYqjcHb+rZN/swuRA+te/
X7pztQVOLK4wG8Alv+HmczK0XM7R8ilHwdtFOxzIZaE2rKduP6ndRpsDKv6Q4hILi+jbRO1/2LQz
7bXpaSrMUXRgjOxa7clZaHSAkclkJ5AyQ1BrPeZ94U/87i7kxvZyyRKc7RSWP31owew9B7+RPlLa
M4E/mPo3mirs8L7fjKoZYKH2yNQnHuhgXZjNYdwVE4iahIofrCsG7y28OV+69+FXQDIS12bQvqrC
2EKPVVlcg4m7kzMsV2uv4YG4wxMPlO4T+YoY9LYNd05EMyGlj0/un1GnE7NEfByVoNiKTxy41+CO
XbJN+dlTPNzd6pOb8143jJSOctDePr6JxcN4MTnbDvxLWXIH5oMooWOZRf+NDhQ8gk7y0kr6X16S
zHAyazh1j2t5GZ+EtzRarVDYffzUMurN+cg+vmU0+Rb4eluz+5OtaTAU3VgOLOTxU8aeGq5HTVaH
ZWa7nUc2cogwySC8mYGlegh7aCV6de1JY8uAf/v+eTRoA1j7HVUGKBr/gXIGobab3YFF7kVpyLZ6
oSylc2NMa9xu+DSPDO8iZ3Z887a+7YBpaFdD78FP2hhqEd82rpDRwqvDuwJ7hSMGQ+lr7xmIIYII
SRIE/jkVzaOEdEbPUb9QrzfWTeMEidFTltTpYZL33fGsImaw95KxnM9shsmSK9gvWu+/auuM36Vx
MRGo02FH8MEFAFOgt36ux4F6Jt5pR0nK7j6OIjI072z1ZKNX8BCFtmb3LyMH39vQH+7+o6DJu12X
Nj4+R37hxlLbNyFCZKyM6mMjlHCbbgqhApXhmikYu+HqizB8pG5Cvz8VdfUuBnztzoXZi7IdXdhT
3Pg8+74n+vfT0gTZmFPhYXokbQn1Q/Z4RSaf1GTJZ8OdJEc7vTddX8/z6JE0d2eVaAYCdrP6gmAB
ovv7ThC/z+77KU8lIBGlYh7o1VRkjUWrgo6qnG99dhl5puG9sb+bI+rlEeRGHljswcvn+GfiIuNx
6sQBAh6uSVebNwCzdt3DksY0DGOI2Ez4YOaFM7aGLzfi0F5kFR3kP7gipRRYP7rVc0jlfDJbZBbJ
uhgsOK6ANDAQRGfJxew+Fn5BUrK2DhQFN0oee5dLXMF5adAd08/zvSQwyxDhL6tZ2O0OOIDp7u4o
WTy4SzF4gV3duvFRiC6ZDAWT0wvGj+QUsNGo/gWWZGxufYxYCplr4DppkrA0PJwaGhdNOdh89z6p
8RDA+Zp/+PV9+RR5+VOaAWegMeFHox+l/vc4VzHFEqhgM13KG5rWP3NfC3Rajpi3ExOyiIYwehe8
K2ZCxmb1TILYYxDQKhkYyJ8hosYsYegVO+GTRfhHQF5koxJ9hX+/aduae9PrgA0D0AL8A2o6tH8f
fEJukEY7S9pf4pUNVQPMHNfkc0P4I36wL4xB1XRG3+je+XarGFFC4H3SoMatb/fpomm7tZ5nHUrJ
IJP4gB1czq7xx2hNBl22aTxmBrFPkOGJkxJN6yqACeZ8EDoxKMRpCR2+9WPlOg6+/OA1M/6IFD8X
LdeeLMntDeBuLeP6oGcg7NSODTZLuxthpsu9HhmqTJ88/F4+/3ehdKvVCCxrY4hK7QV6D1LLAgxs
3NdoRQaZqfsIPVQIHRGUZztTUpCVs3FqHtoXYgsoK1m6JFuaPeKprnh5z5LsxwRZYRYoBjs3ZI1h
j9Rjd0UppwbliCR2poffUXMC4sDrX3a8ad0rNFCv07ZedE3wRaaJSCbD9ByAkVGhQVPQd2sFcDON
BqRB7B11I8OQF5V8i7ddg53NBZIUvopFmFloT1WiRqN6F6stkcK0DzUs0N9ddrmPA9WJFsDWmYuc
jPBCIVAnjO+faHtGHj52S8zPC7IVwf7UeR3Rb08/Iu5J8S7Vu1AMT1PjBGSnEMguIVH0IIjbUpXh
IxWPibAFtuv2bFQPtBAi+09e7joT1RMJJ8l5kdMY6xeJEgLOewW1QvndegMgxEizPltXkZYVyfql
PLuVmPrygv00zNAr9EXvLZgDoMnEWuvqK6RN+UgowQ0aqdK1rdMJh11lGcp1PodeAL5+YohzyCb/
F1ZUCxNyp+nYc74RlbIjb5Uu17b4t+X4TTpnWfN9vstOPmUAF5SoFAWoUhlOShHLhJZIilAqp6hV
5jw5Zurjn7X40HYsuVHnw0LjrEqz/BooSPLNFMuioWnmXd+WbEOTH0NflJMrNa9n1ouxvd700VpO
uWyklh+mIaRvDxzvqHbHfIkFd8Zxiae/RQkCP6jxjjiD2r3DJeuuWFtxCZ0mLJuuM61fZ/r0fQln
8Mh1of0oMYjm7OxJzYl52oFXAvgrjceumRZbKSWHVxF3H++qMtkNYVDv17us0U97eNsxM+WPnvDm
1zlFjBedHJDB8eT5Ws/bz3TulGgUQlOBwrjWeN5VxeDBlKXymmIDozQKY/PArWl0AteKFWKcY3nT
WfFVLdMWynhnD9e0cg7gzigEeIfI7AH18jdb6QRDH0PKRIhdpoHtegdoSg2th23Kqs5H91Hhj2Kg
Dtq2kyrdtEPziJkMUwa117YVBh/co6ngPNlBsI1bQAE1xJxi6vnZmFVW3yIXV2T5NiNcwIhd21Zd
T/qlkiZNjpvGCXjkLl84HdOinZzCIaLE/d0wncOWf5a0UlXlKJOapnUTT0X4rHxascapJE7dL6XY
ek8yQnMbAI2PemDy+JFdhsMzP6xHwL6HrzXSEcZrGd/1FMeFu3wBDQ0wRUbsBy1HYTXJoBaBlcWy
Kh0PU8KIvMLsl2NE9zNfZ53W8iEe6kIfIqkmUYOoNh3ty1osLzSunZknN8jqRrdAEV26vUPEKjOL
4FeLr2k2BEOJ1AdXyzqUixev0dAUtVBuoPThndnb4BwZugma9Pm/6VcYkGiHfHdyghxO079TKi1I
0bchfvCKHbK27L2iD0rxBI3cJO+MQoBc0CGDbptRnIViZAKV0zJ66scXKecc0DcNnt5X4ltRvmpT
uPUM2ESJ7zNgb6i5VJDfXOvE+SGCFynEDBIGXxZfBZ0eVBazqPb4bcZmSA3doHZ8IrO9ZgBtUqfQ
RJlp7GiEOecMOku71PThV+2c5fjpIeOkMO9TACEpI2g0wJKV7fg9t98nMJ/gZd6bZmkwL+G4maZ0
knsb+zCa1j8PEdYG87zrUOozqlQcqll4agQx+0JtcwEH5PKwwoK3cn2Pk/poXloT7lTNrm/lFY8W
bvSF6TU5ZkBIsF308uwmgNOn/nEnWhjI9IxV6QflzdQB5rcwRY6DhP68+PrwD5J2TGIkIBsg5j9N
ju33FDacChYZLdzc0zMa02hutohX0rDobGRXTXw0WdqoVv/DalN5dKI83hTKQ1Ygla1fG2VosVEP
DQR9Y7iwNXDz/HEnrOJNpDg11ID1lWvxNgOF2GH3o8+JRrhBpJXx34IAxnEel0cUguK1ZfFgzpFo
G4gKg/5R3UFo78Su7nH31stp78m4+pCe5iDyshfgtMq1v5IoGUzWu8ZFswyKzTMB66LzOhtI1II/
+aZHr0K0ye3xn9ZWLdyH3p5nDPULKM8UJXCokK/PCPGAIfsvafatIC2RvzcrCTe6wuevWc/5oZcl
xUWys9UOCbSFQTaKyW0Wx9TEbQ82BvCGIc2Kfd6v2KdWhYm0vYxCkyRWx+pmCJbZnouTd5y6oG9T
J0ucGpiZkY+NmRCHin0ystDs99cTt3yyH3LfYY+0n8tFRballT4eD8T7M3dTlVgpB9tk4f0qTG0o
ZxSRwcYHFDusbUzQVbR3TrsvRpvorUqYCf1EYbRjZ+ZOg6Em/Jh/DbiE1uos5OcpHxtKDWgDTwto
r6u208dJ7md98jMwmpP3wopt2e8v3SLKc8kXFsr63sL52as/SLCJoF7JtvOKAc4tStjITW9mhV62
aQmed8eNesLtRBd0lUr/LEZEX60gVaG0du1/mwVaOgrvLpBg/+l5o6tGnYGGjwRqnGJjSe12yOBS
3mdMd57nXjydd+iElS14ekcYsgGJjSZA2LPWJvs8wlXWMx5ZCtyZ+Nh0sXymtqWMXfpWvZDJbwI5
4le5mRKercvFNkSGKueLgCPxkGuEB8AN2+spZ0y3zu6iCKEmyLezunEHGQ+RKvIvAYwLWGBMZTfF
WNX/7egwuwLnEXJZllC+SMx5mtL7Z9p+6MS6gmyRuGYTQ/Tj91juDWlsUmSIzpTmdsN84GZzl4Dp
D0/wAK+HAL5HmRD+nMROYKQZqQaj4BNPIQ7DvJMnKYndCaJIj69PEN3WYfWkoZ9R/MvN2BpgrCAU
TpNx9mkit4VvUn78J8IGIvGvS+IDZ30c8UNs7B1HYpUFtGEcihJXn/PsmSCpdo2lRwePUjX1Qz4j
uSrEf4a1oOxWJfDDg/SQSQ852cJTiXqgxv0PpkHPEIjYz7BsdqWKqTArfflNlTkrjJ81OBKfb86+
aMhfYA4UD/Dp0/3Kn1YVX8GpVoCOIiOqu3oYu/KYe7tbyLFHB9hcYrVHs/j8bxHWoRrYD3BlE02t
wbpvcQGc5+5M8oHafAU2k7xvqWkvRKm1n1xiwHqaWkIl1oJ14rSXk6iCTK1hjvf/tad3K07umG51
tlaRKc0lzIHK0Zjqq6P57Goo+r94+3YHPc3eBVTYYCVTD47Ld/i+1Xz1T7mUdP+IBPznJ9XZmbZ9
kHppuORqBVX4XmxmiIcacn3LTsBH3FxQq7kJQ3Wzh3N4WojLbWvRmkni1FphuWILZh/p8EHGw7Ib
XosQtbqwwyUTNUHZZMR4um8ceAH74VB8eDL3TbPnvGkHIpYVkySw9gUDP/IbqO0EyY3TTv9Sqh7J
CM5d7mnrV/vZ1EyNiLPzKPEJ0cE3ROqOgFTVzrkgR62yaUpzCDzS6vVA9rF9txxjfdVAprprheXh
hAir4CfKOG27dq9zIK2jVCpmHQFX9Vu1QvwiwM4LUjY+3cd6MkRKCU3fQUguHOx7IS1jiFs6/bU7
URY/oG6xO+6x9qXLx67975yf7zaEBpS9OWxqvrBl9+v7pDLWbozIwmaBH5w8e/vamM9spg2GYX4Z
9+5fi9BBbH65sJd5Q7mwW8TuazCUYofEfBG4cnta6ptl+TPaTowEiXkiEFAAQtxUUPY/N3oXwgcs
aC6GLYXMJ6Kh60BHXMh2ZJ1xYok89014D4QYoctRNLwapdWPcKdq+s0d7UH6szMblj+NuG7En31r
vvjiThkZoVsVWeDPDRVFhLiV5rSz1pUXi0ggIqNEsokh/ta4PgCbSSosM+piFOxqAFSceRlblrqj
6niPvqmsibmrC0dMtxcwOwH2nj3KhLHx+LK4K+oOibwX7p1pbZdYZX63PXcEPkZ2kFG07sWKlNyP
MCDOKcs0KjgG0C8224i0rmrhYPFDNnoMbZAE1kcKrZrPAwb7qW95RGrO8Ib7W22E7z8oW4vj/uq6
0O4tj9/BBgyGtzd2S6mDWtWPo/zBsjfulpwYmTp60YJCuSlgTsLAkN8FryDtzKtQRp9pKkSS3Frd
srpB2/HUWQRlAPLo3mmHc/LsbA5t6B0VaaHDVClnigkbtEuvw31CHw4FfEsg59Zd3Awunn2Rvo6J
wVX6l+NTVsRzteTTketvDDB6ztIXJNYFLaM1pVclnE7nAFF4A+0mZmWiQwD14s7ChZ5uA0PR91yZ
gEKflRFZfBCqxqNEemC8X1aQAIyz2I6uBWORri+oyKT/G9s5QQiJpYlqTyx6Jzj/jj6eZnLeS+zP
jrsE+M4EHjzYOBr9GAc6mRzH2GUyi8OW/7jSPgonbABkk0Cu/Dzx03u2AoFsCKPq6otawnbKeijG
gK529DpTvXHRl/U9TvOmC2IDnPsCY/rBZrMD+q0BDmangJONZZ5vmn2XldNgzFE2aAxB/8aPDYLI
EF7ckG+e7gQ2slsR0uDfcBZJEsmCSVqjLqG/leLdTKbZPgQWIgS/Jufe2QXIKMXYDB6vzwE35DMo
Rf5bWu4Ta1cxL8aAOcoRE1iC25/RESX1hWnVewSOPwJkl+iAbr0c6xs1t/PXGq99LtEI9EkuRjjS
B46OKLdVKBbjXlrzgLuyyWUO+n0+rb2Iuv2ACz0LShwcVvIkVB4Ys+TkjH6WPYg2C3MWJxnqZTCC
54l4jO3nDxppKLetwn3AZFfKoa1fOdaR/4O3+75bkge1eYjTEERDAsMZAV6+y0NQC/eCyKXFnV9C
1x0r+WrnY6vM56F3H/q4M6+MSgzuz+uSySpj6aOcn8fNQvwlHkGD/HuyysD3FmQkSx7kgqqEYSho
TrdZM8slLYgdZWn/dV7MhvV1h8gi+IV9WdEGUmhWjcBGsJ7zAQIB2ZW7l0esfsMNZ1itWwtmr6Qz
Dry15tOcFuCrnPPuvm4MqS+z3HGydgPg7bJj1bfGOMRhZMDSPlEOmZuqP+QU18T++8V0mJq1k5ZC
An72Svip1FisI1JtRk1BiY805qRfEmev5iFP5NpjGwxg+oJNCHYQa0Fo3gdH4zLXQY1un5xDMm67
isVpulTzNPLN57C/tF+ERKcy1kf3dBymbgPYzvoEcMVAdaVAyE6Io536ul2olECm65MEz0Szd9sd
oOs0PDJKOHc3xuW50nraPcxatzXhGZHRf8QZfrP+VDhakzuXe1ufsxs6Z6nA8WUpXl7PPd8GKhGd
oz1KXsmHlwcjVqMIHJJp7YJ7llGyi34qoeGgUE+eelthrHTJUH5VsM8AmoEdad8VehYZYhKZ9FDF
QbfdjL/jz/pXRE86d0mS3v79mCVspWzS6gQvhWg5Hy0k+0+eNpGswj9zDVVNQ9us/kIuiP5471tF
tIYI89wCdrHZQZ4e1OKPUc4+Nq8D9Lw/3nvLpZwDq6MrYRX4tz2ncyaRkAzYJrRiaf/CDZT84jGC
PGpqpihDkBn4nMmsqj3a9FDfsLW2FX345Vyagqub1ndfiIPAzQSA2zXJ2S/kgUb9m96xDr7JSQ8b
sqp/vYTMaL5mfBpYx2aiFfBxYZAfM02ImG9zlsdWZg67lOGOr62wZ+e2o8eZ/PRkUvORLPb4wHqn
vlm2c2rSoDZPUMaUQO0nnKvVrkoVW+fWU3iZfz/olKwwNLiJNGLHxuMBCACsDaoseq8hCm+yb5QZ
IRcLdQcOXWc5XpQGj2AvNOmgTni7GJDiFtBk7e6wL/th6IJF/Ww4EBd/Pip4r1EqqNF71Imwt7Vj
wsUPBuXFy6BVb+ocXPVPAMCBNG8MHMu89sHP+mUkKTWYlcdwnrhONvSICzPNyfqdVS2IcEJs24QN
CCF/XT5BtDTezez7vds4fairKqhb+bC6mA3B9KSHRIu1c7xOYq1sNDLrDuLAal7FEkmMXwGxJwEU
y9lB0uqpg0e72IXxvseA6LZZ6gEJWmpAafkMLUSKkQnY705+JZ0HXfL9Bf5UUh0oshD9p70351GD
nHwKw0a8tJOtBOTjEO3WB/q8Ba6ptZ7Wv1zWNRStY+Ch3I6WOCQ7Ffjp9lRGTxQX550Uay7g9eJA
Mx7T4ngAO6ksatLhzdxUlo1y/Myq9lskp2OUBOky61LNkAW2S+HZsLLf1Tgs4TLnx+/qTkC2tnmD
iX5rKGOIddTn7R8wEg8YKySMmn74+WzAo0e7BLy+hBo4yLdugEAG9D/O8C5Eg7w72EFEtP2PTdAt
3pQJcJct5KfhMNV9QOJV6CsEOzktZe4febmxKzOyQy+jmtGYVuJlwXV1TUCUOudFq6sVpX0+adqm
rTMZwbAikl9X4cLzAb41U8MCmI5oL8as/SqBGmNiy2uC/acPV5X4zZGcL6rzv5QEAvR+l9N9S1Up
8iCmvZLfRkhjrauHtYwj03hKR8zHy7W8iGBTMwmyfnvjHE7DG3NbWAEUey+Nw/TsuGEY/Ga+QdUR
vzG0AnV/K+rajugcGIrSpIaReEK5kCCBxlIG/v2iUJRMKVyTJmOLon3KP0RlLsnFBZVwYcK+LceY
I9JUXI/OCaRFK5JfbsgUHsGcbc3LVb1NcKdEwFG/ZaAHlinF4F89zFZug4cXpHvKqBcai1qdjoPh
SW/w7Pj3M5RxJxBehPPsUJlg1+/PUt45hePPRTHtASh5XheJHcmfziv7WNQm7AeKPYMmyC9PCO69
POrd6CN+cjN9XmW/EWQ1BHkaYkqVnRco10KmQqARmOrAUfx0MVWkZBuM3sYvA0TUzki0Lh0rIvpo
baGOCZS3dTBSpVAgJFojDdj/SJ6YIHRESNlJnw+8YvDwlY/z5JkCPZKBOoZmxirTlsMEUCakSHrk
qM/q9rDQFLZ67YE7GdYUYKOseMpT3gE3Vr17SiJnMX+Z8kQgeyGVRTGVM0FCHrDXMdyfd3RbU0KH
fZm/5KzjCDWtq0GLYaOycXyUtkUioBEiAJ8eW9h7ag1Ihqtj9FRUUll6ZOYB8jDU48C/ncTYDxeH
yQGL/mF3Jx0vUQ+3GQyVevJwGvXphU6knamjl47o1Pivuj/d3YlYT7LaMwDhAenf4YpnOKJXIMvS
R8ZJT7UXUeB4ofb5OQwXVuHG6H7Wz4SR4vlbNNwaotefI6nfQHza8tOKlEVLRJfQEhjZ6bNNR7zt
fuk19xBBjknHM2A1b2XSxZVFG9ZDWmDH5kLkx9J9Xmi4YOk2VRApu+LhkjfdRd5pYKxYB6Ycdad+
nthFjahAVCHLXt+6jKpq54t1BNLjc9GIpkeIA6ekcSQVc3uoQeZk22bCfhiC2nzrdIenV3cs3t3H
W83Ve7Z3tnZtYDtW9sZQu5fcp3cImoKd1+TtQfgc7HFHoT0veoyCxzwQZ2FzIkewriZiG3oXrF8X
ZeI/VnPp0mPQQOJImG/5DhQVu4tz72VOW14jhsRJ/LMkJgS96hPS69d2GWd1mFuoRZ781E6m+ySF
mrirO8BUTSpbEnItNoGA/mH8m21wd7pipAN9T7XZzUWa5sIwUXFVyXT41N1imur6mInIbme7R0Zl
QJlrvxJDj3kx0TM7yeBWQyIu7ekji68C9e+l+MtlvD/gcrmas7FzLOi8MLqlEk3y4m6tt1SR/5zY
zg9wcYrcSOiERllOWyzz5V4RwLcNETjtRnYevo7wrh+KvrWVG0lPj/CY/WoQAXyRMsjA8WJkjQJl
Sl0zke4ileYACwG2e9OKD8Wirk/9HZV/XxuAYU/+dPK0dv/t+9GQDuT6pXXiBwfzTHjV5203JQlE
YfUa+3ed00LX+0om4dy43PZEiyYTgfVopYONFmXZGnQsDDC6AlyooRZZwOLWmonrxNH9dVTRwXYZ
Jh350QltzV4tzIMGogqOv30A5YahyZhfqNT8EwU4pkPJNeelMFrsrdGR95478kcQNE74tKCPUdT1
Eg9VUvX1OYT426OXf5GToyArkECS1qmZjXqpSrlrw6YKR03VR42YJ0E6ga5losx2bxOVyone8NqB
00ZJHqOmdILnXR+AorK8tc26wgWPV0FPyw2nzw55EnNko6QSihc6vkSAbVlIPY+4zI/EliZGDxA+
xFyxSG2DvxAF8QhA4nFnPp4LwUox3dv3qBznhQ0Apn3jbO19NOMVnAxoqDoEGcyV87S06riW2aNO
Wafi9X+bIh9/KzF91azKD6UtRfGJ80m275GaXSGl5fhlIiyhFe4FQOpWsLTxKsbpIUYjmEzhR3JU
Tjc/eSJZduGRxwZe4uuzG5JwMRd/oSbtFpe0gr7mnWMok4u21szjAd+6g7kaplgazY6F
`protect end_protected

