

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QA13xX+R/ACi8km79qumYiCoL95/JTNXmw/Mv/Sollu1nSewLnwk6qQvytLuy2zqP8g5ZHUfDkXy
dYJVTyRzKA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nii8tC6PWRY1wcl+Yj+dJQmorGaa82N6txtyUcQdtmyxn18ohe6n/SpcWdMXBCN1HiV+XVlZhDEw
KvXEmx5H6nBr5/f6eVRIc3k7vZjXpluRFM7lDsLgIpfE0fW00UnX/0rMYgmxn+5+4dG7smGpX72S
zm4Z5q7tYiBa+z76ex0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yppU6wpcO6vEUEaOZTTT6jS7XbaY+e5Jeh6nknICBRlkmT5DzQmd7eWK0ShMWSlNt0Fv0kuxSdt3
PRQVKoJayZoHlh1UH0U//6ySDV8PrR8ZKYbnb5G7lC3+6hAsVS0WEHoXFsxe3QTXWezPX8OXISSE
YYTVzXqeBUtBDqueK1cvQyMM7IWnXgyQ/0dRh7UmnEpiOonlQALl1eEnWSxVZ0L5cd+jDbcSlWqj
VgoBh9A+IbjGjOjE8FOaFLUMzvKXmpjNiGzhwyN1qXczrRlE54AWkRUECVVEGR4zuEA7VTQH6H/B
e1HQhNsFNtK03nDJRyhoiacaeHGOBo4yneyZRQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xoEHrB3Q0Yfcf3MYYTBHkrbmS0WN00JVFDeAhGuvxPP5kv5812Q+oIM0e+z8RwGLEwQ4F0j3UPw9
LR04YDkbyd4XfjRJQED6GhUyhlVHkeZ0vYn6D/hB6y5zA45LPFz5aqbLudigfR6lDZgyof50XSaT
wkqaJ1dNbsbYXDGYiiI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SZoZou8zrLQYkyuoYxGz7q7TKCLXDf41gJHR/eNOYbjhVAUcJLojwHpmGq29Knnj056DtiEpAnUR
HkNwqIIUQ/PzBp2ZRgLcYUhgAGFauW9u5fA3Qe79SJmVAKU55R6eP+5h6YaMx1oo7Myp8ZHgv9LK
0atkww+rNUFhc/kS4ivaypKADJgY/Slv1X55We59ldg5OMI3+jFcKD4Ow4Gbs5tHnIUzKQ507yjR
1wg0oIoTMEm7GhN3wZnee1A7XeomsW7IrTE+3/M1cRWhdrj0rq5nqrI9yilbmzqQyqntfJK6N8Y0
QQNZFJ8oCjr3X+2kFBb+Pd3/scpZe1PtOU8TgQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20896)
`protect data_block
L/+ND0YcHmYknVxpg4dM457RF/TW6j/2EQEimVW/Usr7lZg7si8cxwHc6Wh6MX/Cakj39GkZ1GK8
WmVvNvza0VpHwE4cdCoDWmKEMt8nQglbiq6rqtJTQd/xrBbSBr8CISLo01OCDOhmu9euu/iASBWu
WB20kXiXB0Tf1pXe2S5ObG0EVC5/rdGLu2CfvW0DkrqGF/DMsY/Dc/e8QvhHC3oiAqRpYLkLUDPu
rAri7aGAdQnK+bxsGJ4TK2Elk8rGOdO3PgE9HMqR6VVTvD7U/eE1L2acQ8SwtO6UwXwEPaDPd5B+
hbgjrxQWap4efmeuIZrVS/+0v8pUyAOplgwSLUtd6/YJO+K9MNNIm1cQfV0pvVoUKF/vsF92pLWg
mPjGwiGmQFS66Z6ZhOTh9GXYX4YMmFAc2ainCr5TF/RuhvbT1CnFoGhJ+mCJoZhzc8H2hQRas+oE
J5MLKcjII/s8I5PjTFkv3aECyzuxBaisCEPCO3Z6mmTgas5dWRbLBQoboojR64WqJ9md0tTFxfJv
jFAGoUFd6i8f1LdycfL1+nRtsByRroMlO5lrUbi2bGxR/8QBZR1lCi8iYQmun0+indshEssj+yYH
7vm0SB1ONAms/YMsh1q9Ab8RUJpik1WVdqEDHcwg7zjP1VjFPEj6aFVK0P/p3j6qJW2vORBnWIvY
d0i8fw/PUUoY+pO3XPe5hyigRMXJacntrBXNrDXsxZy/QmLXFEqzoGjMuixwmrPu9uSeKtIn5fk+
AiLU6Lomfphr/PFqeDGJNo4HpOfeovfSlP/F0mEyR6h4254Kp1WzLBNptxufrH2+Ya7VN/IQR/dU
vqToP/64e3WbOtpZuw2bB1s3ckBskfvO9x7pY8Zbk3/Rfcp3s8udS5jxMhSaed4YKuHBvbuVN4Q0
BnwfznNTq9Ln+jj6XYv9Tun45OtJz/Zhase0XOy4fU7temJl9L0HzCteWj+IQJiKPzpxleweoTL6
1S2rVKena6ddkvYG+0fsHVIwGQlOQPM1PVixCk++Xzaw1PKYhOLGoLCciUpUoFo9p+yEJcPXFujc
g/1i6DAGawiyYo8zc4aR57O+eKWV9vJYUlBehPjXquMMK2AojEH0BJGwxd3EuA2q+nmqexP0ez02
dNZ+uce4PrNzXDsfLWmQYXDK5of2VrybYL3FojEaqzh0FEwGIWN9l6FYkxV/0TlPX7XwNjZPcH/r
Aei7nuXoYLqzPpq2yYlgJBLMaK0LXrPHQQeoL1ZejLaxbheoDkwyxmPTTDa4fp1lYw/gB6KO7GN/
lopJmQ/QNelMK+3GABU4E0b0cB1iFhwiDdHWa/N3K/9kUpjf683elkCgWdxI94FrHzkpZwIOzmek
Cwuc0GOnn85gVptxrV2qq5ov5oGIjxnLwS6O4RPpx8QfX5iYk4b7BQyQqT06VFdOJc8K+rnxzQIT
BnDJWS2VZEMNARMPpACfVxAILQmrs/F0AAaoXeijbwNSq2jx/glLk6mtShRqSLNBL/zkV2yxosVj
YrdPIPsHwDsKNQEoct+FOISxHO4yWU2sAeM29C5Azqu3veEoKiA0VUhyzQEhKBovcONvsGb1/f/C
SJTqcwQmYw/Nti/+OOp9gleLWjjoVJUMFqCrS3iX4V1940Mr6HR2Lhb8spTu5yvvewwiYRC35e/i
ymn/oVXotbogMsBbDr8s9xorG51vBHmtGTIDco6x68QK9A2c7Gk3kmuYvU8mmCLFmhoCgAtiZ5XX
aWyJ0uAZD2rpZ9EYkSuKf57YuR/5msisoCBwKU4ciSfmXAUlup7bJVGRAZLDlOop2TM/Tb2vHjTI
rJxQ9kgOUHgvvm0BK+SHzGjkcXcy+MEgPAEyvwzPLYpZIMJTIHvjD383lPgYrTYKjtpq9s2y/AnG
yBq7k4AOGW2Bd9DnlgCK3vIccV98NxTYRwzpK3VRaJTNUxeRsecgMCc3J5UtnOaTPhA/KzOAvbii
nEPor1qySzoG/j2MfFPHAlYjn4oiIgPcNqPfHERyTa+ln98+836WiQM9pafMytXceJUQGBOpU3Uv
reHGfXEi6Ni3NZJEJiHxASM5lygJdc7AZ0GQk1Q0RvVxFw1yHr+Zk2oqO8vsO0MVVG5JY7IoNx9P
/yaI1jDSK2GrkhynMlwTR85U01zc2KzOlPgkJY6njNSi+XK5D863NJeqgUTT8MaLSj9aJcNrM9f2
U+Z8dqQR2/e0xWpDIliHc4c9wgq+1t06fXOEtsVm3cnlBpG5LIshQ1uqdvDqzbiwVROE5TDRM/ye
TxshQFgjPPTB34NpmgXeIm+YzPk0zK9ELVYeV1IuczKq5NDd9gOIAZeVDTeFy8w6HJtY2tf7cSin
MIkuhykdortda9M6ktyUnw/5p36+bfaUatJvmmINICGlXXFYFiPMm1SSEulgVq5vXnQXrH60SoeD
AdzGyh/aH+pCKyvJxK3XT+1mq1oOHG6LMygtPH6bfoL28VmjicSYgz109WTD3LkQMkd0dSVc/4vh
3bBo+pWWyzDuSWzk+ibiFVxBju7x6deAK/ZHJxGG7xZbSm+KSyPS7FSP41GeLde8gaVUwpYZ9Mjs
gMDLLUP5If2UItmkSmME3m/l/7eHJBunycn1pnPNWpQSkYf1tQWbj+3SYtTWRJ4o4upl/nhsGf3B
jr2dSxRXhU54XrReTKcSwCOoxuPrgdbYws4ovfjztefYxL9tYZoBBeJ4/6nZQkUfVkKZSs+kyfcX
22kxJkQRMKrDOF+Q8IFTFXlBmSw+tZO41L1buMGVHIXwwTXCDigTVCGnDqucPzFz+vVRplrDTJog
x2xJrGYLKdvRzVscHA+f5yNTlRfaGFns9U069xXa+W4ese5zy5rQY09CF/hu0s6XK2kFnGwDGEtm
wNBdp3qZTHvBtQz4ZDHe97/U4PotnM7hRAv0LtQ2qrXiYAMnY/og6Vrp8O1JU8+SRFmS0KXeSRVS
gLiSq/FbTa0n9Vt7V41RWwX2koOGcNDZCgZ3tZV2p2dYmD9P1xK3pYoce2T3sSJPA0URKieVaJks
PiY5X+pspa+p1I2Vf3ZqRimc5Asd66KJczAYHlVu+HZfu5Y6Exwne4tgMxhRbrCj5GPJJuLV2Hwv
TlghylrK5iE/eiIMhpIbT+y8rGR31o7SfieqH1y6kb60B5WjCmqm2/zEAm0DdK5xgHIwfJ40lU1M
P4F1kl+2G9KB4dA0zQGU1cjZoMxMupNbXzOujsopBZqkNS8xtT2okNipWWCsajbxF/pWakTH6Gy/
DA6cbHrf4kdzJsisaB1vHLqG1VojPinPRb80Z/n9h0jDHo8xwwFFmVht0bC3+12tCPhSZ2XLLzsj
8b/Zd1khkQ2nchMlBXtYWk7uKv6LYGa+q2HTnEZjKrT6q8bluDkjc/IEf4waBtOQ+23DpW/cvrJJ
hjJH2K0Cra1b75IvzM8g0aKBRBteupnCEiFRYV1MvB21aCyv503XGiCaqrEtDMVSuilN0aG27Dam
U6YIAbHlqz6DzwAyuTcbpyFKiQq8dU/q0sI5b0dci+xEGOMkRUjYKor8J5hAdAemwJWYbF86zCyc
eveNRUaenpdB6JMgZUaI5LSWnkYB2ki2EhWU3BHZJ2qbx0wUcM5NQOxVQxI7rYbeJjhZjOgDL/y9
Fr5Omv35tcdTEzp3zPdkINVK6go4DoWCsxk7EnfNAk/Uq82D8Hs5m9aN6aHcVNlKQbhlk3d/jjkM
KW8M1QMD+xJ7zIyqtB9+tcgQ2ADHxz5612FtA+HTnFyJ6m39s6ztK2BtSr5NCnzB4lWEXBpVsgF7
kUQLHhrjT2PF+PZg+oqIsRsujQH5NrXZFQ8USMGqXBx8UxXSyPp7W3JQRha7cjLgQoGP56GdsclH
a+r14q7fr6bOEVSRlVA5jhY3DT4bhMhehsMohiL4qGJQy2pYkXFmIB4t1mJIgRi3fP/2yp11v5cS
QPBNiKyAkaJl8XMTm8R4r8bYWr34QRaeEUtQDUchNINygVWQy75wZu81wtK3DJ3mXJwYkquUC6R8
TAj7gzUWpczHkNpP84o4Otp6MHJyePL0JnV8st2IfSGRI04AzmlC3pVaVXQNerOl3iR6RxDKNXNE
ALhR+sUOgrK3F5fGG+IMMgdcm9hhjq9B3gRwWnCP643nOG2xEjnUUSKnZfYS1avcpbeFLE8x3C2h
p/1nvTDZ+AaChoUhYboaiHHiitn7fSQOVZmcF/s7999N/3g3auK29LnhhxGH/bREFesMAIt/yGZ/
PCoJd4EiB+C5IyNV6UtuSXbtmlCf9v5XkIGyBhh/t7GkFnAh1rA6CoZGELbZYNmbAsjOCSyrMbby
FwGRAYuYdef5EJxV3MSMpcNyc4Bjuy7GWLIltzaU4mAciaoyyXHw9ykzAKneZhmi0WxiscliTZwk
Iy2FEEfMjg0ElwAYeF5mx6zEI6AKuXfiKJd4cLdSdFaM4V9nYAdA1uTIaw5vxnBB+9y3XpD2I1zp
4BFEtPzQMNtxi2dke+TwNfbsx7zCWRxmkCL93cWnqPfxkTuQuRdNwWxCXe0Pek8Pn26Bg3636gUq
xTSkf28HP/8V1lSJTTssg57MV0ld21eII5idZ7e6IrppspihNPyEeZ/SbC3uFQo0WiYsecbi+ENJ
Rfu/dLhuk+we5//m2vmYxRlBKk4o2NoXrNJdggDkJzYjIuhxIj6r5JMoq+/Vt/swS0mi9mFhu34f
SUGy+1Awq6kOvhIt6xpYzL9xQVsjcfkuGnVjGM4c8YAh8ZrCCco5g6WBzWq5ihgu+Btd3aRTbt4L
N5Tf384bSYcaCvybcCgceKfTb4hmR9VwH1Rlx5Y/nqZjCDi/IgsPTptZ/CPqNZQxjWAugiei35vM
Or6HGnKVh6AjSuELRSDnwp9OKPs8YnmAhKiS5tF+OW9pXKgPOFCVtJHZguyeqoRR5ygC8CifEt+5
tvPYNpiGRbgXPE4SIbWo6Zqq59BshXOgoVA35++TUfNFhqFHM2WhTSSph3dLlimt1aXtVznoFv1S
pqkmXD8bRFjLmWSYeJdn5KKJWpQtBuWeJyw74DwXf/avlULQwNvu88+M6QqyM8vxKnnRsmXGOq6j
jVMIO5Pb3Fopfr2UcnKxs/Hcp+1GZS3keJH911KxSy3qiS+zxTbfwtiLpl8rf8nv9bF9dQot7m4y
FifocOSUDewXxR4CcKfaD+IHeNrS7lCauYSLfDEpmfALHFTO23xp8chusaKo5S9me/Ad2MhtaTXL
/EvJiYiaISQ5nlh2OmWQeaeEV62XOp86okwsTR9mWyKmC6N9IWGyQeGUbtaWMDToqfX08BC3359k
dJoGW7lvMWmPKvHa1t/kWoIPE5oiI+eCDCkK8G/vOaRSHUNb/ES/ATrbfBhImv6H5nLQv7qQPGPt
9GkgU0i2HYcq3MyYLj7acln4bZNe8jHHzL8z2OjDj+1s5pwdm3cPluAuDFOhW/eYEPszUjQZ8hNp
+eVP6U/F/KmH4d8NdVcRsE+iMPiZUgd0f+DuF18YFbM7BGsQMq6nmv5xlfUEUjxS8j2egX0Qcvfr
mCm9S4hOzPFcr8UJyWmEsoD0eX7eKfsNYlt88Ocb5ZVfH7bLnv52Z3KMiiM1jZQmptsqELfpkNVy
nPqhnK0gwseU37mnupFh6b5y/3jKhDWv0VmnMVz54nFUA3Zpkqhx5rYvskWmCJ6geYiMstsoxIBR
kc3chMxgoXA+TozOYcL+5ERa6g0wfvuy3bWvc2VVQNePtBTTyPD5ULYC3QhTDMh/LePrj12EiPu3
gpncmOy7man65XYYqOEc3hoU4x5TjTxX54JQyPjB+wZDAMrxYrIFeIB08DzJ3Zg1yAkgUpiCwAK/
+bS5YXzbDForhtv1/AANTM2M+43VUKLP7RR5QqgDQHSGcExUj5hzUbvYR3vsK1sWOoEB8/mhbRKh
G8Hs6s19O7gTPQuSrkpDBmHQjQYfECc2etDqWV2ckTK+QENiQ4ZhjwPhgYOHvm+7F/CWL0G0Dxly
J+EE21aZahn4njdUnn9cbwbAkh4HBWRtkandL8E4J+xaVnWLpOFByX+pgydKjSVeu3ar+Dn55Gzk
qTTgGxADw9B3Wk1aqagmrrvI5baMdzCHi3FLrm/YLcEjh08gQDT93z1xq2j5Rlbu4EtHKCGpvxGh
vlAytGS8/nZq9GZqyjWK+fYOzO008d0lPI9eRI6yvm2hf5x1O6Ono8RRtFStRJ/xKgnbZpINr+ft
rg4ME7l9X8529y+Fb4nEFjZYTrbNGBv1ha5lW2EY2vJOXghxhVNJ1ZLv6UGxBpVsH9RWFYjuP6hd
tB7TIW+tLefREoF6l/uXOHsdje6sc3WiFfpylDtEoj48SietEQ/3eFH0O1cGF5GS3vXKvMXsT9rB
YcZ9ZYvNqb9VZfa+aUwUu9v3iHs/mx33EkF3cj5JdtQMEWL7Jd2biJqsrLtcsDgd79P9hDGsy3p1
U188b4g3M6BLWpQrf41HQ7fDb+xZMo7shZx6scctiIC68GxVl/sJQoHUUnudKAV2ZiJ9tNRfZ+pK
XfaithyjQkctE5jHZRwOpwqT2QSWFQasnuBEuZ4ZISRyfU0Sv3O+n7FGYIpWnD2OpC05ZCB4WrSA
HwieAP8cAYGhe0itx0fhwHzt8U59AHbbIO6LqyhdebHAdWW86A3R2h2HC+lpJAhAqFYIz8GyieOE
d7tgbYxcJxPHU1XziifOmBnbNzdqPFHuWWiUrobY2qdrLvPamxxFAzWkAu6+AoKsm/02BMDMwcY9
2wOjznFG8oHahLkYyTL/weTQ5GF/keMfAolBI6fiTk6g0uPabQl0nYOZroQtqroEkaUpISF86kD8
c3hI9rauZyVXXKAY8zCGggkQj0K/vEpwSxk3KdPb8jNyLqALnpM7X8TgQPHXXu4sSMW6jtdwzLWW
xBhEpq06ku//N6V5FQglsWNJ0RTRgP5JHjX+8TD5XuYd7g9Y0+1w3Xk7uqsruIrb/eQkx42o+M5Y
SERSkec8vHOr12wC5+7iqWb5uV7aqgwVxRYwxlbZGkBeHd1SFmsIMQTY6FZB65Pcgz0HIKIncSAD
Ox7oByQ2XSot8Vg+IKfzNCcZXsPoqZ/M7gg/xX2Pxa/WWu4cglASlca/pINI5Rk45nKnNxARnz1a
9aqbOJAq/eLnXzP65I/xrkWrZRTOO7TtuCsq2xMpBkUet7ICGCTb+Fai32eqAoLQuyVanuXGhDhT
Cu3w8/kGpgXQtL9v+5HEyFz4ybnGgTYQSHJDQYjXuB2Hq20wGADWAu9SZaeHYRJ1ToWcOVlZkPHb
xqjRPc3VLezqMdSO/QKWN0f7NAhKcI5kC4+adg+MnO/4kJafQOOukM9hY6sve+FjNUHQSv6bw3vS
ulteqALVgQapcX2cnVXEqykW7Y5vmowxw9goPWTCoH4SIyImVlblez86HnM/ame5EbJXlnzYakvF
jvlj9qf9h0KM0mXQr+aF9auuMP2kgpUcOsJqA6omr3PIMO2f7nf6Q7pGJXkqZfTl3bddHlfY6iRQ
slDEF932VsBz1lONL1plVhqia2xZ0L2huF0LeenXQOcVOHRPtBTRPmfU2A70JBnzKMRttRplk56/
TJR9vzTGTsGtGt27/HG95FZ0p4YSKR1a0KxUSh3MACAkTRCYM9CJX0/qMEzyvaMg2P8WV9pCeExJ
LMDtBsNIf3Jf4JlZKcONLIfMXJ2Neeh1yJ7n3mTa+zGQj4vdTT5E5tCEdxcxCmPJdi3BbOineeUv
eloK+Nz+1rOFqKfaSmQ5C6N1xk/DfTih1G3+KMwCKeo1kn7JipKNzQIwnT8P3QDGL/ds6zc8TGTo
98v71n/RSi9JH+a2elRDIxQr3bkBuq8CF7kJuUHrEaBVC0IV1aBtFM3+QE/dd9brTnvtoINHd77x
mm/YHUAn57n43fLjRwrpYIlTmxj5hTkRcrVmqdEXWsgblNis7akYF1PWtZrhK8KmB0ggUOsCbk/V
0VVaAHssakh677ck684ZoC3aJEr836jz8PoqZnQ17Tn5pkIJNszKlxqusnYNsHNHkCuUg24Yvy6K
2J8otwkK4n/k9ADa75CPtTqzOlXREbsuH717Iyi0ZMEQSD1h24ybHkX9nGxeMLQ3QWHATlDJA+gy
2R5/GU03yVenQQ4Cmd9CkvG6tx6+yp3lku8ZGDjPV/7zVMnoRMXF3e2ZbBu/eVsDL9TgBcIZqhSI
0EC2rmgncSrodQlK9PyH8BQXvTJxokdp3V1EO4+OevVRyLlUG51q/NQ5/rd5waLzy1OuvyGevWP0
BI42rA1Qd7W0id+QPYx83l/n61WpI5Tt2T1oXtxX8qsgDqtSh3uCyHzCFWMjjo9plyHdQVwGNezY
osloEcd/LGF/WTP7BBP7HExMtzXeyoZuJd3Ggz18MXO0WhTzdLKwXHfK+ox1dN0eow++3/ex985h
6jq1NhBZAmewjKvydZoaWOZL61/W7k/HRUoMH4JxUbYkW1deXrbgpel2Dr48/TtTc8TJhdkvxrfB
0Ca9R9EGxRBYVUY3tkw3mJ3Ag5X9slF02Yl5Ap2ejY9OgkWFyNT3gcOrHYhT2rFMVYMJPhNo4HhS
vuaeTtL+YoXS2hqTmoCFQICui7H4s4rEZhpxA0Sl8hkDL0VwWvGJVDXI+gc+Cv0RcU+tcQJ6WSIl
QRbrpJ4/JEOtqB/NKwP/vUQ91IJ5BiRsUI0QolMIt8rOzVT3zeKmujBf7bTHGGz/jOSOf0VvYWiK
coasL7+xWYTdaxfQfvOY71Nms19cDVIPvAvKY3A6dAtMOGBvABgg22ILxbEavKxxH/5rQPRHVuUe
YSxEpzMWIUqwYsnBrFX1E7QezOTlfTwlEQ/gn7kA1qdagn+8ah3UkyXm+o0NFMLNrt/Jksup1w4O
r1JPEDONwD9SbTGAJgtP/EikGujzTTTJVqw2PCMdDXcNtgGtFTxey4l6rPH3xQQQAULSd7kDqwB8
mXFlkb7/KsXZxvLgcbjDgvblLWRSyzsj4ErQskhSUQ3k1fo4x5MtUFlpvQWQotVcURLm1rm6bi/h
ZyOVHpgAJ5lngDri9lO9ViYMv630xtesevQ//9ueHcGdFWhBFiCM8akJTCuac/LNQWVk96Nlpwmy
KBBwU5ZLwtCrVb8Nrv0uDEeItXL7HiWvI6D+9ddUA41gPi2vtG0mUkZ/HWMvlqPUuEK3YvdDTGKF
SCHa4Ezt+floddlFbSPQSWk/WwwWvUcLGsPjG2Dqmf5WvPWJ42d+DTByZqhL8bbs8GK6WuJuDWIt
UZu927yc4NrT1/M9XwIg1+kMs5CANGzacM3Lkss4CRl1muavbjR1+WB3BufBjG9J6bsQvD3BLbhr
2W2yxJrNBPiIl5lMWL2/4Dj0hzLuQMvI8h7w5FIvdW3E0ukMDIktdslrXPRLv0oYGowzRoGILXB/
VWlllCFn9edzk/NT1yY/DneVXFn4eSRuKnzWK4eLaZO6hNG/P8C8Rcf2teR/hh5TGI7YV0H2tse2
ahDfyBtwGSyhyQkN3pDCXR6keFs7npuGgzhwps/1dGPHnyRHAzfNpvR3j2vHzxBZZfzRi5ZpAlgw
coFdk919TVxVKNSXxR4p8WT7rPd+xJJvJx0G8/mmhWAhfRdGyzDKms6pUD38dD/focdhfS9mlGIe
kN5WGxcZDD2mZxue35h/9ONc0SXxvMgDxlxZvpI7uUsBmmdVK4YPY52iPrOehuAvi05HIlEp4sxt
hBMgyCUtWuqI5tLyd052gHtI9AO+ncZcOimP7aS7o54/eCwJLZf0aIHO+23H9YfpdpzTqQ6lvzsC
tsGmgdtAlXkKsVqfNhGqiHb45yAaGwJoXU46oA4+/wTcsAt5ZULpFIkUiKZ84ghypf8/0awigosZ
OSxns90+IEo8buYDdQeZof9BG1S/F2RIi4t7aq/E5wSjSeLI1mHNCZdfCpJ18rzGXLC11QP+A8ts
hPdCIUvRtodT5aE4y/KsfXBsnsDeEKTfxVmUd1Zc2V8qNK8jE9IDn3of0CuM0VZ0MN8AeL8RryZV
n1VE5MlMJY5WuOU9axtaT4m0yKPDcKFlYNu7Z0Ht/ulb941pAxNvWGIp0Az3KdG1F5WXcRQNXFwj
QPEeB+UdcnE4HvuDi10azS2noQXp79zT3X0rVOzHn5n9CFu8Ay1nCdOAJrtleTj2gqOjZPT0wkkd
JMYffjg7KeieW5uqcU9ih28c2Yor4DtlspFr4DijtN7gxfb1xt87erBsCHp7awgdpvODiU3wsrc/
oo4IFC9sFEZsuYuIpwpmaJNkmAN/yKotpnY4cfn/UHvnFoSwgnWkvuLGEn3gKbX+4BDjBCz5WKSH
6gWPhAMIdMotvLDLA8M8BDZlnIl1Sx5L799qVlV5t9ISs8xMpnc0cAgRHxK1a/VFShmet6g76mNT
B0u4AmotPkriBbgNkYRHzraoU1ppV0mnwBTfWDUi/X0kAmp2a4KOXoLDxnkqlUb0gYs2Y2rYufa8
h4Dgf4AvVeH5vYvb00rGvpFDsA3yxdzn+DZSpMmLINu4Bc6rHptLCyIiFv0Ft28RJyFNubzMZmji
i0vPuvF2/7f0BsKzwhfFp3B7KDSohWHnIRf8VIdbBDhcQ1geJIftQxYDmjGOpDBo9/KKkfXnTIrF
XUQwe/mPLDD2xXkk/Ngf2B0pIzp6l9VL+XyykxLMsfOSKhVJ1rPwZAiqmx+ymvSneKDcfeIT5SM3
m4DBZuALjR02BiK5ZzyhjJLix/uFFG6tYZzNEx2oVaNT//y7VsybIq7J8d3zwsZ22pYdZljw4HHE
q98Fp7UTn+w87sVr8jJLFkHkIFHIUkB4W1+wVXQ35r4OfV5kzWeK0CMcaBzfMp6cSGR3BnynIHS/
ACiLNfYSqQQ3B3Diyvv94uLpxi0d41sS+XOwopC2aTgojSIdsal/XgVOZBn11xPYFl9dxzQJe0yM
/YZjfxFS6i65O38XvIXUvO8iTd+5noTmsKBbPhgkHwxVFi8RseWRfJPvueLC49e98V8ndj8eDiMx
wRHyEn2D7AzVchjrTpN3voFp0bijDZYKyzV/V7TegEDMQn829z45sVDzaYdVnbQKWn41bMxMDKLU
rT/3iDO58WGvXetf69A3wU4bEpaX0rsguySAJd/pYq86yzKpP0D9VHoirK8xbpohGGYDld4QxzGg
OjF75JPhjIBOG17Nx7E72OvU2W4F2XDSTf4Q4Rd9PbtL/ZSLqJRYO/fdGVQ2KEH3u5vV9SNYZbI9
raYYujhVNJbA7nHEj00lXB9zFi9aN0XC2s7dSoP+ynlgOyJHoXvE5pw5YNlO7etBeGt6sT05fWQd
Ob+n3XrCZuALKMikEM1WuxOwjvCZyUMQDj2HyCQoWYvlKdzy3ZaQVPSFJ9ompLoRQ3a2osg+QUbq
szTBjXq5JG/3DZhVz6vXTOKGZidQ9ymRx7W1Mb9bWDzGPw3uNTEBkgHUVSESz4viqowTZy9fRDeU
T0g6GH81E7UH6LA6fIuZz1Tuboy0e2eSQ+qONEPrmhsENOe10+Z1Xx6FV6NZQmepRS8bCc8L4ste
Qn3sMdmqEw1cc8mE/ZQgMb8CzcaiKIheSNZOarw410Esxe6gzkYVqRaF872vXWchpaVYuKUdoDGo
hJt5cia4SMz+y8IlaL7NQXSByGmZIBKZeQ36AipnszNN2XcwKmKylNkcFzweh0FQGJI47iLRaclE
mFWPJnjSoX1WEKlmKciUJ/BlUNqE7W4+PUgG2rFY/fngi8NQYtPrPmqRgh19ReA2dLA39ORcbVoT
MDUkeWOc9uqi5KTxmnk1/345ZR8+AofSHGtrJU2SsZfo2Q95XgUll9xu60UJGfQWcw17yRSNjmSk
K24hYQEjFUZmVxTXJ/IjAPnko+EUSflWcl6C+oaxprCjuBLYVcmQDZ5b/AC2hPiC7xyfORwP4UgE
MU0mRlmYvv+TVfrkp92TlqvHtoRGtvIpfnUVW9V/En5Tlfp4nxI/tXmZilVl2ffUD2sPZNt/fPNV
BMbBfYI8gEb004Z/Stym4W605Yv2JWDW6Udh8MswCLF6Rrk3Lc+1we6wRxXWlq9tsp0qbluM/Tvk
XUP4MvYN/Sj3AkqOWhDwgPEcQ+tagJE1PuFEN+OeCOGC0pPn+dsozVRHQ2YPaIE65a/6V6SnEvvD
7BTR89m6s6ZdH92q2g6ySQ9JV3knmo7LMUaW/tHjnFjHMVosa2cf0L3UBRDKyBsec5QgX+gSuXnq
gigOAYun2yUgQEDyH23dmMAyBUZSfPCayuQpUS/0CHEZ+qUSnBnQuddvVXhIrG3anTl2AwKK9Y6p
/6URe0CzP34ljgAdWBUGbphPDltraLbho8o6sBM5kxCMZFLLXMvkOF5VQyzKyR8U1zPn7fLNtKcS
nm3yApSiQOd9y0bT835493GJ94MJtjlyJF3IFfVLA4i4JBtHmdzrCiM2Efjcq9zmn8k3w24EGow0
pg7ElGEGy83HKb4XwHC19RGlGy/RkPn2Ypbc7fiawyvU0OiqX5QeTuZLjLwsnO9Q1xb80TYz7y2B
WIQ4RwqkqxT/vYOCT5Ty3lsfnyYy0R17+QU85ytYjIno1Tx6xNJ+ZqqABvgeuMmwQNhF3rHUErqQ
dSXvfgNgOLPr++f1xA/d9xlIqCCS0uJKLhI0zmHFw/wh/nny3eNBcm+UGaqzLLyfeZgEBv4t1TvF
CpExb0Di2kI2YTTt6IANF/4GDxtuLto0byhkPxrOKMwC7DmifCEoxvnM9PeS24r1OmTTPU6rqDn0
Mwtd3UicMuKcmdxc9d8IZU9VIN+tFirL0zqeyYTF148yKUj6NxCMHwucgKhMFy/Nm8kQM6IapczY
e4uczs2zPP0K5+P7StPdn8sv36nZWgAyNl1sUxGpJW4aT4LDire0tJowbxO2fdLiRzDCh3ZN6ygY
xzhb4T9EL3PCVZOFySDxVDDEbbqAfNte4VbnOI0EKjw4g2ZjsvcmVkOhRTDsVp2/c/nIT7sUyDVB
wU8FM9a0i+Gw8hW1XE1Sr78DDkOy/yzqWxh/ED55wQABFouPKF5thl2c5n/PZKaaFDfTxu+MxQjK
mz7tGQcBSiD+ydEBNAteLq++lYX2+TyA1H1Za3W3FBrKo0btlCYqme0F6MdBADZLh+jJ7gGqZmrH
SDvMP2IjlWIDvshDdWiBQJWdplBp57oG5QyK911cPDACU9vmikax7y8aILW05Qxb1hHN9s3XMnoH
WqyY6w8fTMd2HQkVa64EskqdmJSit9/nP6NTO0xbn/s5U4AkNTEczy9oXizNSFKOTlLbYP8n6FTE
rc401O4CAYeoJa+YpPRRhhETNPDB5P5YN+HrBi5UET++9x0gpeSibIDdS0Ym99TdlZKNtOrfzATB
CMlvvxW/v8M6swF/+sk4NX92kWl7g10eVp01TJrM7bpfIqCdGAWCMRpMbl/Rg89q7spn0r8PMaJ0
s0w63/zoDEnWjev8WzzqkXclXoVf+NgMgHK9g6KT1/jZ9PABaE37kOkKoHaLvbdKpN364PyRM+rf
+aLJ1G2grHbMjIAcGGV1kI1Z0Yhil7+6E+0ph9xppp3m9UpJZhXk41RngwczWPJq4cIFqPrszqLC
5UEJCcjKWEdYGIW2zy/wWykDDpBdvtTlqZ9LO++iDz2vqKwGyB7PNFeuhbiNHjMd1pDEfm+5bNjg
Wiz7y608i6AxVHq/RA3vlOyGa39bmpjLSrcpsCovUlnmSu239weH7z/2p6Onjh5iCciPgFCFTeiO
V0ubhLpV4WipnJZsmMN4f1qz3CLG1ibD1Y7rGNy84kGyOoUQk7xbNwU0yuCmO3wXecbckKKjacug
VDUmqTCIs9xmEcQ3zqZ5oOLUND9o69ySZb6n0tetLJgS6f2Ujrpw0dWY8O9MBsSNMKYQwxPUV5Qu
TViTuANuMRcWiQl5oi45wJ/AAXOwbj/2OgomWGH4NlH9T8nF18ouHoIAiib7EzIYAdd4Rbo0GysF
spz7vCBgaZ0xxdUrOx6eKZs9mZboRyA+E78KacbbTUx22Q/IbpnlBqH4m78+5aRRv/OuYBApn0ZB
wTdXBr2nIwEAjXZxgfrWNJR4c8OFKuc3vsM1F4PDiYGQQGYY6VSolg+HdfrsXsT4KnL+iEiqX4I7
C64HvNuD0PIy2NJX0Nly2vC1mE/+smAPM94ctlXcuxrwCvCZ4wtKqtQCgptOA1cn3QxlAJfihQAZ
BzDlobxTQju39W8zMjAHdp154NfsGuiH0ocLXk0ePSTo1o2VBxS+cHTb9OkbqdQIr4rFf8HMi77Z
ZEIH60zPyAKrAbVJ7IaijEeMW/xezT4+2RV6BbJgbzt9mLGfOr7xjNb6y/gZ3UCJ3f7ZZCmuXMVU
JWNQEscTCGW+nNPxV9UAJ/AAOSdSgAlYNGtXA+CIuMdbLvkpQdLOtAkHxYQrS1KKHPe1/FclMN+B
1/kiLxT11P/Z6edVK07LtiFkKhh1gs7KF9zsF+4kOD0eW4xkd9FgQOHOdUwPR1Ku/wlOtN4JMpc1
8cWb5qBDgwDeINbf3c9KwpTu9wGs1yYtwIvAk7UoSQ27zEROktT89fJQhfeyliFc+SwH6IQJg1A+
NLcFgE7TOdE3S6cyHaIyZwFyHT/gim3GzJ/bUh78uQy1YqnH29oIdCgZvlDDObHHWmwTVG7FDMS7
ypyVc2TxysFxipAvUYbD5t/525ZDroTjiHfSdEZiB8qmR3mupbO0R8nOVxF5FDNVJkMewyzoNrmU
7yrYHbqk8544q9RGx342yWFL1h5k/FZ/WXp25wOHjgU+MNcN5qJY9ErX3Nfrpr/6xzMnzA6scls3
lxdebtYmuwn547flq4GqwErSXCU2m72MXtZpOxzsvu+Big+L5M40DhYZlwefLYXn1cE8xvUpLn4B
1TJjR7HBkRZZQNmu3rWEJ4h/5BLnTpchG0woTY1YzD443Jq0chqHBUGqPyV2PRHu1Phm1Aa5oMqM
xJQpl4ATDawE0ig+6zTZZn/LkkYDd2kK2TRs/gTdA+LnTZKw6piI7wCUK9pX1tITFIIz7DRLH3dK
i4MUwGK9F1Q/QMP76QQnyCby0Gi0ShCt4dq4o+8tIhIJmKOt9JkMJ1J0JtHHyZ3VvBOT4a6CMRbX
msTq89u/A8Sznk+OUtgfAUJXJMjkXDSyq/PQRzkd8J1E28WnA2GAaPF0DmIBxdEQu+Ey3EyORjmX
6GTDhy3wvHZNGpAiLd9QAw6ZuR0t1isTJfoKyJVwW3vwsJojDCKvUgM81QCWqcwbi+oxiaI2rIAP
RpkQiqbfikLT8P8pe2p70oZoZZhIbxwKf6G3LDRG1Pt11YkOiCN+KZDT6r77/ba/kjtomQYD4Oms
syxmGkon+uJi/4f2yVS8jYgoDqEGQdxc5hyXFadXWauS/u4Mii4yF8BD5uCSRXN6hUs+4a/zXzZP
si3L/XjQew5TZuHHly5pFbGMMtJ8yEqyMXW443+sr12yTylIzdSzOOpgRjwuFQnCYB0zk3Vj1xek
o2CHiFTSMN636BcrGKEINHDCo13dLjDGc6tEfKLuNqjmuesYi1MgJMgrbzIaF0xiM9eve/B+7eJe
5G1MQjcIXY4pJSvvhIZp3oyyXFHnXocWsOJTHqsIetp3tA6dyt7wUWo02HRv2raquB0lXqBUV9Q2
vqZzXkaVzf1nhlm0q4zmInUKL5TP9HehqkFhEIJ4oeBTHAjZQnb1YLOsOpzLFJ0EeS/f3akyMygw
2ytIRZdV4yEvM3L9IHL72+hdJHo4rHF8CKisjs5kwUzKWrxq012NODi7M+T0eWV8vg5HY5bpQJaj
RlUa3TZLthScGo1Y67hhiXFzy+EYGTTFETUBwMJ6liFb8Thl5daybLZqKit4Un41zy0Mt8IeFuSd
whc8ddKdsH9XGTcnvOQLhaKRxIrAcw+UJ0WGfh0iqUT/mIWnN5h3I7A1EBjQGp0IQvh/6HRlyJTl
pOrVDFq497jjWsOkusxx9USWS+hsrKQsQUbDDLciabXlW/zZl4x/guNBFtAoR0hv+FURrnQOS5IF
KY/Wrrmdmavp5Fkk+wp0HF3FZWkZWSHpWm3k0ZPG2MGXyXkkfVKn8iRiNMDiWEblokkfELvxRj7z
x7eYrSFmAegRFcAqfHHhllQDw8lB/mIVg2rnyBdF2yidwddnPb8jZ99RB0Uu3IrO5Myrcr3c6iME
xlo9WqwFL22StzfedZE9Zj4mgZflRjD5IsWEFcL+Bc0TCgTHm7oD+ftLOThpZiqBRmJYO6fK6QX4
6hJjHEuGV+k7xfPSOEADnLhBLJR1+tAHEmALcptQRNMlrNe54lzkIDKzVuTrxXNdThWKyZQNvN64
m+G87Asmv/vkfbJ2w/QNAJQJyk2ZNpP4cln8Iz+z5tVjGmjqdM5BHC+szNsscHED7Bu+1zC4ATF3
zUwj5tON9yxSic38CrnwmPwt9WUD1UIolSzfQ1q3YjADzY8EGnZ+6BWyfAfKMRECDdBOqdkgAJ7+
IWbSk2EPDy1jelE/UaRP5GOg7qaluZ8vc3TAE9wNr0eZ3czATukxycwDUh6kvuDODR1WbrsKTaff
8xq1Xfn3ZcQLw6MxrxHlGUAjJoYJ3Q/kLj1157Rv4pZF+438VStwrhD+Bbnqb2jBrCpL7yZA9n+N
CUazpPtwZKUoh43sb+ifc/d/quzrOmffiUm8ecidHkiLoGWnaj4NHibK0vXJrfQ1pRhD1jOeg13N
qod+KGx16j3WiNJ+2OIO8grS99qD83g/ym3+WV9kTOcRpWEu88C6QYInJvuesaNPgarSkHOMyNdW
guwGhgw9hUCOgCQyiDFNOlxzFe4PmoD939rdfin6P5AM00jjunCDEY3jxVB9YYrLsad4Tf3qCLKh
I5IYy4bCn14KBAJcS42ndeOFrqNLY5MXznJWabaLMRox34Ur9bTzibyFcWXDsYImWsmu9O7NaNov
XzpVhQBYUYNXpZAN/8vYMH8/+myR2A6xR82Z/Txrw2UHJYYXzs6Fedp+x7a/q9TU/8tqivVjxHaU
CMET9wfi1BXfs4VLHC+yGAOQgUFqIX8gCokCSdnwvGMRi3J8wkhP01FJFES0nvy/PTHgZ+lozJk0
q0MRLOIlanzcAU8yQ7XLaqMZNuWzNKBCwBo9mIPntlS5DA3dBD8WeRZiZxtot05RuBxIY7BQKlFf
2rV3le8jJDms80uOK/+HbYXruhYJuuNv2eYLBg9Ds/fbntMhIpKRiq9liw2PqoKxtd9P2Zz2Yeg9
hNQ9STfYVXH8Z7sKHrAWYzVwIqDLwhc1505TUUWTFIFOfaoSu0UA4/oaDIPbt4YDLVYRbaeqzoSO
IMKODTMKFQOCVZgE93xdB+w8RoP9JoncXm2r76zCtKqSEFklU0I0m2OCClrhtVOGf11MWGPr9clX
BqGLjqRz+Cw5CIuL1PglAYXT5G5E0TDz16XStPgXv/3UMnJTk15zzzug9mFvFTPvbNgYM5ZDozT8
DzL4yAA/ILnm87V4EiMZZ8sUvurrOIxwH2ueusWFCKvyG/0kr5oha268mQ6fwDf+HCmsP4WzGYYJ
dKfW1xW6Ok3C/PuFuFYC3r6Hb3brz3qaQiOgl0DgWb1EZU1zWkVBQvX95Hjh8NfIsUi78DlLWvqI
SuCPXQvEYud+Ua9W4FGWyDh+Ak06jfOB2DMcmMAJ4tMUAeE/3dpfuDvLMFytEZlGmA4yCeAIedel
PZ/nZZsUH1RnIEstSgfH16t99Lq9R+Ip4wmlsIReR+nCCaY35XWBrcMht+kghqg3fSJXCvTu4l7V
LoOaxDbaoG6tQln7GnLDIHivToGIyrUldteqhWdepxv71S4+Tl71u7kzWRZBhDGAugEbe/KH5DHz
D7uIJ3wDysSmxdcpDJn1t7kktisUbx6hu4W8h85e0NXIbutHKi3tQ64KJ47NeeQ+NHAofv9gJcx8
+rzBjsk8XwHsm/5C088XN5cn+BslA6a1sOfCO2mKUlPBzgCiG/1p87BF8Lk/jELfHNcZblTcZe5L
3xXu0LN7BvUtuTyARjoWH+iw1mkx+9fAMcljiOFVgDtHzNxLvch6H2nP6k2DXRWBzB6yWgDS+PkT
E2jOGZAudwBAf68+4LYSm4pqgJUBC2TwFtcHu7KokrIsUIuYb6cofjhhZoQgMfJ5SUKluPiWvf4l
81x16TF7Lc5ckGuw6JLlbNeEGLk6Cf3NvQ1ho0CBr7q8m/oW/rn6nJ8pdfk3ZgAHRzp3B+f2WMCt
hoF6Qg4be/eY9/ul9gv+qDRWrciB4SUui5iwWcFaFtZoVoZ1Rtj29nktD3h6h3zRbsbjQw/2prB0
QHjPWmxOl5AKrdcH9MxnmnZ42nhtiuAWjks/8ZyUwqRTwAhvqYZq68DFErFKQ0lbr323f3mIZOR9
ZB6dWW1XkLU1rxi3lcdZXb5OHkaIwtQd3rb7iKOe21sIreZpfR2sh6R5AidDzAvSx/q8G4GhCic7
CLod0uwrmlO/CR/kP3+nnEyYYZXyN3x/5KsQT1HnnP+mD1JtmVABGNLXQgPkOCXaSHrEBrR4uLzO
wCMfOzM8oQ9nO3ihFluQx57XsknnQUlO5QvgEeVXyFL/S6uumj9RSdkeKfsbtdMnVWSCvzetm39G
l9Q3ROF9grXy8SHLn/+DIPShS1n2o8bqsJ1HvwiAIsPZ+LUTA8U4ga85F/BK43JbF1LGdyUcg+DH
dNQONuehNhSmj32rAqcwOBUxDzg/zJbyjcE0Wf47Uv+sux2TV00KPPhptiZo1D8vmVSD1e1QAXu7
ug1ppqwKaohTTnPU/983XbZw+hXPzQcpMPAMvppvjXikxb4re0CJFp4drIMZO7DEl/RjI8Jo/Gjk
AfZn7n9iTTnTyhk/TCljXhEnKnAu4WkmF4qcIqYQ2pNxYOzwVEL4xIRhQoFrAgs6MkIt7FOwo0DB
/p4SfaBShV0aZgAi1zAR5xZP5GKIji6XR3RlkrL64rqqC680O4A2N8ZmhaIYJV+u0+R4mJwSp6Fy
lfj4BB31ctmaESlKyxTIAWHKSmZeNn5EoU7EzYDSZ5pVya7P4pQMCiJqdPp8M+cW4olooRK/78tA
w655dcxlf17cyJxwqDHxI6N5Bk2mMP7aHtSKTdiC+7ZSxiqDW3YJn61S5BYcN4N5zvbhq7rFtcuR
+zMW5Q2GGl4BJuSNWehFB5pjGz252tMYKWthmg7cu374tW+hN7FR6O+CLWvfQkdoyvSbGtEkQwKd
sQR/5W+k1a+FMG6uNz6QmgBLtPon+8BM8VcdfQ8mHuM/myYIgfO+s65fzGGj6qAB9RXI1ajb8SeB
3c/8L6nUbt1v1slWe1lW9zyIsE492mbPkweYXMbYvn3yd6Ve6+x2yRXuv7yg3F145kCnnYMEFauj
KRBWiQd8Q+f2kgXvORST4htJ9Ek6iScytIaYUd0wpWh8ZTczwP3mX5dh1XS6posI2IGfsObOOvCC
/5ipgs0opRRjnTTRgTyIaJ1XjpwZDWsg+U7UPKXqqD5e7yNr0dkuIEPcq9KcHVuNUCoKd6BCPm48
Gej0yBHyhMN7jI3UWj9BGresqaoNOTxn7UUSjkGo7xvD7nz0XkfuerTFq8IHYmAC2UVAEdU2n+4D
m+2175i7AGTJAnUgmIDhga4PckHmMXhkXjfECgHH1D893ZinfdWcmHqWGCxZM3Tn7r3FcUddErF6
VR68287sSOz3eCIEHc/ZcL+UsDZ27YBVLUpCh1umWvyiI90JOM5mulZXgyjRPFvvPSMg9NcervaC
2RsFgKj9vBSP6Ok50pq8OoaAnT2W501YBsjBByKopxXH+AxWTSwvViq8u+03YYNlxm1Qx+LXhFFh
bhk+YcRezRSybG78lGYprUlC2zHwEabc2OBwxylzNW9TyrPpwiKcXS7expIG53vnprbVQud1jPuo
imyMR40k1dKU0r74WYpqS1A6qP9rSzkRTvTN8BWepNbYGt9UjX0TGtxP0uRo6nrKIpIuFtSjchI0
6ajKFa7cYOpu8gTvF3l4FFHUXV4EmnBCQxSUxRh7qTql/wlEd7jsQaoepzuJi5N5SuXNU2ugf7dP
873QsF5Do25MCW7KbD4gRBAhLRR0OE4VgKGSAqPhEFaVkFfcJwii40RGv2l2tGixnsqa0UJpN0ag
6GK3MYK9QlFKDCFevXfcKPryzPfZkpxXE6o4UdXvyWnn04QwBk526i3xgPs7LMz62rjow9u+gfo0
kLwWa52xNIHic5iZClbgknuiw/JU5xPm9P21ztQ8nOQTsCqnO8hiQTLNDWqbckNHvsOfCjsTdRpE
LNWS5Uk6rylSNGtDuA9l6tHj0hKfk05l69RxZDrHdJqn/IUZXmK9aWhGVMCmMnmMGaHgZcevCuzB
D0KDFvrunf1r4EShU4wb/+CUBh+0QJCKmvQbS5ricbFQGvNHwzfxJgUM6tFrOPy3BAe3vlEWmzuX
RAPEw5CCZ+y4uzZDpeK7Zr9agzdbwIRaSzh8dxvsqeQTqfCgNjoci7Rje+zZbXYARQTnxfjfbmUz
xPy5BbWDGbplnUWD5GPpq2YuC37WToFtEk0Cc2RkF2FpdIzitONc2OJGAChs5muPWp2+jrAPsduN
qHGXBbawFIF96z8B5ODmrgFuzsCgU+FvBeGFpcUMAJouWxRJS1fsfzKb9wfecuBx/HyTgJKVrk05
eZfa5tH5qd/a70czyZw5FAkT/uzE6+ilCcTivHFoDV5XFcGAJlruKEdEXAsX7YTpAF1KunkP3r03
UhSMBg3X03RWNsm7zXz7h+ooyzrkONMR5KSup0F5u3rYk4ePQ1goTowWbkzgHr3JHttMFT0v1IAX
Lcr+9BviPA0mL+5sTYSm5yRI15EqgfuJ9u7PUhfLV2Eii+7bw8VQ1AHjz3BQOXeXs+9GgdfgoE82
qcGuOo+s+FFxbJ4uSC+rHcQLkIkseGel3uFqiIp5faG+74sJJAiThA+7qr1GleQBHrSMkalU7P2Y
SGr1ZGuNbMitlbvRFyVVy4W4GU/MWQzSWM1/0rPmj5mvFkXlvMjXNtHVwS8MEp/EOaesaZzCzjdW
wRTDXbowa2UHdDAfrhIDVhcB6q+4oN+O9jMvXlR69xxs0ZSXUQQggnEqyz4gWOgyy2mwUpyTLT+d
Cp0/xmWHFRXAhBtwPc0HAQA7skzS2qx390q18DCDPzvQQSrlbI/bYNcgosvfIsdwD8HJmJLjT8Je
onL+SoSVenWyMe6DRbVDLmb+Pi0yeXdvSjWi6sC9bwdnka78tWvTczQ4y8J82X9iaUP/15H2Cawr
qz5Rs0LU5gIOSdJs+87JkoHXrglqmh1VywowJ2xpRRxYf02nca9ukhGeFmfIByUvOmx2c1Pb/T82
+5ABWRLAHiIFXNb9PMXH2naW5h7X3nyY/Hm60CBtSxjs4MnKD3BzuDzJQyK0LCAty7YW1zTAKG0m
IYHMstRnFpSocFb8/haE7eg8zCliN4h4k7vHqq79vFaIROTsvPzqby5HGY3+zBqKQKRu4U8rIaLS
FjIJUu55zvzyWUT5imZrCYlqkw/9SDRmx+5GFWmmHxpMkDymDV8XLBNdZY5ke1zYXAsjCpKuUYEY
aXxmSQH01NHmZnNtot2q5YT2ME+0YiDZxJdtMenzvI2zpKFqsFJ2NxBcb4EEiLM2q5I8rSbcFf48
newQSBwKEn2ZUtkbfCQLc5ya0+sVJqAd0XZakYotlmWfHBaukFDpsbiua8ca7r4rUbxbW5W24Jko
mEcoRsPj+9cqst41AQxr+/h1h1lzMgBKO/gjy3AvhOki6b9tCBPyOddPmqxFTE3srkSKnd8+n8H/
1dBUdQxmrNCmYdogn6ZhKzPoYuZwyFJqy1yzyO82gZ1YIpAc88iLILBRqm+HVM8pPxAo3GzBQ3Rn
rplZDPljw3Sh8iiN3yt4faaZ9+zbgL+mAAlr7wDbFYqo2gYfEi4tBl+PSTjGPLzHMyeTOFbalYxq
F6u50g7jCOM9m6pgtJN8uEfgqcU93G3UFGMbqDKYj/cxFP5kTMkYHrWWofqtfjjsKzgISaGsSH7Y
5y2JO3jZmOm179x9sXPYAMrWTV6Q7Zb0Y7VBQTKkhgN+5824y9tPFX84eY4XZ/kJjv0qoxRoTrDI
/I9r/DJR6gM4UE5zwXQBoDxEtRBWz40IJVo5LdA7Rl8mkUdvG7XBX6P4MpBFOSGSAKxzYVBCOzPM
ifnFhXVElPStcly7csQQYHb4n3hP0ckRW407taRqKxCiEW8n9E2mGEKJPUIY3+MHIfKfjjP0jWjd
CTiDzzqufSFNQ3L6HyjTYXIsP7o1aB+moOmBxp1U2/NJn7XSBuAkg4v/7rKrQ3mFYqm8h4TAamaS
5OWY/OBQxBK4Lf7/tR3Y9eBDOeIz56Plbw6iudw7eFaHr9tMpq/z7yMtRHpbtIJcStezZ1HexgDT
w/Yl3dUEVXOpJCf7IftjI4z4BQ8wFSAodRRq5/uBuLmOs/5TF94fianuRxDtbiNgEBXV5qn3iAcM
tAhq2+3sXd90oAQolYTk6e5z2Oq5vW9XjVNoQj8ijZgy/LvG0yaakd60SMEC2rur07o0H+BE9Kom
HCQiIc51+qOpKz4Zp+G4BXxVUBBYRq05ug0UZgl7i2X/i0jPXhiG6A1ou/OdkfdtZ1FvvJ6C72PN
yIMiwcJhFQzO4r75VKUhN+awFHtQpRgL6g/Lxmfw+v4oekJ3brEZiCuODFukgcSX8jJtkAlEQH6k
hgu1oAkCU4f0A/Qwfx8efPtU76Y8Akg/Bm5p/3iU08cSL+R6vv1WJETYiu3v7ZwmGj52dLf9eW1k
UN4/AITK6fVwF34GFwDXJDceBjCJx1s91bM9RWXZBDC/QI3rqDhkW1qx2eFJ1pB8t/vio59snyhc
QFpt1vFPPu/4JuQeH8bbbgr6eXgX+G03ST7Vq6vDPvUf9918Jb2DZxAxhbEu7wh7Zd5ZDwNQFXXz
GKRmv42OrJwbPOizXuBSoWdNipYN4ICReCIeRMBfVrsqxlAgWcloHbv2uIVR9jyg2RS/IYvXCIZq
vPHEV84nqHbBR4QkxOwnnTsftUECQOp79WXoHgC4UeurgqK9Ddd6zV2bEAVa4DfyqJZpjT75oe+F
uxqX/LfgqzoTxOhVRqql6kC+3aE4Q5FNEt7xgPI2wwr+Hnieqp+ysEQzvM+DglVLbQYlSH/0YOFN
umolvdJrql3jdQSuJUj7maeffPfOQV+uzGxegcBIDyMl9E7qf42nmHmRcuH8Togos7VeL0b0bofw
pjmZuhIhctoZRWgzVveEgpfTXhSfJAc37otY26QFikaPOSeVsDymQO0O9acDy07l+ymwRAbf4Gsc
qmkVdRcyDQoNxVTQWJTNEFEdGBpetvEvhBgeTJ6e/mY9zaddbAgUjLxK/Dk3dUQqfOGIZ4M8hSZW
d23Tq92XVDONfdi+yGCLrh6yCDxutDNSbwl54p2zgtMtW/vV4xvW09lGeQP7+jxmclKYl8tY/4m8
5v5IE5Sb9el2UaJg6e0VuvmSfWi9gggk6AU7D6IRhE9OTn8oedN+DNWngu4pKaXkzLkbYwR7ts7w
LJDbBe5Im7VYIV2xer0hUAyTi2OY8mkmVOmAKIXfjV8xeD84mBWcN2oRV58oNrBtsqHlUfHaFL5Y
m86fDw3B1uCHch5nFYeqopDErzXPSsmOPT1O8gKkvmj4CYZ3zBcUlAVYo44o7zCGVV2H1bfSoCSR
E5COb8yLODP2uXRm+u8TKhMTO4ec4uwwK1K3J5zD/vI5V0twirbyoagw4UQQtkqN4X+Rgg3o0VYW
kJjX2WCkrI6fZkPrkoMEejClPg9w0yyQIS3lUfhHbSSY2DSmcysj2sr4nqZkCGYQS3m4R0rFMGGm
Qe/nSE6fBjsA20LOfl1Nokz+4bs/g6vT0Nw/O0ywjsxqGvzdDGHtySy9UwoV0M6fL57n/3Ko20pd
N6I5Z4GGfh+WFcqny1rNSTS6bXO3qua9D7eu0O2jXhEgxuyJeWHQdq31XQcu4bI0iNRCdg4kKtnE
YlZCrInREXrWXDLAePbaIJbMTfttv+64uG51rZzdzdIkhvWkESz8m2n1knQ/EjS7jgn2LzvcMZbm
CBIz4byIyBVxKyNgJUEVdmvWpSJTv+NwIEJCpoD0FweR7dPn+0Tmg7nUDxhr0ezv0669kCgANZN7
23HCW6tbWtklF8MSZryAH7zciVCEGXDDnk8sUdsmvKUkq6D14Aj5n3i61r40r4L/3lCdAWIDaKJ8
rg/UR3ckf4Xsp1xmHDd/kwZF0LAl9lVfdKXbCT4ZQw+oHALuzJvWBOzHPqN9qIMuLIyZZsO9QVdL
u5cuOhDnl9wEp2kEbq9Vbzk7GhRikVSybDSDcqh1TyJ1jVdwbioOYxwDCJM64hAFA/J0sJTWVsFQ
ReoSFbSA2M+Q01sooIDcgf+NC/7Ub0CrDYBG/g3P9ALganPME7crYNbR30A0F4Y2w6XcJBT7cckG
UAo4MF0ws3GqMZ20k/+vYSZ17bHoxz6of+Gd7NiwPc5HEs5vdYoTT7RsBTcTQ4u5Xw6UCKegGpq0
ROvPcUmN1SS/SUIPtfHW0tL1MeMFIDP2YZuaUPowzsLHUkRWA0qlXLzTYuMYIt5BWRdsm0Hdwo4o
Fw8aGrVckSJIUwuwvOJXbS76v4xxsoLIhBfDd/Mp7pcBchSzg7Q0uaLK9sUrCHG/oqIN7BMvvUgU
UTxunYZ+7GYYqlSKJcakmbTN+tRevnK64uwUe8RfLhZ4WYpQjBXJgMwmOvisrPHklX951tYccKJZ
SLt62AQp6IeZZiYuFnZghH3NfdzgS/K0mLoL8A1PzncZmJ1zlHFre4WkyOYTA5gtkn3L2vIDQt3j
yxEicd7mOZ/Y4BfTmCbpS/N7LIso3JHnz+6R/hHItANbv3qP0YUPWAFszkoH0k6RQmnhtCrJqAlD
9Sfh71Iqf4R3dVDD27kEmR6BJ9OMS2m4XfCRedLHDb7SWkM1QwVCeC5zMKQ3RvUDCI3NVizD/i9I
dSY0a7TS6x2NNzJymrvpLdJSQ+ucSyeeyyKg9hORZ88OeSyo3BcQBFhF0qvr8KdFh0nJyCU+mcTZ
khG7UYLqg5bKuPQXgrdstz3OQKl6VpDgfVs+Mzu2BYxVLEoFc0j6mT39oLzVL1OChKNHWhRUydi1
jKoyE2wNR7gP0u2z7DvtT4mKDbeI5WV4SgGNidm5U+u4vlPwPBGyd615xPJ7kryBbJ/MXptIP+RQ
R4Oey3d+E9qBM56MGcZmJH2S9yAuKzGdklglbZ6YhydHOXCbb8r89s/au3zsb9NccJnpH6NP2PxA
oCgZEhebXJd4jZLB/qovvl6lLr6qupw5FRfTSD3+49Jmh+EaKEOz3DdPAzX8hGoZVPNkgrWZ1/zh
I5YcvRKRmEBGiXIonflDwkM2V9py/pC5qIj7NRVr81CHzxBfNgnH74TAeobKUlfJhAxmYjcs0e0L
4tfUG/QCBEDYgWQ+wC2g444FkU35qkp1hHQzkYGzjeFaz55IdGOZ4R+Y3avVPJ7IEHSFgLkfdILM
TlhXaFv+eco2MFQqk2wyaIJKsg3t1UTVuUKVm3XgpmSg4nSBGUUbGjeNPvEwNKhg4bFv7tE1NQpw
AvceJ/8BAihoQ40VUOrqlMaCtxDOff8HFq2um88lvD8BS7DQfyU35F82iBdd6PkGo3WlRERoSQwj
aCnJ7SUpUUccg576xffh8aTTjAHfWOpBBflCGYgskf6QE9iTNvVRjc0DitBJnUZC+Se3DQmZHjC6
www+TxurFa5nB/K1m7yppx2ehRW4mV3gvfcB27sKaoBhjY+Xo1+FJK5siY3128x/CnnUrV/Y7Tri
7wrB0D2zq5JmZBsF70JlL6sCJ2/C8Og2zgJSRr/W1H+1feiN/wCv5z9aZGtbmA4rrtVEsClYBwwZ
DHOnN0pYPPvox4Bb0mou6Xh6LHFcoEAPp8uHmXGXELrV4Tg+LnChyLTB4naiD2A6gUowSe1VCTWW
nR1hLRsjoZTBepFc5JFstRq+OL3tUE5OM65Wk+Gkq/20//mAxE4/b6UUU2br1sEinmwh+QtjLE7s
EKiNn+z+5qEKV/imiclTfXzinAXoruhO/VuKy0kzCWHQRpsDLumk2uN5gl6Xu2ASH7EDegd96aqc
1Bow6WtzNByyx0c5cu66UsVrRAShWPAACQYRJUpvSNcSr1yWZxOFkbb58RxN85JYKfQDV7mGMgi4
3J4fAu9QniC9Ck1OZJ1rmQdkor6Qt6MfWM6spCGia6H3GOwQ0zWWs4B2ZWma5ItkrFLGqzzs+bpu
qnUvTUhsvshYGXnDTL7vXLvPIVO0Yk7jtBD/TSvzwuXHK8DbLUDSac88jamnMOS7v1MpTepx+TLb
6jZ/k+NdRwHqVlBFsRREohC9dLpPsKhf0zGUxZDfeP0BZP4ERgS4ho7WvgqwTA4zp1gx9dBEgvuP
0iYzB8U0S66DzU1kGgtBAqnhr2e+03aqlXts5QfwIBltFe/wpYu12C0AefSXsatTTftCyvbfKHx5
eRh+++8Rc2NYcuxe7HkIoe3Pf5D/yiTyEeo1TvunnHoqdfutD3F4Im1jxYGHcHTYDIamJZ1JmooM
467XPT6V09oNPY29S0Ej0a4THZE9V7kQ4ukEVoBczdi0exwCdVgsDTyPk9OOSNvioXIfWEj0+fyX
yCKxP9IIoSs/ELuFhBjFACmObFa8Tg6ZuXf2pc2d5IslndhgPTXg1oiyGL/Xp69DN6rHnyLdXBUH
KckVMEyfCkb89ueZzZisb7p/iZ8ewC1tPkAatkHPH8HRa2AYPyoOxFZnwEar2M4GHbb95hOScSQg
JqoZakzTR7fvXGtubKWVKWaYR5M1NokUsvcuOx8SL+JV1M6I4dB/D4p/Qu6XyUvZw4w0UOLKVLyE
bYYVFZcCO5duDk4+fquYtj3CIm+sZcqTqjsJ2IWkv5uU8PtNFqieuimFFsLBnjv4jcSg9EpOz3Lk
hfeZXD/gMiYpjEs03iMP7j8xaarAByWynMtcfH6vghleGswHezFVtTthp+Ci++mkagmDytTR/aFr
s5qfOgkhbAp8cBPHjwh/zL7EaozhKlZS7AQ9nFd0hSPeo+4aDLOX+uxudJiz8lX4GH0R87CQWvUV
fU56j8T31FYffyoVrRptjzIZSmJe7g3/Np9/hI0oFCEg9xtflfLyY5FjszgDDjeZLjILihuLxwvV
d7d+8+fc6LxsHxE5Fe14lkhPo+LwzaWEaa6fi3ITewcS5LzaxJWfbqotzd6qQnzxTPtfnPR1aqbg
Hw1HtJ2pONEn95yigi8yVSUOtrYz76RYpiklSQLYAjCYfp+IvYi36f9VhGXdXQB2+r1sMtXJekoU
qS4UBu3rVuYwx3kTR7P+bfv3oERkvz7pvg/ZdlD42OlYMaazYyYT/yRepkk2WQDRy2essurUrfND
XfbsSKaRruAYXIcUgEhQ8jJHFbysViu6G7nMQ4V8VUjRFvxvjKXfyLyKJHPXfTkoJBhWJbKID7w0
Nl9wPKBgBn7mWNVJ3Xtk9uxFnreGr5KRMMVg/V5UsT2he6rTVeYLiRlvJUzEY+olp16FRAuvVTc8
N+Aznf7ts/yrICuNy3GUlUPwLaMTSi+WhooUglv9g53oqbvmpS8LKhQ3TFsCdKms/N/KHv3KsJmR
kIG8ST+uGhPwJbmiTuF5m1mh3O29lTmXl4Y6uUcxc23UEETxj4/ZZibOWY2D/WyeR73RetBbcS8p
Z6Ys+33/Nov42HvnHjY3aXUP5VVRXd+ngktWhCSalLZGLi8jM4qy0lG8CXr2p24DFoZqXwfUPmDI
tG/TGnjbLNKYVRKAnZL9sjLcD2BrBzZqBfbkJpY3mOcnSw==
`protect end_protected

