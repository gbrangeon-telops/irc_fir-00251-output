

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jmxpJaVr346lkZ1a+LoDVE1gRSFGUifNjtRZEnGV0oAexMx3qGrmrMofcjVsktZm1VmWfXDcztXM
2yFG9i0kgw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dOSbcKbKyGmwastHjwhWcvg7mo0iC7nVbxSBuuKDePvzqRHFROAJKKkq6GTW/pekpDi7EYOWgoc3
vu3a7xd2BbB8KPxJrQPbDcHKKLsfi9Qu05pG8kNfZPTmVPdeph29tJwJuOY3Bue31aDGpBx9n97J
il8TNCf+vPPl3qN1O1Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oj1u/InDUMUdQbb5KKzCbe7WKv0Q1mJ0hkD57NzdtON+OYFVa+iXuwhtetuyEkD/RFkOZub0bzay
EGz9mYS8JrDX4uhqviZ/lNeQvlGcy4m3aXFV0BaNm28dZ3yofXU/BObQHMb2AJcvSvAG3+NK2bRe
O1i9rDUCI7L9zpBAsqwfaKowW/ytJpmf9i24R0N1DPpd8Du0b8109OjIyuP0B6/WOaUz59+u6rpk
YBt+RO2we5Eynllzej7EOx457Zs2AfpyYb/scT1J2gg+ITQOiXue3l6rpuOlPDO2s8UVnv9AEDol
dBES1PgrY5H3iIxtkySbQdPn1RgrbUXGoP3Cyw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nf7SNu0SV1jFULe1qPx1Us0aK2tBb+6HkavjcQAOW7vm2bkkBw9TTTcBYW2ZVktL2qtI4SdzYqok
Ur+7+BvPVL9Si1NxET/7Dtm+YCiSnZRDjVxRHT/nOJoMkCyfwzbKJ0c94Mhpx/IIVydS9opk1YOK
norD0fiQ9NScYfnzaaY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gGrec2cOqGtm9E1Oi+bdp4JmEjroHrWUud/ZaF+TGsozi+qUj2kRQyVPKMhdue0iIQELWZ+mxYUS
eLZifl90wtAXYuJxD08Z4LzdxHrYp8+GuCF0avDcKZR6UMS6GdOF0ZR2WdDmkxgQdaVnCHNmLABF
3DC4E9wBUl1YKYXSRH2xT5Tm/cD2sgS0Uobvp+lTtO/g/wUBgQClX1AYzm6JvXG56K4a0tlrJqsS
O19bJe8ailtvTRagvfU5lh5iVeppPrENq5fwhz7scUcyvohRe2r5jixGcPz5bVE78eEpH4EwzJTz
GDGFrWw8qJ6s5hJeVjOB9tgbpdnAFcvyrMEGaw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16464)
`protect data_block
qpHbUod2h4hcGmVgJhvLxo03SjdFPtpqNNDg5QDXAnIv+5iPvt5uhnDiM2NSHSwdUpC6NPEg5FIH
0Pj4YVwz3ew74YXh8dYTWRLHnRVn9Dv4yRQGPkojNiIaPhNy3/sEIGmNaG+xqPpzkm6OD2kG7IjG
3tsHWsqB9DehT5BxAu/I6XadreM1YccALbB+/x1uDBE7FCmRV8UKCRpYh/Fb0JiK3k1dOpC0QxhM
GGcbvQb5EmNqzQZXumbBkVvdKTnRWLTB7Rmp8aChp9UICsce9Po8yNKKKCkIdGjvZxKODh0MjdTz
UNBgf805NiToETm1GihkPmLo1onMq9jVb5I9MChFzC2i61f46J6//yfZtyIMkocfxSH+B+fEdbuK
cOU87ODcKZ9/am0nxeA2szMe+zPIxWiscxuutCvSDWhhWYnph2/yriFs+yt2AeJOfFfGqb1OOTUT
MxeQ7x82Iu7foEz7ydBOSc5IqwQpeOOAZwQ5zJYOLHSKMlUCw7iD1GFccF6ZWU+giOcXda27Lvc5
iWJh/4nSzokZAOqIfBsjWYgvDJ9+xjj7Jo5XJrfEtndJD3sPtm+/rX+ykKw69WXkwBp9sZvZQany
CipiJ8N4jx/7WWFlKxGs6Q04WhSgopd4ZmiEP9uY5lL9zJYnTMs9Eb6UxSRKAhoXQR8n2mLWC6m4
64Txh887itY4aVypeMo9YA/o0HmrmD5gSa9KihbP+R4PK+Riw8quUpM4/75YLjk5l3bRrd1JFXDT
8aXLPq0UBpOzaAV6Syiojrd9azXve/d3R9OLOQWitY4BOJSA2aUcCu7vvoWTmb0xtVO5abD+uX2b
GST+PU7l9W2iw5ONuJW25cYTZQdUBBbNoN9/I5ZcGD+I1oIcT6hFjGrbXkHtSYm7vrFf9zvdbZzk
HLYwKx3pwpDWEOdUDlNkmsB/Lg+BFG2pwdmQphrSX7TVZyW1Frn9/05ZJZsCkNAmaCEWzbpNQ2xi
ynLWZzWe0QWXeWhRLblhJJfvyWJwmEMqUUIiWTT85XHHRSqnBLP2K47Wn+pUhqRT44ot4tB9/o0a
uQifeeXdXFA7QJmrKfjJnnyO8vfJgbCjuWGmdEHPHbsn/MJaontclkTZiJoQxEvLfY9QhBflo5j9
aMLtAkhcRaO0T7iT2S9Z0wT9JCJleFIL3YSpuCIaoc/kVKdb8wvEzpCD9oDLpONXj8AjpHAHkMof
DPxSrWqaDSNJ43B+Adl50XXUie3sGaB2HCNsW4CCVzK7hyVWvUznt+ICpsEjBy1lueATWba5TzOM
cYoYCyxJOsQHkGuN78Toge5HHjp4T9elYI8VS4tR/Pa6IPF9bYidwZVETTST0VWFp8yXMjQOB1W+
3WA+n7sRrQIbGiOhU1tFCAKYuhObRO06oMVbN7JOKXcJgGytSCK0fsUUEkpORcJW0Y27zuz5QTY5
IfwlOrt1DOcWNMdWfNGZQl7WaeWKCZVElKF3PdymhhzC4f1IWDTEm9g6Y4ALEG8p15JuMI8HDWj0
mXXcOM63e8F109dnwGXEJLBchb3JzzwpxhO5KNirIBnEc3u/+J8V1Nji6niqfGd9xw++hf1qsih8
qvOElLSws7XsMopZmo8+Af8Yr9Y0PURCpu39rI6I1+YZlQ0k5dZlVggLs0rSj5J7u7oTO8NhiBaf
vwiXED1FfZ8OYC45dXfBx86rfg+MDrqWYBzGIfkU6w3Sn4qzdHuvknA8xHNzuNX8dTlah2drYrMU
g9/WtXkT2h8R8pBNJm/93DNknIVrYKrBEZjTxQrt/g9ps6XxlGXLwbaPjvRjGWntryrvWoQridDa
KnCk7Uu16RuTiQwzhYb+/5URaGZo34C4dKChAb5PMl4cF4OAQr5/67dMj1ZtDB5WnyLDPAkUyMDp
QR/gGItZ2CoiG7LJq+463Q86JycjVXnpWVCg6KZjG8tNGlbalGaMCYB5K0gefKPHLaEzx11aumlx
x2Yvrjc40vnJg/3e8H07Y8MXpJVaqo4y8f0AXCNmKyBtXAkGQTotivCLQTJ4u3sJZbOHlqgNcbTT
YExBhdRsVx4RmKNV1kT8T5ramZgImQ+EQMq6P+d1jy6f+dW/CJInZi4+x2SbmPtHlSHgGl+1z6Up
207yALjJX6GaEpLSu/g59kybiINXsmc6+noJkWBudAqONuudwejFlW+cDKz36x2hX3QwuYnU84U2
q9mmOnHwDlRJWO+0fa6N5u0CpdDd7tHMFTjs9LdWCVkApcsDkSMXBC/AZx1XVi0CyAlhWK+KaBXA
k7LKpCo2Nm5ZGpV1JabIrQxcmxh7lUIJPl4CCZtdAHbPzh/P/+7cem17Qf/WYISi7jNCFScgKJuT
Q0N5lVYOY8MiptD10QuFPyl7nj4Dp8K4Cb8t9n0jgQvXUdEBcY2MjOY25p0i7TQKxrzJPXLuA7KW
+mGh/XL5WwCmjFE1FGLD4EBVYLnWMfG/DPlxnv5Aajifkp95R83+a+SzpoIcda9ZVqbThxUWsU2O
1XE5lrVFbIko+SOA5PfqSYH4pf9YyhjZpoHiKUnSNh6/Q9/5wM4LsztvwIoive2ZYSJdzGR5vRHA
yGznJLcQHILNdqieKkmS5tn4RVrnpLTnYVSfpjC7o16MS3XfBW5zTXfsTJD/yJxqMGhlD46Hu6J+
5VKk3I645pviFHEWqQJgnA+eHg/roL/Y7mQzUkyo1WEipllEUfw/FQW63Kz1PQ5Tbe06T7gQ6zko
hirqxkgkBixONoo5HRT9fH2KGXUFp60NzoHRBjaQktmkFUpXggBfVePSRzfVh2hZLHCcho1+eudJ
JfarZTWM3VFGVcVwO8HRJJG4lH1Dc54EiAafZi70RlXGT5e5VoVas7UL3LmjVkTWvoVOjuxSC2JB
fJSHerSM2ZNlbralUvGnIwo47gJoVJoiFREgO3FYf1EAFdfXDvulcUOzGOpZ2fXl/s4xudoAzQ/2
VaHLi+uL66Tq9JWQil57/KKbntVM066VMzeV37AWxMWjcbNSxfiYuBbUUPIykX1S9SUIzmuUEMUs
0W7tvGOh1cE1cfp18xu+DLFU8XhAOLABWbSunwv1Zp7C/ywLVcAB7IpmSmfMJwi5UEebZF975XJW
ZkYOLUwo++Y5s15L5IZ0exAsRGBNdI+f8fOtS4jr66nDax3R1Da09ia0gmR2y3YWWUlMjXtsLHq4
9cdaXlnXaaVsD4Giw4ss90LU6uCwUoUgcDDjY9hzCp6SrX3xWdp2r1lg1L/yFLy/IKVDjbGoRW8o
q1lPRv2bd+MHzKOPzbX92/fpDVYeEtWF6DcVFg0K6a/65LjKnh4V/cKNH7eLptr86fJI0OlI1O0F
REjTOvzl6U1rWlTRdX5cqrN/rjt/y76jokXuoonzf9A4Rz6u9gMrNK6GcRUHWiFHLj3sJpGXXLsn
r6zb7IyLw6rQOkluLUH6aqRee6EHqQR7WDi8Tv3OtmEQUcjT8Pj9Qot0/ldJ0wM8fO7Rgi4gHQ3x
PKbkmQ6kZC3iF/tlAb2s/kxuZRShTUJdACx2s74WX5atKlkpq8xc0lOY6HazzDE3H2B2wEb1sJM7
rJ4Ltx4XpXqs2HvYIEys93DLM2OdZqpOQ4n4KlKw77JUvwtVUuXj94+If2n776RG0tHL56jYjNYc
zPlNTpMFt6CNwBDzFiH/D0vF5OvIsApGVMDIz+8xPed+FD+Bq2X4loo3h8duEk53IX55xJgfzZ/g
hMFUyk/t8Mar/8jjEXwba9yCcl6GxdtFahc735EnufMSduZK59JGuENsoicaNs2R+V70ICRMJD9J
MgZRo0sE8b+Qokg5y7jqjvB7lRWm3ADUYeCwGlR76KYaIr9VcuzQBgwaDU5RaqvqV47BxOeFIk4t
W27NhzXwDZ6nibCucLldeh2/5gnFYmid5nzy+fd2JNkwdM9B7LAGy1CxlcBtslHf05Fmyflz2ZvA
q15ytHyUMveoaqh4OiqwYKc+NroYda+rFuVpsd3EFTUG9Tupm2VLy9w2an4DLjzibaCArSAyesMw
UwYYI53ysh6WNe7W8TajeAELe74oiAUxG5qExxjvHJRsYdMp7ErftjqWz8zrSCelaHZOl3Byu2+V
1HVD468Lc4g3dzSQIdvt4xSxqkXFp7jLaKxX68qFNksiaX9VAq/RH8J9bMMnfdSBt1IH9Xf82VkQ
NSLcxXWZpAnR+zSFvOwwyc73aHa2Uf4jFonKkDB2+S9iBB+S0yOVqbqDNwKml9VYY/7J0XhIgf8l
hQuk7Fsjj+M4dYomvGqwXjE3rl8gdnHvhG2NcavBtGEYl2xVn7EhKJX0mYq4OmUR2mzspVd7JBlG
fWUJxvK5DE2imSsptNG81GwQyAuM3S4TmsKZZF8BX7vuD7j1w70q089i0Y1tbI6PebanAYSttoK2
Ao618Ec/cwo2SRsLWsMCoGtwaKOEMQ7tgoSBWnyJIqcM581N4sogv8gXPQxYV8KjsngTT/TFD1Di
4D55tpc1ovJwk/y8FyVhk+uEsKuhukU39geyDRVmxu4XhBqXRDoIey2aDbJ+4OfrW3D2DX9CXGTF
Ni+/iFLHkHxZEK57Iu1TJMV97x9yNfeapcX7Vn9Oy76mrnTq823k9F3/JPLa+fIfHuxpPFlpiTPH
fauNzBPyx1/CU4+KK6w2K3vCogIRtTBndXK/iCbSMOXyAzE5V50Io9Gplq+EO5TUomeQ37S6P0wN
95bxDZ/kX0+m77Dsu6EjV7xsn6CCONEP7bychicbTzU2QIKoT97jzFm8+hJAswlVR0t07P6ZLmGG
KK9DypuO2+aSnWid/vDN6HMvWoMVVvmgSsJ/cpRLyJFDtgncvoDbuTsr7jfqWTjb9s8U57x0F4Ja
f/jrf20pwPuFEyqaIuTY0vbfUfXZXUEL5WgfDeogzjuIBHcxrLbE2+Nc1o6ABFH0HF1SCUJbb+Og
r9av+bP2SU27BuXSYQIJF863E1kvhAmmkLGiybUz8ia6R+J9OtZcFhByxh3RA8cMtxlljKSPTLaf
CrWikaEN+2HVP5b3KX/VAKplSr+rs6hW0v4XpbmO81u9i0gtmfqPyjjy4CPp+g+8hEJSQa+BBgN/
6tq8mW0O7Sxs/SvkTOaZNxH+yR6FVhSpeJg2y02WvjNTBMVIn3l0rr5/iZnoVUSDEvceLHV74uTz
pSoZcuvpRzu64EPWADgnW48ajtxAf6lERT0z9EFMgJpRlbmBTMXgy+VljfS8n5sO3IotuWv2lomX
HDZ+E448dTXrmMj969JEiKZNByt1e3mli3IXUvKsc4Mq29QeN4B06xu2rSi8sVc+ZOa1ZoxEqSOd
v1lxWzur1MvNnGls7Rsy8kBUiOBX2HbDN2QhROBNKq38izNiXsvfXJkiwYMewuLEGTHkRXmRSG03
mQrbm8XUPRxMijU8tL9GpfxHl/MMOtz8c0eRmTwuIMXYSRPLjkKmLohzxlwjP0ATrCLfNL7w5kb7
BjaSg/m7XsV3uA++DV+nPfLMlOFGAfpb09bFyI/jR+KUxHK7YSOl67aiim2d0Y/6ktlAIv854wse
MU/qCqgwbAtnJNVxJvN6BxB96fSnL54A9MPCxdreumUjb9qcNFNpIlAk3RvCDdQ4GJ9yM/5Bl7GO
orEqQ0TaYW4r7ItZxDYsa86Yi+pK3G7beew7o6htPEDb1r2TrB2XKfRu4EnYJaiZG12ekAGig503
ZmFuLckEY9CBNiTkkMA2wVDQ6kOw9FprpzMEPinleZ6cfNsOTMuigHGjGqv6GEiEOOXUrOu9Fm16
6/TrZPF7fei6PEEwvL1KuRVY5XNscP2LJaas799uw965qnPJ5b9GkFxIruHKXglnaeSbSQpzlQp8
zoDFtgo/N52R/6WdtccxrEZcyKA2scwlsONQ/8N8PbcSFM1U8JwIxL+60ZfZZ6zB8Am+BuEiGNXh
02TkNNZ8aQdCQm4yabLC7g1KTf2fEUJsaRsiujoJox5BK8FgGbZHZVQp6Jey+P3suFCee4H2Hz7j
rNeiuybObiffTBSkh3cQ9w0N65qUEZU/gjEIXqVZcGgimdi2fe9D7YnitiesnsztIbFepn7sRH9f
wJUTn4WoZcsxsfqHFxrX1YoIdFodxQuCWmGERt6KJvNZ7j0MZeVpyO8kHOQQYnmGyU/kemq6SWXg
w5zHKZdfMu5oO+hzeH3VuEZDWXQ298h1aAw4LD/+9crrXuwG1FFduHV9rkBIXVYVH3Sg36YHxZ1Y
7HaGByoRGBkaOUTzPd1GEtqigCaGEabO3wQimZf7Ozr6Ri64HuQcAYibmie2lPQK12Y9Lo0HLvCw
paluGpTSy2lKFrFul4jNL9xb7sxDmnak7obONzCwqjRehLeORgynRVGEJWwkrFJkbZM9pwkGSxiv
ftzjJf5b7XJ+XQ3wx/cms7ct6zpwFpwSw3ATdMQR3QgVrnNvrSiJL64lNGKRj4xg6md90bJMSve7
flg3TzkwMfTispPiE1v3+mV352yeurL/W8ml1LRHnyF4YcORKRqddF1/5aM5ikBwm99u1UI7weAt
6p79p++yvn+Hn3+Q/QztJo2M3brPngk/xNYtWPBYG4IsA4p98zlF3IGVumaS/IWEreAd0qWmwrII
PNP7qXGY/skcpSXWoeFMe/4GKJDwCJXmfh7pDGIvLD6HdXkvobVj12LWfxGFqxj78JJpZuo1te8w
ZH6dzSTLSjvpucU6uJY0PaQQXCzA4O/rxJw4421V1oWhIM1JqGCZNxLy7ABkJFxYmFJhAwC9fDEe
D42dFQnbPWsbuXnlye3PS6gLGATrsjed2ENtfqz25y3KFgvtbd2cv41kg/N894Oc26q4hYDJ55xN
HpA3wg3Z36symfmD7XXIhFgXrh17kdbNb820uOzKYrFHQKgmKQ3gvFfheGStdaDk0ubDnIzgnhFU
Ws2tn0U643HtQblcPywLJN4qSmLZCcaR/0+Ndjs/lCL2Mh/UKtRF2HsBJsosBZlKkAVZ1HyPPrMx
Ds6ubc2y9hDdOPxHQ8aWsS0wV/ViTUoQF22ZchSK9gNvNUg8PvcIYF8MnxM6G7C+uZWdPySRQ7QG
hMa3zfCcD5omErmfUVDaqOll77HUydv30tAwAxnliWH3kMn838bV192SGhvIzMAlvm7uRAeKOLHh
WTEvfG5mf1+/vfiey7+Is4u1o71PJB0vd1FJK47g0f/Zhq9mdB84O36bDUpZIClTGPhbBBPQf/hU
7tYrEH6uihpKn6rY76z47BVhpAOLI/vEnTAx+bTzzapOPrfGLcxACs9CrC2ex0gXN8oBeUjI+Qn8
glXLsht1/MZ/wnQTMz8pdAkE2tkhsm7T3JlVgIPMJtlbYAVn39TRrCEvNpqGEVuLG9yrLX7TJoZI
0HMeutbwPzHg2XJjdSpw3b8bScamLCG0ZythkF4s0NfR8QeLjZ9mSigotDLXPy2vxNCy7oUnu1hK
5HJCy7xwro3fKM9vBBTlS1/eflgdQ0JTt02vMFYh7Bh501PUofZ7ECIczznrh33YXQgF92Du+W2R
NfPVMpx+pITRVwbH4GGn/49DclgdBF1YKt/AIFG1FtW+rMThuXKC3+tn7duR6g17bJHY99szUWo+
K7lAKwWmj4lRmGVI9NugGKztwpK758H6yED9yPvMp88Wyt+BH7G+muF0Hr4PVJYWGPccWmAEkEr6
xN0TBhKwpiXkkB+jySpQXjf/1vbnHWJS45Vc2pea+qSYpc1UDiWWEutcKRVGvLQoRRkWvCZEIzec
t+pg8q6DwwLWdIQYjeLmclOOCcUg5kkVmXrp4eL2WY10C9rCg+w58Q6ymK4H+6A26GaxZdU9hZj0
3r/kAnvsMMK4YoLLru2WdWZHLiK8rrbIcPg7dd4wYY+QWES/DBicZdykOnv4KwAHZAUo667/Qc/Q
ThU1oV2OOEqK4EDyXIAW3z0d97X20FS3PoAH6nOc7Qkc3omE+dn9K08I4MFSb3etozUC9q/Tz+x4
hxLQIxfS3ZcxiFZn3qW8jy4viHlSq0cPIxcn19rX7qdx1aLkBhmE6uZCbRsIZ26T6zKXUp4ZPcJl
hl0cTKF5eAAThyYvhKP82zBS5/6jS3rYTIJKke9sHuuPlosY3VU4XfrroznndwTDbEYEQ2qICeDV
ERNn1ut8HTrZ2y0WpAvOQ6Np68IiyX680vailS60CW2RQLTsYScLFzngc7/GUAqjwLrNu1nX98mK
Q129jPrtvNalVRa/ezy6Tqz0zvoNmuuxsLxGxFzPNEIVkbTjn+CsLEHYfMfZJvuDqS/i/wqvo0DX
5y+oTpOMxr01BZxEhRl3Cl2xbsO7EXiAZKeTeB8tgdIzISymUO8fhAVUnAmb51gM5EKZXLIGo/5Y
9kV03ZbinFCvXaqA2bpmGkG3dpz7k9xsTFuFobodotHnXjFJmhUy3lJdCFTpXOaOIQqKEeGNDA7u
dJBkhscd88cKprrUQSbwLsfyByZJIOqzvP+BcvUIkgKlwFTPlOaM8mki6vxoeXd6uNFSycGM3SoG
7wh9b89GrVtomcDfwDbcPf95NEZ2NeQx9Xt2p7aMPVPy3/Pc+bugXeMfXJwBpjWqOzAcw77WbE9k
IJ890CuY/PYKmmxkKdZvXEoxLvY0lGFe0j4KzfkbJMReqUlLgRMJ1oTjtzKR+XCJCMMYXZXg2Yoi
Rs2c2Q1cW6nDq2TFDAQdjAdR1zHy4aK7IyBC3w2MtVMOb0+bhwyfm/IwfOx2WqXvPPMaJXyIWasb
rNOaZIm4ZfylcCcRt/gDh+S4u+YugNTIccxMVEr99Dv24oWblFqPgPW7A6GhLNANtV2OoVOGNqEX
J1NhQYxr9Ru8t2+c9R3DwX/RxsWIA0N68tg9QFNBCbG3h6ZQny8GIvpeImb+k/jW0ti1foWFN9Ee
yHfyQwwOrHPV5qGyFQd1l+AmRtD4O20oDc5FOqwZD9oS0FdWlScpL/otGRjnyqgyVeb7j6Ev0VGG
3idRPpcfZ/r1co55zZ1h21kHRpa1brW6PgnrtgYNxjdSnZaPqgv+KFooJ3LgP4216Btp3Lo332Oa
ZkWKabzbmrGtAmNil6ylV0MsmVSu7f5dv6npiBijUaW2Ue5A+76uXfA4rkYLTAGcKXV+uOU2GLKO
ZWuTALAwZYwcwgekZxqVlDMyGgV9Il16KIp0DC0YcA6vFRahMjhdhm4VXSmTwhuAf72gEIaYhWJ/
2k6n2AX76Uk5Np4bU+8ykBnUveaUS3SFXBOhD0oV3ZP6kE8rWIJr537zECG2Vxz4COMNcKYP+oW+
0EBHYbKWAezNV6drSpYp77wOJV17kou5zFXG90/sqzFEqpU7HYORs5OZDgs76hHUPYWLtkF5gz2r
JblF6oz51i5NJKWq03v6VVbYT6b+FIzuT5o40zWuVP90WxeDdXbVZ+pIagD3k0NEBvIY+X7nxB6j
x2KPTJ9lWK5lBwSHfiimpL5SUulTM6cndviLrYMSIDXkRB2jcdIgupDDblssn0XEjPaE4uNPvCF9
FIiHiz7QUwRhnEyNcI3zffhh2eLmXqdOrZvwXVECVkUa7L55cTfJhzjzKluSq2EPrgbCyuouwD2r
ivfhHPQOunjTbHkZMxCib2ZUHZgr3Zhkjc/IagorQ6qcX5FUutj1Gko9IAVei0VSy0hpeyQ0tlgK
Ly0NUHwby9WnS2tX72NQrzOj4/DHZugUD2Gk4W0xoenEYRtkZRX1mSNggsfSpTC97rRRbraguHMi
C3DKIeV4w2hLPh7EsjobDsBIhkLN8ZMJjPVqtOItCO5V14sYltjhwXWo5aP+OVd13+4j+Nml30Fc
T5xCZ1hy6/Lt5X71Kc/RWNYDbwYP0xLBON65RBpj/vSaOnxo+db8uVuR5VV68Oo41fHsA7aU2vq6
HgbYiZ5USNRgJZ7oEmqjDBb4n6DqLR9NCfSVdICCykm5qKCV2mkxgmJRI6n/xMy6YQqX18zgBq4Q
vBoQCTjgmbl3BxE+Vc9wwm8tnsCryssRlXEDrWxw7I0ZMnexs7QN4cOfV1OYGDwX/mFzBa8/kJQR
dqZtqAs8niAeSf8pkVTZmHoTxD42YBmJAdlG5/ICX4pd8TouHkgh3M1yAnb30r8/E+bAARpqW4/L
OzTG4nc4lIvM57OMMxJmCbaPC2JU5gjLr31sNgT5Q+zw1/0NP8C1d4IMkhYyylLCLmqdSslY8Y3V
I7GXG+umQhQeYmwMnsi2Hw2hxIJk7NKXr9YIQc+QJSiytkTPmSdBoOjkTvmGXZM5U2+e1KjK2Qf0
9rtUkgaBsOJ25bdIXulaHEFZOpPN6dGSXY38zX6cDgCm9BrLuTyvGsSwTVbrkgdIZC+y0m49+2EG
eIWwmqb23bSnydZ8VegjTtbxQmJNKXubNiySbAxkkTP8fzuB8F/two9Qo66tncp8JEgqjIhFVZVa
XAm0kgOg/B8Alo531Fx4vnlGpjjTwAAlL7xjXWbzbcthvTrRxSDBe7HxOQK2l2SmhdQWQYXjNZ2L
Xmddb6dZ6jHnmXxvdktQZHlqQLoOPtLiUxWyErTFZbEj5WdFbU8KAs0JMdKsYky64ri0I1ecAeei
fJZ1LKP5HbIdj5X6/jT3725y1/uhKrmD5l7zUFHk/R7sAotKFSv7kC0NcJtRZ8OUhwyg/f/eJBo1
e0xLGMWyhy19BfUStkurAWHm5EYkwxpionChsCRjsOs9k1wQZiFOIiepBfnFD3WpK1Nl/8/+uzob
Qb/Vlg+JSQNsqIlXeteu+BrL+bCew63Brk8MyzCJxrEqzrsaRPsDageW7txvnGAgPahLKSAvREGm
h+1taytNn/k9BghHF7dQl8wXQIeSogx+13Phf7IebHI/d26eoZ9TOXG6Eh9txx4BTrI1BGisTP1x
ucigUGsJsX7DALl+/eslwTYnz0cm+J7B8wnuuE8TLRiGHUPOOi+IMBEugc0AIyrCIGXELxcGl6KR
N2xgOm2j1iv0h5ROdo93U9aSWYgFXM9Y3suzxJ1JC+7N5pdWgyLgRAV+BzbdmxWVwCewABkM54T+
CLyLqOrRUDE8Omqh2wTHLtjyAroAemqquznxF/IB7VclANFG7LHhRVDDaRS2OdKsqhQAKLXr69GB
bHyI/y4VLFL6nAbIMhpP+uiH9eZSATbEBAQ2mHje5RZEurlLXZx+cdtyFL1LRJQgnwMx/CIQwCIm
P+8oLTr8eqLl4a7YXmoXPjh8GykjbYI5M3Xl8zwjGc//Al1sALsrXqnXUYASUzeJkzj/r4hJohHx
CjC+09LLrpaVnYqH/IuNvqCjPa4sSDq7gsiABw+sNQPCph9GOrawbPJ83kLxVxtC81d5JvvZV+mZ
AJzBbxkO9f8WXVihFZ/5jXYCh7wcLPuRZ7foC9cBP9fXsMlLrww91S6Tesixu6bB8ohR4RylADoA
Sqodgk7X5MIPcfK0oGyx2upOOpCSmstAoev7AMO/naVBmQ4wdR+8vIDB/sPlpziSXxm2fK3U+oFV
ySzwnVGxFhamYzl4pCqExSrUvd8OEUKlwHIF/X6O3d8JTVb5aza1YffA8qSZX2aQF+deBsFjc7/Y
pBNeb7UGi8gJmADev6EabY17OYl8Sw0RkB1LPsHKJ8q2guFxrlhbRQevwqhAOAY6X0zov2zxZvpf
0VaI/yNbxNPlBcJf4fywIktrcwbPGbqa3W9Sdy6v6mUeMSd14QwyntP+2pKePLQuntsqP7+io73Y
d52fq61eBx3RQnmlZo5op23NbZruiZrUC55H1ACkD3jtJcNOuVzbTxUNmw51hMNSLboGKIZXSZCY
wW39hteyL5rtE6Cu5pTCXq7i9W8ZkHeIdyR88yDQuNrbzwpLsWukhZuG7z2iUDN47kxxw6cIbu73
b5NLq9Ui97kdSJ9OQ0wqMdfnUwYB5oseoYBxHCu/6CWJW7HqP1ARdeWdm4+ymGq3cG1nAWBBsqQE
O8j+SomieLCTY/BIMF4JXt6Y05G+J5HIxP3DCJRCUpSQdjoG8DSGRI0x2cvbD3iB/o8gQB1Vb2/d
FfPe7OPwqNzV0d9isY/S+OK/7rV8yLPwtTkokZWlD6zwJ8fRVneG+JZPVShVPg2tGpHM7Wu4wY6z
nNzJ4FcM1XBz5cNy8KTz9u2fVps10jQOyLjtEACCJncriwBpRyvfZA8lFWTDSyO4fGJavxroEJBT
7/lPlYoWsuxkLyHdKMfIcQ8g4cUau5BS9ehvjOXgr5ob2BklrkYTudGSI7C1MzMhAAxrDbuiiMK9
X3eybHcy/pyoBE1KRdeZQbDtySC7r5WNkcV3mIiCF5G7La01FTWgjxoOZg9pNu8+pGK/7nO00WPl
RD3I0lchN45tt2wTsBU73/RAO6dexP4s9iZ5oVF5lD94OZBlyHrQZH90I5Y8Omd5EDelz9ByV3mv
xZKY8NEqTYkCFfVEVn4I1/BMD+wFolfAX351h6FcWv7LuAoxMUFzJXKUQ1y93xaXbkVhLNlll8j4
nbXOIF5Ltnt9/7WM//EEKRVgk9srKTSEindsLyHkpT2MmGq04bnRchKkQugxqUfQE7l3ZXgW3cn8
/GFLt2ZXcV+xpDyX1cPFsBttK+GA+3BzM66vZaI/uWucxTlU37YAl4Zjohsqz+s1r+9o3A856+nQ
0ExZX3LeXf67cYjklVhieV8lZayPdgAJn8XqlFSC/+U8bTcPKKK0xEW2yhNaxZKcKCLPZqixVkMG
Qf1EkMb/hyemZXqwaVZMIXP96NkXI4Xb7R7iHaZov5joXefY2IsyT0mab2aPIW9/FEUOop4kwLTe
3bhOVqClByw3vumT85B6MZkNGTSrU6Qcp02QLwBdtEts2g+GBne7ttj2x7/5tz0s+SjfVL3Gv5xM
H/8ZnkvWUiFULycWMm+Y9uO0ONF9oGf8ptRCW6c2TNIOoZD8GAkNMi07VJvcp14VnoOMixG88gqw
X4eUleS2w4EnrfJYPp1Xbk6fvrIanAEw416bpog9rt/cbNsQCZ7IxpU6OHoAqwaLXSAKmRxsLrFc
rFTa0EUEmtPIHM4lSP+9+2YpaFy+JoS7aZQFJexVmvRJnqGiS9hhLE7ME5JjkxN2yyJJm15kG5lM
6yEErKKytvMGbwxWkob6wJ2rl7scFT2FJjV3aILY0HO5twYaaAY19su9dZgdOrYyztMUKjrenZiU
1dUiUF+kSvg0t/qDPC+RbNipT08QXS6ibzKICL85khZvxONOIrDQtpaxnF+2uRsbGgzfKSsXXvab
pqtihnyI5KIkz37wKr3GqrhAOVZnDfhfvIvVLQ5hysr3QMcW3h5voSbOMSYUghuCWPXzk2yPcQ56
kuSG9Y3pH2GpG4wQttKe53mxunkoErNzwscGso5lNWK1HNX+0bbThYNU+HF73STzq8p93B/A1RnX
oY8T1Jfu56I5dWz9Kd0hQM4kEpg3FC9TUBpuvbA7ToC3Au4BeiKFFmkN+aXaTJYHXFUBvK2bVfp5
ChSrQchiBaG88DVg9SX52HbV+zkOSCjqS6YATKWYjNUApr+XxZlpPn8zj3ywOxOzb1qLfdbLkVjV
LAmWqxodTY8TZF0K4oQOmKHJAoI6DhEu2mN121eFmR12q6+0U8p5o1OGpnN19YvJuIB5y6KQilcu
qAIFiO/vb1dJdRE7tlYXEY2fX6GpYyg/D0EFtiT1UwD5JrUgCW3XQvvQVuZjDw+j1iqoUDatz0N+
QWVm1SX/PCSwOu6cqGwa1IxAQ4VGouPru3KAAShiAubPhc8uhmM46fDSelmatEYMp9sRF13bwHKn
fqTAvBBXOyjfr0fWycWWEwqhEWtqYAn4xTntBzINIgfQLI57/4Oyl5CewpihlzxwU3EQk67dcDVr
gZZPIHGkdI1QXyu2Oz8rwuFD+kF/chaKh0ewHWGaY8UBvJYYv1LHByuxn5gOJEyMyIPlMBdwNWMx
mcrUkRXiq8CoKXejWcKgulMDqC5QQCE0iUVLFDyGesCb3Dip9sseG9VKucIAezp3I8ef+udKgNQL
CYPS7HGqlI6AqdrtnNcF5edORKxIv1Oj3L7qf2343lgArm46jaP808j3wlo1cHO4KOQltV3FvAfH
3uazZiBQbgdVV8jnqn/wQy7uWkwl2swuv2bxaCYILyjaqYEQ68lw6eP0zNeFGw0ILmlYGAAt08pA
C7Cl6V49Zf92XgeStf9VwG0WhbA+0zx8rcmrHn6u/f1lx4FPNcctl/Un5nlUDgKKPFm2rm11WEiY
w3b3oHIsFkUSuIdjsgGo0+lWhq8P8PPsA6Gk0wtuy0cMn2afBPSCjNbzCR9woUXBkn8IykGvRpAB
/vX69E3zbr6TepebQgLkGeXONMUhY5pcVHDlOp7CYzjy+ySpbu+l1ElaBvQBwVWDjIJBRPAxKMR1
GI2r0cmOW8s5PuoeFMr7PiysVxJX0VJT6d1B3y3HvDb1h/UouLtPAddfl2C/D9WLC065kEXfTvVJ
6xCX6hZtVM+j+nEveIQfnxyZD75r4F3qcrRr6Qfu/HWGeCJUXHXiCAY9amswf4wP2dfGcwd74q/A
byPmEkUef4X5f/M2UKJfwwnGFhEL150N/lW8u95/oQfra74x+7fAMtyoxV60zNipiPvZLkYM+0hz
T/I1u6u1B9H1hsD+pAY9WHvuBIhlelWQSwgcwpUcr2qOA6iOUNZLcKsZJGQkScDsEzMwXU2llYwy
ZkpdYka9rMG++3wOO410wJ6J05bwJxHjXGgU6RC8vFR/Tz4ORCvRbD/ViQQ+ej8+nlKdcDIR/zdD
ZX2sWqc4zy94ZoYyPqvGagRM7O4JmandO2+T9J2WiTBp4+sRW6/JrhSfhO7m74kpKGpnhaMDQhx4
DciPVL6j4PjAfej16ueaZ7spKuosDqd9b1RMybT6+LPfdQhlf6bjlrGxLjVXhi4k5eyCHu2ATqmx
1vhCNptCV2wat/tfL0PLvbLJ3KIiraxEV1XzYbEeHI5zV7IQznYr7L08pQcTTSF27A25lG0kTe3P
WvihhuTEdj/pS1ht7kvVqPdDT1fLWpU0gsWdlv5CUSBWAmO0+DjGcdMQ2ip/D2qvE5fSTCgy9KpK
i5SqYJXvORucDrGXuYz3TZhLarZTmAiV9pEmhzTRHw51moo9dazF60ZmudN6uEIY7g/m/bTYIL2G
VBglo68nF9Lq5v1nlqpGvQ1gw4bCUCmBmjU7j5dt+TJ9lFtTl3bJSivKenSO6UfOQTk6VWtToyob
AtlKeiyCWydfimZOY3qoXE5+CjkAqsimJBZt/CZ1Y6PJBcdCAVUQ797QWCDe+CoMTUb8mRUudhpW
UdPzD+St5qaTlfnuRD5BPokDDGKz1MWUIf49gbnTUEJ3ODiboidJJC71NLK6ypqMLAOaEKbak6tQ
N8kyJtRSYq+hbtBXk9VPm/I9Cw/cjvpPeAaX2DBllkZcnmXsGclU32AWSIdivBqvdwUw8PfyBZ/C
oeV6mdpZCDbR7K+k9uwXr/kQzIkr6JUEpVYuemT5K1kEo9+tHICM5pQ90xX5n+Hrr6PnUYvexdKe
uoIa6eBFQYMJi2lk8nuuUY/1rTl13jvEImWIJwHSgSIPKOoDgBVmprY5WwYC9rhrhVIYRiAsPIgs
eRrjB7scCI4q9c0rHRBrUvizTXh41yKcm8CQUxNOrEKw+J6LcnbwA1iWUtpty+H3A2kEPYFuapbb
0p+/RktHUmA3wPr16dYALKhStX464U+bv0aqNmmHrXS9NmmBF//q74vS91jl3iVyBwxwrE3awmZG
NynZUMdxbHsZno4btfFHatlJVFrw6S/crP8iLI3Bd6BlwO/ax5pgE6cfZe7NhWbPvXqDW185w/AY
7C25oFMOuGOtVxYOkqts7X5c+uC0QQ4+ccpEg4YZabYxuqBmII+qIFAcbrhyv0cHyP4MKiiz6u2z
6nzZAaCBU1muTlJGpyVf7AsnDGnIzv/TY0YNvEciGixZgBYM+stUKClQtwlUG62xlZ7ygCSJ+9zb
tQHYfMpmW7Zgx17b8MRKb5ZbpZp9pTOlEMGNrcpZ+meB0TOzcfCfgw7IXVVjJ3v0e3i1TFfvaCya
7ICqsbVihFt0JMNun5WhwvpH4BGQHnqB90tWrDqZbfRW0nYvNmbK274MGmBPk99UQQrU+ljV24G6
afFtmh1ZECQ4cUp6J9zYVAvwVInsp2SuW74ogBUiM/W54V/BIPXQX0/JRLlUB9fc2Flr3teYRcgJ
G4Tj8aWlJvK1t3tjxeGyl2U7oEfNj7DtZdpxmvUXvmA01tbAV7P3xU0Dzp9CCeInWEYUOj7178Zb
ut510KH4a6xJWqXDz1JdVWElV3KvxS85tmZGCPtDqgLeVpuyXJ2xaNQ2XkDlh2UNhcQOkQke9irz
i+UhuzWvBuh+oJhW1nWrGZDWBsJ5JUYSMecqDZO8JAluMU/SfAhk26PZuh6zSHudXizm4i+/YWx7
rSmEzY1wQt7pEfGpR1ZzxVBSeQWoR86TeR8bW89vO57Hvs9zWcZRKimOdyOi4DUVIXmYnV2LMJc5
0wDOsmf/U9tDXy/9OYLCZT0fcIxa9pz97oZMvd+/Fes77WKBFXLLmBLkp8ht+mIrxVgon+KCkv9h
hf/tQQAYcagQsln6t0N2/Bj18K7UAFcZnltZqCqp78ICueNW0Jp0Px40UftHD8qVIDXehSTcYOts
rEHwqC+p3crnxlpgRX6Mf4BP8hG13ffd2vbITrKzkmsuod7S4tpHNlgRqQmkJfd4oWz9eKdOvzuq
0oeTxKf7DJ1KOmExlVtCQhUMXfA5OyiIBcQuLfWjB9BVcb6LuJBKtEuZBxqdCGswAl8XptPbwhBL
MOWTyQ2dFZ2zY77T3DOQjuhE8TKhfruVA4THdCbRQHdynKOh2ru8yECeLc18OhAMmP5J5EuDH6f6
RtkHV04SuFifJ6xmHKN8qOaumySZOKZQp0s0kpYPI9xu5AmPYNg8+WPHwmdEU8QMcys4dgAGNSuh
dNX3jloLgJTa6Sgbb44qosLDdISRBKyR5gaAUi7EbDksEKCgT065RRTC+rnlqP6jeNt6oQeCJAxn
lIF1jL+qq9+N6GVbYHYUWFidQIJbnEOt9XviPAkeGeJZB6DmGm1WzjIiDES9B5by3uyr/zfIO5IY
fwru8AJ1pBeZmLFBGRrGLbVAYKh7pzjG3AbplHRlou4Kaa/kLgt05dddG6Tqvlej/Ci7whFKR78b
QyXXj/8PoX99UIcZHe50t5KfvDHvJqHEc/GS9oDA66eQwfgFF11HTDd6OIsRVXD7EsITCNyd7y9p
EClgOTy+zMFxp9NAiefVapdOveYd1FwkOn8eZ+zSuoeehTO4pa05RnhwrF0bKyTPxN/KMqrwaGDl
t+2HclDozoUj9+4Scl4vr9pUsQ2NxFbmhkE5JRtAgIh8Q/moHzV3ExnpshHYA6BaIayVF6cfdfiZ
lGlxJq927qqat9DkTsTSLegBaiAeGSctbIpev25ZlAiJezAHvdQxPr2W9mTRf314z1P5Ukaw9EKv
qTbR0yqmWsfcsrU7hHrK4x33kwNAV+fIvNKsNoyEHhhxRO1uYahBlLiFyWkhwlUpu3PrN+Z8hdFX
ltP8qVVqF/H1toIoYQW6I1lKGyFp+WdjG492FFiT4v4cVEDTQFHCbGOulPF808AjnRrxvyULQL7u
1oy76ACFrrAQl7gHvBWQngNN8cPONusIKJm3tgeqa4OCk8uBQbFfqrWOYQuimV+QESFxVximv+MD
HAQjqgDbnhflrBJ3vkVC7usQbit8hnK/xi0gvYAjP0iLqETsJXLcu/4URHrwc8GaOuPqeWJXgPIE
1rlcn4IUhATXhePrJb8Rj2Ucr+HkmQQDMRNTBZJfmOIbQeLYKxeRQYYjWceMy5GWbMUCyuCttuDT
H2zcnLUTZ9ZVWwT+tt0dT4LYbv65bqAQaNamJjDRPrzYq7WMZXG7jjOFSV+Sy7Ai4GLFFxbSlsMa
Mb8oEqTluv0hr2jEDj4T9VdNnL5NsrIKF4EKRP7xheqOhHZ5SQXf4n71lJbX9Wtt3QLGlZ2Jd38q
YpChc7gdRhhRjuffKParE5KHCC1KRoFi/kYKHml9PGCOc2iElXAXcdPrDXyuCt/t+saqzv10+JpO
TDmqIzby3r3mPxrwjyHozicVoS5FE7jAJ+JH0uGmR5qsUbZGzt67cvsRGTwSBPH2mcautTlHo4TI
0o07XPjEc7tQbd0ZwjHzHeC7LL2y5Ctc9mfI2sACTGMMnyGbPz+SuYs6/d1eTe/peuPduUrvS9h7
ovaDS/SGE65NqdjuBpsUMHw8WN2ooyQSHuANaxc/KjX/QXA7m0lmZCEld3XOU5RHml1zWc9N28F1
YAFTATH+FlDtdSzArffKii7iOHku7ynQAaOiIy8LLZxzaFLfpAgPytPN6/zuFcG/cerwzbjm9Fta
6/JlwWI7TcyFb2W81Oyq6XsWY4p1d8T8mteZbzKqwAGpCPCsfM/Gs9Hw1OJmBzc+xZ2D6jCfew3x
XpxRTqT/hQPs7z00cMnOmkcAqOW0cYUQ+AaTCebZi77sD2YkzgOhbI0D204bKL33i7tqnh54Tdlt
yYvZI/lr9/zHm1oRddfAZAim8Q+B8zUqkrHNkHoTGuUaOFPd+wZsZTSV4vsYLyiO3LMkHi8EiFC8
BUWwxkuliXguBzjYyYUopxAj527KY2Y9oxSXIknZ4S7NqkYKiVUqcX/rXdn7zX7Z/xsup/trkO8e
MA5UAVsavjp7mR6GDstkHcY8yjfqSwWt9SHYuXeKnMiErJDeFkfzXxI2zpqYj7ny0Uoh/b0EySfb
IpX78RF2oXBS8ijaqD4omwmJrFBJFYuoIhROMo4kEVMfT4gV3y+iyzhUWMf0aY4uHIOE4xflCM5V
/vl/TEU9xGAJM32fAM1H9MNgdVFTFSiDTzqDbEuI68nLPxwKm7aUvVlrBalJMROmgwrLNi3R0Pe0
0WsoRKbzAMCY0CkQmJo3gXAzf6sOMniFKeG4Ers8OVm+SHGSYn2RnUmkE5CiZGlwirki1clCvCr7
Xdy0Ihso+iyZY45E96mANeqWg8sAFMkdM6SXuSB7sY9D1L9oqouNAeF7PzCzgZvSyViqggxUTVjr
OWotDUBw9kkSkBUao0ZtFZBKHnD6fE+JTBUvvdumPgcxGdhiWqL0wiAsBcybUju3AbABAp6m0AvZ
/CjHlVFnQWIJUEzOYf2SRwio24fQk83Rii2MSQnwANe2AzWDVw8hU3+yXOzsCxTVKiiXWRNfqpCf
dx3HLQQmrpzsa36RLWg9Q6KY/DtsEY7/7YemTvXvmSn99j/4fb771qdcHxF0AG+3VmNYILjZ8k1r
tRfO0Zg62OsTX7NLKX2QapqftFIlUsNt8UdB3lwoOPJU4SqRw0s/l0UkmnWkgoBsUheia3Pqnw+E
yhfXwM1FvzEcoZRbwf395QmIwmVX0NiyqT6GzhmZrwVmkrtjitA2D+ut2t86nmXgLJ06IX2ta35s
55+BlUh3VeDV6ZS73HBMOTPwRyJPY2BD40Jm7ZlD+4DP1PUFvid9rMo9EKESqkfEjU1G5SlOOyLD
6Hi0rXmv5MQ9az04WDkDVEU1AWLL4jFO1cFn8Vcd4BAEy+2Zz7gQsKlIfbWzPdZOcn2MAC2CnIq3
CgdmMMhEMj1yOAC/3pXmXa4oNOglaX9RSUfkMqeACV6SaaHVZ3+ipUb3tvCLkQqx96JgkeIz/Hyn
HRUY3cry7C8ncBq7EhELKL9r6PzDv+z6AjM7NjhZfugCEfWz8fsSnASqHcs8QRxIgv2caHyQ/3OY
WDbNrVPh2PlYtLP5UJ9RMmvfzvYPPkkHusBQj3+tK/UJ3beB/rYr/4HIODb7OJ2MO07MK1jLnmnL
TiRkCBrnKbN6RY5m2adXWIsq2NBitxmoF9Nu3Rcn2GjRiUKa7xLq7sdsnRgsSLkPm5YTdAsH2VMr
MeWaY1KykVVmHL16CuefJPngJDny0j+IOj2KIU2SdRE+OE6+hs2Xkqp74YKr41sB3bGSlihtevm+
obYAOo2MOqe9salLcSvPPXKOb0A9LWRq4aPjVJaGhS7mgL/te13Wb57sWjyn7hCCnlSXudcUVOfz
Zirs26d0xmlEX6prIa0Y/qD3shE5GykaP1JHhiw0izh1scqnOsii+xex8npwpYDlhh9AwdLjbPnn
UdWv6vHuvA48b3sHdRcMbPuo2YEMu77p43GwRwm1bjteiFb5+qZWlK+9+HWaCESmOR3RbKdPLPSe
UNxgHZVMYsAcws7PKs86etwRwrmZ6C3CfoPUeaXrBL6uPSzkqZOR2dA2SheNSQXuXt9anDXuZDc0
shSGQcAYLzYPrUIYeU/lfSFgu9QMFVlA5fNmQp0fVdPNif/5ud2Kz5+jJhiCLV297ZtUbBQ9EGwF
SfmFL8P5suxXhyCFToOaF1diQG7/DvoSJ3uN3tMCMqTXMJh3kLxJGSrOVhYAeZOwQoqTaqCkuIft
PhkWsDZ9QGg5b/Xitn4gRq9Lq3BI9gjw9BoEbVVTbR3R1lCiP/hd6gupFHpw232dg+vFB+rHujeK
AElWGXOfD5Lvynxp0aMWrLf9k/qdgTtUHMNEXftNkatYhmuOty5+GDj9YvKaHKQhR4zmjXWbtQPT
eC2TyFJNHe9Y4EzRf32fM5hTE1pq50QnHIERg1lVI0HI7I6oQUlvdTOI3A7vneekxY8Xb92Go2a6
qK4xFg2eIFoKpeAvWO7Nn+bpsDOWXzZAQTQgnGtpCyCMgPx3OZEZpWJLBDbspUN4mBQxXj7G26dI
dISQGEkCAT5VGOXGwRFzL86bdV0XvlpQvwU/FBFg2enDZUjJ1riWNn3OUPEfb+GJCgb+l4ypFk4C
YTjnyxBiAAQY7LNQc+hL/9JpFtZczJN0+rccEeDFqrtfDUj1TgqRTQ1Jq5HXTBXtTeNuZveMsI4J
vqHD1WQgdMIG5YIXQ2joUm0CY+xKhASabdq4WqmfpdvogU3SAljmhQIznQ/U4j/SRXuTlh2e6J1y
lNSfnaTEa571QyP2rBHvw9JTbv+bY2Ad2ujN9N5Jiz+YPGHdS50+xAKLLGhhLL28Ft7dYgvijv2d
mDz60Fa8yLi1HzoyZGMNmbIJP81e+26XNatAWJGqXvxQR1wtoilHPebdfzXo36oFscNukuXRGtmI
qEeKFMlYCyGCP4KHlMVUIjRdpTSbaz7UKl9Gi28Vte07odDhg4y976O/YtXerQ4at/i2saCJrM6s
oRH95S8CMwfLvSrkW4EW4TUKqGjtkZ2IMi8s4gyoOf8NlfkvTtv1U42Wdc6eXMN9hrU/jnCDRSqI
4/EiriSdB1fJ0q9YKKDBwjtmdVBN5P8wJ2n/QYiqu5Jb2mnGXV2kSH+XSXHm3VudEYeEsnmMdNUL
XoQ8tWx6dP4ZD3XxAGtxPIZanf+htJRmSbRyS1gyj0781aWKN2jQA80k84jiFBR9GGPuVm2TLNQv
r5NMirrCAazwxnVF/AhtpC+ReNauDdTpK+/XI1cgmaWahHc/2lklafbTJ9BH9xRhnMvy2qP5pbVO
CUED6zjcssQDGuGSl4t1GPw3GBDkrziiZFzD7iH0Ung9a+BDB1sUOb5kSyqKd1CvQ9sC9midpaO3
s/Zemzfd9vKgYVIWXwQArjqlIrdnHqm27GkVl9bq2/iBCh7UYIOBnSYGC12aBfvgrv1hXzOFT+Ju
bT4XkDb58cie/PThlpCAe5qSnlsnPWJcG5uIC1gJhlzK8glynqFyfOQYKUxkYAwN+RVDTnwqE0iD
KpRb8r59xGo51D8vYbT330cTuPtc8HsqHCGc2RgKpj61m727YaoMdHW0nZddGPM440XkDllRYpxX
6Uj5sG61PuDOo9tZgff2wnmS6+SgZ9ERh9mbr0LOnYBz+4PhoYmvIK7XJJ26dPhIob0kzcyhvpZL
PqG1pk+RKKNDJj53BBUzqaFZp+Ztz3bMxjgiWFAf+LrUFe0DFH6ioqpt4g9gURts
`protect end_protected

