

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LQ2vJKYKktoZrCpK4juRqJANqbtQy3/ocOY3ZqWcaeltVJ85vibXAMA5tlVvS0pp5GAf58wutyGk
pEVV5Zv68g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oMuoQxHU8xamO4YIRqVhC5y86VVKXTIB4hGEIvLUCrdkutaN+fgAx1w1DFW4AV5UF4/dcrqjOzkY
K71n5sVp1APv9EcDNy4SK12rfM6JNEmec1W0js2v54algVfB410d4rZG0ryxf2jOEEtG3y1R1uZT
docKTvmf8ciwTam2vyk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RwKTb0xAeUUC/Zlh40ZbRUmoUjB02ejSjmyrw31uw3LFcwmpLfrEGeQFx9W8nBY5yWIBOz4idUaq
fc3pMxhJHFC7jCdnh3Y8hC14pp9rspO1hZLfCOxHKu7GOhZZlRDfFJE9YTYvNMQlQ719mBEfy5DV
yB6StZ3JnfaWR9muuKfjZivHmkGfCe6IBabrX2L7+LYnKKp4Bj89EkuYxLdjSsxwwHL5yBSzQWsD
f3NymUlojWqzg7COUuAovEX4Cr2S0yo+Zr9C4jJ43pknI50nQ+b7CaiUKqbCSj+K5CzuK/dZ/FYE
aO9kMeHqHP3vuIYIBhuz7gnYm8SB2OlUmalvFg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yN6ERKfUqtxcEaZPhTWcKmh6+v/ubkhs44a1yogYIxw8eK2NURIBs5ApjPyj6y69SFt7ufKFYnlE
zs+yxTyZOIDjE0iu1eOyuLmYVN1yfs8OFxlynJLngPXQyLVxs9254patixjWMGwWk4PkkE6mKJuY
ZOkdptcpF67u2/mYpXY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t5IcFW6UoqOUfYz1GOxoQECi+9Dv8vBS33YPIONcGWTXCbnB+Rky6dyYF4Y8M27ZqAdkRtAsKEP1
XbHsYeeN9tcVjnhsAEW+ZxZyVmGkxa8lAjUHEo6bSWwd4akFKgw3xIpbktgKgaV0fLwj4wfHvTcJ
XEKHWYqSYc/CYMdUUlUPXn3ng5DzustWIyUHmy7pVesXYKHPGiFba8n7HX/7Kf+2y3k3y0XUfQRM
e1vWugHsLB14SmtA740nmVJ5TRRb/gYA8FobWc86Rp4qtvRHvVvYBe1XopHUWeY1WEaPGutqYtgU
FjBA3NC9aJ03W8dZxVcVFZhyW8E1aSZwJp996w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1517888)
`protect data_block
XTqxHHcpmOLe3Oiu/cHyVlNT4d2hegBS8fhpBdXeRQTSYOsamtn5ReIH6xdslcyKOMd0otKk2wBk
ISUNI5fhZlnUgKZ3VB3yNMFOHCbQ/44GzLyxZZkASdmFkRG2ljSKUGUzyjc+7yejWMm5vxlzXBpd
2bVY4lcyLcqVVUAypoIU8JC/DTGFPAisol5pSgDFgXgLJ/qSKhSanNyYia0y9YWw6ocUtkm+TkzE
QZSYF+KJU6sf8YKeT8DLTk2D0K5zWK0vEXLY8v4vTPqX4m+W7ROJOTmG+fUPNsdz5wJIrIExxm17
0jyBOopOWGLcUMztVjl6gglpm1Xp9i/qNyunLTtCC26yC1IVMStjfTrigbcNQp5WRdDDMB3fMJMP
QV2IcBEEJMQbA0PmQtD+jsGENf6EQHF5AvI4HC9kiVCG5tjZdkfhYm6gUCme2sS4q1Rld7DDpOGP
pe8B5kV+qyS34YDjnBHFBbESAuzkKMES7ECTjJOUEB6+LK/PsKcPR8+at42k6T9rxdNdYqsO/Uvz
iJpjaEoyGyepzSmEDnn0LpJNh6zGVTob4tX1Ogn/j3F2O/lzv2u4R9YdrsCDA0bD4sp3jeuCFr+g
FIAgH5CQCKHL5MdUEUOm8sUIfWWXk3tN0mt0kS5+Wf5ROovsSdjdkRuOFz9X+GKqrkKmmRiGx7T1
dS+GWORmao02Mc41uIIp/dgdiyrb4s3ZnXRm9k5ERENEFxd210TK1E1yRgs6UXBhMkH+BkWZXDOz
eV9A71AfX49I51URPT9PvLV45L7OIuofJrZ7wGTOWw+cccPWZ/3L+6tjPm1tkp/2CV6Nx6C8laJ3
g473s0PqIULBwEaCXf9wuDLSdr3cf6VQXUJg+2JTIkvKG7LSeenxMfZvIoJ+PyaU6l/3Q5EmCXNh
gr/JF0qmixNTBfVNrMoEasFHpYv7AKpVvpk03zvb4tTWGjikAoMXY9tFEtnKmjBETO5xMlyEsnPh
kTMnP0vLMpEI6tYQhCdVztlssesN+sPpYBHQ+bMTPN9mRZbkF7ynm5UcpU5qvGNqPKTdMCYu1MHK
0m/brsUmSvFRk6Sh0+LaSflXjED80mlP9cutj83bgYNs/YIWcI5sDomR8EzCLkudPCA/9uo6Slx0
HdBT3KjmIn7EQjWsBc0LJFK159TSgBchpNZLl+qZTm4FWA5l3J1j5Ys7cONgTMBHgtUN4SlP8k+n
kzUF2o6LORKi3Rmh8syX/r6BEW8eu8yL0hkG/JPJS9hoionBWY1exX0JMtuAL78uzik2wpCwvfbC
K3ZM5yPNkM/t1g+ZUi+N4SwWkF3OKih0hzSkvTJ9K0Bk/ts40gRsHW0wnNbVNgzyZgQ1nMTJmBAy
RroDIhgvBbyQix6sEHxYu6wW+dD0QsrZRiO5bs29xoTYd/7akLsVyy8g2V+nla6dxuqWi3n27IUh
NcueSPAyt7ViDfLV02N0u+VPDqnPBQUr3w6u5HXDhdj5bNiZl5RXIAAbBrbLgHf2mXR7LKtngKxW
hwlgc7ehb6PnbKz37zabBH5QT8jD6Ol1JNCCfBNbloialKhgwLXbvKAdYZB3YQ8/C4p7GFvgMWde
Laet9PssRukxTSx0ikpuVLI0bgwdfymEQhj+TabFtyPMBxPSddMwc7fpwEPPsL2f7VYfVeoLQ0AJ
6R5Erepw0I+v0wB7yQHiY62Lx63Z7xKs9qt844Joi9JsPpeDrexxL8O4b1RiJCqQPbgjoSaro4Fc
YJPkvEGAgPBLLyRFfGd7MvQJqYTyPTNThCxfvkhsxli1ri39SP3uss9wVvj47SMTPNe64tn8sTc3
QdJCXX0XnhYKoBp/WF+s1Hf/tu0gKthZwMOqJEN/rV5x1nRNSfzSd5X5kpnNZ0TA+Hlt1SMjh4i4
7UG4wmJeoqc87vxE1vKlny1IS0uTRhuJwGLFBrKd9hEEMSBtw0qQBT1NuDMWDWOgozSKNuWlKpQh
KcrtsBwfyUh2tK5LwAUyrJZLOEvcOY4gtWod8KIDoYKMWb0E7NdpqE1XS6ydne67cdj+ZH31fKOK
L5ljB5A4pvPN2LUVdw17R2FVVctFFz11jBbGL0wcf4LK7I+NsFuUv4g0qXkHeCsWjteWZYP2VRhH
OhoUGGC5s2VRXacSa8yNBMIkDFjzltlG1sfz7CE69MVWArFZmWLNxmfxqq0UXT7UGpo2LS34MeWu
dd+NCLftR7lnBuvcTATSb8UXDUiGlO+vMasdKMzc8E8aUmy6rbrV3t/BLsZVcN8mu8pNy1l15VLK
EXU422jbNHhIoeLIhidMvnD7R+Vo+p84ZXrTStorIQE4/cuJgKpTtOm7eJC/r73q014VacPkSarp
rGvTRzC64ajGm6ztUVUtb5mNqgxmQCQCOAz0STZaW57izCeWJO5p4x02nR8GyXarD7wA2rCLF6p5
cLJ1lyTORV8/l6hKMl4DRVogWxQ0v1cRAblyqceQnDiww83HFDYEJETcA2u3JvNd1ZxC0cEnWZSQ
ctQkVAP9zOZGzTysu5Dfx8MSWhACZTn44zSYKsdDys+4zfEo88QKO+D79MYyusG8aPzdDB6sJj5f
ORl4ukFewn/u+D2TQUftZoWoEQvYRwm5WKMt+1HvDEju+vyuIB/+njHZN+P8wlec3lhc+gikfDlj
56DLgIKZXQJvHcMovRa0mkyKCCIr9LIRBPk2An8GzKRXF2KmpXEyoziBjJE33AJVUh4mSeDVx+Vo
juQAveoT5dpOWW6GVky7nktgFgNcnWJK4qEZwlXyTl4/QOKS/vSDaTqNqILGJwAafhOYtvylf706
7zu4NVwcuxYPTzrXN+wqHGp3Wr7Ki5bS6kYsWIln1Bj8sDBKx3rDVw3R6cp4ZITXRJWvyAnXfT1S
fGx1Qe0o4PzWaXojg+mQ3pdN1Am4AR+ajnwbJBfWj8bBpjYaAdUNcHVHJKgRw38UtzvIRnrZjk/d
Ofx4nr0d6KK9gbzhW2f+PtEUTRYa16Kk9zA8Z/oP4n543s2TvyX0o7w48GG1o3GM7va/1YdhqHYy
VZ9fB7gJW1Z7w/ChAinFa1y3E23i5S0ewRNWEmYIgcn7N6+RB+xRKEPlQYmiaaQQ+9Pg0gRLtY53
wFRhIzlR6zIZhZ10f0J6e5i4+owXfegMHooWfoCi+A3+1Rxf0igBM+nZOdXOGylvjVAITd1WY5k5
dT4xK1N92f9x8WnYB72b3ZpfIFM9nkp1LOoa0SvwWxNqLvCTxFpa1ci4ylerjDY2hsrT4/MSZ+wA
IKKOc4LfDunlviX0i3B4IKusS6bpJBXMWQX6dk5BRW0qzC9Hf4CfZzv3njrcJnsmJmyYQOgyjbMh
7LK4a83KHoCPUELjWcBjidXSQLlACumjHNj6uWZLsCsEvVwmuIqbGHcUc3qLgPaiNBt+ijKClTTP
Flg5WqFHZatuKngKQ0dmKlo0wA1z/Dk7d9QbWSOS9+WQ4XT7MGD6VNwgL5tTkpEisoB8mtCFXcKX
ga+8LibBdNAqhmO5OMm1tKh8fR/JRjF88HxZxqL1gKuHuhxRsXDpwVB/Z4IEjTVPORvEMNbRCYsj
j0ZTArWdudcJri5fNTMwx5WyMUolI7DmHwBe7P6uhzKzYDRAhyJ3e7KgWU5kzEXQgQQsSYX1ruRE
9gpIyiq4ooLVoEndPkqK3+OCwbKvKqD7hJr3SGIflHrg5I5kDr6hdT9H1Eq3f0NXeXcnlv5cKgaq
WYaGUuvfsB2pIm5KYE727ostHBL5NiSnnrLXU1tCF1/h7lkvZKu2gO8pZ3WmcigtwgRgG2lgqpqe
l5apWhsBAMH5QxSSxMqw2538bfIAaQlgfT+6I7qqMmramRPWerpkvgAJBucZnv1P6T3u3F6TlxSk
bzj8/RJ2I1ErDynaBufae7gDdmfWPAJntcQSLHiIFZ0Rqcr3Gd+mS60Xg3cFWv9nsw0Xr8GuE8+z
O5ddpg+GIFQzjP0h+5G1Qy0p9Q3+pi61QAhzXgmJ5VZwkWP8ssjeHMQwIIo9xrbp7/TPn8zpTwmc
8RaMFH8w4kcf0FhwS1eQ2bau4mWhCvnPnHX48rMHD+GFTL13sRcLHLLg8fYnXfXlVC8PQKMEe2Pa
tBzS1qqh88YTZU908rFGCiRxJIAgF2qn8F8i9xizpFHE7LjqXHggjPwylIMg3q3W1WuJZlPYwWDB
ZmzXNZ8prC+6o93lyoVjLzKaUovVbunTKtQ5RtXGvLK/Wf0mmPZHO5xarV9BlJf43WExnLkbR3Ml
NxEUSy1sI9KQWP4d2joMNgf5EgO+J1uk6T1RkruvTVauZwJx2e9IWHMCiGc1PjlylpPBA3XLiW0V
XRxRP+XUZoBNJcnEm4gn+8IMdRK1rjYX2vCoFg6EVLrxGksreEy/hOZKt0xooC2AQT8YWhrbVRDH
Uc/qzuPjXqapoSuXOZJOT2DJvQruvYF7k1oPY6NNWxrlzwTz9VhWhzsQmgAYGiutmYSu2ihH6qhv
kJ7su/lvjGPOazTsFdLCbLigDhyO1SfMTOhJj+A+OOsj57tUcTQKqmD+Bm+dXRytVwm79WuwcKqi
pn8XKeU4+RTcJdmI1b8FrbCka0kHaPfBlZ4kdjd7nP2u/EZ9OMfCjlutiF9ANJlhjovWrESqdupu
orafbYedrVBqZpeFARxHHOMpf2DBq5N1Uh3cLM9IHa4F7yW2o9fG4UJ9b5LevlUQfqgMVMLYoKlA
NzfGfPsc3SoFf2066g+GYycyjcHMK3cuOxJE7y3VfCcpOse6xNN5wCk7sh2AddljqZ8xC2IC+sbs
4IPcEdB93jxDX3+uIWtnXGTvM5++PPacLNfce1ZfKP6mcwyqeoHVoG+9XYO8tuyb8ejHvNjU/hcG
3I0q5XyFxey3iR4JqVzdRQ553obVAVAec2sVBExaPUcwglbXOQfEu7mgn6Mggn5GlozXOGkNTh+B
+qB0mT3rltvn0Xlgn0nUxxvb7TY8l0hbVqmsbg+w84k1NV6niFoZvCEGs6I76o1462uB5yD6MgyO
9gffdTeqWKL29C1E7Vqq/HOc8LiVXfPBb9PixTTEdPeQ0TB+Y5ZnRPjJTsRp14LPECI1p55eyS7h
23gJJC0R8gDGHY+t+OMrEFyEPBRo/qt6eHDB+1mHud4y2Dy0uMBXgu9b+D5Zd5YbgmoB7EH1HAAV
K9TYeTgDdCp/7CEjl1GHcgLXRvKrGY1AJh/36Gaohuod2WYcq9DjiBDy1tdpFiqCRV2zzmKAUf23
CALXnPlAtXpSJVYr3Ct6BhQkO3ZGzuR1tuzsc+1QrtQ+6+mxq9/uo5NYPcLfNwWlauj3jnCWTT/V
QVMjbJyIu9NHxl/QWWAOJVE9IVe1PJ6R9hwxC/JOvh4mNGNiYfZV2a3+MK/Q0VULLo7hKwHZC7HY
xC63YZHKPeM6Hx1XEOt5DOrOVC0V+6A2KhPdnajHXmqJVC9k5XfznmhWTE8iJ0AShtSmXbg6Th4r
oEeeAPoY8tRaf55YARL1F75XHcMgCQALa/vOnLCKmDB1wl4Zufdg9CJ2zUtCf+1AJ7bROMeRAOB9
FjHK1yQSk53yPI7HMQEFLYdSMhnutxkGhOSmWhz+HUkhNorYBYWe71Pfi21eMmEso7ycT1joV2fM
928zJniXs7UfN2PnAj9PqlcnmFg9JLSAsYAZY1jxvGfBTf3ET+nuHJ0fjmIy88GwPAtYdmc8xI2u
r32wbkdi3uj1EdSDclEEiq+CTPbr2zp5ndzeu+roDBlPXn2vn4jFC0Z6lNQPtZIjGOlwWl4QS5gq
rq/oH9hQIk6J0wgZ8QFJQ3pIvaT+4DyIO4WbmV775gdtlpseKR3Vzlt04lgZKNJGgwt0yVHOLRxX
TQBO3dVk1sqxGGWpSBXYOk4nU7Lugw4fVFNmTujXmAZ4TpUiLDwUCh0OkcXjIi1O+c5CZFNdkKC4
LpanWtuDc0X5MGmnxe7jVLkrp3FvLWDukCcuAs3Y5uBUaDeqORFR9+zCMsqLvSIc0fnaS1qSdkVJ
SM7XHSJaF47NMYZXFtHsHNTAHB2KtoN4FjJ59yjYyPr3r8wAMdR9M73k1Yz6uxlaSz+VAfPCL0kX
CwKChQqK9AJ4ZxrexV4N7N2saD/uHjFtX5e5R3AWoPPbUutbcjJ7rDrci6aMWcN/uhrCf7e3FIor
9ct4fibvFJFhUdRqBodRJhG5+ZfV9PgiiS3qL0pTmuoZBlTr+WXnTHxRMdIgJzVaZw7rnDkXyK98
HjRtBJivTMkU42SLhcdMktT908qrlAWZ1WoW33Ibkn67EIK2jaMhKxf4eKRus/nIxMehpqKBxGmG
rOrOBj0S//PJYZo2gi88e4k4aPkhTYDuoMXOeyHCaQvgmDfU5FFU57S5GoD2C9k3V9kp15Fc4L2q
qfUSUZLzSaCUQ0dqpBv8wt6w7u/gvyMuABANVf3pLLDmaOfMt2b7YJAk3bZzdzL3igsRx+Ba2UtK
0RTYsszHu+uJUlNLx+sq1XtXfnA23+RCoqN4riT3kAhYdKnzw+oCoT0I2KtUhvQjH8gvMEnVCu9G
w8AsooqY3hvaQ0/6RMt9+/4glD/01vXmcRiD+86WPs/E8SYc5/mkndRIGVrB5BJqDfIDAJruQHij
XqcMMStulMsmP9+78qYgPn31CrXan48FXD3LFsDfxP/O+LBNve+VVoCPYB8R8MwH40uskp4Ln+On
St5PK7eJYwG8ROeeh8j20KPvNcuPIw1sAaSVJlxQoRpRAF8FJqRlTmc/PKmc2t8YFiTRkMyOjZh/
kT6dajFcTmjPicotfzk0zhpbQcapPR8LVNSKQZn1fvUpvPlzY17yt1Wm200mrbPTslbx18MO4J6c
2XEqF4ywStpdshmspxfAjDqgjCQUvuFIrvcuzJAv8clbWcv6dlHA7WIv2IdCbuA1YdmjO0boIvdo
0FTrsrC5KkPPEti6UhMVnqpYvisQvTFVgp+QG4G1VgKAk8ZKaZ92wIDsHoO/zL0Xtt1w/Iwhzzeg
fc+jHGABgmOVLZTKGnoGzOsNW1aKVMr299Fuxy8P/CkUv639JusRtI2Rj4AjeYnER+YOXHjZB6KO
EN/rLEAeE7AW1gbwkBS1Jw9MGJWpZfNmhbV+jQjP8XYqQvqRNyDQYYOnElIZlEiC7klUGaKwHUFb
2sBPnb084eOhYr+Tl8AskPs3mUaWLaxu9UBfxwERptDLOc8CxUr8Jq7T+W9xv/82Rd7zNOEjYysL
3Es7t8R8yJpdi9sZKFhVVygRCjBvMZ2UDpBM600zLws6qBe3fw44E5POZ8NKqUIHD8mnFKUqquGj
P2jpJ/XL7eLbYN5+ZSdlgEWuz598cPGh3FEm3eboa4mbvcqQRFFljS5kmTYxEJaApwjClAmQHStA
mLvHZl3vTsRVExxj6yZzHBW0zmrgDeL8UjFLvh5c07bIyWxcSt0lXPTNJSCN4TmyD0f3uuoB/anw
xYsU/ppWF7mlOe5VIAyzQHeO0Z0YXfVrqCmoyWbOTeupcY7cipSX8UOlGWsk19245aj+vdB9+EHc
ui3CBOLAiMbkRNVIa0WM86RzHfSImoIQphdf0z4d/xON3Qr5WQVR61CPK7AgZvNAYP+38oem5jfj
XDmaX12jD+7yhybDAw654i+a/+qrRR4RR1145FpCB+g5n2IlCKIinnuN0TcsXNquajVO1yiG1W1A
tF89y/P/rmbWC6K5aSYdU8RSPmLjZmwUurhXlq/3zCpj8/BdTH0uYbsP1ETPsIpN0n301insMgYl
TXgv3IUInid8KwG/FhG7jCkR3SU2t/4CIgBqaO8PgNsWyjnziJS6JiE45xq07nGgkS4qztMcrPAP
492MMYjhUX2KjKFiAaMYKS740ufL0s5yR5O1pM7HANYmVc58aabIefMiql5W44AhyDYRs3hB3uO3
GjdNQkDbK5r92JrDGrsilIY2AH1LgVTp0JKuUll9wSPTqOF+uYhACU5eJjKSahFitTeIFkL5mC0t
7x68I53wsHtAmEkagcpGn3EgWf6fLZZlZ/tjMrPRCU0xGa3DnsLLQM78qc73uGCVJvWp5fi7PYCP
1BDovL2l+zWqMG/JG7GjYvJQGLmElqTO1E0Cfhh25WlOU11oMwpi0O0w1luSj/gom3aZY5jo6AVb
ZeB0i49drfV06tstriqD785baR9/UV4jrg2UmCfmVc9p2Gs9mQ6ctvDs/Q9ZZxD7IDKoGb6/x7NI
fVyL87GcGfmP0KQo50rRhrvOnTo4nhLNKhgzHJbw43sJrbi1M+s69wfJ4LXDCgyuhq3Dw6SJSDCN
AjBdMRoQlG5BCXM1NJtkz6KzMu100X40eCBzNsAWo+eoIuBxEzbDqV+B7tUvPit2V+/L3M/11eWt
SHOAhFMJSAOiR6gEwwCPr1b9sjPGdF978JxD4Ef9fMMN9obMKuACrgbcynspeypob5xhi/HGSJfe
ymDhq5dFACqEHyS+KJ4L0shtqU8pSrO9RhL0ous2U+A4s/C9CiNU3m8quTwpMJmIwSiflfHInpP7
bYSL5jjvZUSDuZG8VFuGp+e+eILomX1bhtmB8YAEmG61SW8c/sMMKC7Ab/yeC1CWtOiwG75YXnPM
FEtL5Xw/7LKJfjsNgLaX2PPdCQ4rClTSLhOzlb3I9OjEbInMRlOOpjc7pYH6tyJ4oebJAIdINXGv
3ewr3NjkItE296AnsfZKOzlMqEoxsC0kiYAGy4TtCBDIK66Oq9m17vXYPDrbqxXrRd3Wm7N/S+IE
pfegMxVDg5OwH4DrStnOGmC0xn/vD1YUayZUq2aC7G/nv+03PA42koP0PQs1Gjg0TRP76vO7RCYO
cAGyG50HqZSjLMCavmBxKh5lkU03SIVr77zVi25qDghN0+zjGPTN+jJ57TbuWmWibPHxuw6sJd0B
phgwgvEFEph8xl4JbmfgqFa/J7E7Ps4Pci3Ld9ZiZjiGwLl+vgq1kxiC+6xalxjmzytQq6jB5Pbz
qgR5WdULvocaSFq2cXcTIXg1LgnmFc8yrdSWQCuyTJGtEWikny6eK9Vzd+BJ6GWH19JSsIyqdRwh
VbQ5LcSYc6f29pqb33GEaOYDDRMwEvuidhBzTlVzpZmyzSXsK6N0hwM9hgXUhDp/TC3Cf89SyyP7
NYn/mpDb1RYyQVpeefWSqLvqN4hQ/3XYelUG616w5yrOAil42uHjUGyDQMXJoXxsSabiBA8eIvQd
0IchLG6AgXqw3SLK/64fRzh6k+VhhU2EZfzdUKlDK4X0S2GQFaSrXTazcFtSLJbbs8WYwQKI5mjO
I9+pSgOWuOjiscg6VpugXeZG+xaccFuxXDZ75M4GyyqKUBJXoFY/FIFRj/hl8bCcvuauOdIX7cM3
5EXGt7diCFQFn49MEXZ91YRu/nwXNumgp0ZoAUUt4AuYNFhAcLPpwXrAUJUHJ4XLeL42doyhNUaS
Yj4Ski8S5B3X6sBbr/896ohAQ9TqJd1ILJwOIPYu/dCJOmcysmfF2eUwNN1gK1OsD7c4EyjWX1Mw
ZpIKI0tC9nmI0QufmolnITkMi5eYhvv3U3+f8FpadCi+WTsOt03/KJ32H+k0YERkh1tQwfWBpExq
EBo4gSavaRSQ+n36qkcI0iecWOG9PHL5F4bTKs/kzv9Wunx8Wnd7CYQq9OL+XqoRhYlUITzpmx7G
2vXVPFv0VFZgdSyy+s/Rs0OVJ+6GrvFSLuH7T7XY15eYMsVsTECtJ2bMlQ+E6ETGeBqbqW3i6VyA
0f9q31ouaLzTW5RpbeXjAK8Piymgsu9TOcNd2ZPLAJlWptBtEOosrjt6sB6VrSpHnbYc6juQWJ4u
TRJaSkWci+qUqKypnNAGNZPWMPWk1mOwkR7Ejuds8tRvaP7l2EzraFdbzvjHiTo+w5+7XaBnk2X2
jMff4oOYHC8MvgRppVOR75reKaHtiGEYEmkCFlqXLX8wAVjyZ0HvPxYGPARXv3d0+v4PmHtFmRfR
MWwHmcVvzEdxq29Y2crldKgtOtAHsAGGVNEMuZ2az09fvj2VP7xif1q+qKrvMYfbBh/Rn6G4Wz/E
RpcRLK6UVeeMqirfwOMGHSBJg2NZXKFtwpDq6eNFybwaxHtPhJV6joYavEeGMVMo+rLJj4sAvAMX
pgPp4L3awjOa8F1K1I5mgdMMeyJsvb3J/0tspAkgYOPjn6c1Mn8wd4zuCX+yYE0vtwkGQcZJqS9f
gu3JXaMyyMCFJhTd+56+iQ4zX+EWMvJY+5E05XkaKewV3bh8i7/hKG2/a36UEN2QMN/uAPJQMi9W
Gh2mJiur9QyE0spD9ryRURbqO9oXutFBXpxACSEr11iE5gXQfJ6//al95KZSOFSZJGhiHjwSCwKZ
hT9VpP3A2b1XL+sz6qJ0lZZvqV779P18ool6q+zgsdqpa8CZJr8NEKbJjDxCTBEksDkLqZBqB710
XQ/REZuaqLgkPhJPswyOYxMpNm1V5DqkZm8Smo88ycTleUMeNagPTrWrmBJcrfF2zzCRmzOzV5U2
pEHdktk6BdKGXGMAC0ERhTscwKt26FPGmfRnwXE3bR0FrUWR72egh05lNWC2IXq/xdH2edsDIhZv
KcbYBJJ13mVCz1IJCS2iSNfOD88zSr+tKzgCN1P6ZjCg+0gWTSU/+z/wFtGxL3TuVgPsruttoj/x
7lyA8ygHd3LX9svJViB5mLfa4+qd8gxsngxYxZzoPSimz4/L/EIvjyVr2hYm4ZjxbfsSkEOjDphT
dysrEIRWBI6OejexG/g7rbIqyXoQKGueG6p3OBTaJOW/1vHP5nuIdcQmLNPFgoEb7g0OvJ9Ww720
rKKIE9rO7UnKHDe2Y15N0/t2wmR/d9AYeW8QSLJjrHTdaIGikMh3s28RldWLCoeN7533oGiYEalb
11mpCQ64biVA7VgxmSL5aF5MW3mpa2pQG/fP3LR/XVMecIup5DG3J6TfAn54j8fZrQNN6Rmc1irM
Rv7QWouakbpbRhdq5qYtEWbtfyycwtKjQMUhniJ/F9yWUjlgFFx3U0eYIX/rF9iRh0BM0HpixhQU
C7OE6kSr8ADZeGqqYQX2p1n+g7+vtsafMawQ1w/w5J6r34uO/NeZk5YMxZ2JNebt9h/RVQ6Pp5Er
weF91waS2yz7CWTkqyXv+y4R+y1rQjvzv2JzgRLzPxOdCOt33gCn9KWhf2UsTRmHu0U92om5PwQR
GwntIhRtDfkSgK3hwF30+rAai341xNguZVq9M5odDsDFmuME6stJGcP6336rZ8GDKUwRjSCBJFRm
O1UqgIb5PY5Zz+fD5gDXewMslfR1m6rU4lY/BFxLcsmp4IvocNuoM87DfnuLI3DIhw/mZMM9gdkP
D/WQgVn6XLL6kJhBVydvy4/bEnGoSxxds2Mm79P8mEhv/EfaqIEz8tfvDm5LCbOLpkivT1BI7tnd
sBeGFQ6oq9N/IpwyWfNxEBx20KqGVyVWskmcD9njeiDXkQSkxj4KG7wHQrBaKCUon5+ZfETEZas3
l5R9uaU/sWQNd2YjaMuSbkCEYDuMQyA7dgd4G27J+/+u2to7rT4a/NRRcVkXzaPRrT6m1ejUdbNW
D789ZdJp4NbbS9LsWa6ULnfGLhVSDcFWgaEkia9U+rYq3qzFOOBcJAjjs/9hBVCvgbTjSXDVyYba
nHcI16wchTNwwy1ln9HpALESFmgAnP5FNH4lp4u/tnLytE4KdsFAVfIwXuIHLRbu0lskiFs7cNEq
RWigG5C6Kr1BxsUXuUJupzcz352FdOQde238vvKY4Q0R4loFJIWW9XBF8qDGoH97/CsJsXroX67v
Wwx+qncSbVyp9HCCQurz5rC8tZLgejaMcUGvvEBdSCxm370zQ8fB+w/CHhi8ZbXHwQJ7tvirjuFD
qcVEUzeYkkkgrGGvnL6IoGfjNLHGyQMvjkgGQ1px7KE7DPFlIB1Kn06goHalyGiyV1TUx/TSjc2T
4mF4VsmF3m2zufvpsFrPLtRSv96nTCxTZt4wwaH+W5hhJT97c14h0Sm9A5cglBEbmk0MwfcK9y+i
nUPTigEvevDwPiqLFxVzubDzmJRoJNs+ge0N8YtGYa3BSIwtbsQqraOq69ebfMS3Q2ptowXfx+hM
Qkk49KDIbf1ExneQ6ANiUAIq4vQNuDZuF4xOJ4qveOTLFgIW/0GllmNA2eaOtp88Ghd9T6ubvs8p
WlKZ/hI5z5TdF0pZS+DQmfv/iudCc0V/2xxgebjnMYNBKtI8NHzszZM/dlm9WuSAFdnTl/TIeFIU
/67sJJHDcVYYmtoSQbp0bsPRCytWEtxC4L1EvQOGPJkaP+0WRJrgsZOR95t0cSP+tjOipwPaintG
fGnjanthP53RDP80N2mYgEwZTTDZzZGNhpHwCDhr0EJQHpyNxJthCxJvRUzabxpT84fMbk9B5FXw
F9CS3ocWQNEW6IK/Fb4Wa4iVw8BFDjadNm+IIVKwGZvihYIa4GizhlaNUdaBGS9eA8ZHvlhU+hzU
QYzDoG06l9UC2CzZHBbdjEDnS6C95jDPrQyuwqSkSQ321zpSWxwxOqMBz9Yd43FQ1kQe0XXuBxBv
nohrVi2uyAZkqau9MI1iTWU9kzpGFdIfleTCJziw2ACQhgUqCYY/S6vdAmFpxVExRwSLCQE2wCEv
1mvYb7IVNUug/w/flUeY6XxzoMsihg29Ej5XW7d4+WUJW9DIBK9MD45DI+6yvgsPqXTP8RCWKptF
8i9Qhe79ER3+7MbqwJILm0EVt5T0cVKii8lGj5it5MbPvrRU4AeL1gH4U5kfc+sbwhTfU3jg4G1F
qRv2+YRdRhWbTc9YMGqUnm8zypEP2D9tS0OnAo4TKQFEYVu9/KXuAHrft6UaW4bKYl/EZ1peb/Kp
lWRrcskEisNbk7drV/ueiRymXks8cn5HlwhzMz/eeMbqf3xq9ZkwHmznaKT+xZC/Tzmr6X4F5sfB
6SlQfJscDTzOX9Blc5NbSaZjO0tyYSX/zjKFnER/3d2gjbZ9OTDYRQdH6OIWs83tiX5Ovoq3158H
47sxcYJ97qmX0XaCjsqP/KKMFdt7tz4wuHy4FNlOP1mkrCV8HM7KJCZWukJnTRYQynxN9FdJ43T0
QDhgQ3u2abhnoZuGoQTBhSCUvaEBfi7xGOVxJve/1TcNmEjKskelXwLeMqVbpRg7mIsKc3X+MDrf
6pQTkwDglVO2mx/AFkWzRl9Sguxs32ZSMns64d9huRs/FHQbMvNiih1xPhWQbh0iFdRQu0SEXn+X
AWrASpOWnXbOXELvDCVYe4c9wQd2+DBMxkn9r2MJXZEsYIjzbOuIFGATNiAZoT6HcabUmJZfL22I
kZafV7CabHuOBmr8Oe93h0Q1+Lk0lNFD6K8gutMILleSCs+wVGoZaMd+cPbtiES0yqBdSbACb2rd
18BIU87sQmiD565YI4idaCiRBBau6S3jHTq9nmFp2oEh8v+Ha82xWseN1y2j9GCqNzqlBmkdOG+4
pJI324occL04wAIRVGxriLF6Fwr0Pkv781uuUZEkzspRNIrAQtkVaUEu/rwfy2N3ACjMVu4Dis2y
s78gHwfPvwU59+RtQRo/j5nWIvIvHHn+7h0XLVNHmnC29pJmJortSrZsjGOjV1tlnXd8byG9/5fz
Kg/JAL7GH91A12l7JjYYCid7EuINcbRrsaxpvLXtVxMiZxnJSVg27m5mjKy+zmGUJ8wl8H9fVrDq
Gn6quFoy+8KpeIlFKZ0jTQX0P+A+OwjUQ+LoFlC5/ZwCfDhHqg/sQ3x+PI14yfg0OhsaaJKcpJNH
xmh2POJVrF+kxVqBUlNR4JzO81z4r8e945TIuuRqYoEse7bidqEZNHkpKeOImQw409cYsQDb5BIU
NO74W8xwmUOXyPwQB2LnjT4EbzUlAs9e4dtChl0aZ3aKZDlGviViMgqKeyZS/9rMg9kQF9m0+Nm/
e1p3MHzaT/28pq0h07Gt1vqsr/ViO5Lmt0MqJv846q+rvfLlc6f2bBzB8b6JZMIBFO/MqSnCt6mm
kUYN2L+Me/bxkLEps0zT8tMXBGzvpoEy8mvoWIf/xxKrwkFXGFnVw2GOprEYaaNPoQ93G34rAAnr
sRerA+/pE2/ymv+yqyj38dEUrZ1JNZU45StNYiyf464oZj+PI8Ra2vixobuEXuIWn530MBIofX/V
pcWaInXw/KWllUySJWEmtYYozR6Yyhj5Fq6LK5mnauHS4ve6tl313Um/se2Z63s+JTI/e1wrW6ZN
yGtFT5LTFFGGFz4dG/LxyMwhn1fnPZpbA/FggBJvqaDjNVYwpDma4/8a+ztpdLFiaRLin0PiCejy
NF2JmPQumPRgFCon5J7d6+fFcmq4PWGQUL7vZ5EEc2ZnIO35hh7NSkl9xxr/SafY6dWowte7Irzz
L23GYq8ugDRMtx7mX8EM3YtJpUaQZ+42ggA1ffxJstwa+zix2NUX7e2VcCkO1tT6UukUoKhhsQ2h
NnKDTOG1PMiEHVSTkHmCNqZzDzggsH2kyj77SmP/JVH0DZvrBWInWOBK7QqT07aYgpBmkB/zeO1z
YF462qoQZJpt/QXFA7sMvObq7H+rl4uRF4aA4O6i1gTZ+aOJhqr+VkiocEDT8imMnBnZlZlXIfcr
gsY2iDj6tVnj6XQaoY7jRI0DJ2uM5iHCme4AYr7GUHuv4sZUHs7Dsz5bstGaOQ5O548+B1wnzHFQ
E9aZ1XUgpvPw97gAho1CI9BCw8yobn/Dk9433niLwWEFshcMlepz/ac0q/TUjWIgAx37+203tYb5
Czuj17QSNd103xUCHo4XHmfdE0jVl1hvuvrE3+PrLksbAfoMjYGaX1xvt6FGffNq2TdOtbmLPyh/
pyTOCuxl8ymw8migrIHWBK5Nf3LPx4tU1KgZdrqE59t7Q5IdG6AHHTWL3xYgtbkH+VfqDV6hHQ7d
gITOSPocRvYY33GNwxpKLeebnCnELM1ZyLKGVhz2+qOJ+1r5EtdukBJeDnztmfBs5658iJ2wyUFD
kHizUzdq8CC5y+1ooArXx9FB97Hht+qdwU0/FkOqjPOxKdV15lVReqN8+uWUCsJfcQZNy+oIgC0/
akp8PIT7m+NTFELTzWAIduSExT9OWg+xLGT38lNF5dLpF8oBzZVuSDQZmUeDHS+Rst1f5lLK7sfP
kcR9so9ydCivGaTYwD4JMzWa0xFbNK5MDTXxH7ufIZFLEQhhFkCQO1uTivn1Lycjr+VF+oamYfd8
jOhSiDD/FlVlfCrTvjsUUP5XWSi+5S+22TyCkjeUSaf/TYtHwTEqiyMlBeoTh4LfgbbkldlUTXFM
i86Rt5UeZLWHn2n9XYRUABFT66Hc6Mztah3hFBeSqu139Sv0WdHen9OcX9WUApyTP3g11UjaMvCf
tYqeVlsRyNJlMu0wN1cQEq5xkW9+3yF1fE4dEgETmIRcoOqnpjLfMWWsvgCuyWZnOpjAjq87yeJ/
cTnfp6wt6euKqLNN8+Nfq795cTK7VjsiT7GMqBtgNvvVZwlFagO4t4cVneQ6ZhOfanPrnp0HGoi0
55hf5uno08HDdZNA+muORKT3fKI1XX463HQV9Akq1k5lvzuM9FJP3Lzp0Y7K9yhAY2rvnfUX52nZ
ZlwXjlFm+6Ut2YGLoj4mUPiq8BT3Vxe0ERl4RFeFx+iD3/K/kFmXa6kFmtbM4ftz8FN/RzjV1d7n
yU422ieVDKrWgeR7Rne0y1hdorwMnlF3euQV+p10UcEXA7lSvSDopEx/6aur63lbOK0nmxsmCyhL
tVddmye3ZDRx5Iu6BjnQYqGSNuNkK2oWGLIFSPXTvdhccxN3ryPQhf7KoDwBec+bzd3qpHiL/84z
lyjDgbAjTG96+e7YvjT6F2ySa3wi5zzz2Q3KYXlAnlrxLoAVh2AILKWBOMO1sDvnGXkIHsA04Zrf
t+VkP8X4MP6dITz6CGPk7DQQdPwZKwPRRAJu3LiPSs40vooWB3WSOaYlM8QHIvBKA/DtJZHE9Kk2
Keb3t989C+9EzPD3yAb3csdec1x2RXTk2Ux78OH977QbRXYSt5JsvPprarhPBtrlCUVW1Cni/+Mb
13loKUzIMtce4y/NqoTR1UJxGPNHZ3aQTDtEMEC5P4VlX/O2Mw0l70T13M+yXU9vOTTNrt/Z6Oue
tkewLJpAw0aV9SW9KwhbG3y9ttNXeeQ5KGVOGZ6QA9fHMmLnPMJIF+Cr5Mm9PdQV+U9a/P/d0eNm
TGAOrZq0V+yYYlBBkCeHdNmIB3myXOIQyNLqv5V/yVJs9lKYmfzTRzS7oDiUvXkMBryxPaTE4BZ2
Rf2hZCJth8gv2OgaXGjAJufbcm4JuvKa7LcXo3GOFYFvlKdDVRIHa7x1xwz1NJg0wpForSKwhREK
66bOpQa/osOZRKA9NFEhufiRy9quXVBwtEBQp/XVWahvKCRI64HS7Zzav5WT1yi3hyWbVbPYcXq2
WPkm62FQjXT/Wpu25BpXmL5RyyVAQ1/YlJaUlNM8eIGJrSzYNdNcFlL5vmvzQSCHDmrSUCtWjcr3
JFFOeFxdPxViZYGkS/y2368M+2KN37DsZ0v3oFgwmm47qOBkjORY5fjXEyeYw5Lko0tKtnMfR2pi
DWo7dzi646ETZame5yrYjvsUO0Ujn4DqBOHKn+IWduvbcep6TbEfl0xdvpFM3JTJC9E1zS2sHpkd
gaVPMRdionyBjm0kKMj7qqv2TVpgDb49GcPgmP4ONKbDy3i6IYsecIFGgan8Y12dlbyT6/A3QB+U
Glov1EiQy5zchsoBeeWbfzMD7qLy58W95TFEn5JVv7T+STgMeVwQdU4FAMAn/qUy4lIoVmpk5Hen
ceTeEJGmVBh3aIv8SlbEYZAUa/iSe4q/BM1KQiHEP6Tzv9eYNxmm+D1XFdrLDlgDyto3IHDovh5O
93OzPyZZSLHkgGTmgiLMyXoVMXuBuo6DBYPzOx8zib/Ql8815pYE4uY/DOtH7eFfu9jy7bmn/ioc
UBeV07UzOKZ6m7ZJosnkJn0tPtApuLxLuc8BZFoyf0SbHmPn98/BeABdVpYEyG2OVSX2nHwIWguJ
Uo79cbaq0rXzSojA+6Ed8vvd1i0nkVaR+pIDSwPDuzA7r7G7F6Xhr8x0eNaEWiely1WIrFp5C8y9
8WFywuUiIeeyNE3H4QZvsK7meiNGEAof5JxZGcehAhjhrCt+p61YXp8ASBdlFBXErPreWwysrZTt
3bpoDW0MX4j22RRDRh8+hsUvVSN2MjE0j+XjzKC4X1LZhzyfXzCg6Teto4yXx5po1jpoNJV8XgjJ
WHRPQRXIx2gNZ85Vi68GA9Ca2LGKEhu2kIWnvGC+4HDLGP25o69KuE1Eivywpv/qXXaRcQUxH6OT
+LcyLPzqMIMK2I8BdxKVMVp5vioEyCeWPUtisIQoIOZars2JrCAp0Al9xYHSy+T2QkpAHFn8VULC
odQOaffxQ/CXOC/FykHEAc6BOk5B34KhWIS0MMyc+iONi3JCTOAKmRDRYVMaDa2YiVAPGuX+hOVr
Q/spfscJddHtHhpnRIk1yODFg/xeql3aZOuCT0ubza28PHuOA4HSkfo/3phbeYTcubHf5l1DTsXK
DbXoBgi9VL90gVNQN6TvmhvZ2AFrPkvsRDzXL1/rC6etUwZCMikyowC7d57+te0z3dMVU/qHBC/C
dloIT/sh/UAPzMn++SrcFJM6ukrNThQIQQFjbexrfIqj9aOfGuRWvQIqG3exOpHkPAIV9m3jQqwr
CBa0TQiMkWHxlfaJPO5KCpcywZAfOVEyqfASe3Z7/emIY28GjBwwbEbINeKXXjeBp94k3hXWCiOJ
AZjML0mId4tUqaAkg56GKcrcZJa0OkSEYIcTkZWb00mfB8lq8Y8mWANKUD2p5R7eiL4wkEh8L+8s
G7oc4z32NV1NtTzdyW0t7HwxFYTOpSC5rzk0CHebubN5xUcQFC68yTSXzhGiLt9o7HEtXWjAMYV7
08foUpe7fGHuUFK6oViDRLlOQKDV12i+R4X+kyBUJlASIDTqgGO5htQJG2oynOdxlEXvwMLdGBgm
LKKdDwVliIAxUgK+Zd4aa32W5fifyCcbop25rgx1tkp9UcInhPN/5HY/R0QKr+as9QwiJnHQcKCC
HoNAL1yDsyd+GiKhSismGRNzhOXds7hyXDGoZTuM0qpq/mPygk8OjtD43dr0mSkai4j0Sdg6wMRu
8TFlCwL7+kJc2K1uNJUKqQ0xLzyfGY/vEt3yB4OCxY59zfQ9112q78zos54oNcPyqrhMNDMM8DiA
a2VlXRK24+KZ5XzW9kHplC0X0QqK37qRvfiwkr3C1PK/6JXPTS1aj57WV6zVOnDQVoFhY77A+Zgn
dy2MMEzDuEjXAbCiiCo/Fj9Oq4FP0pghSzOrDEUFCGMnMW6nnGQso/rctwjWuzfE5ICJJu+ckQ5L
L91nwRpakbXx7Q/dcq7WZTseb/UHOQQkViRRJt2oPfbWeJa+CYGasYvn1j7j/7hiIeKBuIJNiloC
D09vFnr0VZMKtPMJlFvuqo8HDPQy/H1Sk3lDYKQveXYPo9g9VmddK913TxoCXQfWTyFT/dJijNNF
Q/z1NNfFUDJJXxW7rlV1E7mASVtWJDmvEBnGuoc7dTu85plBRZ8x7x5kUPuT1180S7qq29nui7+A
OPkkMEUpOofaGJHeI+Z4hK34tVKuO3fNWlGHMU6Pveq1iwPrJka4jJTvvVuAhxV6TLOVcM5ABB9l
avD4Ia6erD4JwgQF/YOWuzS2Xs2A9RG375xAoyRKxJVpJqosvjzJnOIEx2/daLhjxMUB5f0bOtML
jZOCAhAjWpx1PeSnINBNHxHyFVGGWufgnSZhRkypOqCmDPBafuNqllhhNkdwOZvrzpFLhFLyN1vr
G/rtTiO26/4f3ircY+2/aoowQWUwNGuOYS8bSFvROvQd2lshjBwtoqMOzeZFlbTP8aFGLsoSStQd
8zZ22brA44j0JBpFWWtNtdwN/Af92PJYWPQfb63XqPqCuXeEgBiFu27tBFEWg6mZBkyotoAvbGIi
tYSzaK2irufLczbhlEjsxl+p2UKE6te3erA41ej6HzAE4877rtIYacjwQV+d32DvoFifBW+j+Pec
gNGoEvyou3k9hQ7uXKAudvXSV4j9PFY0uHvphVavQ7MdzS/f39jdUjmsH9HhkH/QmrlVcFlKb/vf
yMytphuQ5i/Z5raR6RD+SZe9W4sFXF945rF0UFt+hYRFmPQEqthnWJyz7rkB06117R/B3br36phq
AuP4LH6bmdL2SjNv/zLPC5tYa54b5Egbse+hu98klZQnEhaV5vjgMvWzxqxuZ+r4rwX3FKZqxt9C
1bgkRUk3VSH6jIuI3O2qs5U44ewpj5SYUNEkKmFgK13WnUo45qUoGRzoXzcEloEwwTU2JpJyocMT
7qEP3G1uzkiJFz5Rg29f7kLuZ2xtNniw0C6WBUtMW6Y/SWAH8wAyyk+l8lt5AcTPigd2WCJrXr7F
4D7ol4Z9h2vWo8QWgNBgBRwyEeh/4I2KILrufuKVRiDssEniOruH5Irchi9MMruKhrw8vxSMuDb8
SqAs8tm7I90ViU4JYdgg88jrXQL2I+8HWnw/h2LRh/ebTrWO19kJ1kYtKr1G8a/AvSOrtO21VGAb
rXqXbDfqnr5ybDkbv6kGAk8eJk/GhY65Lqm+4DHbJrp+GCfCU6SoyKLc33LgGZSo+/6ZAjGNBaZO
2C9DID2D6JHdGh5Jsvv2uBf/0VMfhx+GIVWS0OiM+4VGVdHIQJWxZten82RzjyB3GpuWlBheZ3Gu
NopenYiIqCi/G5vX/7EEkd5svQ+5RE9X4dZdkJdFenRvAIZDU+MD5vqYkyKYZ/fAtfgQEH8uxJSK
+R/RzntDH5vI7Ag3suELChflW5OYUI3d/wp0VNFrNzR9zFplm1fz6T1BBpH9FtQo4X7YpQT+Ec6w
c5nnG7IPO9COBeIHnJpIIYpuBEBw0w8wqUX0JmnR+uWkdePDWTFbZlTUB9+Nu/8rAty8HeVdO9vv
ThHpTUZBoB6L1gto+FVcGvYrwGfh3ejtxj5Y7r00gjYaIbQqNQ+ihg6L/PXqPUEB7l20eazKc8xq
PxpiZgCHZ8CnQZlTHeN0OEdNOervNeZPVlJuk1PyB9EkXH1vz/5TMkzl/Oe75hzw5DqaikAcQt9m
3olgaj83RkiSPb1dt289B0E3QIHIu7jkOV69thUBU5aUXFyAZD9x3Vs0IBe9E3Oen6TTKEWccOi7
geVgfGp41yjbcV3/nIxZbyc3T3fjyLGsSYFuSNXcQBozyoifC9N2GfgM2CKu0BJ5pSmQ/0982kXH
BljzTAHd8slpxDnwTDp2dOIOZgh8PtGe/uV8UC1UD1bMuK8sHPtWP7EGcGRR16otBOGnNo/INv+U
s6fJq7XYfpS+2zZ9rMiDIlRV8uOv8WPyKvpUZuxmX4N6OP8vZy1072LsSAYkyvbrhpot4v8cihd7
kixLJ+JLkLI7ZYyk54zfrT5iOXzy8eQeYiIR6xr9p99yHAg+GyshHlXNscQL3bvda7Vnm8Z6t2L8
HQ9FlfCHE6Jzvjf80GatIEbMnuxOOGxjZv0bXiWJUxTICkzFACEyAiRM9FeU4Cw84UMCd93WrTqa
Z7looLdgzPgIIlmPy/iFR/SYddZ7aUAgPFlyRFqRabHWD5oRUgaxHyj5Xei2k8Ls+zgUHGDK4T3u
tljPfDvk3rFNyw+nh3sEMv2LPwibYslalz6ue5/zPlawL+lViM0yEVla5bSgdY1TH3OfvMxgH5Rj
C63CiEYM5LH/oxiLR9yr87ieoje7+qKfxW3HM87Mqn0EEYtV9841GahAjCDJpq6C2RBKih8kvLd0
4QnuS1pi/EzLZmXT0i8JRikbaf8zhEUjBfYHgVUUh6V+VbIrx1/oHsxh21K0ydHoUSsvMpyosWKH
hIO4sOhVRlZR8FRS/KNi0UHD9ngpRH85dMmzZ8USbXNbL1CsW9h11BuMOuExDb4cgnyFin59otMD
Uhuv/cdrw/vUJPS9zoQiDF9caVLMGc9AdH0XXt9hTTPckR843BsJ+deJrMXXxbB4g7go6gZLLmv+
axOEAls4jMsKntMjttB/9gIh2TBBg221yw3PwjHdUXan8YIAuEF/Ua47FNDjPjPXCTBwK/Nou0Lj
tP9LikjnSbsBso+63yhxEHeDKjFZlDem518NH3gigmKHgotsTcJW8RWqcytA+l3Z4/+LkDFEtU/R
jc+swm0xrU0gg+65gKiFT4+2BxhRedFegsvtK+LPx07B1+Vw7ieTc1qH6RsLM4rm9N/vxamriJdd
Kwz6iLrhKthGwze6x6DhbBHqZIdYcBvjmFvDKe9L6SerlVFibkzTqkAJMWDFIQnYc7WRyu++xaTs
X9Lg7w5EIlgIC7603lZ29OpEQtcX5BlyzNOn/XHxSzWAIzztHv5uZJaeWp0afEc5O1zKWdTP1qUE
xKbCev36mBXFH06E3SGfiHqrBsxTZExZNH24sIvgtikcSBq376PW3P2DPFSPW0vT8zqGgFw0vcMr
rg9kxLDAEgC3thfYUUzQjSpKnYYK9+7jcKJAIY8TItQaljjyCzqbC5ojGq7CPC6aRDd9UVDur8pm
yrO48N8XKWSQ2RKe4AfOBHXiTmy5rrhchOGitfC3s/DXivXc88S/8FUJN2JKcbhwMj3EHhDmQYTe
o6rbJpuBEDFv2ELHCjMROPMlTITKc/j8mvlaBXL43wQCnfDSrkwGvYK9kKcXZqbGt4FsK7RVPwWz
sd7sqKkLhI2HWfbqFdZigHtM1gwNo2qQ3G6IQkJINvEOMZ8SGpMmexQ3bx5+GQYV1w/8F+JWVdZ2
1+3MlfdsIY8QMuV2wndnL/fzx9AdgMBXeu6c5ycu6ZlLExaS+yLqYexj/qe/v259/b7Wc5Itg1Tq
GkB56/E7AcBXdF+iovDnPfA4kxe5CiZBQMhIHxbhlkkERO5fhy6ICL63kcxiWsa9fd0WOAdMe5x9
/pFuZiafSrAHaE5lZbaBrUgF72hUoQcMFNply8LswsqJ10z5i/SbJkU9kD9mewvs58PUykZLWus3
UYEr6sg6J0iVJ/tClRGhS8vi9T1KI1/2X4Gp+IqgAMBZ3yNWLidAU/NcyYOJsrmnmdR9Zz5ardcM
cjb8BI7qTPAIUo5dby9ll2G09fWRG7Ni+Ps5Mxubnc5kQgriTYq3IcFocRfHFRQABLInl2YvsMx6
2kh3FiJyjZcqBMEkZCoc2OwHhlcGGNgXAlvlEASPRYIORp1jO7OS3LXfceko9cBKsP9ysSWOoSHD
RZBf94hvV17oyZID5qLlxeRV5iyt8WP8oQ9GbBsu7cH69DZgroI3gRBxcoAisg6R/MseEWE0P18S
jbfpzM/zchMbd3mjZTPlCK91cs7eL9jXqgB4/8MIY7vQ1Rmnr6zbtj4OBW9YBfrEwtm3MOk188DK
61Dce9rjSBkmRo8PSwgRdB2OEaa15Bnw57AhgBHSq61PmdO9tGkKePAaH2cs2GkV6tSTfGxBXL23
EM0SZRIZQwymb71ycINTj70ams/2LU042R3YUlt+OMO/VbAZikLQm3KJ0dv1nNbulJNPPU66DDE6
s7B4tTimyWFnC9dzHGtuDkjHHE1iPDy1hDVqx+upr42P64oqryWUbi8lRDLBZX5wdkIm9O4pUmBU
fKnf4DeMBoBdG7bykiKVUhUQvBYMrKCkDf8vsfUXkUhG4TVgPX3GBLi+mCPZ9Mryo/Ok9xOLZIfe
bhBfVqSEN/Sx1uLJk5f3Od4g2mp1nbZBjs200MGaGaELvPdXVVePVoO/5DOKpOv67kuHAjKV8fP1
/S/KYcfLBhggDbnBVqvP/J/O2R30FFwpt4fO2/C2FDN5KDfKwtcPGyepNYISq0w8WbvCwPtQM5KF
GIe/aacqL011fcpNMgNbY5hZi5NNIVsuTsPP4gtnRR3gPVX0fk0oixwSpW6JOxlYApCPYSqBBFcH
xZ6laAFWiJJPE2hyX13LWd4/GQKmw3SJ3Bd+LfOivv1lmec+VIStX7FaYSoe4U/nL4u8BjRMzuyS
e3CukGBogGDqDSy5U4dqXGNIAYv+AGu/O2AuEpKbuWDqYodtHgizqxt3YwnB5Qw6AWk3I1bvfPiu
jfVU4CU/H5IiCufFIijmgAwgtdytv2i9QbnLWPRqjUE0kZo1XrigQXxEoMgs5hzFRQC7NJ6tlBQy
nvHQzMR78oFwpkMJuSbqSlwKolsOA7k6l04mRUHrxTmG0AWvBd7a4ZVlelohhrTQcDhBk5EpAY0M
f6SmxbkG/kR9HdeAtKKp0yAS71Xb3Iy/XH1W64fZxv5fhMu6x2nLf+8iYvLtkCpLMy3J9Ianw9v3
PSufrpwdTpCX+PC9lA80taZAKRGjCji0d7Lriga1dyU6mNdQg0hmeUNy5gshbPl6lKFKaq4gmQ1I
cxl3Dg3j9cP7T3fCP7xMP6gBZ8mdWD7C9eoC6Lncmxqa9lkz0ajbdr0ygszL4ZSWMqIbmEMAzYEE
lb2L2OCYCmeuW79CA6K2o62RoJCAQ4C39WtxIGRQ2r9Z//ii408PG9SPLtZBJhz8ayXNkXMSV9ab
tJjf9nnJrO00KgoMbGoxhsmRxwOdLHag2jgsw9kXiIWsfTKUYNkidNz0xZW84mkyGfEN/LxyEBNr
48BvFDqXd3XplP55nalKQ6Aes7FKOekgSxonthSR4YBrzQLJ3FPhgmwaiM2x3/6plzRKSMFIeeUS
u/ocv/QiAXC49gSGK5XJBXK56CQ/O4FVpt0J0XhxlCrTsY3a8uZhETvvMdL07tXNi2xta+CFWXYn
1I5unn57FMyW9e243FyRN1iVCkP1yHhcDOneNrrRAbrqRZ6q6xAWer7LEY2+yJ58yj/gNl1Tfe4p
Em4zDVrhGQCWgCxl+re1wuS2VnvT5IMtRejQHo7ehToqs3EW38IE0myGvzIdeISKnixgcJnttbQT
7q2koWZUs8iLuiB5cuWp8/YYzrN6xy63cpdV4GRcKmqgp8t9ji6t+zRh4JHUSsHUltrigfFMdX8K
U8IM2aiyiDsr2VDh66J3680orqFmo1u0G1O8PrrxnwmLuwLURtx146THO6uLj59XvmguQVxVPsfn
vEshjHWGNRjk2PzdUWG0PYXPRzKbWcIaooveTaCY7Zln6K5y9vkNT1nc07tvkiUuDstoCKUEiWJn
7H29wlS//Jci4IA2rCCqQBk18+PHvSDomtwIs08vDGK/8GoX/lqX1MEn/IwL4RFUvWL4uQSJ0Q0p
hN3E8ZXVcgfR+LSPxNwypaHfcBts3FY0zwhtlJZr7lJJUG7TdjP15KUFSLfHb+M4tuAUdOsNB67v
+Wt/PpErOtJpsA8jsGVcDNH/jpJgDuHQv+RZgVGGK/NOs1+JkKU6sIn6qZLZd02AQjlzJVdPEA5V
RKTFDAPIFTlGfZjTODJrrypmA/EEgYL0ZCIRaFzE2/YjH4JZDKFga2xepub+oEB5MDY16wXowbGv
EbRy95kJoGgHw/aLpUxcSB2do6AaxiPttPPbdhhe9D4nt5fy+vIoRnGCkXT2MoZtBDfgNI5CLkk+
W3r/nAzWYJyvuMcpbSpWHHNwZOwXYz3ibtFCLtnIUmpU/KyzagQXx18Od+xADgnx4hoHMBsPu21I
3WpW7XSv6wdGzCg4D0jBpb1yHeZTv0qyn73AYwBb1lmS/GcWYG82o5kjZjFgvdneuW8MnnFUOS0e
ZUgC5pbAojtIKjZMsEoYI30goWMtfKT/nlL8GIoPUphTZzdwxMWouf7E6mNIdJ2DOF+aeQdhQbUa
xBH/0pb7qnKI/jJN4CyOaq1yJ6K/jU2wLQDg/iq8ZalGHngfBCLbZ3OhD+/Ahsd2CK2GkV/cqvMJ
05bvwJmf3rHiUsICaqAeWYv4n9n1IJ4Yvaz0bssjE0pD7x3Oiq388+YZcvTdkJC17a8OAwfq/0Db
tXZOezQfbQzUgLcSx0OoGI8gdyD4UyaEvt4C36YMKaNdulQJpm3GXoaFpeF8TxPOKO/XXXZBjT92
ghyew+cw72I0osv0gJoIMdZ2jJOb1DIaMNC3IX3t/JUwOd4R1q43o0yY1+rQv35etWSLlNCXI3wH
WwS+xwQXtkhgiebAT+ZHoN3AUZ/W9RI7xHNrz0ZUn872T6O9jnrAkqII1RZ8bhB1Aawz21pU2ZL8
K7jFK0vUDdHov9EMNzZwtgshfG7vMcS1bVGPB044hgCFL6VT9192VRKRoJhkdP50BHUCFBBYrv71
l5nneIok0504qisUOAqXr2cScHBT05fbtjbNjQlYAuJgyot1GPIRkOnhU23tLyy39apqGwe96khm
ocWuaF4REUxJByWapkZfrkkBVmlpF2MvlYSINE9h9UUs5lLH1uC36iHTBbS2eaj3HRn4JIfUYMAA
F8FoLFPqc5UNfcAoXAwLjFlUAkX4Yi7PTHcv21GXlWqldcp534JUnM7vzTr3VsnfP/+QQFrBZVBL
5WJdDM3kaN8pjcUtPx8NrNOXTLLkJIWrOQj8Olqsc5bceI0Jr1tGkjZ3ZYdIcYGzHjNP5s5s3TZQ
TE8MWZiWIjRus+rHz/+m9Fo4vmqzqogAwY36T2yFUvy09af17IvNQ7MfeyGzZ9YKW/qR89mau4pZ
hvOFKnhwkcQwSqBu6so3ZKLYTCmK1Sj6cOsZahy4qwtJNWvpdnaHbCHkp/ulBxpyjodmvTYzn6Jt
552xEJgGDmo7/5VlSHP46YWRMZ2fvxktk7aNuWQ20HevHSQwbHpxdFl1UdDeVNqsZqcSSsI1HALK
RKNDROCeLVH5dJ2o7H/DGKjKDF/6zvQm52er7qvgvP+Nn/iOIlnu4jXCcc4k26xrWIstdkKFJHq1
mFIRT47l+IFJcI3Etz2qEvU4cpHBxQPxGKITaewzJ5YM/WhkEpKwRb82TLWgqE5pfl+6Ud9MG5p+
akMGfmI4lo0Sx5+jvs99S3cDa/f4omNmE3OzQfAU00FSmGRwAf6dQhxfk8vyxk4c2w4dZR9KtRFC
6E+9jv81M3M0iEXWBD6IgiJA1EZ6hT/cFHF9chQ99f2tY04TYJ7L8FgAXl1qCqXZuwohvZcn8TU6
d+JToaI+5i87gx/xuS78jeSv1x4i190b9DR3ths0ZkHOka577ADe0uObYdpZiprZH3e3XCMfs950
X0sQUwr234/Vo/a75HhCtt9ukFvcZy15GUoQ9gt/m7m0yjWLFwQ0ofzGCuGgo7uX2ZpSv8w59GrF
iiM39Zbl8M8n4KT8AsI9lK042Tkud/xKEsxrHuNTEJz1W3arKGaq1Em48YesZX80bIFl3Twd45AQ
iK+rXcndXknyORmIBU1WAqxxquoxj/X/llfJI8wY6wuWnuKiYLY2C10ASNUq8Uxz+uKFUECjrDNL
4uMx26IfGLLz/TwTCR8Cj2UtjhJ0AApCuHqRybBmgtNGFI/FVINwBV4sD0FouiBi0CgQ58ADyp6f
VlIoypo2VwYkVXIXMFJA7FqBChNFLd635amncpMBQSBprOobEeEjJ6yFgXlYiz6I7Dt77yB8Up9c
L4k7EjBYr3g2nFlzFWpXz3HD7fAyAlqHihQXqFh37vsBrkyKYHf7TTD8zaqe4H+Us8Z9feCH7k02
2zvAzB56CyudRIyIf/udTBSVBmH/B4SfYpgAc28rfwQNIZD518o8Hpn8WxZW8JEPI5cuYC4brpO7
tuPAMcpgGrHmK6QDtle6REbjAYMLSuflcStntMSJmNvjG/oR/Obs5g91DEgX5DtCzQ9K6R8d4me/
BjS2WLg6ve1JiPMD0eXgWIZr1wm/0bnUw2o8rwH5++qHPadicJH1uMPttwtuQ9qnt67H4EwMRK8b
pMhRTP+td5/0pvPvaPtHfZHIni0EAheFPKtJaydtTcQHYlht/QBFeBAPul6q6ksCjOuGrJPoMLT5
0dl9zGZfQv7RR1TUNc695XTuqEiGrIMOh0qxUZgZIr9r+wyJmVzkZKMXZYNquR416bR+Gw9G0TsC
ptFbJFrgNxmjNvLfTNhDq2Tttg4JCjaSq9OTrjoSv2w4s5ObPH2lQylLzEBjZXD++C3+daiqTcwj
9XLlmqj5jPOKcizLrt+fGBEveWj3zjMt1ddnSvyYyuhE5oK0baTS97jiDkPy58j8B1acu1VJdOmg
fjCe1IOZS285kARNSSSQYUKBhlvaN7hCpbyJPtf5A7mv27YsXByQcPk8gNyxCOM3y56Y7aGC66lv
rkxvMncMSzfXmadW78TaM4toIeTIjUnrZFbx0grmkqCsm6t8I1ZwhUXjqRZkgOgxvJ0BfC3+H4bB
rKEj/YPRCWhy3HBkVK/FScmSJ9Ne+FY80glBc1oTOLP+rUM5zAIBvAzx3jNmMZCkoM69aiaiZSF/
40cTWAKR+jjpPfVIrSs0MK5PD1/T1OW049IaTAnhsmNsju8faz111kp7ElYoPrq8KhnYkwYDnySR
ZLhXK6LV0PJ3gVxYgJy12oLpjzeiRIJQigrqpkkkwELlETVWqmynnXIxN25O7ZGCUaibR51JX87q
pemr4w/xv58BEIU3lXLC0h4Qsh4cmV1D5OWJGdlIQ2rjq8D9jdMaBHTFxq9lfqZqNTcOupUBH85y
QMnLLC6XJ5bokEvqrVKm1uNXGd6+c8nsCFoPYgfKDVk7EC/vIuIWT4/pYzeqWplcHR3WK4duy8ZQ
f0IturnSOLij10zA8G04pBkIgL6MhYHQjOMGCiqP5KXABXIcutqYOPqKKAvLA5NA3801dA8ut8tM
9mCeEbFL46bBWeBemFuQxgHg7wTSb5yi9hSmAf8WCrzVZzp31aO3gRt/2EUg/J8UXuBO948L09im
egJS4SpymwwFRIrzgNSbuG055Po9IywbRbHtBU7trtV4M0l7lH4EUOuhD28vU3QU7N1O/ADHzK0X
ypGxAkymbUBnw1pn8hfARB8+NHkYpnUQSWAMrKbzbDky99eBuAkHO8iC59UbrVbXdhhxX3f17OB+
BNjDabfhOaJQmoahxsmwW3mESKPDOCs/H1dFvmLuxjPSFdD4RT1Bntz/+BdP34rcwgy/uKOWQPGY
jI0tuVVDpZaqejPd7KpT9CUmSTFzGsLDGTXPevam+2gpeWsFm4MFUk8jeGCBZSnw1bq9xpkxfVzE
rQJZ0iObHIfSBHABpRDkC0n136dTd3IQOtulkrtVinAheAkfX9nRfITDyZkeVseTInVTfsEjyhMr
0QrChErw5pPOX2UFUOz1xcc7n0bn1FobNKn1+NNTZxz45VlO1Nti03KLKrLVD+uIq9MR/+FGVWOU
7v1jYq0ySl0AFOlwNl1GzdGV5AT/V2y9vAUjXdGkUxaBMweF0CE93co5o3LS737XVtUzstg5hYXx
0i5KXUSlmQok7q5oxNfZw2sVCv4nOcA0DUTkoxJ1wZx8UNOQAkNK4L+cISW1uKAMCy58gnAGFzuU
7zZ9+C8QzdT0AuObszlXsxWVCijdAvav6JmKCNEL95LLfTdUlJyfkS/a0AJlCjKBASyeGjUWenJ1
YEEtBP48RdMhWfVFxc9ZhXMS0jYE0bTF8qZZ/dUzwpQyVikLSEgvij9paoI56xansJRIMPYpEx1C
nof+1B2bcjqS7hgyWTTfutJAOsjYvyMNQPLZMGd2JBljiz837yISzAYUw0RIlvMSrGc1MmtoxAiS
ugW2J5lZ8krrqDYL6u/SVQ0MC31FtA2HxcrHfkad1cL8xUcLbXneKcersqA8ZsRjQnU6u9EBJO9h
FBu3jzQmYWlmOB7h8CS9+us1ojxFD4JoKUr4eAF1/tEY4lTJDarrfWgdAGb6HW7Gfogj7EJ99Zzr
gd7F9o1DFR7EOlP7ASI9lGAgJAvlYzwZjXkRKn1m1Q64ol/o6VEPYCWTAiGGh1zd8jyzRj3HuceI
PKN4ZL59nCRvQaUtIkzTFS7UtvWDh+QKeCqStghBGxxlS9IGg8zKXk2NYYfpuPtFFnKsEDx/TPZG
Z7DM4wwC8c18f1FyznSMjODt0Bm1Ey/c9k6nWeiYvqXV7XEw+zHmdKVH+i51JfgZ+O/Re+V3TRNb
asokt0NlfMtDbW1Swr2ac8Joxe1amVucOhvTWrHEWiVuj+Y66F0k4R2br7pLyxZnV8x36TTVo/Ho
ba2BhLhLVRA+cR6xiMfvvowa064BQFySgw2FS0LBjtA+3KOGbgN9bZv9vPd2T0AoYP5Qi9wPMFl7
wy3vNfcfW7bWMhpp/LAuOg+n0cmHZLFo8R9GnbC6TzSiZ9riTr6fPZJFwineM6ERyIIB8P8Iic50
cHBgdxokH7qHklVpxyaWF7mpocIeZoO6aijvK09G0Q1V0zWMTOQA/V5cTv4sqgEjir5GXuW62XVk
VXJsK6mOmktE/yZwheNpNjs3lluxPg73g4AjJAih6BwDhKJr4tZHrnxfdtFTA3OU4yyR/K5QT6/x
pFtRYy6l3sGrmi2Krzz10KTdshEKyipE/y/K6BZXCcKaT2+8gEGTURbH4qJbbOVibwBXYXNHm0ZG
xv6aIaGanOofBsz2ERX6Z45Xmrc+esubE2/R8OupzKycxDh8W83M9t368xBBZ9NU8jojFg0R8SOQ
FHqQt9oChAyzsCR37E5aU0v+K2lp8Ccw7jfcXi4nfgWgO8noCOK0onemgume+Vzgg+lQ891PXJQF
vQf1NnTA3VKaqtqweHDGDIl4svkQGKc2bxPOsdRiCCfKRrbAPb9WVT0zAobkpSUamh1T0XJO9ZkP
RrR+by6+baJOVqMdEElBTRZBn8lAhUy2EfmfMVhqANtDJyMJhwmq1kiBkaL06rjVhlcq6RXtcjjx
oQVlYDCi5Zbp7LeahkBJLbiYw2iTZQ393+zjywhHehbK5FZoYAJXkiTx+QTwq0jZu9655jv5zUPU
onni8UjQBSMo6ibr9JismJNrrNlXrWp+swQp6FMkJmXRL6L36veH57CkHK+A5fXXtnVdqjFyx3of
oFydKs3IBViEEayINrfpYTvbFJbVVTzRHMNJNMa7+BCqJedRWF1330wtxOwkzu4TJCoY0Kv9NwdG
oU3wLLqYWCnLNkJgUV/ovRm5q59XZoPoyjHR+1ULo2Dzx8Zq8yGXE3jTfyQWz+Rj800yEJAEuiU3
Egmkf73gwT13SVcJkTv70n8fRkH5Y+1nBOgreUcmzcRfGsc5r7B3pWsitWHCV6DJnhLDTD/XD0XT
tQQSG1dIhaUT9uniu+XktLF7cTWaWFS03wIvdQMTAgCwsR13pmYH2cB3NWQEYRZZJWNCqjgVjYSr
yDNnnNZLtpswKWe0QJdzNgbzijLPCsZUQoKz1vMW7UXL/3Werm1PGAPZBiGT76NdSKiEDp/sI6fA
ZpF3pOgl+2MOhS/zeRAB483DHJBce9hw+MjVN4p8XKumq2GHm6uIBuAlanaZCzP6a7IbQ+YHIKLz
vuUKh127V8/LiJt8i9vKSf/ymlOKg1XOvV4K/TA3H/a8at2jMERpqEUygM4d5pSeaC7//D3Jd2dv
35wMvPAxLyFHKrFt/NsuUw1Q74cHDx808oG7cRC2shxED+8B8g6t/vIip/iQ+5KUsm87z/vscnci
fxkFxV83c/8kx5IBA7ymSSCJe92++1lhNU8BbcMF2E0jkUJei8rS6jLjlIpzxz535blqDu2ObUOh
odu9SXs0bANaK+UWbSySpg84Y8IEkMTLy2SKh/dGNcVHvI0FDIABklpvCXQl+Jb4uV/oNao+RkUn
WrUwfuVBTNH6xkGoLcVI2w4ZW6HOCi220d38OeRHZiomALUfySFlg4vYQXdQgJlgWJdjaavC5cuH
tqMbYr2C0WyubNI21OvvPz7KKdpHUqPqja3BWZFYcCLWJmKj45D00OL9F3kyyGpXoxq10JUoP5z4
S/lPwYKiTIYXBhTdH1XiviIeTtPkauoytpC+nad5rAuezxcub2LRPNi1edb0S7MCPo7TTiyX0uCB
xVG0f+oN4dt7edKuvEfYEhrJcXb2U3zhEpmd5PqpbwpbK2F3ZP8jJ5ZkS2o/qZ2Yn7h6YaYXnV8M
RJVcSUZ2irCgCRE5QdOyWBFEW12esIb2fNxpEubqWH6DxVRi3Mn8TW3RMGNMqO6wmpIDkZZwHh9P
03Blffhgfmdb02EjaE627qXkIsXkaZbRAvq2TbPjCNfH40CRe2Z/2hf6F0UPotFj4KEnldR3lXBY
iF02NL7gRVdOAxwPdsJDHQV93XXv8sTJPEPrtyAWNq6UsZY0y4jpwHsY6ID8Wq4uWV9gvGi4Lbjf
hovJrQmVeAnNxhrKA+Be9jI+vSzyO36VRXWlPM9iEoeE5QxKA8oruUJzq75ZB6jSYcA/BlRN1uIF
lxrNgx9biudYr0kIepALvkbCa2FmP66A0DrajqDQO6SRo3yXXKtDPRO3ikUlRZXg9HK+j5ky+7Nd
yMdmnRqrIdUuqmqQX8f6lsp3D5zXeaOIrYT8TtC691sHL5XheK/kcNnnD9s96xpaeEBUKoRrsF8t
H5076Bmhd7AYDJTogK4txS48hQNtTM8rnwUdob8hA3OEln3B8GxVpT8YSYt6miRuRMx59QP6ta9z
jyJDa24rAe4tUBsFddqSEjMCKWYcwwSFkgDPJWPVzwpmipH4Yfq+B96Ul+4EcB/lkARQC6TmjGMF
Kfp62kkBEGNmblBMH13lDBa39uZTZlXrhi/MWRY+yF0ohs4yDP4A8mSjgdhuXTh9euIJ6lnvpAuy
4P8al/ehxalfkmM/NEwByPIKsOH0rbgvthdldrpzk3euiVZQGkP3aEPtSyF1221W9vct1Qm5HFi8
W1d9Ed/N2/B9CoWTZVW75i4T9HkmMZ5NGTcwRri/CHbxDhiWjxwYQKyGmoZ9mjPJgYy7yAh5txRs
UubjOSiRXx17F+HO2J7SfXTxNwlibI+O8D0XKGd0DR6b4ZsJAr3OjD9xxRj3NdW42qVVHw5S9+sd
YfVZyujl3usrRrHgzrD0ZbAryAuh1fsNxmMb6qQIljHj4nQd9zrKrNpWwBFQ9Wo0zHAPSMaAa7WH
rF3VveiU70YniioizH2wLb4AZTr+bl7D6gtEeaRFgPTKvwJyTapB/FH4cT+qOySNhOLwgsztUtki
I9Ko7T7XZ5HeKa6AUI4lWDk9vK7qs0pJDywFdmJVoFA8dF6dLefPC0pqm2cg1HeRurU6fyO9ZP7l
1TwDkubnBb2+Oo7TdWRn6XFbPmjpZiXLZh3+orwPjHCslUc1++Mm2TMe8XXFiVkf07whY/WdMPAl
DxZEx6UvMZ1xKg0WLubXyaqgqVDuw12JG/tLcoQKzTOu2IW4hnDlqTBxjWJzl+KGa1atkUzhAcfk
W8vK5H1xm0wz7qo5OL2iefh6jZtfY/kzOBl/8KDJ0r1wtfV0yGkJ5QXzgmAx1E6q5sHL+VUGvXwl
4CTpb2rJ9CsY3Tw8Arc4X3lDBL6dNaRJy7g/vwUUwfBB6DoTWOqmpa9JLX0nog+UCoLVIqAanPcT
Ouwwq8jN3sH1utlBphKMCHlgwSeg6vX/D4N6zwV13Zw5FuC7f+fXTHYRhT8xFc4aXa5cQ9cSZQrv
SlKrg6O2N1NtOiL9AM+/jsI1LPc+Bhu5GV5Jd1MUT+iVXiT6wNi40ysemPj1tClNVrqAoQdoClwl
RJ1vwiHtM0D5uakYmmYh7hrHtk1oqDvjmTSgDro3iL2ITifkOC/Nut85ibiL2A4Xw+LhTVnP6gtO
QHC8/LQf1AfySG6NFJfvqQHUujLeDwl0S9k/IyidzzwdGYueSQAPXLT4t8YLtqhaD3ygBx8HW/CR
zIQeBzXCfiKqwSe4a6/1RRi8PFJQ/MIC1ULGRalrosmrUAn4Mjf2zE/ELqUIVqr4l16OPbga4WAM
ZE5dq5azj1RqAZGcXezEgG/pHdFFXwDlwvagv/mKwcbMyybs8dGL3ZIp0wB0xrjmj0HkJOiwbbyb
KngH9eF9SsvH9Zu7mvRb1C/ydvX08/PIPjr8r3q3AVqyY5cdjGVu1ICs4Z1IHdJT5SnjdLk5uzKf
AYcx0dc6aXjyHVjPI0kOW/NsLzgSR2sAXllzvGQBpq/OFyER/hvY3PxTVsllk/7iLhioaWWRRY7q
mFFvPC3au818p4eigR+2OOz/Sd3k3MHVCEwwVoj0o2Ibp0+VbcJ0pXQf2z0zquehYERQYiJowpVb
4urBgVn4lmh/32m3zpc8awq+Kk8lj2EETXq6L7CJVG1OztB7UfMvwuuG6VgD2xswLp19vPJ+4X/D
POsxWwuldhlybMVG8cynnIUMMD2g/+lcI6TvB/UYN3L30LwyqsaRlJ9iAt79N+wEHsszFcl3EoX/
Vhnu1AgAKEuzndRQYGro/CJs3jfeULfnADZ2P2PAZX4s5l66oa2d+bSEFdoVKFkqT9Yk0UT7s3eM
n2jnTKyGvikryiRxJ1hNF9ktJOlLbHgKhvwDRfrt8WnbgX2NIuhJ3hpf2b1/ZY24pNxkDioW6bOc
ijuxUlUVgweD7z0SgvRC2ij7SQAPeZAVSDqiLNMitFfyi6vRXpxZkMpSKjyjGgk3LBG/S6K0kszv
lLFAJNvX7eHNiCL3Js+V+Irq1n2oabllyxO+7qe7Np7VZBw3WdXXKngv2nNuuK34GlVsDeakWp04
DfAT7BPIJfPDXcNhbVvTKcLqYjEbQ+uEkjgSSIaxa9+dSiXy3esqeL77XT/KEfCfrMezUEc51H2O
GPQQotZzQB2puGYLY/8LKHzrb3NZDuNKuLLvN3dqd0G8tEEUukLwwQWMIArblJR1Nr/eGmrXeVPO
HtIDxBwaIawGy+8kJm5w9eXQXJT80zH9ilvNIAQNFsCzE2zsrXAUIdRZrR9RuDCQ1Nbp+Ag23M7R
bvhtiaryqgpBCdeQ/pxdKDQwh/iU2OMlFehQuBSPaYEqmrNDy13kFobpXrab7BQeGQ3ium/tnAw0
u6UIQ3clxi074K5LsYd7y1VhrlCFd4xXflpgs0J4v117dvkiiRsBrwhissnW9EDpIZ/NpSkiL2s9
OM5YEBXYrBM3ly2VjHlJh5DgpF1/AQ03H+I93s8aZHGqNui8coK7M9Z2PczYLxt/Hb7nzb5//pg6
H51GtTBhaD4+WNtBkXi2nXCJi1PQWaKx7gC5ezhYlzEhq4ueb7XeTU9JHqtzb2o9Fkxo9eioUEhZ
ljsjdsQdJNjY0fhZCi6PSg9R4+MeZThK/EGcMGxmMQFM0u4aiwQ7jm8Vk2boV2sFCJrGJWr63BKL
I39naSDRHtSKzaKnRT1OFLLUp0xSAM6814ZrxlmRMtcvnR4wmWvqfzKuM3UWYOTmmi+DHp0DU6HC
2wQ8BKElVTuNgYagWL3CyRYMEQLr4dsLbJHQnWaS9hwbDcN1lWmyYCsW3VXoSKzSf+YH9aqgaEbb
tzifQd4G9CJNwOvssPzSJHxioDIn2gyq8Gvky5RC/z+/ag+RLIpREx12pVEoyfXd3kmk/YeZyVa0
otX5VSnN4d9TWSlR0F9WuM58cHrCJ7ZJ80b+vNnTt8XSb3g4/j0t0UxwqsK2wuKaHBngAAZRSL3+
kwD+Y5CFQgnr6m2uE2CJfPaSQGRFAuo698/xf1nlvPsdojKJxApNRXDzKnj81rA7Cu+4sBKo0PrK
K7He6u+Cmky2atM+5n0ZlZSR1yvSZEGXhJbsddhXGLFP0Ay577vMqQUha7S5rQ+7VlyadRApgCnv
uaTqeoNX1acDzi2UOZ+65XaCcbsv9zRCjQr1Noo7r8dfUTLcLqFxMTnz3RWa6h/iXV5tUt1DnmBD
h4pgmpBvM7g5qjEWixfd2t4q47JMpDzJPZu+BiqqwewWUliD6lde95/tWM1+OiaMSwD0v5ISpO/k
5qIIG0hnzn1sXFrlS+/ZVSU+VHaozEuQAs61vd+eqUUee+CqewcvtYjdOFpBKyxSoUdss0jKFsJl
oB6IrND6muPQVryGEzu+JoPg6zSo5X9i06tKfQbwQfji7Zr9K0lOHL6HaJ65YvXpRHXhwC3wzycs
5Pmdi1AScu6drR6SToN3Kiq65VbdWW4pNGliDdrN95Xl3hhrEBKqLhTUQVJEzK5QWvIfGZ7VsHWg
/IZJ1LJDd62VevsB/uwknCHWIBAdL73inO9WDu+cml312PaIwfrDvfseTopZPsf26MqRqSLbVPD1
YTP1l0MfBSJgZchHOlJG3/DH0sAFWhxlQG3WmWQImZ5QPT7cD7miACWw1S5fcPWqQ4b3yWlM0MaI
JZYH5XjAdJM1L4H53HzI5U4S1ls42q5dkYbmuBojgkD1iTEKKJYbbkhVcxvMV+lLXgxxagWgbR09
LScac5tuU4XLKMhuogf0fltgD9MObpoQsvx2883aRca2NJIe14KNf9Awkd4Kxn1KxMiuy/8fV9wl
mZEfjrjX9ZHz91nRsJ+u1GI+zi9GMwlL76/e6dEzT1FzadnYC3VJK6aq2/8HSfpmwlVXeqk3Y4+N
F37al5OVCgAQQliNAKYEcriP1hrupCTASN3nIqEdQCd7PfAMtOxfXQXCXcY8IB6gXoetwzb/FBWT
H0WCV5+uoVQKlvd2qpe7YXuxqP9Y3h4/slCA0NsZ5D0qyu7MU7cGm96HlcFCwtLLJdXQLRzazqnQ
Qw7nlqBGqwgmpd080XiLsV8rUtYmzBdOZPSflqIz2ckhIzfQ/HkUEq+rNXLtpRApQ5jF89jjmQ4P
Z21l0lID8Zyuc23x2Ykpq5A7tez4UAs0db5aCHKg5U7qy3yf4IcOq4oJ7i0DUfxUX4b1X+ibLZYq
dAezVhk1+t6JzB9aE/EJuVEGkUXRoYsmSCWvac4BXqXwOYOL9MpRRptKSnSTz2Uc07cY8h8/C3Xe
0J1pbvXTrtmdT7fNTGQiRQpEdT8af1Wj09C/5zAuj/mTLMjbeDuO1B/G9aZ+YV1NAkuTVAgLBqlZ
SLoJKiU5TeK3WogBUo7tL3AIO9XOzKzgoDIHUPt9H88lN7O90wnG0TMsnK1tGRlKf0PMVADTj80g
YECG/XU1RkfYFrrmkIR0pqFyh4hhuBJKQNmmXv23RAuxhURZsXkAw/+s+PfHgA1t9L9tmbv3NYUC
I6XAfjJoAvsDNRj2d3q07L2WMrrzbfan/o1Ndoj9gy0AMZacp3kMs1flmvkMcfQlccjE93qUWZ6c
AtWHYFYkwBwoHWskQmRTeN95ffMlV/+q9vQXAx5lGZ+pfj6IDkQDWgJQfEaH4tP1RdBoX44F+KdD
O97kp5B8+ubg4IC1fexiMQ/nDoviDySYGJ+sdjvmWQJ1csqH53CadFmNnWfn7E4JLbAGTwmachEX
lTYdK4Rtp5HSUp6qHm3IsWvOWh2aQI/GzJ1PEUGY2qzPwKtRqKhTIRjFsDAJYGUkqiCxtOY81cL/
RJvUUJf51KftruBAogc0+kkCWqjXGP0LXa7SSvxV3KgfOrXmbwYZ8ursSRsLuQJI2TL7UsbCDp7b
5z2cBlbuMzMxZxH8Xj7r4a5XjaSfGwhOylSAhxy1HXHPw13+HmQnXz2SDedYS98FXS84Z+gAP+EF
o9X5F7WTVW6asAdQNmv7nfxx9XV99m+zi+6PkS8g/XQn2A8JGdtSnVIPQeWXZejlhbht7d4yCoha
O706njpQaw4Ki9GqehMg/kK0tGrNcFfE8zVGZl7gyLQ5eeyic4pzbUfUfqui43NRaYmPyC1xpVC/
y7HbwEGD89gn9yaYzPSFx5TQWrm0qZoG72+TrNcAmfUZjhIIMky0Y0Gp0XU9Yb0NP1Auh7zu7mkS
SY9pw7rgujH9vks9L7OeLCYKxHmlVjKtAyd32XmKvhRgIz87vQ3AGUVX//rerX+oIkXNjSHvsMeZ
D5EilOisEZWkOuHmq+SQhWiUAoPXTJEY4QvQbC7gFXqgJnZQyhC5t4FprvKZ++UodbUxsgLsi3y7
rxJBqsGFfuUj3bmjpxOqLBkctNdP9pfvxQgJZuDtGcy1ZsAHrxGOq19e06vwAL8U6WRi7otuLqe9
UAVIG87PUQ3zVwnp3ayfBrDgZbzdVPdWPODTjvQ6B3SjENIgf4JxqTYNpxLao3qL49CxOCXOnPDq
fTAAHKAMAgoSS/SRjgl6G+BbdeWm0XJkJbaOJUDgSLXJMBCROFK1Pas7umi8dVsDbANojLFIqdeq
ZrlWZdIbKTATmbXi7mMMNtkoIROaW7Z6n1aCyiDu/vBYZE7FRK45jUXam7o1QDdnmzaUizrlI4RS
Ivy0Ssr8eTpwqA8LDsYpjYNstGj42w3m7kcJP/90FUv06ayqtmXLzoWpj+MNjIrg+1dijItr731M
FEOLDbj+z7qFyph5en5IE+7IggboY8GE0S1XE0CQb4pRBg5IlaBdI+bWNCOBVwDlwkbSbV6Z18qG
iuo1SB183GtVXKWUzdhVLXJBHDGX3rPinID71q5OnGux48fovDjf5osicKqA2ljEKQj9Y7aIXgbf
WR0EwUGXFSHoNZF6SY3e1WsNON83z53EquNY4aGly5ttJetBuh/izRIR/Vo/M8FOpGJd9CfMR/IA
xfrT5wpTqG9I/2sunAtBLxWsI6Nh3faBiekVOaASWDJ90xfAAjH11/gTnmC2eFer+XceKj6+xgn9
P9fY22iUClf/am35gDqDKtexMi5rchIXk5U6HXD7fV8oaPNsh8007wM0JnDtEqlO4af+UBGbklf2
hzKTzpeBOcaZi5dGFk2Wjfu8vEL0U8R9V/XvKPAfpEPaUFnVDR+Gh4+fkdZrkfKgoodN/wWVxGg9
cfd4TypZyTDnlkKfwzdhiLDHo+nqil+xXmiXgAZeyzeE34LtBRFkLpZ0D2i/X9R8D6IfdpBgI2Pg
3ko+rQDQj2pVOxRNr6NTP8324tAIVW6vrVXGDtE2G6tpWWVf4+dkxZ/NtxKGwKLih9chX3vAxPJv
ticvYC53jBK4OAlkSplisqRWqz9RMpFfhISmaS2MJ3XcpnDCaT/6VJswIITxdJuoujjbYDEI+uUx
qbxMAIPqL38/U4bqyH2m9GekOk5gZrIIIO6PjB43eqWGwnr4q8uRgiadksMwryFhB2CULNdSlaPX
mdiCRwNppTcN69Ybfi/5kC9EcB4QwqA9UgVMDvAhhh7J8spMTAs9/bYkjyNZENdGEIvu3m14QLwF
nj2Ic/95S0ywizJ/+Dn7rDpYC7gIFYA+CLYWORpiERws8BMTl/LOagCIDoRGan5Y/b+p9AA7jl+T
4zRUUZgHysvG5Ic11sUWsen+ktlc0ynhho+7mwOeqIPVzaXjKiuluelEgkCEodtHZJUJTU1j619f
00tewuq+51kEDUkXF/ipgYlyinCajA8jHMftUB6TjGzfTQ1ir58l/wAAihJg7g+uORYU3DlTF7nk
KlFNvHdmWP2ttvNNqllbO908SZHK0P2tgiUET2h/VnHd/CeeQzYepybbbnIGOjvfsb+JBOTXqD+1
LT+5H/oY4o2NmbQrWG+/vYLTrT+rLndBAacc0Xk9k1CCD0s7GKZIyEhFNZhXORy7i1zisklaaqLb
iGS9rPpJPhipfWAL8IKnhCCR46pbdkg4XyZACWmjFo9d4QpUl008dulHnFexC01NZIUCxfKo4Pnu
XB/6E/wquBUu0P6knqKVOyI/++G+KZPwu37eyPgVovpwuVA/CpDmNcXa0U/qa093691IorKoYPtK
oadT698QEZm8bPpeKMX0n7oxoYNbUWUiUPgUM6XzUKN5AImSuI/vmwtU9gM/PsjTPlKeyiJU8tlx
zH4FPLSbf0cmBb+pBGUf3ijKbn9BTTUpx+7mTJLB4jBCbl95ghtdPSaQvGiBd43kenwtPcayLl1P
N18aUoR+ucC30Y64+JKCEPtEicxfFhBhUS0ygV8nZrKgbpBZ+T4Ze1mXeUqeHYRAg2d5om3Zf6JX
KDAoWVQA7ZM5YEtZwfsOHquMLW6aC1fty1j5s+bbl8gxtX4IYeh5ao1EowH9hXJ7YaAE6KdrPXrK
H+kgP59NUugL+xoy7Cjsx0HyY39jgqCBurauvHXg7PTWX0ljrCohezlROLY0FdPQPbifhL45Vt+T
qCGaOfzEjNMmTiV3GzrvycPGQOs2EUSvPW1sXdPr6Bpm8wnHxkn3cnOZ6dffkiXKFdsBrkIJJpl8
Uyhd92G/P3rCC0PrugpRgN+G+uTnEMCvnYXY3YUeAei1KCDnsO2mbFShJAOrCCbbp+q9dMu/OPQ6
OIB/EnsCmqBnVzP6maAigCKqJXI05/P/PHoTjNboCa6cAAKsyaUEoL6T1X6h2KF9/3OUD0fEl66O
m1hIPe0904WJJVjaG31zsmCixhrXt6FwSa8x58vul90AbHxcnYsIFKShKINBLBvngW94/UkmyTQJ
91RdD/q9T0ydV3Izc36KvcgixV05JD3qfgTK2xUpkEbs3Urb/NVGvphEjGmgxP983rg7tez5Uf7m
G63d33ztTU6pvJCKVhcSYttsSKaC7lSuQ1p10QH5Uy+yIAm4P9l7uKN5ya9z7+AxdgIPkn0BBdqY
rHDsCZRWOkkeaXsm/76zsBPEvqLyh8M7MngkuveQIxB6tW+iYXlFpB84wwm9avuBnQzydu9TwaJf
f6t+0Q/gaTkJwqryQBp67EwfmxMyTZsI7qByEQeG5iT9zFO1LbKU2qS6MjxU4qovZrdlb7H4yAlD
B2ZmCDeJDURTTza/ITNmVuQBEq6HZROYLLzYwvlNmBQfh97vW4F2Lr20GA8Xgm4+SnIX5BhwkH6g
4YtRByuNPy5MbNJFNOfLZTXklFFj/3auGWBFetQVsmrZyshb4PLzllCI3Ey2JHWcRPGp+4jdXtDC
Qsrnw8iOnkMEa92piZ72VohzZEXcRNRycLfXniV3P+Q7ooSN2rMH/ZmoLq7LJ+NyI6qWunAxbu/P
WLDmiu6pYRQTuOxNEVs/6n2XLGZLhEy6y6S5kpYUXYvMmRp8oKxLzMrmHQXQEyrBHGEDhKWq44zF
zL0aKdUWqge5hywo3a91A0QKShkddrLyHnLD2+BBOsADSm5dd1r+CQMlAEBG3XdorYIKLWkOSCdm
yZj2oCXzJxPEavWVaWojAtdOzXZEpSIeTNaZnQJj6FlCb0NSBE8mJ6wlfrqdYBAgINMw7W5zLE/g
JnjfHTSTkY33bh9KZS4Ci18Zc1p5677WJlCPpj3ImhPV5xXve5yP3BlTUlPS20RPz2jxowf2ZCRk
SOtZG9OBgLtiBc5OS2Wy0ex8h4mCGXzcYkpblwTBRamSep6ueATnsB4x1i8V6F8qIcv3P9Pglz9u
YWHH7BwGw+rs8LyCBHUqRn8kbq6+SdYE7YU9aaTiE1lGGqo6/jq7AC18yhuxkoiopgG8qkRBD4DM
RlfzhejK0oRnw0pGwfvBdqvnlSYvQM697IYGnXbdZWEno5g1KdIgErJAVpbxUEmIPra7WCTGOC6c
EczGigXKbpMk1CKFmw0Xnq1QVeGerIuB50Ixow/YBzdOBblpKao1FwLN6CNHDvnn9FcjqLdRMH1g
vqDq6OdLVGmdI/+UJ/8d1A0nRncAEadC1/CIFDsO4ioVS1ZXZOX6LJ+PElE3nbYf/7Ui3upC3JYE
juK8bRD3gURrtTiKGmF/shEuMuVexR5QX2Jw28BZStuq1H4QlD5OoGS/b6cJCwDwuVBKIUU5TxT3
xZ+E5fAw9XW3ddqfR6761IJQbILiHDqxYC3UGDkqqOI5alOahOSAjV47v+eSwq8K0L1PPw+izz2U
yodZT4HxAwxN4a9mBsNa4kuPHm/a8sfqVcDT98EPx2S9i0mlI5/T8+zoMNuyqzTAAeBBNqkj2Dsr
Cnsa1C3SQNjJgC4ifegY/9BfIiT/nuozbO6p3XnabO+ng1FJ68Bp75VQipawhJttoR/wvaovGj0Q
tfvNKNu9XDvRPQ2CfxKfrDtR0szxUcg3hjk+Ua27JgxvUa802d6MzjAXxGotrQf58+Qx8fMItxxs
tncAi40zy0XEfVS8iu1HDTbyE+wgGUF84q4NJimC89LWJcn0xzpwGv0ON7GsQ2+7VC38WRL5Keo4
g+VoHOv1ny86nFjmwDBTanHxaT82TEgKzaJPqYUb06pLWJgdcF6OyQPUlM688ISNZKWxp0sUfMTV
mGtXzl9IVBRQlwKfr9c84+iObHeR1IzOqLBkbqgYSiPy8qng2O3HZfcofGbQE/0ykLTOoNzpoFdE
b41LgDU/w221yvv/aZ6aJA52syLh9A4AjlDcSU9Qx9bduWNcsTGMe1qzGptj7BK3ELAA+Ihenn2A
+JKjBF5Pas1Lw+riZ6gYqsyGcVfj8FgcfkBAm0FkjHYlRKiWZZjnWNBNnelg32TUEpWMAx4Ngmkz
DTImU5vAzK8i5JHCK0Av2rRfMKp7aZWZU2oQiSAUxu++4XZ0m0Hn4sMh0/aKW3WnyessSbxnAnSV
S5kwTXqrL9V9aCIaNea++JG3y8yE9NFbYXiCFvhP7iEw6JUNam1f5rImpeRxs8IDL9QsvtEDTBQX
T0s0SZWHdARJFOSoNEk4cuL3jYQgjudXrNOSKoEcm13Ri8nbQAsxMv1reIKuUrY78uHW2k/AYiJL
71dr1LOgdteNrlzBus6cMoPQoFTT0cFxWT+dDv/V1pnjeoEZ5t/J53zZW2SIvC4u0I1+y8YBbm14
kldUMbWUyP212BJnkChWRw5jZhpmsnRiuWo3N8wDkKV5wEi3E9OHV/6bVILMI8t766WI1MLyKXrn
3L58+E+dvKiiXG8/L8XH65y++oKO8JX7TWbVbArX6eLkX6st3oCBvrySOjbdOwFXOixOK2SZXYlR
OwUlmFoRdPRsVQRwOxad9WS0wV/Ku6CrmD/PIrYA/LSPTAP0We0WUSFmAcw+iItWvPMF87++zeoL
6KkfmK8xIef8EoL8j9nvYQ2MPDaHdkgH8RU5qt5nlaKpzNULYUUK6ZhuwqLYMuXfkaPjPh1KjkPV
szxq8+o5DiOg5B+zcenP5V27FFYXOC1Z6OMdqIUyOeCGrl88wo+I+XAcwt2id9PBzqHWqtpUdMal
dd01biOFj4txBRUeG4393FcVu93GOob/YeszzPt0QoONPIh781gapbXn07o8osG48YJQ8HCbdUm5
uVpiv3kKuwoJUxg/3zB+q78SRjEHMksASXwmLWscjOqQENT/9sHCXcsIl1c7uMUtvQU+psDgeEW9
jB0/0lNi9Wn/ggEtXyayH8rjX1qt8FsjZd+Oefa3T04rUjGMj/b5ODzcBezUVWdRiWyT9IDgAxOP
9vYokTPeSEbKhJmzTjNEu7Ufl9Y+5K30yZzZegSwXdWahAI2OZlGwwwTYMaKaeCQvTG5VhQx/IhI
eAgpLiSRxAO1Dv7r9BZGkVeMIXotp+mOL8sJs3LQ2fFY+47m2jVD9qFIs9Iu63wXqOu/DEnKE9eH
4egrSOwZUOP5Nz1rLrwE8EgYB4aZPH6w+Vqvqf0HZ1/5CNLScih0gjRm7jEw+24U3A9LJND/fSVF
+BwZrpV7qW3CtzWojfaUMUih8/t3sXqxbThDswky71LzVYcnQFwbj8zbxjuR1ihh7FZSG6SBeuTX
J8uEgKTdPiQXNbF2JgZWJ8wmorbIb5vH07t4NJmjCVHQ/UxTbUmr1GOZ4xrH9yWQso5W2pX7WEAD
IE9ZiDhRs5khv6HxssXRcPvv4DaecuNZ89H/6gu6nNkAvYFKCnPvLE70cbmQccQwDdwsiCKUrbSD
7pkOMTBario+F5zrZsZrKjEyCUOsm5bEGVBDPdyuq0fLOq7OuKZMkBQyE1pdLZWyCWXhF5JTPWdC
IEhdeQrInTysQR3mdjrZR2oaaLflxS82FWdZ9/SgGV2Ay3L2+IU65QgeeC53/qJXrElZcBDu+2n+
QL9DSskC0cojwt71XS7pIkgpHg+L0QbW5RrHpgkdzWcIwolSg6j84M1SwLHDkvRiIKfLvA/B2OXs
LDIeJOF1MJkPhdw8y664HLZCyUrJ+Kpg82uXHy/56sd6zi7TyvCziaCNdRw/9Qgz7H2LKm2zubrD
rB8fwrjTMymHIdvjzij8nAEDT97heZga0FFS84inmnHXpCSQ5WfiqCFRcqw3clO95ReNspksFKqR
dDZ47YB47iFX0/NcQygFPx1GmQy5SSBR5dxKNV0/cN84yEEzoFEWpt3hquID5rOZuMYam1aDCcdN
xsdhfXsFS46AVpZ6cGolZRzOKUCnqLlKhktQ5Ypm3Wrn0F2jlBThcmOu5Ci0vj2VV49nv7t0IuWB
Z6ri8zWBTCN6x5CF2puWChby03q/oCfxUx0x2g/+uE3ZEI5UyIntZS9YWQi2zV6YOP+Ly5i+56yY
Q7KmjG+kdIv6gEl2hS8tpcuchYfjv8SPdNaSwMnluaTO65UG4Y49Zl356KEUJmK/92MqnhE4Hy5f
yyWjS+H9re3RQ7S1tpiw3Iei+fpSY3v+dQI6tTlV/B8D8O4d8j098dalEf30zqLWtNwNH4zM4IlM
6cL15ZmLsbrsXOhz1u+lJAtg0BDdeYFMDx6zVdcs4NDsZzz6bzLl2BBnUnQCOXdACg+dtQyYHZ5J
mkMTIGkvm9c3cDpD+c2xNSO6Bwewb/zzKz5cfwINgywSxFiF9U5OEoRAqKa3u+1/kZMK7E9OgCf6
XH23UoUTQe8VbNq49yJ/rwK8He3L/SAwgqgPjfSU+Ss/2DU12sFLUyfPusERuX3mfYDWXwaoXk3q
JPI3tdu40MnPkXg3SzWv7sBDpEJFjcjjjID16hfq/WSt0HEKG0e78h8JIPYspPiZ6suWVLQHoWvV
Tgkd9i8Z4dQFFEjFQMVDZ7zQGppHQYlK5om3gRO9ftOWM2QIzyEIXlWuMKOyd8CI2XorVuwYGNAP
8vaBmngSMhwZ3J0l9OUHMk9HyQeW6o2p8sgDTuwf+P4FzjW7U+NeBpjAdZTXtMxMD+psouCGlhEM
xavaKn5IJ4BYXalcUp1bu7lpoXEq0BsJX8jN5dyhLXv7msodQyPPcULCjZHmRm4nNtVleX98NaXa
dQgBd5Jh4KFW8/4T/Q45SxXmrfv1bTU3LrSkI0g1sBUzLtIel7rwB4Kc09L0kSIvMDQ6GYd8L83M
MTsWMGjS4+dSXqSMx4lYSPpnBww7TWN/XSlCpvqydkcPic9IRqG8O9vMgkXwCPDW1SZk76Jc/nHY
vXkhNX0iGaQ+E4N3C0GxLgPPz2+oS/3NiRl1bwwV9Zfpy2FYX7QlKe0+bXQHpjDW1de14+Oh9wJB
M9uAkN6msHtp/sZF8q9jCEvV0XxriqLYOpUCU0znumyZu6aJYB0XHkOEDkm9BLu3fm9MGBxJAEqF
eRWQMEo5oAX5y2WljuHVf4wv3rT7uLOJIyTofvonvJwv5z50Najnw5IbtIi9yWZ79BAt+Vtiy8k+
/RW7+AYJCv9avOtro+gCvukRv9iKUUwzh/5o1wmjJegVZ3LDYL2WSw+k1Klt1p9f6H7Yt7ZzU0XE
+Oey+klf9mHvlHTG/o6rUbkQLpdHYH6GMhdQ0WE+MOe3zmfjVGMAYf87DkcMX+iaQ/OyJOJlhlXE
N6cG9pGoBHevEsUOgNoumN6DN5EqECzQCDTdbJkUpGuqGOCaI4gqth/RPh+1ILKKiUic816eXJ9u
PsqYVRgdn4ZMoFUECnj05lJpNX4yUYWleTsDp230YRSn5sCsg4za+MhlAbVkFJVAYTw4bbj4S0Un
g7/RFk7n4/BTBIqsyv9SCc2RGQjS2O3jGHZ//Ri74RuJpfi7+peLZizj9Brj3t5WrUn8R6nyI183
1digIXNL3wwUGNljN0bNBSpN1Os3ryUaHlyy2T4q2q1hUSCoDapF5tChLzoFIbSA/fnAvjI8oUCx
1D01zEzhPQLlvaxguJoWl5BDiHpcP+G9UGBtQza4ZkJpUFvwXoRF1AKL3fDHY0RAr1RefJ2Vrb9B
poaJLSC6UTaMSXjieAY0maYyGKMEC3ku/i8+3PzyIqutZvLYKihvPA7vfQV3mKBgVRZMWTo/+dE9
pW9Fz8saQIRqMj/J9Rv79jvzyRvjRn6e/XgwgLoL0IlpBmI5em9xwYeRFmvEopnWpDyanjEsoGI5
3EJ8bc98mOifE6E2DBZdbD34Xln1N+dempl/WzZo5P49RfgSw4g2LL+cOJbmjianY+xS266RV7ro
AKfWBbDoFy2PA33luFiWlPE+MhmSi/ZmQWul7vdxi5w6ILoo12WOUHu4Tc6qjJGsGlKH5Voq40cF
CPEiJ3zf4TG/hChX7DppKlxDy3IncEO6Le4GoyGXTUuEx8JKSmjbWBWsxn71utwH4XFqOTII7huo
AUZyKels/4SnP+kHEna8hBaBn7r2/mbGqRCvnZG07SN/uw6KJHzLvwv5N9rLhQ/py9/A9yN7ZRkr
Lp+VfLvkWEjVN4QqDWQolefJK54eaYL/k+1RNTL1HfOq8HgI6/YiOx7BnwY8juLPqfM5Irm/0wXg
JREhjudDRT3yucUFDTVNUPus9FCrMzFzpnZeDgDRy3WdzapkPH8ZVctJSYvEO6MEVxk5K42NI4IE
QclL2yXAMkbMeD2DOV+XWSLTgQauAz4v1RltfoEqxpid7lpk17rE2wzrYxUHOFnVfQ67yT03Npsg
wJIlkrqokf88yF4U+ASm8bdFDwTwhg+lN8G64bD4VsbqN7rttmO6ixmkjl1/EhKnX8Nt4BInu6ZI
Rdro5Ks29vSiXxs7iD5loHBdJFCJYgCRCVSYW/oEjudk1Vf1cCZz4gYFlyaSbMFHQY/nqZXRSBlO
klXBtjSLyVc2hhbd6OWLt7vQbpmawtVr9FKA93Tllv0cB8ms3DoSMBqlHhUFB/JcHVm6W8WtseR+
sFQ8KvdPGrapLTLGc83IAPaoBrpXljnDv9ua25tXe/Buii+zpaV1MXYTOJUQOjqf5S2T47WFpsvv
CntQ4lGgD73A/EQSkwKibCPsVM26NudjeD2n6uwXaqM8tbseJ9f8ry5QCNbbjzme81BUU7qGPiEL
6YZzvZVpExS/3Ru4j8/Bjro0XYxjWLnLhZmez0r21JLnDFXRJoXaYK10fcseB/H5rghLtICa//IE
If+++Aby0TVBBx/tEibjWyHzJ2Hm8YIx0ytnqA6+2SacM3YzCnFGggWf6TYH+kRUY2Ulu+6d/Q3j
wWxUDHOY1cFeXIxQsI0RjSq8uNmlIkFijviio8pOQya67kXzhjkM9ZpdFtgv/nasXJvfDDAi0lMU
trA2MK6S7VF36z4z0pFb4rnEN2K+x4JDhsrF0y7W/vhh668bv/bI9cRGgAsPm1gMY0zl4h428Rky
jciXUdTyMg2n/pES6dPfGeiAY9dhFW237DGgMqS3fxNsOpVMQ9QOUJL1eGVawfBZd3Ays5MO/h1x
4PQvVNkGTmr/vQEX/xQOggMbgHLBK140lW5wWewAHnAFY9y1wdGILBnui0LPuKRTxZPCyN/69T1Q
XJaItrmHEPTBls46c6r15mnsVWX5fMS9WTw7MZCxqr/xckoEPyYWPIFCmthjd6qZM8n8JFw2Q8qP
OVSAUjLAc/csUb2rydx1JOBPcKvGXIFgoe8HiroqfGTcCZcpKAvcFXJfPp8QYRr4mkTcQO5dTDiR
Z7npdj0hhV7RcpPzQHY7PSqb5J6Q/AEUiTq1txG1wXIQ2ZBmXrhdmiXCtH5vRlpUm41J9qAe+MD/
pR3Zf+OLVYSjbNJvQz3+cTsqx50TfaFHIEXrugNkBsklDVyd/FN7dz/pqXx8ImkGB82ft4COm4fN
Rd+fo1/QSJoxyx1VLdZVEHazH7JKIq70n9hkiBJnnVwQRA9oX9fp7W8SVn3BQff4L1a75w1DXLFA
LrM0VaDinSKQ1wlyqI7pkQI99JOmd0tD/y7TIAoBARPqknKuBlARTad3AgxOVnzSSrCLiKyAkiSq
0zzZNiqWjkNH7E5nWrRQl6g6kGEFAJF2j5xjeBy3+tQKbsmWfsGG6vDgzeVRm4R1YcJzHk00PwK3
abHs/mp5TGcWrm+g5O/VyFTFuDSG2s7Gy9gpeCUp5FETmFJfEmNbk/P2XTWCaFy4+jbO6SdISJf4
7dt9wsGJHBctfcstuMjMVg3t+Yc6ynrwzHICxdgArVXtKFD5JZoWdSw7J2grIHJmeGnbrBaeogQ9
6BWfXSRVs1GGIwHh/kwJ4YU77iVnMR5t4zmSRSj7ecQxTmd8F1A528l4VhbmIpyIUk2QGeHumUvY
oglORi/qgQWO7iTicS+5Nip+cP+WIMIVpA4xvJfm0nuELf311ac/IJzByTj1ibc/MVXPSZMu24HY
rQQ8lVGr8fSLtCeOzllWJj9IDt7dBy6Zgr+dW/MnlXmXd6zQeEQpDCuRUWDPM6P4e8sRO7lyAoKf
OFrsukbYCcKI2UNYHICyecggfYYhXU+cAV16B5JCoIs9h1MH2klg39FTrsgAokXLDfkBRBMBPnb3
I6S/CGie1mLlQitgS6+Kvqwb9ew9Z+60jUbgmrwOHksebRo+ojwVoEmPZe6Rm71ot1tDHO0t6nDv
vRtvDif1IoyEUNzfj+8IESS1B5Dno509nRpk5zcJvf1Y1xWZ8BKRs/PcMgfj/i6obQ6LXWEuQmEg
TOX02vMDjp22bLx/YzXeir2p+4twudk4uwIf+bvR3oFwTyJR1Xt7Ntcx8lMviPA/Nhc4aTZRFUWu
P3w3zpv5cPPMWsk9accF8Ktsy+yGyq3lKRXFetBO8vrnADYPSQ2NmwerGq53SMl3PPzCIR1pRRLk
OlCWTAUNzFroZTIS3etZTRv3OCSLOQ9nULbZGw67OXfjsXxMm84lXJfk29D+ZxbkhZWO85jQ8B5W
vxggWpWI01cEEVo7TDDruClaC5EoWMMbclyMHb3XHTTvan8ZdDViZddr7EFriAcGK9xGoq5y1yWW
ItXjMFElXwQeIfw2A77qDQLcMqfYGioCHi0X/xfrGWlzaI/1L03n3csMSfRHZiM0RRjM6tQus7Nx
vSaQVeQpjHYAjiP4L8wICy9so8Q7fRvSFL7ybP8kOHJ7biwZ9qvHjcUY8fDv2Ms/HrreMxPA3C60
7HVRQcXZtYsKDX5L6htctL550f5F57MJ0OK5HkHShRtzZ28W0MmOGnqGQNfIy0MjEcmQPCAziDfG
7UZXPd7lAF7r2jodhIHEvXySMCmCS6TSoJ5CPRkhd3HMv13n4Ila6LSJ7RgUFcr9qrkTkcPeu9Ax
aRHeePsvwQ7BGGuJOq+pnTxHFyAfh/9f8rafXabm5mb43OZajlVjbMOgefGiJcgchSMFyOUtv7nV
77pfhEBfF/PsGcOvNgY+w1b1+AUJQ4gDJX5vXQYWHfTYQwrZofcZrKFeFZ0fh2Wx9ouMka3IX1Wm
ThnNjZWlzgIVVBbFlnH/8B2lOrWUzdbAhmwJtfiGCB8Zhd6j8P/F20+o527TNuIK3dwdtVWZofwy
egBEdsZB4r+Ug5s+gF4vw9OGv4KLm9zOrLDDmiOc/Gh6b0neYK2fxU/Yyk3AQoZ6cwndnPqZ2odP
r7VNowqskKZlcigCuVyNWLXE9ELvttwaxMlbtoDJDeYxlr1Smu7k+WAau0UCts1makMaaxj6Fyrh
NWmljdD6R+W4I2CkxhozzBWBx8m9wJnPk61/Ea8qnhfTrMgNKtppI9XQizXZd0mD0OPQIeXDhkjY
HhGXFSG+gIQovPdMgvyarRI/RAlPN5oDNer5qDmR0sqzJRndSwuIs+j/Kbx4IVRxThP7rz5e8Csl
UsHHAtaFvketHb+PqE83HKHe9PNVdNNc6+apWqYZF8GEKVoC3cpz3xNNcgjKIciuuiXT58FrTt0x
gD1YFJFvaU1WPQvW4hro8xsE7tvYqKMeC7nV8BxiE/bfaledJxbEQ3+ApfSPg+0e4n1/ppfgy8hj
wRkrGxjzi5VQzkG6Z3tkgA1oi/JZJZlQa+U6gBvpzdTkwbUenVSRYNlsnp8JK9SJSCVUaDalxu4b
ichk8Cs2JQB4BpkNQUmP8jhHXi5lOBBnQipC9hGTDzRsfn8qeKOMzO/o1w4BlfoKUWV/zv+ZGj0O
Z+CQL01vT7+zrg6i8+sTwsr5C3kEZbf7qFfgga7BRt9P0fCvDhbQaOFVzJ2KkzeCyxTytZE3q2kl
6NTaf3wFlq99gJNxA22KjHwdfirDr8q/H7OSbIgtBX47g1FQvnZPoU1BU5oPwL88ut5D6IVKXvar
IucMGy0jj8gz/3L8jLPb0OJ4XsN3U8t5qzCdJVSi6JQSU8sm0hZqKyapoJOiFAHiM7Zr8R7yOvZP
Cz8mKMqxvm1q6ffST4BPb/+R3PX/3I92nbEN1bxTHzVEX97MYvPD1qDUEz6NMTtD/49zHliK/e1x
qB3+2T6vP2lseKC9JLhXdqG1Ku0pMzIDwvdfDAz8kHZlBq60z5nh2o/NJedehzqbVw5+me87qyee
UcbP1YRqX2zelradLbUrUh3Wo38C53IxnRri2UNvQhuVZUTTRvoyQTwRJc4q18jwAawr0QzoTogw
wNRpCeRGuS/xJgUCEgQecIqV+wMsSPzWWOjNeViAZj3iHFzttyd/a4EXK1JRRlb30lA216eg1nDd
2n5SltI6s1sZrxelXXCF7NK+F+oetoa3/SZptbsLYfCjFwpYJLPyPysIQr2EjMnGZpn3paPpTsJN
VIg3AJqcAoGHr81+NFz++P66kXOd1839wJtbXrF+PQ8SWqllxKAwH5v716MBo6rz9bkBIxzjw1jA
oww07EWShe8OkUb7Sm3udWPThiR/3a5Zd4xAJpXF7t72VfHkH46R/ejj2pfkPuAuOPN2IOqdIEvm
lrifm/Oi9+943lqJ5ESEE4GPw9ylZbxbuwyuf1uD6iUdeIh02edbQ4hpojoeXgR5VtlAmQjoP99O
gO+L7Yt+JB7jd3t5yWY3y92tA5yU/nt/ewLTke66lh9TPPf1DF/gnlTiTyPV0dztC6UG2tZG4owm
qVh1LjIfqWbi8SMh/2xflppuvtLVUi02rCDO56/9+rtCS7UEDFxI9e4Ka3nXw0IHdGG75vx1Fy1Y
CFaXdXftKvK+4Kn5gd4PKolg2eea1KQ66vsMGLk/9Oa0pdMuiNJnY6Iy3QMCdP+jeJ+Rr1blwIWx
xfz9muFQC9RzGwcFE9T3MRZXMcJq9ryJlhmQuy9Z5DhjfVgobSrwqoySo5BmgvKUMSoBrQCgYmtm
IRSfhwSySz62jMJ6HfUn8wa7s4+HWd1LTkqL8D7i0aoXLWvnvyqMEPK2MvDFIRO6hlW01ecgDm2x
YUoxaxNqbbBvjc2ht2Lf3snP1UamMFhfOJLEVs/Cv8k0VLCIUcwgy2Ij+j/XKEu3tabcv1QMOuWG
UXra8UfgVLALP1h4alKFT47HTHyzqiz7/iOT9YEeQHJkishi0upUrLGAx7a1VZ7vDXBX3wYeJhny
tP3snLJ9sk9z9ZZhG7EXz/TXTkqvj7EWagm5h7pxeY3iZYa/clozw5gzwGJouJ52IleNcziT9aaN
qCMNA+lDaRpK2IRABmf22Jcvx5mOB90OderaUMS0TzJ4Yjj/doz+OQu7kGF9+nr+WbvP9o9/tymP
We3mQ6+p1f9zrH+4t6Wk1UtgcYx+0vg+82rCXPWrkjTGyN2QXwAcoDetfrjoZVrIyipqH3JaVncm
bKvOcQROiVafzCfh4Q+qJM6nEq64JB4XP9eyiV1KrhEslBuK1ZRyR0yKqqfILjKwZ6wEF7GzIm8+
ln1AJQSmCMm+xSa4/iq2CSlM1PVmU7O99Ou2b/oENCvBnY7oMpje7nkLpy84st4LqeShQVJFU4dz
ZypTg4+wop2kFNFHZdxKXl9kjOnaZsl1kXjTtPR432j8K6FZNSFsEc5fGtRMZJNz2ojA0g1vMhXh
bNnFo0Ac6GOEmt2Lwy6v6xzSVi6UZk9E6m1N3Sn+ZhSqTGE7+7SeSkHD3B6lpVArrEnBPN7IkP40
eWUuqkaGkQhx8vQc1o/jBTv3tnm1x3cy2+V59DKmBrhnNT3gu38hnhCU4Y8HJhUqT5D4CFn4vwv2
GmkGwQBeanLL3dqXEUKpnmp8bp5oXa0+aK3Tb1GP3Ckt34Y/2wviSsxlezd2i02jWnARuzvJrF2P
7p8a246IRR8yF++ne/oOMUpx5EXqe/h5BOnltJ6o7ejFdnWSYFP+yencwrX/6j/Rf6ESzpDS7QHT
L/anyOTMLOKC8b0ilKmbKAD+zbpuvqMe1g03abP2xR6gDKruKouu+SGvcutm0pHCo5IDFNchIxlR
L5SJAJOeqYp5zhbZvV1euNLakXqYuQRd14WM8PdO5T/+6tUxgF2GC6rLVumD3GQr3EjkEcLAJwC/
4U25kqC0k4JQ3T35DpTTPGky0BVQCsWBcSItK1jU7cSL5t3qbiCGty8KuE49ScdrYseIOfAtQlFz
eauV/YqIB9hu008BhE7NCF28MtnKDmv33Di0/a8Iw6k5hkHDa2nyBoJnLPrZpFKcU+PcGSwSIO0d
XfMxlC1YSwCT4/O5oDnlFgLh8+y57a/qz4ub8coz8hvXHECFnGGD+U7HBF+b5GDUujtbxRNssVEb
RINxJuwtCFYIuvEb1gn9rYYmJPInXbWrBe7ouUSu1XPmh9zwBSw4dA9kFnY2de7edqhEk8SKn0TM
ZJIclxfta3jdLfMhJO8DFYThagExCbk47ZE86wZgBMeYuUMuOtKFWuPVpxJOid3wFnz6vYlXsv+Y
ltc7g4LBI5IQu4DxH2EzmWM1EF70CrdrXwpsIr8gCNbgxkH9YbpOOCWpwNJj3+dmFQmi4e9ue0rC
j2y7/KfFeGYsmZiGJ3sKod5Ui43/fYwTz5VR3HOoqmMmf0Ea6QSf2DxkdqreEyXxr8H9poGDrQ5A
jhRyqYobqkotmk8BkHlc2X6LX7f4G0fVwf56qTMzE/TAACZJ+JnNxVG38GBj7YK7eu8GbYD01uW6
0N3QWCnn13uYva8liLTWYUZF4rctKTqYNf+LHr9T2J/Ew0IuEspqwifYcy+2fsDvXx9yC18+Mm3d
404q1l4c1F/Tdxp6saWI8wDw08P9VZcs93tKhFuExxM0cGlkV3QLQRrXLQ2ZXrsZgTU1QJawNYLd
nQbMl4I3GlrqFRfwJviBxyUUfr1fTWmW7UD5pqUyMm3FkucUuAbCyVqaGsOuXJNrjW1kjyBpop0p
w5Kst4hpSEnG+5ktMHD/XvjluI0jAQFJ6FDZbzo+HXlBWEMZBa72l+rKjYXzE4+HGZYhdAGSWmxy
8anDefMeqyqRTc32P5QeEIBQHg8zZIyyzN8OxEZOA0eFFc49SNWKjwPZeaZdnXiZKRxzb/IT/h7Z
55FtFtQyrCMltbY8NM+dkjb+Q4dMaGMRPMkL6Meo3dpL9RKZZlXn48nipGj+P8M1LWxa0CF6FVXz
atPXTpVxS1aqXCcBmkyolIxHzfcBzyKtidUDFc8wLnR7fdo81wseOrtKR/9KoA28Rik2anvYeGEE
PV2vwNlboB7RfHsMDhAvaAdE8u3kdB73kvZ7GwA/6WxO6Tg7oWtV4kzreDwUc2kafachXULekFzo
zoCUolxln3istK5pApSwXKi52yYp5vKaZTSa0992VFvp8v5apD58UOCGyooMy6aEPbwCuWxJdARe
+cOQrcVfp9Tf7hq8B37rggX83EOjLLkc+cuSjcGyBJRuPGL9TupX7pv4xBzYy6UaJd9Ia8PZRblp
INW72b6oFBSgKFKototRH1R8SDh6WCQVihif3DizK9MmhxYm9rp/HhJFuUZQQt824Xik9Qu/CV+d
ixOHq89ahphPBDjMqn57QysDPSskPU34sfg2L7evjdyG79bpIDGzG2zucK+WecBQTg1lnNtuu2AI
v/akwXVwuZYCnnRedtnYQQXs2fiMn4cfwJHM9rC1g4vQ8gMgt/Xsl69nKKW0NUnMMFm1behvVia+
AcrgrfwX7t8k3vOojyPxLHZLNMwTsYoJsRxmeNfltq6ks1SLuFrQBCklyLCgymuxt5zehX8m+JnA
dZZon9Aekf2p+0F+H0GkYPqNCKxpXE1ah/BU/NWBDhTMnsU9HaOK9czB/OP3khOiPKxwEUsC9z0w
dhciii4C2h3U/L0TGPQf38qapBTkmB0vs98BI4xwENE99MAd3WQUKF+oi65hpia7eO4hwpyGSjL2
FHpgr4p7wN5uXzxQwUyXgFanc+5bl/jYHSNZW8H7hET1mgYyt+9FGIvcdIu5C+G01noyMmh5Kie9
x4WKMvr73QV+M53Zco7sDey/nPR+tRIeeiLiC/e036WakwJETjIiReT/gZKPIRgaywpAueKHBBBI
35jCQDIv38a7PlRIfdyjA/2mszayqw4BAm2M++dsOlhF7gfIDIHTlfQtudDDbFFxbjn7m+2hC7rh
y6LPYxZKNx9Bk6gsV8M2EY5WPl7JqxIrf0M6z1JWbpNMvOZQmWrXIRhs1Jd36Gtx8svQvdDeTEEv
GYnOzkz6bhUdvxPsunQJgLoUw6IyQbVNlpJazMS1dZ/xtx9pOh9pp3N6SZKnSss2DNPslnacb0e+
go86XeGich/AHDHxBGVtHH6BxH1UNnx6lVGrWA2QccsHVzqS80mSt+eUzri+pGClQMBcb4XqmTlb
82lFOUqyaXs7iyS3tKEi1AGcxTJ2Z+9T2VH+vjHBCUdDzc6cun1VpkNqpuF4xX7yU8TQUz9h41wW
0sJeM2gZVtFNoC0NoaY1lygXJ8O4ObKrXwL3ICXVhrp6y5a0mSgWDZr8G/B/5I0Q3rdNNryvDlqo
WZu/lIKqjpR+S5TJfhArIerArWB+6K3/kM35FbJpLD/s73rtpfLQEkzlFCZivAFQH/zedTo0MJ0r
56+gRmwx+1Ot7U/2dyE0OSKQu4IztwW6NGl9/ln7RouraFa5AyILVZodMH3qZTQA+bSWLSLBEsdU
UVdy2W1guL3uSgBexZHIHc90eKLT+Bh7L27AZ0peDF+drlZPf1CkdgTAY7fpxIv2e6genwV132db
Q1KT6k4gyIMUebVwbArympl9VCLgZ9CeMvWAwT5qnwt/TjAsXGC9V8tnZPQWd85jRTbfRT1P00pi
5pnrWyPKcXCLtDF1NG2ZGt0W8ZvpglbjFJFxbNPZ3SAygGyus4zJk8RrwQl5xw759xv2OMPggAWv
suRrdlNTwor/lEG97ui6VuQd8bgperGY0w8ch90E5+dpkY4JzoqVz02lrrm0ff1lylL3/71BNr64
wWbW2S84w91Uf7hZcjZr00/tYnKsM60908fFpf/WEToAHEgzGGUpp+fnzBcLNet9cw7RHsPmKl3A
AXuhjTMWOh68IYgXUO/tkrWDDTzXJ1mAJPchqZC4V0iRXS5rV0YAd/EEcdi0x7wvLVai0SF5BXaS
iH76ZGosCa99Jao7WU20v/dtOFUO1McnWkJO110eY1+OF45IhmMVoMizfdOpN65dbgj94SSs8TE6
G/8ZDK2L0oSIz7EnoyGRSZLhIydMKUa6bdraERTEEubQ8e6P/lNlzkiM1XwMFQytuLW/e6FDplxa
cI7zOoJ0cXXhwDJOmyLPBvHtk0NKV4RpSKT6JZEFol0tzJA4ls91IQV0TPrlnUa/8I6zuMHJzHbc
LECCBnA5oC2AMZVcVbo6BLjvHImjno9N+Cvj9bVDwJg52AcYR4OMAPV1EJBi69LnfV1QBG5Za0YY
EHghaGmpNoYFmOZY4zXefIW7VQoj9pSqmylxQVDSXM0JTfOGoniGmn02QuQBY5hV4mbbey/4bCTQ
+BLeTtTzxladNsvCERYWKc5TBwZggvpmFG4WffqckxkOusitVH6AKnBGnEFAnG7U66SbseLyAsRp
+RvmHnClNB4vzpWa1iHP/1O0vsnntowOklsE0PaRskA037+an79k0ySJAtc1k3TRZX8KOVoPF7k3
6WWa+LCX8xCk7+9GwGCiMwB0Z0JNT/SaVa6Pb4YRJdSkBaGl6Q1Btcs+4nRqSoR0o2Mb2mCKMuzg
f4l25pbmCVWpVnG9eFaPBfCzrnrApPuuZCb4esBETlnVDWCyXP0V6IY8alINCLCEVJqHsD8ymgvw
rpUyEyAjRF57YwoBiYcMF+JDiTwDZH4KZhMPvlHRqGUnmAxiSw78u9Z/Ry2sTZidUSKQOvr2lo6C
7vcCXEoAFBRV4vtIOCzsGYxHpBlb5yMk+ZOyGfTcfZ0fiOYYjBP9u0aUNl6hVsieQhW+7uzqIjJd
WRZE8furjhoTUTShgeSi0OD6WjKbDUn4SGYuiUCYPK0bBZdYJ6pjP/qbTpAPELhHBz44HkwA/8od
OwK7UMszJ+DLeLsLdgpGXlQgMIvqfO+L1hTMyS24Oi2DhiaqKBb5KIgDCRJojoZjYxn2b+j7rVAi
6MoWovLoH1a5sUkxcFG3whbs/YUAHUFjVJyad6J+7LncAXTF98L82iIKvo/XEbvSMKE9eFoEH88w
4RXpq2eJEI7CZg0GBIrdESEanROP4ThMfzn34sj0WvUCfieKKpr7ICzju1wXA5pIokapEDwz4ZzC
8W7Ao11jvGYJy0KeE8Uabx+3yOZKdUwyIZHkH1lTV9PTu5SvwzdrvKwY4bGSmzjfT6WtL1i/tlZP
Xnix6ebyQxbuUcXrt/n6HqExO6KzLf2Qk5Qdbo+SGNsNeZUe2hvV+STuJivgeubpAiMM7ORAr/K2
ELT89AlIjoSDXh2IedCdGT7nsAcQUcTbRlfhBiJO2JL0MR2XmIvwE4TUvDLncirXwfdqnYJ8qKgH
FDya4BchQSrPtBgQpPYtX4Y8Sp4JeXwQA2qd+eY4WOxGzZZnENafU6gDlu08W+uzmMKMgGgEV1es
OJyK6SRW2O2GWau2yUzbuChxIEDTfw8MLisE4XphzfM6CiDJGhkzMRtmNo+/gAZ8fBYpiH7uIz9y
OxxwF0rsRw+O2C7cHpAddd96cm7KFY1pDHjsXrvXOlZ5c41kRjHJJLnDHpOermUBy0XG84wY7VI/
WTAsKO1bwXNpIwp5WULLlTv1E1IR113CQ4VMaTDNbvl0LI1cycxtd4V60Mnzgc5wWyv/rhFttRVF
kKqNrrSd2ZB+AN6yMMu9TEfgDTzPJRdA1SrBOwA8dJTF6Q5Sx+ojxRKlGw6LxMw3WrWDPyQbAgcw
WFuroU8QzSU7ofqkO/0SYq2FR+JoWKTzRynBfZU6r+Gu+PPOMVqZYYRef2GlZL29kUM4mepgAumW
+wznOMBS9ErdrHDv+zauxcpOXqApXpiSYXZZCHU9UkN4KUBBAIdD2/WQq5JEcYE9itz6S+ueop+g
I4YjOmR9pJwLpg+Mvpel8BHNZ67D3ZwVi0Lr+HJTtasZOl6+lWnBPI3brQVZC+dqOl2o5zJKrfFm
s4+Cz2VieATP97m9UTgHaRO9fuWR6t33L0RbnA8VOuA7CxFFdO4Nh4Wqstw+qC9S0OULSSPuoXFd
Hc0TvR0AU6eCbJSWJAJBwWZBB2p8GUFzw7T6/aRcT87fGSzzCMgnFt0I05RVXByYm5gqVbQ4bzyR
C89XfOyi9TywWOSjeO16w1SXRJ8ZwC5wAd2yRe28pa2YXpwJZ2505Xaa+RLbN5ykRtR5a77KLCyr
Mlf27vCJCPCIHvtd8Sjm3Vy5EOcvHbPJMJk1+niblbn8B4iYHD5XLdPMJ/Lo3N5OFA4SZcXQjowX
v8pfnDlzYhCkNHF3OR8VEoYfyv5alf6rb0h5neFsdSS0qabs0wSTXUsOggcFOZ0un1COxoCgwuFl
trclia7CFRwwiYuZynpNNGtHrVfTOZIq4fklbQrn2UZdMtBnixwYcjmDIrfpBXpwZ54Sccjr25zU
EA1U9BVsz6x0MYFjoS7YLQgkeKDEen0KnuzHFvT77wqKjtx1F+tPhaMB5w3gXUyLRqHchqRSOnur
DkFPwrEPTuUWUdEol7l+cJoisVOxXXcafsG8LvPXFEfSgTN82WTgeuKtOpHyWPMY2yltBeF1K7TW
xUsZIsgxlP05qWdHNIEhoHl1JbZtYi4dHducjyfio6WsMZQ+TDdYGDnlb6k6EYTXY7XXvMwPYkuI
zEvgC+JghYg71BPsxuY1sAV5dZtFSVXhwrZKe5alK9v2urkKqVygggpV3KzF+eOgj9qUruC1tjR4
PjaZ8Ni0bbu4E9B+rJ10Ao22TYhg3iVLCqCCrcgNqD2uf1FF7oolSJC5uTOTIxm4PNi/F0n/M1Dp
S/dZdR46kp0i0Pk6L4oRFcsAiRM9k2x+2ED6umNhgLGOovUoMdWLvI+e7cSl9ZPYTNabLw1HSVM+
aBWp5+B9tpHEoU4Wr0li0OIsCezsYgmW+FyWCRB2NtZ/L/vF6hTjUSwyKD5nx6qu4484B7TqxhP8
glgd/2q1zKwbboZnMCFUxCJBeAyvJ0n0MU0NHnNXFe3SKo3Eth1mFAeBMOUCizxdw6qiH2MAT2Ko
yIz9ekTOzugQtJr4jbUGR+k1jvH9WUHPesR4RdjW+cIQHbis7trGtxtTyUu7RLjaTRYmJOZMiK8c
6tk1tNK15MiDFroQF+JeS7WX/BkXbzTdChvnTs4PNkPqijowdRo130KqU/wWekfrRiDFoREDEEoX
ZWxt8srti/34OE09k2b5K7TEzkqGB7ELcBsTxgUt8ahHo7h9ABfCe2c5oGPRjeiiBdmhl7Gv4Eba
IP4AaQGXTSQmZ/KJCrLZj5G2xvHPi7etcZwxnvLxrNc7PtUZxgE1kRwy2KIbQPK3c0/hvmBOeqSJ
bZmaqoSqufM2cPfFhOqs2RXh/AfPMTDmkO0ttt3Na4VLeySDT3xJ5s0ZoFhHlTa38Q2Py0cGrnJs
1vZ16kt5kiuKDsR0rBa1BW2Gi0I8jlEuHFnT01m5mVCKyLBTrjOFhduC+i0hWksuSqL9AaMKbxTz
83pwqpHWCsVOdoTtuFjB60WTvcBhrbSVWQVwmbs/5ph5pV8ssc1p28qGWqsieqFyoSdjXpVC9kbc
vOlA6EMP2859velntW9DNDWQCnrr2c1tDJgg9nsW3XmBp7d4bb4KzWDHM5VM3tCp2nMtQo9kkYiy
4gROFiT701tPmop9wk4DLUPkcoFjR/bHSEs5dWzvz7aKFAnekAhHQPcjUTYVrzWRne+HuPVxZir6
R9WCsiIB7lNoGj/R4v+X7vZ8ZhrQojB3mO+dra8phnOiWWY9K78vBO/z8/YOexiiFFpJzi41/oh3
szp0SXEMS1xxZ7YzW6ODxW95r9ULY3EAUFc8M1j7CgGSOiiewsIJYwffwiRQ3IZgNA+CaZ+sSf2p
f6z1KgniMQev3aDIuQQ0BLGYzB2aLpS/C4Cp/4FSx3fU8CxISNyiFqgohkJHlaG4jfgTvxhpM2op
CoqQ/iT5LMuCLF2gy1DpkMj19Oa8cIqtcrwGsEV2MiqA4PBbO4TQT7MUSgqN7Fben4dejznbub1G
CIA1YT54Esi54hNf3aj5nEwUm+t6Syd/FBNQ7Fozgs86ToeHrysNOkWORnTgrFOQ1BtdItjR6hSW
PV5XFzxE8ynDl8Aub2CuHnOVsxQbLDjXK3a14cEG4CQvu5IazB3eEnwtW5hIvUfMCHuaB3gBDsPw
V8lHZG3ZKIwmFIB24U/vlO7+vIS4J5nlkZ3qz3YgIPC1iwDJuL5WTQ0k4JZRXnSwuztrbKjIKK7Q
uututZ0raOMdUDdZ71osyXfZr4zj8/YkyRUZ0/s4h02t33dZIFWiDHy1uwHYI/0yNsL63ikn+gS/
wp2HO0HZEhRV28BeK8J0qA7FWxazq5FFAcoxBzKNW2OMO+7+kT5ugqK7GRwrG4Pzt5cFOLcyUcMZ
D185bEXHaBs/MDKKPZRQjmC2VH5hVHoT09CLfy6Vu5FaN1E/C7NuGaTYA7ccC37wUdfXLCri7QPx
Tt/upuXyU4207VA6EWxdAJYTjBeAQ9sB9uMSQWDfeHkTXVgRmE9F/X8+fuqxsyIip8EhmLxYxmlR
Jf7Aqwfk5gZ1P/M2RevQqBm5dfKk/qLQ1bJasPr9NhXUcC+iZlhJ/hfzqAXq7X+Iu4eLmY4Eqs5m
sG0seN/s5UbOAq2fEki1KAq0l7LTck+N/kYOTq7eauHc9N6Edbr3ndkggf0Hdf5gTprdPmSm2PNe
dyNjwq8IPq9dZRu1ne08mbuVtsnUoQygupN/CHYvTT40n6UpxQTgraJYLk6vQ0hgp3Ffu2/jRGi4
eFvBHy+A6hRQfGwdBhJjZaVknwEU+9o5RfCDUqJ9R/CMJ6nqIxQ0LX17O7krY1uOOJT1qyXPNHT1
KdCDAiWWEY89SpWXvB8K1lmUf2W0sHHCgNIyyigIcjrplysnB1IpcikEFxidhGG7FfgMgskS+pny
AnPnNK66SIvYUGgfFVf/5qBn9vsRRypFIf+OU38K55INiySmM0KWZaNgm8rpzfWpxhiSIrgRFjN0
UM1ZwbLGAFOXqskcg6nvLnsMrpeZqLpdlfLYR1D1NClFSIE2GYjtROwbxHL9lMtscXT79Gee3/yX
R+04efLgAt/P8brEJs+GeEL+WsA3xK21RQqXRtSQ7zr0s5UdI95WlhBkRNvyFWxA4Uv0a/mrQszp
MEQnbvEMxAaaGEzWCKJh87dNYF2iq/2I1QoqqyQI+WiKT7r9sJCeFU2CmP1XhfGv5vqj8+7P4wMB
FdCJqynDGVQPyFnhAX0r6G2YohPzq7gQf7WMqnAW5XbSJQMt0h1DVunMcOjfoAhrHpKRnU2e5nLu
Iai2Ff+WN0kH7p+jQtB88fVQm5CLO6m0/cQcEpZdpJaqy17kxki0zy0MnkOBzSEsR+ayDWtEU+0R
9LfmQT8IWCpaS3hRXemgHQvVcbk8FFvEmkeZ8Ixz/mLocTVLUlw/EZVahi5n9NBSUXNzxJav7Z+e
9jbgkR9i3UKowNRTKgb+0EaiHO068+MFboESGK2XL5dfk1OYigXs5QVXMfQzjFWpldCvAxL55O4Y
3NMs+8QK/UDP+TaA8tVUhzYUIAD1HvaoJuPXOa1NpBLyVkwV4ZfvcjJHwzkFTz5D00u5PKAJZl3V
2N31uBje/cqB5eaijnML+epzWNBxgDMCpWPfGst3TaHkVFmpZybDkZtxNmy4dgEAiCe7BZdF2Tsi
DS+c7in1cCyUtnct3BrcgeuSarzosfBsRPV0dwsdjXkndywLPVZLeeDadTcuRMMXhMjXxMMEGItT
HjgTnhAtnVzrA1p24XfLCb8xGhLtpps8fOBRIvOIMjBz8WNEcQhD3/+dmQ+7QYvYesWnbMZgSWlJ
/86RgFTB5iJXbDCF/BNwVmPiiMCTkp3R055YLZLwchuzCogKWVlXXoo+UxDyY1ZcdElD/xkd8zMc
MnLsD1XsiKGhnyaygYU2VkQ/p1txjvLkArIF7QRZ7j2Wsdqy1VlLc351yUwiFasX/H8WffPK6t51
CQSXG6DZPyAZZXUExtSxy45UmxKQVMsQLst0G8hToPGfDd10tN1wpmWoGTZ8maE40rQ/isNC8vp4
t7exhvBm/tBqXmP7ukiZvQS43DSYZAmo/IwzTRtzf7jRQ1APIPM/JZeX8n+5U90i8R26QgXR9uom
me30XNivzsw14m0jfwlen8gwDGDviuRJLf4rHNIf0RUM+xst6xL4fSK3gdz0RsfDTnsZEj/CBiGR
1oot8jbbCAfMDK9VZgfMuIqotS5GCpOcvzjsk8kkKhMSqQQYeDXSq/xrQ1V3QZIi2TYNy4Y07UZ/
hiBRkiq7WgigvBI+D8EEGXHfiK29Ccjw/kM2mFXwtf0E6BngCJKQ1rJddB6DGF5xhGmeChqrCqTP
xS4yq92wbI8uLWC5pZNXOe38N4f1XiFxY28qosC4HKe45pZn4IgepzUwb5OVz++fPkEQSfMjei09
SP8Fg25SWmoPa6R/cbtR/dM7X4hSfGuEL/0JlpTI/UmGMgftWHy33Yu6DxMa3sl2Quk2CDXldDH3
Q3cUhPoyGehZ3zeFqMAYh7jlrkxbY+6fMFSgQ0Td7nMB88DFd07bnqQoB4rO6eB5GhWxdI66gZ6w
rrASFDGcU2gL57wlxTCVbhQFHR8ivOL34b7E5znALdl9Z2tFds+UwTLEcRlJK2Ia0LaXBCDvzBGU
8TdaLe9feZndYyf9HHs9fUOQc3xBXTeV6iBa1cTRsZwFoyW0p02nUBVVk8c9q3VJiEN7QlFTU5kJ
CM527r8oIRKAsGD5mWRcDJL2Bd1AWM5vJfs7eLBAiXHauM9iUmZ+EWR3xYBSOzTj5swqk3PxnNPr
Xp7veAGiKTXUJ3UaGLtrYDnhlk5tKDIDvVwc2dtGMO3s6V9AUkxpF1heIwkI0j6jYzyhKekXqlcl
KMsxS+B+wakMIJZs7ARit0tNfGt0C+8Qo6wh0OUbC/2RIsV4ql2SnAGXcXqwnTIBI+HnwOLvsZ5I
S7aaohSDjIAcLsv72G/qOeni0cRUSmNw7DiiDwqVoRxp76J+m5VHa6kbbHOWcnHZ4JdbJJEc7rmT
KDV7cHQghaYnUd8EmGy8SHdd/ns6/jDsx+DMURKIkjH3Rnjki5aK0Df+UuKbUtuPZDOsFwTePhKe
WdoIbTL6I7k+hh67SYHihXV/6X/Lg+QAO0sKsidzRfvCjh2m1uleCiZ/4uB3FW0jzGOasv9D6AtA
Pz8aRKDK4dcRjBIRGzFArhThQJmi9p0s6nUUV4uLOgUzF0f8ruAlgieOMaPM8OczHZswQRSpwtoO
TbZ8/w8lIiXeBhwaX1fIkifBsloseOMhH6wLjhIRlXo/Fem3F49QP6IHpCsxKLfDmxduLsp3pgnr
Xcjxm878SZ/eLoq0rpeHHy1nVosRXtqcH0FmxucxcJBvPlA5A43klWFXZDeIEvuwNWNhJeGhbuhN
3Dscb6VF2DbmvRvbmayAsrDDR2jATGUSTttSsJgWEpLYPi0kEuyRVBSKoCNPE8XLNu1Q56zyBt6h
0CoIbqzJ0RImwRXacVtJpYuZAfvyx8ERJd+ELpVlAAuSfxSOE376qav8im3A/xNRZ+MmDT1mcEaG
pFiQdEttuoDkwwUt2MvrljnaiYpqlVDkN9Svk/jVHE3pqy+sEQ25F60iSxKXZEv2dwW8kMLOtekS
xoMPk/X1zH1AnGwh4fnA2GV76AygEpVasodz/43oACeantedxP6jWQbUwl7KmQzL6GarUbcFKm8K
mWazCPj94eD1toi7uImvq+tccTmag9eZ5gvlgiqNBkAeYbpmUub8rMleaEZMC+Z+GmG1RSH1rIt7
j7DIllEnzQbNGUEcKpR9W8n6/b+UpTtekgq5CX/krR4AfjUgSzuW1K0ogy9SfL5QOpyn4c/LwRmF
EoW4cwJiYpKOAoPH/B7BTA+UVtG9ViCmMTTY4kgXLZ8b/b38VaF5PNI0s2SaGof1Jb5bQXDh+mkE
Y+G11v8T7IpY2jRqEWLSmfvrJ2ZK95Ag0bFnbVhH3+/+m8WWaL2Qo4ss9aPzYlyWBjxYaJahXoQz
AMvE664P9f+tKX/E1moeQCMOEe7LFKvph2yO17BRNJlDildnYqW4W3OxxCXgpxVDMqm+LU/5t1sb
eATqq8TlnCMqdXYnmjk7t4jALZd2UOuHFECa2vPbLkLOoE9RDMuCit1bVcdP/GeLXQp5TeF8YaCZ
2Z745ezpWc6DRb4x09+8M5/bikVyKGuq8w49Uzl1Kmk1Go8/GsIeICMEttRe74BCGblWJ/09GYeG
ktzxz3ZVdctTGAT8ROP/wg4qPUNpC9ub3xoe7l8dPcFeYeHQo3Wq33rRdvchtLgN508QAn7hv82t
BmUJxIVPAkKzJlbIA3UfHUXt5UwvYIdaiLS8uSBipaDkS8+a5KtxANyf49LdiOYmHYQh/GDGqgoJ
LeSJ9lVYt7OXlDc0OLH9r/P2GIb27F7WETRyLzjCsFGvzMWQjoPg6N4XYWElr16kdxp1o3gDgvmE
obzAHfhwwNb1ZQgo1unFQtaHdVE6k5/0MMzxRM3wjG9JWO1mvN1yTylxQPk8GgC3307cWHBBtNW6
uuYZGJ1dfQn2R4jvrv/9AqVmFAyX6NI2LERSmPzI4wCrWQiI447RBA9ZT2wcGiqDdmDcpfhQGyrE
qYKXhX/lnyvS46VzVlYTNeNoLLB45C+saHP+CUT5GGJ82skkGXEFw8IdFxYNGfIYQSpF+ZTWGHrJ
dNmUY2eUt3YDnrqCbbba7fF7GknUUEeXpyWAsJYin8tvYICAsNtJ2aIrI76Ig2C2JX0/3fq0FvnW
kt4yvTcpcPVDC+iz7miWakSNJ6IsQ26HpYStOaBS2BVUWkma2eqzzA8vMUubSnyw3HrMWh6LPqV5
gN+2VQKYPFD4bccVnbhAdRhVzOgLiWaZFSXzEcJP1XWpQFHUPmzljOMBBTURxfE2KemNvUBZdAR2
EXa35OFI7cXpLFgfp2J92+80Jg35Hshe1/l0SjwHBUdxRiF6x+HCfkOVqlgPazvv7WDg/KP+qZu8
1lxlQQrwb8WVKC34SIpQkqpJRiacd4yaFfnK3a8tmMPKPYi7A0uTzPoVs9SEFhogD1dEctWLV0wA
JKksxoSeJaMTjdVJ3f45MBS0ltx2O9lgv+T331hCYz+4NCesfnJ96SrS5x+mz5+kFWb3NnnZm9Sx
d3ayJxZl74A/SxGVm/laHaMuLDdX+rqTppmfrMpJfvEfFWoTYnfVcq15TBWxCZrXGhoPjskBBbQ7
k7BH93f43cGlvXZ7aa0j4dYRG8CVhR5IkpnlztdXFfc89Do3J5ZUWDB+Lihn8FlWRWWfVGMThugi
NxNO8bgSjfHKMGqP12wgBG95iTgEHb0kgP0gtOCYwjTHRfoN+xok9gCX+m6Rq7bq+1XqAD3K0yS5
6NQsWoR8zle9ZrJPngETfzdfs9iybytfv18M5cPt++dbggVz1IGaAYdxn6yYIhjcebIKwaRsvu8+
PevruxBlUwW66k21QdEHI/QQ+d9q2g/uz79yclqtGtrjDjFNbn3srhXjxYoCXzOKiuYqQHR6jYq3
RjeDKKw33e7DwUkRBgApn+4R+NookBlI1NIt+xA4EOUKoxUwzK4BqNAsxY9YiLTuFA5TV/fpbjUu
rVxT7tRLrMlKpMvsXeI+YMwPcfnHuGOLlFcIYaqLeRD20W/6qrbZAaukOejYKsXk3JOFaEYkwsK/
XBhsyFej0kmg/+nKbcFFPKbkFP/d3EdB0aO5G7D9LGTeJdaCf1Jlz6BPZDka9dH1FltFmBta0Wo4
tBIKQrA82AjPjcBTHKX8C6Tc4vlnYTQBJgvfdWfW0pY5WPH+Tb03QcSlVS66fq35FRSmhHJ5h33W
BMHonmUDertGr05iTvifjvo2nrVCnMsfZr4dcRar2zV6VxK0QWYJ3jzkjx/AhVSy5KT1NGgcQP9P
8h4CecgKiLZtP1NGcYNk3CYPiuplZ3Qv5yXGFNYziwqOreCpCGyVqlWL0ThPaPWFmhhC5USAgjyV
NVGa3BHEx+dNIXeYFHQs6Kvx4p+LFn7Fk+l/NIK+GfvxpuojizyMaXtjJpXrXrbk/L2uW9z6ywdd
mF6MxGQpvxSsmEoMyFT2Z9ehVyUNrMcG8fcLBZiGN78Ip+fgWY2AvWFT0hDHAyy9JG7qmSK0QlbS
d67JCmpK50mi+q8i+nuiB+u0lBEHtXIHCpyR35K5fBdlQhSiEGdsCNuDDtMQQpsMjypNoyAQnky9
PGJVkKC52gzTlA5lBZyku07N6Q3v2EpXiJXdd6U1fZCAm6B+HviqmD6M9EKN71/HB3WIwJYWG+c1
I3jvbaGKbE15HRLlz9fTEi64d9Ro1RM/VmOjGjSG37l4V+XGNjzklpJYgB1j1DP6KMon1XkpCmCU
uOKE0k7qi/VnpWtoJEo/VB69rgxh3F1BfQSSNVUb0JEstasDGaQNrkotjQtMuU4Z/d37XBYG36Co
nzSnienfS2dT4HRUjSgKf4ym4oALVM8XVTcORXA5OXe48o6rIjoRl5/rgjZ4KQIF/SzCyyxakNqK
1lGmdir/lUV6KbreoBQ/skxXnULzKpNUi/AOnQ0NvvXMPXuN64K5jxmn7m0QWJ4Uhexomaif+jqI
6F9OZYigfVSUteOSBkZUKQtyVETQ9IK4toaim1V1GT2OtamsZv9On7U9bbV0jJ2bc2CFzFz1IyMK
0mEmufCNGPJIBNvZ0yYqw+76eID/uR3iv0QfyJB4xLfzQxBHCsXQHQ74NAVJtR+tT8j930iYbaK0
Z6m6aQj91IeN/8Ene5UBQosBcdfjfONkFWWcMUXIkyAnZHqJHdVjSUYjs1e1xUpQl6g9wjp2ck5K
qpqsqivym0nPllb8rYQ8lXba3JwT9qrhmEPQbGSb40zc17nfqhlotIz/iOdqpPP/EDGRDTulwsve
DQBTlOIy8XJfeDZyI/qHHObg1TBpjFlenzDb0Xn7m5RZwDNK08dR1kH70DDj3dhUWfE7Es9YCI7n
ZrD3nF7XRW0Mmhnj/S9p3PiPV9u0bvghfYnok6grnzKsJKNtASZrq4f4orHK8FosqjaP5T19BTmG
/LTl59ht5SrVbCByJMBdzWLuMRWireKzuxrBfYMySUo+1f2dpgp0okFAPdJZFI2eFZ3FufHr/oED
c0U846Pw0Jc87zdJ9UZtFXrbd8qbuxn8XvcY5htV+QMblP9yEsiTI82MfySEZTAQDRlZibCOxYVO
IRw5TcLsgt2PAjBv0qfviZ7aulsRkA3VQ6xpifCGVpW2Nih2Od+l4bKk6MZGeEj9+wkxubTpuhdB
Lnx69VM1nMygdJCsmPZDf4GbfACQh4OqV7oyHPUOwwha8eFnVVMQI5BBgELksN67XSadHRhl+OD8
lp4vEjlERE/g2IYHwrQ/B2IQzOrjLisaratmrysUwxZMMY3OVkEACR7mpr6rnmgweTCnMdKNLxBq
CEIW3XXajKHpuIWZb+/iJUlYeKrI/lwmXl3dTTrzsy3xMPS4W0RUDg/aCQm5N72AuxcD1IKExR6G
55QOsxx9Vh1+1hMw6sCkCIiB7BtzMN7zPWoP7YJB7LfZsKQOuMn7sJUrJK8iDn6Xy6G4VafG0sCu
46mC9XX3+uy92ee3JZeUlaZ1yeWpSgwNytV4aQ+8P+NyP9LjxaAhtC4dP/tm3tAPdMcUiX3uUufi
IlWzjsh2NxZNUWod5DRdCJx75mn8FRN4fqpHktT8ENgoyeanyfyCKVR8pevQSz8ywYrYNqRo9zJz
37NwUZEGoOGyL5iLbTKsmiaveZ7yP+v/6ILmwkUyy5UmUC1h84Vpt2jzYlCpR7V8R29HWqkaKmiz
cD5o6v6TINmiXrNWR8SVfUlXNlvNZr/VOU0ctDMmMFbB59FM+Pqg3bqSyFR9E2P8jWdnxQ3sgsax
EAnUIR1Jb09naAYKp3l2cD+wmPI3dF13mntjT4CRNfCDJvBIg/2Zm0+B/0pq/rXzkjSTj1OswkbV
Eltb5MuK2FqN7bVvDlOh7ZGnv7iRfcpfUzIp1Q0V+nkTL+G3QzUQal+XE4AYHIoHTLFJOG3FrYH7
7b1ndi4AWj0befMn/QOetXESP5fRcq7APbgEk8jTPJ4A6MpQOPWJvgrKUqn2Mf/SwQfaTbSVX1db
m8yACZfQn2byTikLeHHLr2qFh4wqxCf1vAvIxVGFrK9VhMeMjnxbZLI8VaBMISRScZrAg1574E86
gFpZVXeLiH63y9r8xiXV4/jIqt6Y8cRuGN1G6LHSp0M6Qf+WWfjIK9iVcgYZxIwaLRprgCFPbQiS
3v2xrCCI1Bl0W8xKSsQF5g8lkcANigPmN05YS4+8K5jg85KDR3rgZN52tQY6WixhXGOqow9OIno3
VSRbTDIvxLC1rco1yjI0LQluAmTZaYtql42OvyThS4c7g+DDfuHAyZIYoTF/Irbd/qHMR99hmmux
YKDqcV4Jx4J+esOPlOsS619BjSu/4WIkK4Ncga4BatL6JV6v9EyfvKXToxqghPzmDjVF1ZN6BNXd
bcWpCDdq049pK189KonHmZ6enkCOGx98rM4jlMwnrsySAJt+7Fbvk/H1zgLSITTQOvlZf7keUVsF
GLhhaDb2M05zwoIsApgBgsJeFgh3k0PN6kLPFRXzVBvDIV91ngGTUGz50rE+uDLEwpil27gKCvS9
I9fRj8NUaTX8Hc0ClEDErmDRRlZAUJxhLcCCZjUM1jrTU/XQ2S7uUXHfK9lzwYWAXnEjWleYyP1r
wUgjlOjtiEtAzWIj+nMGUIk2KNoU3glC8fopc8nUOGJhncndX0v4ZEdWJUNFC8Kf5qCcku/4Toh/
8gMlX0W+8JO3DsfAIcbYfYX8Unt+geioXBM3rB+joPWLGpva344bzUhppqhtyvd4opGo5Ia/pmPY
yylnaLEupvi9buXgQHQp6WmxDZC6ui9vHH6lh5SXnStwWJth4DFjU0eQ0QbDbR5RXrxMMWj3B5u0
p7o9jfHSgYQSB4argwOGzXySc+22NLLSMw3bv0frz7VgTrrEqwZTl9vlAYRVl7wKftQ3HKpuvkFY
ipftRXuwzZN0zNkzsLTNaSt4+9DknChNormmSUImRGeq1lDstekY/Exw6f2usDSYU5wz07mePSyx
KE3xb8iWYzbM/yM5RngokO2Gqsm3lijjx4iRjlOxnHKQTxtF8RpxCp8ErqRSU/kFvR6Vu/iwG5bn
MGoucAbXwP+1s554ISIp5JpAT0rr28lq1sDoJB4Hp46gOFypz04unISdLZ3gdIR8JnBpvmw98jlz
pmE1wsRwI2xAxzZ5fLnJw8rmOOk+8yyImhlmqAHAGUEzJerVHr9C2//4WcHNYwOVGuT+vkXoSk8T
hIQvCOOuu7wDOpHc0dn4hZS6xqSHhR8/HembOYJ8uYa8i+T0gyeEqlgGKlAgr8oMoKgf2anR9Unb
9NUA0JYlTPeR/83RLlbEF3mfYz3wYJq8eChIIeONGzQTQpfYKXFgiogAgXxDkjLjw9P6IHiE1A3L
taMVOjzkKAaJQE1uJqEWakni2tKDWnRDSTPHK6HKNY7WRhPjbPlz2l7aobSfkADlc8VLT+pGtqep
4M9D5qOI0V9VUfnzXb2pkHnP6H8EMMLn47svYUvFrbZTQGzRulgs/iFp9mOS52VrOm2ceHni0HBq
OWo5hW/5mZJCRlHgqSyxJ7Rlk0Q/8jKb/xvKzJm2TjdpMHYdFzI61cT5xGDYZJBjE8QBgGuh/Aqq
Y79VkJWTHVSKg/RqzXvuq3/Pw/qW++ZhqxPVhNGVW6uRMqJI8vUyrCbBtlakK0EWCGmYYL+A8opA
RrgzBdNU6sO0FpSsNC4N9xJIOk4zVoeHifn6YDD7tFvTxGenXACcr0jCaALbTrGq9L6iYYG10z/n
lA9Aop5La5Y3YLft/BYSkKLD/tgppP/WChctk7GFq2ocVad4Ix2Nv1TzA8g+SV+EbMeTxLkTQ4t+
OEdbnqbcKnfs/z5yjxyyOxHW1ciKj8Z3xbL8Vrdk7rwlPI6SG/N5+ubwmlG/3bzv+tXS8euImzDB
UKKhFsqSkVHEuxW6AtHBQ1cn1Cjyqi68DcdbIZDCuhETbTBguLdEnpKdvs+RetA7+fjgGsGqeJpN
5lfDFKDi5o3uYVz+ZMkzGKiEQoOH9EeoeuXLEHwnZpoStzlRzq0yTyPQxCTMbJqleNn0tSRoyDs6
lwueoF/WI6sw/roZxKJ+DsyIXe4CLicFvC7FTrhGk8OjWa0z0i0H5EyFZafi5EaHrkCVeOnPR05l
BBiKJYkifeCbZ0OUNFSwBpBFq6oWxhYx6O3z3WNTTqo5nDdLeB8ZrqZ+y2MOs4JG1NyBkXwd30Bx
y9efXQVIO3l6+e27b6SpsNoTnj4gP554tC7i0FrclHnc0m8zUkoWBFa84XBbKo34LjPCL9ANWK51
NYjNsp0dJmL67MymsbwiBbvBvLroN9Ifc4z8zQpriB87APNYxleLqKoJGkagxZ4S9tQ+uP09C6ME
3UUcbSJW8RYqKuaYYrtsdKykn23Ti9zDtLiAM3Lzeu6hP79Uv8LBVeW/G8ckhplbBU8UhsUbGZLx
hmCcaNEdV+gnMI75PchV6sZrmB10BU0ASs35VvPRWeTPaIznrWwoLLwzK+yLImO1mhUwQD1elZVj
vRyG7SRg1rjyNxwzeCJyUom6SG1OfYldFVwdhDyscHv/qjyQrL00kabOX+C36Q/HEJIJ4mKOqSWX
ivRWbreUx355GNkas+NnjYOrij5v0oPRpJiYZrUBfitTN0Psmakpz4xZu/pvrJ2IVxqTfxfYr0/g
BZqtmcQ9gyWMT2yAWXfTQcEbe4kEM3J52MKFHL/E6GdpXmu33iUOdrt8x9aoLfo6k8kq1xsW1mBm
ixk6MNOpKImLL3xvV1A1STLTBAJek8dCWRZ23Uqd2AaHQxOXuDYxqasSN36D1N6h7/LwAqeuqtfe
xlWtwmOwD5Nnmp+SqycZEUo/fuS43eEe/e/PC48CdLjsMFCq/cuvnROA9SEOciGQOBNnMrXfDCj7
77wIAsmK2JA4/lZ1GaD9JaUVH3FSgsysIP4I/paTVgEh4wc1Qbj5mefr0ZYtr4+x4yhD0v1Iv10Y
Fr/MhDZzknEQyBBFFIEdfy4zE/DG/sVmHX3CGjxI/CqejNhTcJu8SZrUUeb8XorwlRgrHokkzKYE
5fpfFH+KhSBbBGhXbz+REhpTSNClyB/Koy8bvHPLDNDDkeXfcAyrrPWMYKUGohklOPuhPdRpkF+U
izz2xWNqLD+zhuY313W6K/t3zgPQ5ESLdHZ4+vjaforfpbkRC0u9pgCp1uPlr9RcN+BVKrAaEmq+
YBNblAUMX1mJqtSxj+fjh/k2IdIZ41xHqCjBrEti1GguKckZGn8ebq8MWXDpvZ33CkL81f3e/v3B
/kwyCc+NQY8y9C+YjDtg+CS9DbXZmqqo4lFQ6OMtWn/eU1AgwCjOmoxte9DjXojG45E3kx1SyHSS
cjsQo5All11n5R2CSEyHFRa1znmsu2dr9Yh26BBSqS5c13YNESVWf1FsJYhmMUDhUWgYUvcyEujZ
J7F81PwpR76ds2njSAjvazZE2PqTm0D9c0o84Uq/0M10plPpFH6H/4dlMoimR4ShkB/gchwpyvlS
lAk5xN/K6ot/QJ7c2tsp8bhWHqQRo46RSqtphOkwh2Wcea8HrQgdsLrGM1C9SF8SMhWdAxmWV2Md
bWubpYw29QeFU4HyT3XBzD8EryZqfaDHPeoVmWLYlzpJObelkmz+StqFBb20dGEhG9hsUjLjbzyk
ugvACSVj39C9lwesvhZaBz7ZtBEjYamNeutK1M5hk5A1WvOHGfBZ/lHmOvvh7DjgAYuRcnlBBsrb
Najswkbdp57SXJISSRRH7tgqVn2O0rdzAiGosRbickiP6h7Rw9d06qrtkTnGoXaKBT05xzBmSPGD
r7UMrKBOBvb6KP4lKkEOXf6Wtqof5pjz1VTL1f8h8L+h+8YbanJURaExBNjGTSn4qIiHZ/GC55A1
UJLKAp0Qg8qGw60BKTQbWpQz5fIE0zzKOFMa+h0VeTVBkxuaS5Oo9iySW8mEl10NoiuIZaikgG2N
v9/8uZd0rfpKwYw5aNMDtV53UTg15OsRGPQ6n3sZ8wRcrW52oqCAxrLEG8Gv89+nFJdLsAqHDYTm
e7rAeM78G62L9Wn2wLvTUPx3njqV+FSE7Khh5Bx1cRjJqPiDdabiHUfsaRw2b2IYXAGkdP9pEQiy
hd5k6bOpQC+RDvNPLvYNPZrgzMcuQVmJgaaxgZT2xf354+tsmHUtnZ/naT5uukg3GGVNPo4FQTDa
cEgiZPB3QNhe3cquNNmuNjz1ZzPO0sAGtH8LZH8nMUx+GNKYB4zr+9nwKBPFp6QwZxKAvNq5b6Uz
87jJynEWxEfA3LPqErmVH9aouR87UnK+QTHNaYvzfvcTHEi635LFHoAtEHngx1RG1rILjxRHNYY3
5UZ0goKinWiOkX/KluCLElMNpHNkv5x2aYj7QQBbZUJ2HFpV/E4oEVg0b9jGAErJAnW5aksGG9Kt
czpmqBddX3OD8lRmcKQZyuEwkc5ZahwTuwSpIpG2O6sQe/g+6Mm6rTSU6ZGNbtN4ANhhukdedKuj
WVtzH7L3sljIwf9rhNpzLN11i3gpgka8qUConmPF035QFF7lg/qlNVWjiQyUEdAfweWN9rcQAhWN
4Go5pGX6W5D2Xw50yMHmDG1nr4nNJrNhA+l/M2pBTi80nb6BL9xi8fDEGKKJaPclreqVKWl/BFr5
c+4TFlSzZWnRK/YPNo9PGuk8H0zhqZKkcQYomGDRqE78KYqLloqV4b2xzTL8HTqbfAA3iJARi6qH
c0qdt6FCaAMFgpAWacBIP5zOFu9rdMyLjxlBH8Upae3UZSgsBjVdmTSbdiqvK9CWiYUwbRDCH7a2
HZq0NYaUBiBWTu1sIDFR+c6D2j2Xe/F1CHm03ZeKKWJ36lFPHSCl4n7McIOpi5wg/mSuU/rlRzlk
ZqCJK6qYFAsYRCkeghpZsBh2wzofCNMNwMh2gmCIIxSXGeKuQBMhyGvsuBhmlZfWhB/xVNdcmU7b
o1Hcrg5k2gm9n/eyYH7YqjixxgMj9h1gLSPnUB/9RJo6PPHSVlH8kM6gTYqVo98C+/taxxfXYTa8
uBImRGA9vuJ+zI6bOyHHBOSGU9aToiI3MJH0u25oEG/2/a4XtEzFBj7FjygzBnsQPnYr+g45+h5O
EVZo0nyHoFwaHOIFtvmoMRo7cVvf4Dpf8v3zvTADiNPS6HQcXWZY5+70JhSBBuo6pdFaZ9HkrkHq
QiDH1tz9KXYFLi1mOKJHXsLUk1LrCamS41u0RR8NSlAsihSUBAHtBw6jvYE+fpVuIqJqx7i9Ag2a
+0RiCcF91UIsaveJwPty9OE0SsLxjn791WRTn0KWD6b+Gc+8WHiMsP5Yjo4xYU0Gbok5pY8NSCMN
HQ94DAU65yIH6k11H+qmJG5yunfHdAkc3NNOhTfKhqy0zrOUdsHrhxcBesp1B/8Zju8e5/77qaqg
nh1FFMsNI2EqgtjvSslYZqXW2WgZHuxIL2smx7zMWXiukCyqHAWi9ottzdkPGPHG4Vd7INpvLKS1
AcUM9Lm4+8kyiF6NPPuVtGK1ESm5812NmXLb2nNi+CGBxyeJF4WyyUxn7s2Z559qerDGaKUHzA+2
u8Nz7HhUQk4AHg/+UFl76RviC9ae1KIssohIdkFz75R2BO+ssToVVC1iV9G99vBHb3kmzLL1VAOl
EKl5R2+TPwVYG6hsfCaA1rizuk0iNuuCdCWWI6vC4y/IToA/iDTp0k1whLiByrEs/1OvPdtco9tX
o+pKBDw3hRqSCQqZprZ8lcLH/E/sDli4WjmRx1coi/NvRr/6jyD2KBdwKWJns800nwqYgkhzch42
s+iwEHgXmlG1aKgYJYNvDb7Y5dvmQDjagOI17WBP+n34E5RwRfYSXLG1ztvL7u428wMhVKL9OzVY
eq6tDcYfWKHUgxc7fHLbuDerlM71E63/6cbBH1/trUPnZZ0himZwTi9UPgwf3btdviZpTjmNggc1
RbzPXE+EVULMCWeVLmoak11FfcpSLd/ri1LAkd+lzgBskLFk/o0HTQM0GkPv/Daq8iTbd4BHinVw
beXTgVl9Wf6GlYlHwz5K3ktvurTO9QAuB+0RvShdR3w2+ucLoWROlaJSqFPibpVRPAE0RIRNcqpS
+Fglwm1B328XPMGN77avJ9IsPFdg6om8D7VWG3e4AJv08h6s3UGjaFMCCRxvtgHTH242NnGT/rcA
X6ZMyuwyIsQ71sQb2LbMMYWzq1c5Ifs2xyvSwqV84/Q7A2HOLG8pbkF61JB3N4Z0Mg0ia8rFuqmV
Cw1R99bTadC98uBKOxOYYrHojM/Yh9BAvmTOi8kqQr09CESxqruKAIwFcvbmyzdQq70fps1ZdQKd
y21fVzM8jQ+k7CXFSaDQJw2eao8H7UAV+M5hcROGSBgtjCUPN1fAPmjfyPaUyHYsF0LhcFdMMliM
6V5DikOlUs6X3cddBN6zmgilE9brX0IZQfyG0rQGcLzCtGJQ5PylFTulsBemlYUevkFLnvXeoaX3
gXXPhHVYvl1E7heuwsSYdz9BCFUMOIxP3Zle7wU0QUGqp6ljWsGQ23Kg3+0v8MUgho/AsyRCACG/
ySxumXYQ9YSszPHmnXu9mROrvnIF6u01BcQ0pP4RstRyQP5bxCovcAYySBqspRm+L9N9mBpGXTEO
Oe44ZWHH7WeqUmQqESwpF3OYYt3xVFuomltCckW4+LZtqeMygz12G6OpPrRmZRA7dPhvUMKPcBuM
tKnKAKci4CInj/piGvttwZrO8stGdJDPrhgFkvYfd47IgOdGH9L7nhscT+cQ0GnYr83lKtgefEoz
gY79t+vrBhdCn/guU87hKZUAZEcZ4ENeNlZ33cQXfRpRfMoY75W4Ei4YoiWF4S9pvNnzEC1g7VyX
ZZB7HwWjhijsV4cfd3/stsnvAnniEhoQASciEfJIhbJVl1k9zqH8ml2YvYYT14QDSWNyc8cUsJHV
0SFZQhW3SaFju4ijocx8DoXq+3+qbP8H5MLkQL54L0ETLrkROvuTFaOwLi9Tipc9d+kMtR/tVH7d
krl0AoVUqZJxwQ5ykYqfq3dXQ4J7GecuH/D/SOOS/7qWqPAKHRDS8VJhh5IFsi4wMm/15Wz75GTp
2Yp/+2GI2bzsJ7MoJgFldydLLxex6tppaWgN+97zrgyJV7T9RkztozZIojE5Nf2ik+nt7jyoI/Da
c+i+WjFuA2Qk0mZIvn68De8i9TjKn6VukYSbEXcoXMbeo8mUXrBUd0AENfcMKuNCSbZmG3dNyEkL
3Y9bil8GjSPlbJs8+JH65wcxMIhi7amZ0uwTrUgn68lkXn35buWmJzCD6NesAFXpLLpxRkHtNs5N
F/+52gsqQF2eNAGaFMU+u/fieLAO7hqKrstxUu2UWa3MoR7VaLdJoQ4pUZSivi5UNRN956RiFiGB
ZIufEi7JLfGq0N9vFmzSpvBqqbTYN5I9UVy4H/+UfqYy9HjC6ZbuV6XsxHo8vsmhiZSqHKy/K3Wd
qBX4coSo+v/AZvGrrg0zLPDKOfGlJk1SDO81eZ4KKpRpK5EvzD+yxKjciyz83KBbD2j2BVRiqu15
CUC6MmBkOZJx3oVB+nNsbJvUnWmlckSHUldPoEpF6kGqkL8zFEo9B2wbl7MRKUAiPccekifNYiOn
WUtIyG4DYSXDawyw0GhnE1wCJb/rv2FuS75QpKaH9ved1vl4xWfrt+2uMyYTuJnuBRC4d+lJLsSj
500RwQXZvKi/+N9WFn6UhRXru28HMnfnztNc24uTsdHx6IyXj9QQ5w4cmOeEzcODCcjKAsu1tO31
9kiVYzLlTBDI7LFDOLQi0CjSNEUH1IRGtOa0WiIQKGr6zstPqHnI9D9PE0NzhcXHHCix5kLwRXEA
dZv7fOU6oPGNvrrXQaO6gmlY25XcWlHLyCEULzpMajDI618BEedxUz/aNpB8wJIyqYBWrbnzRMCo
fhbpvV2v+HwYlwz12cWamcy3+JYmZetHJqomJSM4+3PevKdq7SK0sT/g0wDBYsyv+yyGgQKurq8R
ddrYa7z+svfgo5d5va9hTrmMz6BrHWi2Vvk3bQoZcSBKlfxsv4Pod09WuoVnovKNBYAT/r+REsbf
SjhIjcLdRqXfQTYASUPIBXj1gbtaFcVbbrQ69hAwgNrn24joBryYz1MPQAqkosuwYYiVUpQyNtbt
AqNGNP0CpVAJZByNsM0bpGV6FaKdt5MG2DCoV3AsfrF7WD5GSotBsx3nAnDg8q4DbUxc8MTm6Zfc
kQbnim3pkF82YDrssxaG62TxuQi2zKq/K8dKLPwBxFhB7VR0JegWaY5ND0+LmbXjg86v2JcxvJQW
7LDj4kV6TF3JjW1ezWs8wrbZ/p/5wzmYIH7N7B+ueKztGFTaiU9K6v/3X5+6NIoIj6htJZQ6KRX5
F7v55AC46UfzHxzXxpvkuGq1chOup3CA3551IpQV2HSX01cXuHgiOhTRkpwKYdqcQ1U9C3IBlb9d
23w7GA8aCyE41ViNyvHNhQ4gh/fV9URckP35des2gnnc1BoEL/2sojVH0egmu0dLU13Nqie9J78x
VsRl3hRCeFKPXcwz1Ap5sCPf6bFl+lU7VHMh8AMNonxZNOSwSJVEyIRpcQ8AN4g41fe0ABDdg6XI
lY41tGnV1Ajfq0QPXFpkHAevFlBLZqhO2CJmezVThvYx16OIOxgUM/d0j1ZJBmgKD3ZWsP4bdCeO
dow7BdBu6Dk7D8nngH/8tNt9Mt2SJoSMFeECzBDv1b0b32/Im961DbkRrDfbp7WN991GMSXh61Fs
OL/ItqMgBdwbAtMKRLrq+tfOlHyXBdWe3AYZickZ2i1YpQ0IqqwijgNErXIy212heLyFv+QM1F9O
wKJ2Xv6uXwqPb07wb+BdoQkQiadJohfsxFBFw+vSfbb2Oy0l+f7p9X2EsAI5dNPLnLDrzsZbKHIB
RTghs1FeMC265nrt7WuegANaU5WpD/CP1ITkfFxl4mRQYD53Cmn37rB2RlQlqa35WA6GS9ez9BoH
biOiGbHC+zsCidvmODVct70zgQODSz5Y3vWJKf3K1MvIUVo+pq/tygiPJu6zbNIXYpAH4e/Od13U
zZdcU6v0CtF87p3BrKAdoM3v0AnE2qwyXTQRVvU/WGlGcRV7QcBt1tf8rk+fSLiHnjKHyiZdbDqd
FGr/T0cLZbVvo49+B6tL6Y0I6zAEgXmQR32cdpK2yk+BkpcRipNJvDgYRMMLNZgJDwJjpiKKMSNp
eDd1+J4II1nFU5qaw6ugj4CSzt13L/6h65LGs817b6aRMpEGQYejnILr/hUB/HXvgl8evduhGyzU
2vp1pNaRpVB4BWK5Q4BeHTch1eSYWl9iGl8n9rWa1dXKeIT3KOCTZL7JtDki/48KVJR8vJOBCzem
65qpoKoDXZyB9na2wKGUSmt1gmSUdsLdoHRuOLcAICYPf0Dbd3XKKo6BcGwaftbNGdekRh+ZjAii
he5YDdl8JX+f4+TTUu6FUOYBB4gzYaj64evs6Sg4oD5Ghx9dCa4TWXl9+sOoyD1o+tIMfqLOEZGH
D32OFlZyD0uTp/B1ZHscMftXwJwrLMfeTEbfSLTHm6U/4GeyZbxFV6Z8JY9e0LS6onNkpaUFUJy1
hTU9BMfVw8WQ7qDxI0XakHoyqGJNDemhS8djhkKAbM00dDTlxKw3jScaUdUDWI8vJtTl/pBBJv9i
4Tdb268o3pBImqdmhEbKqVhdPFArZDuJA2YzI68sBJf9ROhxP7q/xBQuqKg6iR/wweSX3CPuAQSQ
27oRo4nh+mWdqJVs6DcIDRovVl3W6wZMg8aOdktuqLu+t4KHXgCtoMbAuKtGSOBuhBHXhqlQhPlR
UK0ix0JrokEOswuTP/g6xyc6djOtx4OdSqrgEGGymK3dgfZb6O+xYp++s0nBeGp9OXcXskvzo6qN
k4sjJ0TqG18RgRlwrkRb18XYBT3WuxbZmFGUeOG2TAAj22tnssqLGurtCUpb+VNbs86wi2R9grM6
godEjep6Vg61zZ7+OY7x8nX7n3r/kIhQ/IZzUtROt+spdY/Wf8hJY74SGXEFfpym693TGmz53xPF
ao6KizpLcFEHQHD9BGgHb4qwqBeMFqCoaHDTrQFXY7B5UDm5qF+LwLpL/7JzmBHqhbS+asd2q0sf
RbqIp7dr7h8WKdHCtwkUEUNkybUhA1XLjts3GoX1l2BvKRpegNIF1d5moUmqChayf25xvyhSwOkq
aifVLSjnTjUjAysXRBAgY5gAjNTv07ocrHyvGAc5dcUh82Amrvj+FvmrnF4EqpbB70+hTqngxfgH
6XuT3u4gg2544PZ/1aQqRxrkFdZLkEahZa3DwrBz7r9aU5poeGfQpd88yJ87JOsOC7XBExOWebXf
FNkvVgpiB+Ke8XIx+qv+cZFkgLZiXoYtbPq0Z1i4nR72B4LoOKBIaukzx8i+CjGI54MqP+jt6bgd
P9s6ZT1G9PBaSiot8Fd8DY7lGR7kmdDJ1dvDfwA+hbZ5XOD8pzTDJeb16IuAXPNBUKhrxf6fThqG
Zp9MLymx40aKhVYNPbhCOXkNIjzYmV5i95BZSJQ7CuTs3x4kCIVln3I75KP6gNqEvYv7HOCWyQUU
YqhH4XC/fr7APBAsqRc5sWj04bh9dUVEPmzf/hZGqIFYIXvtkWdI1YCXkRUYQ63kGXLsj4lMPiK+
WCElEB4Zv8BQhJgPun+UPMw2OJ6MPQmE7AE0Is8WwCp62ncpIPWnMG6JopQArgW+AaICrSpyfZvS
e7A21Zi3RxczcVsr1G2MoGkg6EOzM862hbSk+Llvl69kI0bGoHkYEEjMHfFUfHtpG2lv+WHKWgrN
gG291y8ShMKqCXITC05m9casflHf+88NcVh4HjsH88XkLDVihfVzOD55HF5yWLJiHKMoIT2lnV/m
vTiTvx6GxHgpkkxcGPM5epndo1JEKX8tHiZ2pCz+spqZXm7hSVGoByvDxV0zBtD+URQmbgQaWrWl
ASdb4ohm9QW6iUEV+la43QkgR8pscweRMyGPaxtAYq6pvyzGvCkNtstb24iwWceZHbsv+4usHi3g
o5Al7BWE3JpOTppLU1Pg9UirVWXTjVOXyUuUkUijxcLkwuzNaq+upe90U9+58eg5/LdlwBO2HpM5
DrpVcEK0pdZClE/txSpggLHlCRb9NUnfZnPPOknCw4cChGpVSdq7Gk7/9N5ZmJ4UyjwN/+Kfktu4
RiWv3S86fPc2DuruRplD4wvJk65+k13QleCMa7QgWrk9jlyiwaIIeeyNQ0LmXA78JwXOZOsVvvez
QNhCvLENhN6h0C8fyHp8jeihgMjjYz/ecqUoKSjN4QxGbZDsID+BxF18GxQJD5oJ5jFzKa0ORx49
1y3eqGogMxjqMOTkMDxN8w81oT7jMfgosjCxS7eLnpv+UyMnOVDUYLwur4Sc9XcIrr3eEP4WPcq9
XV+ci9916+wNLyWDSGjmBxlPvTCY2OiLzNzVqYzGCHnqU05ux22SMa/fOOLj3XGcqMkIN7ei/4F6
OEb3WvhA+po/kx5lXhvIaSOdEvyVtwdy0bwp1dLE1D5fOq/SzGS9I5iw1lSETEmMpL3Lk7UOx+VW
TjNARHTU/W4yUtsHsfCMqFZsFmS/gmJyZtxHVUdKWx/epcIXl99H3iwUlUWfXf2aMydWVMqD51vn
5DGcJQmpgKEPHODkeAaECOzAj6Clqu4baDveGXcxl56eBFX43Nnp6Wu72tUzLVp2nEqNicLgj3gx
mHuSDs6cUdWPQSXryJCnCOVOmLaS0XMCWodWAQyVSdK7FDYQdbJrrsVrKqKDz4/+PpSJ11NYFbp5
IHo1bASqitxE5bSc37xmXtnXEI5A3UuZwho7IYFafwuYTgRivSfKxMduOsnHnuH0T/Fbqfaz4vXo
ypyl6aQ+x4N0bkdOn07F7wOWqS+gL1a88uj8co2B3LHeHu1ckqgj9R/9rfDmmgGbhCZxX6PHmyac
9G8m5dSrxrx6wj/fih5ssa+THKR2jrQ6U3+Y0PlAV0QC1iTk4eYWdOh30TpGK4AbJXkl4v9g8knc
qhGcMPxYBt8dyY8arZmHaW5u/qwU05f4pMZP3+ufn3WzETttLONX8XA7lPziBsnV2jQ0q8f3wLYM
NyYCFCMPBn10mF0+xY+GdV3wriYKYgFRUfw9g2C0E3RK7fMsLP+FHHGgk1Dx2D83qQOvoRXGz4/m
Y4DGFluS8BSenbP55QAnbqQJ6SVgETPJUZg8udaAjG/RrG3eRT2qTnkXDngD+M8py9ELdYfSLkwt
psA4qIkBOfrpUDNV0ykPdZuvyagTq2/RxFouAu+SLP5rGA0QADhGCQy2dWO2Bub7/B/pbts1b73c
vMu99ZJRoTos1abNVC+Ejk3+ZNVRX/iFE6IK70z8sIxOhQIUEfmxQ8QDPR9WAG6GY6xJ541Sa6h1
XMcei5j7DgC6nLNn9FiV0WZ1m7nQVbZ5lEUj1E9ARzrH6Rz+EtVA6cH+CZM1shDO0WnF1CtLKDlY
6gHri0Y3oU7t+eZJayy08saHs/SOUnQCfiM9AuiU8wpSvK85u4QlHDHaDsbg76IvrCDt0TN5cYl5
+1HoXZRD1nhLVqiuQ2cSImOc6RXqfm3tbTj4Yo4ntljIdFcNc7QePvjdfXakHHJZgfU5os2x3SAd
waarA6OsRagX2Ny5YLmFtK6kOb9KqnIDdApU47KU+8zFY+Yi4ODROLtvqDjXXcOx5TewwDRyFw1C
Zc8K7ua5VAoMA0puOkkFep9Nxr6OCpBbqM3LhE/xDsAnWjAWUcjKYGZAhUqydDzryxZJCIncjh48
CLPDL3E1VQZqMQqTFFW5Pi8E2hPOLEznvWTLGSE80gb9cVUUQE4rqaf2E6frgChbdhJ+uRcnktCO
tvaeM52hvxlgYumoxrKuM9xiCT6soN8t96Lm50924tBYYLW7jW2doQROH9WwY4qPTRqcZUVntoSJ
UTp0jiF+/LQ/J+YuAsYfygQ8BQ1iJo7bmB0sogNIqk/zM2DBjtP1Z2qQ7xStMDPHITVZq2f0kg4l
IPY+ojKV+cRTDp4GJSqWflqzLP7nLVkd4SzPsoWsn5iu0bl9k+GK/3tVfwVOd8bptTLr7JOLO4s8
vztIcn4QS4qKEj9vagj7VVnvHYkx+m3XrgJvuu1m1Yz7vicjAOHNYhbOgnvOmnQZEfFgFPE3Yd40
DRumDPXski7ZJVORgGGThumAyRiS857jpJOTWL1Fbt3eRsFaxCYSq74utalnaDGrxvel/ZUUzzTP
ZIVsl1PVHdo69D2e8gdAU66Hp6ODuyXedjwRDTDMBFdqot0B72p5QBEMY1iJ3oCACC50AJpALDH+
dzPTv2bA4VQGoru3QbpZYXM5IIzbcFkA+8ovL/vFIoCO48zuLLwOtA+AUiCu0NsVh7BKy8PXuUen
xJz117l1Y9M37umnkHP1f8xxOr/0PZGTokGY9eK2LHArL6nqnexYnjcGlp9JKpNQrGcnR+pcfh/6
WMzujlYCW+4Quc/MAcA3Wid1ojb50C+u3W7lwJpK8PFZTGWL5M2W5ALP1dY020j50V5ZffjrpJ8i
BqdfbtqyGeV4e2KYVQfB9ALKCIex9emvXg1o+wo9q4xvjulu9lgUeojgCFxNLMA5lZzAOURn8XYg
3IdCTl/Swq3w0+x+gyPCu5x7w8jKpJg2M6OP8L3uXS25ZdXN8rUlebHf1TUTROcPcsr9l9qNcA1Q
E1esAbs4Ajsm7PCKXpSfl07s+9os0Ri9XnRtMSip10DNnUAPrhkwZ2RIMbMkZeM5Bp4EKkiGLKXc
64u8/i8kO9OM7fw41Nl27Zv6nf2Qb1rUfOcYm8EQmIjYcA1nQdE9C8NPiLBCMHIAue1KR20ZPUSv
fB9iyfpGZeLTLHjBTB32ymDcYmiktzR7mLnSplhVDBgrchbikIFzRgP5WVCCSn6sIIKXE/Q+5qT7
sFRESEADkfQvNSkhGBl3k66DBoRTCxVWk+ixTD/TO12qZuWFENdaYQNaAUkP6yzndz5cGM7YSf7O
QKDYQW0H3nZ85mpphbADF5nKhftvdlFBgsQE24x6ERF8CgGrI9/NwlzYKoDBW5AgucgksyOgiELL
+8/cgbRNxjKUVMIJN6taN4SFK2IVZTlwC30HxzffS+oSaBbXfIL+o8fRQYPFUt6Rxyrvm164p5HO
FWs+ds8w+ZZgM646CnkEu2MUhwqUINHxE+5UuMfYuw5W9Amdp5lUEXxMIfdIqps1U3m31i1pLSzc
CqBF4fdrkdJYhkOsHxg4abTtg5TD/FIcIOMnCEyUJc7hVsZCuaTfTgOFidk6UvI5zH5az9j/ovrI
FcKLJD04bsHgqBmjQi8NC93lKTJP4Pvt7T3D18tI0xNg5DaWRoJ/qMz6U+hOU/+qX5UtOg/M1cHp
HwndysCR7vi6p3zMZEBSL2SILKf5TDqPQMWIFXNDFRBQ9gAMF3jNDKgnTGcDbdobwUrV4QU7f/yc
V8ndAyTAtXbEVNqBc4K+rCpg7/5f+dPwvMTnGiV8Vt+Goe3KwX2d2tfrLB16C5HnmaPfcChTjpzZ
jfYdDAXCMjGRXLTLYvkqhmX755/vYwgDqBo2W8eWk+ASlw35voO/XFBBczxzQomGyT5ydM/RNnDR
gxEPgAtMgUyrgdJwjQ1FKom2ohBC2C/1VR4rNZiviJ4pahATR1E2JZdmCmSKPIfQkO26/+wHAmpt
JeIeg1+NJ4TJePuSe3GOBl8zmi79Y0JGY6EU8Gr2jYsulqkjaA+8hoTELfT7WEo5wDHZtE0PkQDi
Z0f119T/CNAay6RmnCadkbxzBstTFZ6iGasumA7Umaa1nHmBPDJASwc7Ds6DOZO5FFz2MYNU1azU
macfqXZbyQznOr1sMUSlWP1W+5nbntdJyIprrjDJnMhYX1A2gOaLnQ+lShNtMpHQvohwzZSufMNP
GJ8JXOsA+rCOXzGHIL2kaDbL8fcQzo0vyWz5df6hWbYKhsaoHwMdjNxwy88plAZWTOGiSBJYFntY
HB20ZfD9OgjvwaIOgqz6jOEQPzfBSUyRI46HTt+2vSVijuFo4b7x57Do4U9eppzAv3e2Iyq6v39j
YDGMqmcWpqfNWzTLyreuNhPy3B1XdRzewZs+xGhMDoxHxNlhr7lZTv9w8YDVLo/IGYls1FsYJsrj
vAnggM4JnPm7Bbu6SscMTwJyhlBx1HRjAXswY1b9xnY/GEnVpfxxmEH4ZsAMIC8eLW+mqPvYvvnI
/0XuP76kcCm5fXh5JmGjFuD2XIgp62eed7k1Y+ISVN/tGl1nxJGt89oBNtCUm0p/vw040a1kVBWF
BnRbm9uDz1X80t72m2sEPm1aj79rsUD6slZkvdenMnW2Ngcd0cimN+oKyByrc/jy58+d2g5qHAbD
z9tDIng3rYxYL/lPM+q53NTlJHDIuEJCI6kqO9hFiSm3MVFTN3a8IAHIZXWp+38ulfOSe2sIC8jt
CT9sTtxEoSqtsyAOLVSxCVsLSQvBKc2ikwv1T8nLMlSlHCzyvUh2oS+fjGgtVO13o6FG6217iXrX
mxc43Mv8zL7pZK3M+5hiiozx/hbMABh/dPe9nQA3N7cwppbySA7mmRMFamogoxS44rMkaJJ+68Sl
4OvN+ZbEJ8t4zOW+84KDV7GVVfxF86ILwBknu2cC+wuwbrjJcGV7//tdlo60K6vU/YaCiHc2j/Tx
sLnUBRsrcE5rYzssKUoFBY5p+e1ehTJxWL6cMcsEVnTaBd23Gu1ZPQSvg2ejKz8J/y+YGklc+0vi
UgtZNqSl/V49YenfeP67q01XSEIZzUxvIBR5k7m3IYaQYi+MRkRPNv/D80wrQg19cV046qUQNT95
gaOeK7jIydrX6iv+oRIXNHRfBgv30U64E1iiIsdYBzjEUZ0OGXYun8Nh9C1Avgh16+saOKQio6zf
WDPbp1efkM9HAmmf8iKVR9Qr8scJ4FI9UXe3kuAp07Csj42vAIxbytCXWWsaWR8dcc5u+03f8YcS
610epluggM+kcQkrfMVeVt0WJXEP6oOvZVB5sjLZ44p8IuYM4N9XIrcnYwjVt2E+il805FwUmFc/
2SHTTz0cgIsmLLHKP/RwQqdgR5rOFYoEUShfg5mEk0JNSvc9so9az6xx9lg4gMstB8NrMpeIl+0U
hGZHU4I35AGmduQR0BwPmKJrhb0/d1KiXj0+k4RaGccdq4OLIh3Cc/h1Y/nU4kd8uE/iCZMIYq3e
ERdbE3w4KvnhrYAoAbskLW9h1FupWWkTgk2X+Q+czlgSWb3C0DQaNDRnoVLJ/qU+2fwzRJElblJW
mMzI2kTJ6wpiKRK+XgCI14OZTQBzzQumxAfIyGt+bifYpo64FOg/Yp4IOPRxPMa81TCOmAXekKo1
OFfCNgClDl5eYDREfSoXkuVQiocmZ1+fnpccnvQ4U+RSYo7ENo6ZDr0eZG3yz7yOVvmpRmGu4jzo
QGzn9McPqxOQ7mnHHLKcVfXffeby/4yAD12MlJ0DTRsur3LIWNAj7wxtDG1uHhZnzED8pBzDy8Qh
7tqqWOMFSqBdlAw/iTuB5Wxpo4rkohMPOHS/GjDo3oewX7xVSO1HJOqBkaCasm0Vcy+a21R/COij
Q6gzITGhX8Kfn6+KuWle3pgivTD9LV4f9IYJXPdwzIumsr1K4W/Y4/lwY++MVuTMi0pLAB2xNKFD
Fv5g3prrLOUBqNgukYY8Rg06J1TR2xk9CQnmrwhVmj4YZlUulg5pRE2nL3sH8UNYLdj2ASqnDCyJ
MzQyStI6JL+TlyiH51c8nS/6RQU/LctW3ZFRrRhxE9loRyzI1VtF8h5PUeCLTCVxAOyfpWX6obnx
iqVNXAWQLihiSA1ol5qVH8v67UdC/LMCbU3Cdji+FUpx+htNER9kcoyI9LjA8NmeJ89dl2OZlsKz
U2e6Y99jrH82elfFbacIS+pYGXNe0hpyrrK1uGDr/QJ4XiI8ioqRxWsLxMp1jyHXn1C3dXaZhzn0
+UuXJeTiDXlZt4r3GUn9ntmwBFcQ0YOylaH3wqWMYIK9oJzLyQ0AflYOIjFQylIikxTQx2yZ6PjP
fy+F74zD5EC1LjRuVL/G3Fb1AC2lK5W0WUEwD/J0VKClGlnFqXHwDwCJYPSHr7RlhkxSUr4ASLjK
vd0zawhoVVfZZ2ewJsNRZqIuQpnU+56isjNwjoJlaGJ81uvcBjuFiyRRvg5O+s4dsAKz8biPULqh
SHDDOdykuFukV1TWhV9NAxeUNCLsRWq2RmBGRFY+pS6jvS3t7NKsG7muADsdxijKuqg71IG9RHzm
H0P6aKEd4cWMsHdsclhfCuT/OmBd0YL962q637IH+EcX4m1WpiIZ/Bu9n70Q9TC0ZqkATUyQmJlu
ugrv2rlFTmqxw5KB5f7DrcGlZ+hTBX0YtH9L2YHBstUIVDiedsQ1lFR1ZRW4oqTfl5RUQzWrbv0R
sdaQBQTv1y78Ic/0rP7JPTEIS2Huuvvr2kP36Wk+un++2/9VVNFKavlYlkvEJ6g4YP6BybyssaFk
BgfiVUzchkb/qV6uf8Y50OZw7299ckrgdvHpCoPEDmxkyLw1eZGIE7Uwo/DCHOxB4FCQSpKvQtQM
aeCS9P4B+nPhNTf0hqWCtGFDOEchlmcYSUWdIkjI4fQIi2ymmbrg180OA6Hy7t+nE0KumNbXO0HP
j1vHmbVrpATqTpNvh+LmGDHyUy50LQYVdQzvZNtJ/A4FEWhftJj2v8fMndGr43aoBZ+RQJpxgHRO
OnyVxwUvsdVrPAQk6dSnUj879hYo+mr3cTXWBsjDKorCTXro5XqVFckFsnQUl2f13V3+IAtoss4P
IWkaWVKL/9BpgxrDXVAhf6Np9CnymzpErb++PU5TYfWRJn/7BQdUfhgmjLWJOwE40jh2eUgBbclp
kb4NwaiiMsnx3ACqcHnEtLWtT/7A8RmZ8jXcDYy8ZCY3G5ixgWqPXAJvEnF5C2Vnxaw0yUvlquTL
5wwitkMJPN2IAcv6uKNzHum66xCx71uEmkPBEWH7sUn3pnhju/wY9SuWHle5RuTEDRkaKfykqsL4
7R4zbvLonMhkW01w6IOXqMTpI+WFPe+CjR7+OyGD++IrXKWolgGMeNSDkgrF6qZMCaCZH37bbCvw
HCJ1rD/LmzDHAePRWFGbzditx7Q8HCBIDxmN78/EG4EdhR8M67Whv1a38YG1x6zM2T6GMekaWXZv
EXecAcbjgf74gGR2nPUIk+V2cAV6GHeNHgFsQksnXg/K09tGmFZXdwH54aj3hU0WEaS2w3wNLUPK
9irsKAMvifA5VmJpK2k3mh8GKTm9AMKzg9UZQNgA/eBdIm5VKNn5eD/pw5OKvpf2fs5bQIrEY1h7
/dcP+5pjaCNBW5KFKfiS1ylyCoxnvW30/Yi+Z+eLCDJI2YTtNj9CKVFbDLhUZHm87UagxBx78KoI
Ut7TVEpdD2ZDqa19EyFhKTmX3I26t8RxAXmn5UkFNYapTIyN2hOd8lBbf3CvT/38TNdnORMyGBfq
1mwzp6cFkBE07CGuYHMYk3CaafxMv8fgVZ+NksuRlnBRdSw/5MXON5MfbBZkIOp3mrAyPSBcQjI3
UZJhXcXaNKx7zMn/aaevz93l1gAao1Jpui2bjrAPz//9D74GHHIlS+PGFpqkKxpo+o9F3TtHYstk
9usN/xE9XtCTmqzZN5knT8NliOwWZA9d/zXtdnTsNo65SftdjQzfqObZNf042Hk/2mHG7dRbQeF7
eoAz7MSytIvclA9+z8KcHqoLiuZGxxRkgbRZbJyLN8ADqddqMsEZkHfZdlgF79BDPz5GXrPei/vW
uBBWpzad/ACBJeGGggGWKrfLZzYnuEic6aw0APhWdUC2XrezrWIPwxT3E0pDHMUr9Sdlwd0FgDQ5
70tTkQFWHuhw3AUeagSa1Rk9IOJNwCpzS63Ae+ZAXkf73QpcLj9WDkHATbK1Z+U6facXwiWmN0j6
vfsF5UZUdB4aLcLevNy0dTCUG7Bxfrli0Qn47gQnh2XkT/QPooLwpPCwxRt1VlNRFYLCqi97lMl7
f8lYL+vg4gJ0rpDPFDYR9gxq5VVIN8dKNkICAjOwr+JdfYeGU16GkLYK5D8+5TCw9d+6l+/ormFy
raEaXNPvxXX1arZB1UYFlfS4oo+XDdrhTgPpJX4vHCxGEsCnZtPooo+iXG22NvYvgCQTDllIVhl9
pcY+Kd8D9qNgIqVJbv+23dAgd1UA6rYXFNULPvLXEl6pTzm2Nr+rYahMMKdoA8C8PYBwOiHcVNG8
daXpFtc9RTM5nkQmwMq6vSPB1DYTfreiOwYW6YWwW+0klAKgf1tSeUGr80yRXoU/QsHUF+I/cRZ+
ZF7mnkIqnFhoiqSCZ3ZsOTiAzb0Jox1lGzL+UpBbK8xfrgkTc8kGZ8uVjsYIHahAfoj3TJymeOK6
9l7Y9tfpZJBbjeqdEaEivIKFW010Drvo9OW2ecvshAY6Nu06EwbWKAzo7nKPMdl50xZnOEF9WQh6
vpkbQbV4yVWF4ZC+ZUtfZMo1/7RVs8jiZsSbNer3i+82XbzX70nUPsBCwYNzvjVjBvz2BtDSB9KK
VgV64CRVs2aAhEvS/GVu462BsQNbESNcNMP+263aB3yp4gYbu45yh8PCwliX2NGcX8tOu0hsRqTp
kNN/I/6OAHL2WLRVNyjJTh10zMxaXjCnsKf6NsTvC2iQNx+QzUQ2XTEdx9ZpwpaqUSNI1GWVaECC
MaEiSHdV+Xo8eNczfSLFN/DJNsN2WUWQAcxbVoEyDpHg+oH847VjE0yRe5zOiR86Cqen/akqkMGl
SWBANklfEygEa+MZkXePKQJk3e0SGS6HkwVVS/FtEvsypd3EvJCPyLmZ0K11CSQWeJMigfafPaZd
XqKvfaB6+tkG2CF80pQcxzQ1ca3rfgcdTDu2D+YVsGkBIyAVQdRY7m6Wc1zBnR029JfPUlp1iM6U
uxEG6VK0z6qNAXcX/av/r1UBK7tsCFIIKhqBMp9yhtLcNoosl3B5oorFyH9nVpO32owOwztoSiAN
DoUk3WxP8goluDUnt3wGXrdC8EBW1G6rETtb7xaM2z7iMwByeBkgQTyVYmZIjDOUr1qBUg+TUXCc
+1DiT5JVWHaa+nxzeORfCX6HLp38zdXCEt2DS7v387qy6IVbW5H8SUM1WPXcy3yEwO7bAveSUvfB
Ga2wMB8BUzRaJg0MxfLQksQCkCgxfSerUfkOgGVVCf0ZlNmlKXbCMrneaPXuPYotSM4MoxOIAjm4
FtJHJ/cIPVc5iJzKGDjY+9KHOsXHsqsY8INZp7+V9Hg7x/dEOhA4uVeSgt0Ruwc9iNVqZ2AG/rB2
5kPESsx9BzVmpM/p7e64ARZ5sgOApFZl6+A1Mi/W97mSnWmN3XziP7c56a8y7rUktZ/uk+6foCSb
B/JdSuDnO0GtmM2rTYEnK4QbEGb1xrBWlkRFSfxoDEDYhPg2vXeN45iX5AANFtu7KBJSue8exmFr
CECRhklMHU8In8BKilnchX9RhO4/zaPW3ggPYGQhXuZwtqB/i2XqGbnvBvlHQooxlFngfgVLrJtL
2Le8PSUT8uBdwJwsSXmlvMDpdcaxd6cDBsFYCUA6QQAolUomn44uy6sawPrrLtb7zL1+PtqOGY1/
Jswe2h/0RX8MbbvtkV5eotcYxJr21SPsm8dMfbBN6bawuDXV5Z6XNq8+c3ICN0M7uASFjQvepaCe
FBpEmX6IcYSbL23hNaQde/XA4o6MAjra0jyMoOqQzO/c81tGwDM0kdg1j7YRMus42yaqC4p0RcxE
NRBkE1j516ZpdDfq+OjK806aT3/2EBbaitiTwbu22HAhWSHFdvAUEhqlmwQkFlkifWpPPtcI2fnY
LAZ45iHoY0xqQp9utqGw7Bow9Ang53l7k64qQ4UKtPZKiVLFaI7PH2JMpWkyH+Lizyf2spB/USUa
UAJrnNKwdlQfDQ8gqnlGyQc8XTGZUoC6xFqr0RTCBvKNQEvjTIoiDod6XI7kR07H9A64u4u4ZD7t
hjYjRoqH25/OTogDoclxbqxw+7HQL9hKfKBURJNFPxeEs0LV8rmxbjRWa9YT5zBlbVxmWP/W8jXt
98fGbiI1eJscFhBa+BwoeqPQGC9QCe9pEvcJnMQFo8+pq8+yzks2uX+zeBVbGwcAVVg+loRjSi9a
0r+srrpgdmqM4JCYT62I3j0BtnePQAR0GL4DBJPMPX2uLGtiUCmcEZrNf/GHay5vpVH0q8qHVEw0
1Q6wkRNYvjojJBZCyVYp6xKVs6iWAVnQAT2M3c+uo4r8ewsxXCCZwGsxI38ZzYYftAJvc80J6fqC
ttbkyqatW4XLXPa6sYzGrxRUz0QsvB8HfAW32SOy3TcISpxsNmRSubXHULmXqRzbYem8gXTa0aH+
WexcRM8+0CIU0hSZXgi1g4aKljY/rqirUSnuXpIMGThujGGeoNqOPxyUw2nTh0hcWsDxgyDdSgfr
k0lSKtNfuKqAvSf6IO3B6/j8aSfMzhuF5oMC0030ifhM4C7t4LufkV/37LHKaEddZtWlZlIcoHY8
xnwf5AX+M9BylPcgO5zCREJCOnMumES/28o7SoyMOGQ51VhCg6yDp3JnwW4KZ9anzsSNJ8m9rOTl
LLfdZ2mrQ5G1NJZslYb6WZuIkCx4K+g+5xyLKk1M7Wo4alDcS0zC9oDqekk+vdMyHYC1miikJ8wr
yXaKBDpop+hxmpglbhM+OpN531ML38s+j3zTicKA0rW+/xMujll+Z65EsPy3pug3Xk5srls25oiJ
Z9cCYOANMu+WcXPe9+4TMbDO/6NBgd0odCKxp4taRMYeHavkFFiIDWVFTDTCbKgLJshF/UuMdzkD
LvZtDgIMcZO2RUNKM5jBOcvCFhqd1taC13h+KUHJdypA1fPVBVI05kCP7yLP2t7wcDGAotxkSm0p
BgIbxerAUT4JfFh7M6SlHkL9eKH0fcSP7H/NzzC9jFrTFlv75us1M52t/65v69KC6O12LHzHa7uU
Wclv36qf82mO07d0OruSwG/lrq8Q7MHK5FIk15HIzAXfRm8Z76gyhp7Oyljii7eBgtWH64xvyOWU
wlct55hVlobyeTOB3LUAmVarf4/6aDqideENi6OrinK2e+WWKuSP7kPIuMGiS4e3xIVngedIJsF5
ZOclbbpo67uuqHegX1k61p3kdjC97XpY4svCRljB0YK5yOqIPDiQRXWx4JRmsM2tLPgVZ+sziKUt
si9U2RKsTU0aqIe1zYqC2ArFDdz7MUCdnx1omJ21SIBzRuMJHQ/OaqKKLq4tYNZYQHaVFw1WFug/
LK8+nrfebsJCgKeg4wf4VUVA3RuZ3XM/3RpJGz3ofg7/7BBfGEfSF8L5w5pzN0Rhr3U42Rn3ZaT6
7nhWQkurQM6q426gPcN5nTGi/+DoO2YNm3fONyKjOGtjZZLPFOPMJK454aiwkzLPt1VMEYbZeu9k
OYA65hld7jZ662n4U+s3JhZiJAXAyd6wWIrC6blqLMJMfYTWEnjYsoZMa2AM5C5XYEXq5SYLDNEg
eBXUvxshqaBMc66PKzqO+1WkuLeZP6kZvjW30C8jZ/1Nicrqc2aBM3m6MVWK92DS2zMz14PiSj6V
/HOhC+jZWKMeGdUa2JDsGtpyj0i3FVLqyp2K5HxQsPosc1r6wu5pyLWKe+cQgViYP55Nuuq1gmh2
jWqOG/Fxh/1GLafWzsSAE6+D+wxfPZcgSzTU5ennP3KRjaNX6/fmIIH+gtdeItanFNIZfwopsAnu
DQQuRDt6Xfe7UWM0CBr6WcF+4cSAoDC5e0oBZ2DCrjsY0V3klReXuK20s0G8shp3uXLPojKwOsFg
zDBU3bWyl26yuWKseIZ+u35+hdSHNDrAP4PzY/QULBvyD5U0c0lNy41SszurhGIhsnNoNFGNG4IR
tIYMUqsieRwZLr5xU3YW82pzdiHQhzc3U3NRlbWg/zDbR5iYfWhcqT6o/4jn88owfrl50qVfdiys
khHhkjen6OahGRp0v472BhiDKjDJmk2hd1uYbsO74ASNVEkftVXewYD7N9p8dpGjMweOiUAaQ/Hf
YdJqylapWnAux9I3LJYdYbQwfrl3cQO8sCo1TLjcipRU3IPcKiC+f0K2Glo1EyPtxwsoLLqhXNBI
EBOL6q1EJWWjbogeeIhodmghjDR3bvc59WjU+YSz1y9DpvYKeagoqs9+t2eLlOKwTZHqxDBF2EwQ
IDOLBaErf5YWRiDEYAr09GpCb8YMbKBT34AcG8Io7fp11S1a9qLYxch6SewurDTKxS2yIqe6/VE8
68eLpP5VTB16lCmh3yhVsLQEw9W+VJV8cwPj90VFwhSJ1oDWk5taNfWc2uOCc40jc6uvawd2jx+l
6hv6v1ZAy5WTOF7ZmKobj+b/5dhv6n1/9+50zwBYE0pUDNsP5ZKBqeGW97uXFqDmFaAvDX4Z1Vgf
j5PyGGaO/8fdEqwJmCYW/iDNEZhhf4bBEJg/PHSy+sq8TVvMfnG3HP2Y1EiXPJQPZZVLJCx2pXjv
4jFEtJeMEvrPIksYMeNVMCC7XXPqa4HJiDCcZ0AVy9EkXq7eFZfn3eRJ5Dfn6qU12rPHf7EFuiGE
9GfwD98vsl+cMtFH8DiFdCm5zQWfB97i5w4zqvwtCYQB8L6i9cFNk+w9f3PHvMfxKPRDSS03teH0
WiHtgKtHeZv/HL1SsRNh/Q73R1+7AW+IFmkva4dDcPc8x4g7c2tIzyMvo8Uvrpz1U1DWP0Vs/MPp
7iVOmcRha/bxav0LAKQrekoRHkeh2LRl9RaeB4aln+Wlq1iqV9rGlgOv5X08YyVMOOdeXWyu/jiz
+9xZx0oACDcklHp+YJ/3UIPFFwB3DKY4NThba6TDBDYML9Js49bRw2AZLjDtebDS8HNyVdMWFXZC
5IK4dheilBLfmu0tqoMdm7SWspHa9J1XrnTjG+i3524fRiph+QmvEyu1Bf9Un5QJS/aihwRUwymw
rjbtYBZkwhqtdO8YWjxAwa67PToo07tW8GF5oxSVjJ5lW8heY/mEf1Sc7zU83zBQrjFF9Hv4oE8H
nPkR7IWOMR4+DYLEDvtHRwaKc2vee+M4dtnGNFtG5ECNw5tZdb+R6WtHL9gqqj0xzwTHMGbyzEQ3
uaeEseQ2sqprdJO0xqJ+S+ecFHGpqmhVc4ZVU7eCmZlWXA7Vll4pz17uq9SY9TnjSFLgss4wLs6+
hKe0EQlatgvE2Tuy34geUU1q12JMzNBsjd7+FKXk7aD5opBiX/NgyqqkvkG5WYbuSzZoczoe+eBs
vczL8EiUVnBpzgxCGzA3ZKh3gbjs3XDIB2zQ4gY4ABJlwsH7sS/wZd1Ulj4P3uEN5PVg83M49zhp
e4h9hSe1OJ4qaj2/uTrlB2Db8uh4ioSC4FcBRVKpki7H5DvM9wDanJtqjs9dGLaVKx4q6eGy8vhe
zGOhcy9sswotcX/W6/WSnx4nNWbt1sdQwTRugpsRZkku8PwCmwFkpaoMYh9sILpRKJfVdRfJN3Y8
uuUvUB1nIWUzyYlKa/4iR1LiJLvkDJ/cgUY0Hb2toR2NIYp6Y2ZwiJa7gTyDVhDzM+5cuebVFokw
COx5OHOd+FilFE7HICPUrlOAvAbVrFOYWW20rCe0RxwMCwtvUdbSHE2vieKaor8fGCGCrJTMET2R
2oV8FbvbazIQafbwi7pTX4qgVqK2b1CsYYD1inMXjGq9Yn4jPTIlEX2vNnHrB6VPHMmc887AcJjA
IKvVy+2EjDJWRtw05XQY8pUG9vkjVrkW6loQyxDFfyh2N5M6LTfOpvb30Epe0HoniG5FmxSMMZFh
jeFH/zExMMiVhPYjpm9Bb+RPbn8jHQC7ck1ubiL/W5NimZ9hdjgxW4Ssms7S/UhsqqtYQaNTOvgD
ZWdqG7RGS6pF8npBHsSj8I11E46D2P58XsOyTeNOFWWLj0jPV1g8sKn06jh2OqnTBm7Gd+SmhMej
UnN6f3KiH391Kqztu0ToR6/OofoVUEQQ5SGiOwSOLB7H1yfsByAJCE99fbbwcYZnDCPy+koQ9SBL
vOEqNXriKIT9wzAH/VmLFqfkB/wrPF3QJN+IVWiBZDFJUwgUsSZeZQDT+A7fMU+W2IQiVnz0z4AS
yQ3DCCZl+hpKeTblMRB6zwHzWL5XgXoE+EHMHH1f1ngU8gT+b+00I5FWnfb19eetFbgvAEOhaxTV
5ZDNevN8hzrQrqvVHiBqH7XQt5+1SG596QSF5kWGRXHzviC6mHBME3RpUSoZkNdjHeJ5oJ4e9B7e
acRaJ+N4TfXmKHb3ZCnOjJdY8WckSZUDhyJ7HvKCeQ6Ne5TKNbWi5c//ulfh8jtz9gfAcmM74nj3
oxStTWEy+2rRL4SO1QNazfoWzM5v1WWLMHyBbC7Kh6A8EKqCZhX6/M49NHgNPui/DcmtiU11yuAm
3quuqlKG91blS2v2FGfslDps6VXhsB+f/W8g1+ssfB4UH4GT8qXgobTNXZ6AmFv4kqCuQJTKosz0
lXgPkJqkFakOQMspaVj7XhOdhpsqq3RbakSubdaemNGUh/HJPwIg1qbPacgQNtW/WGEthEU89x8W
orfI4nvaXtrsJdDEAos6OnXznExWEjb9XDkbaUZzeZhT+UqydWSkwuYjUKbK9iTEZXeipnu3B1V4
IfEO8e/vE1TN7qDC3dbJSjXri4lpRPD2WSr1/QPYAu8Y9iQolLegKlxJcDU/Y2I/ZUQ5mNXxcofp
C5lxUZw8V8xHOIz+IqBeF/8cBfNQkNe3T4hWc2jqCoNX1MVTBv3Hq1/tYUmrHBHHXEoP8B7Kt+ds
uQpsPkcZ/uryFTdRuhvfp2wHCNWY7GinNyJVpdZDwsixE4s7ZQxRplZx5HyoFLC1J8fjYz5f0Im6
l4HA0H+uPpVPZZbNFLxQhIywyeGVP/Huc4rjt3wI+dsTV7a+ac5Gbcb85YPSCV5wGjuObW8XU/9s
hWhyBHTwJvIxBJmRe8vfJCdlwbcOfnLUo1yQlyl6hdX+kTIxtqVzDilo8tQwfZ8PbBRiU1u9cVVi
VSqzyMPRSBCDNQwfzQ6Tg66QKsnuIipF/6hjDie8Ern4P+UsTDjnjk2OtmmvBG4/H86EzySHkxq6
XV5aKp60pL23yeqfD5E5PeafsDbyacF0eMAJFVtkncCnje3I5XxvdCyhmk0PbVPW1yds49+in9T8
ZTdxTX4uoIeDMjoEs7KmQGGija1c6H+wNM51eZYbrwKOthttJsFfwEFZaDdyOFQVYGUyhkyBci+k
fyuc36wPZcEdCwAz1uYQeyPfRo7OmXJm+u4AESM0F2rq0RJqRGPGghwSsh3uSWy50DMDYB5Yovkk
6vsNVAi4GnJeGER3j1v2DU4S3Si9ufVgkRRuP6dpAWHnBPQLiGm/tbjZ5Ui90B89HIoVU7cW5olQ
a5Yq7pliXgtJdDOpeEFu/jqI1E0E3higBGERroUVRJfYJvpsw2/Eci0QowsXUvkW723nwLSNqMfj
jO6uG3Z7uzVnXU12D+CoPnEVbVLGhlGjCB55AngKmotwYhLDhMkjqQk2utl4ndVhEj3lI6kdH4Aa
xRuvM6sevn64zUFJmPen7QyLn3XJe+enrpzI0ZWzvS0peZKMDzGNkCvAXmQ3AxgqFF8YoGTJraC8
lZB3miBaAt32L8YfiS5/bWrLfzM6GaMR4eWkLZly6ca5Y2tweqsoI6EGdQqpDywzXRvGZqKiq5KZ
FiP8GN8Wjp8Qi+c8S3Xr5LX5qrACgEGnUSNqRd3BLMSH/VNkpi1ABbV0EBo/NCPJ30zmh5jnWqkU
PGIl8lsREtxOBhddEt9rCsmG2C6FYe0W5r7JbNf1FXKEtiwZwWVwWRHFOUMXjH3T9LYPZPwqBVIj
wWaM8UlzFFsG49xUt44wnuxdkLUXs36YFzFiAHFMEXMb5uIp+9CpmxKZ4dT7BCBdx4ZbTQvBPUBd
Q0q/SwJSQyGJGzeqd+lJrC1sp9Z4fRM7aQIYEcINbFB7b/CLmLPcmZxNlROAY8yvlbEQOj8R+tsL
ZtLvultjtaHY1l1s0fFNoID4eKZS0UGBGDpPBPdOXU9H+/3xyN5fB/5M8o8jSIMR6RIBXnscnq8N
MEJt/0LmZqjGgpI9jKq0dnB+fWLwyaI9VgF8KCk8c6vuIQjWSdOa3+N7ec+t/sGdEM8k8OSqOdKH
IHpwkBfNPV6VypoK/WN4r0FcD1yPYqA17ZfmafH1DkHphDc1HZQlB5Kd320kodkyO3qOkblu5Qef
T5g9Wb5EIJ6NqKQNdr/M4679vTyXJWg6TSfdj5tBrwr34IDXH5FYRVM/Dl6nhyHfPmilnArsvQzc
A2sRb6xh9LLanTa6p9wfmkZz5jhnT8/K53nUIxCF36amKysYnm49O8whnObiPL2md4nNiaAw1nL+
fIkjf72v9txMvIKqCv1yC5dCiub8dq/hPjhBHpqkqKplZlqBi+xTTbFf8BHSnIdIPrWJl1QUIuSw
wx4XzH9sHR8cCQjozA43qcUa6y8DQZ7zNkhMHnWMLncUR7jGEIkzNq42XiiPpTzgXLpIsnALyn0V
K0ik+uDkGPJatqU1JrgJAchzQt4qr9J534dF50m3S3DN5japSVgjSoZR7MCnVomhBKQbTQKQ2bUx
DFcNg+YKZAHvjoJk0H0OsWCeyx8Y6cyyjzm1QpU9jC5x7zwyoig1Nx8HRk6LzP/HO9fkeciJg4c+
CRDyhruGyu/IwIP7zxpZF02SNX/sO7gX5FGcRyxIfN+YxCsyZO+K+SlMn7sNn/jkOLb1QCTLPFEb
znn0t56B5bvKuY2zvCodF779cU8ZsPte+XZUQa9kiDBc4jpjNKTnm8TpANJhHtGXlbmDVPUKiB/Y
Z5IXuEznUAiW09URHxIqZ8//KJsq9y3uUVnQtv0fkAGmNa9SVtmEd+hCKUzfA4OC6Xo3l+msqZRL
gAldMTDuQ0OTzZy1LP713jIYgQewoV7V0pzETU8i/+4RcOC7WEAQ9OJCq2VDyTfiTYX5F8AoFiuK
+JjOvJdMQfjEk8Z3kyS8jRQROyMO55eG2LxCL0Of61tffUA9ApnQbIDxcd9hXglCXcD9v29izOfn
CeTOeBvCDGy4qy8s5askYfXslaKYHCWe8MKFUQg8dKqJ1kvzVGvqibPcZTblGlxDpAw/i5NxnG2X
Gvp9DVFiF1F3Gnd4YdnwqNHvLStA0cZyq3GlortCEvy2kEZn0Sggac+l/fGGGZcWNDJR4W+JGB6l
PbOtA4XeEoKau3SMYMjCyVbvFz/3PlBbFCHbN6St0GYgYzojvBj7hiHqyYaP/zdeUtN5KNZIqGeG
ariqC+tPPSQS8xwxGFRkxtO4GJWSpY8PKJB7HKahJ6h24c6ZsDhm4T5qF+dFTs2x0nj1JBCbHISf
WyZvkXOHMAcRI4hpYK8MLaJT8fdQg4/fOwBNWE3bAFj++6X2FXLJqJ9VZAwSCLiijO+qhCoQW5BS
8JOB2M9/4DX1Puguag1X1te+a/5HMDfb09D1JNgG1JHOG6RGwHMVyp1SFLpxpnctmvXM6GO03QAU
LCai4SXeu0+eXQDJFL0/apEfLfM6ieRXgxQE+jBFrHaElcKOogn0fRpYSmmYTHX+YmvW0Jdzznyh
65LugiMYKYv94N1qPy65kr1Vzp9uXhgOgyI790AOs9SE6I2xr49sad/L7DVolh5A1lbUHCbB++jc
YverJ4OTQ4MiujLsNmqtqDE4GlJccw9lROwsvIsinWKssGnrW2GCoTceByvvABKD8QOa2/AmSdJf
yN/P45XzgQ94IkqVsnI2cc1FxxfPq4KpQclPV5kgqa6oj9g/CQFR3JVV2WssYoW/xGr0OYusB7v6
H3fycas8ERpgrULq7DkGnB1xyE7HgBvVYT8VTusG89X1yFl5mRlI4pZiaWiHOwIh285dqOa5EFr+
+U4kuNc7BwT7roNpFbYlkofJY5pVH7tigoTROzTw2mM2mJxnXr7YorU1ESCxswOatcP+IVL4kEtF
l15p3HImryZifWXN1v3SnDmXaR06vBkfjjTA3cNQDllu/2jk/mcE2TlDo6d50FAXiA1OXYPPiC5a
LzgI34WDRoE60D///f158RbIP1xTiK6EAi6A1mp/ZgQBPSfh+uDuCfV5XUqR+B6Bd9BvHRAhI2aw
CJfgrFihcAGoLiX5qcftt+DEG7TTiTU0ivcUsr3iuvYZdhgZ0H5jHIOSspJ0d+d/QFw2qUMIgShp
MQkEcRD5x5C6PLk/y8kAwDRT5l3o4gdcIZbs1eC78A2FW8xhpbiKr2UXats43iLcxea8s5/hWk09
Asht5wAXZWwSoq2M59toqGiPYnrVAqNHUR26PRqEPyIMul4Z7O8lhOBbUR1aIa4KYjCF9UyHhg2m
i7AkghGsgjhY/1drt1L2H27t+rdMsr8kj08OsyEKGgMCc4/f0/VW+RK/M4WFf4yxIoW9XxbnDOe8
4MPlSDFEZmXaN9cchk+fq9P8rYWUu5em7ZdUqkbm5FR4LbPxhACQOboO7ghR8gQkUutNMzvFXtxh
ScGUfgdDjz/E67P0GIWBEzOoaouneYM5RBBcBGNGsUHonfo+PA8yMdB1Yr/paOJHGrtiDSAj/gs2
GbnhoTBg0wE2zmQ7RI2VQv5kjyCyuh5gnA7WEidxnjaFioJ5TpY259doOD9P7s1WK0rIG2N2X70/
nfr8vSc45cX+6HlIACdpG4QZZ428WyxgAEwCa+H3uljf0nJEjdYtBJb1HtxvJRgDdhZfOjEA3BOD
jzzDdo0qMqhFpZPeTj0mz+T7dLG75qEDfghU0CLzsYTLe/y9dGN7KJ6iLjHwYHkbipJ4do0UipAv
EY/zBXIn0GJWQXUlGjfCU49f/xo6f+YeIsHCzlmNP+hOgOKktYDT6WnBiIrgb2YELCcoVJtWMAc3
Tjx8ibn4nYkGneizuC/1Gs+QBtHQfAkBpszjK7joXnV6+SbF2k0hlsNk8F13LDuU6TVc7BO2HIZx
wel6xnVJp12IHGyAxZ4hTW9H+2F9rEshCbCsnFX4SWfRKwfb8zAtlGwXnT25+X0uyxhx68JEhK9k
OsXZVQibKXfmzFKNJhrAoDntSMxsexh2TbfRAfwpOJqB1DekIslWGusX8Cy9wbOVZXjhSmv6pF/n
me6HU+8kROUT+cE9XgjFF+BW6FL7OHRMNqr0Xete1Ew0M9qCt/hofYi/Tg4pkr7R+jKvEdJX/Lv0
c177QVdzubX4j9onA38UbXzs8+K8YxDJPpJTza3vLXfucIagMNk/ov3Ro/CMQr/pu11FLzN1fxpM
M8BoUxdlmAT9Hr92zH4MyiYy9wuaojDNQyX0N9kJEHhJATEUlRZVGi4qS58cB3Jxzv312NJT9gCF
00esk5TdloQU+awWxWbtLdr8i0bronVCKyD3MWRCcXXVn2dgfeV8KVdtNRQ3L+jHWhoQvApays8i
w4VotJ7dKp4LHU4ImQKkBED02mQwo4kzVFNWQ3Z0OKKJWmucxbN8a2I8UwdHABSH+9Oxd6E2OtoN
+pqsnwrCeUMzOCHH3SJrAGlVyVJHKHLZ1YHNx5Jg6vv7dc8l2qwclwVEAKRZS+le+cFvsFrKZxkE
bCDZmIq3QVDmJCxlSctpU3JB85OQu5R5VZMadp/7c0x+CwUvJHOq5wvZ8dUWvfiZoVVOebf6GDQb
+KVWFUU4IG1eKJl2Mgxfg/ZH9Y/p4izm7x4DojGWsSI1hMFDEiFpAF9abuqwVYUEpEfMu/WShhe0
Y7POyAjauhnlWVUOq8/IfjsbFnu63qP1eDPhR7AaHmS2Zxva0ht/tnDsuUULKvhkTvQSGKicvI3m
4rik1vDdHj+QuUwcgPLcwFXLXWgYcfgpXXX6PGTNx0dDpJW3KzguJD9ZnktD1Rnb9x7Hmcpzx79n
BBc42lTBlkLJqxfRvAQuKMnP9tuHiVqB+hx3yzqrXjdfg8RgbtzM+Fmo4QYN8d7zDmwpgoX1b6nc
6Pe0nwWUXo/nIR+AhBcIJOZPSyN32OX4z1sh5C+c4YltxeJUdi9jqYLOnXrcXFNAsUdQjfpGRLBL
PJkUGSSJ25cqzqU5Ry9uSRhMtofmISDebufGj+jQF6wt94+dGfC+l2HtVXftJh1T+drL2qa7Cr2f
K9h3ERSJIhI7M87mwr2pfszcEW+INaU4AXWaD9i5cn56n+bj67e9Dqhfx6tDAJGTf3HmUUtqQ2dw
7nO0WUqlB+5YyNaWDRdOy3Py0t68Eg+fPW7guntK019tJXg7JnEcLThZcC7MFABFgxlqtkhQhhxf
LHs0O5r7zikpO9QDC7SNsU4YSksCDfSIC5g1fneQ4nOBxRH2ABy980KcuN1YyzjLQ/jSDhxSH49z
LYv/rOp+UmlyiW70A8rFrs34928myfm9KEWDu9+KSOXmrPNs1A4DtVchk/J7Ow7ZTXzP/hJfWtb5
ku13aCUSqacUyZMfgcU4W43sTU48yvHJ6YnDDZkaYgZyrdr066W8E26nPlkuj9QVrXZ0IYjKiw2z
CmUa3A4hzctSbNTDiG4pbi0stPc7LSdHVTRIC/PbaXDmOIK3vDdbtPvqiKSCXtN9CeReX1kbeTks
uRhmYhK4cGYXXWTRrZQDoMov+Q++zW1DqEnwA/lJMQk+hUP41y4FWtTShR1gwhs4+o9qVRiSFVue
npwfKDFqPj3hnIk+8m1Bep3fV69K5H6YAU55b29KFw50LGCTqrLLbG63kuX8UcsY1GWe4RSiTsen
D1LhWjLnUjkzJOGczp/dHkK+CVkllsKfM2kjrPsotceXkebi+nTmCmNUyof4cisq2AAQKebLyovZ
RQyLQgLa8LpJPKFkYgQ4k+8sdnzxu8TYUXuH4HZHpIM30p87Dc3ppE5PLVlyA93wqCfF0Soo+TUG
6gSgld/BpU/Xj/wcoKGYOvvweui791U3sc6F2b1AA15orrXg2lOt4InlqHS2jrQNWuVwE+BZl7bI
AzCXKxLlLN/Qm3mO3SRwp3sSdZclWvN+uvqFJrJhI/l/wmvqTmPUyy2LAk16T13JrX47M93Pwof+
PYxi1FNaIcjEHfxs0owCHJ4o9c3KBpDnSX3bY6R8eln4gRrfZiMyP2qDTKn0bx8JcvP8r6jRjpYZ
BuTIkmJTICc2OGE0EDMtXMnDK8uHNjPVM9bzvAdAWDYyf8Esqbc/Yuz9Q4YuQSDbExKkAsMaGhBO
qLdIFy0ISR/jhkQSeV5l3igXs7LveZqyfcuC3+MY+svZn4bWhpCTzwAw/vxKeHgq+S6h+IwMbB8V
8g/NzTwn6iw0Qnlopb+rRvBpJsYLlWfKgZjU/De1WPnyfibHrvlAqJLEX5juuuBP//jC/syBpFUd
jL+dA8Y/u57tx1i9f6VlpuKtvuVRjde1xqxlkviwr3Xi94mLaBIdIr17jtyuV7AGeQjFWXNVdCJm
CEsKAh/QeDEs6q9FEwD4JlXsuaRjKPX8toYuSu1ARPEMycz6ocjzScOX0PFzTChurV1dp5UK8tYE
EIU2uHgoT8QMOru5Pn9zfg9cqJ5tRmjeMBSjI23Ml1VwkFpjt0WYX6KY9Z4GxDeEb4y4mvo/MkTz
D5qAc79TqFaXYhBWzW0t1tAsWgshP9PO0A1rzlZ3q41LF6FP53NWtmmAN00yXBUHIoz8NZsgBZme
YwfTS6Z80ddLqxpdqqoLlA7fJqI/nbBYRuCKWY3NpfLJjB4fETtdRs0gGNBsm0i0H0agxGZt47zO
8JWy0qoDQduMT0re5JjZDQz2lqp4bgQ2gJXpNOb1Xo5wDgh5vil1jnsep14JI0lNwRDacE+hlkGB
FJDAJMJgcneXLVEnG/Bsi/pWijh+D9ZHZLybrct9QLxxzNO4UORyXIpONloXjPmx7TJKOQ4PT3QR
WyZgBTkSAEBqznmlFlGO4NLrsq9aps9PdpB54hbzZjQPXAUKqQwiqvNj6sqXS4k6am1cxcYbRHs0
VVATXDp0BnJ23sEIMVvVVcP6/5KKztMm7tAjsZvHoInilN3FXljtnJeExUNIjxCz61wSxj85A7IC
EXzUMYkLM0es3BWcNTV3NOpIpPzSVeAwc77tK9UnnySgNol5mIg04G9mEDqt+GLV+8ZmaPlXFiHu
zAHLL6JEfFkjpDIpJGkSnZVoWojnSmH/J7z9BYaDyNvXeSYR2f/WegZRsJ73QBlgptFkz/5nujQK
Yse1DL8Rhrs5ggI0v4QsBdLUs3Zwn0rqnu1gGuSIAlhfItsMOXadWCsb0ZV7CCIaqIna33XMOY8g
GgOyVDJpe+bz6tvV/Tt9DiDkg3uVvKH0gboQQAhI1TBzyOFUnXw6J4jbXdrVJkiUtjlFjprECigy
i2oZvAu7hExa3fmVIlpsJfOwlYpnNMd8jz67Cr1a4x0i+wmT/XG+nuCXzgV5OgG/mcGEO9Y7Y9M0
QlOH8Y6+UEs9/p3bUutjfFGpWiwwU6YGwUgPOp1SRP0aBl22avaDJmyJ0SXDmr1DlZhqs1OmWz25
WKyMxWjrYCJiBLELJbLZgD3HR1LpJ+9thXm13VCZU1O8FGxwXAHC/XF/qw7cGO+/Xg7GvXRnLGpN
nR1iQjt3Lwdi0YFJAFKS/PK0U+Qz6OtYvm64Mm4xz4gJFKUk/yxiddkxCm1v5I9Z+SUeRaCdVN92
zwlSRlnuY3u2YZEBL7ScK1Ge0l8X8alUoHBIhTAYKtlOUB+MqqirAMvUXoKV11tov/q7ihMoYQod
frklBRzT7Fi0PSI+uJK4dwBMk1edXZDUTPBek2xALMYKkucUBZBSj8s6/IEavStWycG2kcYDMmNw
PoNB7KLsBH0H1po9gkmNTTIsqDdYWpv5JHeA8C/yxlaMZxIyc57n7rOMPFVxJ+ZsCh8NCHAqORGu
sEm5I/ByECOt/sBnjRXGtpouEljKnu3Pgkfq6QoCQGAoHJ3uhO7Hkay9YK/96pDbIhY/9BkwBcVW
0qsbyg1DoW9wdGhS22cBfc85EkdRDgwkS7qrHxhfWWq03HylHb6Pu+rizuA1vY2kRYLXxwgCI2TU
sfD4SmwGlc/s/tMUb+BdLVLBJcysVcPKaEHw0QTP7Hvu3JfxylRs4Y8C/sai5XYBDdxU0L8izVbT
9j2PcJSANiSrlU93IpU22Gns5WlVY4igwZKHXLNURagT0dxg4YlVC4v0BzrmtwmtR04IuCH2YJfK
P+RKTR7QjPckt08rZW1VAyRjM3gjdhnHUGED74HED4qYtBcJJastgHbyfP8zqwbw/4zI5I+qGrqP
e8/JUNAQoD5C02CpMlCez+nUrbJClEV2hwpskVrTuo2qBqv1umNKZfSZXZUbxcfK7ES9unUY9M3U
zsnK0uWBqxDxJrpxZRYmjD/59mhtUzU8XawrF5uU1ztTOHXnzoWc6DLy7UmdxpOXI2OdhtzA9poH
j4ANmMcsexYbT8CERG5MxyV9QakvQyhrg3UxDkPqJI442T9Mf3DWaT6JHw/iDqxS3gzrmKtM4X9v
bx1EGVrRXullcCtYe//GqmdLRM1TG1BwzBHaIF0XepUr7pufxGDzFS2EXKzgEZFshg8bwXr689iF
mILyAObvh5Jb5ERQWT1K/HuP2Gr1+o4OWZCsQAzRQuReFx2wiEKCfJ/bGTd9y2R6A4E+lkZauLzU
u0ZfXa5FPuqw4tiNzpT8tQw/rZxCfP4Yncisf0epDytCy2gaFY3NtGRkEZKYksrZjw1jbX3DToAV
SaZlix6ujINHkhHZfs1Lgisty/DsWNu01IwW/oBuK2K6BTscQqri96uPtIMU5wfG2M/19xZWkgir
QaQjrCeDPnL7IpZA7I9K6r4/1IYayXjIZTH3SderKnB3kx6I0fVUXE1eIJ4HLVgYuJmY0kdmWsW9
/voWFEK5YfGEZsFzsoJbO3ninSXODbnZwCegHJm/7lbVJQcsjQBo0Se748LvJJfuK+tdCB5a/Ml0
ZCorNqwlJgVuAvB7kuwWUeoahyHVs6T6RNZ9QNI0weU/+lktQBpslnESjmDk18s+YYeDrMr/nD7u
8ctm2CUKoG2r+/a/zgh1GC22UH71wh3VTqs6fFBj5ZOLZxLNjCBEhBaftvMDSgmP8cKZTaqlsL69
//zy4zmelzOrlzSXTrlFluI5+EMAXZlK/qkpjjrxfszAAl5HxFSwgA2y8YWRfb50sLvF5Yx+BJUD
z3pmWdGARSNV5J6JLn7oCFICudZEd1A7/IIsN8swaaLRsU7U1o1oikrqtFbmRPCR6oY0Lgh3sSc/
ai8f+izI/H1WAk800eHMJbqZlQ4vNBeA0MVCRKwyf1AmRFbzJZLwZZRjdVM3Vdq4I2GGi6nZb2S8
JCBxLjw75BbisdBoZg7SPNS+WgDFOJjQ2Qry60hEjrMcwrbu1kwAM2a5NAEDx6FCRAbjExhtrXjs
ZZMaI7en/qQwT/+x1UA2xn1HVjnPk96Fo+D++kGka07yzwkQumrVR6W9YLPA9cNmnYHedZP5qh72
M/KWGw1nJbKlVGFAaneoJZvl+I1rLjWgfJjQkEa4DceyCQztJvJFOBALtb5Oi/wtWS3tEG+5YQPU
0Q6Bc9elmcsmyJpLlBboKl5jha8OYonOBw+HKPvk2uYCEmOKwQZjkZg87Y4HZTu4XvSZNFxdNS2T
UH5cXD/TagSV2ZsVJV+FwYmmHOqW2zVQHJAyMm9zdl/KM599TDUBC+LUyyTXwF9nZ+5vsXUoqd9/
pbIubeUyVc0QV1wJJMu8E7d2lxtbQBg+rZMU82WCsDC+/jyszA7fsoS2B76U3oFKXmV61M1Jgj8O
VXrA1cxp88Q9rBH+S6kSCeG/LRiMBN5Bq2PzUvmRQI8DEwQ0ySlq8rPpDwm7rVckKUDarTO9TGPj
FIsLKwfPAhcZTA2bWS8oYXnpDnl0MokuEiKgyfg3QN0Hzi/biVukK05HewIomsJ2mDkUmtkdM/6c
i2x0/HpIbkO4GlkqNx9vnukcUGFqFZLp9LGL+KuKhqjx48Pp63whN2U9i9eZaP6sVO8cufkfPBos
pPh9I34k9WRfZ+gqBFNt2ZOe80EEMV9WL4FMMxYz1Cv5WQlfmD2ICoJATpiPdTD+XJaK8tpUIj8F
qod8U5ca1YiCUZremMJAf4fby1OWWdWZU64Fzm7JlhjNxBEHMyYG2yhIrq36j83nU71B7k4UjSe3
WdixjSEajbLlidiaV5gCO1IzICqnsFi27aBHYsxpVUm6bPI66xWOMJSKyUF9NxwZjXt5tebsFWX4
R9XVZYXbbG7ZI7hkNKu9yjNqTg6uNqpCCnABUD1KTdk0LF0Gq4xLIWEj+xGkX9Wcfy/u0+wh/pUy
k4d0yRcBFN4wN6ghNzBk45MfyhTfcxgAgCoWWPedZzg3EVKIGkQk/pSI97cFnX3zSAXdOprosSH7
WxtjuFs3wFOzJEhn8oQzHj02pUr8uGgsyWGmOQCR9H39gXsJoouzJ6bA/TuTTO4q+NFPNwt+IL9j
q5+egmp0H89tgJpjiPY1yOV3f/Tmh+z5vxMAfSfC61Eu026rhiDXKT/KSg28ED5CpCm6y02XjR0P
SYHF1WVy+Zdis0I0kPByRzJ/3loJ/bf0SFhZaZpQKgzLIcI5+ec9rE4+TlMMd+cj/AflwPT4zC7a
Qo5pEpmviKKW9auITUDhD4wXKC5Z8PZnu3iu/UKJ02K9anN+xInKlRoNMkqzARgo2fZbhoqKszBB
20Oglr/o1csxkWxgMaiAnC1ny+xE481faTRFbHvryu6/FyhmwoLQNwTD04cCeoCy24EkG5gJA5zb
70UmycmzU1YKA5Bcemjo1B5N4kwZzrKj8cVmzofGzjr8Ofm8U7lY64gLvI4xS3BXqcCc6FKeNw9A
LUXuBQth/UdwBVXaT1GyOojJz9n/P8wNlZB3ye+Qmgbm5pmtuq5hRy/2CiRGeCknnxm+JWPYtFrF
GkTQuy/5Pbu2fAFzkd6PJDYsshCm3Ij9xQztk/RkKgBHE1kTCz9tXQCsZuC7z+IBg8q/l8Nixs6Z
7VIEX7ZIlQ8HVwNRqhR3tSBVvnAKsg71je9p7w0XNHLiOpfGvKVPm9V7xuaux62i+ll6RLFA6XIH
dXt0Vl8Z7IkEPa4Nq7aEFGDe/Fxh+0NmhygHcYVw+VLs+hCcdQLONpAnasw3sFK2ZldrBPNhk34R
1zzRxE7djh/UeI9C6t9pTcmGQstcfpUMOEXG1o0cOFoKQp/7LwTPOK12GhLtOIlSnj/8N1fysQFy
AFOGjoan1BalXGFBQePO7GMIsC0ejLJUBndOBwwjxrCndvQkOI7Tm+j4fyoXbfKjk5hDRnW1eaQz
QrgEFkt3IR6CP1t/xyUMbqVdEETJAWUNDzQFOiEp0YhM3L8TWLKdugTpfHqzGtSqz2pvMifzFT3n
/7sukwambB8O5sxQJ2uq6MFzhrvZa2eOpCFRBAetDbXo+5Nff75VNO+GEJF1IOfOAUDCRGEovLN0
bAaeAFEa3NmIq/LzsMx6r6wBGsViZSkLVrd25ihPEhyyC5dhBHVGtImcY2oH4i3YujhPceDXLyOh
9XRnHd4j7HDsn19n7lyWw80zKCsk1L+dh8kNuBV8CRH0IIrJhVxqVK3vKOPCEIkzty5gOeL1juhm
/zuer5/h6vfYmLwyOIy9+dQTDGoOHZPDEWSX4GEI/hPuFJvlYe6D1YNoMoJtzpEfLCZyAdPaGbha
VUD7iKXGLXIkewIEx5a0iJERZMva73+G2cAeaNBk00SaSWCDksjigs+yJTnv/IR6DuAWlxtt5K3M
XLaWwsIrQb8zHYCSP8dteasjhiwYu+72IEpvBzXx8oQZ9jm7e12eDcNPqJ5plSPrG1oyfxN8d/mU
TH5jS27Fv644uszfL6brZxsfsxq0g8K4LFvJkuyunDEICs2Bzu2ZP7XCHFrWbkguHNg1HQPgAXoK
TvC8NyFgwisfmfY8IfAUwA6lG8BTgv7hxlZdLqbh5Weh1eXhUJ5FDfOT1ZG8LvQBZsh91kAkmuZ0
x8MzYNT5b/XdbeyhIVtkww8sxKBY4cFhN3Q+8m3WoCUjCoaSElOO6LKExROStj6uIVMLHM6RNsoX
6s4ztwERkUGg7RIq7wYe4GsoAWKaZSedt4WKEmGh/hcpTL19gExZ77W14l7xfyJoXK98yQfYVIgi
TOw6PNEZ0PhQ8bAggOzVcmMBq1fRRYXqJ4Xyp6wlCF2AAPd37gWYgV94E/pEm/mq87spwzjQws4J
P2dCfp87RVGZx1ckowcBlOIgxfgoYktpoFzqrrlqQA+ifjO4kF/55zZbQnNe/F3Ap8EhSKjxgKnR
2ffZDaXY9SffVfFgxjld48unfEYLfX8MxvV82P+uTsCWZn1zJquz7Q+Qb2Fk3Vl/aZTFPBKC9rFI
EtNOOCMKep1xLfUOUbWvsKCW3zgo40W2BorlTvMICrmUPSPbA0eLEP1VCNAKN5/HQ3ursewZGzq2
qw1daJsGf7H235Mm9y+QzeSv45evvy1HpXwk0gkDAYfAWZJaXeKuitL0Pph+SpdGf99usVdbJEZY
dDdpW2CvnG8BQzt8It5yOq8i2T18adNDg5+d6052Ec8XxloG2L5PwoIo3ZOfaI5mDiTrdXn/HyQo
81UG8mvG8LxfP8WobPcgLUfSA/fpkUJPMsFnSzoI6uKDfW0fWEBLdQVT5kgEeA9gqC/+K39AQOgw
dUCa2T+vzRFeHXWtaK87fLfRgWwOlcXZLe5co8BY3VhLIKSj8hbPkU5ONU4t+4zkCeLPDM6EZWeX
MgutMn7CJp8Hb79VYjYtuHcEGI554u90uLXcr9uBOqCF49OmB0d9SAZCeto1kO0E3PpZjS/rO8Gy
T9if0mHr4fcpyQopaMVn4mK9THo4E6IcXMvLMYylWDY0tJY51ASJWhqnht1xpmAr/Z8CxzPeifS+
dOFl4q1FodPlS147870FElpnJtfTvfQ8kK13zihY8gbI/efPUtDImmiw1Ex88MVx2CGKpO6RVqvE
NcfHJZiDrgk9Z+ot6hvoKj5jpWXjBKJJ8Mo/edy5Mx4wGiWY1eti2UlzEK7fCFhrl1w44OZEBV+2
HCGZHCv9U0GsOfpVgRsU5JdCmyU62nfWb+WC58X/ceIopraWnjvW/UuaTntpTc53xvclIUU2VqUU
+4WxB4AZ+wlTBIWzc/ZVXKWOrZK1eQ+wpt/St/ym8iNNMG7lZmKUIHaSaz/4gOlJ6+YB1WAWKMxP
xsLYkTQ1K2jEpb6d4WOcZCSGe65RhxsW0U+fq3kxYmm4ZsbJdNtKyUXfHYH9Npg4WDbVEEMh2Kbo
CyZF+7cNgiTPwipuSN58FXzdW40UC3GU324ewe8qbZMduJGbhqFZExtiv4nPOrfwjdNQxdxyCfk0
zXL1CUICiKj+AOiHhiezWNd43E2Z5yxJpFl8YE8AoNA0W6eDpfXf0fD0Qaxn/8GS0cn2zNIQWuAI
IM546/M8SbdiCfq1EHPKHvULkEo6vOhpZM7IAZ7HsnUiIC222ZbLTiCxcw05IrzjU+IM3V4JyKtP
s6LwawONcmruz9GU2djviNfbIw4VYXIw55diV9SmrBFQuXv47ylk1mgWErDicBy5V5VZH6J/+x/R
ugUbJdlie9DdLJFWU5yTsE0CuqKhEMEw48Lmi186pzdMSXbRPwOdPCDKDW5rcLRJLDD37SauKj5G
9lwSStfZ4AN5+i4RyQ0Zy4JgOMjcYsxBfj7czB47dMjOZEPVYRovp2XUVNBSHtPBD8emJ+JOMHcj
pRLE6F/NtjYLjqdRANIIqNFa0mLIC5JLqS7R7JNcjZywPNk7nf01daB5+c3nSbZsvN9No94SZnlU
P/aUjDIhyQUjoXC+SGCjLwY+AmjwdtsKwYFXzV4bRrD1OBQNqwkNt++OFs2w2/L+LKsTHzULNcRV
uQV8sGv4At1qjEqPSFBEFP3SsUNCPZ5UbMl7OJZtFzRsdTLNzxc/TvXpev+ar/68cw6CEhqWF8jp
hVmc0DorCY9egRAggIJHBO5LeSitWmD8Nplz/OXdlnhO+OUWKSerhTM8qvAJPZDaFhE1Eit+cFtH
B/QFibwC1DuU9FONZilgrPV4kSotkAxLPubUQQhy/FUXiYQEikIJY88IbbEk9wwGbK1t10so2UfA
WA6N5Jax36y3J8VU56tUqVzJMLmwUk6U4D348SxYMO0Iwflk/jKLX+EhyyQg4pZsb2eQKii0oY8V
q5ZObu/9yWa3ep8L1I4UJPwAZcLDeqobDFIrqCDozjKHerKR+1PPzKFm2Z0yQOqCBvicSNzjNl3Y
mUjAgVtwEqaozq1SO5iB6xNrvheajQLlOmYT4XLkyc/ucT1dJ476tL8d43Zpa1MzR3sRlhlLQaXZ
oZSEPZ+ZVMVJvp5KpqJfg6Rlv1lakSR2jaea+oMW6/g5GZlB2xNXzzaoNXXOYniv7Cg5ClxD7rxG
aG/6G1sq/BBsyRC7xIUUol6LJib+UUaKP2FzBPszC0LvXqMyGvG7INEP2wUcKK9tfkjQADiNH59M
alRf9oRdsYBMNGXuXX+7pf3fK1JpTD+PyAHxkuKdqLZF8aXl7a/zdqC6OoE1sD3KYAL0mUhby8Cj
3BrnbA4rDybGUvjfKm7BfDrEmg6mI24uQpwpzSOYwN7tzToTmjY/13b68H9XZPR0+nBgjBWNkQZ5
Cl4xyuBvmGH6c8ugSzCQ7UPjCcJikupbf2dLn6T/r3G4fkDBCgOYoX9GSosXxKPRkLghObE/Qcq/
ex/eKE3XernHaauf3yCDD767/hNINF+Ltz6ycTbZZzvkpwhpoa1sXGbRrgltZCTS3hZ0OQyVeJ6r
G0SpiVYqiyrVLuXnHORyXWE+SLbMvxUSW8EPvrjLGZfFSc3SHlSBb+gipp+6mVZ/qKNt1xlvkeyb
FuV6BEa7Sz5LkbqzSQO+QBj05yncLnY04JNpXF/YPOoysPAIlgiRVDDfovqvMknOFqHsMCpn46sV
TsNEwFVAHea2a0huPP2rfxtIn/4gc9UuUxN+KctEQfNVuGs76LeYpePbkwQfrfedlsNL7NQO783i
OZq4N2toe++IOo3i8xW2iuBSXQw9wbodkKjfIf7XOKDiJAHgFRT6AQqFOPU8+iYZF8l8DkzQKGoi
WQS7L27md+R/ooSQDB1KHAFEnM3+F6TqxpteTCcirZrWVD7HOkDehWyChCOFbVqKDh7VpOs4ggiN
TbL/n58sBAzAkbkosgQFHw6CCZ9VUGwYVUalxhoaimDDnD/qeeq5e4igvzsQ8SWJRk96iaC5nHCN
CD4YN0c9ffhnuOoyZYSzcNwOVBMGBLZ09aaP8fw7zPY76RdjtTNyYj5euL9idzsr2YDjp7ECCUGW
EL5USqhhhSdmKJnxsI3yqOyDDRYClYV50vyZN1yDgo2RC5KrXx61AaaZ2h3i3FX6E0YlUWbqhY2O
gOn4d2awOLNubxoPWij8XZJFkxcCntH+32fBcgqCZ9VUqxV5/txT4QTE+oaJ7UCiifMGqfuf8iEk
4rA/V85I0Ablqs9iusmNDtmZXl6JFzOO6jiiPVUHJoSmcM/4uLdrcT3ichDs0Zks5qQUfHiBzukm
pr693/0pLX1ty0DyQnO8rmnlOh6yQaOTLhItr8uIPeZa3z+qFkmaufS6Kd+jXh9hXAFfnzwKuwu6
jmCXBqhPZpkZewgU9lkBe51Ou5WCttmrPVIS7pWleKLsO5cul37VpOR1YysUEuPG1OVyEUZjtsNj
I7dhlFRFdJxLi7ZDw1FxjlvmRiNWbX5H1THbic3wIbtoX4dWFBWOk7EIjfLyKL78HRSJ5+v1dqON
7cBcE8WX7jX1zVzXHRcYmpQLL1SDEPibYGT6hCnSxpJOJeW8vXgBEB/w6+m7JZvO9F/JL0wdsR8X
dTGzu6J9v4zAXsLQe5TUfwamrwYAmDiSErGS2bbbhH6xZotILc1sHyZ27Xj6yEYwpH97R2QDIVTL
hnPL676VJaaddiiCCG1GxaokOXtrhbIcN4/IeNZeEovgdRei+O9zHbYe4bvtGCTjEi84HIaQa+lP
xfTZpGUSHvsY9eINzRTTue15rxRsJJUCLEm7LzkYK5jGqzRcEzclTj/tN4apCXyKdY7mF+wFVoOL
UKPnt5YtgSS/9LXxgTqX0Dzch3TmcAQD+9ZgmdG4tye5HDGYjLAe3MKanzeSHmrOXimV2Q04SNlq
3XcFS45LNmwmJvGMyZnfIYU1cZckeuui6pgbYS9/Ap/bIC4+Tum8cc9M7W3/G3YEvBsCMujgP4yp
5MCaSI85T10sgMgCLPhFVb3rO/DovzRTBvbNvVIF6JHqsNgVPQwm+ZKR74zStg3c6kLxbtostuS5
Q2S52sdcE1RcbSkcledxAue6erWTpgJo19AfN+P+gJ2WFRtCUVmjSWifZvwrvYar5iGp6/3Mqbw6
Ba09HXNr9FfsVXg5o+EktjfW7X7su1zT7sJhqTY/9XdQM9l6Y+xL5RwvnnZArYABZKW37DjFFzZP
j3bAIoEtU2nVjaI3bDAdrre8DLfsZuopebqAn69reLMkcy/KnLVHPJsmpiLY+g379FQJCEqqQzoW
3DaDf3qCYoG462Tm4DBVRBkPqja/zhyv5x8HiaoctLOmHoZqlTLB92QSFiSNv99UqpzW1U/WG1I8
tdkt85uBoeP1vRYgsU7+bka6Qp5aM1Vy7r9KpsDo1o4ivS6zoW6j7aAtWw2J3kM7c8S9hUwhhrXs
R+k5EQI59QljxEeDGxroF8Sqs3Nf4OsdtSI3z7AI/NK5b9RthNROIjjfSNF58undpm/t10VcrLGB
GfQK3c/Q1KkwN/j2udC6bvV2lYSaquEyUf44EYICt+iqr8L7t+3FA3R8CSmON062dPca45Az54eW
gVf8PcydVhOTmZBTtXfrlIouu4DnzY0uFXdXbixHn/iC5QHHzNn+sRLOon6F58L1ZHIRgMexSWBu
i8TleQnYIp8Lr8Q4ES05YJ2eAOGRMZXQq2W6E9H7KDq1Czt/3SC0wUvKjF2UYAnJegj9Zocc4cts
G34g8zz/n/O7G0nILtSkCugT6gXEsmgwtRlclN/WJU11UWRR+nbiXd7Y0fk+Sx7uwbVO2jPqcgQi
/kIpkwz+C7c0XKaFe9oNuXGqzhFF0fkKWKJSGxwvECQuPrvUwHOjCbEPjBntw4JBT1Oj3HAbvhgm
y4MzGyc7S1QbmfFfZ7uLkL4MaCU4IBH1MaePJywS2fiUQa+vJ9WLkPAWksBVHzltQeDHtA1wTsND
m3k3sxQ+cQRrZGpErSOwxfWyVTjbFSd0AawqBeqeVEG8XsceGnAbE22yAgxAcb7WZs1W3waHy7RN
RVmA6GIbQMf2xYdCsXy+83wviTeKuJtL/g++kKbAQRT8JPgqPNZ9mhUpapB9URXlJqBZdWq4r4Af
3DKlta81XBZd3Zi9wLjFHsJD31jnPRnDY4GKO5CMN3qB0VkMnYwz21ZVMZV7p7LibTKEpW5MuyXD
DCxhx4BQNeCYFE2Fds1hfXgg6bRAQZCYg7fn/A4UZnRpgUxYeJFgLL1DxwR53OQb/E01TW6gDqV0
k1ZX0JtUxFzCuX9R8jhohdccHzTw0ly2PgZyuewpXiJndaMtn+2uj8uaVR6PA00sb6O+Z6pnrihp
hQ8/2FwBGNMgASQ80cvA4eqzYaJTf4USBjy1+S1SDlXJsJErsjMgWfht1sTOsivjgYRJQ9vYjY3y
nRwvf+rlKy9MfMVMh+cif0eTPXwtgXZNtlskUhkCt40AwL3tx7Ic8zrMsNwRIyeYvix/9yKqYcTI
uVTWOVtQVzrAYSMBbyRMfp6X9fC4vMY9oOX1lDdip3Ibpak1VInqQu+mdFJKQpVdJn2qUfBjXj7d
HJnib+8PMuvJKxXduzkKnsm1/bkQ8sdOsfH09lg7IU7zMBIoUikRDIVV8wI9PvmwgJCRfIG0kKfs
GvtaM/1m9utbySEtwZIFa+N9mTqJMHpdpnYo5v4MqgTQ44bF6WCqyk9HBgDmlFBCDDDQPnL1INuA
JkmbkelUC0y68Ugcsswgv+5NyauYrGCCx6S+Qjwg1ra4iqc8erXRwvojaDXowMVqwARfP+mzUPxx
Xxzitv2iPX5BYdY74s2rCE94Ecsx3UC1T1bzJRLICZpb+hcGjeY3hNfB6Lrtcjlco6WG0rmC9nzr
HPpymw+c3aN/hwcj+oWVMro7WqAUdLTiR1m1INMV8ogWGgKolrC+AOUUmUKTbLE6MDjgEXtN2gtD
9PaPa8xZQgWirkPazJQrVVgfQbJslMFuT7dLmGdEL9HOIE3vqsu5JwsuIqses0b2PpPeTt1EcJoQ
qNNk7nmn7XHDT+lbYGPt5WtM3E57KttjF8hxTRWb++eFy901Atut8+fc+hhA3fjpOaCLIe9OdVPf
2CHMr1M4BxOISqtV6Tk3kcKfrEoFEzWZ1XanQdl1lMeyg+GzuCFxTnSg3uSo8BjaEcvDp32pFrQQ
9CBwFyXHre88jsTRhNA1Ju9j2zPMADVL/cSVMN/rRndboOHkHOVsAw9HRpU3B8No60MHP/QK2qVi
J+CfT+k9uqAfxJvQjtULkR+mR3wg2PnPcp6vSq9Br+U+W1Z+q7rXHdkEAMQZKWoqn+MbK5OajFVv
aL526iqjCESfTbLy4daFUsKI/mMMx2+4E8fmnzliHaI9JY2sDeXqyCoJDD6oeJqbcqmKDB7XGEsJ
E61QuBnKdiec7sAQiR/deYV72PWWZTV5KbtRji1hrrLKhUejO7KHHwstFQC1KNx9b2NW5z3qEWiw
Mqd98wpeJ/svK3ITcjsrMCA7w/KE+pRNlKJBsP80heuHNtjcqACZarTHWhdOuynDA/GGEtmZ+M9D
xu4fMaTssMvROpXCS4bTPi+H7AFY/WJvctkvl0i80MKayuEkVzsWyShVNAmLwjOYDh+NXqc5WCKC
mCySfl4v7dsCBp9yYbRh1WzxNOjLVXzNYcbqomr7x97G38NBggtuGOgjDLsvklALtAWO0CKSvbns
AjXo2aD0m2f8HFA9V9dsI5LufPUcxNqBR1t19nvGBC/Q2Bys8h4mH76SSi/4tl/bvuh6Wmd8sBGS
d83J+8s3tnSe/haJma9yDCQluq4ib6/Rt/58hVJ0M9/uUxkOAscjXKnYAbRHvBlGV4juu0XwAA8l
2wZeJR8M6YlPAuTHUzwqacxQCGfQoYQ3PYtAZ7LGjIHr8mLDwWzKtqxncLYCyDi8rhFnek7EfVfO
VIZNHSwZIbLzMzkTLOiEwzAAY/GcHwjqnIS0cTjzPSFJQRp07JFuk/CuUMoOQkqF5wKqbNAeaSJd
cxNG0uCfkEU3j3vssLlY2DvjkVQDNV+ETmx/ZKYJtkw5yO8H+xbSBZFttMvO+w90wnjOg4Yzwf9r
VTZoGmn/pkosZGwAHmRZdfXWL7FrKSfQQZyIWxVTMHahsl+0QcvPy+XsmGcnjs4z9SXzodFk03GW
VROtYeEbbN/djpGWI+FmAK6lQr3c2D3T6d8CUXuHzCguXcA6bzfKeawahpot8UCavwKSL6RkkwL1
xi8S7RpqRQbWAgGH4r2DXrH89SsboJlxyEPP8Cjff+ib15d5KPNRH4x07YN9abQkmiTo7j1tSq7Q
S9xnxPQ7yGbcOnOR2QRBIlkcDXhKtH0veWRU/xcifYk1oebT4pxdhP77dXjezHoD2nlAiR8fosOi
Fby/8MJfrM4MDp2Iazw1LaST7ZpvcO9rqdEMJdnfu3tGSZIFh3hgmrCZ2Z3cNoe5kb8D6eisPI4G
PnpR/AG/z6rPLfmfc2FZ7yKqf3G7dxqFPvE9Iqeel+vxTVPBmHUH2jOSL0DpehjN0V9SlLMwT9z4
a56uWI9MeiQSLrThiv76qqqZ7TjRUXWvtm8XPEQQW0FxEiDiy8Xz8BP0tMo5PLOrOXyaGsNrKpfZ
kTQw0Si8qdA+cd+5Q4AcXnCdzrErMJAI+0c8XDp2EIYXTJ5i9jB099TO3548qCP4qZpYHvKj8Y2d
IS3IPS82tsaFRgco4/3msRG/oyoZNQLWTyJLb+Zz/VsT7IAZqNxlSs8JhMrCw9nCvP+Wp5kjdA40
CxV7Tf5yAheKrgN1qWYFZAm8LxV8Kb5LvE7Eng1PZOoOgZQ59wQHvkKvVNB9mQ/i7EfWUD/4hQ4a
MPoUERtrSH/n4mGiaX5P3wB+o1Vr9sHgG2/VI5J1eCSpG5z1/at5tANshCdal7y08IT6+kqfBqG0
XpLKEwv4sy761o0zjKVNwppMI12vBvYKEMfUOmgcCGT4tQ4y3J5AeBPr8q1rZDuyANS5uyTpyEQq
Z8wPycZzFPwyAF/K9xq5cQZo9hY3OwIDNNXRDge56uPclMumbugzv1mqWOs7igDpc1J4J1/N5aiP
p59p+rVPx0dD0JnGr0mSo/ne5kmyjsySRl4Ig2vQo7LP/Aai4xHtI/F6JIR7fYXsTKf9OQoRGH45
StVc+JcjaUKfz92dMhvYU5JrwtidEtutYJcKLa/qxVOBdlhbo15/OWCgpSNWIQVZwHTXVxZtO6Bn
KUP9KrDt7ennbj0So/62aLVOWq8wwh1DpVG8LP+Ebg1DEN9qzq6KLarah96z2gh8+C2fiTLI4SaW
1WUXW715CGbt50dHem68HpCw3NCS2T8KYGPOjDE8HiwcJZa9RR0RpvK27TnMhDxgag4DW4wb+WR1
aV7feb0KbBBXMuZav0BirmThACEe6otcNo749WN8WvCjV14api6eKmg4uYPYN65zOf6BGK2dgaRO
L7QaTjj/8EetaBYpRKQb1SKT/VLAvH3aur+Hs4DYFel08gqNRF9lqo1Tvmvg/l2NGIXd25em8G1j
kOO1FRLT0rg2Ut817+e9bf/5yK9iMm2rO+jiS323lgwpKHCPGm5gOyfQI5SuySL/dkl2kWvaAQoR
FicNgN+/WOOzR0afs1NAiHwNEEhvjOx5Uq1Gn4a1JDO1xqTQ8ppfj/GqdAQuWlXbzMjfqVckPJ8W
O//NMqDPCavyCYROS7bdbT2pFJR4erp+p5uBD/O5HGsR3/x1tBpEizt53BEsfZ6eV4B/y71rDu4m
2nw9l4w8+kB7mZMacRib05mXv+DH240n/Q3cDiom1HzVcKzaDztrVcH24v11bUA7tSSCYnAs11ig
fvj2XOugn9yTKe4OWLNiTNpj+Enu0zMSmHdBxIys2Qw0Hw5eRRbwYZ/NAUOslAMiMvnTQlrDaHDo
81I+m6yURd5/vuBZ8sQAvmLr7UOM18x52xWaTYUffOiiaUpqEng/pTwrGwDjJGgHCUmRzBj1hYGb
EYPAS77VuuFf3KQ+larRjgyvSnVb6DrLNjg8FQ4aZPiGMmD1+vhtNxYv6Ypj8qo3/mv+GUOlGbmf
Ru+n+nwOb4aKMsSZJ6LkwfMYobQxjeNpq2JdXghXf5NZgQATLpp4hs3hDUAm4Wl7FusqniFkdch+
fFR6KVjV2ODxc90uXqUhVvaPMOQqxyBbscc1J1x9TnTnlZL0iJbEkM/LB2pDp2ooGasWL7jtpwz8
MZBZjfjzdUn+wtEkSoGETSqS9UtTiMg2tiHniSSeIJxaWHhFCa9WzynWOBaHJhw8+PqvJaR5QY3q
Y9mG44ZlU1fpXoQKdd6+5LVTtaGjVu620Mdzi1FWRxt2ArQRLKePamgGdWi2R1V7HL9AxnvWbxpC
fb/VyGg0AqoAwGrslqUFM7fUfBSa/LtE//RFnrOMA0JSRE8ItrEyrxEALQ8rtsmhs3QaNriZVuVG
mB+b9LouXRdGe6Y+xzF7i/7OLe4KTp/kBf1EXJJDB3f0Dcomrcxq91bvpoT3SGkt95qrU4YrFfOd
6i9mrgH6ZPPlaNrRsgXot7yCl2chSTfHhFJzqtzTMRZbspY7r2Gj4cIDy6lF2bcm6touSudbyXJH
CW7iBeLtxxBkaFqcfNZlOoS6jpP4S5qmyVqML6c8RuJPfTKiYgrb5PTfausLBUjBHby+X1Juv4Hl
SvkidI1m2YjAoMCfOzrmGBTnQnMLeP0sp7kAvDD1/0vGyVNuRPx0L6QcmHUuFhf7dF9L6cfUq8Mo
EpTKTQ5qL2To19qHgQrTCqMVOZmXs/eAJyJnygSidIURZuLLXD50XRF/KY/e5RkGZ+0Oviz+Bejf
At2hbubw2tz+LCALtB8mxEiZSGnTGMkCzbzQAK7cDbVrVZZZVHPbBj9LYdUeP1rRfiahPm6eeb4L
FOfHyNnzlGR0j9z0HDol4tczblHjdjGpR9CvWPGPeD3Vf+EHtSLFrZjXNvurJK3YwiFJLQBE0jA+
iweghpP4M2yBpmxmDfE1PnfueHY3VybwYaE3RdMACP+3NmohV9uN5/YtmpP9+cBP9S+pIrtUJqXi
/3tG5BbM4Wbj6w8x/v/nDnlVuK06Oltj+D4Bi+bFGwEjfky/A6rRuLAgBAUIHhqebAA2IZiPhd36
BGJrZutJ009cR1Jd/Bd1LmWIw4NHGm9phzXrs1W2wgucWcja0Q5mzUIWbidQ9GNIGNLd723e7RVc
Tr3KKSMBvissU3vDlNKsnw5nMZejDzPU3v5tH6sbsSh3IXgTfvKQuCPvZr5B02YKMVDLxFgwxvWI
kvQbDOXmctS9bNj1H3jF4kxDg+MD+VTdCvP91YU9nZMzh4cMzA39CcRe5HO+WI4K56sGfHyZ6MuL
+gornSzKh1/NoKpFL8b85Cst32qAFNhTAFJDh/vm8Cq4uZurRMeVTc/A4ERCzf9+RQQlSvuOuvSE
2/VtOqfgnYui7H8w7HJpkzuDNEHsE43AvVp0gK6CjOUGS5JxFvtOEhsnwwl7L2RjbobJMw61fSKx
8NMmjVm7xgeaYJMg0lJ6/K4CSgYWauJq6rUwlkksKI/44k7Lo6WdiaBn+yGT8AG7rz1sj7glk8tI
+ttx11q9StdgNl3WONW51A8SEqZWsYnYeY4pxQZSp8Sk08QqQMjbcLXWlJB60F+5iuYB+JRW0A1j
b/CiZSYy0sfxBTLSJXmhj6GNIHlXbhRoCzGQDdlgyFv3zeue+bvtDfDHKjP2oLg7N3LNmVKXanJO
xHzKdXC5MmyXQGKEQ+As1aruRJLqsW4EzIeY1JdzVxfQCvByzhmcUZBJnNr0uxuLQonViXkW4gIV
gylQspN+50Ep9E+GFXStabX6EIc02AdoBHWKwL8J2OtAkKphFQlSKO3SWFFP+BDXM2otF6oKGJaV
6CPceQsGUXvXIzghl3FiGJ1qVUAT1ljBB3Bo/6R/bqEVnX0Fv2+e5dSM8KXqmBez3G44KDl/liCk
ro+ZbsH0+opJIzaHcT1IxfZozRuHybrNDB6ofoLfHpITurCE9aNntG1qe1N/UyqA1IAV1wn6O2b9
ZehnC/wgcQl9/roId7fZs8rlENc9d8bPw84j4psJkkGTQHzSSg3pyVHE5QRO7qAgRLAv1WKofxgr
mr9d/JVkWnLyy+tmqA6+kluHFkiuyGc3ZxjRAce5fVqgajdtnAAfZ6T4Zr6n3/TWNRgQtAKVPkRL
/tLxubE9ead/fwpGe5tEzYAVQfZnWfz/1gtdG8I6f+TWpn3/bozjpNhEtYUG7+26F0PyVSizkSgZ
jVgA+sj0urlNy6OaJzGFQCiuX5h4iO3YWoPRxiKyFY7M44Ovp1ZACuMaStErDMbZBSCKFjcA4NQl
hDtz48Tyli6ftiKpXbL+9illzRK05noAAiS04Q+2jPSgwpraNExUwbnpux1Yld4AxvSzJpy4e8gX
w20I7dSh6LgxmPj3v9atocfNvABG04QVW2G7AVpUKPGtQ0kqoB/FnQAaNf/2fOVdb4S0tmZjTbXF
K9BTKY+tbUGlUx2PR9Yr/b5IRFDxP7mTd+GYwTZDyYBUUWao5FaHdlTD6k3llgwZrvbA/9JAV63A
4xQus1UNiNk1g+rfAb+SufwdK6yl1LWA7UoRegfExJ0PAZnLUJJPA948NFrffJZCdRuUh972PyNj
76ZS0bElebO6lN+rGQjXUTgzzb572GqkWzdUjFxtNJNMtmocdB+vW3nENWLTFRq/sIsPvyYwG+/z
HyqDrR5++fVboc7jzh207TEVSW2NKpM/i4/ipxfjcRKPeIcDSiJfcce+OiCMYBRLVegu0AT/Z0Hv
RXmOO1cjkLfKLfK6K19Ht9pn0DxQOhdew1MCgmKOhYi6q7UOgfWtO/DUKSTXzsOPR9eK/oKiDn1h
OOydwoo/JzFe4XrPN9+E6THH25FXGIVnEWxa4Vm5awu23sfQZnbrnIH3kLBrLOyS3VNT4rytuNBS
HRNbVvCvPSHs8pYOSjQt0in9EWmAtoFJ4NIzd1Y5o1wiikDjdRRJrmeu/KYREJugvgZACymD+l0T
7wcrTlyFVJJuWzXFfylmgq5aHcyyZL8mMtAbs7KxmElnyTxOP8qSV4sgG6pgY8iuSCWxzKnHd1v6
nkrsUKzHQ013KH8g4l7b/+dQSxQTHzu6twl1yzO25x5e926GnSsmcv+x2DMztRlxlkIo7rUG1Ab/
UzYmoYIEmcRJ1LJ7VCBm0nxc1RQBy6ce56jETnxNMiLLH4L2YFwjC3QH97Y2osIcNQZ8sCw5cj6I
6nbDbBZH90DgaU4n2s0EaOYmq8uw0H3x7RfMZKxwese5hm0I/Sxi8uVqx4dKiiEVZry6UqFjmV/Z
xHti5xPcvlb+Wj7ob7V0dQ0xJ5bnpLtIl7b+Lo19/3JO2XNzcWV8K7Dwsv8fbUdMpzJNMTOA8Xzt
b7LessntXfGlbPoF7B9cegNyxnrogF/KSxfDXY2X5bLEx+Vl+BAKp1RJaKFYzmt49obYwLoRRD1m
NwZo970Kj8+/0d7r1SJT4KhykU+VG0mP0Gtqaxd4KdnUM0bYE0Umh0dsAmym5weJvVLZaFkGJR/+
oFDL1HjyuoG0sl5F1VjjS9ZHZypNrFCkIDGhIM9xIq4+jtG7bPJNFQfDnPEg3gWORyhkMmdV7U52
lRFOZpX1ASa4fcLTRjwJM9l+zBgtSg4pnDG1E/BSbdBQJmCVLbPgUun+qDtLp+Ok6MF3mppy9L5a
29eGwIXLRX8zEomSXS5/4vDUHssKEXPO9uc0Nr9cjS4t7g/eGmdjgLq+F/TZN05f+aKl6sKiPM+w
a6YEH3KHVquUS3TY9i14bcASggF2zNAWdKZsfQudyB7sPNktegp0bDS8oX+J7EkPhuT4EBdeRKUm
JyGTVLAaFjp8MC3m/OYzhD/WVZMQaBplSN1V5ULPGmsfhutzhO/1jYNzEZxPqOVqjapi9Y13fBb/
FVObU8QyXqJBStm2ejUw/1yTV/4u6STgy3odPd2zg2JnhRoykQdVSOCOA1jLHlCV5mRpbT5EpGjR
T42kHzrmKfOh3BrpTrkpwdG1e0PztOCbccZc2srJPWzpDRZpQcf5ucfIMLhcLGBVs7LAUsroR1CA
4YS5OkHho9Cz8lTRm3CYxwywAPUTW9iMiFQLfI62wjPvRQA/HX+me2gh1kHjNUAzhyr5Mkygw5Ua
KVrLEhnN2c1tLZ6quCorrOLXAisucSgOolNPUSTEec+K+/cC1qlF0A0dcGXGd/Hej650smdrD7Nb
+MaY2uVy32TCvp3z+2re4j6J9KKVB/e374KRaRXJe8+Y0/QIu6H0UOtZysZgOer0nBFTDS7Hfa3a
DQfp+BIsiuiJVJ6/j1kHPI8Dj2rvDoZUYC16D8OHtHmXbltBYmBbAwTWpA1OIsnSnP5+Lea2shYW
QaZtg2QX5/hEscIRWejG40i/43MlXq9YAOJs5ZO53yGaWp6pHVdPb7oaWNb+LptX2PMPk4t5d0aA
Ws3s0SiADACCjYeX5Xa9AjAjzmnkGLX8DoAdbv4fW970qhD3wAnHybr0nWPYQR5ehJxE4iYfRGrZ
c5gEj/mtiXFqFwjdPoisIwq/W0cI+wemqpY3PIz0AHlAYS7XTF6DhLTu1vzOHBdKUbz4pLz1TYSi
b5Zz3DHYKonoVdlElE8wXpWxPqCnqPGZaZxnoXsS7jRfcfIhOdUGuboSwzDzPrxyHO1LxoAAtrQK
5NUEQIn+njQApMSn91qsCq0E7S617pA/kTWRHNzMzH6WwOXRZs2MpQUNNoxvVqnK9vff3x09Hefa
DaywIf5WRJfndEOMiOjzqZikgoqKlLbc/uxT1UB66c4j5uAde0ktiNmjhvwQoGKeaiGY3f2Lq1N+
dawG0Asb39EdGayBEhyLBZFxqj51q1qQHeww/RJv58o53RlanyWYcAAMR2d93JnvXnwO4XQgAzOz
aGH/td7AQyb/H7T5MpJqLnAqmE33uRmM29Mw8S/pHBhQiW+wqbaeVNd9ZmcFTAzFxM4Rh//6/Q82
EM3pR5xd6QQ12Xqb0wZc1xyjRQwOv6DYE80rahZdzE2DLRE6YGw8PcSD3f6DaKDaqc36KnZxL1BL
vJ39WWEp0b55cLZutQCQRHdNogGYlOSMmeqGCmKFlUHa2eGaZ4xHPYZVja1cVm9bEVcx8sfjN861
HfZYYjF+Lh+Q+64ybG4MvnM7QRSCIa3Bm7UZX6wsLGcO93rmKfng9H6LgAqcSFVc2NBxkEkds/3m
lPyy6h3CQ7VvI1cZk/7l0P3Y49JFx5+CUzmsQlERXCcB2OEI+0AQ3Lwj9csXiWL1Mz36xTnI0x9B
7yQtifn+qsWDkxn/rb0pfXw0Nh9H8AAebE84wLoILg4w3A+TDH5QxHrWFKdR2Ervo3VjRDCMR5nV
MoKwyw1HlwAqnqSMHhmL2/vr/kcJbBBd7v9jakjwXsguFAtKRUJc8TJBdOP3qLjove7nh51hEuRG
dFWL36U/itPEy9Tb0dtyEZJQO25mzphysXT9wTXWsVmUJyH6Ld3LW+lmwbGgHkUCiLgpONcmrNUc
6WeLo1H17nNptMGK0lF2rwZJYLISRIBTqA5qNj8q9oAlug0onG111BrhRMjO26MNUUzTHwESkqY7
05MXI5TosHAlxiRURz5E6VlrTxsYW2qq9UWmeja7AmlvPsrbM8W/AMRkTrtkWzu9sRur/KDeTJ0W
crKkTqaQ6UhMQLK4J7ZYWF0dObBtgGUbG/9BwWKkSv3qrDfvIAeHG8LE/h+88zehCSFf7bUMpby4
2B6ICOxwOB6/hukEPCnOH88n6JBEsG+V3Cmgwpuqf4r+P+msvkMrDQobZtFH6L6DeM87C4cNZ0Q/
H1KjJ+k+MSFHWSARabLzh3dm94yxLtuLfjTba1TM/mfJ5jACdzzBrxXGSxX0hIMLsMJnKNm9wiAw
0UdvU+3yZdPLijyl32EwuKSwcNb7vhlsSObwNsOk5seyj2yxUgi953B/3Dx9/Oism+kLGwrNP/bA
O6BEoD8X1ms+Inbq9ycv2WlVLjy4btnlF1v3A4SZfvQEEmANd938rwm0KetTN+c/GoQjFVM0dcCx
4OHrzcNRQo0DubF5dELQ69n0xwa8eJu7wRhGuCSL4tva2j5g26z1olCrsV9XYm/gP/BGMefbWoSF
FAzsMPWP0NiaTXhE8SPPeuZbXV0Zc49WEqC2iMQALwb90+9KR30GdDxo85EJKhIH4K6b38Wn6ZMh
LrLB04ShQTuknSjVhYQiurVy9hOjix3sX9/N3WgO2gEFnGGSJPpuI8REsl6Jt0DrIzlhZ3FkVTp8
yzmjvJsh8xcggvV5mu4rjFH06pglNJRE2LTGuupMk9L5YTugcvF8cYoa/YS07oCSl23ZIHolllv+
RoidMrwpgqNNACZz126WCVw0+n+j3M5J2wbFdZ++bh9b9fGhRViLs+AWa6pr8qiqoF7/nNkPDXnb
ZIgZHzhcjK+Tqh3D8lxVNz1lHnMdi2UF4n0dyPNi95BjIEd7L57BuokW3foKGa18F5zpiw9DhnpL
b4pD3jRPunoOr+DUA0+vyvQW6ufW782MWrnctchyztEkkpOwC0z6ZrDLiqOCk1yj6fdJnZo6MzE3
djJlFPU9lszuLGpcJ1gaXwvArw5l2tGljpXGjAVXUOgkabTZvSysd7gKxRYGnCUx8GKyHnRjoGmw
ie8Av5tJ4AgXfmZaPKEhPxFrMQWW/G+LKWv31UtzzhG7QmX91F+I3PotmQRq1Qe4ad+GuzgSrMsi
ABig/gA/VhL55f/c+uqBxAhOCU5ZE/qd5yoC2yPuA1AeP3lIPOMCjJ6yvCYMHfbMMKCacM2PAFEG
qEtbejirTobgCtWqIDt4Xzu3D1E1BVMpZIzvbsOaBlykutiCidlL2YkX3OZkY7uJwaFwQ4Rd3F1G
SaOzt8mtXIZ8EP3RJMDkCl72DyArS9s/FoU1I54Pc5tAQJVZIGMWO/+gRNO+c+ELUIdabmpqgwHy
W+5x9b2xSCa1FZDA7kygsfbEiICsW8iB/7iSs/J8Jw1lYkQsGHNKVsjj0JntiM7/6jqYRU8XkDT3
JQu3mAYqEXwIcSf5we40tHYOLsWNJBW4bob/RYhiBy4mVehOfAY1LfMJ1u8duudLirWwEnezZKaH
mJ1mXWcwOIfzHHTOb9SOiQF66R6byN7Av80d3C0bhNlq97Hq638qYSsg1Mh3doHrwaSDP2DJS1oa
wU4QlkuSqtOsiiYKAhOhQVsYfRUBAg957zq7O8dHZQjgUu4BdUa17jE7Y2ci8fwQFOglc8p0aqx6
X3H6c0L2Rvfpux1QXGDv6zG5LjzTbx+9SIPTCW+2iiQQo6beKnP7gdzG8puLDIdyvylsCsB8VETv
L+hoR/v5o/EeAbOkG1o9ayMJom7OBWXjRdWa4DlOadGQL253CgTLgEpUvrdnTAbCJBpC2lynrSub
cEkCKhuU7ZCcQyp2lH8QH8ZVMvESZtogEr6xIJ4r0kkd6u5hOmY7QbdPCPjgNFzVzYSMpnwWQWFq
zmVBTRQPycjrgyitVFXFPjefsviUPDno+ds1mi2wkX+vPME4pMt6hPhHphZgJA6o5ZI/8+X75q6O
w6e3ExqFKQ0U46hZvePCzg4v05YZ1fD+uDegCS8BWUp9HWZw8p5PLi5FYYUYevcludHUwUAbT7eH
VP8LH7o3Va/z1zeGkjDGXg8OW3Gm8Ei7zNSmxiDQ2lJny7nPdym/G+sL2xdnpIlCPTxDLglftHfG
ECQIP05qasgep7FuzlzOhzP/XxoTEogjslZzL3yyBbYdoup9n0Merku42jWKgQ/rzmW16fJ7i+MJ
/3JyZ06P73xjYkNFwONKYqZgk9v55QRhoubWzU6tznuXbLpNUZSO0zhvoULhAOF4xkk8WCkNKYjd
dXVyyDluyD3IIa0gIF+PWzq3HpFGwaCW28pDVuIMHf+3ENVcXN2q0Hapy77B9zAicm5DBIuhsAAE
dNHvSGdKVtR8ztRmmWY9k5F4/I3QgPBw9/qp2msxHFfJBP3tRTHw2TgFneirIe5Rv6aTBGRfyv+q
/18rTLPrnbQuxdARJ8WnGVhgw3VPFbkXNO3vF8t/oFcUI8Gsgu7s1CofDJTLV9kpceCJxjB+bhwB
Ks6AeioR3IQiXZxd4ayi6JfZydc6yYMtM33/x7KN+ERRxBiR6xfj6/u/pOLXeSIK5ceOZ3AEHsRv
0zx09ZpsuGLvD1CP+XL/O/Aatd88y4CC2cG31u372HCsTJvcM3HqmpC0h+iUytrqCjexdUUAjdUW
Gf9XHFkjZmfFoNcX4ot7H46eukK0RVKF0sEn2bwye/Fw2zwZ/xbmA1RkAB3IJIh1vDl0Cm+Cosae
6JEdmFdNUTLYkHq3k9jx3uI3CWyhSzvxy7ha1EsIGQ221yitRLN/Pm4JbQR+be0ZDVO7h3IWRJFj
mr9jUCcbCtWn7+peipoLpgqJe+yUNXKkJ55PAvUuXSgLsro/IQLtQOKJIQC2k1ehrab6rpaL0nEL
VcrXodIn/MUvXGnYJ2prGpVhF1wIXV2Xb++gMoP7zxiinDBPUKAIH+P2UCcA5L9BuZzl5CMJg/OU
UunK+a2TzKG6e6iXwGiRKIMtF1KndHo0hoL2tDCHmPnnAkObhvRl64Qc8bdfRih8g0WwNiNSiCH+
fYzfoRdByK5g3ffgIHRvAtpnhNiae6qT1roV8ZbIeHuETYvwdzdKk8RMZ3S76R/aU/iJ1zFvQcpB
XKzFKZmNP9I6MdWVX2HMmq43eUaGkEwakaI2iSkGDSQweLIdcAR3YuwGLE1WoglVhwY7dH+Yl8J0
VYwDrth6NQa1+TOFw8ovn/Gut4CIVCrUJeQCo0kryaeSU5Ac4SmMZkps2b5Or64Hy6K7+i//t41S
1J/5NoF/TuIaCqtWI17MnldIQ7j9lkuRkZUPxPwaF/eysPMhPNKN96NRngHSd9Ujq7ig0BMyCB7T
rdJhQjdDMQ2OC041enV+g+MI8Gjt4kOwbX6P1CyN0W899Hic4WdlpMnikyWOpoANLGpO8ylIM92r
5Pu4An8T5YnOd+w0FwoNaFtlWG33oPmp1teJzgQ6JEC4Ev+p5X1rRCJPpYtvXT6MM+Teex38d7u3
idIrNvmFD6/M5SpZh9Jfyi4AuVINBAOFBakxyLIu1wFQTm6djMJGlTA6zoP3KtwlTpoOBmSsL6PI
Nkb2KqoA8wAde0EP6Ey6p6SF6AXtdAVNQ2/4funLbIUGATO/gg9Dtk8DmXvGaeut8XnsZIUpQW7N
ZzGunwl9THSZe3F012OCH98ERWrWbRXV6KPe/e2jgcmV1BpPQdiQYWqV+t75bcmlJmSbiWQ6SX0f
Ca7s8rXY/6Rkr/V+X7V6K6764fQw2ABlUkrf40C9z6vJyhXAwG9JK5Rc9KORWjPt0vOnEpjx5J0n
3QOt36kDIDeVJf4isrruFBQtfy0VoNiChluuba0wQLcXZW5vWE4PXTvUWXVTv3XiNgGdhg6xp4G0
Nx0hCv64H8kw2e70Z6lzeN2cZ62bhRZsFElYIe4lkGGJdtUc24b0Ga4OR00QrDK9qagnHVgdCs6a
BXEQ6xSkmIkCRgLrgKJB0qEXjDunr3R9qWJYS3GjiIYa/TocWXk4HpMndAqxXgPCtukfhXG+z7mh
yIfGSzO3aXHhkyCyhZqrPee4JvneY/haikbl4ZatWO1koopzA7qABITNVrTrsbMYbPQUCkfzL2xW
tfV0iMlJ8jzzIldRIhuXF/80A5E2Za+CdMtOpK+9ncp2eZFR0kMGyZNAgx3pzQdzdDxXqbT/Gcvu
3gazxV8zz92HTRya+Q8MkfDkP370IY/ivh3qVL3MFpnEShOnXE8e4cwgd702PWCJyTonOyaD4xwS
vfHrAiTuGjo6K9ynGPMbQFuCwclscpSBsbhlbMwcC/uWFk7SP4DIXyFoVnCDqyDMxDBfLFYf0BH1
s/H1Rs5nonc4ijbg+BoKSNVeoC+/F7fm2N5pM3jGtvzZ2I+rGNit8EESKtibdMeG/dhNddlqWY5i
iHdq4RgY9BcrLEoAThMp/rEyQsIdq5scVSw86BvmnF0VLU8oyk00BqhpbNvhz2RgQxt1nOmAoaUE
202U0J2aJilQoawYIpqws1nDxKSH4gpV2Ka9Y9148oANftEDG8Vcktv+Fb1NcKyWVMnjevm0Hgmr
2gNhT5MaGBWFM3s9O+FVjQqVte2GDnMpbqEQhSFZ6eM6EVaivCfToI/56smV2t+su4JiIR86H/Fx
3OiIXSlWhQ+u9Y7d8ne+7tZeIMcHrMoZqf+PsFkbp9V+Qdt2V4BcG/dL+iaqh53+uAPU1pkAeUmX
9apecTFB8Gq+e7D3nGxy+w1FxmBBb/4cyu65a1JR6MZjKlz5Bbha/Tkbu+KhQERihPo5WGFKJwDv
el0P66Vp1c37iR1A4fm+GwgEZQq5WoBKDM9FPhYYWOjjZ63nx+NX24ZtKnS2ODvKq7RC0+WblEfN
c4bNx/gygh/uvrlsFpCjs0hHfvb9vkTfjstLKv9hy/pXH+9iTB//gm90fds1Ohx83NB9w+aoCUva
EsgGJFqkuqQB7012A1dwdlrR1yfOqLG/Pnqc08tKxR4M8vR3/gB0Bq61VIB4AvbMKea8bH6utNmA
4+LMF7Jh3VO8YJ/CONS9CgCLSkBa9kmk4nXnhOkGtC003YH3QynGfjruFGtofo0uHeXnjRt/P3fX
WUZ1JT7zIuD1hepSWjbfq/FOB7dpODZaKydORwPlObyjVLiKyLCXGDcg1S2WEqPMdAjc2WiIPNVK
lTielITCeNxlOSx0CCcBD72Lc03iNW2Gytk4vCCrs2uZlsZPpiykKFrRFva6c15nJLZq64Q2OGe8
1ObwVKsmKAw62Zfx1WyHWlyE+t0CQiRx5Q1KzQI+AE/OalxmGR9KCnTMU6zeJkxWxA++boPxTTeK
Niqid2bs5mHiwYHLRJtUnDlPzS5FkJR6UcPzXCk4Whhs6S7HCwkITQzjJJ4XhwYrg/+8mH+5w5hu
xp3Xz7BwkQ+Ydz/DGWBp7U2EAJtbsaMjbx6xfL9z599XskkMRfpEUDLp4aBqZZNBjFH5Sv7mab5n
ARlrkv4YEeFiyXLH2SBZq1uNg9EJYdsuKpeRGNVSblGJGcnJlZ6rm7W+yXa/jTyMK1SWQcoDa6QP
lBBAPpx7XrBXwwXvk0k6cKvC6MI1rGtDFNcuqRPfAYd0BOTra4E7SzQPymtmCzazJ/Lk8+vEes37
1ykpzQshCsfMbZPCQNdLw5OQ43JLqZ841fDq7MEMXD2Vg8N2PTvZlx+BJKjinpZPyu/UGj/ZfNKd
xJikUi1AHRWbi6kOKljqoyhfqJyXg2BpZ8nE4eY0VsVr4eAskjn55KobY87fS6tR8Xgey9dIdXkQ
TPbFN3J4s2etiOVMw8HrhWSipznXZi4ct7GyW+rmR3Is3YwsAcATRWhA4IpkNOWTi5/F1h9SVcq6
58U0wSjUsL0XfDWndTdorbww2JLKdgnS3zw8vsb5OmY/+c1XV5zT2DJkLfj4GPqsszOId3D02w4O
lZxjwbSRWE4IsNThHqsJqi8Qqtam3iJZemwenVh+VSqzGWendsKSt7PxnY44qtMxphC5FQuyek6+
zbjwm4FxaFmx/12WLF1T4MxVAL05HTeQauVN7/fccPDAOuNbkHkoGdBWdQ+TC2lJm0dVambs4VbF
9o1p/wuxk3twIrTkU+cGQQtyGr88tFVEnvzgmg2+phgsY/Au5DWkGTdQCPcZoVxPZijX/p34IxDq
F3IOHBXERoIsJxYnhh5GzSLZClASTI6bgBY1R3/rgbN6ypgcR/Tjc/W7vfUgo/bowD7TfxU2NQul
eXyv7Q9gBzvxnqBM5gfilTiBxL5iMFB/Uaceb+o+q+QBIXohNcbZgIULE2l+eZ3MbrMYmRBd4/as
+VGTym1SwAcCTqx4xgnoq6Cr1/9j2s9O9J+zgGjI+WHJI8s97zRYACo9WF75Bg7dOgfhIH46S6lz
vR3GXaYnxBgMmyRc2w46+aR0hjqMutjmA9jUYc+ToCNuVl+9YvxViKfNESxQ6g1yKzDTNUwhLULE
R9Wt5X9p6tUf91XRMnHPO4ANuzbCEH5rad5mMKaZa34vANehtcB2U/H2dINlErNiYzNSluRz1yuJ
OooaelkodZiwSznTf5VcCEv24w6+3FTu7UzoFDybvQ776C0Vhrgh0C4c+E3cWgLJf+VzFM/6RNn8
7TrWyllEjuWeMvjklQ1fg4ai7IEDUeK7tcX+ABPFQgbSXY7gfYnzDCpHffIRd6zdjJI2Nj6iv3CN
3AmIVbZpvazqRadz/NaQrnA8kxyABg7OdWwGx3zr8fxSz0ywpwq9s6v2n2DMR00Fa76Ail1tjswF
7G63gQcrjPxBDxs0+TDwc2T4cdlnBx8/qJwgreTB72JV84b/qIBtoStZTIYJu1SDm/qu0E73Mkw/
iLpeFcodHENxAtG2p4pXO/+NTSZotwRV3SOH/3Bzpinl4rb1bCrK1gtMF84Qk18jGFXjRI/Zvj5l
auHuQAs0UCKKIii+Vm1S6To8sPKVsXCueVUC5s8jXfS76iKNF0/9iDIdVKXpM++LRsU/2kXaNM3k
/I8hR6KdQfF5SKn2dJtuyq3O+LOpNAepH3jc8FRXj0ElEXIGbYAukFP1yxyn7NdtRpQmdvpRkSZ8
7wPeLbvjDqTkoC+JqqYhv0x72H/iqCPDKabW9G6tVQrHlPe5mWdNg/eoDCjLGoTF/clEkT1O77+A
VpWDakO4/NouSk8mogw8A9q8jf0jXxR2YFmnLylbSkKRQSMdao9qlajoL5wsOrWrXKH3qI4U170k
OzFspYDjBzouBbDgci61tP8TQFryQRxnLrtqQBbdSgAXCbZkYsv7oime7RN7KV3t+Lg6Xf/V8l8Y
U2/GZ4sfh+iFA/VvtMFaPD6xZt/UftD3ylHfHiFiIbHJ17Nk35kKpJa03q6cYgc4lmFm9fV32LEb
BmYPdjjBcFCPLXVZj8Frk/Y1dEIdHnJJgNdmImDOSpPGODq7YxjzsScaiHbOcwC5zd/4PDUxQzNs
/QKWWiOoIxs7ZS4/96U7TpI1k6gF2hmL0Bp5wgQJwSguHIuA2ScaVO6zloIsNfqf5Dfru3CSasao
Q7clzKa3Ng3j1nIdiiUn8OWHHGoyyzyzuP4wLv7gooFvWGQbyrz3kniBIZfJ3qSNMk3qsTfNJuP/
YiYm1vtmQNbpj5ZMIksXxBQeN0sDK1m3wC0MCvqRYOoj57IfGW0WwFsACi/TbnpEbnUIyHUx1zFa
gHVbA8gMQ4xZ+sgjkcYmdxH7KNjhHDqn1vDavJ3b6mXqMVUGGcNU5v1z88ZVeyGkJwAmyhiUKw6p
7BZWzhUep1WvRAO1fxuYW6G/LaxaabdxSch+MjijUQdSs1ZfQ0PAbEJMm1VRO6UO3eAVpIGdu+qD
PmMItmb5NeUkybAGtMSbhOu83gPo8G2PBU9KLIyQ7DeTOB6tQvfT8WwBGVy2aL14Kehy7/meq4tw
7by5DqJwoVHDJGKkdtuSDQla0xRMnSUtrJq0P4NDbXm27EePclJd0rD2pMJ+xf/kgDhsj3gzuWjI
ThI4CNlD0CVFwzKZTa7FHf0UziQzdYWmgK70kVjrQ4CTjU8EFvq6FIfJOQ3gVdySkbop/SdCEG3k
ahUTdcDVocBXDmW3KEn2SeUPi3zV+FbcwiruLiCVWiC5/ygU2dOxLiuJNR41i96XqGulM07PoUkZ
cDSRjvl7XT8A1pgnIfN04J2RwDw4t3/WbgqJoLnzYcao1gKQo/bZ7L+zXV7NiUQySCGLOofiCRE6
kWaFA21+5PFUMf8sNLvSZLTCpSneGWmMm9f7KEZ1zYrbeXHaEzGY1E2Q3VZvjgkQPg2MCPMlhf1R
dmwpoUHas/fKaNfAW1wOiajBuJWNtHfCq9K7+8LRjAaq+aAIY/HUNk9DVxEyb4dkyC7uV/Xb1XTR
3MGIww0RKGF1cMQ5PVlBnl3oWeRIkD4jts9WDAM9pdq6bKJd/mwfZoGRCS1gu2TdT2kYAKFFW5Uc
FXG8NSo7Ya3ixoD/kSnK6XoiSmP/IVrlPDEdnTz/xxuB32pWP4OZicNPFaUooAtI+HZVZnEjV24s
OtVormx/FAfIpUZ0i90+nkQ+4D8fxk+rHnWP1uCv9a3Xs90k9EFSK48KMCesYZgjacsV8BPVeaoM
qiYQ5OAmPTshdojsBRbquS2pXypBtIfOGWtHQMQoUBQxDHVtNYK23jX+QOrMd4KlcTrQtI9kKvIV
sv7cea1/+dihm5b0RR4TowZ37/v6IU85RdCiFg4UckJXr8THa7NFTeNL15/tF6J1tj1E82fZQNab
mXP4/jdO58oZFUOzIYv6f/c9pSyHClOmwozueiV6/7oxcsg8YgYPeQ65RnF85GFClkA3DAcF+4/x
UcT/Qh29VzAM+mMyhHlEaMtK60Sb+X3y1f7Kn/HkY4dPOKiK5/itcP4kclfJwxNMmVE8LzAsoKJL
HeHyfg/58ZfwhcutvwEPTnYAcq9TDH4qc57+7tCHyD+wg2gumWw1vfl08QzuhmsydvERScyzheKT
0cGS7l9Ae06sXcK11zOaAHcGJz6FOCuNfLTZtRT1ieSwL3tJjOn4k/yJWAQhCMSWEvJQ6irFey0F
AqpRyifuYkosNaqgnts4Ncm16l4TCg9L/NcIkqUpVHVAMikKAVcBBmT2x70eFCN9WdV3IuFPkvEo
FCipXPQytHooeO0lJ3HBAr544TvTsf+K37YQmNAQeZ3Nhwe941b2El9VmlROO7P17YvyenOnBadz
eMsEtEnruyuFSxUviBMiRNnCMipg0DAoFrWlZhvhbJaDqBXSX4Nr/ouHqzec+hvDXO5hWmys52Cc
EBiiEZWzh4vdkv6zcaghzP+2uRLVWf6GUFSagQMTrwTpAyLt5AJHSmH8MbUJlK8IVFwuBHJjLxQA
OgXP5+Swrt3Z5QPl2g+ZFEBBPEi1q4NWu80btk4N8/fToQmxEHJSYTJkv7PaaA4FBHJzdvoeEPiE
RQJO4wXzBvNvnBJU1Ngfk+nR0IuIigYlQUnhaiN5DbazIEqHLyhYiQ0wqsjgwn8vb+3ew8mZIEf7
p9VKjCop1yofxvQBNzbgsu9994Je9yeJp1JYk+BZnaRcyE4+LcrK6QfxKKPan+XTaTrlKt+wKA1B
0k2L0kHtZzxIVUeYxAcIg313zRuzJxx5OHzTsTaOvjxNfo/aDrjmh4aabtHsX+vPDqU7Jog6NWXz
PMWXTRsAmL9gd+z/JTy7nER22SJdOfT44nYm82K98XS1MA2bgdhFZm2faHzPFQ6BhdJ3CmbPzVYC
QjkUqw1ca+XQuOUSPunhVnxEg8LKO1Cyvkt6qwnsYl2RYLH5OGxk6hFjMcxMHTWPEdAc2JwP6lfE
dmWa6v6A6x/hIevI2ayZ/itW2hUqhGFjPt21j2FB6q8YFdJZw+6LHhYNwMGLoSf5RGRZJvgzB3zr
01rL0oxHpAAUc0EUvKIUhF/A8qBOhvxYXwOwFmt+r8SJI+K3i28bcsxvyE4Ve+vfE/XcEzXduOQc
gspefAqV+mZQcGwUz6guis+F1rN8mKvpGQcCBMwr/xYakjzYXUv+2Lca7KvWznh4Zdh9tltTD40K
PpNQbTXVV9qMjo5U9ySNYStmucBqOWw6AG02d4IHE2Q0HZsn5dvshGKm79YtRTERZflGG4uxIurA
/nnytq/oETnjqczLPLbIjH7oDpKVqyhQhggKVR6/Fj+RLeRAXlqOS05KLJvlIUXPtCunWTMH0BuX
geBV3AwEAhI6WxqYP2nk9hAtygye+Zf/smc710ButwAczn48WYhXRcl5x20dCZ/kVPG00UgdmcZ3
BZ86dw7PjBA3h4oPQOJuXxhSck92p/TmJjqpfoOQmU+SHvZDmeDf3sCozOVF5vpwVM0Y/IwzX624
dIfbNh2+DubYgPxew+rQCStak9wlyFVM4u38WuxLoUmJF1x9fRlsi6i/7xuXee6/mZqbhCF26Gb8
pvTfaakv9gNUoxV006SxwSmeChGA0QJiY3K7A85J5i5GFl/rMS8fEf4HPEsc72Ilmu3rXwIXPMba
R63U6HSedT4nU5L3cAR+P0LCWAy4Hk+n+pemL6lALk/Cwxl9SazgFrng4+uPK5FXmnT5AWlbTQa8
Tib1F4hz9Hg7IeT1R1IjLd815vgw/lvP8bdQ/dzXcxRnWtalzKYxnjB6o7UzX8gE/FiwyahESIif
bIa3ZHeIhHTd+OpSGK4BnjvQczzFfnTO23T5gDo5Yw9vVEPU7SwS/rCprQhbe6BQQg75mZqsRlQv
Ylw5NI47ZM4gsIFZaJBi7E2MUPw/gN+dILfVsTckJ3gdFbKi3UD6gWNIepFqeEV3IOvNzP1rsnf0
8muES+R/3eea0MlTXDizbiRT6N5+1Gi1u9qCTHru+NdD57E6TOvM/ARkUs8DoiNtpDDCjTvUzdi+
BvqyqmorQvdoENjdFHPbRNAfY6kEKLGQO6KuuHQte52zattS20aqQBtGY83PE8zX9m7cgVh743eh
3X9HOCARQaHtJ97Bk3vHr5gJOz/uQSFmAbfFLTP4T2kXY5DWV0GXhhn7Dgt6kjmCGsHskBVt3crZ
HwWmoyxQtEulOsogyuMpSXzLG2dSZrco4ROH3qCQMx+lN8huGW7wrHicM+skTTroZBGi5Of6AXjT
KWDwSCtd6tQA7nQEpqPNaS2QXTe5JEBWNga7/VqIYw2rUUfsMgQh45V54cP4c4j2JBESs4BvKsbq
WdyBpTXY3RUoZgcnrOjSrpzvqH68oXj5AvIpxSI4YyscWtDrdSrUJ/ghj82Uh/tZ3XfqGt60OW+g
bTh+QhFAnGc0t4ZEMg0cT3G4bImNR6fHL61lFDyrcact1FDRgF6dYsO6HtQw579FwkBFtyJJx5F3
r4/eBpSnrTGGSZpT/3Ejzx0YtSck0wr6xKvy5tvE3xBOFav/NhMNfsnRIlaqtGevG1FQnZoURYsX
baMydxnZbHL+fbbKrG4KozKLFXsncQPcygbeIhKm7bR9GwVKHWeBz3taCiErps1UhJT/FHLIbgtx
qYWf1I0JE+qw/3u4/njVd9jco+uhOCqiiR33yuFtXL72DzMkEj3C/F6GlmN6wZERROurB+hu6WdM
ojP6RV0yaoBS0lHwclrNfMdhYklPh0IIYOQWEb5orJhzk/3Imlez+e5DekaAZmMjoyb/i6aGV6TC
F0squ9m37tWN3HAWONh6IzznG1IoZJv6TBM/WrAWGjWregk7cagXAUCpSLlF3ggHIGb0QHEuUlUn
Ot0Eg4nCTaVEef9Fli5TlWv8DtbeUaLnV061Tf4+mYl+Ivh6lKF4w7kkOn/iGrhAtfDQ6hniwtgW
hTArW3tZ365vkv6w7cBm8s76S4yANuR7qD0bDb9t2ir4mnI3ih3ZmG+9XXaDYStf6CtcTIlCckPG
88GJYFT6P1EXaaG3jDQ1DEjupmmr2WZ9HCVisvVBIPB1WuZwqwzaZbNP4NBa3843bUy+zHeFmrkH
rVt8DW9UINeRMkf3/acDaeNWgMLspurouAQWh5iFM5jjZxtYv8Pn8dSr3xwwlN5U+YCgJY5N/W1f
cPF3nP7GRW28H/7f+amScRXpBmNIyKM9A1cFrcpBMYnwxFoJpT9+BeRG1bYpNSKmVzQ4CR/82Kf6
ivotZFy2dAW5/6ELxJOX8jgVbTI89jT8hDBCPHPccw0QI3cIWQ4BnHvtHX61PKU+dc1qVLInhpIx
JFhZc4wqijU7xuyfzLdh+ogDKlmZdDNlpjaNmu/B8FDPy1U0rm8bQlTc6Zp0LI8bez9GdcOykIk6
GICmXbCJr06IGXPaV3Vdh4Q/S2c5rBf+qmvTHz8IwqPV8VyN9kpVN2prGJNkFYgPg+j+MEfP5iM+
MGVV7fpMRtP8xHoOuUwCGNVzskH4F3HnqoXBUvrbCAK6c7SanYq33LqQ2jWLy3gpRUOb+vKSqznm
IoAuF7FRpJDLkypmrCyCBjObUyLivy19LEFv248fojmgMPx/lq/H51+bunmLZ1pNxvAkklQIXJ4b
GJnc3fhT0m2bz4sqaKCH8xFt1fVgwVenrtw8QsDd2AZMMBW/K+v7xxqzIVW9tfQW+7vMPjsgcv8K
v1o8GMXw8ZGg1S3XELU5ucvgOLwDSz1HjqLX7WmAhPmi/mMDieCQ6ccPonLXfIwidKU97WRe+zw0
T+yNT05TclFKN+GrXfezbmpe3RnDZ2BHqZM4LSiZAUBlw9eRo8m/6Iyz554/VE9hN0ZkBHylEfci
pC6pfmFpmf0TN645KCY9JNM72IjRDbceO922EWtEK0Npq/OP7bR8vMed4df7GzqYS6q0V6U/z3bo
f7lZm1sKwl9csIwwZYW9bW2A+KLUjwDcuTPK/x+U/RgBk7OM1CPwxyHv97/5X1vPpPV9ZGm2aAOn
CyR4uk1jDwgQPIplP27lKehnAoM1e490RzhW5SM8/X/tY/FfUI0NwOZCI4U9UjN7S12PME/DxpwT
aUjWQcIimb/f1GbDcXU9gnInFGvVRWrPMI6mUz2N0oamxEb+35DcgzvrTJ22GVWaFbrRPRBh4/A0
N1LYlNPzdIQHZqF/hiRUdxqDsyC9cousWOhHuqFyABOHwhf43Uqit0qmlcR5m6QLyq9zRrICCb/g
VclFlATc/qtU5deVZDDCfhMVaLmLucUaBdJ+z9GYWcUimzUrLVqsZ8us3y5lYrtu+Wv7qkB9vMmG
7PE8vRDvTeK7rgO3QsEatBkWzcqi9hHJLNaitjY5LNE/ZK0ljRwjttlUmzNF+apIiLjTHmImcDI8
9ThN1uYHck0L+9OyW9lclrR7CHs2MpFEzCcVwVvcJVvURSucbAXibKRbehUh+a9CaJJatcfJuJLd
CP2V7QEY3t1vC4p/wEnq4yP/HFnsLeY/5ZBapAw81E12mscq+UaGtf9U3bjsTIU/DP1zaMbidV8w
Bd5x2NxS/+YZXrEvD0v10FNBTRmfvlK/+aC5vpEWlELs1y8RaqRZwTlG3n3I0JmjPdt6XGe1dGPr
Rd/VeBwJAe1km9+IxeJlUbYepkbQlEUgl/+ZjPjVBRPa00vvmKT/Eg4aFriLQ3z8a3HtlrpBhXde
WzAYMyln9VZeRQnqRC3k+ZUKDuW3HS5Gh5c6wlYMbDY2Ix8TEBqhXrMf+JNuf5KEZ2CVO4UA1iRO
a1PXR3/PvJtDc5HaGgmN8hvn3KalhHuQC7Nwb2KmwRU+WZ0Fke/HZE0gwRQiBmVoEOWi4iV4iyiF
q1w1PGUlyQucBCYsTMMj0BfQyE9pROb0+65bbYLMBAIbEQBAk7OTRrDCrIekP1NyxC7UWVT+gQa1
+JLebttbJs92ej6TPKgOIxOQYDqaipl/fU1pbevsodEWzrH5djLh0cIkxJUvA+mObhKpeeSg23tG
BYOiYkKxJwfzsFa+/mnsJtMTXt3To72ps6trrJJXbGOKixnZdrbsHioRDUGfsF8ColkkLSRKZonj
PT7MeYCpDhCsSLroWbN8y+GJbSY6Ho+JdhQgFB3MFIgsFySb9ZBlkdu0TI2eUE3CaxtniZkafcBD
nwJLQnV4ajNXLiJ6y1yxmd08zwWu9FvW9pUZGv5qiP64cTjD6dcjSeVzsoF+4taVRiiReb1eEnvk
OTQack18I/uucyyPItJ9x6mbbnah7Dzebl+KqFhqnP8yHwZ0lf5uxRCI10LkLKE9sqWLA57z6a/H
g2D4Frbv0VJ+aEuxQtmLQAFfGIcEK0L3uEDMkXEilxDHQzBZPbBF9wkmCZT0Iaeopz7fa/4Tp/RY
xKA4HUWNrHT6N1qUOt7ODHnqNvu5BrOjjTZ+ieZrBZw9KPM0XiyjOaW5bWn/l3B+Vv8v6p/M5IcV
JxBqf8UvLk5keSltBfVi6KXLYI4EZodQqt/TVpZEGOryCz2IJDSOCGBwzhhI/J4IWRe5uw/RLNtY
StLPti2+ZgpI3x6GsgVT/WqNP5AABpRwkWoq18wa7YXIsjPc/RWCTrqJNxdZ/8m2EUXqVf5WcopD
swIPr8PA8SFCYehKRYPVBDtQ54isD4jqF5gIaqYe7Hltc+B3y6NsvD0Id/DZgrBwjzMiNMdPQfrI
c3X1uL+MARNdGsxIf5ixubzFQ3xCKNwfmdogMJYtl5x2hQ6mK7NroILVIiZA03bpfb/0jsSVU92E
tm0gRFfzhOQ/l9XhqKbP2uMYjoX6ID4VdOESOmzDtNkTNl4KpyJug/UE66mCpa8v8yxmz59OJxbg
T71obQXoqb+NXRqSMfgUOlkP/VP8Z8tkPGu6TPEK6tFCPRgHdWHRIehCnvUilZ6IKvAcRUF79jbM
oSqNTKK4gQAXH1TeDrz+Ikecqo6OC+FlWxcredpPKD2LBu0y1q5joZmESr+6haBEWJzibEW9mNaq
XEbnKu7Jsiw8VqKUYJFkBolARu+3dl24snn1rdU2655GZt5mSvg9M5NB+f90tQyqbLHbPGFHMuLB
xKnFJVQrpyRRBV3COuI1Ty+sv0TKmW7xNe2YhnXVSGgYwMViHAKzQGgSYSalw1ejX83tA5P0xOMH
GetWWoYju6LQa9GUKgYFyCNTq9YcfFpW6EJ5F4M25y1eqLyv9N177WYER2MGJTSIeQ1/LfwdRdDz
Jo5tcYS3u4IAZig2f9xklwAfpKYMr5uPtxxjoauHVm7pOOQA4LnSdSno3YuWlO0VpVEzvSmjQv2b
gnRlz9HT7K4EgP9wgl/O5wixU78je/7wySsKTSX1S3pSOSbgDIcrTb9sj7MHQ26ZHxCNTLkxHua4
Jq5dBvKRX7WNr/XklyH7UAvhIcg2K0qs2pggGwEnHePyr+EtVepgrfQw8l/avjW0o3M2Df0OGQp6
GEFuOY7dJAmsfzqLd5p5uKafBfHQ1GFcHCOrrCrGeZgpkAiY6mwf+tKOORo6/ou1wbf7xYCEHCyd
j21eAI1lMJHsPhXghdg+0oaTkDV9g6IVH+UEe81YTQYwRcchWGNPrY2qcoGNlx6uFdSa6ZQVZH0Q
4GNp+B5Napuv9vul1jRcVUny+3f4v//ASZoxKlII96PdS9WwNypotbckN8BLG1Es0TokRp6ttYPl
u1nRs9NFTXTUx0SMGvl439ep+op3/dF2GGjEsBningFXSTTnkF+E9vBM+Z20uJjF07ySiBb69ZMW
PG8SoDppM5Xx4MRy7BC6u3wHFfPWPR7bFBXcHUr2RiHLZRnCIgVDFQBoKFCA+sO8PmZX09Oo4Ptt
k4DldqIVAqlbrIJWBua7b6PP608zP5fukYuy40N5G9zota62nDIr28yNkSTTHnPPMJOcRyQMhGDs
iYbUXgtrZmV7F4IcIk5Wc6S8u61m5DOByUR2cmNji9GUMNL/eDbaq+gg/O3b9VHAlS7dYn4QLYUX
mdnFqh2eZOH8IFEUcIOZlf1pJU71PRpRWhB6llkXm1C5/k8fpm5GsQZIUngH4KtdLFAM7eMK5Whr
HEYRsoDpxEuCeTih/K75A5olAxy5J/VJCOJhYKGbnxRS8yuQkDv9vM7N68Ve3tiYZX6pbozOIeGQ
RcxQVBKREHKAQRxQHocMCTaQGpjbL7T79ap7WlTuE6tudGg7DkFP/fG/15JAEKCrBzSvT+1CBIC1
Lv13bOEeeM55fFvkecrq3QFu25sH08r5F9u1jhovh3liBCCCHVVwZtFIe6VGbHeNx76Hi0mzhuFx
4kLZ85pUJW4Oz347gRfHK1YC8pDjw0gi3N1TWisOcEE6qW987oJTjLtCPDPMWHzH227ZqfoGUyrc
Li7aM0GFx0Y7IEimRdPeAbM5Z38gyCfXvUuM+8e3Z82YvD5YetcwJ9n4VjV0Y0bTnIjS5+E/z1RA
M6f/dZDV1knK/Ph/rNm/E+kl3Y05LCmW8WFEaxcrOFSOEJeWWpy/PwpFXlVovqDeU2a3zy48XCED
Pge0SyF3zhq0oEpcGH9t+ttw2eVHsojB74mc81c1mDz4V7sPWqNBPCJCZ64UPCWCgey8LGJmTe1j
pVErJ4rLhsaZ5z6HyWf/LGJpA1/ZMlxzSTSv9W1lfGF+Tt28HShTeUlkIpdRX/oWvCPHHBI9vwdG
1bT6JNyXnc0lNGhOvNZ+cUBpF7eCoqV0jO6C7dSyI9QCILQpjIMxS8F3md0ZG7UCpdgCMyFWk+VO
Yi1jl3Jur8KKL/CwsNSFTn1z+mIjlqJZ7mPoADpk5eQslhD1H2gui4hdbY4H9PKl4mTUYOAkSBgb
Q48uaSCmDNUT5eTzut3D+WY2rrY6epSvp674mOhuz3fw6VRvt6q/uBAw5XgHYR6WhLeXt59CwbDB
7xfNUEg5sFrq3Kxey3fnhDp7MRjqt79qy6tYdKHMy/Ma8s/h4pPlCIF7Gw4PpXdT5MBD/trk1zTf
IpD0r6fCMUwAdsW0knj4itnnu084ApSCMNqIggpBeOubVRzgWFvZbtYQSaKRTZ9wAtISVCGrntZr
VRPZPbVFybkEEo5iuXLEF1nwgw2D0vASCWMCuVXMFDnhjxWNQKPT2OC+sSpfsBHkCGUhN6iJ1lPc
1rSZVWigRf0QDKpqEyfNkkTe3F0aYHwY6FI5Y9h/V06qBD6wwqy/7JVq+iFa2ko4wMritPBXct6S
CU4lo3B+MXlsme73mvQH+fzpyz3UDA9MSG16mwS6hED+vplDut2Vbt70n2vDtwsgya4up/BaqQ1w
STWxiGNcHouZCT0oVPpzjhBBty2YdavBadsEUL7SAAOqSrxY7ZVCvNddEGaSRFu2iFWHLbHJjwCd
iGeyazOTTQOYjUD137tSEqCSeDAMJy2r6W3fp+RnDoGLP5kUH4xvTI+kmmsGGi8pjbaBDeeIDm59
A4lZJhYkelArWixRWY6IECDiDXuAmsiuAAVVxc0zzzQ8s6AhA6YRAApqTlohVZPV2BQ7y6xir5uV
t2laT3IlyV+HRg8N9KkzLLRI0z6R0BXZRbo25tye5xGRioYEot28pFO56+E1FQccYEwU8x0q55+0
dA3jxBYWnNUL3LsqOSrtb8UApLeX8NwXuz/rh1SWdlXAcUXVHE9X8vInYGQik9YvxlbYa+4gDn2v
LTt03lGfrEnBAl6apvIqd6Ojoeh33vlWXJrLJBlF/JOYceqJO6HRyc1WFQ38A2d/M3evmJOO8nyP
Stdc/Ir+71CWyW3/uuIfUSyE1RAIseDSbn+roLSChF8Pj32owzCqiCkMCOmKSIANgza4yuNgyTfV
GWqTM7cihmu7PFmMIfMFq8pFj8Wh+rk3cQYy7PPU8CP1swTpluMVDnH7ho7xQxMmUeWL8WQOPVrV
fix+TwOoGe5KSyL7vHgn5IXrl9qV2X15ECLaDtpWOJpNTgSVXOPZY5r0ve/0oPPqEL+7rqIJsbOI
+KSwSRwJZelQe80hl8HsUllWzEwWeuXiM/vB4tT2JZTuxL238gY+uhH924SzoYtcmtuWEQqkM7PH
zCy5gk/HDL3+5S1xkm0V2FpslJUEkiz8YWdyHZ1p/85fuzPLcYBx2tHM3zgK6kVgZU6+rxfWeKG1
hRkjx0pchc2gzj4Gl7Tzn2gU0czA2c5VDrhZldgx3nbhDVU0XzjlbcQboh09cW+DL3eZMC0OFNe7
pNI3MegrPmUsHBNnT4kVD6Nw9LT2Y+OqEMmOAlfjdN0mMhC43tvyJy86dQpiVdmoxGVouwSWlXW4
B1DNZpSn9rNcvSsTYb6UvehlUg7RJqD2136/M7nCDKoVFYVtiUlMkHWuYCAjTEbP9ho1XnXgC3uh
8I+C/FEo6qZG7ybCdFVEXBHPpcbm5J4tffCkYFX6ZPqzwPlb1W1766AAd2d2sgK7wOMfP0twfbjY
ncFef5f1C22TcwCIqGYPML4zrp6R8ARuxyoLqcr2CLHgb7Ipn4ZQdlB3vhD++tmqcDRpq08xnZt1
oAJ+fgM92on9yj1TukTPChx+5nlwaE3o2xocy8dvd77s+YMNMpQ3Xc5ZVTQIKQyUBJRT9GR72CnZ
8R8ICibZem7rx+ouH6jGxLXUkItKjJdlzzZ927snjmLr3tQ/WFxrhx2a9Uqc766M3oo0FXZDqbSu
r0rvWiWQrPKdmnBuhOAX7EdSl4zRYlx6JLgPOIO/+k7o87VCQS3b38qEBom/MYdfIs5IV7vVDf/H
P6sMBYsyQm4xuQ51c84jtJZrRgToP+iI8/h5DoqIiz1dV8EizLX3ETKpEHnETPdBWQxgmX1xSMh9
R7IyuavVNzuvXSS4czeRiMgpA54pHM2VPy2jvVknnfegkfR5UyaVEapKY9ydeZseWzvNbK01EU3i
bJztyL8x9Ml8/PZVirlD91+lgh3qnO2C36lp1hjZBdhtMjNrSIQS9PnWvphsm7RzIHrn+Uak37m8
ZlENvCCNAv1hy3BlY/OAgDua1UMfqyyi1mlXyKXPLmpPwLLHtWFKzT24YnprCXAFgzLlmcw37yEL
MwHlzz7PrGsPNLvORPP6G+7rVnibqaWfsUEew2hjshClZ3XSVzesLAY+hJRbGdV3ZXwlKm/q+bz/
8v948cnIj5fdGHMVEvVpQdGaGuQ4o6iVHMJyw7/8KZvWD4VT7omFxmzWvMukGLGDQYhUqJtwOPlQ
XSOry5W5oqAbNTM9MHq5j6clh6AJ77OqN0d7SQXSGfuViwMS3op+89Mxf+vE+hMjdnaYC5hNDhTc
uR0wh64ZPBBoR+J3Jpa1N3s6lfnBR/8QikXpo02h5u0Ik4pe6f88Y2JLF2iufvEZ/hgkQlZTPpOe
069UgnGYckZIBzKX+cP2N4hOWAxSXu4SlB5r0OMLIzJOk/IwvlfgBakTeYVDDqmY74meXmMcrQvp
2KPdAyeSDXuWSkh2fPIk2sXC7g64uSbBEaXdqILsDa3amubJ4pt6I+rdNKRizUnzacnQAVNlUwmY
As4vtjuYJMSepY1FlfT/wenfypTJJXolXoSgTA4a9yCXIvwmBGIacanFjlPaJZzahJduqE2ng8j2
AvtM5ZjpFkuq/b3LI9SJWWXqQqVOddYpQXkIvKc7Vo6Kf6LgQ+SinpK3Tkz8/Mx/V4+JF2DMED74
SDL3Cv2yBrLkOGCcgycrFoF2aD2btTkaSSVxbAdi9qvmU+gUuYd0gY2r9FqsNEwJQAzglggfmJx/
FABXV2VScVTqg2ggAXOSYRTf/3NQX0ZVGaDih5NakC/ALUj8Fu2FJFmpp4vMQ5YIaZD3Po+Cau/l
QvWqOZeCpAWSUQkH4jHbqO2KhI5+PU6ZU5d3QYtdtAniiSbAbj5SUnPtW1qgrAbRmOiEjLOoP9tw
ZIr/31UMsb3Om0P8fTdmvMvZRQRdxsRvGJqg8Mw709NgXSozvfldhHc1pQHJEGqDQqaIifOt4isR
jVO/TDyzoLesrvIdFjbv8jjRAmbGH2VtYMvmKLwx16E3fnF1zvMgEmXHJ15t4tqI9AGkp6tz+uqu
IDIH2xvWlbvEORQVafoIT6OSkXdayDUwc5+oLFqYhivanc4kYbUDNftw4D3UCkJ0zbpqy+1oBsgO
j7L4bIQjmEw817ViHTU60q2QA1mE7NzmA0XGXzOGhya/J6BskOysFPfaf8sSOR6nk0ZQhPSo3nll
OwjXTMHqCb8Pw08g/FjxX3ylekpwElK2GtOSXxy4ZrRH0SHFPcBY9SNJEkQg0K0EPmdPA+5MXNqs
DA8WhLbmEWEzwEuJ0U0xshHdOW+3rv1IaQ3mzKORHJjqaPUDkY5sGs+b+s30ijHJfhoFyE3aleLE
Pe3cc1eDzY9owJ6QVCkAvvHEGH/MFJvhV656yQ1f77Geh0RLBhA3QuT48QIwb4e2oE8mammBZyo1
JkajcC5t3JN+hrk++/Bu9NwKug2JsIV4kiKAYo+hzT8Pd5I5jKWRwkskeGaZcnkkIWq2Te60YPc+
Ge90PNLswJQycKnB4iMKxLKiHnKW6E7dWKll8j71amoyWd8FM97JKiaUzwbbI31M4qkgOvLRrEN/
tjfnw/KAHnK54n6+VsyTjnN4+DPh2pRKL47UQNMOh8NV0A6i1k87a2wYAB++EgKnLZR4CSSbPH2n
fmN8aQSD9wpi7UcXuLtbQM3qA4CjDwK0NtGtALM2GML6ME+rC30y0mxeENvtkLh3ckZMxpoMExRW
ExOPC17/gxm9jsS7S9w70lxkd8DQuKBTZwZkACJ4Yre+FvGEvfBBJ8MuhL5hNZzjXAj+qrSww7lR
cNohsA6+gP3l0HurxViBdpGCH3nOumSrPjzm3VAXPDLR/Wl3m5z0JAYYeCNwvtAf8KR/DTRZN9EB
gRHJDJkHcjDuRLf+ICGGGCF+SPPLPM/w0iYhksXrXwVLLaiLS/X0sjTP5t9ZlTFo/1ItII/ShAKv
8r3IsiO3GkOt/KuMLP0QjsbDxbtcaC7so1U9VlAyyEKc8M+S/+Tt/8hjE5IW2TGPGPa+5YMvEdXw
mwP9bWcbqw54DcsXWi311vI8nyqMRjlu8aRl5BC7nNpA+htN926EcQ9MIzDThSKrIQoKDiPzFYRM
Ru3OtimrD+9ILnySxdJ4EtnmYwJ6LAabjJerZpFF7Zws6ij9Ifusdd8zaW1mtX/0Xe+AzOPJUmVH
NLAW0DZU4VZmoRC/3TBDSdFeETc+OCQdjSfmM4yTpnjwFjQnGFyouPyWa5a9vTAqeNxB/UdLQpH/
NN+OnmuZqEQXKZewkX26MdVH9h7/EJpxAirK1UTEDQLd5cx0RkFdadw2/Y05ICiEp7LLqFu5qkqZ
FgmoFp3gxrfzbo6VNWHKsOqEgEGB6F1bepMz3fZFKtDhLux+zmsxBZ5dlHDAl36BmQw4nJQA/DW3
95Xayb71mupxv+htDQ6oeGTPIORItdkq/TUpJ0PqEH4iQOYpNeIvycJRaqQw3Q1LmLqYkTbi4tZG
unX8Pv7AQEEl/cTETpjq7wtSh5NReroHnR2jmQHldKZEgbjPtdgzFU72eRcKEG+07ITgIHaR4Hsp
EW8Es7YEf86wQIHdmM+Uq9sPhm84OKmYhAiLd02H9CBDsgR4V8xs7e5hsjsRmuyUWUDSANM2hj8t
SycfcUCvLeTocOMJWrmLGVfx4YLENDO+/UMQxKuYZm3X1TvU2jDndQMuoYHskCbayJehxQhpfLnY
WfdokLwxw34fhzwHnUPkXqHcEeBYx6PtOvccPn3GiD7RmyWaxomH8XhrE6ihlcMBrdH80qaED99o
K5nEL18GZ8CtBLV8pCCaPGsN/nFwVUBx6tBmPJ18QtV5ttcfzJZSEE2jGwpIhLF+0+r8R8aHLY8K
3WOHVLgqnGjKqjhZV4e8v2g8ZihUhbWmNGYRG5/LWznjwcyxdY5t0sn0c0JHirOL5PBcJqt41Rwz
29buYHdVPYPvKHZbbvAMJSOT9gG71jIf0PlatZqLnarZceZtoTCdDWZwjaR9SbZIVgxY/Ql8Aqg/
C35TGZAOD1yax+vTEaH6mfjH8XITUd1RaeIoHeMRpDT3NBIyIVQwESsn3UFURdYlI9wOh1oHOZpV
X9J7CA7jmOonq/GPvL4oHiOj71x/QSw7Q4H8IE5ZT5c6nYEGhovv32p7x+a4nWr3fn6fAnKg9pZC
XH19Ulpala5MDLTZSSB50OVOP6XWZpZMSPKGhgxyaV56HrHRophSYDqWCALtqEZu6znNEar22IeA
ycjeAfT+13lIenhQVTckVbFC7N5NMxr/ryivEHqcVOFqIgDxbjQr+MwGK1W+D5x3UeKycphLgTeK
xOD5D7lm9nj6n9DVIXnLOLS7a7AKegqABDyZiDapX02quDxcva0TZ8aJ7nw7pspdpA3B13fEmfGC
iyh4uI/c8srwVj0DfdRi+QELnrbYLWENtGz84vmf5vsX2nIrmk5xIzV+TNVFZpYrU0Odcg+v433c
kjKOR+xVnHrpT3pobcRfxTTcUPen1FhBU9/sEk6gCwKq7CqfcEpxaQ4jWD7kVLKiq3Gkn64GK6e7
YlMtc6szR4VyJWjayoa8AkiIBHlNy/xVYspYtJ3LTFE4NJvPkLSABfuyfdE1/Ar8ObFKDRolzOj+
Sa+4UREoEXgyCvE/kSiNyICV+NoHXl568Y0UIJ3oTq7Su/y2Vf08Quoc3HLAe1HX9RNE3VvdWvEn
U+cRHbTNJYRdqMEDeRTcut870huvDiENKeOchtly+ia2eVAwZDGqJUvj+VqiNLyCuEfjEY5+EpWP
I87uJiskfvBxgQsTykfAVAuTTxWNsG/cRIoveweOpPM3Vckyf4Dkzq9h4g82cAiIatPNQCpDk3uR
vnm/HaxxOu9ZZrJmU+Jl9F974T6NkPqLmiUxBn4umwfrRFTYHvOmEftRhrMOqRNKpnQqu6zWKH48
+CW3VEhd9krgSonmiX09g9v5FOeTGar0rH+2FtwIgad/P5YuAI0FfqN0g+oEybcee3GjR/qLK+BZ
ju2eQ7gkiKXPJgZllRo1c2qBi/5/Y+UW4Ah8OgZiVhTcoHSZ7RwSkJOtN3hobxVn0yJviPXLq2ze
fv55Djegjrqbni2YMVRMIlh1lxshXD9gCF8hpsS7pkvZaPvrfg/H15gTZ9LJbNVizOmqk9SZJFXi
KFWt2/jxjx8s9tdMbg8ikt2qJ4LloWLTxSgaG9lpD02naP6linrVXXVc5a1NGatTvVdWd+O+2U3m
krmd1uDhoiAPEqxHX7hBCxrDYZY9zcIVJHcAD9L8Y0Dge8zqCatOhDvN4he8bLuv9hBN/1BVNpBh
1LiSIuq3RKyvu9AQ4HHUcnNcUn4fAKlV6KIlNeLHJb5Tl+RVpbvgslpwWyk8xa871aDxcaJr82mf
lRY8NiN0ArJd18JplZmtmTHlfvnqTDxf5/X34htq8MnxP798irbbnm9f7HPjdUie1awBvUBe0PVK
RcQ0sXqC31bIEPIkCIOYQ6rFlsgfP3x+CiajOxBQdGFppM/S5lqNuWVYQ89lO9P/zrhsWmpeovSj
OBOWe8Ia5vRCoJitFaUgX6MTc0NocYqoTDKR3hAlnx6fCf0HVam0wjqVcfWlOOJjNIHvIcNWEJBn
VuBsHB6UYodLoda5iY9mIxD6ggmOaOWnjpMUadEBkoo8n0iualVyLjsz4/c3LAwM9VBx2f5oCqLG
/+6sU8v12nrVIijEeMa2k61tux4o8xkmk0Jdy6QpCbINsqSyvQt3kTi4V7vp0rHnztE5Ihiv4PV+
Yf8i97ZGe0rP7IaJioXiBg7tJLjw0H7hed3cCHkbl1pApoKL7eDtVgB516LICeqb3FIuHUGPkTHF
ln58DEytMHg5Z4ev0+CAMWyxyeGUgdf6nCG+zcDY3bxNYu/oM1lf8lbNL/Z71So0QAday7OSxv1I
Fkt+G49AJ9OVL91QAzm71puzzIArNKlocRzUlADj1JgtUAHP1vSc2AZF2E/KuCs4LYRznPwE66No
V9Neqdx1hAYX3MOIOpdb4oRuVbqGQ3rpnWqUFuknb9g8Qygp1crEl40Kn12nG/TnILJ1AlOIx6Wl
mDofDI2x8NrhomaKIxouK9zgSokKY4dFrfEw54KHZvvcAlZzw2WK5TrZrRSvZaRsMN6gdyBu0oP6
1/yRX8WKl43gP7KUrmwudinAl5PkWcFSsHPig/WJi2l4IkX+dEJg2RpSgiCX+rm0zk+CRX89n20/
xgDkzLzTczVtWZFSSyO5ResetCknJlTyhXPqJMtTRwWdTvDY+FuxaK0eBJ/ytm8cunmYwnCBtkzF
i681yyablOAHZ9rha9wZchWi72+EQHCHqWMk0GqR/Sn14DhkkgjdZzA9J9nGb4xBykVOmwBxgYj5
my43Bh5K9B2+ayhV8wOxBTqHQ2Y5SrWKu811C0uouGMxPkPWrXTMMV6e5VIjMH//7AX8uV7irHvA
kfmcETEzFvzZu/6xrThQfV3qREa96w31bm04yaNVg7tNE9eWnCmg6F3ZvfWADtXJKC8sVCIuQNDN
4BEyPk0Lbb4SgOXttLOQLUiQEtBSmskuG08+o8jWZjZNiQCp7drAPqtcPalkDOtJtvEzNYTpP0Q2
KWKzGoXoRsFliEiZotvEugdABzAS+aR15UnX64ocnhPbqnFNcT9nWo5qs2AhWnXFBkG05xHFiwxf
vboUu5Lhebz2F6L/eCzohiOYBWrCtbpTDqGQZPDN8tcNTPM2Kv7M56jC++4lIEwljFu6hKapnDM2
USzYCz0IJCbGsE3eT0FgMmiH82L7RlMyP8pOLJqjSGNe5ez4LVZA4absRpMcWjX3ZAuKjcDbCEgH
JRAYshfMpadzx88oveYtx+E0iT6gS6Xr+jT2BEouDALpxhT+HDzSSyOhVKlZkAjypcESunCWyPCn
oP8hpkeW35IdqZK4Fy4qJ2cKqNZgC6K9ZxUcyARpRmSVir65R6QECtP5QOwKristFhwkqtl5VOIY
A3Mg9o1+piRxTPRu0bIFuzbTSjCuY7LEh4VrRlnII7uwpxWID67flczEmipr6yJNvX+ltOuhI3C2
E1x5+lTOxeqkQXBY9+Pinpgm/saDSJndaUB09AbSGYp6gMLSqZy8lHfZio/xn5WZVgQzpdAMNY8z
xv/3ik3TA+GzmJz+Km0fz6rnO1h6WNYHQE2ifMzSbWx/JmMe07cMcevjEPN1WSMeRqgKITD1XW1o
s8h2XxqaPNeZ+r5+ckSzZzqBWta8qHC/T1NhTFmj0jRok78FQxqmm3elPmk/NcHe7ecLF5/CdlgM
jNJA6x0aJftte/KKQCa79unovajqLEPngwFwZDxNLD2REXWjCQeY1ckiHlRz0IwgStjQFe+wJ89A
63j6gyFXsOFdQgvY5X+eFGSDM2Ry8gQjPAVhuW1rfbA8Ys0O+ezi+uV5CTcSVF0xjWSGW5dmW6z1
CUfUxmewW5BvATkaPyrnllUcxWuGhpbqYeWcmmqFOUznVqDST6JSE6PEKIotvJmDSKlmqucAvv66
TGYDF22gaX7kCB0Bpp70DnDOZgjtFYhbPvDLrcuFBbhwd8yRexVQAxTbn7uA0II6W956M4VGf0wx
Y1gy/V7wjo/ZxS7LOiJKzEfa+s4azEyge31MqtHBpPyhL50oTRUZPKTDYR5Nfg9sBYIUEebS0xb/
yjk6yx0lP7ER5wesosYkIWVaLa5uHVtn1oCS7SNtYvYNChdJICOqZQAI/ZItMFXJP83/cbNRvWbU
cuRm7BlvwEkag+wm2ID/fhWKipmJU1EZ9KPfpP0BWZZlEKNxCYP3mB62ht0TmaczOhiJ9Tu3Oc+E
2jviD+1lN6EoeeoCDiXOcvGt0HAWRd/bI1TkcXtvJrJQPT0VrDC2bFlNhxHuu6nZUg4++9xf/ur+
21S94CYyY4K03OhOv8FJCwbJn1T0pAbHDWSK+wD1W/z+qgpOOYh5gd+VbJBAh2j8RSRc2UwTLLNE
6aFGQTOi8SOWQHG37n9S9jy6+VCs4wYrDJtxyZct2ygAakNnB+z0OkHXHurcTWNQZEPChkfOynLC
xLNKNx2VX5mGXLjMEvTDRnLg0ODFZE25GSSs0mI+NSPRfeLky2f5fD9nXWafxE2VilatvWuf2go+
Y+UzeiuypQVZ0j9A+FHBrPe3/corHo3TfjLtE6+FTXiaEqs50NXluHazUH7MBElLQmrG3GHkCPzl
8tlsQNEQDa0EXIIkvMSZUm2v3RyBlA1PuyaJQJyeUOnnK1OosWZ0DZjxh09e/0zyaPv6KJkKYU5P
VvsFTx7MbuvjKJP3HkS42QYIii79c2AvTTgFmp5f9Ytx5S6raiOjkq7EDuSK0SoE2LhQi2/Rliky
Nd2JnvyiYWGdWNzTg8NSdPOaRg35UuJgjaKXFKsFFGx0JyesO3q12sV4/j0XqwDJjFlcvx1T2a3A
4NgGQJmUMT5+zO0TM1qaxqOLaH4BLsoXXSHeO1PUYVG9ekl7oV2N0dRAY/havTuuv+V0pVii6HmR
+WF/KbAs+IipxG+LJvQeRxqLG3/VPmHKnkSuPdj1UufACP4ZvyOSYJ4YftZvui7/MG6gcfpLLgDH
5RUBinuCJwN03Evy/dYzuroNGtPj6PC8VktfPTUSpZe9Hc1DlapzOhY8s49cerQFsjUC7SrinDFo
WaxMLohVcsH9b/aJTFv/I42/m9E99kVrCDBbtGNB059/3IRfLFtB14BdLSFeQUyOCQ5VffzqKngE
Xg0TEEqjS7COjOUCtZkKtkTD0ATE8WbWZ8qhYL770fHpGt8K8V+wUkBHVU2iNbTvFgiIHMtLashY
k0Xc/Xgx5EIYAZNECnWkvHf1j/BqkjEtYaj/X/quV5u7yBXyL7qI6PJ0yD20qOSQcElRtrI/wA6N
+9ONeCdH7rnAItQyJE+MSN0vs82/rQmUDd1Yp4h4OAo0Z1nQK1Lda7YrGcptoHpYzwlFw0xywBBB
QpfmVz/la0GgHvwF3iBNZarppHQH0NXPJeL0fvPB0k/R4L5SmUtBG1Bdcm7iO9ztSnV7KfNQaY6B
3xR/GhKC3zYx/0/NaT0BhaOEliBQOjb1VwW+alNV9r7PQDLY/lEt+RR5ZFkQlc8Fob/mPIrw+oR2
KO/rblWwnM+UmhAKu1tDtGO6J4vl37ojE2eWk4SjXG397I/sdHPcdiMaVc/PHvyJKvyTIu8QtZ3E
P4C34t2c/Y2I/KepZLGoisv4AlYpUo7mjA3uqZIjh4JSjzAhLrYHUePx6yIdM42NO8MYFDBYxKIp
X6NbFDp57Yz1DHJ9hg3fiLaLgBWTn/qiz7DOtCEhbduzbiR5O4DpK8A+zHv6Uj+k0/lHtIuWzw/W
hWuN6/TDM5Bho/j8/bP+NUTqo7l1FwaJJxrVjIirm2MbDBO/MWXLWs0oF3JSLu3IUmbe6mTq07l7
taysLW2sbxVuNurw7b6Pp5Ed097znVeQE4DIz8Kc6O5dlDTWw1prgubzMa93IhaB8x6v0jmi+oRs
MqYACl9k/npV0uHzRTluXSAou71Y1VHfCEDdz5lPkbeo5p/M5Vfn4hqa3QGBGSlhK+2Wgz//zBRi
vM7+1LysD3nGK1EGkhVJzlbwSreyA7P5jlYSQJX2E2FDOLACy8Xt+H+Lf3zSGrJJYJ7b5zaKSal+
Na6EVoxr+nqypjkuBHEX2n4OqwVi3IUEddi5A2prYAIItk6bWMZUmE6pPYFXoP6n6szl3B46YZ9+
ih1EgIxZ1nZQoDkmX/Qfxn1pqKbktu/HaCru1Vfxeq6amJ7hBgnRStaiOFRwn5jLq0U8M2/fuY2l
vGM73srSpcI9hK3xpIgQKyxKnubV1bhTTjAPSvpdrsDCIZzNZNI16K/3WzTcsn7SJMMFeW/3xMr4
NpLu3QtbKN7pdpaMHTwfntY/ZdUYwGXqQ7Ox20EH0jgmruGo36rvslUbybQJCrOPdj5t3n5b9tpf
bcBhkZuL0GxZL9Gobs1fUnbTzKjOfzUiWvpM3BZFW+nYxUSXBwK+AyydhUYonQudXxVR8HGHwn9b
aKVYGgVA85jieWtRjg3bSi1aoeKZAyx0Igyb/1fLJ1v4D6aofVHzcq6Ck8UbU4y2F9QfaR3Gf5RZ
s8ZR7xFAlJ3KBCEIRNyrV2kynRrb8USKpoJgeKvIu7ACDULvSzcj51UbQOKvXqM9hS4rtlUkY8BQ
uuwCwTze3t9cnu1I7OFhwxt7CouLPW/RGRSq3KmySm4FnWu2M6xO+15InvtsvR2NQ3FIqWkaEVg9
+aRYwQVRYZNotzF0rlpEcEsb7XTFDLxYd0VvYjolieN37hdBV/QLinU5QP5g6qa6TJuapiK89t5O
6lsWRFrEPTVFt7vDoKubeatt/zM+yZyRjuBo8X8F/iGFXwecNg7Gg7/6EroaGmm3OaJh6lCsj8VO
SD2gNd2DkvhcR0oYsgjXLFZpU9I2qgva1mFhKpC8JNBtr3sQo92KTkc0YEqiUYGvLfx2iGJ7SvNt
llTc0WDBK66jSmSk2V+iT/S0BPJOcaFjnWSw1nG8Abnr7ZfaFKeh5LSl+bbKVxXySkmJoBxQ6E9W
mQnArHYTXY9aJfGh6Vm/Wi+3TPXbnBg9g61UbQjR4x4R7gDDHiitbtCNKiylG9Cnr/CPPIM1iGIV
Jhd+LWwKaAnPx7+VxWIiDsiICxI/OrhvoBdM8qzMnMb+yeCAIKPqoUXuPZ2GxHDxUEFndjkwDCqJ
duT3WbtLqMAjdalFCUXDb/SRKwK8Vx7lY+juGkI+ioZI+J5vqF7N5+O1qNe8niIX/+QElt28a/4H
J0jtsdB6n/pRywGHPvRYG5qXT4B9FvTYZtgJSKFGgEblhOwHJS+edU2DipIsncI4HwYmw+FnIAK0
93FcFu74Rt0giCS3d8GJA0xnMjGDpPOf6AQFpJL+xTrad5aGUimHOigMESzMzXhYMKigOUI+uIil
tmRQj2yL80FPH8NBB5Gz3GGGP4qMZ578MaiCAwCq9m5gLCm0pBkl2y3wPtCnVqh9nZvYPOkkiZri
i3xZAE3co5242RHLyB+4QFC96gyklz0n2MM0ZTvxFJJuyXgWFtk6AkpNF2p3T/BeiXsgHEVXdqt3
SYki6ahxww14It7ZtO6vp/jDqnv/O2E+FpEhTTwi/tLcxQAcHRGgic9fd2WYXe32AEBk25Io770I
/2vKp8Ts7959Ezv7E59SjCGAVDPJ6VguV5Jepim8IcvuNIE8FGhPLZsJJBzH4e4LBfiLvbw5dxN3
PwgLguKF3nq0nK8qwqpgg/8ahZ5hpjBhbfem3Bw6PggUTE5Ftw4nSVDwKIsfk/Y3cHKk9g28vTzs
h1fqzS1Y+tW0VpOTtYSpt5w8s6CYbiysrHNq7lt40Akm3TdseQV8QZ8Sgol9C9fY32PLtE01oB4F
iFHU78lVov+vFLyqNwsDol5jcnfGzfG34OhYIvP1EZxWYJA0HxBjh4O9P9bW8Gh4fiwhSHpG+j3f
STzFYnZ+ODeLLbNk1Dg4un+lLh+/IH1uFG1yOUS5rRFQ+syGdkgBHEwJbOFMflUNqbfN2OfH1jw9
YeTx8C4EhWey4BWAjqzvtk0oCSRMena5ChLWGjI9w2K6vGtxaAVVrKtUl/kyH/+4Ywogq+x9UIHQ
O+pNmpW/qjmE1Dn6DNHIOApvtUZmm7HQBuL9i+MfiZGtux3A0P5qIYzdBQpRXnKeGHB+hM0DzCPz
Q2D5eSLTctxNw782TuZ31W/njENbb+OEWXUUIbWSarwcd8ePQDrHlmiCAbMuOtMYk5IRE7unfJ3R
iKz4ntbIOKElRuMTCo0Pfu2D596B0xksjcfQBDZ4ltVT/0YuZ15fac4x9MvT421wJV3vk/SOOrF/
2BBKhHks27hentE0clHwrfxWc3lyYtsop8jrdcA1MUMZTEa+VZD3viBweTPd2tlWH4X1mbsVc0Us
A8L4zVPUVZEYG9gw1LpzFXHzjWzZqU9ozAX2jnj9mvUaCf8F6OT5ahYNz2iXoQlzMsFGvneL/NTa
mXvN7nAcBGZ0+ZK7d+nBmJN5bQdQUcJBKcYUx/Txy2mPCOWY1LOrMqHKbqcf8B6cG59PIWTBcOV4
hSsM5S19OPMxKoy/zSWlTH5J5FCDrsH+XeijDJ/WWc02WMlZsAFqMrf+ok6/qeEXzBZbAZQZb+VM
M+6P0PDRV4ECGwZJH7TFmYfb0jHxJRr+CQ8g2I6FUQDibduqNz7INHBg6/6JlPRh3tIZ85Ug2zXq
dJvoZippBkj7nTZyz13FLvjqCYjlMIvoNEqic1Ugm2rQYMyQ33kHK+k7zDWW4/X9/tdEIiALfJPR
StAvtsNY9tf2pTNQtb7u2BvWbWfP6Dut2uCBsVo3MTFyuu8zPgohqF2jl301iLPAgfIA5u2Fz+Bd
GvVhJaRO9rVej4SA2P93pu90SSHyLMxX51zyliMpfxE4/Q3LE16zFuYQEeDOS0xX4q+HXdh1ya8E
wQcLUVDo3WKTBgvJ+MmX6ipii/akIjffdEkqQnftzPswjz4zLFINTIYra+adD3jukSdoDiAOz9ZF
MK0VhDEKmMPJJYF63c9g66qavcwYXur9Ogcpp16nqXyvwfgKXgzOO4gzyu8nQoBjVV8AcGQVUoXY
+RawxibKkGBQ5VknHIOi2RxHQoIRlZR82DtYrKhU8RWGwW/O/xI8Q9P24HgUmZD1b2qfSqXEJDly
MJIxT8EATArNnoZO9Agscwg3PSjwdepNKRmX+FnnpmTp588804YQ/LIUzRRGHJ1fMXBRiDH346w7
URptV82qZoTJK8HSTpOkhPdQPT1XCesiaX7e/MFDc+YlFb1Mntl4H7SbvECLTOxbL0RrKXxZ8ZWY
2ZAW0EuysxTASk74wnb5TQF1N3kFwSqJhp7trJ2OVsfS5roAR09dWbuh1kZQ31/UdmMUOlzcxqeT
8r/wlhZILhC6g3d0NX7j36HhGceojFN+/7GU2A69MLD8kNkkfwAO16fWu5l4VEDthGUuiey8p3ku
L9TM/Zaq6Mpgk7qTksFhUe/9vQmD0IJ5agocgiyj3eUOE904SPO74yz/ns0/nWYwOzc66AZsDLWS
2uy8R4SHMHqHDaXVEr44q++l+YIuhhkPWfQCWrGuj2TdZehDLLidDBc6oWc58Z2wq0e67BFXepiO
lasvxXGrtqmUEKOPq7rQ64dVTmLql/YF7ogs30jdPYvJ/FVl7zuwped0bhC7Skz/uCJLcQMvjxp+
JTERTfaXDD56xbw9kek5bYY5/2S/s7UegWvq9Xxf0gnLGcJDPjcsrMGkcabYqWcXIJctIZHT/6+G
2UpWQqJ9otK0kZKfkV9wuPngOPvocBRo73hVU1E3C6Nys3G8Hg6c2fiGNYc7TZQawbbiyt73as/N
DsYTlFNQbhr2qCn2RFQ1PoEasKjaAvRA3BwuMbIv0C+dlF1UeCowMLzi0HxT8zpP1JsLXwZ7AbmW
0sLR89IcMxZCASCW9Rh53jUXTy/bidb6Zk/dBHskd9CcOfRa7k4RsURfZulAFasNcmQwOTPrrVl2
R9+LvsT61Gd33XOl5gxpLQJiGw95BWgaJZG0AOqoqFJvo4TAHdwRErKwBrYkffawLHq/pwA1qAH9
K+YtPoxDK93uCpZEUuMCPbRpiz3ajuR1faJ1bHGjlB4vjFPNE29P2agqof+N6kNz1He+G0FHrFCF
dy7Ps9Rd2m+mU1PjGqIq0RlN3/fPYPZF8+n/mBE2JcoeB0X+Pli0xORBhm5tGQgchLt11KAzwHfc
ME4502apu5B4GG1HEkDCwBTli8CA5yIhXurVmBULeCNyhk+uoAk9A2tYCweWNGWPxYl9quQgTTaZ
Ohjtfx4+LG1/moK0aOuTwFLaiu+PoLgavt4/Dk7K5VGbqyp5+5ww/DrGarZpJFrhBk24kdmp2Q+L
RjE+DLQZP1x197BqzEx9FJTBGx+vPGRcR0x7RE8OYbrAADmlcAyV7NclqiZ89XM8jKG8xG8Jti4u
TXttCovbOvpp0g7u+JeV1G45QefAtWZGc1JOU5U9n3yehTIaRPcPkrB63KPqUOQE5xCMbtr+buEh
+qn0FSEZ6bx6YHnxgt3d22V7vDmFAvvZEdR1VFJHkzGC21whesmiHWgmFC39mw7RZO7ig0IrntCS
LbG4l5OjQdM3Ct5GO1Sb2Ik4XFa7dKKSbiJ0B9VVYgy3flOaIXtJ4CdjESUoHlL0/9DRj3ZbFraI
Lv26lsHtI+I/1KfwDoB3RXVNH+OewNp2nZl6e3zpA890e7FIKhpGY5IV0M+SzKTL+OotDdCBAUDW
Ki9fMw5rFOEp/xUIg75X8VauPUY72FWxAt4RA1shbMHn4p+BrMorcgE3zOc2AJH+QJwgLBluS6Bc
6Nyx218/mr2Fno5swqboGm8HVjCFFYinWinzDq8jlmSxytQzuTnJpbAnxOzVeBecvY8+Sg7adkdh
IgEnyxAoYEmabMjWo2t22STENki+RW55jcKrcHvRbUuE7MHKV61kXSo5DKgedjlY4YhHgG9QgCiT
FfSk0I5NIgDRJmFNACS1d1Gw0xvwLSGGtYDxlF+s7DNW+bZXro5zYANKuLG86B4KATV/GA2yS7UC
zp+hTdSTK1g2nQ7toOulGMHplwd/qf93bdGda8UGSHHq+Zv8R42e5UrpU4txIaSapFAeXU7nHwcc
vQ0yiJ+b7o6zOAB+PBdh5iHb/UtAlpzXGxiZe6G/QevLx6dLw5rzRsvkETR3ffqtN+r9SQaozmbB
iwtTU5bszlTVoPq6OKg1LBeG8Uo+PBcWWRMTK7SZQzoFSiVT15/1ylXmtYIKprNt4m2A47JcJFGK
zil54IOqYpGcRAhkvJte5RjSAR53KRLWSm/LFXyGOrW/iR+E8Oa8UJiZBgxT+HyqCTLt1xZZinM5
ZPpkbkKhiz1ULGi7FX68Y2GdXZz0Ny/Xso7KKkPWVWmIKmayjGESbPp15ZWU4+Z2JeUBPHdQioAF
w0eCLJcL/TfYAc/ABW1hxOCXLrqLT65cX5OmYNtp4XIkS+3pY3qUDdoBI4OS01eCxHpawYfHZp5t
VF7vG8QUBBU4H+2aTR0OrKCvsdFc1uM1n2XE6m3gD0xohOAEc3tGdBOlhJmpLFaUANfd6c/xfjQJ
2Js7cmeOWWZkc3ZacHK7uk7SSpDZi3DDi2faKnvxn+Gg42SbsJA67xCWc9glDjnJXZ+/szwtHRYB
q08TDuKwyIyMD8BDGLdmfYtVeh0E4dyiCXtwEwBiiPxgMM8Ki4HgpVD/alMDx4O+D27ycFP5IBoA
Ms1w1YJtgpk60z4uGnS8t93QtztpeFVOYl6JegK2IRUqwLuIMte3BZZEpWFduBAT7tEfIvSXAeUc
0dlKvSnwhb6jiPbqUWRrbj3tNDnS7qXWC2XBMj7ixArWvuXlKGUDzSOPFO/7OSBwFRKqQIOBUYX5
RDHrb0RhNxbwgTVTrXvyVg/xbDkLIXI7hIGOlFZK/hnZMUBp5nHwMeLiSMtWLLf5wb+bkMP22xR5
lbb5bPEfZZBO8958Qj2s4jZwpxAlolsVbakg2vRLnH+Ym7fZcpLmIGMqrEvh8ne1+3tC4BITdvyK
D/t+5qg6sBYT/KfkgA24fK8/fC8uVvPjHYfHsLEPkSHVsjF4rlw4cA3f5GdzS+Fjtoas3y0P3sYw
CvUrggjMfSdQOfh92pOZAN125FuhW9+FjeTh9W0NYMyiqgZGHkz6TT/qqk4NKMVgbGrryhT2IwGi
BmcYRf0019CSOcc7RmSI1BhMPzZxJ8+3bJkvL38S/L9puVKKnSpTh/XKaNTb2A9Sby9rzhna7jmR
iDbvQ3JZWBOgmZOefz7FFh4pF9dvv8jzWY7WZ0cyZCxvwGoNu24w4W0L7hS2CU7WJ9N1Uuw375IN
0l6yjOI6Qu2jxittHvZT6UdAesPmgr6lbKylYI26N1buANfRPntoG+WqfS+yagVyGJckcfbh91AZ
gNYULWblaQB9ypbnEszhSiskFz322bW7eSWLBhg0Yu5A+AXLPvZv6a11afV/7sJT/RDE7Kg5M4bI
fobJfbnhGmrc6kakgtWPX79U9+lMlU0MOaPyl1xRxEkP8UmaLog42YYF/+Pxi+giv070CO9lf3BD
TAutWRL5j2MrgWVfwTBHu0Wv36QKlpusHfPwLzPYrNqTtQUsEKliYI+rbGEgHVNWmSXU/NLz1Myh
ZVrpJRp3E5NUN31ZOlNjAYZ8vYfKj2wEm9aDxm0+YqpjgeztCvJaNhJ0CcGv9FgiMwteKFp7HfDa
2PJ9k7dHirb5IVEjKQ7CAqggxxQhRa1hzHQn1YASeOQBq5y4PWjSlOLaE0p8ndCbFbJNn5FwZ5ji
lf2nHzRPPeFhibjHrjfpt4D+JFab8KuSYcpQj+DeyjAiazFq5cVYMIPWI/kTNsWlVCKhvV2JnVG7
CMBffcZAPZovhSoy2OE9nLkrzpObv+uJFuEIPKeKymH2NujhGYnTNstsejaSgbWhzIoGf8IgvuxT
xg8M4o/7FdsGnOZgxh6s4d5JIDedj5o+XA6FD600JxHkFsjpg0zJY8LjeoqEP8hwxywWjCT1ZOdn
hAVj/YFFx/EKJO8SlaZ4E3tEk0oHnaoQU/lGdw/tqA8BHY3iepkI7A/DvoDZBnxbegogIunRJ6yC
AzkW/hLMwXgXV1KvN0Xf0Koerx1Qrm+bG+L5F1ZbaNL1XMDHtWuxBS0/HGO4GVuzPkD7bwUPCXzX
6DSzjtEXGpeNYNG4x+kMF2KU7AfOjayv4xUvXN4Ccv5x8ppcOyM+dXrNLIPGuUWUzLd1ZcVPHNX6
ao3ocXiSJkFFWW1gF+1uc2qHBnyDvvmAyCAIsIxJJWMczrwA8B2ht6fO7r1nzyiK1fYNCtWgRa1r
e7mIHBUoEzfHrL/8lUVMFSSgjO81KyeGX3/cSQ1+AeutMViiqYGftW+ryh4Gi12WkWmvV5IEVcW2
eN4/rH/H2k1ePwZVFLGZwwg4Ug0mnuTAc+Wj4GBwsBafq19iyO9plhXTGDg/572cILp0LGYu51zC
vSw8buHnnEQrC4rVBF3mwU1Lsp4gWuvlJuJ8GJ0SImudIZCi8MI55CKceraWg1WSoyulq5U7yuUw
nOjsXii3Vq8Lg/Px87Zz6bA5N7sWgaFlXcuUvJX7T9LWgzy3d72fikT70kEW1FNx/npnuPTTfUV6
2Wf7fslfC2v09PMl4wSzbwEHZbgqbt5yh5z+/KD+ijF+LCR+dDzp5+UyUwH5Zkuoy2I8DHwELUge
iJvUd7I2K/JK1kxtwg9WrvZKbSCqaVBO5GH3wjdfad73SKzadVmJz+MLY6bHTODxUYH4w0Pzu0EL
O69mhhXt6i5xAc41pz18Sf5GXm8CRMTarbu/wghUiBuv1k2WMyTBweLys4AqSGdOBPBu103QmYTM
JKdXly2dks+iy6tqwQ9LoxdtjX0CyNh7Qk6fK6STOvuKLJ9is8VyCqQiZRqY6ZbCFTLWIvJbqn+y
3zVE95EH9UXooVL6aRkZeyFDWHkNX4dXGQ3oIMynpN5P28YNp5d4K9Q4kaEi2BBk1450shX0HV4o
rW0eWVLnRfR+HW2RIwSxCAuxuY40d5M5aafIQiCsE6jvYx2VPwsqy8XG+iBnuErN7gdAdMA468gE
u/y1XW9BiyaZN+6VXRB64CpuLk9LjlPUYi/fdKASFk2eMhBPjmE/SLEinWCq6csqtvExAIm4NOpG
KYe13P/2HvpovnQTfJPinZWcwY7MObMZhDrReaTOlefDWYofZthCIxEwYX6JoC1Ke8UpHdB4KY8p
39LPpF1AhRexGO7PglCy+yc0fNZvgA1wkIV6LORFByP9N0Gnb2RPG58e/8sZ+o6tK4qI3oTFQ9Gt
dpu4QRwhH1ZyOzTU4/29lXFfb9QnTp/xjolgHQuafkBNdZ+zZqDuDVQfhy4Bpc7iTATeiAQ16Ju3
q/gMXVt+D4VsgZHK5tS8AgrYtN+sFExt1tfKcTlqmdSs8GytUqlNRYT60ZQ8vjlsPy9x1BaUgmzf
k9XRDXCy8vXjd8wKnN3PpBQ+m3u3yMBkIBV3RUnjWt/HqCsuLNrO4r08wvgWPrqZ1uR82lbkKAK1
14kbS3i60BJcvKxY5p/TijTMHLGBwHAD0bJX82JQoixktvpba0ly8M0VsssPJR4AElJgxpLg06Jl
q7Qp9Kc3rZ1gZCp2NqTAvWI9FJMHOn3M4mrrqI21ZlHxm/SynccDiyJNXPP5XST2evnCc/b7K/E2
Z0rgXpPSC6vVnm+2kZ/hGBWhTnnlkIMNJjTzClQRvucUjLLbfJIi1vGSNucHeMC7SpTS3RnSYg1F
+AY3j5Bm19d20x4ZykARHb2XKWXoHfitWlw0uOeLURdJIhdYk/zH40epq99NCXCEjKZng6Vcnu4+
5xkWEcYDwZwhL03OysZkdxOH7odAV1JWb9cZ+bxu5g3KfsoY48jiYj5BXWA63WUl4b3XlhEDWDIB
lts1bVyjUG9iJPZDF+aYujOwQdGF4kBX4L+w9lK3fiYDr7UrxlZptlONVHH8h5stxXX6iY0X8zCr
wRVcFXQOlZuEsh0M4jMlqKZr/yTxG18w1EhvEf+8MlQRAcXJwss9fU195HDsFXqxkAZ1BMPbHV3l
Pze5uhSBEKeZUnTvLVEfbqx1ZOpfyP8g6dvVgpCB316glp5Bk/ttYbUm3VXqiE+GzIBn+4xRDcDG
f80ztS5LMZ2PMAKmNEuoxRyxx6ngKUELxBV9H391Bzd8ukQP9wrTYswfgKKrISadeCcQYamuS1HM
CCrCFOrKCSV2DfDB0xAm3WXyoReAmhw5+wZZGvQHgVqJnrfbi6ks9JC1481D2A40bw9iTbgIAuoX
X4s2LiVY9nJBceAmChpAMMNLAiNeMN4xmlxzL3dp/YOISiyysc4GvhrS/88+onAZYznebCqaHNbi
A2PD87lVe13wcfWWs7jZg+CKRSSSMtHsHO9uE2a96myUmMWIhYImEnisrQWVSWr9EOvi4+1lNkI0
yTUHl1qUJBQD6k8fTSugL6hgSRykhqpoR1dQslZkreZX3c2kkrHFFMl7aCjOpzr1AQmGYvlSqK99
WNg3/Ir8e96++vzYqE6J/+BcnD5g6yXS86JD+149Of6xDXGqyNuQYSHTZ8U4GwPN9EH3FLJlLwIH
JjhiNBjJ5Da0HdzQsICuYPsPz8SxgkLEOCeLI77W23GHud+oCb2bmKlO0JitIFZge/p+2ScbTj8k
x2AXPLPAcupHIh5GTCEyVZCRUXH+wx287Swj3CuRPEDH5+Y7e/6OcWNg6X8xpTQSf1D58/at3qC7
mzYcCQRS4nDdq3XC2XRFSjz/7QV4en73u7NrsgYKy3aT9zX5iw5iREHl3cGb4sOmaUQ+Og30oa8h
MQbKWDUmkGw0SI79jQfjm3GS0syB8oDnJBhLCkZzt1eYRGkya6iwnOfflK3uQKyijFTH7oeSSYwP
nLcFqpwTReGbvyIbpIdvV1siP1KcJg2ujcsi2joB/ZskpS/V13K4ZeQ/o1HTijxrWvANHyL4Jc+4
DO0L29OErQyVKektaI/l3NAPQbjWjPIfxrFblTKFwHU3V2qoJ/vY6xz/tViernROkzMQf7nLn/Uc
i9O7dnB/9M95wP2ga8tWPeyCah8zE11k/ELjIR6m9exhHZqlwDaZjx6+fSQhMVAVEC8y0bD69dyE
1Z6cJEdoTlLtsWE0gO37bR+rffrGY/8zQWqd9ZfafJfk/pLX5shMFibMsDOloXD5ewaFUKTfkbNd
d0aLFSkzYgIR+J3MvIWYMZ9GTZH8Ps17h2WSwsYFOg5ZCEMznJw6jfX4PSRtsmOn/aJj5wlI9xKO
TYfBQVzkHvmQpR/DCkWyRcKeg5uFDmFyPqbDd9HSpFFM5epuVBv9+57B+TRL7wGLFRUGkwO1zfQe
Xe7PzGm1D/vAT5BRoo2QlXaFCIslvhLGRECnl7z1otWmLPdMzT+c1/S2c6xS0Hnxfb0a+GdGVfb0
engbXFzQWOxUdreUzqzbMdmv4v63dtiZZwOlzvQ0yxC15JjKIqim4Tgqjs+k0xJz1izHWmWftmvD
5EaqzH+4DOvpn1fWET/aIvuxD1gy8MiZGyUk4gUfWkXc3vKTvCbVYkKQb94k6KpiJtVtDUBKm+I2
l2TD4QImMqBGeiyb918PqB1Ebw1OP0oHo0OqX5wJGjbshAFlbGKE5hXnto/93t/mj0dc8Wyf5cFp
qlv/3SB2nuc5oegecyTqKEeaPR1FqNkS2C1PK1Lp864sk3eFPyDOUTVr62PzYyfnX9O43O+oocf0
pRfhhIc4a0xM5j+lG1H9IpuM1f9qX4LokoylBky50k4rFObU3LtJX5qkL6iIkhB6m7qXo1UVgMOw
Rl4MObGQQX2VRfqGVrsntkIRF+5QYbKaJ8eirbPmYF7ffu6dBr3PvRYvXvEHL9DYdSpDi8KxFb3G
cUvUido9NcN9xnc2kWWGI3kTnzYFBjSQ9H1QKqPrgIvX92XAW/XceQAPDzEV7EDzQLf6d6vDDxMp
sXILIx9gEPHS/kDVN9xrx2T02CzAKFEDtNL6EAfZuAFn7G8tdQSGhMOtPgrrhmEX+eHD8FoHyTxd
4XRFCWYOUQVI99TXOGhNGHdSotOFCN9LdLKXXhLfYKXiYvJR+gyYvL+2xIYoQbhsfRI0561/A8Ni
C5D8/c06jmyNSijU8XwOSmYZOMX1PnHMHmZ+wD1JTcJtJ9sNTxK9jSpLQh25lq2opJGBfdxeQoaH
uTXC8HiDL7Ff5LhZhNizUETBruL7QJBGoMrZrtL/d6m1tNdhjKVSkXH1zw94AMw+sxiWMtXQ2Vsl
rBk/yu1xbGxwAt4stILhwMHKKO4ew8ba7zgECfWSykTsrvZ0YxXisFjiyWKDaBGpt0q/+vhCI+O1
U0MkTjj5LcjZw2ageHY173kvGd/gCss5Dzd/4I0uUX8HccTgvSyb8roPG/ktQgqpeesuAE84DPjD
n8e/hCL2zRAGJVG7tp6fOdOhr75aa7qPF14unizBWTdRUAwiopbjLSCabCqI4W4UrO+HfSBz3qqd
FP+rge0dUJtbNPgYKttQ9rAowjWpEc7/LnOj24byOURWPB7rn9PWVe9Z9Vm/Fo+k1m7ehylhePQD
mLIMVELVHM/2Bt2/JcGRcKNgstxnTC3ePVEkkuvgYrL1N+cXcsf5lSpvxWTS7ETYYeW0N43pKAxe
5qR1ePSBoAZCuRNp11BWcC/XGOvnHzGxordOj6VSPCnApk5wqxmHnkGbCaVqnhz+yGlDscS3Rxpn
7n8Qc34fdQYL8b2t1VMuL1YgLi2IAeHQ5Sb+NuA8aZ3xsRlZ8JBQawZLDuvObXcKDil6TKnIOboW
/wBsavPFs6jBHk9VrHg7PXwzeohdutjXi8cMg+BG7oTF4kf2ehk+lc8GgcVrAK0mXePuNrfWL3xX
rhQwycnNBT+beiJgDLJ/shgmsnulWYnSKC2ZiNTjwBcKsJ1h1AvREWLweDiYyAiF0OroNNJEtX55
0TYGWHCa7U2tnJhDZTp3hCbfBFDzPiH5roW2wVghS/nm8SyCiXU7mFwv4jtXwf6/H/FVAjI3Bnn8
ZPqcylNspw2ZsOx9McEy0CA90GOr7M7QDurkTdpxBTuVK1jQx3b5GsqusaeZB+yiOAhLl4xztTS+
W36w8HofloU0n2iFyUBqFHeJisTdAoxCCw+q0Ac5WHiD/89tTcxU+gii1eS3b0X3PL1yuFLlGTBI
0gYNuLVyC5J6cs9+p4a9qtViE9UeDpvDrKFacfNv3ozVMx+jRay9xyKvZr5rxy4bq2jzTdQO/CQ4
WsIUnmWBPRp5eXUqQHO91qTXeF2Y6ctYs7O/5fs1c7j8va8XSq5pgvZQsJPaJig5xy/KCVcBUJDb
7bGNzLNm23L0CPsNl+5Hbj9FK0ahEMb8s2wXsjLkJsw29m37zoTR750OfEDLSPoWi7F8x7cFdmmA
19CkgnGj4kqyGoPi5nLbV3/ok+RtX3QrhQ0JurjTf2EUz42kmdWlb+R5d4oT6O7BeD25APZkOBog
Jp+TxvWpC1cAU03itTO4o6CyE5OIJqTjrOVOqSmIvmJFKJcO2T0v9qSKdpNNarVfjnYOZqgno8oj
2fZIviIi99e4NL8MAi6exZD7SiIuYw/dA5EaD2SEbPuOKBfhrbS+umd+iE+ZAjnsJ25drNuamSjQ
noiF6W0RYLdPG6Ujgzc5C6VbBOh7NcUVD9ufep+LF9HKsbBnXccuhOs6rM7n1+DqFNzm1/xjcwH7
IPHUU+OfbwHo+pxUy1bSpCHWE3azMNVHGreYqHO68NsisPDW+wLkrrzhKgFj4Tx5B36lQfegm/fN
Xhw+1WptPmGqzX6czqL+JuMA8rLOqqZkhz90Ft5SEJeoTRi3fpQQwkQVvYjWnsgoST66q+gITylC
rLKKWbXmRDx4YIbDt9BOrS2wj93guEzleKqtrDjko8jWnyvfJOCz8lD/t22uorFCHp0Amgy94e6Z
7WzqEH8vM8xEGu1E3fU2MY2L48bDFps0OMls+bueAs04YN19043Xuf34fv1doiq1CpZvDq/FVBKP
j0E8VmeUcqNH99vuSUlQzI/LUnGlvlJU+YnaKcT77doE56LRbOB7W1G3Sha0mRACzro5TH86awhS
hNBd0zo35x18zzipXxAHvNgcXtASmmF7+uXwwHLt21iJfl0T0fLGb9P/zmVp7IHz9yPb76Dmto82
rHb+hIoOordyv3CD/1ObpgD6Z2uf2inXyCEVLUwKHwi0hgx5dakBa5P1qpaQqb2xDiP0DHsGrlht
u6/uYuzTL9EM3F278r1VSsw0YYy2BleH0avkzvlIGO8qe5nMYLGY9Yhu5Hto+WOts6Ixzwji0OjU
6I1ZtBWPSU5MTIghHS2r0fsCTTpZPdWY2Dkp6OrMwRPyyuFaSOvteuF7h49OXTCidstz6djZPcJa
RJJJsCy7DI5ypl6ezfZ5nOgtPqaN1bOe5FEXQxs6R8TM/KDfGsVYyThdXkwHx4KD/oCdaaSL4D6L
Gc9zegEaXUEZSTF+hA3H6DlxL+GU3+yGkneB8S6cIxwlREzbuM6KQiW2lGw5Pe3rYYOO1d2OYLO2
WU6lyGxH4KchJuAa/oEGXagPQav0B7Q4AbY0wQvk7DwMk4bgB3GfKvC95zfjj1KGFaTfoLAb/JE9
Ll4GQbs2sOIcPoNE/uoNUuekUQELJtUFJfHboVqSesk8EdRz70W/aezWFW9O10wPT/OUJQBZMj9O
ZKCW+50tW3TqU443EIZ6nj2QY68SgCq2EL8B8Dijbl/HDxpNd7m8o91jZh/TNdsN1e4Wer37fbRJ
c2ugoKDdH85RdcIL5NeS6mLo7C8Tg4rsceBQb+zb73m6u0EtJ6Y/P1dTXTXoSjjuPTgIG/7CQCCv
d8COdbcTuVy85QZHXmI2oDR40Dpl/wCZpQba+DBWDOYzHl0xRFHw3sxXPd18NS7yzew4YHdY02LT
jjRhORpYvb2IygzGFvR3TQ45Egr/3DgZ1kW1ZpN6p3u5vDZg5VzEeSoucLBMxFuUOdHwCAUg9GRp
xtpuBDfsrvkJa01mirNImaWwpp+n8UZyVcNiuzwEku4YmTgycpKgWYtQhJqwHkhGepkMKsFOdl13
DwxzzF9vbbt2dDXwqMqYIqnf13JYOU6P7qYJAwQWQtBC6LzSkf36c6xu+8+mnweM1CgqokEhC4t9
fmC/c6oZAtu0o1S0rTw3Ef0LcY6ThAXEkMulw9mA8HMyrwqEZdP9dbsU8CQ35xsDNpjGiqGmLMGC
mH3IBFqLojHRt4ZhtHR6W6JfzKPRSjoUzGFgGNrScSje+Mis5iwQCYy1WaKNxG/SbkYe+O9381KZ
64gC1qYcvCc3vxm1702+UiHvV58gQm8nwyHTgpskr48DHvs9d24vjWY4vOPTRYi3+NQ2fA+kDeL2
+H0z2HqtMwJ8M2A1Km0BrbhVZpTN1/7UoG6UKMNKYK1y7D7TsVAnvEh/xkVICleF7Y1dKBzeD3YM
uiNzvHesSJ8tGOUpAyKzEEK55G9+/duDjlBw/h6LE0nQQEmvHXoBowCg+us4ADukqlWOFS6Q96BU
+SEXNn0c6blBixvTgxshql4P0zzjBvxTusJAeKk5jpX9A7x0Fby5s1jlhP0Mny+Af7LvP0mkd+OS
y1XWyzVCTFBXfweupKVEnAaTYGqWHF4nqGDMwf11y+wZTk5X8Y2OoV+XwiG9f70wTV2wy7TV11HP
ZlvXpA8O6wF8aV2u9twByZCa/L0iVXOarUYNknavU9Z4is85g2K8SlYl9gSQ0aAl6L9A9QWIZ2TV
6PVfTFtNZ/xFtr/fmTVbi1gDA84GF1Bvs14P5+YRGiHz/d99YuPEzIMDY2qfjsSwYf1HzVJk0vew
dz9rEEBX6p1zDmlr3cYfE6BP+wWM9GF/2U37JAqiZSHhzJ6XL1Bi353m6x3w7lsQheCiqy/FUQsU
U7WLJLI1PY6iJzPromSfi+hBDhNST5WtdUXJPQPwJp0/vuzaWdcgiYelT2QrgulH9lCtim3sipcv
gbPeBC11jGZGhB4fg58gnhVWgoPVRvekZndidQelD4NiUCyLicBv2Od6sd4BRcwKi8EUNnnTfx6a
pUpZrkmhvB5K84j/Cj1tImm7zjNxzieFWS0KzPLBe8dDBFJKfGBS3GSIdtAr7QsP62sGZUBp1eAq
RjosFIitICgoKzLBiChXqxYTAN3Ck+nL4YIFJAeG76m+TMnWoYC0s07Wyp6xIcWSIMvDRUne4Ox5
Uj3RLhDccDOoPJODIlJYIvSBHUyPhSRLR+RwQZ3/wnFsoCb+ynRdjvds2hmXpRMVevmp1JjRppx6
xup1kuRjNkFqimhuO4N5enIysD0atFZSw/QUr22cJR0jWJwb9b3Zt767Wcgpu04eqOAjmLhwQWrb
vcud3KEsY1Mahb79zBAW/Bx17CBsbLDbcb4tNGv6UAqNPJ7Hh0XeOfun7NbU57h9ChSQ6G/5wnvt
Micsm+iFldEc2DvCifGN7Gimwh6imGr2fVSbFGFlQDekv45Unu9V2Yd3sArG1oq2Pkz3Dt+Qq20v
mfi3R1olM3a8oZi2kNdGaKQKPkhoTSvx0L95hwOEiCMoLinrIaZ689RPIaXuvzb1Ycqm+56HZQRp
FZlIhNCtu0LZZnwlMfkwLCCoicOb2njzaM66eFrL8VU866YBIvmMTBs8V/nOS/dZjDxrISJ8kyx9
eB7hmI6DQVPblO7J642sHRpY3Y6JNVuld+QR15lDzNyAAKj6utk0TM26sd5qSZWH0wZJDjKqw1Mm
HZQ8CiuAEueuObEV+UR2FrUGzgiLPPDln0YWdl2+Y3RnyHKs3am4roNKUR3fQiwHvOYQEgeDhR0F
Pq8D1vZ85F2LdNLUv7qTkI8dR4A3lo4TBbxkbFf+Iq7fnlPNmJflI96fYrTdpHmwRRNbHU33adir
flD/5CZXqayFE8HohWckLDTG+wC+DBeXj7V3/fGpFjavmtQyaiWpCOHiz8I9onm2uhDHuiKg/1XR
uvttdyJylfLTh8D0RMLbcxXwD4gWdlg8isRgCadHMPdhWkPjkRpDVqxfF3+7xs4cb198nJwGEdu/
rLfJaTQT+oJ9kmjD8jcwh7+47TpDDC5MeoVsN52SnwHprM0vCGULOsJX+QQjXrNhvRSz170piR98
Dk30aMOMtp/x15B/L1QLZ3ETeJSdRgGS/Zrqb7I02tqCNm3iOh/njYDsEN8iMZMxpzHUYCi71J2A
dyMZ+RuXBnd7Y0VcSPJ9whSNp8Nhl6qU0UpJ5FwGYjHZaEEtRioRQpleWmnj9DPEwa8LXRxzfE2d
iYECuOZsRobeM6C8KeWVR+uIEeeE5FQ01Ak7Pj3GYvAMjLVXD8hlsRe+Qkx/m+Jh61ObvTXIeO+d
Iu9cXJoVNn1xVpMNkIHH1Hu7/2feQ4u15msESGUXxemCxPAcl2DnohFdVuDXE0tnlyZKE7WO+UrN
opk8tBr9A6AXbLb6gceuzLxNGpvBInNySRLD1093XR9vMDpIQkTZsamjo97uy6j/Sanrrxgn+qXq
2aPZCtJGP8pHoV8ZtU3UVZoqw9YnZkJk/Ja0aP5S9v7nAB+MfXN/3HIfqdyV6fYYRoYThdiBq5fv
zLAJY83jLAKADz+yVhm98jE0a0SkcyIBKNikPThAQ6JC2vzkC9YzuB4nwJu4J6l013grdrNeLszu
MmKPC2MLMUgJMpW+nNT9KApdZHAlYrntlQKlCpBLcoaL05lOzqPrd2d4dC8JXyfep+/4VFVbESI/
HY+AXAU670uZaLPoUeBz9e5EXrebPP+kQBIiK7v2jLT+f5UsfCkpnUHnirsO/KIsRfewqy/0qtiW
Fun3eAbsCKG+a9IupA5rloxKnwZrRzJAm5x6dza2QzqVfaRpinw473MykYfdBCXMWjkc/o6u/jH9
YwbTqyXO2NGZ7ER04BJZyEhf+2JctoidyoKvNYZkVPBSYXmDf/Zq/yW0URKLOKI7pEXcL4+/wXOU
+fd2ZltBnUh6vFU0hyw8vxWtXLaxm9iEfmK8XfCaD6V7qpvjpOTWUnPibfC3spFlRrcOnMvYuWL4
qLXzYjM9BrgMdVsEd84u0cdQrIDR2NDKP4FEsjbPPZB3jpnha7CdSKWbGbaYcoORoWs5pxgDCwBI
abz8XiSKnp2ZVgmA7etcyCbPIlHUrSr1oeNRicMJy+WqwLYByi55cosXlgRItsJAorEuJl7oFQCp
fJDYJipKeyPk8uaNmj0pBIW3mTqiTeDZfeQ/13sJGUviut3/3w0ofAp/RPVRisA+o94mXtXN1GRV
+faPy6LTNeFKHWMrR1E9XcnFch211UJaNl02jRiHXycwsTD74Pgd5TNyljBiA23fLCFteZbgp8DJ
PK65AsCj4Kn0Vpit8+uz92R3Rsvc+XwsBY0l0arBu0bzHDN23TXEcUlwndwIpg2NCoM+vCHbij/2
qhWqpPJvzeC1N4MmLuSplRGNerFgU9+YTSzE8PJ3YuggeKcYe2SkgHUvyK3RxffRP2cfySXoRKCO
az3k8N3dU+m/qXGFQF/HnVzrRZd2Uv7TXAM7ZSbHR2voQssfqwDahD1dj6tJB72nu2fnJzNMJCjp
0CA61AutxPty4xqE/LiaV+/NPZxObqqeTm/drXo5YpqKKD5oHAPPMYUuwMnG4qEhtOFtdDXWqoyD
Rl1OOgQeF3lISHHxrToEsPQ5T5QBT2jnQjRXoV0SK7rm6X3BUSGkHCTaxpZ0DV51w4cF7dLFVoQk
KZ1F+GQwTkSLZFvoFeFfZKm6R6LN+TSGjjlSz9KcqOyWT1ZaVOiHgAJsT6lXidN39gntmExfwB51
9F4rDoez/gRlkLgr9yGO9YdQHTf4Yw5HGv1894c4Loig0b0Jjf5wS8i88E+fLhRkEqzv5dz7f0Oy
ybxAZ03R2vtbmhbvvkMwbwV6uBTs8+ekdrV6s6uKFqaVvwMreneEhNirPU/YW5AHDFzgUkCGwDDJ
u9U8Sv4ave8juPUVWvVW9QslGC1L0FsOx6mmOfAwm4tzLLy1WXrU32GPi51rwzgL/lCsWbT+h0Z9
5ZxHN0kkSGhl2gCq+zbKp2au7KjDc0XFQHeDg9J8kXDDw2ewyWhko6xR7wRQWi8BoIXmKH6dcGaU
FTOAZ2mGpu3bdsQuv+NBiDJWosqU2CswssjF1p+tS15dEHKh3jsZ0CF9x2ZHiD3PJqpUwP/OpQ6U
9omddLGad023yDD0S9+Bld9rRRIYa1fVlUHDGgdi6Hc0mu01pj7RZOP9Oj0ukRZF4bcaET7Sh7+9
DGQS2TUA5fY2xqxtYaBMRGGqQy2kPMvs50Kr9Y0Jp8dF8aXzf/tjfFJfh238qnpFVNDOtSiwPXDa
0JbkysfMyzD8Rve1w9V44sohsD6dHLU/+gP145l3US5htiLMUi+mSCfmADEeOHm9hPdkw+qmVwjY
ZymgkC6+row1lV3TisODtT5Bg4WMDPKdjmuQhUbRN1jJcXboYv5CNJ/wCtXMuyNSdqiHM3tUl/dy
t5EbV84tgknpZ0+7/RhX+bqkFj0nXvaLQ7dIJDnIsS5nAiMYfoW0lexJyLCVyAiNUb7zeb+nJ5Fc
hxsWg9TedhCw4/0V5EmRKRZ6biM61Q1G7S+RvShBnQIiHp602NfcbUz8TVIsI5y+mAUThX2W1xpT
5fRFdBqRuQwIPasvTZ5P0cUUYgJmbA8TA9/rg7MBUYAuamBRybIsTdWHX7/7gL7zMv7Emqz4YXUL
Rv54pp7aqEptQBKh0YH6SX5JL5ejJBJkvwYoL9QTsU9oqXPB9+qAVz1sMdAsKkWuTNgGAkMGBs2W
BaPfafyCuNZXhB2Xe5no+G7GYis2lspqmUoW91MEgq4JVPqHKeKUnFV7zI3qg5kb4ZXooMA1yNip
xnen60+Cx3CBPM4iL+5MtiBIQm9aky/neEO2dnW4fCz5TdfymkgcKJepdd5gy1V0kPNDBrVQl8+x
s2dYaWcoWQXaztoS/wVQYM2BnMI0SZ1B82ShFaIHErkQkf6v4mbH9L6LgGyTD5866swgOu+pCUeR
KZcrUTBJSnazyBtMUq8QAMOwyLjX/HobxsCvhUDxLtMcYwgxHdwRBpbcR7NYCrzLUFEcTLXqvtpQ
SfVNjZsQImE0yjn8ZrPtaIAJJIMrZtZCg++ddC+5Q0qTK03TqrKkym3VrQ67w9NDdFIx6uy/AL7e
X5nefwu4t37Qwyu2siTNL0MuUQU8lTnbtJL0WkxsqaoiWVKYOpbCaXDY3ey9XPXXQvq2wHYqIiwV
mXMgM85MSS1vezFfEjd+9FpCZD9KOE5G3grQ+rX8TupaZkdZZdgL1gsImv3cgnwtNhH2/R9ECGIq
lBiWYizGFLhdy6mCuAac6uFiXsCNL1zSRrcQGdZMFAnnCvT5FoDSRdhiv5GkDXw5nsVbVyat+laU
oPa5dsV7T+qyrG77PwTA0G9IvjgzzmGttwgpRz2vY+4ITxPt9ibSp59bREc1n9gR+UjIL+ik2QKA
TDh1PiPePajjd90O4Psnm5zyYjpduKgjE8ysIiscsukdobVwR/n51TtoJ1TpZRvkt8wEwEdLleDn
25lbNAda3E7yVHe+iJ3gm00a7xHdM/TdQ7WCM0p0d7RY6+LHqV7XP/ruTj39us7tJhIvP0Qys9HC
XR/CXhvdt9oePxbfL7kUjEG4aQOXCF44hjAVYx86mecs8D1lt/QOhPMFv3pByRT5/+8hFKeI4mZn
K8uRGfb6bD3yE0k487irrYnDbb8Rb+PKbA2w/WapgD13Ve7JT5ifSWrMhwBwIIy2zEBi6T74MYLJ
PcD73w5XOMvY8rI0Ohaekuej/r9cDFIsZJRwGvxjnc8l/YHI4fNx/4vJGxeOSynLZVMtl5pIoXnE
slMvx4BbzZT/bQdglDbD6Ru1PvdC8nXTeLGBn/5A+z0Rg9/Ji05gfU4IFaFebSD/MVtk19Kwk3mM
orDe1STDybff9y/sFuoHmRJ2XrDup28WgMKASsVhvAgmHMDEnXbYauHyWDwk6bxTc4IL0FaxD054
rrUn5IhrvFGGsZt7al/Tr6ICdCxHzss/R5iItsT/iXSacrNczM1HuLqZpiXZgOVIWRUwOgft8XdH
GlNJhUtypUmToiCLUTk8BG++N/kR8N9kRhv1Ke1kUQoU4633bWjs10q8013JW73BMYN15w6A8l5b
7d/0uZO498ZcGXQ+B10MOXmRCbSPqpM0srUofhac7TbS5wmL2X5woARhaA6WVPqhHNUveOo6pXwq
FbVRGCYbwLCQKLBhc9D4bOwxFju4CtP7piToKikh8PF8ZaRGrLr5yFF46q5S6vjwrrqWZLUyeigy
eAvuupZxHxPlHB5pFLWOAoHaSEiWwPd2xEtOa1lk+Q6HMPM2uWjrrGAI6gM701C4cDf6dqY44StX
ZbUXgibWaEVGp0M6r8Nq3jUR02p4klNNjeoQaM4983b2y9a+l62ydYsBza8E9NhoeeAjpHE47nm6
9IfWjgGDbxfC1PtN+LbE/ixl/+/VrxPoWpm0uRFEK3tJfQxCwKaSxU8tOiI+gOXcsGNArg7EwcD5
sDcIFtubCyzfhplVjKF15RBoiAO/nU8Vm1T/C/hetxZ4nF04rqds4QhlGvsYEApN3tNvSoJ1B7Ue
LMvMTb9upFcjguvzY5qRt2ZwpHoDuXCb04uARJ7Jwg4jqWNdVZKpffePgjrEo1852RkF+LpBgSgW
bSh/uIHYcyuFMpvWjBsktOOsMWYZ0QGbOGaLBpfiQQfv8wzCsqjpWj7GM1Abrlc7xCw2QIMfOMbo
yHvKMNhkZ5zvYLHC0ZNk/isvcOUMrg8SvQoOicUDisHww5XQXBYwLA7s0d/+7h6cOZfhQtSOIs5V
qhbMLy+LZWFMMo9AJqSHT/MlL+ukqW6sK7EFtd2xQxCCweGcKTFBA55u/SecxPw11yUgGhVH3zBW
eSCIVBYyVyrKx/MwTmCl+r1sZAAlqX9o0Poeb8EpNyjMz11PKsSw2DO1IQmDFXa+vnhNUFS8sMuJ
t69LbAkmvt0EacUYjBfZOKT+3l8R3UAqUXWEmYQ5/9+NilvtLLifs8bmSbM+sXEZCd8ddJyDUqJq
rYzOxXYIF7HLNZaf8KkF0XQzx/LA0DDPTXakRrnsBma0S+dkDSOO76jHAkFC8c+qkGao3f1y4DHP
/agWA1L6tnlNkFoDyd1hO/5wjyrwLcTxv5gcsYUPG3Bvmtl/++Hgo1ZxyNFbGPdF6dWERGbq7BsQ
UnVZdqugOGkjUW1iOcTrLdFx+qkXWjEK6bQCyqkfsBToBR64Ad2MuQMtxFu/uvAmackJxLOHnmtc
xo7QGVv3qyL8JgehdU0jxhUE45nvXDC1hV01dbh6wZGQJ8DafQeOrn5Pm3vqPY2WdFhypFYAEstM
zKlSn6/KnNMoLvB2HwZ9Iu7KPl9qSnDg7M1eDdluSYhwh0ipSJJ7d9mCaCmHRM76yc+BcQjjALZM
/WhD+N02E5FitzA+Z16oFNYdaP7ykNdaCfR8/CvZHO5FV7YLmhXw28OZPBqsPN9/8Ih3N62VSOsv
Bz4xF5SQstBVMewPxN/piYigaXBQr4LaiKXBo5SXI8xmWS4sJzMX0jK5/vOU6z17Xk0uzb6q1xZK
eJ7dW57eTnGclAfZf74SmWbalpH1+aAZOcMb3tWqTFhyILLgvaoI1taIR/NHEwBP0BUMzlXVEmIh
1APosWGJs5Aoes44jQD+zJmsOVzvxsLOy2boTF10ry1mUGZugs50+khwb6szKqF86xlNGwyf8jLI
95svqbj2tKhdSBcwJrF3I4ikblSgFGngWAHAX3Dd+mof3uHAvTJRdTyLskFI0WIAQJCer2r+s3pK
WAtlWE8Tjf7/9BpScwGuC7QA9R3vgsEP3ZEhH1DwRF17rPm5mQVUZI8A4TRVyUb4ZFe3Mi8p21J6
r3NKm09QevBrh/M/rofqRr3/omRrwhGVOYO5EHnAvC1w6E5gjmRewA9GI4MDrxngPiw3pxidKYT6
A5rJUorR5B4qA0pQPBMt5U7V9idlVcyK5adamP0YN3bH4CiINayZ61kSBChbl+P+yqc7cLz0zmZb
dQOSJ+bgC+aHNy8yCRpFJt+/bdqbSNgqzTnYU1LwS3DidB+146icS2Gi94NDVekkLIFRZYbrgjBf
bw+Io0ykL1Bjzg5WLSvDqUcGhIxLL+nf8byBjP9tlta1DNbpu5J05SWAVaYWI+B6li94prmj+sQK
i2slAjXF+2aPyUA4RU4CDSPZ4IIN8dIZatz1h9BApN8+JpqMbnTn9bgo0x+peYU7RUdJIGkUDnMs
YzjoE2mdfJ2VKAuUJ3qwV4Lm/Rz/3F+UmnkvAqsHBw9nqh50Q+cHmepYK4REB62t4KEUZ6XJplQ1
xHQI5mMeXB5iKattjE6ko2sTY+G6pgkphLpsjxhsWQZPck+wm4q7Xp+rbiVBFNJsmXScLGGaOKdO
Wig/L6EzT29Lq1KG2JL5d4AYj2ZSfcVmRz9+kHcZ49CLhi2ThZ1zT1nrumEYbUsAaxHCTQAbehtj
uBsEEbPu5q8VzjQ1YzsBXNrYi5/XK/wCFd4AIg6RYQOOGkVnypwFbCgk9vk1pcQnzZtDKjCJx4aV
+b8q9UBhvtB1lD1tychSo0R93jF+BkntAl3nYef8FiVDq0qIZ7ysPk3gcSq6HsQODw6i9hNZHz9/
VlgOnWw88FsOYRgylSA6uSNNOhX6a6F26/atOi69T1cuZQERktdznBWVo8npb5AnGCrY7cmeV0qg
28HoTAiJz+49XmH1f/Lr7FHZpIM7h5cYyz0A3YSOvdGNtyIGfTYj9J25aLc/vdy4nwzPEW9pQj4F
AV26xZ7Fg8oqT0EE+Yx7wxUPnUbTej576544jAuXwab8cJs4WVy3fqj0nKJPvAX5jXU3rcXOpBhN
oAq9LbVz2TWx0FELZ1rE/CILor2HpuTVv0G3VG8yypC2HWYPC0lrnw35DS8Asz+IZu+o8CUm9Kqq
xWRvq6v7lQbYkqkMKNYzLFKd+WaVff5NiGX3f3uSViF/DlPT8w9CpY+qPzmKVt5hep+PMUg0jZIs
2V3Ng+qdXbuX7C66356r7g7tX28KE8T2ExNJreD/vJYt0CPfmAJZ+2ZAlGz3snawfXPAT1XHxluA
zjBSo8CoMI2teHTuKhoY0kRVxZAZx0sZpGJWZ6foFkswfZGjDFiB08xOXP/m5hjpQlAO/G+G+zCY
Ff9fpuDgINN5QyvlasNjZjnSHUq3+cORdV0c/3p01VpGu42nUbvE4sHdeFrBqUB5YeifF140dN5k
dOBs2pX2TV84DD5RaGvNg9uNoEDwa5W2xYMxUV2wrjW3mB0Vvbk4VMJQ3ZaP1HdpCwqhlISQEpre
GjpeWGOhf0yDB0ZGlz+AY12kI1by5bFOVBDSTPd2aoNNB6xO2jKw3tgzQGnCAx9dUFi3qcKQqJ9C
l+sboJn0e+0Zl1cweS56yqJKVBc3Vu78qbIHgjEVsXdTo2YE2d3NedOTNZdpFyDwQO/R1xGoLBaZ
7bagY0ZhhGK+7ctUoedUhtQptxKOpPKPAbjDi01DAJfctWAOJxiwXnHQh2/ltWW/riBuKrh/AztV
fM9seKlXhd6xyF9kt6ewM3hZetZKFh6ywUIAfzXeLHocLa2U/2NnQSD8Kuen92v0PL5dYee8aLug
mknZQQ/sVHs7bXMkdqyv8eRlnlUyq6fbejRVmFXLT+YVV5gkb3V3864vhrBhaCouMmJdr1dl/hPi
toK4+mq7hnbpuM3zY+IuyzLlxwTI1iTyOcwczLhgf3JLg5atW5GcntqS7x29Fr1MK7PAHsWGyWS+
IYzg+oDwoUs/vxGqEP0Yto3WlLdX0b5UYW/cNHwkFkcwyNyJrHCizLD4ZZHRdoNPnraOAGj5nw1E
RbreRRa7kZkiV4Ff0QfrURP56FPv0AJVYeWiVXktQkyXNa4ZsoLR1gCoZsOFDR7qW9wlWemLZ3IV
5+cAP6uZM8Kq1BzD4oO9NhHiz4xwbwbz58fGBi57+FRgIO0q7ZXzZh/4Z+0dXlol9nmzphkeFAeN
iLkPtvsHPTzESyzQMwHHyOhH7ZTL2ZCf2Flk+9VU3us3VVdVubpo/YxEKNRpWn6LpdEKSNvxgpV1
9m0YOXL8yea42mu5FG/MBl6iCg6WwC1OoRu5EENkfxA+I485kawwdlCW4S6L4CMCudetFEZEb4tw
dgpNKiyY3ocgRtiCjo0MQDoK4eoFhi/FPIqcJYm/jGFGpopezsNHzpfzLlrknDR41/TehT7sB/8x
SW+8lRKiqZWxcBtXim393QDRHRR2fA/grFwXu9R0BEqBB8jTu4Nl5yNE/B5B7kWLDKr1DGhEowew
xqighDVrtxUF1M3zJxsJAYGKhNqMpdLQJTHgOfT79pU+fexzYoqwpEv5lw4BTQ2H11d9PBcyQD8d
BuooZYXG3jncMCaXzyuQc+FFxhQDBvlIN5a9isNs9tdjCeMsEYbeXxtyWnOHEdn1TQnLcJ1IQnMC
MvEmjoEPQl8UeN6ym2QI8x2vRRIZ79iHstJ0A/ncHLYLTcgc9qTwRQOOtnsZzWAJIJuIMTynt62j
5QP2PvAuffFJezkNSQXoTn3ltTMfgs9TgZzIK747kuSg6fcjENPiS49Cy0ltFFXIMb28nH1pM/im
BDjoWeC0mOdTuHB1yTs7lQ2MQErxp6+aPzKLzC1rV7jAYC1m5N+jiglhKVjR7ZT98H2Ino8qhGLV
q5Q0E10WRzMfvVEMJjvaTOKYhgDoH7+0r65TDkO0rH3y02kDM7GpNrWzN/mYxBXLVunXiYEBcxnv
Yw6PUfrHdDFImUDxfUdsauT0tuknmiNM5R7KbAb93d1mEg2/8YTDry/arP5KzCD7NTZj/Y82Y0+I
CPc6NSrcjjt+80jtv1a91KaCbQDuiKJUYxk7uUGWA2+BkspbMPWV0hgf5Jj5kyO3iBhuCOHmIC3n
6gKwUv6yhxBFrGlGUsZ1J4Qscfm3V7dtfWxAEEkD82WAG7AbnLNDrcgPwRGyVaJ0B4O9GWpypz61
e0mKVYLd7YyP0HEoM4h4Bc2rw74ubxv84C05g2OMGHY0XdNi20OTO3JPtqyMLJQfLTSSVnOXWbY9
vaq+yk7vhFGPTsHXivU9GWfETZUCYvqYfnlD9lHqt3qi53sQu+VbvXFL5byybfWRGmyH5zPpJTHh
p5zOBwsGjzR2MXu8l7wuj01nyFzP/POdrKDH177VdEJw1aBU2FYFCOMYN8ev3euqYV0jgBFTBzWC
isuFlPoFBNrTWni//QxyojnZ/A++GoQsETy4inLwmw2lTECjcKNT9oumjFb1uBASZmySMMePnxxO
8FgtA5+8kMVpoB/qdcwC+bLc/C2M5YXfSTCDXk39UBXgUnwIjAQICJTM2hzW2F/hEHJELv/EqeJh
hAu0c8aBDyX+JKQie0P/eH6TkVInJj5EUlkZlZe/ixHlkd22nJ/2fjLf2Dg6i3TO3eVbnzyaC2YT
6fkNqm92K2BejkmnxNyZqahDS8JNyFrxGnQMTgHw8wCrfUKfXdWKmUoEaqVikVxbwttdiwPIJ4eb
hJYnTZ63arHAyZWvt1fM9LY0LXBc1AvBL/6DvHhXptm0YW/PRDnhCeqiXYwYpo5GRaimTfOrEj4x
eapsDBu8At3R8qVXY4zhA87N1kvW9ZVh9qV7++8ZUTtLUSuxOw6d9Q5XbNJS5x1t8CP0rQGaXBBx
8G62V6ZSBXV8ptvklGLIIrAuhY/WHpXY0IcJtHTN2x6b5qH/uvbRoSz5MZM1h3f8qItm2YCH+SiT
fAiS/xjvYa/rH3GqW4104ld8a64e7eyZdznXHLjnNZnYdUnXLpc1yBHAAtZNsWaX8lGSNRmUDiKm
3MKmKOorem2RlJCuD4NdLlePlrTMkYU6qjVCZOjP9uC4bwLwwQQN7qeeXjci/FdZqWvstQONFp35
SKbRaCBW6jK6H7LZuZGI3HeuBGeANQE970OJ4FgeIBgBTd4lo4JJsb1Sd+wRiGmTX17IKM3du7CO
i5eHcJK0xJU49SoscutDErE0ynNRGU4RQ3+k+Vjyqc/mMjrSdgov4JueJ8+KQ2j1DBGmF1A+Ylfj
KaGsyHq2vkkNaGoj1VncxGp7iWWgmEt99lR4ivC7JkeMNwmqwS+bOidYsnFyhCuA6sY6rBek+bnM
Qet8Pcp6CmoW808vESbHZefDRcvQag0I41mU9ohoxl+EZJuJ9ZDqGpIPBXIKs4EFamHEuG9GQRI7
j0tI0lgq6bws5qAtflHmS+ADOppVk01Z++7SFsMSjtDqLfqcCM7ZrvLqvjTg3z7vLJo1kWnOloK0
1Bwn6GbDTELBwud8DgsZigpM1jwcK9rf8Ch5PJt/49um/0eRC5WRyacRpu5Sd4MpBYphyKkmMy1m
3GWQPodKjcGMWJ55UQbDLOFnjZseOXzo7kE/xTCjs2v/3rZeRr3aP94WddvC0xr8Pbr2NZY1DJTS
ekaOLoo/rxzxG5yvAkMYMoyvr5k3GBa/YB38obflHWyN0/rGUgdHx2Uoh0GQA2a44n1+V1STAHKQ
2hCBfFOB+VmX12E8XDEPsw7EDYMjMxEtQIUr5p7biOIHO547NoQTPXfNi7/kaymGDg2yeQasYeMe
J5lIAK/CZhbYpOealq4bXinVlcOxSZnjFZJiq9mkb8nIY66avuES77d7jcDitVy1KONF1Drymcd2
/QtL4XMO5pLDNI5TglcnvIVGHR/l/gr2dckxd7ZZwyF2QcVXhpAxnc1U6rHnichmb3rCTuGOSAEc
wzjSia3F9hTNgfT57PqztvAWjuwDq/KgO3MFMuBkZsGoJqwxML0UXZnYL1kw6MUJ48NHdzIycVk8
gW7xfTNHp1QIO6rvgtkLxVyU6r0VMWEuWrrRvDckXPwdSEuHohygkU+WQbV1C4Vu6pO6xrofNl7M
w75TM2jbTLhfXybUDpBN4xWny4RVToLFaUi5zwxQixhd2wIxaf5d74dTYcysrLwtzC3pBLhpt5Ad
tbsbh1QvY3HtT288rQhO/xhIftLdiIDFjlhU7NBOlj47TmIfqOzkevFLM5xm0cK5Hz+cbUAsxwKU
njU7gpaCDpB4ULPsYr4VNfc5wUaCRXV7AmDl2CtWI1iBUzC7w2SphL9s8Zjqj0CczCMuKpaLqwLA
968qEtCyV20wbUoD5ix/sTKvgWCDpLvj4Q6pqbMVUERHkMgC0k6JHQeWL6l9IuZzi29pDMonbVKs
zT/K2wu8/OUWaAzK6hhgQTZsgUj5wLtTn7eygYKQxMBFesyEk8N4yWGyGOfkchBrYdJjmc+uqKD/
8nSOHYC7qStS0qqTOqSldB/kNsmGWGKn9XkNFdBUPr+fCZuDcTslBU16fJmWVaAEtlZBE0uinzpG
Lh8mavm1DnElGLMAGgJdRJOWLk7bLjmCBQ0b5NyGqB7UwWsWz5ysN08/UfVRyV4kUrVhCwuQxvIK
WgEd9kbekcZCPbhLPD0Dh0JzUrP9qRK6ahH915zTJVXP7YH6LYfDsDbrdbA4DXR2PFOCgUd+9Y+6
gfy2vWTy9U1vXhTrNRo6cG0aN9jkAh/Uar1qWUaQIFs6z3s0f6tiSQAgZeKdC3b8ARZ5DOfXt2H5
6MpaySbRNm9B4ea01aKFuUl+PSCKj6lgzWJiGHSHU1/at9WxcEGIFEl0pQjGQ+EvF8uhv7opk9Ms
Gcz2XiLciAnnB24PMp7dYoUfPhnDeeWFFprWTV5jUlRl0Qiog0eHt5RMGXmfU04DyLaadBWYtMFZ
cqJnxK0GZjvGi9Lp5ZM+dMdiLAxxdvn2ZRW4RwaTIJLSW0T2Ee23O3C09ha6iIPYTTfSQJ24REdl
5BXT10nSoZ13EdnHpBRhloW5EvwJ83KxDNDIBE4lxJNZKx4OtlZfovepBdP36KWBbgaBWUDbkS6M
aGzU18Z/+v2p+RCm58gaksqxKJHBe00CS1QWF8fQFSRW8rgprkU1/T5B4IfaldrXxLkszVBm8R7q
K4Hm1QN/08WAI/R/atQM0tAcM3+oa90/dLVDhHfjjCyrMsr/NJKlVzQbTLnt7SM2xbKi+6ptebGf
shoJ2CWfgb6Oi99BV7bcpJKpvmZEiasjPnLaF78qhxxiD0jQBs0u9Qsq/mwnmaOxQCiXnA02l9tl
NSROu5IEhzf0e1GpZ0KheWf8eYSWGaCBgyL+SyJ13sZraxuHcYkuG0rkYt4e0JIyT6zfpBmimYkj
Dnb521n4WxoHBgHUCyV7Z4Azmz5wwNwT+PoDy40jdaVQJvTWW28vZS0qZLaDMIDMKCU1/IINq7+y
uC+3YgS94xZppRv5lxp8QwUyNIypNxtZmgrblCp+t6sUt3HgFLACIt6RHKgI3K4VwDvVzOsUyfZr
FizfAPxQZpSWerdqdZu1+wChB3k25WKLo+wMJ+FtkGaesRdlCMebFOfG6mYJdGyb15YJ9JO9h0ej
EL6CQmPc0vVRrzCPWCS7N7MUjq8nj/2V0xw+HGIR9soR1qnLUPH5Ae2QwkQToFQdRKfIqQkCN5jK
gG7Gs1viZYTDjSoVIxrB6EGwDQyeLGVO6oqT7YppMaaGZRwUXzL/GC+n/bRHB/LG/6/NWQT8Kpt4
nc6/6RfR27wFDHVDnyQKgwHWYlUQUbMPgIDckiuAE5KoW8nnG6DNnwHWXLtx57wrgbtWep/vWA3E
n1W0EVbdqsKQMWhKT2nArU4TMT1IO5kHikjfhSyjOWxBg/GSDhFXZ+hifpR3qJjMfuIjKG0c4c+u
URXVoyDbBx3odwNkjm5mLnBDnZnDN1QZUxaTzlkc4hKgSxotIxKW4FHBC9hjRC/mE5Ce+0HZMli3
4XFKSUcDyEKY9jp3iDil+rjtp50Ur0hdzZuKXnMheMJthC10eM6AzDrCiSwGfLRdb2/q6VoJQMTN
jEYutaBQSJmHxXvpFrlz1IodvTxTt9vAQ6poBEtAN9onvf8B4xEvvYYVgg6cKFV93DLrGukWzbz1
Plq7bwAL/UXhqaP8WExbP1kQimB/C7HTFs1NYVL55dYKb7L4LICyvPEV8fM/GzHZPj7XSeRbA0G7
nm9PQ7WgxaYbLSCA1MMKfBXq5uiHrrm7YJ6ac6b48p4RRO3u3WV5jMovn6yd4Fzub4TBdC9/pDta
vcC8FiO3kStvJ1w7axcTvKmEO7q1rqOblv6HdWN1h80YdRIqBRnm4aznw8GK6CUbovOJkz3+FBER
fmKwKT6Bbh0nvVXHVYl8v+PizyxhAp29EJX/L7JSbezHtykAn6TAxPi5UdEdx6xgliAbZipvFYLS
EAFR4NKvZjSiHTe4ulJ1Sqc85rdvtpY0zibjWm1aNlnv+53QdlEs1nqcSxMRX85UOMVw1Cwn0GRP
CB3BpzKXBRqgbk+Jdyyx1C1dsfT8DITaOXKikyAxSedkY7guzpST2M0wt6UT6jFUdSoL8SYFMnO+
nBmtcIS5LKZMDGSBZQUSc2UkRCg1gGT1nxhXlbqDyr/XXduuEvXRXYsb/a1CMwWlOhfLDFRjH6WX
iF3/ffaEf/zRzSw2nYL9Lf4pQwRXCZsd86GUkCvxc+Ua5cuPXTmhZpXfX5Xpi7QffA5cKvuS3MgP
H7HH7kOAuwDd2d1B5oBqhXGYosZmCbdJW/DQKKA00RxRaTRleWLj2sPIRV4CWuiyhbp2HFG0GJnE
Md+zFo11zQYq8IXMZvLK/tkYGfYCxOghknNgaZdigL6ApSBe5rYfVFamiAGpfjXr1OgAlKc8/SHb
uXSIHSabRfWsUyvzIZDWF2VgiwkRiD+aB87N8DlRw+tRuBYCzda4WqznSlu8cNYyqC0NAeCpuCDU
oXVXdnpoLgokqeOVvToLBINL1wPMxB1H6813yI7ACnJ24c091GhEZ/okOZ3hzyZmcsReCmi7g0of
nOb5RaqcolvKD+f13KAAMJMjQtZoYdAiDjlAys3vU3lJ+qc1Z2W9pQHlxih1gTDU1Rwkt1ZE0TF/
nGgC4Qzg+3RR6isTqCnw78zfamf4r8mrgkTiYPxilo80WabiBTpr4LwebyBTUR1mtPZdzcqlOeGy
01uIBuum3v/sSRJYlqPeTgwmSnMjQmdSOMeWRpLH9EsLZaGeShqpwxQXRFU2eN+roAz8C5cY0ndu
gPtbpzO1nYFG5zDg9Gwqjg+SlY6PovCgiyf1AAy8PlNJWpLEkc/VnxYeunojNGwuAXJIEGNWTHzU
2vnnLgvEDcnBY5dwL2BTr8vSwzB7XJJJOje24jkRceelwImjHFyEJhJZXCCLzDRliG5sacokp7TL
Y0nOIvwCJz7CUJyerhXWaKGY0qbRqFoqSI6+UHc47j+q+JXJvhWuEGc7pEzVnpmgosWZJMW5VyLm
YJm1AY2fuRhKJq6n21Fj+k8QG8Ay/pyX+AZ9JE7/mhNQzYlAtX9SXIBTFPaThs3Ls7TdxXWRo36F
Qr5X3cMY/ar0RKa6LFTaxD5PrBJRGOOVWjV3CC3G4U8f3///1We2f8wdiXC04TpBi0dFfOqCc/Ga
xxQQMdlbuyG0Eu3ITLNCdtOseFc8P3j7NnKEpayEjmuDLOpems7oV0L6ZCPMpQRMBNEgeiCfkja6
soa8blSB2PRHpBtouR0S0gPjQWMrfFDKcRb5mBXy8HJp8RIQ2wn8Cj5Uj2zBodGqdXhNfkvqWS7U
5nKvnRZNBVXjRXR+ne/RBdzTEoBgZojUKHiiQALh4ivrY/TFPGn1+sizXbl075aWMQT5bvJovttV
vUCCvD4At+9n4Ays0G5HlYuNwumBvHLTk6qTl67heMqjI7iUBuzwET87qgkZdmLl+be8yQmUUPZJ
eUNAICjxLgIUmg6fzk0IHCTD6YXJpEG79wAJj4kGzDTwT6SfOAobcR0zW2L5bGhFO6x9WKTijzCi
x9gc6Fp4EabqN+wvI45Yyb6ZKFfFFnt0/N+5LLeU3J8gwPLvr+OO6GXw1M6r9jEnNWxuysoNivkV
ff/AIMlb0iwR0i3qnIIgg8uTJ1mwpFu18CEF/9I22Ma0ANvM3i+zHvCq8Lj4L1ZKPCUVccJayQBm
D6HdmqNodQ72LtmMSUQi5d8zPBA8T1On5p8SLVAqBKmwmOMucSFMVD/tnk34JuPinRkLsYG7wlP0
k2tHb74tppLSXioNoKJS68O1t3htXpsySrqCE1As94QPukHKYP1HBdTbxAdydk4SPxGwP+FB7gtm
y18U6maLE+ugqTul3cQic5gLIjbW+06sNDnTCKV6nItntlQse0UFz1Ukp0RkGiGAygE8iH5VAkG1
ke7m/M4UgraQBb7oL6lTrln1dqa573kz6WwE2BgrcVyShs6ImcOMu3Py2m65DjHxBbv7nT5i4Hmc
FL2smV2K9r0wLwCyiN9ML1ntDsNDqf7U1EC75JJGk6r5Y9iegufcMDCr9Zg8KQNMLOs0cgmfqwBy
ITNa8LoH7o7lOzBd3y4ljTvUzsdAok9V5jsddcc2qdM6/5l81BDke0mb7Bwcs7O6z/aCEfVv6iYC
KhhW5wvqKX4L2FcYw4UrqlShjUG2TF3W4RwwPWyuleZc1XBKezM/wzgxk38RIPXXlO2jvc5iYIzz
vJYGu1OeDWallszfeEpJOj8RxCVkDy1SDaKKaKa9eevv6SioN1erBRkSuq3qhSwa93e3PhxilMGj
GV/FyNPFrcT8rTlJqaY5oWHTvWpBdNsZW4nH7fPunt0meU2iWdNVW8YkeGbmS4EQUyU85LRJ5CD7
ijBuK2kt0ZsZ0LQRzJIhnaTfJag7DAN4zgZuiOMSMXQ0OwPuaQE++5vzgACHZkR8WaB26bLsFAkE
ibOV8YnabcznZ3yNtKRJ6tECLM7R9c7u9ByKqcTCk6o0PjZKT8C4a39GHl/EXB8hHiKvT52M0mmS
8LBJVnEL4/zZxXcg48jE/tB+2IyYgk8sZxmRKI2gMjib8c9PDGszYVoddPKYb2vEWkZv04HKnRmE
jU+i93i+83y61PAHbf92XC3N+7MdDi8FQZnKiHRqxPH0V/bwscEWtisIaYnXygT9yLluY1j7OYco
QhOdJucNNfJlatWwiMGixY6PyOl9iOdff6m+xBkh6XTwiFg562QdA4xJeHBecbTECig4Edj54vsM
66hP4T2O2qfSM3sfDxJ1Jd7IIsyRcHhEQJHBHTr2JliUigMKRWRcsCKW4SCoRtwJi7nZEFc0Wr9V
JAET5S4mz/AFi+i44YN/DohND7XqI6Ad+A4OmUHjf4EyVEDcrN0PgkS4fdh/su3w6Cym2AeF9lf8
piUv4cf+Or1j3PZeu1l82iFOmQEKzwKq6dgeX0CHyJcJ0MCdI6hatA5Jel0RerB7FaPTMnD4uy9v
1xLsI5uH6leExBqnPWfIgJY5Va6Ohd1pq1vB3p06ahEjxRsCjCfKStTAj11hTmAeVWcM1KsHcBOc
Lmqxx1oBbbyHwIEEYPaH5+CYPCh6Na7+20kQgsbwRgWDKNFXmKHKV6Q2IfjpVp2MPB4uh0YMDhWm
gGSgq47WPP/EGJgwh8zZulXtHt6s/iUR4bsepTkLvTcUoiQZa6Yyy4IJTaHsxsasGfmCuotveniW
fEXhMG84ogYIV5yp4qEYPTWnNfohmuvuq0Kf4XnY2CJ2ETuS8Te1StlI43JMR80aGq319nGKa76L
lYlDQ6TZbSJtJHzX+PmnhENep8PiP96/6Z5SNT/gTe2U6IA8mWBT2KCt7s0qY5jVJnKKFOuTuB4y
4aQ/+ZFqOFZW9sfIdl8Oe9UuXuT/nnuNEOAhaWfcn4jcvWTJtZIw7cWwiK7ki2QpTRmR1Npl62me
3DHV4Y2jrYrL6fPltzUKFhGV6fUpXFbM80txn6hVoI47SCT9Ky+Qq1+DPXC4ZHFaMWUFUM1sOBN1
nsU6aW+JD9AQMe5/W1wtjLwslrrpT5CyqaahIY5Nw2z8Y2xh4qNMd/gIP02u1o0UvfP1+IwubtZH
Scqlwv9IZmNJsDfaatMHyHpxg7e9ggauqjX20iPaBbD7YI1a1Jh+id5zSzpPAyDeXLkOusQhEuGw
O4P5nK/6N4AtCiHuiICvGeCepPxOgbqbBip+xvdFTbOlq6G3HUTvU8nfX8UVKvbGyKCSUEI52uBj
2pv7vVEnPCXeEzv3+u7YVeK17lQsICwhb1yqUkuV6J/rCt4j9MK+hhpng4Lm+ncNiIYYApkVeVL1
F5c76zytXCXGGuYhZQAgN+wi6HrrfxXodV4soTRHBWDcJ7HfbWGECq8mXWooiqXkFXEU+wXh5Xue
xObzo9dY1H7+gCL0LroVDvQhoiGmvADpou2YWTp57pLj7AHuVdIbbUzhlQy7V3o8B/FU37pEyPP7
SRj9qxBAaKQwYZ8NKabP8LxndDBXMp7U/7g+2x2ILQddg8ZzOBtSln8bWJaDbU1+ItEHTDW7gJy7
upq7kf0KbHqrTQ99hJGQhpTJ2kPyxiqj7rCbNbdPKPILz48mIYgLX0J7OxXYjhJU0w1xRWHzumLw
OtRjcgV9S3ehJe8lUtSx66h3ICsCG9m8y8OKZ/rznbxH1mIr2EOa+KMeseIF1Bt9T9/RVFFjyAJ3
Fzt0AmmBCZgCMHR4PMvBYKJLqaimmisgHrZwa8MAL+KWu0e7LXREjoXq9rVWoTfnOwrk4okW0urM
UrL10+cryTPYg2USyFbf2If8FfaUTeV44aeJciv5oc3Cei1HCRomVpzcB3OccFpaJEUEFH2XQXXS
SeWYly6TkaaNDF09tvKhKaedtBhOJdDMwv5Udh0Ptkogwd6rcrM4cRslpeIp02+iG7YvgN7dJKV+
nU4dNDa+uFEhaKhtynpuJwJxu8qi9axHJTierPtsRAjA2uJjJ0geJ4ZhvTJYcGiw/yGL1UVBIpKL
xs0utOLa9Y1RJ/hz7Ky63jwn3DUHqKTjlIBHv/tUnuNGpU2BaLtGrOOTnb6LVUzmBwqinhUmp/Zk
f7X0ehCjTCo/pH/ik6TUsfTQLqkjs20/lTYrc+q5SWqnccVWTK8KvEFN/DPbMz4jkwg3DnjtDI1J
j4RjEqO8/Fqpxjvbpi/JK8AABHF2CqQO2dpKnM5IOPzLl9ekf23lrHEdkOfwqF8MT/fKsdggEAma
a0Th6DA6VAG5EnC0J5G66HrmWRCLac1gsdrMd0PLNDBOiZpxZRqC7QlQnSVDZz1UpKGQDGWitMyf
TPS9Tyf12edGhNJlKAOHTy87NxuEYsil7cfqYTWRlS4bdy7xIeQzMsitgPrFVW1rq0vuJFAfHJJU
Wvn2ZxtNasY+7+6Ck+j3KR3J+rDBttpy80VbnBiyEmy5yNfOUZujXNGSzaItLbYCz7BL3+rDHKiz
NhyyIL0B/ChjAkSOCzlfCD9svuYwUpYCxoGHWPirK4pRMr0ZHwo6SUQzdQTqy7omSO41cxOiK8J+
LIKgGbLUG1Jj+Q6hrDBskkMNp80Ud27taRmjuF+o3ZV34zSYK1KDvDrTltrK8nr0Mkrctxbj/6kQ
3csJq6emsHTiuCEgOw5hq83Vch7PbpzDrp+m7PNv1rjrtTxbjbWndweHchruxhofl6t6LbYRpxzH
iRbFE2Z6SB6R7ECfx1N2fcppNpVlBKLmqqGL6dfCfen8IVIIMYq9z38vPrPbOytmV6NFgA+4Z6FA
1StBLp6PD9pp7BpYJRAKKzTHP60xcjGitcTrHout1dBe9iNCT8Oq3JBBCM/cIuqaoO9pr+qUCAtz
htJ1DWYjV9h21woIuw6XuBuf2/1QfxKsv0Lyzwyj/PjBw8EYfMPyhMemC5+gP7TtQNERDuSQN0cI
UZXJTVbTOu9tD55OKkL+H6WrbfJihRG+Ajt0yykh5q0AUdU0cADBRdgGeCfXzodoa5pCFg8kcNYN
309ilcBIfwVkAH+XdGKyFe9DIIUfVZ6uNpe9lE8pEhzzUbJGqCBWt8pJtcGiW1Xg6U1E63IS19/H
y/Qps+C85MYCm+jaJAJ3OH3pfeAmC8audvMUniB7IprvFSfTG2Ni8JAapXGSB5KGc4zaesYbtTBc
TVroIQNcRutxpUOoCQyO1snAsfMsozMlF3/PKZW7iLjTPZ21C/p7qN6LNHqTemAitsKpzLVk94AJ
QpAYTMIYDYls40q1qY4smpJd50IOgbwWghIKN/UBX0ysFO8PcfULr18WnkfCp/chZINNiZHNqE6A
JahQU7foPC5LIBmnYb/4NbROzrfRtMFgDFhRIcJCQNo0S7/IAST0zB9Rne0Z32Wo64cENwTkD57U
N+tyGrnUpCtQQtJO7GMVXQNb+pkh9gtnqc1ZcMrMhv//ZdpbCn9t+lO+fEWxJ+3w1+E4UlavRPfm
4MS/tIDqrEQ+frXDHg2hinjyyiaUmq4kcB29Lc/PFZyXiDrLZ2JIbRjbbzkmoafneHnllkD7JD/6
uV2cFPYSbo9vpemQtRhW6QPuMIW+YRr08Tm7XjWtBSX3CQqOxo4EhLqzrU+1TAK9ZawlLCCLFVLF
7NSr+jfqrpgWG8D+AkbQZXQjkf833Mf58+2JSpiMyMG4JEzpklDpGMki7nRdnqanFenfL3mIlsVG
1kYCHGFqXjjVbmtP5QV0yC5Zo8DAAcv2i6ilHAcvHe9GjJ6YM02vOvd0s90WeT8NpNBYB6dFcCDp
tVHwj6B7WUfDwAbP829Et/v+E++5NHkIL177FYXZcww7SUtobguo291HIlU8y7S4z8REW+e54rh4
xzghoG06HkY1MKdxjgtIT8w7w0ijI7LE/ZJBRfqBcbZSTMTMWdIOhcsTlrIbY4KSYAYsKdU/yaZk
QGBntslQECQ+rZDTZVWR6vWc86OyNkaeL4OyeP8dMuGn9aWLzdWb153NIT4wVr1az2+lqUskOAtE
Z55q1AEsV3Alw0zjBTCslsyZcbkutRq+TXeI8YuBVOvxjjDcff5PaMcYWQp+PSS4hP4kUIHaZfHB
WH70b9+BAmOeg/oR0P/b+Gs2XCl2CVEQqyKCsguGf6jgVQp2NmDt76L8jUZibj8aDZMqwT6sPpqo
dugB0Bz4zTxfSnIsEkEVimGonuWNjLna+1nIdMvOh86W8ZmPXyb9bcNV9xNHQeFSNb9ixEUtUO2U
FSrw58ySlHRwloakUwfrebyo4vA4oX7xr2LPF/B958ldGbV/Ri70eQW3pu05Ou8UektUxx+gIeWV
EIy9mX+3BjsxRPPSLIeseBgkUaDueDeCV0/l47l2CuTCUZwApz+ARqZLeTqWyLUHY/s6gGewd790
1OPJhRs0AxGwFn4RnD8Lrg1tLzG/0fxc9R9EiN2YFW20NOiTdusiKsuu/A0ThIp4hoWiMl8kie45
PJ8mAzB+d+Lh09hjwGLoqbs9dDECblkYCi9JmJKIbF5s5E5smx8PFmRXfcE4Y7zUK5Phlj/x9O7a
rDMsUlFzAk09DPmrwWXfKf4CnXVA8adcAVuLQvM4cgi6t56x2WqKcZBxYIj7uwUMpSeLHDSIlNEa
e8wFeeacEEfo9YTfy0ACx0sQWlPvfEJ63jMA0rKHGgLq2NqYy6UYiUEgLWP1HBijghth+TJ+VLNu
mNV+7lvZcsOMl0yv32FhXm4y4UvFVtGwbMpjS8pFQNSVTCZc2yvW07ApSVilvl2hE/PueoWMuf8Q
vNVsrVsyLsNIjJnQQq7z72w/pJfmPkrZ02LWZ55f/smrBzd3Kfj0WceRM6HCBp3sy0O7uCtS+o+p
hNaVQwcv5Tm/HR5qpNMg32Uevw8KJEVdwG0I23E1I0ECuJSLXh7+veKPKqX6B9D9cBkiZbAUwiEf
jtd9O7xOtBU+/DQpLS0sVsfEqk/iV/Smwsf1+nsy4jo/Nh8NTRysAcAaYBKapcFX8WbzVAoPsImJ
UlpKM5Q6vVfHAlcHQ6cUnVyGSv7UZe8+s/kTUKouPlUj5azQoCytgd8xLD4CGVS18Bw2uxL5NqWp
UXCCpjceHEiuEstU9a2zuL8qwNB48vsIDrCUjdnhfxgTKiZV5PTgR3/O9exQoR5XxEqbE8vo4b4W
PfzayzkpRcmCp6q3Qlv4vtPeQQSIwCLNifmfOhc6j4cd57aZYEepK4FmuR29lBcBu69WRrzNoOOl
O7SV0m43NYhgwh3079mWAMikq288bDNcq47umnyV+UlIRJbgVC5BmyuaRbU3MALRjURZ/XnvAr5D
+g/eTNZ/D1lLoB03c2EnNkcQCrkwJytXDoo61EbQnVDsMHL2G/VZb8dKgIhZrhKDvnH96k8QU2Bc
OT2uv1REKRvK4YTQSmtEfjVe17rF0nRruTvoQOXmn9DKX28IJHF03PFGKU0gS5JWSvXhjNBv4jZ1
KxHerVnheNngWbhMNv4VgvapK4a1ctPRRy4Ighnk0sPfJeZu1GiSpmsJTttqqyvjDlYQR7/+aP1G
Qf6qyQHEVB0gvWtYdQlGX1gyhvwvXjPaJAT/wSU9Mb8m+wxGT4a/KuuydlvZoB8Kv+y6Y8p48C0m
HZ3ENw7R5g4tF7hbgb/iDTeqwUDEKxsPtSBHz6gWRZCO3Gbnc2gFDs1z5fMYZYuUKX13ZEyKU4md
5Y5D8HqaLH2khc6YJxjufdWgul4NzwC9wzIHAQtwZFcYeb3TnHOTfpeKwhkWPgnht0/VShu/NBPk
IDcRJA/oDd3AVFNAvQWN0Wm5ISivxXpbzoWxR5OM2wHuSZSjVDW7cm6wthAQY6rbREHYFe/u9iwj
wx7WqgrdLf4Td3dhgpLrDWyQ3QahCag5QL+48thiHwU0ZefFDUXW0GaCyoqu2VT/Fa1Tl+AEs2PX
VCn4BsTQX7UXE3fAqJDXWLVQGJlp5WAmedfHfjJuBwyhSxeQAYAs/hU44Zp8FmLiGTpG3ewDGYoz
ta3az+WTP38wKYOZ5mb/pYwY7q1XJyn0dswdlupzf8MqqRh1FnwD+mXlZ5UUDgu8aKc8GUqNDLA+
wZ4oVzMyoOTuecq1bb4mqrMMS39xBT8E3+fGnWrBaVLvEn6bPV8NzmtrvcTWM1+a0dWF4xx7ibCA
LzFZxVp6sdPv5LQDv9IqAr+kJMtuP4Bkv6VkB4sfHycqy8b3H+qUQVCvbIM8Oq3tdowUhjPcrJSM
CS9mzz/sfI3RZsU6DTy9E6tLFMO3IdsI7xXfozLElGPEk0i7EVGj1ZUwFy7c/qyovkEFYzKYSdJQ
xyvdHVUwiWRNFVuCPTC87Fx3bhdQDonUCkrARXSH/Oda588fkboAlGv/C44gHQDOEvaSGDBDwuGU
2p+1F27P0JNqVjiyTl6e4OwzSiUf/HJT/z0ZIPnmfyZeUSSL24rHUbA+JY/dm0U+vhQEYYYYdfhz
A8s0iG7va1FwzkOcMbBhGTN/C/++W8tWMj5i8mosmPUNN8Aao//Rs+GsyrefQt/KPs9xXYTV7GKM
qNs7vaR5oThp7c9ZqoDj1Z+ppjPkHCo8JLJAfHhScuHFOiEEeHrkpf73OV3tBH3ZWt+N9/+1K3UR
uL9NnSPsbftuMxAIjuEY6sLVxIhvCDGPPcJhwT+6WhZX3DKLfpDyZVoi1j7O6NhTYpumR4Ye9/MD
efUZCKUCUKqnS/Vk7M4EIszBMa2HasiXFmMyNLOEXPEA/qoExGw1aYujBQXRvnDMJHBLkFBPd2MB
p6dw+Aj8CccNEdHIyT+A8CVSdZk4oephcwvi+YOK6kM8jlEnxbPVvoF65UY5j7MyScgBmKKcnCqs
BKXfO83VuFgHXHhAXeazIeS5sUdTO8JadDDj+ya64p3GzmYmaK+/63r3+WXgx5UnEAYctNNvsloV
GrVu6/vpGsZvCKwV7K8Cb9KodC5PtDDlLK6nLx9wmVwd7vjaNaYIsY39f0uQllpLgmCFQkiKaAfo
uHj3okSB+ejvuvC1OK2QOHgZ8R0YY4/cwuBdc4KEQoRB9fDQMWILXR27TPgkw0AzLQAYqr926lc7
oPcE8tMEXR3jYkQiYtCmsaTV86hAfA60CmMzJXVQHpwpUWWux+Q7GdVzeVAZoxkFtqrst1l97mcs
6YcjcLYXhP7Lb/XpZ/9g1bYPs9myQk6mh4M7osQRYt62L+imYK2rHu95OJrjs7CeEbGJlBxOeUbN
hPG+5DL4n0cn4Dgbud3ha1HxX9LI5khZgs/AdZvLCDtTarmLGcQdnhekOhFuNi4asExcNLH3Zosw
NcqWb62D4MayA+UBJW8Jou1ik0bpZ61cd5bAuBDK7eShJKabZ67bW076Q/9wTFZco43I4HTW1Od0
MbiJtlEtVR4i8vjtPsWLshriOLTf082fOhW0sYlVNa44RHuhXuAJFXQktijHIYXvQALT97k5e0t1
91Qe7wWLtR4oLxjS8fvkv7bSN3vRcOZrotOxSymJBq9v6UazrXx5G1SWlJkEXJe04EAi21bfwfK8
PDejeC/2lozcY8V5g2Fo0Q8iEpJZESJQMIgHbWOcG9ioPuyHR7XIuGInJRb3mjFHyawyWiWBaVjG
W6n/vvFeOGN2O3qyMUCAb+L3lYbrgMmvAwRTUD78mDxqZgpAB89sxOG8W7fP6636JBw1z12feds8
vIF70JuYk4+aQxV0O9rahkCOBzTN75d71PxE3gCjAJbE+RBiKqu8bYz66c9eorxHgYmZGkOHqnZQ
+62/77mpVWj2Rk9BwpdMKyckaqHad5LVf3+Zn3zZkQ5z0UfuY35Q5LHZl5OOA6EjaEzJbzeyU0KN
YXXo4HrTvLmuswO1/pe8qwRMKuD8+3wkb1JLx++QGwOf8WY1b90ndrNeo7NFaO2wFAzSYsOdftlx
AEshIGtL3LJeYh2oeeUEfXtbtbKCIVmxZyJ/VIRukZNcDohakJh90RC6p2Zw1m6OJqQVs3ZA6/fv
aGIZIEnlJZphRfQ/hrkLvctKUk86u5OuKAiSKM/9O4Q0WwIZWJjEFuVFXgHCCtL7oqJBYizd4AE1
WYZVlrb+vug/uT2NZIQG/fBnSy8rRxWBftzE2dWqtJZEg8dzGT6yhMyYfhHCH5qNhwGCsx+eIAG2
IJxBc8cxvqvZN09NvWV0NhDgspsO1PQ2VSJCRbWdbp9V4AaCMpjNYmDgjKOvqDWs0o8WDkVgs3Dk
ipwNpqbujmaIR4DTs0PtuWEhf7ZCJ7GqFSBG0AjE6eSbnn2V925l7wRaRMjzVqcJjzUFF0bUVgdy
ie7WSVdlDHhcSSlNAtUlreZfT2aTINtCWtT668pi16FLeCcTXNV1+4g/voWoLUeWOQJ4cfftAg3m
59WMISfvv3716nufUbmJrSJ7yme0+nTrmhaY2JBeq+KxBPupbAkUgdJBQdd49zP+32aIr6bnHSnO
Rcy6yQN6ez9khddsTJGUmKpLXghOgLGCi+EwqzXOnpn9QbxKPHfO9lXIoLEMoiHF6BSpQd0ZtwC/
k3nN9k0+QS7RP6eriAF/nG8OjT2sjUKO9Jd2irZMaJ8kCRaEBYUlVJX815DRm69BeMPHHgSSr69o
KJBsu/+UwEsYqkW2TB/q1nR/TkcM4NLz2WAFIgvZ4CnL6saBLGqji7J4I9k3Nb/lAxla6bxNyZon
HGl6gzQ51xG05ANtXvfRnNjqm4Qo1drOrB/Ws7sHl1ErLAYGtJIsjzPLFRwJ4KjJkxpbV2WbIfX8
xFzP3jvgaYzwpy9Ev3o3PEMPBp1l0G2dBP3A61sxjNWyF1Ij1mOove/n8QR11FZi7Cf4MiwvEnVy
tiBtZoTEV1+e9/uBVhShMtrJwO6y30ALzBfEzHSFSiH/pX24mc3f4paltVTS635V4Ili6NhpVq0j
JNHsFGhOulWdjMhTmFfSwTnv3Uh940BSoKLiE/bQH33P/UqQK2irZkC7ttk8UN5xjfmNGp/VX38O
yYDZjCFasdJiJUhHeuIKWov8WnpguASMB2mwZKDZu6I96oYkk6SAlxQ9JHZfWOZYlZ81uBTrxvWF
sGVx1IpVIOwrs1jnK4D/ECzsIzmOw5RfvDliUjBl2fwOLMl54Q63hToY/VhAdSbMB5hR3dhUxNI1
9OEYc7ar/yZo2/AhE4Bn0hKJa6FbUFJJ6B5DL04LFQI+vKkATRZMmR0i5YgJ4p9pch6Eyq3+ovOc
Ld3mp6u6RfXS8wGD5BP9lvCE1iqAzRe+eKHbhBizFTyAIljWBRghADj8Ifcj1kJ+f35A4LG61lIn
Zu1U8LawTSdfngxTdPnHzNwIhaX44751bklZvnLCamUmj23M7/qyGX3Rje7RE4NW3wD5JofkMzTJ
DgtzCFroDrPeJfkwj+TnMkWalVnRJUg30UKRfnJstSpaYQGO2SzN7PxIF7GXpdKIb976fT9nMFpC
Rc2LY7U10CcuuL7LIazmlOfC6Y2hUdQgzNwQN1esvn+Ov2KJx+ZtbBmSH2fg9rvYRH+jH9XRDITA
4mOi6sWPIYoJwNk9qfmqvv9m6x2EqA7aKkuIhBzfwMlnkw0dFYMFLsZwVGVquWcailWtrRKMMW2o
5t45MCTakwGObUfr7ew58XRA/x1rVgtvzGnlyFjcjVLxUSf9N7iggYQfCZ8mGSVvGum+INEQRbsQ
c0Vbs6rwsf0DdRp6CGfjXK5pXqM8JcT1rkd/DuNli6VidjpGXZnXtW9Iyue2TnrQ30FPcNL2RVBt
d3LC3a/z5jVIX+mTuB+eRSQEo0Te7NMdch5iIi4hzeYgUJuZxksTMcHyNME+8gYEt460VUyOGV8A
GLFrAG71LkGQVyeu6d01XTpyyxDQ+7NitvgvzfBPwVoi5NYkbA2BEWqJPhjFiP4nuw51tgA2FsYM
mnqoVIJXpxhOzi/yybEGLz7lhvGWpMekSIPlD2mpoW+rMtL8mS50/ZsYnpt1PhjBNkzfDKo5XquY
KT6pvdRqjLqQqwB2kbvGvQVDCkN/g0POhA3ZElbEDrtu8HLKaBQEMLqycDMafJWHA2Fpp/OZ9dFQ
ir9jTiDJAZC+DG6yJRnGmE8RG0e0T8CUfOYXKvZGPWA3XAqbDjUzYts/F983CktWU5zkb3ng73tn
UN8ZE6TLdVbwIYuci3redZd4XQANDmc2IrLGvLy0VoWPr1rzjoNTP/PajBEqo/v0FSTh1V+iI+2e
futMhghBaF0DcDaHZxdQLg+DQrk+iC/ouJ/FWBqcLubil5Z2AzZx0MNtqNpXPme4ku0l6B6+0SpO
9GMt+0WO+JtRAraMYBxt4H70vAaTV7LnSvuCN1Px1ps4qUQFabGZAY3ZfLjCSOnjI8RygSvaMhOL
3D2mZAVw1APs2dVjjVACedl+pKujZCVtP2zZGt/wLvH2h/2r7G1g5rGCJArGYh5YZmRwJ5QZWGBp
w8mD37iFLOHbl3gtxGI0kxYqX6ddzcuOK3pUlQpHvI1IlSi62Mzpqitn023l7aAoNcXMNuomBWOr
iakQ4MkSf8opLepu4ziVKZCwlNzfCu8v8gEszScfJrRsQJ5a1Sk0kPcBoHSc3WvGwP6dP3ux5pFQ
+/f2KPU00ipAFz0qHrXOZKwxBGE4twl3qeoEH0OKaVrf5K1uWn/uDq7ixaxjpMQya/OHNDVAlc9u
Myz5hJTKxhFV/b9h42aM7AHYgTsC12pWUR35ydKboEd86YuIRT86PFxGcZb34rP9m3f8gsCukb4B
+AWxImNHdIGunceG43pznXVmzKTrKN3omTs08E2zFBb2F4bc8Z2GcptrWaLboVTmajsW5PQz348c
mxSGpKfSI+no+E4k8yCMUmQBuIEMAcvFnzz3SdJtwdjEC20n8apmBrx4FVylyORGPMlMxlyrwizW
UF1hWbCUV7KadAG/qgVlg5tb3G8GlAFcEkiGkYEvwmGSyRUXg+Z49ui+8BQCafwlAbkTU/y6IHvg
UcIkjZbI1nKGbSHGy44ywLDXsQnbrP6KXhqFMOQBSu7x3mHySisydc1BPnA3Ggpz3nEwVe6aMxNM
OVtPNBA1NAcoh/A9nXlKUV6i6KsZbrYdFXtbJU4D55dzZcPWBaeALzWh2frjf4lt5VOH9DZNjk/U
LHNvFuPsOxogc4yY3apzS76lnHXyRR50GZs4jJlx2raQk51clBAwMjO8ix8y16btKIMdWCVExAHs
ToqgVUV5aq6fzmGxSr1EC5NvPq8GDWFS97mQ8wkRlqwx8RgstICUUBWuzF9VajoJKhFE9j2RtY2n
tkRxgvVBL8i6zjchx/k2gKaEmi6xMjy62qyiofiHK5MnFAPX1o0pqMW8uyrTnvump+phm/Axh2HC
t55hG8YIrRk20dGakpfbfW53EjJBjqHhtyHQcz5qi8p+yGFeIRYPqW68EVKhjx0KRlf1tD0y2UFV
nDiBdTkcPeQztPn0oVJuAsvc88j72LC1g9atbGHRzgQ281G+EMuebVtxl2lK4aiT14COEt+DJD+p
+pVR4WKbDHwjyLyJJ7uMV4MZ/Gwn4OqpCpH+3PMUnl+V98HdQjpcjigqCQuRMm+yVYhe76Gkb9vD
K6iF65x3Q2kjSfRG+fH6qtRzHfy2ZJwULfign9vXu3+JYZiP2t0G7btIiQ07yvRsZH3BZI0E+dnO
zdBcmwgOJMQjTHCaKc8V+VI2bbHLuZoJkpnsgVuUmKbcYZ+7PRZp3LCaKKeGaIgdRwdrOeUuTfPt
jnq47TP3UNqM2Eh7E/jG+CNwwTFAe0kKCSnAwqdftyVEnMR/ow7sRhH5oISLMWBqXB0V7PZi/8iv
vGJWK70ZN36k8vkglEPtQS9EUsNIHkdreJ3orbm77z6mtgLRrqrElVawlkMfCWkAKeS+fjye/Jhn
fzmxi4mnYYjYx29JUcP0FWPDiDU1aG88TOyjB7OmfIV3yD+DTDKcE7PjWRYChn3FjgdCFKePaRSI
qjILyNCcyU+I+yc580zUNoBll8ed2N2mlvZH5i8XxXQvUvb0RPoYQtXFclMlPqfepXI1wWoFJ8nZ
TqAzSNs17Aeq82h9OHKRZMrJ8/hq4OaiH6EUFnpoyON3t6WP/L+ut12VRvGEzUnyBWYHb55ZRN8P
IcIdNfVCQFmBCqc5tDUxkMiEv729S5CnJGfbDVbw/sHSlNTWJp64QRSZiR4vW4Im3x4Cf5ocMRPk
qyQDLS2j5zJXpicRA5RVNfGpbAywI6P/ieSg8KrekIqkXp2YL6o4P7gKJ7l6yJpPesjLlH6ShBHi
a4huwgKKA5X66GJoUQfrjLOIqMs54QaBabEO80ZnlTbVGXMoC8OD4fg8l5OtGnVtzU0Xbbb2giPL
81Ktw5hwa0QG4RkUGvoBYvmuTuLtyQbaBKTPqP5ZV2agSJZu9q6v2mZpsDuXupOceGGu7k31Xf2Q
orYwW4J9MnfQQvG6SZv04FGw0krFQyL2DxfqCkRfDvlPQcMStLzk246mC+tS5oLE8+Kh3UmKqvJg
nkiMRqp4obJUQ+uSeCtyoVo05mB8QrV5nXA6IAVwdP4irYfRv6fyTcSflNjDcUm3ZXj0XdXK2twV
+Ouqqq1LFnolN8hCNAeTA1bKaHU7XNmGf4emnUQe7VP1YnwanbGTcaXszfVw9tKq0Viy5aHWhqWp
oZy9C0r39QUpxT1SaxyFYPl+WYHTMwAbL0VnxlgqOaE3XrGrrdak6B3GNNaoA88dsUopXX6omAhJ
bvVP7fVedcKEirYaGK3OfhJCF1ImjYtMW+ruXUql1cBuWSmUiTLcL1RogCm0JAVAlDq8qSPt9mbr
xoPu0gG2uCA1GnXFmAZ9VdH2XHi/3hWuFCCCSEfpSMkFU+ln3bzg2o0Nk7E49VWauMi+CJRPfxvF
aGi2fS25qJZmJ/FSpXGBH1TPe06Zyc/BUJBSDSw8j4hMmLIV4V23LA68Tt1xaCKvSQKGtPXQikN/
zWBmUGHyjXLqbG1gHJ/kJXI3WKAgNNP9OGtMINXJhhdCHHwsF44LSadg2hFwKl4LVEWKA/hpyFbb
s6oU1zwj3/8VZMe35kdqZevJ4CFGaMUqPt5U+5m0MAqM5r6AvAYS2qKXnp2Sj4lVBjRXURVzZ+/x
A5t7/u9UYgFG4nWBmMmF4PiUi/qmt6E0mxORBL6+lXUWWGRJaFf4DNOvyMLbAwkNWnpn2WnlMD71
iwLP9dRXREARdQC45hW165bIbvkQtJzmYDIazLhywZ6bElgAVRF7xYSWoBLQYf96WHISLIBGd76y
567IF2VJ2/taS4Aas9chGH3CkhqRD8uPaYJMHxzUinSajqUTvyqLj349F6vFLIklyi1MzouoHsha
4x9tlCjHSF0fhg78zyToSX+IRXQaN9xEgU31ZIWFhAH39mPcej1ns/QS+2nZslCx8iS48suAKWus
ou28Bw1S7nkp6VPZMMq0rhAB+CnOf+9DfEGXze0f8Foyxyi3jZkUW5xZCDHVOwONP23URtCo34fO
tA6DP4w+iYwoweliu1WkPjy0n0m6Ddnu/3mvBvyjNdWcNkcP9tyEY0YDtMaddx4mL94qBhV4H4NA
cfXjueuiIpXoofO2QkkyK/kXqqZrXfo/0x9Io6PyNmbr7N4L9F95qousYdgwasUXDCmpacJtbMxq
nW+sQW7GWll60D8L6rY0UAlBu/SbqmD8CDUYk58r8hYdIkngYHriz2Aymvi6W+W7PvPZKKsWxBie
CWRbBFchCC/H79/cTaOmvS6UG+cr5RgCvGSFgrAnesLF/Ct9W5SkrS8KbE0MKiSIQZKiB/LTz645
qt5lBZHdojtJOFoZOJ3h32RrGKQ+3V7t3dS+Yqna6euXibLdyGQkJ4EQx0WxyNm2k92Dzbl9aawi
5cBFq6Vh2+ABE/wTrmeft/SOL9lZfr5TKpS2+/wodsDukvxuMb3GNFc0NfcmMVSBjCIxLEWlP2Eq
kLn8CX62j1gf7msdkEp/L1dcKkOjI4pbHSlIAFo+/E5RDv1gFXDgSfKquLrGqQZbKwuORloFbnZO
O4m0TO90YxYCoIOgklJIqC8Bx5Jq6zMrxw6xhcKyNEH/urvGkSzACCEyU15L2gRj48jZSNFsbIgN
OJhMoSieqr9N5pvpMrRw6IFWRDNtAJuimhz4iVfwMizRZQA/puGclI2yjY+q071YSCs20rwGj3sS
YM/buTlWWQr2tqpicYoH+eyjFrTOftTlATCCONxP2gVtlSpaKbl73yEQEzJDa+l1Tf4GIfV8Fq/N
ySfAxeaO2K0P2ArlT0ZPuAbZToUoRQ5W25sF68ALl41tp0lMlsTm6qyRUnKrdZdnGKN1kjymoDW2
3JsgfRsA53SPZJFuKZ8A6w3JCUQCeMzUMcUf4Kk9h2WNqof7nhA46zIZwSpwd9wqcX1OigymD5sv
2pgh8RZ/kqPxHHmWEO7RCs4jVA+2bh6o/wfr4sNIjfWtKhY/peRuT2V+bnVIuO8RnhTIVBClTcyQ
vkOauU63VzMWEPpqK6EgbcM4B/Z60LBihGYSzLy9Bs/sQXr2MZ688IExdzWKfBskkb+B+XdjdzsI
cJDptrs6AkppiRhdZBXtt7eZxMoCahF508ppBls8YeCWeaMpC2J+Dn3HzdXCFKaxMU5g65Og7KOp
HAukB3D7gvgUYjZNA88OseUfsaNeO1E7HfO8d0IjCxt6NdGdzu38x9XUxfYp0dsm9dypicgMU3lJ
wWjkgIgoBZN5yDcQOynCRD+HVnH0OZBoBc4mfpwQOfRKlsG2yDWWR/q8acNFnCwpG8WaS6Xd3U+T
uzGxuOOYVr10MAti6LkqcrsfB7CUabpnfXyqdDrgibfKCAX3lGH3xq76K/PfISV/q6tvTwPq8SJQ
2NIYzr7iKDUZEkIH+qCKwAYNFGZOWebbp2FfZpgoyq1JsT6F/E1rQVt+wVpamFygMvz1EiL5ZcTr
98O9CCoJgFn6PHD3FkRbFyNcgnnJNBvk+Z1wbwQRpOsrUPfWKBY3Uncd5WZUr/MeEN9kTZKwJcsz
DvkiAKNtMbc0i/7w2qxIIfp8RnaGwagAiKWKNnvJoTixSbfLk39991BW3a268d7e4ygGRNehudEM
uHVBPQqwYMzCW7Lq+5VahvG+/YmuzkLsUuSRCKDjo1NEB6XyHFfPQP6iJOZ1vPAURHb6Rv+biulL
+MZ7RCEsrAub2T5QK63P2DOxLkeX2Kr9FVD7zjU01MEwJHTtBsP+K7mbASMkWtwCFoXQHxwTxFEe
SbB9b60krGwakqQqMzT6Yzcq7HOoXctLUXc6iKFv6xlyuXOS1j9SzZJRzxnWww2pRp8TeH0vugG4
fmt1O1ZFtfNQ52YCoXmjS2mImLPiwrBmDpVeJ3zICmjQIx6byL6QDGaf36BLUNtSY/r9O4eitXHv
N0PpuQv4O1bBVXuxm5IcBhhRoQ3QGEm9uFJ/AYKoKGMNciDOtf6496GVgy07dAnvDOv0TePEcc0e
x7xomj0wlUoqcSxTlzwIv9I+lFRkVd2moZ1XxoRaTE+1VSS3qY7WCU57V73Lj2KDfMV2WwZcij1R
SSQ27S/rzI2x0yCsndp//u+6jn0lKaMaFVOPO7QzgZzYEZKKKr12o7MdTo7HNus4+JolUmoLZCpT
osAWnB/fQavnCxUPyImpOjFztxPi3KTZ4XnyKBHVzytJBGIDXQExuhGaVt8/6fk0bsLCJ878q9wn
+o9ggaviD7kF56JNt2tQYeH7nf0vLd7WAFrYf41w/ZsX8iKK6LM64JxCYDmYGoQIkFaSNe5de0ST
DxDnUx25XRutxqYSwIgONIectBiwd6eq2QWlAq/Avr94K4HW4vz3sURKeMxeXL9kzxMuJMOx1lkO
16F8CCZbUsKsWYd37NA80O1o05VyFfAHWXg1Ysa71rRX42eCCfauHSAlpHtUdR8yk/bupoLt9F/y
lxQIqrjoXvs/6DhScL/05qjmYGjV5GgYUz/u1+t7WDpOUVuPQBhOJSAUqyn/pFErG0pCeFhQnMw0
e3owieCOzVp5clh3EPZDg39UmLh4sA9OSqNYA1YShLq9gyjlf2gq4uxTcwM3qJ+IjrbBclJmeQ2G
z5aSDV9CKVaHBynuTvjtE6lQ+GVLJ6XCmLpZEykjOIGOOzwUKE2rVV1Sdxe34BNwS9PCZB9SYgOF
Ty5J0T/30+i+G8DXfusEtFtk1dbiYQtNJXW1sS9lSdXyed1ssQkB0WHl+rvOusNSr4+qkpvzrpq4
BnsB5Omcu6NqyqR0MeiD0wSOwSZvZ2jVcmYTWQM8gGvFZT2R6Qg7vcAzxLRQhokSlbXzzCVDvf9K
IOjCTqdv/ULIoQLtTKW7nhW+Jwe256ekJkkaTnnj/jR9ZYxW/d4vm7pcZZTfapuj8HH7/rx5lmIQ
edQjrUhnFoMXGRAGcuuvRYeVOkGf14FkMmSimPaocstP4GMf5kybzMCeZrauN1cEGJEtVwz5AMa1
fMfKFcjZ4FUFb/3Blv3Dhbr+DEC/aDBSnmvPymFyp6ZrjDj+WpN2uJIjXy5NfbS4C1qrkkiAuX8F
fJX8et5guNanp4JTxOzi/obLX/9O4IPlCCHeuKtiRfSdECJ/qC64yLvGy8yMIxC20C5a0TKCCNR6
E99/5YmVS6p0DjzDn8TJEZ6c6JdyBh1TUOh9U7mMOpQjbF8bOHeaQcUQfV7e0EWqN71P8c2Xbh2z
c16MQ2o3uTzPZHfDV3ZObhjdbTKP4/XwgPJAS2VbCLXO3YQmznoPx3XxwQeHSzEWBmuKNBYBAYDP
uQW8xv+ZEaAibcDv8rBIp1f/Rx+gq2/DmEwIY/x7dzP2yVeV7ih+kz/NbvfguVfHiEWk6+eD3ef+
ilnmLqHF82Df4/7FHk+dvaJY94jUfmUibnms5+NLzt6s5sYCiGrSeIPmgXEWfM4Zj6Kmsmco1XOl
jxqadNMjqZB+Tz9NjA3eSoSoCGuICB5NNro5tNssqFVqut9/GjGmqwDqlzYyHLp3Qy5BXQvDyS+F
sy2CbqQGao01nPRC3Xyjbb7dGegE1ZbAJ3u17jSOMOcEZRjO9MPOYLFbNW227/qezwCBdeAJ3N34
Zim++SesZv+zlsLUBCI2I26CoTOrtHOo6Mbxs7m4BGDc5I/CVstYEISbl908QZeilX8aN27nJw8W
Krj5cq87xoeKamVjiRQ/vxyfFloqJXlO1GuvpFDFWBY9ABR3hm7uwVitMYJ2vwPgI8fAfe6qFQG3
D5C0uGskxPBcU7g/fmto0t8All7l3sjSlm+7pXeT56VFcKkuKA0+L7PIVKnc2jJ7+ah5Le8xFCwY
NqivFt3GiwH88Gtxtc7JLP3vp2vpr8fZ7KoA6VdKtoPE2fDix9tThetE7CcdnGdEbRU2YbjHWH8f
Jlv23agaRKReask1j7RqWKwZkG8RA2wbsubAshw5VC1Ixn1F9yeY/xbfdNJXRv9LcQJtLa2ewP0/
t7F2crLni20o2PSfueIfH/QE4wA/a840E/rrZcC6QS0v/EVyIz9KDxknM+tgWssmNJLdUfIk+4+F
Ts1uFbNJLGy6oKXtywbaXZb9XFkMUWx2nMpNFZfVlNHYusateLjbo5JKwQ3+paC/DIo3CgR9lHcW
Af11KLNrmzpR1DMs1pym0zysNlkJe0EC2IonYc225bPMMIhYSFLAs8qGSaXI3u6YBphx6sLq9Ved
gMg3U6YqGNAOtINUe8/3a46ChSsGPB79FEbwpiwHmmryD+lkjALzwRHiiMg6GGOfxCIncat3EmtQ
1rzxNYW0fyLUkB+lBcxZOD6/1EKrMwyvTu1eKeqbgPxgiGGHrRAwycVnQauXOw/TPxCSYa9qr2Xz
dG9FDviWR39PIBelAV5gjry94D5En39OS50Fn3v1TrUzFmjRiqCK5X7HATBha7BHHwGUt0VRNY7W
1vO1+axW2239xT0Q1/TR3olnYAN4BKaDfXcUdiVfyLHzJnGk4ocNGdoBdnvzJ601Yz0SPcOh9TxQ
GQce13NLtW7+UbgCP0kIskT0PiwVVSUL6EAb4GMHQUjpzdraNmnW6zoPf0trj62rJZgZIiKEgiFb
Mfzna23Qs5QESosEp3X2obA7pEB/0VtCMvnBHwaA8vZPKsv4kZrRjpA/MbEJq/EJknOolqdhHBDJ
XotST0/Lz0quKC91hMnuqxBIElfl58GDAgyvDpf/W9/xNM6aCKOuAnHcVBC/sbjqtBmjHzpOFX2o
i6wlwm1mxaEq8v+wEPIV1WJR1C0f1RUfvHFBedfZQTgATN8KwG/KakzsXSu4uJXipcDxsW8ubaUm
wPiifzIPeqsSYO4YHXvXuOgwLCIW+mZR47G+f22zsZs4B18Vmh/nXfVvwyf79Zt/wl1erfBVtB0N
So8aEEF5P1y0Dlxdl6rHvHIEjB6AFctpBJqXkStyupkbGDCS/0ptlgfWtLsSSAv3YW0L6nZnA114
lMRgcyxPZxdC4zH27XeOZC5q4UMai9e42m7rMUg99rSbKcXupTj+KrgZmi/yUlQ4xk+OMJz2kYH1
fJAAAtmy4lSJ3wUV90Ea4fZoNo57k8PeorW7zlYs/dz2Vy6Oji2UdUDUy2QAGvOc5lf+XGYA2gXQ
+6k0/QbZxMq7EJQedAw9vjplQ9fw/YTGA0Ujn3QWZ4HXgLWOw5MY82WJunvTTW9cqbBRmToRk2Oa
yKMWNJaLE0gm+4o6q7omIA+hHf2jNP1QSpguXq+Fz08DqsYaCinVZcwxl6D1TZvG8RHHHwbK7AJN
JShelOLqQVp0SqKCS5NjjYJim7+m1j+njpT0Ch24FmmZE9BvDnW/GFu+BPB0eMhhrWzfI6cUr1Ct
Y+p1XsWT0Q1SL9zBGyYWHA2jHOsE43Ce9UfutacQkMOFA2p1tyqi7yYtBxDRBfO3d6FeuDxF9LfJ
pW+A96JmlWwkI3O1VKC3e24cqnbgwFHUJaddMz15YXbttsXke/uh/lVNFClLfpbjK9TAZ44W6T/T
pakoWzzU/G2AXaLCWv7oQFA3I17mZ1XkbNjq3Qf8kaU8wTpZGwvZHIFT9absxYI00n6XcZdM9R1R
Uc2TLZ9DymwFA025c07qZe4Nkg7JPhXD3OoVh6rgrhF8TKtUBudy1qZtHJAEm/8hHy3u0AVxVEqw
VDTEKw3jxeSFlPE5suBn/fJCnnTbdetHGsEdScSqnPHI8Y5XEkC49vn7rI9cY1q7RKD2z9SBZ34X
TAJkxMmfoD24xaczl7qVx1BAGGMATZ9Dy1O2hNZy1gc3OCsBUsnZCwDhzg4iQSshCbi6Fj9D1UMi
a6f2YVGvelZjrWohYrVrNMtKndBoDDWGie34cb6U90q72OsRkvrUsV4ewyD5e3n7CFvHvj/dq3Zf
dWeMbULfU2vYT/DlOaZ/y9a5FUbPi7ptTzcFEazwAaJ7XB21Q4fP+KcdW4joe81BrXR679UmbDMI
+POGDX4MrCEob+Xlpqg2Jiy93+oTpuwg4kE2XLtugiSGRli8aa+ylxFTikRQcOkt3bCCtSupSu2B
w5mKzdHERmnFgyUt3AtaFYfzfGq7QOppd46iC4+VGwmdm2scwy0SiAP8xscI99eFrw7wp8eVxgeT
zV4FL1jfAgpksAwYoWfHvHMFl3JKdke8hbiQ9WTD0qJNzwQKuItDtKdxqZcR5Na6Yxz0raglFsSl
Inph0JUpLSwS0A9cgVFNKWaU0QfgUIacEw6qMMzMf1sLUi2RlA9dtDMCFQD82CLqIXAJqYZPBEGm
zjzJSEjCrmspVj9zxgDBVyqDmKdJ/jsfw0oh2jVZwCJsEfHT8THtKlSorit6cLZJ9vlsq8YFdAgj
nt4Su6amnIGdDnJJK9C+E7Sf09oynXlQQiYlJAqt2BI+nwIXQa+QD3TmBSXw3wbtlx2LV0sfItRV
lwYBgg83bBJ2lTYR7GDXQjyTu7Gbj8ehRHAsVtn2hz9Fcv3pydDKdFVmvUKmXJyLzwXsgMKA5Vws
/j9uX0dGW3WwjGpPggo6UJCUPN4miyjnyLvMsoyrrBxx4SPjy5LUZ4gcd4idPJQhsoJQSUbJKR5q
ZWvbduZK/DpfJK4m0ObPmmzbniJvZS/VS+XvC5fGKKTKPxffBv6us1hXn05XBhXEXcUUDT/DJUvc
hvyxVLmCPNXlH9yXoORq1Qjjt+zLpH+dtL98D6x5Hc5Yr0VvYr8KXrlohCr5IxBaAFT5vqoswr20
E14dOSjrYdBRNOIm4nJjfFo01+m/kB+DnzyKjAY3gJArOsTeqLndxkYOs5Hp8tZ/itHiCXLP8vlD
jfkKISNMncV8NyF20PCcJ/8wzkktcPSoVcYaNQylNMAUKcfit6Gqbd/One7oL3VwmKtWcfGNsO/F
9AZP01aVUgGNDcyJA00FtKJtswAYPZ/nTAXMwPBZKglfAS/uxeWhSS25Bo3oHYj5O8MTTyPdwKNG
6d314GYC8QwunR/+LVxpU7C7Zwd48XSpUsBClMNGhk9Dq/H4DNMagFhC5bX3fHMGQYnOq8MsTl5+
bue0yQPZiIFAqqz+XBWWQMQ6Fdph0rBVq8aB8aep85ccCnFtwUrFBIJJl9PsM60b5RiO4eMfn2cT
RUoJ8fjtm9SK5ekFdY5ueBRTiCV6M+t7jnIW6nnb4JwBJITC0ppbAQ2nGoW5TpGqc6YciXb5UAw7
s3ZUV0SRkdhkWxL5WqaEIHbMx7FJ5MK1nObE4R6bnfFl5NDI2UD/TxkYNIj1QjPs84uDzhm2BiJn
J8gRE5yad73CPVwAuIAaZJ6r7GKpN5m3Ev4BjM9pWRsRFPrD4kSUUQZ+UfBVg3LIn8ubHRMuPldB
H91qaEpJvrBeZRtiApbmt7s8jaKlqnmobX0jcsEXxAHrlKvWPayEt4C7WCL09KKdVzIx3GJNbDUS
wouK/tCwBRiH2+gPSbpfSIEdZ8D2kA42VDKNTzTnaJyn7brxkjzeqmHuhkAmjdxqI7J/ENMW2QuA
E/oRQNKD4Ba8L386pXD1V33ltQ5zC+Y6TJUr1SnZY21MWRmX1JG+h9sFYLo/J18w72w7JCU5WpYu
fon1s6rnA16SAgh+c/+fMa+A/Ep2xYGAHCNk7GUSEDogFsv4xGRtb5ZKpYwss5eLuZoJJznbz6SY
eMtmImDLwJeJrnLgoG5TV6GYOtvjt13uH6M9sB8W9272d/T9TsCk4gnlUCKmc1vrxtDJpBTAjfby
Uzkxiu58jan199uh1OKCKLZecRNfoEzmxlwpnidIK6cgWLxaGodqNPCC8lYDDxqTNyd+xXIvK2I2
lcJwOzcF59hCkF4dOq7syL4dFQX8kxo2PjwzO4x5gJ/hJ7ZjgDvkzy9pLuDRrapnvucLKapzozpE
XKbhkt/k8d7VNiAzG/DySOeNuG3p/I9B2eukuaNFHB4jhZV1qtrksABuwDNkH9iOGuVn0M93SoAK
StbaAqLGxdjE1yip/W8DAuuRd2ITVdPzC0U9ypHZqEBXDMp97InoG7VN4buJqbx05TAm4oh1xSrG
f9pQ5uU33HVl4olML1BIpz8ec1nplQdDYhhjsU1W5Mx9r6+KLW2xAA6zRdJbaIX7kAPeVvysEkHg
FgIYLiUUmjXqCA1GuAoQSMikeQU/RtoiyR9NXBOV9dtMiDd04fO6oHGiAgtW/BSuSAd67ZZE4Emb
RRLkSlnreAE6F5BxS5eJ5buH59w/FDYmCU8jlhTi5k2HPL/VOjZWkcQTRk2IowrrIv1r98ngQKD3
CAqYusf4ihO/qCjzNolHhBM89YMN1nSSg10+IQ4DsVBfsyVN2mFoYIIDqNESWGzlDLlRdw7qiiOE
mihdX1NA4nbNMKeGiYuXk6fn2iyijrhvROSbJyyuSCGGgfYTzRlsGFVrONdCBbROuYxxpO3LVInL
4oBhNgdPu+vUEEdN3lHaquFB67fV3MCJYwFe25cnGPe5xvWdrmgYopIiB3JLVnCPAQ8snADrJWI9
GjXvMjmJBX2JTD8Fb0Kkl5FnXjh5r/nS7KoE4ZxGb5HnD+aYKqHCAUimNHZAS78U8K3Mx6tL2PWK
SerpPtYqteigDZMNa1t8mrjx2HsBNk1b6juH8h9z/mEWR/dLd/tbiwbcwJG9Jv1Beyr0jJfQqwHu
dn7QfnqKPYw/sd4MX+vwgVX0ZL4tpUQed2SBSYwc+D8bfrAdl97wWOXy3xIb2ML0U0T213AZMXGJ
9MlYAej2XKiWs4poXZmGUUUK0Co/GVE8c/CsGGKR8zP0ANveD+JbwkGgyNl+qrklWl/FaAaEqc/e
b2qwYj+3jrPiQTCq/1FQJqLLLaS7q03T5h4GTyTfwjIkF1OzkGirZyWQSg6TVW5po19l5YsLLfYr
ssO9WuTWrA5ueGxpKX33o1OaKIivKFSJZiCta5Vie0YUqLrxmHIYURUMqq4fBml9hhkvEAg9MuAc
AFaZ1dqRTI1PkEUdm67ER2YMRinM5UW80dtVJqzxf2kN+vjoPsRaRSpYCT1GKnY8Gpv4Y2dB6ipi
FUI8D44XUCJGYotKuMwssWj8IF4A/L/fWxFJ71cSBw1rYKItnN8Zx0vkOCmLl+A3X7/1L3XR9WH2
qQQ0wINxIxIJRUM1VsoDfSOPypTRYWsBgHmSDbhbfunMGR3TGcC0zjnxTtGfqFKT4NHZbNcJOybM
W98ty3H0NwHVI+k0TsedHR6y6bxDPEMLoMQWfsCdGanr2+qyY65RzlyVO25aMCF9irNQGQVDFfy5
c5QT1La4jLwwWyfPxM8AxQJZDrQaAFzH87DOeGG9ZY8yBm+yrz6xZjO38JvfLvpgXHHBOTyoiF0Q
ozNlTfYZJ3of0KJV2G6v0U8hjYl9Y8qvz99m2pioIbFg/dRK4ieGpYcEyBooVWYxIR7c3e1ijk/L
zU5xmRdAibaMoAAG3txn+Pb6/KHteH40NBBXoVuqqmd1EZ64JHKPCuy4+qBCgH8QkSEHD0lnEBc3
lr65ya2D5jiRFQVKsE22wyrZHtg5AviO6uLkypo6DXa2hAFrwHYzKywnRJsX7vZM1snH7v1cTURw
FSrCsAnHPhCWqxZxR4FWPuRub3ErVmvPm0buLn+4x9dhee+AGU5wJ57vAxp/3p4biOLWGzB2mD+F
qmORVJTmONivJKqWnyxS1xwDE+QwsKF68XyzPI1bqA7OHYm0gm4tDaZqv3r4eJb7QpAt4qT66EJU
PpCLpGhRbK6mmXDFMabFIbZfnGMFGq4B9AgPIVRckI7s6cVvU8pM6zXz8vYiNYY5yXABW9lCmqWx
ioH6jTrcCfZHhQ53wCBgB4Aoc1j1qYcBVnUf1sdMkAgTfg6GvvpzvfLPGHrQuSRYca4Vb2wWw11v
9pz5+iPgb7VNOEZYpi5P194YvnIegIFjLhFoPTKll9/rVbosWb940/OQu5yXd9j8rDdh28OREQ2i
BMDg1hwMpsCGlq2SGLPxCogfCbgd8yjIuTUub+0/3oiMYpoTMBWfRqwAmbCqFWnkxt1oNqD0lHB0
FZbRGnNHVHal6XniKxZLrWN/c+0h6uAaeTfjW1vST4BWpoEEEjBYsVJTLzp2eitACBqRxECbPRMS
S8Z37r/pm96nl52Hs6lHa0h2Sp1khX0zokPpaCOw5Z996C13tUsGvhoPIkKV/wZqXOCRE2dJcceN
WSYXv/Z+BfeEhEiEZl7VoDrg+CxNVD9R/9nVifmQ5TeKUSYml8Z2eNvewXTUNYKenHHz9DCYL9LH
R8znyztfwjnHvuGMGtkwHWK/i/77Wf62VypMkDsq5us87qashJZvLbPdAufNfikRr35JWPlSrN9J
8bofaNbV+KpO+RH/BWSKnqo5Kpm/ZAmayIIhgg9Z9546us+3eaMVUxTFUirvXjMunBqR7fSqYgfK
lm3PC+6fpkFcvzKeX0ICLeg9cYoBOgAIVV9WMgz3wjK8daCkqT1zU7uH8GmHwdwa7b19HmES3ps5
kwjdijRqOEEISvVxUkxtFI02k1D137Nydm8fbzt9l4DQo3L1QxrKwwXVfjl0kAepz0y887y2LAN1
JdNoGZLOJGwm8t76j1F2TS5iMoNYVZgpSdqF6kLmIEqrySVmzaZL3jEFSDJoxxtVmKwMJ2tBGUwR
F/VKKIhj6K5cWz/hvJRSCh3waItNYffGX+KU2vDuHU7MueJ7+3rFVsXSnWvJ4dcm3o83sVLpB4N6
DaW1FDaVgyOhGg2wbK0//+ftTPiR2R6xMLMbw+YuLREVY/iZUbfq5dslkhI5KexDYEBiBAktxQF7
CdSuMHMDu2hGC+8xNj9ZNSGP7ha5Ix+Ok9ayzOqCUv6bzGxtXnIVNMhVeMzj7mBTXwATDh5xdcsB
sxN3GBs+UPfe1tlqd66uTOQxNbt4HP9UyvZvkeAB3A6E17wvBJi7kkTYDl9xBDiC3OPdvII+0fsH
DgjbmTRiOcwXNOJjKEMmrfzdpiuTPBRIPlD5s3ruQ0xbd8nv6NE2KNjs+qx4aHniw9xpHsnfJpCQ
VHZDRC8rBlC6jOj2fqyXhmdukS1fmK4iFQiS6pTNbImspolEaIXE88NWsEkAPSpv9nd835xOucQw
2jMXmxjo5HUsY7ZZjj+MiZK2SvnJlwJYdeg3qfsU/UTfNNi4Nu8hb9hVIWFtHPnFE0ilxQdSIXmc
MCZQldXSZuGeeumuaEA5fQCm74dWHyWuJsT0KMjk55xBg+HWX2Cvg4pXBUvhi7HLrdUJaqu6cqsU
JDGcKmY8PmbSa/jNncesqvlbnP8tdqHW4PTG8+5V7UER+JFQSz9VbMxWOw8sYp4Wc8Ci9Nf+fELg
8rB30AErcBll4siT+He+IvvORO/xUFRPgJc7YjwrDPUQS0T03PSHJiE55/8+NDVnB08TkfLlZcSy
+20VyzMmMTbVt68oAjAdUXscTSSfdDAmrTUffuJbpnLqbnvMTjWA76iFN/gwW3TjDAe1LNxDP3ed
df4hYzI9oXVSRzKnGzVX6Fkn30fesfiQU/761OpOkz3KGEqHHV17S6jio1ryRQNpqXXuU0+Tddfc
98ZZx4GbDH35IpZBlYAcQwY4DRQ2E1kcmjAOkDTKgNbSZnEhNLyAyIgwM/XIlzXcoq03EBNONT6p
1KIt6ZHebLrAyEn1jBZ6kRKAtj4HtTGn8sgxeJXAMrEH0fp5+PrqlMnq+xJu3bSIDTCOu/8Ckcyt
0sZJcMfp9aauizBN0Sj/KtBY5aiALVVFVSmyTFUmM6kb1tAik+XqU0iGcxw6/V33gqfTJChsa+cH
jrcwm/fCdKkLSaXN66JMLI8qqWGvzHJe3ngvGW3hj6EAMtwMJEajIvSh+Es5ygGQMU4SwXLIFX3n
IO42qHD1ffRZJr7cYAvkYjKdDHzBWPeRS7cAi311IxGd0uakNXNQEnF1DVAJ6oPPHuuqmhx2bkOM
DaKRAOYwgJp+Ggx8BfWKsZ6BOwaLum85m2WPsnuGOw75I1K3pd+Upx97W7iR0LkrfDnIeESjS/vX
jKn+2KGLUs8ozFvdMGew4M+mVObjB/YHbNBzJDpyV1jrcybU/S6jPxqZoOIEEj8vNNBtOezktbZZ
8JwicpKKq/nuf6buAJp5ievtaRkwwTuvntQp0/XlDvicr4iyJmDsCb2Vo/itkcX8vQCC9U0bHCGK
skD/ym7EfuXjmmV6OUcDh0zw2Uag69RPvcqz7hzESQxJeYFCVnFrN0MRO036t2YQvsxaq9jj55gZ
91ThBSzwfOQBiZQhTY3DgevepK32pItxHqi1DCa/3/UmGUpKNTtvX0cayp0nEEVBlb8xoGm2R5dY
irVKAhcpoOgb8Lj1NcsF2M7vmxm6mLF+hxg9JmMOc1ZSy086SUcT9S/kzKO/UaHByeDFugUxqKbG
bD6yQucnvpuyUYiiOtUxNErTQcd/2Kq6lKPW9/GBOHyR5sC8GV3YwHYpjVgyeqLJCeSCVVhg3r9l
cIdKJmAhtasd4w3Bn71Nvt5KOD9Q+TB68dXdjIhaZ78h8Q0zKl0wEoFyeQejF/DPPyosChFLAPRK
cTV4GVpnWAYK78Sn0lzDZR2368iBfTFK3riKbXLfeMDF7Fkylsn18M7iEpOmSOskOiA1w+WHwjdc
wCSMe/73lWdNxMuDYYL8z3xObo+91e4QZ1We+9ANbgYMoaeuHIpFTUaE04ICdF1pI103Rks5Zwci
uf0PsHTeGKrQmXzg6BDAttGN/S9sHUWFZ9dqkkGQnTfTqdy4ImdHfjpZefXdJ/LBoRK37jnkWBS5
OFcEKrrZUfrrW/B02GK8act82wASzogEsMuYs5ty0yvYq5mHnpWs/RWBXkMZwbQ5MrVaAwnW67bQ
znX0H4IfJsf94XImJThONHK0v5usEwOhmUEdRul4ftAD+rXyIcGRXlY8prLUFd/Ely5vJdQBVQUx
FqBj0pHxS5VniT0iNFOCo0J7LEJ67fYU/RxY3ywqVthQiRZQdLgOeB6CvGcVjiv4+NgzUl0dnRWU
a6P3DBtPA0c93y8IPIryz3vYxCdDqbmZhZVloZxGo1PzZsS036gDAAJJZWbK3rV142NgNUloV+sC
mG8c0Git168cXYMwia7mvmvbdTDMugiYbDUz/xgoie6JpiX8X6crwLK6GR6/LckDoT4gwe6tw9wH
G2iWRwYHEVsrwO2w631XLIr2AvDyQjRvZagWBX6IVoB3ODH5GLUmTalPqpnC/G9KoD252AzAPyQX
Rc4eP/F0W4nNyRli/cdbR6+NxZIYCGEw7i2o+Wj6FhpVVGPtLKk/maD4Lxpm9ml59p1+gkAENmdQ
07x0a8IK32NGqerdHmmThrdiU+arPWlH+FCdhpyRgZ7dwAAGcs4zSgKNk5YzKAa1ssO+8HR1cTtz
tMQN1HXG3FdQIOolzmxaoY+d0lOqyNuxe6XCU1fSjxRcZoDgeX6NnUufg1MkNmLt7a4+KJdcHj90
EW0gpTThMvxPX2ixphekPUYMIyQ16ZrwoInwpcshlVv43S7OTCcyPV5EJPDCVpH40BF1zeR9156f
uSO6wiEkZDu1jQzl4A9ggFHm+BTntXubjfhuvEFsPxLeI5FAbOh1e/EEBqDi3gWSqp676RJptpRn
rnPJaMlbHDNs+O7G+NSR679rf21sZIm//teuxGXhLfTkQo7zNaQWCLd8ZRPbDWZEzwi47MGUrJka
JQXi5VbT/NruV+v4HkLMShOjCzURHwVq4qhx+7Uj3uEzGZ2+qAEw7XpS3QugBmrixbenmhqqyylL
EKesKBjCnONhN1Dz9fkM0b2TyuRUZ1jS3uzsjsUwNV47WRABNmIaPSxn+BdALuqCnXpzat6YNIdG
5rpXe20IdEoDCNkAIrM/JH6usl92F7T27Ow34MzsB3+IofNPSganunaEJiosOjmcyBsBiNfj2AIf
wirCqU0RXsXZNVVRZkj/dWmg6Nksg82VHuBn5dv9A4oZ3OldU6HlJfYdTKL3kfpCTuquIpZcuaAz
+mYzbJrDyFeB8U7DFBjMED/dqSW8D7sOymS0UQpVzvwT/0w/dGLZpyzeJy9g/n2pRvazvN6LzxE4
TJf7QCH5ez8hv7or7Mt02e8WCBY0EjvkZfO9l5r3EhB7aOXjB87r5B7c4SFl2PBBd8BFOi5p0S/U
AAN4MnoflMgurq0zG9EIoMg3ex/muTShvgjPa46ACjCxNOFsZgiePI4CEcbRgYe1ktVx8RrZkkFp
WLhESQpJGAptKM04PMBa+Aq+rkOsSLX8BJDV+ckskCXCpF6MH2tjth6VNOWqkrgX2eJMEx7bW0vW
X0eaNvT9/LnpCic+CnyG+cIVwcN81OKW29UDlblVj15td7n4damoOle8bxbPTJRGy5tRv5H1p6Tx
KmPRBI+IyG8w1YYMme4zskOQ6nN8cyVbTLpKAq8URvh/mW+WR6WBo1x3EzHNFEEYCKkNh2fo0PQV
GQumFHXaBL7n1asLa7p2+pFOFUaHcOR632TK4xhoypyal0xu0jNbWr2ZDrM5S7W0H0VuwaBsjfqW
nAbRFCSK3i+N87eJCskoviS2fmtVkq65uXLaBb/6Sc9TZz6SzTJbrHTLnB1yykEjf8JKb2U7Ck8M
F2ITv18mMyuJsWg6cO5gUOczpLvLNYJQ+rHlSFbKAedMV+LyrVI7BRuFokvrsbLVndwSZQ4AFD4H
qbtFZPQVkS2y4JKsaO9S4nCb6q0Pr64O+qxj+yDeaM2D7MJVHhmfSA00kWN8VphYL2cPZHpf7T9o
SuCad5HOsJtG6x8F888eEV3ISn/2tyvGvaRfsbQrNzhymagFCtCzexCf6aUfmaFPcNvRBFIXxqDW
1gvfEnzKreITUWYzkJplqXUcMm0VW78qedbg3qItSJHxEnEfA8zUoT2WA69phRPHXYIVi9UJnbi/
M1EbceUcydobDfjBfR2Z/D+fRhVHylhVcrOLw+2+rb2tay2826hU9BUtqDqS9a+HdyLCZ/PW221l
i27iuN33rA+Mutx9WNKoEVnsm9xKljd1pjG4ZePd+4uHx3jLy70dTkrWyEjca+1vbgL84qifCtcM
28ZkmwD22OPIWmepS4ewowud0Ze/8XewAHmfyj+xyXHzVR8WpEaGKz6Y1TNExVbM7+eAGTfg6P0G
jXBUdnzlFw3G4m0C7amyHooEHwuBtNwYZkZJn+Wnhv9zNjYRJMYK/YrLhLI9YJ6xtbehBdogahRU
VlvqtF9uksaQv0sjrXQRoSR/7f9OaccM4ul4snrz3o+ijqX12isaAsaDpx7wzCmufL3Yq/ql6Lxg
BZvqZgTKx2U4i5syY7MxZnLfiPOZaoD9Hyx9BqN9gc7s6wuWBveAhXXBV5P/xa/63zYuK/YVNFsa
j1ZY0UmK0STE+sGg5C1GItB6QfUgT5bGOHNHiz/sTUIewgt18gQPva9nHjw8vseEt8uMdNw8XhjW
7AXCD/RcI4h6HE8Ny4KC0HMrhvPTDspTUufWrYK57LEYVloMiLiEsE+LBWYX6e3Zsp3AMtRCBdGz
0/X8W4zgcTjjVA1z9KVkSNw2Q+5bO01IEEYC+KKF7KR0SevbL/dIPYy4Tdp1R1q2CX7MDN20d4Sj
5j2d3Ee5G04dq7qaYSNadAA7llGLeyWWSA6gWGPuk2/t765j7nk+Llp+kTvLlL7GZK0Zlk9R551B
ponWreAqE9TF/UMO/4Y7QGGwLXHzN1OIX7hU/i5IwrzOekMMZvyjKK+iWrk6pS7WnMV0/NkikZCB
ip+E/Nu+ezWyIORTe79wIbCUsWkurwGDMYLf9o+cIrqdxL6b2T3dyGEcTAgtzFDB3BqM84c9RYHv
B1LoLDIzwZ1pQWllSW7xR1RK7+OCqCjcdBHIMKLj+zWXO09hO4Ucuktiqse2DBKMOPx97+vOn+QI
Qd7D3/rMX42PPI3Gmj5UOQW8cEqNwLeJv+37arB85BNQyLxLW5TKkOy4VkDHs6XAkI+wqO1I41UW
U7y1AEnYNWJzDA6Q/2rXwuD41uky9M5FNeQoAjX5bIEkSrzKjxrR5TvmP8jq29Lv/I3XOaZogiVQ
iJiwmDc3U1NdTM36l9hM2YY8+VWUoo+8BERqX4yYAiEMXGxFkOcnEDpclQQOMTMahyZZoPqWFDx8
tt44SFFxeIzu+9Z8H8YMahYwxcZpichqZFhZOiYRNhWgP9Gv1g5cnVjvvSN+LeoQQqCaMhrosji3
d7j+cVlfNVuQ6UF1D9nEvrWfGkuu56sEynO+FW3zBVgybMadB5Eky2qICrNwkUvjHPhgIgLt+9ZO
9nnPZRvL/sgY+VqrO8JCP35VLUlcmJrvMLorb3SP2Om1A/NwQ+yFJvIrZmGBnATcAC7po150c9//
Z867Mz1/PBkUBMnZOP3viGhEpESptXhz57gWo4DN1os9uWvcMAu9CzTERkxMjx1b8HwmC5UDizsH
SrBVkKx8C6gTYAQORG6i5b/0ITcUjeShfUsjqDb1+KhL3u6XDjKVXtqxFtNsDR8pVGPWTdCzWw+r
YJFOw8exhveN3w+C65kwydesrpfJqtHXva9iE7lCtz8v61aKBHnUvIkYi5QRLf4wa0jiOHjGZRis
N00XvZuhIThne5OxadFMQLxql0u0BD92PHtsTaKuNoMiZffvC8Fwi0rA5WZvzWPyDz4go29cQoM8
bft7jWDMt1Yvih0zqIGhZv5OTpCqWLkQzdCOZjRWzcciMODnCW8vuYBbQ7PkUW1f2MmRbq34QTik
wCNl8RXk/fPaapX9Hm1nUNF2MzUEWUwpxi9iQZbFwOwTyYit6eUU5RhirOOZn2SqRATzBr7ALM/Y
vNFGKK7hC75hHVfnswbRQWHrL/hxiY8FwUP/a4ZkwXZ5KowWpggDIs+fCkW9tKlc6uuF7tkfiP11
iaw5VE0cQ5YpL7AtH4KnUm6PqV+3FzM39io4ybA8BYHIR4y+q0CpT2t4Il9kGpHlZhAG/5IiQ8xb
FguWJJTgS/1jtx8W4o2nmIuVVNOIn+iHQ//IxSc5pSMCP2eu+O7km0UZItftHplbc/QlEmZlClJl
vbV56vlm2k/U5Y7rO8rhlC/ty/Uw5htQDlHHsY8WjSyYijFFEOaChn7BK7KXff+Le+RbB3Q0fe/X
nJ5NQT72mTn3dcEJk2Lj+yFtnvWgoTjpaz842OW3xUOtKN9AJRhc/qYKpDrOIQpnFG7tofqFQ90E
AApxljzZM2mOD9xEVrYxyASanurzcZzLfhglyfThlRJvL8xmSVbbnj+AZAdIDSHpaaAcsRHQ6l54
COCNkeC3bGZxbTBI4pbFDBuWv6aNL0LpYnAsxKOPfkI2bAuJxej7XkAKJbKHRWDi6NABM9Zm5+68
aaRg3hUzJG4imK/IGSN1FtuB9nAgo2bWS8qdAOAfQ9tsI35S/jcA2xIsPRrWJzMiIdXdmf/0sdkr
pu7pmqpNIjOCOkf4cMRU2n/zhgZzChK/aRGClkSLHD3RYR201ijVCkQElP2TtzGZ/bfCcWXNtXiH
e2QqMJ4EN44GGNQLWiO+7/RjtX/F3HGW/0m3cayDyGud/EEFMfHzyqm654+oRMjfXtO9sdSLp7wE
4LcWg2cXgJsKK+vhupGAwu342y9fJa0BCVt0i/8DfbH5BD9VtL6uk5CXKlLXHj3vufT31aQ/CbqX
gcZD9RMFvhiXjXDrwpIiYZYhmnWr2yd1Wb39Vdjer/qgQb4AY71xOctdm4hFf62UFNj0wlrec+AZ
7178ETMdHhPItDacULTnzn1aC1g5M4pvS6ckcznMdPU9jIox9jS9YKL56CKXYLImxCPeU3zFws6p
Uu13gQUDGSK1SRYcdrvQm5t7kieTxkS5YM6LHFzGRZinEDWRhGc2Cl7cla2axr9lqkRaU9w0O5lu
utCf7pCx5ARuyxYf7fu0q15ae77TJVLLXC34AjRzND+liv2ASFFF5TzbFmkA9IN1d3btuxwbHjrU
aMLFJ88Xtlw3FCdt/NrUSvQs9IHvZifbQl9sKzTFhyxT4EgIkBDtNdNam39ttqvtah/iLFWwIOHk
qB+HhahTdFM2MvcaRlLKV1dWGyuWZbkDNkPHXzD4/3SbokX/Oeczsgjw8XK4XiPiQtgARvklP8Mb
vX1kdE4khS/XLKyebJW4Isqf7OAVq5It9zpQXifYeWKeRNUkbRsOoX6/hiGXWiSR6IKvEZo9vSPF
Mm2IVmOHWonoYR9hX8gGGgqpamyqD8lWdJNznoWlZltpmM9bJmPAo4+NUat1y2Gbmv+rXXB6c2Q6
jkgYscggO/nxVY4JkF4q89uve80pyIYrzhR3NYha5+/xQnh6t5y4qh7wMGDuytpLg5B0/Ln9/u3s
zhJ8+aYN71MOCYIinhkaibWmi8l1lha2XL9BmvtWFtkbz1CPI9A4c9s570lc6cHVvwqYF5GsQyuD
/W6/Q7w1C36WtdhsoYkO0e6Eg5DNE9/ocj99x28pEw/5ARMMZu03F3DnRo7RcBe6E52NqFsI+sUn
CfcvjnNmpHvt+ibCoKrUY5sDyy3n2emYFgNwVu7+1lUlChJKimFVcocN5qif5ss9dzMkrhzOsref
b5gBAIS7wJSKkjXoWibn42L847gyvpQcOV84x8GcaUkNj94dyNv+JTX7TxCRs1K+q/JdgSMqTdA4
7Z5CrTKyB0al71BMiDU8w/zDqhA4TmyUdSNSk5QY1l0EFH1TKuIEpYxM5mUotIZ35PRRkIZau/A6
FN84alXVWf4sDle5idsIb9Zggveqhb+kR1nOyAc6HjsQXU6aacg0gQsihvJISOtl2vHHiHOb1vgX
lOPzuHLRRiguwjZ+apXWvZe7kxtgY4xAfUR1OEF/Y7WjsdLs6APc7m48EJGZUKqF83o+Yb2M4zy4
VMcU/obVv7JhQDt8fb3gj0JD5rZY9XA5mH4PkzqA9cRK4CSJfF1CPBXisBBnQVfktlPvcne8cr7T
B7rIpheKPyWhWVYC+cKxmXsaIZD+3kgOafRmsUgjOS2nkIw6iJDQzIp8kLBdIeu5iRjF9Xp9ToV2
6eHgr+oirqRMJhXOH+XFnCNUtG9gKc3x7bmGrSbGXZlTav+qcuF0+m0EjUsjhGjLHA/LQebt6749
MI2kG0/hQ0DwxubKP6762d32FfSVkvFw4f6J2R36YzxSKLu/iE1yt8T17+TcewUDQGst6X0+jrfu
VEA7vb2K+3+SWccV/7W25wSaEjq44bklk4QO+/nA/r3+t5dBHjoERU7oHe71IaurOiIlGwbW0r7z
jd5zKMjJPTbd0FX91tHh16BoegHhRfCkp+27h7bYEhNshjm5dOMm0lGMfN+E8WYutoQXqYUEZezW
BT+k/xKOqbN03hWZmo57ScD1lZwf3cT5t5JCpAyPftoERqYxzB6otPorS+BRKoZK7l/QSz8IxR8O
uvWCdcPYWktUUrfjcRv4CmPHcdQXFay6CK0oVaIZHkXIFMv7YohmcsHu1qL0sxDMrBW7YET+2x20
2jcJ6SQA+1t+zxGSYgRl6NQCyuKieQ727PFsBdGUm29fHkoV8uaFXn4TtPWMvfmV5Fs38rsA4L9F
CUQt5RqB/iMQTeE5zXLLsNrio75dL+L0ytRYsQnpinzLGyfKzJkutef4zsKDIgr9wFns1pmlFEzl
IBdsIHpA6nOwnkCCUqKZ1JrDmycMMK9pm6znmWnfCqTb9XXwTcDT6248JYg3JKzoZ4c4syjS7aiS
NCLkd2TebTfC4aSmwXp3d3EI2e8rQJ5AXEcwEKxEwzEsmyBTz3nmXvBBDqgRistM1yMhrgzM/yTl
oDnEXt+rSw0ciz3b52jXuYvYawvatJy0K97samVQ/WzqctsZxSaCiD3hF6pM/BtKshQAXwvp1pBz
Dmmk0U6V7PngJ5TQlaWW8irAiQHUI2GJRLiWHIMMbdJSJMetwOM89eMOYJP6kvHs1GUpJaa9YgrR
vGvE47LgiX/wwAPcpT346iIbWNPP2udqxxU9iXMkDWgwseoPauWyaNB26Y/htAGeEHJSsI2LhFxC
YVy0zhBGnf5HgGNSKR7MKnGIjoOlPcdDxXcwqNQnAcRik74Rm3TcmtpOE9Db4gEkp3HhtqPeOlyo
bVhPORygz7+pZ8xaLxpPFx2wFQUYp6VqL8CPNcbQr6XpecytZx84pgHdmEeXQXPf6wBgkP0Qn7Of
Waj82nkTqPq4+lo17HkBXdJopnHl4RIENjlWLgIQWZ/9nyGPIIF7yFUzai/hjXdlrr/1IFW/cl8D
d+zc6IREmD3Dkf4+2DG6CVkYDa8VLukn5pjj2FXomSoLzqOy2V4JT+MGAUGfwX55+4PUPngyJ4WB
gIS0hcskh4aiQ3Y3SN301A5+Y4ujGTf71QAI7D2Cyt9MWCqgph66lIJOy/qSj2WmrINz7Rtfj6tX
o9svZ19QA65vfPoTircVLQg9Pob39lXHIpcyefdAL14qITo+0B2kWSZtwpudWScy/vdpyh2ymcng
zmjAd1JcPgLedUMfMjCFu5UAgV0nAs/bLBy+jII+FMAcTdIrg3pF35HgNzfPEhTkYgjJIAG7I6OV
eDi1sOpsLfcg8CvX2bApnnuy+M0ojgnInEZE6ypH0N+KgP5Pa8EVUV4wxuSXm5C7sHZNEgQJwLIV
EmaJ87okM38I0od9CwNiYlEkSf2jEJvVyFENx8bZJ1ILbt0GfwiyZhIP6B334fJOJr2rEgsN6VOp
CjHeVC81azqWs7IZ9hDzDtSQk2ERzvzQJXGMANFLUTIMf5o5GLKc5GJk8voZj2ouvC0ssKz0NRAe
k0Wwe/wqx6ntUXA5Be9eH2MEMVQoNpWfrk/S99aBR6+wJ8Su5C5XiyxjbsLKl5nkj3IfO8EWD4Rb
AyYSHmODnhIrS+ZFAIqqksgwkLGsvzR3F+6zSeqJoSMAdy27gZXT/piLTHNlONBFUIzLumdJC0ka
deh8UlMqXZwPZXJ9JZbdcAnjIaf7QeC51SKSMFzh+XR4hvQPeM1TA7/F7vgZF9QRFyoAg+4wT68x
FvLcPogBjN6iqehcX/08vovUS0OOazYzpHq+uikAQ7EeZPvNCDvHxpOUpbHaXD7L4uFQo4idvZwh
tk6tl9BMm3sP8vzf+XPlExp2j5yfPEdSYEV7CU8W9LrgP8T/8uc3uASTHkXrJY2WAT2be7irRpnL
UfxJjj3EcIWRUIwd7b4JiMBJ4bEFfkXnr7OL7hPp1tY1D97TW2/tcjP1fBOS2rgOFa8zJffuMvkK
yM5PwARD1vSig/4VATGGnBc7/PEulpJJJL5yCIDge80UtaltjD8UR+ziMl+JdeGsdOUIfcNuB/gQ
FpFDOy6UbB0nXM+GofcYPnPFSl1qT5EtN8BhxrnsY131PctsETWQtrcQM15r+J8uHGtgHeUJUcr6
K74S/j0PV8qFZPsfj40GzmdsjiP9V51e2Zcky0QcP5OwqP/tj4BXJN21qD8cfZpHB9FpaTWfrTsD
0kl9P2nVIkv27JeCSjbJNjmwNDpDUpnR+6dP5JOU6oaVzDZ1beHtnitar69UX7JmhrzoyfRMTPif
Gkr/IoaxaeMaLKTttQvJzXGC23MWTfF82pNmqeYivzWuqZdNIPVpInNnABeydpCvtguSezozpTEE
qDmyOsPYQJGSAg4ZH8fNQc1Q+wj4IzyNaoGZ7LArusAMxbkiYNg8TPE2In6r8RJuYQujEL8xDhxF
VoiYQ9gmkrOKIsj8z1ycOyTeK45EUfRFAlWZUhPCNodtpSueJamxnNhjqUNvPaNg2flzF+Cln2Qo
LeqBwpI0VLZFVRZdMa3CaUdc8cMuLM11tZ3jVrRGPLXi9jnTA9nCYUQ7mgT6P4Ahgjuur+z2cGRn
kViFQyU/+7AlDmVYBOFF88WEofYwqUkEUueEwGoeHpk+B7QC+iiNooMKfWI8r2VZTp78ZKmL3pcT
qCNDz3nWrKUnPakayIePzsVr4t3h7MgIoI12X0D7bE/rOPC1XSQnmAkN13IYqXFFCMh5cE7dMEko
9Chp2O9HRtbt2uDmcTvbXJ2mgl78P9GPzB1B+38L1KJkNmH4UPnEfeBkv5cxJwM5/e4+ZHvzIiyw
qcHfScuOvC9J80nrym4lj77An4VrUqHgZ7c5D9vDC0cRgzT8jb4tlSmqwFlAzTELywOrahkmPYmw
gWwuMSRcwIul7e6x+fK1OIllJVoXoVG5XzQ3lGNaAQ+E07d2Ukn1qdTENxvySRr/cFANfwfWwFdV
YCN4861ZXuvHPcxn84b0m9rQom+fw05WwmVqHiNF3cF914cM/uRIjuWH97Gjci8Dw50737fwMBPs
u4bV/upV5gygRiYSJAupg+KDYI8n0cMyrkiom3/X6qvoQZZN0wQT8dlHB2Rrk2ofaFTTqcDu+1/j
86lnEseu7LDqYI/zJS0uaybDh3q5K6VZQnl7fbRIAfMZxl/33LEcNv6DY6BudM27axUio8rVn1k3
0SJzFRHP/oH5dTVMD5DFRsx5H/yp9i4P9YSfo6pAYDEGwLAoSh4sToQcVfprFCi7LA4QSt8ivRNj
GaAMQu+IUgmXRY089rsnA5Ux5ZRUZ9zwvY4fIHgrw0dGmku1zQdeMQ20t+/sEGDcuNhSzgVfJurF
UkPG+W3Un9IDHYjLwLz/TsJxY27T5HKJu0lFFu8eYWnc2ZfKITCNqXkNwdWaRisc7Po++u08ndS+
hpANe6mq4NOrpagyrj+JEKMqs8YfZQMCBbjDIh09cKC430alNi9HkO3zlScvyW/Z77GUwwrm/slO
x2cCc/iDjpkqvsxr6Q3UP2M/hDjVdnOgE49om/nMy2jVDDDl+j4bpQVJRuLdHrnsbL/R2JG2tuaq
55GAbMWW7ZG4KLkapGGYsY/+EwrPWJXatC6shR9/0XHqwsZ+1AwNQSNBPPzQ0kJnqBFgI0In0Tsn
c8EOKWtlv0RVOZcfFpisZzDcRtkRlMUe7zgPA2auZNpPGT9APyyf9EUkT2b0fQjKxXWgvBpexCq9
qPO57mWE4z9kWYoHcQ3DC3gMItqkrppymC/s9FF/H3BhNKdgfb/aa7RMykuRbxanihsZ13zpnJ2w
O5Iespc5IX/+njgp1qEAHhMfBQOF8D7ax9EqLXsaFneCs4k+KUvmGUEBMwl82oRSgc5ERAvhpx0K
hFSsIF0FbZWarnmwsQ/crjKQKd6SFMyzJ3mMBWgiq5l8/CTN65MiBkq2MMaDh32kJY89CtG4yp94
LYpfdNY7jKXYvRZcGEDwTn6giHaWZGEKY+QrNZ4ZuMYZTK1dE8dNLClOr3dPN7CnFP8tcbD9gUwC
OLiW4yT/Cja82hecTUvJqos2JRh3Ve2rjIDNDGN4EblhOX9ujpYPcs7RGFQkrLY7NReD+OYszy9z
AXQn9qtITfpZpdPwc9XszjW90a9ODAF5MAGHNwvoZDuuVGWUpuRehKIEh1VNbmjZYEyTvhPS6mgw
mMuBrLUzchV/rRyqywPUVe1+hWR8QtIGDgNXLbVMvwBXSwqwtdu3v6++Zs/UDlLWOdZ8r9mTb362
AOXSvkITEoKQ7xmK2K2HaJLROozmvmhlatn6W6CPKAK2p9BWVzdvJTRkRcnuTRDysK9M5s3UNjd+
/xXM2yT7O3gbPCx/2N3KSedLyQi90DVpVEI4kvGFP9H1duMi9RRUsKpqcuKqC4R62ILuSFXPW1Sk
+5TGFc2BNH7ju3xG46Ya4wsi+NBps0hyFaqpg9tUyo23bTVeeg6VdAL1KNO65cJ4/UnoqX4aados
Tc+A5Oa8A2LbbTWYJkRCFyj8ob8QBWTe9VSOLGAIJgwWIyoIYPk3i6iu6hlmFbMBqm7iEbLMC1Me
shQVHXPGv5k+J1ia5jPdWDe4zemgWT7mGiJ6ZbrodrH2JujxcczoyDES93e2LzKa1oir2u5+Yj1s
gtnq2J/Mwjef9DneXoSLvXLvMvrsaslVYfUlkJYU4hfhQsJKKYG3HAKNQfZUtmbDUVsffDHHm0Jt
mhrbMcCHcYK6+amew2VjuSlu3UlHN1mvlbAwQMEEsrEhVPdGKnEczo0E8Lxb388xW99tnrIDzNFl
fiacRdxuiaSDtigkg22bn0PyUOTyfeBMPkh2QhOSvj+DOQ529fF3VuEhhIiT34EFMgJHWhQq3/Be
nyEOU1Xi25249SfUZfU+sURinxjKZTyxxxfqN4D2QWkWXoz8J4Qo0JqYF3rlFAQAVIw+5WbvoWrJ
kAHmFlU0ZErqu3iSX9QnsUYNX1LFGetw/RAnir4ty4eqNc2knNdfdKcI4DfF5V5YMqfSDmKrxJ79
BBBlIK76jFP3pNS5oQVHHhfU0nzRtdz/h040c1UacrW2w9BHPdFKkbYtMcpG4hh4EYyVO69iNNTU
21GvlCNbwvb5qnDj2DUQp/1szRXdHmXBKI7s5Qxx+QQWPrpggFBKxqD1ca3VFF0Nnz0dspNBRLuF
VmBQe0ikcu45eIW2K77pE9a6kWpGng+R+Sd9eUSW/Jof/0w9SX8wZRQPZ2EPdCAivSbzLgafSNvL
uknT4EJ547NgAIHLK2ejziZjOVWMj2MAoQSesQml61sc5BWYLYqLo/rvh0QOYfUCPhXSB856RlYo
Ogrk/UE7myd2q/R8m0TB0k/8fD8a2kK4G+Pofd6XtfD/c6fvd2v5/p8rnb8IOxZw8H5tOyZzgkIT
orUWwZOOPaBeqcOFWOTtaVcnEgzjZJSuIq1xD+Oq2njSFZZPezsWVVsXap9OnI7fczRjrlIO1CYr
uwSLqv9PNlnmCSRZGc7nH2jHgFxSgLs53EostmT3sXkbyMFp/85HPNsguyGTKA3+LAs9SPLoeJCP
1/5hp90XHEgN8q1xU37IgofgDHMVRYGw+YlUV3W1uHi9QWRqH+dtgHB0UNQdCaEIafs0YbCIeadE
yKxJEHzHueFJh6b77TLjQTnamVurQBA8RaGW8LfiexHaEALBlnCzn/cft+6MHyW+5AApTB/E4Q5K
DDBXOHyxrVK4o3b5JT/FaGUsWaPMIZNnQukgsJpqVSAyv0XwshCtJWbqLNpTZNxYXKAMFu3kYByk
8ClY1MiLTradJaM08zlP+pJce63rvgA7SncXWizaff4RDbVWntNspOtNsDs3Htnxr5hWcDwp7cUS
havYq+AtDyrCYo0+hsNVx69OE5ahSSOH8wSOosCNbUuFH1jA0Zdmro71bLdfL5XhcGg5GxlTBMsZ
cgKzbGkwtq5e8/M35tJ/s6y2Q/4jPpuHSddkmkRGJzMMUkhVENL5Ig4F3X1PPxBYxsAICjjLDxnw
2FFS0Gr62y9SJzUes3TIJo/4UFVa2vusrMvNbTIEf9BfZkTjV4vHVjMEaAYbhNIayu0aMtPiMjNj
t0b4ScBU+2NsCznWNS/eOiLqYNRMFhkYjVdFazpbFvXAXwdagdxH7XQV1TLdy4c6SOwKN961bDAH
LyC/FBD+o4Ed5l5wqBO5J1WSgfz5Rrih3v+tcpulmPLNwiTX+HHYC9deLEjRZHx6OY9Gi0LugouG
qu26tMGq0flkPlWunJ8iRlOyVROl8lx+T4I9XiOiWtX6/Jw/SajwKzxbbvjCbFzJ8FTLEvPKu+uV
GqGWLFkaw32LdDjW9hQJjHfK6/BpIN8BqFAy7mcO5jB8btYTjpNzJOsxb/M3dfdA0TgbWfdelL9o
fm8WLXA7aMN9XcKte5fk9H18uCcTGfpaO+0zJv/dmNSouiY8HVeasXGWXeyzy/cQ+8vvxqGTlrce
ZD9rOOXWfxD2wyHvcAJaVqwBQQi8GOfTrOx2uyfNDHpWecQ4stUdvuL8NewP9XzzkvpmlRdtMmrv
ntECK1X64Oxj9008hc+0pOFo1/iiE1fp11AEMHOaOoSWzGKeaihc/O0bIATsHwa6haygm10q8KSa
h4YHEjAyKNxJuKC15DprGHx33N+1lwlH/d9c8DF8NbwLKqDBpTxmHxI5YCfsfg1vLOmnww+goMAe
wgaOB1h2edsDbC4jK7kKjsHsoD+zaWGFNBYh3QJBhnWdJynTbJCgaosfg94wWsn0Jh17RAOeD6hT
QN4ykVYumgSKtyE9bjjQSDFlIxn/JDZYqlH8lgHrLJp9U960SdYcocKkkMC1UtaSX0f6IDP48+6i
RGBg9RulWAcCqJAT5+DBip/dIOPimnoc9prOMZwyqdzdYbN7P3rXVUTgu1FafvGUZ4Fe+uoU8m7y
wy6WjDXeprqXQRP5LY8N7wTUy7t7I69xOa71A2Dw2MMvITwUHL6hWs//FEZCrbhZe4DohgO6eHIb
Z13+Gb+aYLJ4djHsDJ6eFltKZlLQfB1+nfTLDgAKl4/RujV6oG+KvhHSZ0CBi03t0PFbQkUSx67p
t9VJqw4uCurRugIQs69GMH6snzTvKM804sMGIYqggDQSjE5AfVwlOuh3IXLFDWNYQA23pns5ExWj
W0HOC7R3YmtQA04/XmH3GbAe3Jw4HwVX+gxubPzpf0PR3efjtDWMzJdDamJJd0Z7kj9aPo92FuiL
N2Yd5kpoY9FigoqpFfuyKfJ4B8Hg0meVQjb/pWdORHYS4TxuasRob/QtQqEAyBMkHfXVigTK9XGI
UPljs420fdSjOZ4fWZhncCrmje4bjWExWdUbTSuu9Z+CkXTJ7aqo6XIzSJnmybr2o2cqv+SwcxI9
9/nixn+mbfHNn0ZqPOelgypfHywrppFT+hr/+/cM5JRimQXM1xKlv0ga28qds8awv3tgT09xn+AN
M45gmvKUMsGdGhl/b6g+ggv5D7eMoHLFtcjC7pYUKjVAgbcl6f4BYhLtEliKdxzuCHfGkcfFoHM5
FcoTM5XkPbDx2+IR+JxImfkJPsxXwty34zY9mzEUOJaeydTXYeF1NJvN4YbAyrQy4cV0F4ALOxGQ
GM7UmFawYtnY8XYUjTaOJA4M0XG5CBeAC3X1vhvkKOuQfi1sGuLVWsgIRyo1B+oGZXWQErNZ49OM
RmmkeG8RPzum2KM9DtFOPs+JDWXURiWM3VLZkLGnwoeyOIvqZ/DSjuJVaMyyTCwH74QOWgqp15hd
x3LFfG6yP6who3CbIPVLDTTTQhiSBd7sYZteA2ZFDaQcA+jI/ZAMlYcyx4GGiNpN9qcSp9YrNG/h
5mxrQMcZeX91B6ZXH7fxBy8nP97VTDT0K+qqacAePXD3bKWGG7p5X2zBmTY7lspI2VZ6EiShbj+y
tGo7+ur7n5zs7n0OGJm9XXdGB+3X6DLk97pRifnXrpvHdgtbkDhfy+qsJo/BpboRPMdWb/BcdQCB
BD7x9rSw+LlJ1MjfXmIfKlI+2LL/FmmPuMSYYPcu4WwOIubYqxIbQ59HphU+LbYEP2hwHFfLOoLa
34TifRGIEtWOwzOxo/5wpEuvqGl5L8hSOgu6D0xR1aQbKougHBcc6x/ACJ4qkVwKT4QSntU/s4EF
yVPlQUeSOl8V5w3bERHts6h6s89mxf2rmQTVVsjTiQXaMrrr0nr5LLL3e4p7QnchUhNhDk8sIyzM
2YUvvCKyfGXOJZbY6T7fsDslPQz3kxj7E0XmhaOSKZVXSWjzIN7L9z468Tasuboki9Z6AsOH2cT+
TXtHCkdpmMiaw4rA9ES2ecX5h90j+XJkXAff4RV1f6+oy1M/vGdTmt34wV87/JXJU79nc999FNrZ
L3WiTRJJqAqzCgDHDcWD49QxJMD+ASVkCnIRv0nDa4WNBQt9kRM415iwLBJDsDJIBCSDtcOkCOVN
lw7lScyCLgWbj2HZASQALTBUMiSICeQe5bJYCEfm4Xs4xoE2KKpTushOAPgL/9c1t/bV3ZwL2H5R
ePmObIeyP6lIbfvmoTvfOOGPSl+QESckRjB51XotfCbuF83ztmJhrDl0vPCIm7hxLZHP/tuKadDC
hD5LnFOOTrOLyVY+ImHdMYnxca4Y4QIgu38MNfXHYRZxWNxoGe39Qa1V0I/pQnxzNPUPtDf5LLXM
yHaW0b6kcqWCkz3s8pv78W8IMxlPSiZoke71h9LKqqvBoxyAbS91WZcLWHalgP4bDlyxBwD5AZVb
YUpDiehDIdNP2C3S413Ynq2C7ozGWMddMntEhYtEKgD9QSYJWkBNmqZVrTQldXYCxNVB8FhhsEsL
WpiO6bwKmc/kw0YyFdtpsfxWd/Du0G3rHM93TD0MNnERr6Ow655zMky/kzqe+UTt908168bMJWuw
Oz5X52ML5VHx4DCzxm1KFGx2WwNISRqvAXGP2n/4deV55EH18dXjkg/SB9miMTCG6KXALxbPq22g
IcwSiUPMjWlMZI7ipfWo5Voti0S3PZXDuREfFOU96xLwdW5XCEivcASUrZf/bTdKguhy1yJkMABZ
yMNOAL9g77yCCwwXV4PDxMX9xFfZR4YcUOIuQPFtZ4wKgbJPM87jbxJRRY7eAIemPfLt46KuDoz/
43XX5EW8Dek792ZEg/l6ZOYhtYv6W7TUAP3SJKJJ1mRGncZW9O7gcoiT2fvRi59oXm7mVhyQ2/HK
Nxde8GHgidVApX7JKP4iwq9EtKOCVrIHTU2//kDZkqbA/DPhlxays1CkLc34HSq79QNib4p4x90m
oYD3AkyNuaxROy5k2LdgihNpbEWuOINFGicPSN74bVSAEZdU1D+GSBWp318HHwaKZ0hgAxLiJUUw
iQFJsLveCM9LyKuhxAzJraMFBIgQJRDaQcAx1KJtv9nefFazBaP+xGzii26jM9QUrNkMyUxqc/4N
/9r/9IcvZTC8Ivc++o86v4T7oS7Lw/5gXcncLs3oZyN0uDOB8x5fxhAYz/xnqgKs0rX/EeDLNbV0
470HdtGQfiFbp+Z9lU0nKfVyX1Yd3FGA+tnFrlsxWMHTYCYg8Py3pxEWAbd923H8Navsm+siifs4
ufZiWa4H9xrWAUYMWk91aKd9z7121sHuXRlbX+FWsacmwieePkIqUj5nadZDhlIurgDXodNKtBy5
74DZG5G+VUfOvTIEzhN3SNz8MDZO7OPBH7/Aa+b5z+4aLjU8hc5Mk5JTQz3iBeLSBrr5r6rOHHMn
FMPBXyrGMG4gMbHf2TXBNhLCfUiibEdsyOdkqRZMau3BCrBK2yQ4Ph50bWuAfH3sPuJBWjo/T6CU
zV7pXyAAWZXxkC/43tBFrwOeJuncGThJwO7aKGpflRakyPwViZZB6gitwie5OwVMdphtwun0WgIa
vJunrgQfvNzi+0X5e14FyYPWi0yekkB80fIeBxU8lyFnqCOvVSHUMqsKLK1SwFtwwb8lykQCnGJz
p8+ev8x/8wI45hmnsBlalM9ez+3YykxEIEPoQzm/xWh97DZa6j+tZY+TnuBjQAK8XBhE7+p8UvCd
ENUkfaVqSqVJnV79n9BTD9NdPom4nH2n3/hx4HGU6vxhuleRv2E1TYm6d7h6mCJtn44jy9/8epq5
+J/yieDU8IELTTBk+XzE32rqAEe3yAZoQ38AsGS0vfX8qf8R8dTQ2mAa6MTwtxLKumy3QBh/vozT
vB2C8PV3/U36mRop4WuWYca+hVT/81UlYc1VFYtWjU6023H2ubSVJX3MGICHAhqYBcIAKiTCl79M
wyL32zRV8tS3ThV4mtKwUreBHtoSJwKfRs4f78oIaIXAmjSbrRTuzEiJchEFDX0ZL67p8aXTP17m
LJFCdasdfQ/6SgPTHDiewBSWk48cjtfnIVCeAZGQC5NmxgJgmayfFTAmWWWmBBK9R2IxvjeMF2H7
wqrP+JqF3cqPJBZzG99jfmFskOiOU3Cbn0kFJbhfgqv1VCHuG/WcdqKl0tW9YhEG24VTi23Kdw7i
tGsVkoMW5nRGMd3hM/cUhq1DjicOH3EBMJuz8Q0HgBh2EXaqWmO62ysAtjR5OgwLRz/zzVY6TDgI
J6CuoB3D2IE3J6r4ssBNyIbYb7e04nwJiKO2wmBiJqH3ZbfTZSxNTd8m5ihoy1ChbaOJWBpSwIfC
MgaRC6pWQAFwIdPzBejO2BeDls/jpoCI85Yfc4WlU/hc+KDJ7DM616sWNR1Wy/H4TE4de/o4R/gu
Y3UASTLIu/alR30ijhyO4oazFZRllIXYYAIZvrCN06plc9VDpRb8Nj5kQrmrd0nozP6fzS5tr9Xe
XQ5dEiLZHC22GWIep3L6Cq1RbBX0by9VADxk/lgPYNAmWR1Kr49a/Q/RlLVeLvXRTWSXLpWJMUxP
FhbggfX84ocdVYOQRprwaSjOhKi1UFv+i9zJfSqZSeK7z0MARg5u0iHFlaMKiiMcCkuug41oYDG5
sXLoimlcfeVx6+iMhpL6b8PZeznBsKUTynQhsRYiSNWFpW8o0n33Teia5CtXoC5PXldRfjOqa+VF
L+vQbn4y2ZUhYpIeZ3i2ElQ3cHMkHpMMmdURImyt282x/odOFW+50uJZeuWE+2T8fuH/+aD2TCH6
uUZX5Sv/JRlC8j7+MJFaSvRiss/T+BBdV1uU4La2un5l+0YXsVobuMYMTAHsHj08RBc6sRniwc1g
EfPqNCYGtWTeHnC+XhmaJ/Rw8LmumYIXl+sIy+I6QHuh9eapjVvtNP9DeJm/eMOSY8MdT8uPIxYI
G3+l3vNYslM1+lOKBztq8dePjfdyvOKWjlguak2amC/O93Wl0uu/Y6tTQ9HsMvN0Yb160hsO6Xke
5z0lQGs3pIK3TqGePlRwBiXbW04Miy0xOCjb773++S7MAu5fntNobLWhhF/tMTXGDZuRgRRiCqk/
wTIA9EO/lyntF97NNzfPeAJjGB/WxFO/yabuWgZSsrOYQZo3x/EG/JNM4c8c++2TVtjiSKiLuZuo
Vy/x0OJHolPHQ98MSpq+joHID5MTcmG6UkPXJ9/vhRly3kbrJmTtdk6rr/z/2SEEHb64QwYPtT0O
tUWPu7JIjtN6FuiAk6jxfqESApc0LC4cR/NbGF5BwS75x5tvKkaBlZ6oR7qfI91Ku8Y4lQb3IiH8
jIEHsnbWDEO36aM3dqpF0AYvzSWViltOsHuIuvJkeiX5P4Dn0N33KbQsaOAfiDtUkCzGBDOlQauL
BwgWo2A7kkeUr7REbU3z99gGbw2J+ISHjaK3INi7Z+q2aEVowJlkwV2ImuHdoi4QiIqKZNEuiSZB
b8doegwlggPUKdSeIE9GSsHjn6n64iJR5Ied/Br6V5f/vta2A5K4PPRjP7j1v/+tpzj6WZc67Owa
lakseltd+b2qsnLsxup/6XeWUZMMAHPT1LSprysCxN3P5ErxIgkYGM6pQDEMiM7zchHEPbRDOeON
q43wPccWOZgFdUupQdsbeT9zXC1GG2+8U1wtycB52MaWD9UBzJ2m/XZRMprSij0XbiXl3NyeLYHi
S3uQiM5JMULvvYdVcr3Gor12UPNUlaWnOLWrLGlaRSqiBKCOlbN5OG3OizmfWXnyWI04K/QXHo+L
HNr4RubsVkvtbOf73iN38SjCAsAfXk4F/5YUMe8et2q7YHgE49b9jZ8jkPQU1CxD0koYWuNBPHgq
omfMtoUav2pqPwbbd+fBQlDO2sXeK7Iv6apBkoX+GX4KB44p8DqAVgHg+s6oMY/sX7Sp05CcnC2R
aCIY0TY1OdIU3V+b+gLYNG9D0B8ALCuKKDQ63pamwwfi56gO6NauQbO9mYdm7mr5SKwXo3/dpHgp
UHQKWxSEARPwG674vBz2Z48ZG/Ojj5+zvd6GLXQLzcX/lSgqUVIi8qA9cOtBwsLgFTTx5irxsWae
oq4ZTN+ZkMw0HHHm65msLDj0ZjIgHv08GukeDK3Pp52zzrP3q7GUMsWcfOTfkTHUwmIiGxnDPx8I
rST7AUqWuOVsxq11u9my8QSW5zn+aM271aLmymgAzqx2BO+LAFIEDH0KEEqMK8+H/WiDllVGtups
qD075j7AHobykA9+3fnK210rqk+wEeUOa7DpZi+qP+Phsj+2haONs5P6spBn1PyP5/0dAw61ASt6
uvAy6/1rUE4q1rqDgH7BFkDMYdc9Q3qXc2cCVmQZESJWj7Ak3J8R8bbuh4VoyjNL0TdeC2a4VEzX
F9QjlH0eRoTHUEH0GmCxRH/7pp78EcNaGiEvefTbZ9Pdl7DlF6+iDlDSdIxLd64qINebixA7ybq3
HlvZmLPyTlMpTee5I+ZNbjnrz9Sduxp/g1mz7Rom1VTQ/KJCGy9qNQYIG2vlPC+JdQ7n0DyrpuKD
5zuK1xPz8W4OBg9unaVwBTusHMy/8PXXUfRIYOBmt+H2RuiMXFVUQzyavIXTAXuIRkXv1hqPvrz7
N/kYKoEsZf+x/znccFGgQC/4c1bAkpwlmxhTJRtJNkvosewNCO8lhoT0AuRFpxPKFO0+5hB8HUSx
E1IPWbpp6Wqc9EOOcCtArVKVWJ+cD7Tiiogumdrax9ZMRXv3ptxFFJmzChEzuFzy3gUuA1En7+6t
5xND7IHhhFwgWnS0XvQk/ZR7UpM2aV3VK+NuiiKVRKi0Bg3sbsBBhDLglGtQdmPvQjfPhaLWznCZ
Rjlmm0Q2xMaUtBkZ0TpZzfuZSKL/q/OLWeRucRuLpDdIqljESPts6i+GqY3RqioX8Ukc3o48IyPh
70Wcg0WFRmKZOpyGrM43tM0Q7VRYR1cGmJoOyAxuuLCAKZ6IIETjD9e+w8Wnfige6fhBmNh1iwwf
kQQ+IEM3vRcRuY6nM3YAtZlpu0oUMshOHWBDSJboc4MFmSpN1W3ZNQkuAtdTpUjkHKgzhARDTg6m
Gve2PvRcFTSAotlTSmSrjvmbM6zKQtciSO11wan3ap0KqbO/Tyd7WlgMwOjfMFN/BNykMu9uAtK0
mmMeiTPFmyFRFfOac4YjXLOgzeyVm2XUwSHPl0Kf7bprbvArxiX6SjmmeP6NOUC3g1lpJdeFtwdR
HbANBC3C0DVFMZ5eyYGofU3lcQS9DmX12zshKz9h+w3NKQxDlDoiBNWNF2ekqibXhFuNSIhbBvVb
UxbmQNRqIA40yHn7sqvwlJjbNdDYVhjtNazwIZUGjXVqcljNpIde5y5HCg9+ZfkC8x16tQOYz0hX
LVi1YNJ++mhk1IJmCGvuXy6wSL37FENdhFyTzUq1Ki8wiDPwfgeVg/qOkpesFDiCbvGrWcsi+djH
SFyRPTfQBz5izkuPtPAxxoWu+DOkNvoFBzD+wmKdvELBD8sTjriumNj/RGTJtTiaKpwyPBWlsX23
VUIJVAWMVj0uwgyjw7MUSLcvQQtfOo0Qn+/N+HLGp1UnGB+Ajql4/fUamQ/D74TYrmHyncvG7cFh
3owLhCB+zkhus2OcImOScxuwhf9hpDyq3cmh0QO4Uo9ONGGX6AVPVK+si1UVuW7qMCvZh1Kl8ROx
tUKx6w9oFTsRzzsloUNteGM5sd7dXMV8Tkxt2ZuHmp2m3mhpx7SDEVcXmNIGMYRbkH2+xrmd/RYG
FUw5HYAxZRYo2Ye7i3nrdYyw8zKkYkrtw99MRith8MndXwp+6Mn+oubYp6CKY1BFwyEQmwi+fg8E
+5AsPbYaWYc7X8gRJSy1jbx+5ni9ASrgrCO4c9+Rib2LkFTPm9Euw+VY912NMKL/rC6qO6xLhyMm
ijvnk7RCINVxOUjLXJMpbY3ybLz3o2pEjJuD1RKmxBwV8SafQ/7immumalnPoplVy8EdNCRbAtU4
Trb7nDyMf7O/oSWbFvtszGZF959fG2QHL8oQjkTkrHhGrP7GftTyVGVdVB/XjR5xugjKnc+NIyuF
ypJmVJbVU4m6tucERR7kgA4qvtg42OJvN8pPvogqsNN0KTY/C6bXfJmpNRi+Mq336wUEz6OK1eLW
mnGz9wiOBC6eD2fFnlh2XuqDE4CMexd+dtc10OuHEyHslvvVoiI8s0/XxXDRy8zJ9rzL3Scv+jeL
c75vmRN2hC6P4RYcNi7kZ3OD/Sf98lcQGEiOuAs5AQEZ/FsWpyBoXTBbbatkAAQ5CI6vqQ5QaYL0
vX60tN37CaFvVd4rQ0HUY5IBH4RL4Nh4VauI1VlhQoP3dTDScfsgofM2C3Bdt0NDvdUA0NSKveTY
Vl97OK9zeRi6JRE64T+gtek9LsR9YP2dy2WUZH3k8BnQhdBOJHwMyyftWd0xj2QkXh4J+oiblDqS
nVhDxf8NHzPtMphGVltKa8A4Hn3Qa2v30sV3kUaUZ6s3zeAIeWZtFTQdZc48O0oab1R3ZLAhu3TD
EPQEypdD2YJLJEwTxARxalJhUr8FzNvqYocrf85Gsvx5CihnW4rHiboEOg1h70Qlc52GOn3ZrMFe
1T5WovtGECe5kZIoGUFx0KIBnEUV4y0D4QeXnm0S+kUHGMddHcC/EZ0aC5OjLIlJQcbyLMKVU6Fg
oz4b8MQ7IheFyxVEBHs9z1P1nyKN+ggSt73GS9OwtTGTsqQ10R/PCtmaZf28Y1nuGtJwH9pAyhx9
Hm54zVWXKhbmMIbq8iy9XAhzR7lwKxo8iF7dHR0HnqCg2uxv04JgbNpjdtN3DLn6hHhS/K+kd4H8
T7ZpJxB+m+fcCovhZq8WV5KTuXy/I2szEe7x0RXLTVEncpSRHXRvHr67kg6UmEoghV5setUHpQl7
KJJ4ose6rdtVZ7vMUX+xNGK20CCJriSRI+Zd6iNoAUNZcPeY/kgE4yZ1Hng2zuZZNpGj+xoiCvYh
Pihkktl0t76UuBX8vTzAryKoMXQErkhOL7W1zs95hAWuo4O55LWlxfLf+XOFwg9u+MNfe1qb/QNE
dkcrAxILeK5IY2mFtZ+6sas3iPgHtmRw+ddgSccDQcza+2XoPLN+v8DRicb5hOX3tUUTzcgZpGdj
uZeYruuYzNCNUWGYMP0wKrvJrQ7hOwKqUzZEuyh1EAumQY0Zmu8KHZvXZAtse9TxHXnLxp/peFa8
Kp7X3DmHw8Zkw3DiTislCo0PaGeaMxMTTINb5dtlOo45z7b9jLMtooCuThfddtsP3IUNmAbkOthT
G64k9WHMC7MIlmgw9orwUw3ajwOcNeA2suK/yXwCHnGa/9RqR5GmZAltt+585Oe26Xq6Iy1RneY0
PhNKwNJBufJbT7Bl700JnFohQxkUWzop5Ulkr4kGKUnOvIVsi9Mem5cOkVQf/BMo1qGnEuLx7OBe
THbdTt0BsdNmBm+QZon6MrXpc5wokLRGcFoK9dBid/Y0c021TlHyvgDetGw/QnNV1in6uZIb7i03
xSLu1x3/UF8tVLsEam5p4Mp6XOl17IdPMf4p61rlF31Xg6qtDfS9K9c3UGMJAs6JjNsnGY6ggavC
eJud20dTZ9s3MN9sJMnQC9+cVjFbQEl8ZYqz7UuY0LbuD7ioB85V2FDq3DPdvqR8/Io31BHrw+p1
id0wORhyzM9biHcRGTtjt9UJUla+2iiNqWz5QdgUPxZbPyouqeuAX2VOKfwRtGb4HAHxgFo3z0Zy
Ad1VEBqBOJmg6QRlrPg7Vk3Ra1KBSgZZUwQ3Rw5JVMtoqcgnQecbP/IkqdIZWwI9XPLIxXkHfies
i/ZhPqGRTCVb8pY6JOfTiBzz6+XOgFdpe4p62ECsPXu/yeHB1Sup5FJOx4kFC4kuFNECAjkwUSOv
e0i4GTc4BUoFtVVTclFSZD0/SUBmCZmbjHz1cYAqerAkPg4+83Xc1yPC0qMD/8Kyue9LfNWc78UH
O/y8HMsNRY+AOSYuHgoP4QLUCEeGXV2ckTg6MeJHvsCV4SmsT6eWNp1W2gvzkySi7JkCZNqDyh08
DjXR0Ms0K48ccPtlrkfVdI/QUQiZRxINox715fGx2RDo6Vk2XsVbomPjYXkeb2MssuwHBsjPguGy
RCCQb7mAf8OXr4tdBog7RaYaEC+GW+aQhTrXJAkhm8krf1ME3giPDGKs4rvSJb/3C3076inZgVi5
fP77bAAGm/WZFrC2afYan7i/wnD4kru5ioa6rM0y7bMYmJjgd9T/h0UkTS7yLDbIl/UvCrKRIMV9
t9cHoS725NhGG0TdmTP6a+lHPQK5hSBUwThMy5lY3vc3oCN6tCdGDG8GWDUsG15kuZq0xLnHJjdJ
2HN+n6KWiIpVbTIEXgG8+Qot/41wlEwTggMHdOg/TjYBPd0XNsUGfn0D/JXSXJHtZCIEjrGhIo1t
zkvEwZKUrY8CdKbf2G6k8kiIM9Q7mM2rAE3pvU8GXVWyf4INHOhy6L7u0K8qEqKaZQrmKi6d/L28
iG+z9mR5IZutTuuJBFHh2AeB1fFa4yHXyuoe1CW+QYmygDsRsNTz06TRJ3PNPpmibkKEJZw8+04i
UBQofInF8YW4oCit0riErmHGuQUUg4OOGcyZCuOWcMIw7V4puvz5rOnUKit/OXy2Egyh68B3dbEJ
e26JKmsgP0ymX06m9O3PgJdtJPJSvAckmVrJNekkwJzxAiujHw5SDsCXXK0P0AeTibd/8U5DKlcA
yCmKni3+LBSsxzsVYSrqfP0KVZTtPiyG6QS+QomSkoUNa/xG1wzUOnPQGkSpp6ywkS45qpggifQb
FY26lwC9gAmW0VnFIH74bTjRKt0mdSvGhbEzJwpbNkzyDw2ZR/sIVjyrDmmjGVPGGaX2C16b+7Pi
qmg+albLIuSJJEdTX3beLBcY/33l5rQqu+FZ+NNqdBbND6FkL2ajIeQBhb+DWNWdhWHAdG71Af2O
FJO4tRbryI6lhV3AXrd90obugGQGqc8c6Pg+Am3KY5F9PQMnSJrNRiwhwM/qARhHAP6FLMDbvbz2
1F0DbL03AR2bMa8k94vfofDoMg54lwGNbrDDOROkXk4A9oQ/5H8OXiS9AWwpsmsRCDWdCH3Ph7Xc
Vb+A7qdHJx61uxk5Fn4D/mahK1UQ01K6FT1MwBi/PM7HfaYWeBaDR8/39u//N+t1XWT27cNH+3II
AuFniL7Bsmkh82kfKBQjIfS8Ap5fd0GB5SbVBgle8+sirYPqk9Pp+qK9sPRXeu24oPZiFu/JV8XK
1ZmxJ8E0k3d20S7qhyl8DIUvtBiooBusOHzcVH6SxDRbl+SaBFrFStVw+SH+CPBJKRio2z4MwzLZ
Y11ahiXkXUwKq+9XXt/J0CQOjiribuBwGu/0cUM7C0WRodzYOp14acI7Bc5NClBNYyUAORL40WiE
froUWh4F4sGs4xAGKlzEezyRr7euuAyV7Gp2hrSLi2MJMWvvDR5AwUDxQVACn5ghe5odONqmu7fF
jBELM+8tayzhiCbcdYHIld6FMW/BiQ2hzf3R7Ui7YkaOWZB5/6e21Gcoq03cfSK9H1YVBNonaw3P
cK0JI5zY7RmACWygm7GK40Xk90A3Hk3nmfZYXykTWqeK2eHn8j9z7De9DBqhZXghGu65Lsmfqf99
ZybnjL5+yNs7oCpWB8CPLsRReCj8OnqjpI9q8Nw/+HlFbmnxJydttyGOZ4u9mMFmwFO3NRZ9BkRi
U9ddYCicqDtgFWeuA4qBlRuptD94JvXC1L/9kq7AQm6gzm8L7nFq0hHyuHp2oWVxCVagpvFex1N/
MHz4FUx2e3IU7EuUe7lIVc+8zKomKzacee8Ify6KinVWEUptqmCayuUqwwhucgq172Q9fm99fNty
DCg98wzcFQHUkmk2hGT+EQGJmplDe9M73LltRdtokrDKkikP7NHIl1sTlxsiKfoBhAWDPNhK1pux
35L6vqs6OXqR90R54n6uYeCeoUsuQkm1Vwd8d+sIKKMEiYl8aR3IoH8FiutUr9SjlFiEZX1eCcqn
f+tgYb+tkstUwUaRdknn9y6XR/Wlh7Nbwf+oz4zFPPateXkEPCj9F96IxG5gVAf34ytCZVU0zDJ2
gPN/3Jtn0PBM3vZDGvbbpyAnbv8woDVRyj2h/kLGn4cmu6c8YkA9et1bDcxcWoHGxJW27TK4Ocsl
rZmHSszBgTb4t3gxzBlvT0geU12TlmnyqZ0OpcEyz/GFnbZW6SUzGYcly+ilhNMEY7cFMA9+BJud
uFMHye4szIYbSQdAG4NmHJDHhPAfL0/k2QyhwZ1OKROrUK5K27fjl6aXil3KPIkPai4cXwkPMLdI
zxOAbQ5ePiS0tzEKLzinF5Q9M8SJbY/SKXotxi3eTM/To1qzaYPsneWAhrVa3/3nKyhrpp6RNXjc
NN2Ybt48nCoh3IGSBNohIc3t/gGCMbYZSizIN/6nUd4PI7BhS4/j2xYX91We31etnr/UWjYKwgAq
65475jBFzu3spLYOJycQWxI6+jsTUgSRfC3Dy0j0acGWYHZlxLFxn5jCZTr5asGYYkHFrmEKUfdL
TYBUGUAc8tHAvyinl2Nile5YprSONg6ume4nLqwKKrz6c9GEPfuIBgJJnmZZS7/Paw4cKzOd8aPU
Tm+n1eKDwB6aJCT21Z7oRSer58jbOMb5QMLPzX1UENM9WpuSLwSoJAZ0B7oD3jokvB/lwcHiaokR
3+SFvA6LWtTtHRLYqJC8FCHC8DEn4euMJRMvkOX1Ug99vYnodWio6WGgFfGr4tGCzcqzVAiWSTT9
1zX1G5hRGmLPzl4EgPeio0pG/gUQ6ZfjBuGxXJixo1g7jA6dRgOvhRCm694MkotICT5XCE/FWWxe
rEcs9ojndAMi171gU1dO8TcX4kFLlti7mquz4UY6+8R2p/OH8t3GFw+ETDWTY9N4g+LQI4JrRjXN
QlfYgtzmyZxVWawdCT/CydigwcMuP1nUjtfCjBCniX9IyRNksYh1j8FHnFIn9tfIT/yGmEKb1w1i
khJKdYDfKJvlJwIYG9q1K6rz5Dhg4SHbzTEkSW9kK5khZkkcpjXgAhizZKWnEEhRzKYlzJArWb0a
tzMtAkjYG7GNSTrdp5xQIiFYy2qz7z6Orh3Sxu35jwg7K7cdvieppVWlSvhlMQcAs5UPje4P09ol
FdXWPgqCNARMoImQL/z2kX1U42U932AiNUO2NS1rmyUnA9iQHLAnNEhaFTB148zBtoP6DqZQsv2z
UEvnOPeOhp7zUM1c4iCeH5zLBYVOSydtq32RU0TzOhXfAA1gjccupGPjwxsoOt7eiLYXheW1TO7X
YiOeTx7m3505lMSvETB0Q0oYSq2pYHsGRq7LJbGxBDSxUP+yypOwKvJSim4DNdNGRsaJ9cP4qbg/
X2eKB/VDHpaVP8Zq7UlBVwQBbN73Dg+Q2gbX3kQvvv01p+FFWRibrcslXvyww7UxUPD8+ZAHQUh3
j26B0vvR0j0cmegLEyKsnfOLU0IXWry+gEqabq1ApbfXylhaXjNRI045k2Rlndw/vLMo2Il5YQwX
ix4CoSZ7xnWgg9b8XYXwOJkuuhZdvQwl99TUxwpOY/LFZoIAhvsEUrIpmmKIXzwbspV9KD7Oz60n
Sd/drmDkpSVmJ6o7g5rV84PZmWp/CznyV9Rzbitqc1itSuqNqAu7JPCi9VvU5rOtjfXbfg5ukt6s
C6KLK+eg3t4RTZzK9wdjOrkNRQ51H7sYI2T6W6GELYFHtGYDyOTveXnH9EW2JKfyVWiHQn7JFOfV
wPQdgAIpH4FIPz//1upuJpLlZ7/6m+lodnj8LZjpATv6FJxbnmelG6rj/stryTTVE89rxR1rdiKB
j4fBl0OmLTuhugw6g0WiVvo9FiC2XmVYHZTB0RvEgwEH4Usw/7698I2Z4ugzli0MrFx5qu8VAMkn
WlUMBwW0QmrXgQhbyr6ZoWMc1ir5c9UlTmbp4FNFzI53fZTn9rcv0kFBtkTxiZvypk28/yTyz2jW
5zwzg6TLEYKQcBwQ++df8yz5hokMcZMe5BclbTEZxAXLPathPSTKgIo0PsSfnssHu+7KTeizhHb4
SOUtty9Hg6z8e/AC/MqUS1jx3qJ0sd7HYcrHafdNv42HAGBlo8p0KnxVajiF3hhW8jpIxW7yZWGf
2bOO/y+z7chxUfSF3NOnWhdcwYkoggl1iCq/UjzQr9Qz2vwzkbDBhfYivOxrdtIBymKcCxLWhxxm
QaCZzXcJT08vPR88sJaw4XkiHZTbMNUFE1T+drja/nF7xtrV+WlrpaKwaWi9ogataJmIHez0bJbq
cxvFjinG2YP23Jc7hnikx9MjpOyblrPEP5o7AcAeIiKo/2wXnfIeGKDwK2fAhqTSDECp1iRLz+Pz
lYwPexwPrrAVj8VNKNOFDfqSQSvR23wRiSHgR2zdaKbchXOxrwAb0PMtpN4T8BMzxXYjwIlh4mA+
vsPDNIrMSLdi0RHH4oweN+V65vAG7U3cDLibs+Ll3hwRT181W3JN2US8duwMLglTLr1lMArqDwoF
z9GbSeogOWbVg32AjSB50+aoXbS7IFXQLHVN061jBK3dqbBRM9lv9VmhUSKkbSfhas1UmYj2AIp9
Mdvd5M98zoDIbmlNRGfnIPXSuxXNTkk7LSGR1yn/JRDkz+2sKCyl5Nx+sIkxnVrgcS+hhKupHH65
y/VZNQv1psk1pgvgRXYndJMc7biho7ipyAl+ZKcmxkhSmcEE47S96H4SUYV+SA/xE/bScvHLAgRv
n2R6YozPsRkfu17K0L3atid3D+PhWVMXRN6Ild/OPuTIAYPrLOCCKY6jEuRUiuVVlQ2rfDynq4BI
ItTIaPGPzdJX2OpZaYMsvpe92AoHcnYDljf05szH4PasebOKQ/h2QDVebeaMYYzx1/0HyJENPzJo
wlWMGDsfN6rHrlYq2MUFvvj4fCO7YIxCX6TZbrbpHEzov45ny+1t4bm3I4ICbevc8FLBjdtMzJDa
ZmfVS2PPemNrSi+kC8f/WxoM4bNFX5BaIMLlCNSePwV/+WfBa5746x9Yc3iZzkmhvzhk3ICV3/Lx
IPe+LA6CaJdJLhEhr074MpcThQnQokyCYGDJmqUuFGWkFQ80UNsi8ms70yRnnWCqrpqIGFHn1X3K
GAJw/6REdWoRfGDL2xKqXsNqtpaX8agefuO11Hxj0JWJ/9pKB+XunoeAxHqhVSXVo9u45b36JOBP
bAKKe5RY8wzkE/0pLQaxQ9seXjmUH+LlCJSpqHuSHW9l05y95MES+DDvdP8CFnuj/BRuF8jPof9Z
WwDLSQwMeaQFiJYgms7/oTjRm5nPsS7ZYhjBkm6bxg+pzE635LOnIz6kZAIYv26VK2AF+eixfgGM
paGR2fFESg0es6s9Ufm9muFoCPITC8lop6vugN57v5XW1oVwtkq/0ckrd5OOxb35jx46Z7pj1ZCm
5UErVI4tnFJr3Opndyb8i1BTwUKrVe4CbVU/dE9iQVd/kwS1TUSXWDo2mWhvc7ZQ+kJUHUTyVUwn
+kaoXp1B0M3b/uPaOlKCcljVXEFB+qwld4QyhXuoOS5JnTs7JqMR3tOebjrcRMEhxCIVoKXvCKC3
hwP5UQYgCE/orm2195ok28LJDCGNW4pIFtSlScnlkIwG0FoeqJyzHsXA7hpwm16pA8VAskrTIb8X
oPiTLJ+VES018fkhFYf2MRqYZVeEVcuCs4lhsef5OeWxuWC3foKi30cFYoMMiC+3gbzmE2KOfr/B
K7QQk7Ufk48Ta8EnVLoCV+aN+mY2gU5uD6PuecR98AddoCyBJ+Z8n79dvHDLsGNJbkAURX9D6ebY
kAc6ww9+qGVTH5W2a38FD7K825DKZc+v98ofPYYcpgp5arf4lE1AXTRbYp4NwkaZR0tbbYx4uPH7
BY89/0urf0Xd38o673zotufou6OHZxW0AUBbAIrIO0Lbz04DFNyo+puAmALv/0eUeqIh40fSsIe0
xQVB7KSlC0ZcmKY1JyWNSAJwj2sukDqD0wAAqguVywlvIshlaiJ5DH5HmRXEiXhVTwcyMxWp7W4n
lxwzHJZ7UP5BXygMsuzXcO7b75WmZefKvafj0joyrLBUg0EWSWUKw3B08AJpFIxM1XAKCPjUPJ0U
rwL2zEjHyujrVBWuCie2ENQyY9i+a1e7Yx9rEXfhc0jlhUKD9O+AkxHlCg2Bxip5CpZDToTmzCGu
tqbVYcVwqAzQdbwQ9jb0q4NEF6eVQSkxdwxTFz+b3Fkuwtbh36gOILOCiRJUJxF4xULDyV15Bu0y
r4odCMJhRUdsv+x0WXu7EEa4UdhQtYHo7aEPkc6A6/dGUrt63A4lSp5qJMsowLPo+YesrPhZ2/hU
TNHPV6GMDrPjVKoC5V39qUl1XZBADRyUIdikbWkuSOShqWUvY62j6Tnqpbp9gq+GzN+JcBRlRgjc
ztHTs9G2LHedaCl+UaJKXj7EErql27AgaQ1wASDQ6XJ5mC0nBEAQhWA3g6RHoBQvbbjCiGw5oFYJ
Bg+ClnoV56GGdViyJz96c2yNjpZTkfN75x7wmICG1EXOZe/u83KBTol3wNxH2DX/69wlUineK4D/
Vx61KXPN8LkaPRBIKJxcyJNYYDb4mA89gx+yHrnle98fOYRQ5UXatoZncJrZlHPENs/8Isikl+4V
H/jcTMzKgjC3mgBfa6p35zTrf0Y05243kZIlE089lMybuuSWsv7xr1kBpUKnmLkLUDKKjMYWgrpY
J8baHMv9U1Iai1foY9vKItr8r8XlZeKxOx5BSRGTg+YMVM15WKHA67HWtV1jlsHY1dyNmotmiwnC
z9AMOvPJrK1dbp6dG9RAIv+2G05Ygd3idwPo6OO5g56/+AEWSLVCznLD5RmNBRa6SRgB7/5M9W0S
0u0GEV5Br+QN8+GQno8cnrDmamPEKUFI+0JiFaBpDTgToC+FCVXC28tO0jVxU8JS8kQpWHSbM+88
v2l45uP8m6FaWSrLqpTV5Me29yqPVJ/+RZ9GS8sFzDLBIpdMjiWxDGrquYutoy6PeyguEfAa3m4c
6eVnqXUrjWKNKBt4eo5wnK0mJdJM3wku4JmtY5hs1iRxKnvbR8BiQ7nVKFlZo3OU3Q+QhYS0/ZNx
G9w9TRZTabXrTh6rQhxM87A5cbOPa5Gvo6s+8CkeFOcE/8VnLsBm0QM+ZifExaZ0jWnqCHAj9dDx
PdUo5IyCWH3NlujihOdFaPeap5Mg9r2oTIYHi0guMnSbWl4n3Tmi7hiCV7wn9o443ripDOP+X5gd
GcmAb0kAXeUFCYmMZlMb9VJxxANwQz+O5MTCsdOuWuvHH0JJ/bePJbjri3sMQ5lstykekKewE+sT
LeJ0ONiJrODsojMJi61U1hr7nBY+DlnsEjguxj3/11ezkhMUv9X8dUBVuhD4ZrStyLaT/YShe8ub
8zGSRPFbLEwywcPIbZdpOB3cUVlmy+IhvNse7fjpMLX8Z+6WYDnC/XR45+mJBI7b6wvlNCen1Xmx
EGa/RohMTkzXSC2n4RkWACCNMy80HA+ukbfB9IGxyq937rKnY+T7nc/Cl1x5a8Lv3l5GxSVJTwzS
YXlvTGAkZazdspaR20OnT3PnVUbzfD4MRyJ04m41QfWl25Rh5/jHIT8klmpHJUWH6EArBvA3VbyW
Cu4QFnU5/7QeeNjMhCjpmOH7gvZ4kzgd+F8Z/0hX31VnYhpvkPkFFJ6fGggeMP3KXwqQ1N9l/vK3
RAWAeUPnyxuHWSqqpCBkMsDbxoVCNa7yJTHv/i9thUYgWCEvkYErfFYdlqXX15nvJuo+uVK4bTqJ
sgyprkZs3RW2XpSjouHa2QmA+qftJur6LOXMR63aSxHP1z319b6NZGcVfGAQ26NsmIDYH5OQOM2f
WtX8FfuJmYLETAEC/ZOeazYQyXGLwCZZbovsZZ5uyzcFo0I0e0EqlR0fSpX+1NLHU0dr8OboNxJd
UsP6vtyOiOKA4IsibkfAFGc3YXnbASHw0OyWWlkdQBH5VuyztVI2mlSJYxbeBDDFgdd6wW134oVv
hTlfzQLYSJpV0+7nA689M6jDeEmQqZgG5QTmNnU/RTOkZFjw9/1XiCJ72OFrJ+4aXg8I75ipbdyX
6wgt6dplQID9mVln+Q1MRtWwmThcJpAWs8kBcTR7QZyYptGWm0eXAszM3xc62YMzholfv9FLBHCn
DHqkJAydMjWg5BnVzaoSbABi8sglKOV/JZj4BADAxnv5o4sFFG6mi1s8yKauOyIYD578NNjMnVW2
JcXNxYhXVSyaDhnU6K95huinoT6/ogu3DMCyjLmdRQzIwzJBX3FVTvkWfW15mE4G7IMoauT6jzpK
hmqmJ/F9xC0tbkKRspi0cG3XL6oXT77wMxsCuG74TXaExIYyyCyHGla5U+szdj04VMGW0oWBWWxi
rQlHRKJiNvji+LZlCbdZC5kTspSsvuaoZqBOwqrXQNxUbaZFQ7fjzUw/pAg82W0Lt8i52QU94vCY
9cCGhSx3o8ImPeFSF0of9zag+0vjf6SR1/0I0P0hsq0plHq3L18L7OE5PeDsjzx0prIbRkNQl1tn
OejZF3GOS1SYubOnnJjXStUfrQz5+Y569USgA1d+bOEkvLsDXg5X9EkqZmznXFDy20J0UtN9nebS
lXfyRl94L34CnYgK6s/Hm4HAVtPikmhq8+8je5kbFEJLEotShursSEbv7Z6GGMeskRuR0j5tkEac
d1cPB9vR6WV9dtYWVNAw7/crsoU9kaByVr3hu7dMLynfUBSeskhNxyoIpsW7pCEPlP9a4lEJaY2n
pRmyAS8f9pCqdt2Y3kBYwtdJAlZ9n2OAdLKEVUn2TVj8gwwxuGHCfySI2OgB0p+he0WvC9AGykR8
X7nb7ZiP0B2aW0EjAgLWJeazmjuUAyICsLoI3e536OYmMeOKW/3+ySfULqAQeCkct0oDY5xkxllo
vqIz9eKLPnOfkDWSDfa+Y1nYpSDKf+8tAEFq6ab8ja1wmj9dd4wXCHppzfO2xT0aRJ038RgRJYeo
o9WgeRk4UmcB8pn9jG86fQ/SgOWqRm/3B5Mg1Kz4MRhAvYMPqzESy9BMmbJcyzBNLwTU2PQeRMij
2cWtOTxAQNX0RGHic8YuqH6jzc6f+tvHjvwiMBterYI1n4uDyhQXNhmanFUM0C52fJ6yiu5mL59O
O9zMiMTiQaPmzrSFf5QdlDEuzkSCfoCG+U8rVTzFxnZPTzV4pQEoo5OFV9b9SDiLb0G4Vns9BLxY
qvFR2J4VJFOZKiowkQauZ74Z+4U3FBSUhdau4clt7T/LchOwEH2UsQounLYGjyRRfSRMSfiGEXrn
yDNzqTy6vECGGsinTnGqWjQ2idWKauoC6WyVT4QAt36ZaCZmXXkqKq2UGQtC2nrH4PzFbXiT9xe4
dXZTVjkypPVYARzXjiFNJ7o8t0oZS9YWPezevbZChrMq11eVqJZ8/n8ufQIoHGzlDFOfLYeGZp5I
EqHToW928rtirc9L+qWxniUjkxVdqxlqONU9BkeOgKoQ/oWC6dORrtcATjNQC6HRDSP0MaLHF40H
CDDvnBlgqS/wQ1tdQHQndnXPm7NrldGx1IKHGxCNaTLafS9AuYM/6Vo2nDPIzZNtPQ6tzD60AiaU
52tyXJ50JDNbGBdDE7s/QPmoxMSub1lkKkrTuM+Ygr6Ml9L6ZI+Zan3a1v422CflXYiNhnAUWt7A
6HCTtDNXgQBGCfypUrNedYYAe/8h6b1Xgr5fyBbxc1IwmdcQ11rYipgyysVrg790TXn/YgqcTWHg
slHmPep6Uo9gjhVYnAQ4X62UKhe9Ov/vdpbmRCY8fSM6JB2ZsU3zcPF3gTAw1oif2yC5GQDLYTBG
V75hv592PkDwMeMgnaYcoivhCFUA0M20QM+VeRpguXfhFTRFlOiyfWPcjelP4PJxsptgc1K3Sd1z
kSl599iu6GCgd4yMJbVXDN2dpBNpHOFo10NH03OyF7wj+giJxR9yODhmeEbKmXdQQX5Dy2BI/kLD
vZRMnMNaFDePjcUREjW+r6yDj4VxPEsfhV5lS+KyiaQZhPnNsDQSpAtxmQ9Q8sbGye1UHleimad8
3QZRVNcmkmOQEb9R7VF/ruy221qiLkULodXdB2wwqmPRwEabisVc2xsCpisMQY8iASZTz0hL9rhA
+/W7YfkHO6l/UZUScpZl3VpHvDhpfgxlzVx0HPkqhda43I1HknJl0fFsXIt0u2fH/Cw1drXhWLDv
7a3DIFVcDwTLqseMYJxjLCnbgUS/KCxN/TynCAHJFXeulU4IEUFCMHszCNTuBxUUbBWXGXd6ek7U
HCa0yBo386EmqAU/J5mCToSv6e9fmGUHp0AXgxJA+SQzR+vvTsD6zRNFoCl+jM9o6XlbsjIk01FB
8ek0MqhfKdpba6DVqn8ZLN19Ov+CFE9dqdtXIRnH1wv6YSJem6KVJuZrstcaLD+t4VSTAFUlbPGt
Phjd66ETpuh49d6o376gTSBrStHxT4hlmFp+E4+zghQE/6Zq/hPS2mxjHdjqXTg2zzck9Pbf8K3X
lZd+lkLgilHczfLmT/Sm+mRAUPuuuTtdMupxobNm8U+sBZ1Z1IG0nPXWl3i+kDHCZ0pHG+MKAVZS
zUdWPVRUbOVmEDyBW+as7ObsQ1pbkFcuZaOXkqbjgsIqWCW+r9w+yVsLkTJ2PyDXv1K7/BtgBFsL
lfVciX73wmAHOlD94y1Ch52M9GG603hGkWjxuOyOMsPXPGpNbB5mowhoVzBo5Jsd9aQLzIaiXaH5
pIcQD+q7XpZyI547b6K6/NxVbZ3Gu8s2Cdm0LQhP1j/CBqSTEhSuSgvI+Z2hhvw0JA0Ovg5+zzaR
ISjnhff/6F6JRhYVtJxwPrbxerv2W7hUZWRI60CSYoamwIivRABJPqe3xyzcfPTyf+K6pzf3pBzn
+6/qaFgayjcXF1zH02A+oyz6x3N0UhFonCF7PVNPUpve2pRsCB1B2k7nL234HwbbKI94lPL7hall
xu2SfY6T1yrnt1pBGBRFPI20DAK0WtjAeC1yat0+pkQG+SzpLrzkit8urmMtEJbe7MZUky0Jx7iQ
qDTsvcop3mmcZcq2gDBhSWK0cUPrdZyK/g/ZhMBjeufWnuHp6wV2IWrUBj5AAKOHXapmpMVa9QNM
oCWvRyYJg13ZfYOxKlnCi+p8EnM1LmbidISxIKkbRX37Y4zn208/eReU6GI+bCBw1JNB9TKcFlmM
IHq7+YDxa6+FjRQUJl/ap5UUYl2j1GvmySIHKUvrh+bbQqgkgEAbuDYstHyEzZfffgw11AWCq4VH
IplgQUgK8FAfFfRm2W0/vf9xIEMMSXMc1cl1k5j8fTRM8+HM6xWr5c7BPVMvA8OOBH2x8yRZp/nK
AqdrUraGRznEMloXhmzdNNrMMO9y1lm1SaZn4OZ6S+5Nunv8hzwzhlOxxctZZOcwzXs2wLFac28m
zjpIkzxNR2UDWVYt1AyCByQTfI6nAGlYW+9/dQ2rG9eCUqKI6+BI4qTCfm4sqkRrhfRYiWaHwpDV
uR0UlZS81Ei0g1AcJbCNqq2OzaHOi692jt7/Rzvs0Yf5agtpEYv+Is3UTZK2QFXFCdq6dIEHxTCe
imbBMph5R3Zwu2OWGhpmMKmgwxT9V+TKsB7TnpKKwOYZGNFP2bacE+C1eRtEX7tpllT2lOP14UGs
NiUP7QFrftxioflL0qgWw556+Xn/DYuifY2XsZuGtuyyJDrdG82ufFjDdNWnzMKECp5n1FBElHLK
9tR3QTQgjObq7FWWXpWckwuCoSSrzY8jwN9UEf8YBzrb65n7laR/gpbIjfMQQ/3KPGznAACf83s1
aAPYZQYRo647gRx+2iJe3eDT3Z819iC2W4konc454Tk6D7d4cfi4M/cbPqYVlNUMfpXqqueYtJvn
FH5BzHsMuAax2No9/RdT5JXRlV/tyzTtFA9UOwdTcJQwSxLbrS5QKO4x0Gh2lktPWegiOF+c6M+U
7RTD5dncu20W6CruRbFv35uoewnQitvDDomL9XAymihMOsIAbsdiNcqGBJ+IlrWVYvk2+AljLCvf
i+xFn8VLgY1neovonq0Criu3MoTCtbGtWIc3S5eS974M8XdkBO6Qg0ElmMRxSnQ5jwQyhWhmxy7U
CXheDXZes1Q/kGva9LwHJ62uFCpyJzSFS+9JCmYCOqe3ijcMTsNk7jx0W3cPFcYz/q41h80eHV8A
FVXfK1E8V9H8XRY6VX+6vVM93ufcaQCrXY+K7TVKHfRT4XasXAPUFlQ/MI7Z5/X/hZYdFBRVACWu
tcl/6oAyA/V8zX/dZHNWlioo0GGjDgoj3oUrwfbDwf70httzSi+O8lbL7kSBgVoFMq5Ph44cHqdG
jp2TI7bryCMgxS0B2jgN/oFgnGu968F2q6GEXBieDehnVF0Ab5BS/V+n5YC1RWBYCbucZtlgx5Up
7Int8aJHMNIyISm/9XC/wOZGfOb/+iifDsKkMUcFt0/lHZtHUiG9eX+royJJ6WTuuJNOnCBXqRNp
BVPpGayZRe0fB6p3X6zoZj9pwSlyGOgEPTSK35MeRvlGQnVRbh+5zpkUDuu7sFO3Zz978uC3HvfO
JNceYLWFbPpHRGIov6l92owtGGr8lDi3oQXi+4V1ltOEwO9N2ZSZ29jFIOQ/kMR5pO6WzhaKXb3l
P4wGcGjsdRPSh9S/LecxFm07hGa/SHMvLxNTJhzVaN7dFvG35rLOx2pSxD9lQFL6g3h2R6eaA2bU
uiQdnjZXQBey6l+XNbpUSSIsy3NCGSIDtVTUbYlfRAl2f2ZECPK3HnY3eYBqB+w8G4aL4wzJLelb
H5lZE51BEA1tj0fKxV8sfAEzpYnKDu8PQKR5VQbmVk6nKJZIaWQB8rJ1ByilUzx06IFEHBQRbYUs
XlstFslUqDbavyp0QcAMDFTmP295HKjao2SM1WRDutlePdlnMRmrM1wgiOYhRyMKUySr0y1GsJ5o
j0GSbDh61u/E5/Rn9HJSLNoXrW8SKd6eaEspWz6A3uHp5IUfjLHbm3xMU/lnJNFIIxrX4Oyo82gF
L5HkeqC64Nxuvr9jas1D4mPC4FLfsfVjloj1DbmMBP5f3rJ2q6+6uGUFumzyhmQl/rA4qd8AcWp5
/RAB0LGdlHJf1n/tU9RIi0HgiMMb3tGzUQ6xSpwSUEOlvNNlY9vxREmEsfdxREBHnSbrYWsXTfLs
2LX+VCdmwKlS0hJW7Xkx9ucTtqpsmswNXmygfG0suR6Dr6lgDDx5Dv3n4L4DVsx7X1EelHlxw8cP
WfSQHBHGR50Z+dJynd0ytYlVHGF39fKAxTc0Ji/3JcHaOpfb1+ZfKddmKIfOI/YcoSCklToO34Al
QxYJo26xOKMi8nafQf0CN/19txl98feoU9tRaTqoKAwmffPvOr84yaScf2/3m0zPB4CKtEH4nctp
ZzINRVRVEF1XfCcQ5ktlUkfgQM68nfsp6Kq+iH/o21ImNTeTPLq1+0EVy6arrJoM4UwmPkaPbTZ7
QrOuxcu2yxJ0HHkTZJOhT9BxffeLUKMfjQFH4cc0MOnYWHnZYHNRoMB748FCzwVBajHeDC0ES3M2
kkDuv1i4N73PIGksTQ4gmBCT8fz3pl9Q8mht5Kgu482vRiuxdpH6rdV76BJ06HSow8Hluib0jO1p
5eC579HIrwWq1aM40dpAJyi3qCIkDaeBBNfYj5Av3aRJdJRKy+oRRbEFW7QHoYaMTSrW0o+xvt2h
agyJknFuJwtuRaQw0hb/v2umA023a0tn93Alaz9pqD0vFeZy5Aj+uGMrofB1PuKOBEU51I/S2UBQ
VHAhkHMeWZi131vDP8Zph04/00ggmwwfuz/8OuLOXXoqVq9M911q6EHlScmK3YlNBrgb1MxGWHmT
HtKGr0Qfb8He9ShsT07ulab0igCANkBs5qqdIoNQCik4fyICXj8s7ko8z7fbD1iwCMzYhx0b1Ku5
ybn/edNKXfV7re1xohL05SmB22IZU6GA98W7aeD5Q8pwAd2MUYcSuTNggrgzCiNnd/jfJhQ1IV8w
PZzgVHW7n+XnJuwhvILQji5Lqiyr6fXEExwiQPh9O+Hd8hMQHVo493A9zkFUtB8T8xxRd0UI4IUn
SlKCV/5Cy4VhTKHpTGpjoQG1ZXuVQVskdkGWsBoIe4177ODs4T3KKkID1xmMc6KoMKs10DE8ILxm
GkO7bn/d6cpJaJgvZhjRbZHfb3wC6B2tdNYv1hwQhAg+S5azm7Y8v3N2IXsnymGm2JfDkFCpfHNV
VHnCNWapomTFncAn7WUZjIZuIpGATV8ivK4H/p8qanyd3x7/1Xa1wbnzFhbPMAoal4iaDMYG4vov
PdXkkC0cLqvvEjdjyrpwYVihp0YX827/XyJ625oC1Qc/xEOKzS3NrYj2fyheUaNhmEbofSx2UX7T
u2OtTAamOd7Hdr/yydiwnl0ApWS8Vv9MFlqeaOpUIr6Q2hdUFkxLh8e5kGk1rKTDk11Pfyy4ZIEW
YRznDWp9p5gyncSCQoHqGzdVCseWuamGUDtWZq0JGiRw8Z4DIMpqIHikIETzp1a0hTOsgozCBC4w
OGI8bEYTj4DIMYkXx810rCwMjYltxq90iNkpCWrhIBkxUm153tsRZh+x3ro3NZ+u1Lv5UYrRQsmT
Un27Lrou3VNaeRCaGx5RL61VeeEqz8Q8rBWt4u+09qpou8bg3clcbK+IoA2xIgTnwEs+/owBrMer
GxJ6GzxwNroIWXjWlmH3TpynDnkWREpZVzYGdmMoclGdbyIAe+GSMjOBEsNf+BsC6uwCjelZXKN3
K8k7UxixQrd4+DXekCRAfVxA70frO4RuzQ6io8Ia8FAcsjq2IEIPXzFrMRa5U2wzCvpLVduf7aLf
T0/3Rv/8Tj/VC7HKp83QYWdbMExf74y9tHxeAqp1gFImr6u7oCczlpGsHY/BnIBZJGuN4VZ+Z22M
FR+V+pi9cKcLa7DYuK0/oT/KgPMGquq2JiCv6AXqaiT7Lh8/6oJiEUvBhS94YipSxPM+tx4fuuU8
eM4d7OTqfDxI6ooY/YImH9DZoqXr6MNEIjfMICOXTpOqnLXa5x9bylRBTmHCwtsO26kFxMH35nal
nr0lh2MvUlSc04TaFt5qVB+kCa7jgji0R5U4hgKxuDBNpSDbbVjv3FJz4QDur7EkoN+qwVkX931X
SBJBK/QQmcVVxdFNxtdHi+6TjRiWouE35Gze04DsSNs6CeylxoWQJ8iSdA84wjCiaGMZmQ255ZBY
7r6SltiEMofK7Bs5DaCqyG5C+KX39+02JOXMsXqo6l22r26wingUD8P9yxcQ/hHyQdeY8rnQlwyR
XBgnsFXUq/yI13BJGK1CpGcB57qYs8M68TSQeQ23221pAat2yidRcNx/Z6tb4qUExzvpIbjghkjv
xcB73s/5UJHx8drayyLjriGZ7nj+rI6wYtNWTl4NgVPP+ekhGPYK4YyTR4eJITgodpz/w5oeTply
Ijz3Cb3r/FJax5EX3t8SmLF3h8u9tfDf/CfNx+Z14TqtKlc9q1crQmXDEljKwXByYSkJeO9n7gek
zzPWkiKkEl3S5Y/LFW0swJujFq5yCcBnlVTmU1bd2Hl5S3/QYJpMjn2HZOBYvF2keC+za4OOMGar
Xrj3cCobHtl5NXBxuO36W+gidiLUOCDF/JB8diewNx1YQr3iznUgdnwFJrD+fqo8ccMLJ/B2NHHQ
0mZIupxkIbJIJlUiuY4N6tPgL3w2m+Di5JXimrHjMIswXqtw+86e3gTYU1StZy4ekC00BUtZkkTi
wp1E6+pnmxdOWQg7tWaSlWm3okfUc1fu8neJtItn/NUwMgbaMwoFxIZqxkQFaW8YdpbCteJ/Fxgi
Nl4tDdTXdkrfIiDHPBy9iR203RBpZmggO8Ez6xp0ta+oT3YehtilDg5PBWyfuV+zG73mbItKEwYx
x++exgPP7qrzIRRps7NZthgG6YWCLMvV0Gix/wSWDWzBrRQgRQIAYaCMgSTgMAI3nYtEE+lz/G6I
H6tGUJz2IUrGIpp9Y5CIUzFfqtaqnx7+Qlmo7uaY36RIlstGnPGoFGE9vhpjpv/dxP83Xsaf8p7L
2kaF2BTvrOGYN/U1b7m9lmgikZAdyXu5FZHz5Ilje2K8l0pa6dgLzOSmLNvMkQ3QNc27mpcQMIg6
wEZjU3kPMvvmRiFI2z1bojzFe/J4ZhZ3e1EUE4dfl0qPU3YboNZxlVRmH3fQefGA2MazddgE6EhX
j6BxOVL+E1E6LjWehh+/+5eiyIbTv+BB3TMGRqyEpuSZi+lqBy/f3KAkfyl5ERMQEuRpdC+CovYb
e/40dRWapgxGQShzixB+PNaUk1ivFxmcxNlHz1tICmN0HvUCupGFcBkYzzp38uAuYM9c05edtwk2
VA0NBsE8l2ESDKntsDVrpx9vpv75eT+9VU+Dq5n1gfpyRdA30rwEvAtwubCvnQvWEsy62FY3gBKt
tmkKZ9NF/f0OEPRChmCKMkB6cXMDOn06VixI2pTOmcqs5Yx08E844nRUfDPXKApOzZHGbrnicrHt
xBf/BNe/oS0lloheupAiqAKPhnv1+1OnKDmo29rz28843FEsIuSAxm7KSMEvc2IqnWvGmUkFF5qs
nMKNt1zk4vy3mxmTBK6Di48rVqn4EseTp6NYWX/m7K361mtvAzPThwh2ifZWqHx/XIE7UoZSAN5t
bz9a9RD8OB+5RZax/RxWQgqyrpg0/CUNGp7fJePJGuMF70i02EBy4dD2y6yK0FHyL7ip9ooL30jV
Q89oHs3cCvfrxMQj3gCRzqe3ydXWHEI9hDlO0OLqesirfCVoi1TNOtxvGtAVMzhF+xsQL4STldVz
3jxj9SaaHXywUnjt/WrnA6VcbhFTNTCRC8Thgw3B0XCje1ZNrS8qKjRebNmOXjA4H4eKJuySFCwm
KvN1uKlyTml2Jt/d/h1saJlYrSHoRWxgL3mC5M3bxsbZPGuTpo/nBC9jP/Yepj5dzJVbF1uXtM9z
GWCGoi62LvZ+Rh88WJVs/FBzIg0fjluwQ8wdIUFCuJzGUq09hgkSw+Tz7zS1OHtSlJ1tx+PBKJmX
Q2MKbScHYoxcOt4FVKelvtA9qtdZ0QQei7ixdkh6PBL7jENXq869BE1K7/JstqBJQQU5pgvnt6H5
QjijUJswcbggkHwdKbAAU0euv++iGy80dr0As1bTseEo07Wb0xfV8WeVZ+2xfXkamv2SzN1Etgrx
J+jeN9pd89R6XA9YOgEVrE9xgHw7LEfyqTiVKXX2bRxdgzMvxKQhZDYOhZd6WFWUTvrLHQrZI7LB
ziDeBfUTigZ/VqUB/21mzRJp1JpoCMeFwXahblFUP54C5qxEqHx6TY4lHEClnv6ul5VDxdhMxBjZ
n0OG7pFXvhJv/rv8s7KDkaVjq4b0+scRsk5s4lzldatz5cn1C+GQb5D5N3vgrq6NFnN7QqYHozQA
1HdwWMdfn1IfUyoIaYbV4VJtoc/hu4L8b9sOz60R7tGS0LugkkbAHLaY13RK2Gme6bqVhyaycvYW
dEM5S/M7xS9pJHh2ZQuJNPy98Lw51SeJXdN8kn6m/AwyvsR8mtF4v4V9EYctjWgN033Plpa+mFpy
2RnkCi/eMn17hfbnKVDdn/3eBpLNkwy6tM7niJzosqxG3t/n3M+XMe0chVxgX8kdjBVCVqJelNeR
p5IsC8ILeGk3Dvfq0zMDMPIIjz7iufNzLgJ4TZfI5hUTMxmd/xMjt353EyrpxumL2a3vAnl8R6CS
kyVPVDnqJTsQ25BG5P3S+o5/mcPozzt0sUN0IXJbXAodn9b0sLI4+AOVlTG229PWi+zbU/YcDTgx
Bhwk6cwWYRRTSUA7nONQGfCBbeNMD5+dW6NXLl4BDxELfQLnVdNXm1Nu9TbPhwnSrN9q+OVjEs1S
gY7xb1MjvoHF9mFT4VErT3G7+z3VWpT6nVjBtMWjhUcwr+btzXZ014wXP/LZ5wVAwFqHbfCZ7Co1
MzFD8ay/6hLoFQc0/GIaWa05lPOMeG8UdEfA2JAAt1xMZ1svI9KCPZwo90QqaHb5GvHdAbNgxICL
4x7smN8yO3fuQB+9fXED1AGi76hbWjkQQbTKTKfgdeO81iCnGS0n2nMwPadQ4LyBqlDUS5zsuzY4
HqxmH+CkJktQhaiX0sTEmJQUkdeBtpKDnDRwnSD9FSDXzMBX0uQg+aGvIDnq02PX01u+iCbdGMTm
UNxaluF/yP2CMvhmIFca3ZqbT4ofMA7B3aAfWIyH0Ka+HNXLos1ORYNKoAjX1i3+L3mQzUFgjDa6
rm7eKyG76FVaYilE6PgUaFhljMHkHNceMMcMmCjubdHNDH2qUqFWWGAO2FV8QJJVYu0mYSQbuKNU
JH9V3Ty0TnN/T2Hw69fMjLnVGfskCzRqCqdrFcNrKVXrGoUHAT9eBMrW9+ldXXZ+waTnYpOzUuZF
WCeM/lqeMZAS6ADJkWDTqrE0+U6nD2hnGaSMeM+jiPZUeMj8X9Yq3o0RIesROxoRGXn+AAm9GuJg
PS0Dc8QgIzxB0vR2BdAsqCSV+9iU8wnaio+D56MKqzC/I5eFvsZs9Xd+M/dH3xSeNzB7zJikIwDi
VvhiPfsYoLuorDFpu4K7Gj3i7HzVR7qXW4a+psJ8N0bRGA3a09aYrzGY2Lad5KuklHCf42xWxnOv
BGtZ++TiEpKD+5WR6CP5O6OEsIS6YqpjH8INqXOSxA3KmbwIQR/O3c/petYSjgsVEMg+hwqpODcE
QFvhhZvxGrEN+sFPjfhsNkgYHeSzM2dOn15IKfHEp5SPiaiM8pK+nn7AUydd3PYm+utyeI/dT+i8
9ZgfpIiDvmfIg4L5AoQBWek3vQ3qjhttWpHOSRDJJq84cVw6ZzjBL6GZ5uOCqAGQp1Ht2K+aKmKl
NKRjW4INRcniQ4iRjTs20dm8AS5tUPinzAOpv1sV1j6m7FDkKMo11iGRj1YIZwbk7tabs2JtLjR8
51RWTIzhTasVYd7eb6czvkMfpMUbMDEKxbit70/XRzBglRon56oGtt33j75ci0DPRdH0M6nMEB52
4AunEZt5IuW8hTwXLa8i256snqjgqhljdqf+nB8spIlOYLRCVLKqtXlSTPYx1HmZVM/TddwhGdXU
2pnGOXsMwkoVci9Zth2V3ihdN2Hbo9AYENmARBp2hDVvZGC9/hLoU6R2up7kmALzqmrzN5mS7ZPP
sT+V/XIcTZQZFhCcm9PO8CBDJyqGR2lVbdFpdsv/tGGKNjKtb99GbYlbiB6mXLUF1I15FjOnTy9Q
PwnCi8rR/Q4GndRwLCxKc+u0e/4gl1vVE670dO7H+WDl97BThQpoKAEftXjQGn/mb717eAOtYkYi
qbj2HfMUCMLzLFaiDDsxD0x/jal6XmyQaF/WwOGbhQ+7wDrgCd8WwSwqNMgWj8/rfa4vG588msGZ
9CegV+jYUp+rpHC2tDq0hA4thKVW7YAmLEo/RcpQM9DQmK8/1oAYn7Qj6te6X/PZ5kTl0WE8+Y1G
yKb0uFl2sOmV5uGAmf0BvBq51Zl87Gz0D1rR5qmbVsCJsiVUIgeUUKHaPO6m5Y3qgtiBI625BUPe
Q+o797nBvPLqyXlPgvaVWapY8q0uzA+GYD/QQp7wZa9D2K70Bcv+3fMEsAI3ng3PLy29ZEVuN3uT
eK/oYrWStSlSwGhNwnnGj7Alxy/OHqkOO2cZ0sxQNMwOJF6ZHKAUrlDT86RBCqPk9AvQYwApsTVn
SvdfOp9pjPO7H2vyndRM1FSRYHj+aHVN/87ZHprPNxtXw7A+BYWOVAquXO7pG+tVfQdLRivXww4J
mVbqQdVqiA1GiyuEHWg6fNy4jK1fFMYUu7iU1BSvCkuZrIss0dZXLbxSwmUmbMCCVKnKcUAqho98
cIWwvwQehq3FWuItDK3l38CEArSKKGNlCykyG1gmS4MV+W2nFSaPWDtHbk8syErevMh5aB6lfxnL
HZK7XD5sPx0+L287GDF9rW3dxBhK/aQ5dpZwoy1EqaBYiLyQTsqU2kR5c5asW7m5YiZ5tfdITpMX
j3J2wQpjh+oupRKzfJ+TEmVzUbkA3o2yn8KqwrMYW2KEs1O0jFj0RQgASY/CPHijsFnAAWSSD9Kw
VSgz8PP40acpI78BdxKhrflQAd0gLf6p4Bvb5FnfClWv/e48fXkIe8aLXq0FXeCqu4ey+HgDzNog
v/i8zxVhK9FVhjoJTgEgLLq2XaIkE9bya/QOAQP8WZO7E8LnHCvZm0c5DuJGIDa//4025gULfHFH
ksL1d0zIMFaPhH8I/Eulwrp3uz+QfzzKA3jzaB1/7lUdTtutJtg/RznMDD/L86NpGdRaLitcEmbw
gGBXWzqTfbBuuMMAuSDy1bzmGg8h9m3wxgtjlOTqnpX+1vw7wIav+k/Pq0Tt4PCbLQce6Z1MB695
kvMOQFodPoEkmLv6xovtzKucJnEViX1hb8m5wf7hs1udknqKKrUSJDLgys5oCpXgwd1jfx46d8h1
Pz2OEf97KlXxKKJwrxOwtXkbUriKTB1vwSl0x6g5RlJDUXgmZEUBS5BqGEqFPozmS+ry+KIJSJwP
cFaLhmsM9ghiqK+TTHt4EAqwVQBe3l6qxjnMdfYzkcAJGzdrzty7dFv8AL6xisLSzc1vY0Kjo33R
93nD/9i9gZC0uQjVaXhcvyqCJUVhZRc5k53gz0IuiKbwN6KWs1WSCCs9XwgvIa0hCzyEggCpOxke
nfuA/egkZ4gxHDkjn7KiN14Si1wT297BRZpm/kCRp5rPX2a4hSXlb4JwNSrlrTWUHE0kVDMrrsSs
w3/rXByF9CbYY0H5cMYDyRxwOxnE1AbjBGoWI4OwF/G5uZemcgi92ZJTeqzWxgD3QIcjYJPlHXs/
5sWiyT/eFBdN14kjbloZ4eJW7XBupRNyG06nTbn9hQNfNpIqewnPrxF3OqsXY2QwUFgG+j1902B9
se/Mt0KTxvkv6PTvZacYSJ4eT7zr6zDeXv0wzeATqrMeZuJfTuMDLhNe8hCGHz3YJ0npkjTTFp2q
yNFYn9UVvmCm72u0V2ClPCi5yr9ieUpWrLCDHUkgxuYmrB0l58odDCXtsKusJBrB9P0+CVsPwKde
GnjCXjwv30BXGOaMxgqjAra5Du4CMSEda7IAeGmQsrjbcDM+NUaXBE5heI22nzkJRbw3VPBcjFhY
xbx+9vC1PDeaJ/g8lIpHbWxUvZtOJyWri+cr+75Er36AKgRB8c6M5xL3s69tqhtB3IotQ6m5qjGV
zhe7okhimxUwVzONDD9M5RFXgxHFn7kCYevCkTgFq6qU81CTB/ccBN+tDDQXQHhjykPp7CMNGNQn
NX7KkbrqyS+PtBQk1p2xy4k1xhgSnM/S2iKguFPRIFmNiGjbKFaas3aDBCouUEPQu3SV/5N+gxuF
uMPzVTQmam5ACXODIQRDykFPkiEF/TcvHNScED5E0FutInRbixJ2bi22lgxpile9nn4urlPAU0vc
UDuchiXRXQoaJpjuGqnvfRxLN213Sug+IB0DvlmPxth3c0qv78zQ//3i57Mxt10AbiIEoddBRm2e
n7XxI6u5PwlG4kb5duP4nnIpJ7Jr865Hl2e2KQS5PbZpFMmyuGd9t5NbDOUo4+Ign7OOp42A5i6a
kZsbuU1/bvY8GNyR4vEJytbeRvmoC3LuWYFimZuufupQdVfUj9G9UOUmTd4M7crcp4C32aduVUyu
ajGqbONAAzbKLkA98bPemG5r197NIQVWTleOhFiyjjXvco0r/N9IUUIlSuq2Ke8clxR/w6G0dqos
mHtS0CBArjByUf5POrZDuvMAnbVan727pWQT3FZBLnQBSAnoQ5a/n5GL/rqW4t5+es5FwAO2ff3U
P0f9Sa+w9qYLW9Ies+n6DEDXDUYa88H8n5mScwe9seBspPQ/FSwHQSbqmMIjP0qyuDrWvobH25p+
/LR+s1F7AI0VOOcNr57ABfK7v/S4PDwUU7VG1zbSnxJymkCgnR6g0FCLfnMYKU5iSSSjsx55ut8X
Jq3g7n6FLbH8vHGMBdtxHijtXVVaTJq07jd87CNYhQLRlyVRuE8tWu1hCNenzKiFe48e3PTIJPnU
8hrOxBl3YWtO1135iFkRXDBB4euuXZJB9K4ss2Ng2UfPFpl7BlQiLUfTMhcjUgQelQBbyP8A7f+F
yvxX2SyPx0gHOwOUB/DN0OiucvabR0I4l3d3PBom/LbC+3p1eS62XZ7/BDA6q1emfg5dhnEvduo3
VgboZE3IhKsFZkHin7fYp5dU3dVA3HLYNru0RJywSTfi8JR8XAlzjg5gV5bm6KEm7PYf4N6sgfIS
/IQeL1b4wn/p13kEWukI77rii1aJw7PncBtIpk0XFLyTNj9n1MZLYmXpiC2ua4h3X0lRUrQJ3kR7
jhSmgEeGjwTjuoxsRCp/JSs58iiA0V2zRLTO83GnD/z5I5w63NbP26bxyz/g4iPbsiWjxGwe3dO9
MPhCWSGs00vkaeH26O/KlKx9H/c5pivkpTVVL1WBmfstrdFIH94OMk6+76sdKYqac6q5en5jHQxw
pdbBWNQX8O91c9Ijg8BgEd3OxsDHc/LtZULD2EVDyTyMy1b5b5UCaNdfFhI5804RcFC5++lXFnZL
Q1lj0QGN5VzBV1FflIQZ6cMkVEKvVxLIN3U0zmv5LHj9VnzHH4Jf+D6IJaXSMqWg2iADY8nZ+G7P
G+RSM/E1VUexnNDJZ7a3n41YDdJykhl7Gs3L02tBmoj8TpD9iZWsSyxrkPsjLN9oBZFSkx14Nt+o
XT99rwyi0KF6+8NIuPIPtstTv1WVjx8OUK1W2l2YrThfmafxM1BiTBDONiwlf9uO/Ce27AyQvu5t
ShOd8XUhJfDTfpGOKzsHGEfO/GMCncEvx6lQBX2ymHhbbGhEXcUJyhcZg6lsOahDdyT/ITAg3f+L
uDBl6pX2u2hyWtwBVabIMGWC7uDRHj/xvCRMSZoGk4xXPhhYSF1N0wcZlPNUNCM/kktZxSECV3IU
FfFW9JfLzeomMqAGXqplNl6s3ip/BgYYtcU1QHOyFtqC6kmgPaQ37SEPXS5jyIVcrd/qh9bmokIr
8AaDv/cunv+NoddXTH/upUKlVO8sfaciNsOhRxAlnm5NbYvJKGL/Xl5XNS7H61zgqYTsSCoCadz/
wLHinxPBQUtlfEyZ3WtOPX4glBwGnqQzRsyGqWVEj7SXmH8LW7v+YgUeP/l3cTIcVt3vinksMgoC
UkeIUHFGB1v9JGyrXUaxEF/T6TkVBMVbBjHnZjTMM4I3eeW3i+3rpVbSRXy1KjC2cKewvrleN9V1
4cOySM+37N9iRiIjv9AqhjmhMCgl7duh1JQ423qOVwVXD0+uk/J5eJVGpsOVEV0e4q9HN8KmKZVD
1zpn3ooLeOXj6Qy3aaSbLdn7EZxI8QSB9tUkamyCMnX4VNZVkw0vmIBSRLZCZzCgX+FAzQwebial
cMl6lB7MTsu0Sm0VoOyYjwcHe+6/Fmhul68mZBLOLWFhqEdEMamFfo61kAjYpplqEg0m1lqShVOz
zcEWXAgTzferrxtZ06kArKxXrnuhfxEQ4V+gjn4ccBqermYIDrpruaspa7R7WFqyXMPfYKoxIAyn
wTuOT6GvrnsbZ/VrTP/xDT0S2S/gt191JQzgPWQilSScT6Fs+1oxF92dW54v7HfwjRK+WJEFHow+
zBcI7Y4tjV4uUFVl3E+vwAesLPNdv2JvAkL7awhIKFQBrC/ad0P42q5StPgkmyZETZeMJAHFoWbA
rYUpmbNz5yVW98MX6H8dLJnDawui9x3ER7234EipI0xY1MQux7QF59xugAfVxZAFNV4TJC/xfOnw
1Gn3A0f3g0aCBnNjQBQCb5vgKDsTyti+2OTZHJhjTG+jhLT/BugEdSBA82cCQLHe0nUOsJRDKh2N
8jtB4RXOpt7GXflgc25SBlq1zeiEQ/9nS64pfrT7lBiaraPi4KqtAjQj/E0l3pNT3JCfOmy2uYol
52WkuPmMkbUocwv0BH7X+AtmQmt064wK+aXDIVqr/nZZF1XTDBv0rdPjlG1FwX37WD9DImTPOtFC
euwKrOWJ+AzDiOCjBBXuvyM1AU5zws2iHVd6NkC5wZeretmyEUsuDH/SsHzCMLoUP2aeiDJoiCLB
h7VKXQmaQ+Hsfqzb0WX5HsALEAW3uXl4YQq3J0dh5Bv6HXtSYwYuxq+rqDLdZT366aiZpbJDSUi5
A0Je9LFwKryDdJg/xViaygYITd5bcuI77UEyGLecfR7NSu1hsPs2EUxFz6GBOmKPP/j+wzpNpkJ1
0+KAUE1kL9z4iXBwGBwrCkfQam+lTEMij1acJ9X59AgGdyk66qQahDDN1fiEm8i1HsFCY8N9QVE+
XyYondhiAWAfQSgRI52gY3Kxg7X1jClozw+4F980rqZNovTMslW8XDLOnsBhiNs6OyK/SQse9wZX
XeXow/Ha8+NZcLkIqIR/6I5Dhgl3tFGmGNytxwhWPTnR4XURi1OKYaRkb8ewh5sA7Mj6fON4FiJt
//y1ndpGYcOT/uqHo+oVM5ELWmJ1LvbJ0i6QBIJV6iq9+fb2sX4LfqMldykSaV3tpSKsTJw5dLA+
xDobzl5Yw3oc5ag578wI0yAo/NOUrE2eIjgLqD8yn8uKqxRheRNpuamGFwl9e7IgT7bUiRQPCpnw
xmJHuSYJs2b/kFvjolgvxkBGkPPWsFu48JyrUb9Aq9cr6KtDIOcFtaxBMYR/+dWQmgEpdoQqv+yH
i5ijCaaerft6etcHoMTXV0ZjjCiyr2nNNpnE/r9PYV6b48aqMjJC8/ueHxNcVUl1huid2zxZGAAu
LLjyEW4yjOkCZDecHr34wIGVcwSIcTAI72EX2537jetSd3FQtCYg8LruvD9BG7EeQzglB3GK2KTh
BseFSNRVwwVLfPGKY58TZp3cCQgxblkYzRzT/uDDi3gDIfVMKWU8L6xDtfXNZ7em/wwsiPcvtJn2
3141xNGVBOq9AWpOXIo8hXU8/dLjOLD19ikeOu+EoByRmua9CldZhHkBwL78haZajv4usSRjpKU6
dJ/LEJkdHCi8k/n0NZshi9gQwlh7az89fNfem+9tz2vDjwWMwJWsGWTXMUjiJyI3tZc3fn4OfKYT
J/0XdK5PvEyvJdyEQm5UhqN0WUU4dRsop2swDS9o85Z7Z8+QB6VM+3cE7IZhFBOCDnKMGwDEH26Z
i6nvyBw67G/AbHenq6nUJU6y6NsXOQsPgG/fzA61HWB0nX67ckdxIRub3VCn3p8Q9TwuLX6fcBo1
K468P5DYQ2jXQBBK7NYP5znKfPBzEoCF9plXeUwJN7Cm9jhH7zB36IeqXjCp6MF2eBD/fG2gnaoi
Q0N0HfzgF4V7LcCZ4T4ESRviiUGqUHyUU9qqbAH8TRXvR/WXF0tNE6cuuEUM2pl/+x1CiFfzUEXf
Ig67SH2Xf2oFwdreRKUWuwKVcBQAR5kOEUjD5gZJqyeqYZlWs+Q5ODRp/ErvKbSygb3PUD0Xr1my
69xgR8VlralUvjsdQsU80eIqe6/+eT7uAr+Ud6VoaHsuS1iHo678tVnzDY5QOakpRSkeXVXugjbU
d5dzZIbGjDXCgCJpmX8C5/Tb6feB1PQlNtyQRY5WcmOAU6SWz79leiNkl5b/37OYyv4M3w5IkkFo
8CN4baSKPqbeqSSsduM6nU1o4shH3qkaMV+81EhNDKHs9jL644QYb+Okc4xykzDG+NJ3gOfJH8pn
TvK/QZWjGV9xOMifRuNekm9coS1T+57KEq3j2b12IzZlRxozwHNyyt1K/wfUiXfTgpANSk62pclk
Z8HDxodeHM0deZ14HxgMNKinnr6QXr1nFmikE9sBsZEbf9QjNiakcMzUYUBm7wYLTIYZ/dKO1wsd
tCTEMiTYxTFvqNkkSjvkm5JmTeXzC3ylOqZ1kNFR/UN2s6Q+iWBDjDl9zoPslJX+FW95Y/8Wi4hs
pDNg5/fYS84BgEFVLy7/HuE23Ige48ZdxXlwRuvp5JLC3+cqZ6+/q6eTh01b7wqJgWTPtPZtXqxW
3rzNNGuoqJrg6f6M0oDyoG/GT9nNXbGRP0ETkqvDhkqu5WSeheQjzDzzlNf/RwXozUZm15GtvHaI
nXeYDpOCvW2zAKNeBQNGwKQAGlfO0VQyaT3WWjlQsq6dv3CSGoS02OUm2gfQdlb6e+WIIYzPiqd2
rNTjhJThYYeeQDe8tfXiI8YbhMApCb/rfszCXfHGOJfXyl0ydD5VdDpT3dY/WLYpq6ZIdL1mrTzm
OtxcR4fi5Cp0YuF423B2YlvdlJ9cNABGo9Elq4WEkVwVp0jSN9KxmkgPYTRtWK1mZ2iG+DLUzEp2
oL8w7BpcD9jd2N3bzYkqzdyZdhSp9xfv0bDv9laXNiWUYvvX4SpSttGdALXjN1SS0Ayju9q+OruW
KKNsHPXePn0asNl2e0CVjuz+dnkrgVwX6RUHXgcJRQJU3b4fWR8H4SUPTGi7IhsZ4lCjVcKtW5ib
BngXcBRpKXEuL8rtB97VHSuMgDmI/AKnwjFsNbMERgWV4NV0Ptf0ipRDykvvujEla1kEQPd3BmdG
yUOBmB83fgohTZmBJpi10v22CyFQ4e0mDCtzo9s80uaqgoDCdD4cXuSGHCqzj4RoaiynHnc+j1uE
ujsngZK84Uh5NHQwM9VUl4TAdPt1GvI9PgaGyp7V+PsUl5h1u5sLTuygS+tGrbt0R1D0nAKK+XRu
WoKdbpbvADdX9yFgwZ65R4YD2XSFXkyRlgyEvcNnx9b8GC0pMyYpvSfd5TJcpbCYWbBgJRCwMFco
a6Fcy8wk07Xxg/us3UCgjHMyE1YJsVMOO2KqjFhfSEMUuk+sxdKgXagi0gHaa75rBb2EXPk4Jqsc
goYSmuBQD6Qpgdj0d+6n64j1/Xzp2vdpbVneld1fe4BjFetdpxQfN0MB7NbW9UuvNlrJme3DTQAq
9w4yDiX2psf914/IpEWkPIfkHfe2bIQlrPIau8IAr9WPV6c/wVXbFW86f9FCp2lpDGE/JLLLHr94
UPAiylivtbryoJINXrd7BXyLUB0x0J2XeO/ZLxFCmDTdm3mKAYNE3DA7br5LeGBsRilBkoLwGc2h
+dd4qfEwzjRcixN1Rf0LhNE5aUzJr5kbtT1TFhZ0NYxF+o95f96rh5SMGuh2wCzWsvd+n7B8uI5D
qae2Zs7yUyrcHVia0XHf5TlVbO4q/p/uY6+qhxY/TjQ/IKLQvaEzSrMjZNSEcLwwKb9KJL26U2bU
vJyNMRGu7caUEGfuI+6h65DUnmoR7YanUhHmEjgTkXbp3q/Z5LLntyzsGiC/w5zV5fiPZ4bjzifK
62hblYVN2y82csvHSP0pCiDijhsHX78gZw0kNoP4nVq6lO4hey/NHekBOwigtDqqH/JE17AJy33j
W6TMzyM9i0AH4mF1ICHfL85J3SyQY/BzRVBzV/xSuhqm2BuD45Hn/IIYPImvGLjicjwPhoqGPQhu
5R7CJ94pJUkmvWA8opQN/TWaZNpQBjDvjMo6fYkkhSA07gZHEzdkJTwhLU48ndNYInMrPM8fa35G
sH/tARQ1etM/IO6iq5hU/XY27iRK0wClBR1JI6VhNOr+lOr9fw/8s6KpQjtV8Q+bubqaxn71y1dy
8h+ssEnxtLdPREXfkt45EoOltuTY++WLibvYV/4wbu5lmB+OBxcat80ZkAF5I2W/h78f4F0GWdpq
9rpndVMKlnUwtbebw5hX8zKY9WD+9OqdBsNXs8qLJkqBaR1B/EiGS480QJT4KKANnvv7L0gCDqeI
vmRV80Yh3ogR44+27bZzyu5gGiCAWHtVYNkmSRA3uN/bdHKR6jGVau34K0grrKhIC+mu2d6KFZY4
R03jOtGXj1km7W2ZDxzgK3SDs6EFJdiwMQq2asZOCx0WnIoB1V07Vl2LeyGQ/nCRp9FHdklYjpZl
AAd7Ut98sFcHI7Nt2gC0r5EcFYLZqHcrsLv6EC65QfHHGcgOjOJSBGpTXGocmAOSuDn5E6pkVwBx
wwaruPxwgpnLV7tL/1eq6rTO/hQgfeYk0tuNPpc/Xwi/UmrofPXexnUpHJ6YaBhNQj5FQmnSeHMC
Awes7LEUmA+Df6gD6whVDZBimCen4ZY/jecrk4L2kI7fvXKCxz+TCQdVY27+dak2sTAYq7wYhlTb
c2Whsf8NLrL/isD7rEUlIHGHXu760Qmgo368U4sVz7Bq5LmfreCq4eiFK4L4HlyN87+dHW/FI908
MMmFpwmpDwTvak+vYjrWo3gfUC/0OQiyuJcgws1IVZGVIfRrzpbwsylHiTFFyiFfrcxLikowYq99
OxO7LbeKOZcqEmMOumUDK+Yjq76dMLj/EMQ8wnFTsldh28bb/YV7hrjxIZWxebmZm3kZ+xQIk1KB
EA48xv14Rn9d/prBXyrz94J70uRHE3WTKOo/PxmwRc3EVoztFoh0L8rFBdbs+Bg17SyXJJ3GnWsj
5nWMMb05aCWxKb8ZTnLe/by80Yn6TDBItH6XiqTS2YO2mpMpFo2iGjHkdjjV9vURl+N7j4scYuSu
gfuDRiZh06htOe45sKatTtZsuS+LbwqYe+w0QNoxQkpcltQkXjhWT3LFDntUW5SDS8Nm9ShyEm1j
V4lTiMjEJ/U8kIBy8N9NB7/jWOYqPjj8G+ZVFsHCZ4fIlWM2Hb+CMjjEeZ4tFIx+TCtocSK4lHub
TT1HafcysjEcybIjTOEEfliGUbIvoCMZfVPf3ab6RqnG48swxHhjrYvg1Pe8mRZhKcvf3YAtBEVu
eMeJx/PNsi8SODTW3ObkgpGI3DpOYEDQm5+OAx/G7IJ86kxrkOVwSg+EpZTSF22xU9zfSKEppPBS
BoTJHL11E+7h21rCxwHnrXMyGR6kNet379ZCDWg7VVeU9dMPIlbth/CIUYw90Fe25aqytr+i116A
Xp7G8e8EzjHUKtSY68SI61BQfLmBPza+kWX5UDUSCT+XAN17wHffZuANRO8Cd6/T9Pd0g+WHwY/V
OYXN1VV4w++U7Hu7xKbeWgUNlZc5VwjxBQ87tFq1k1cnblAaaVvUmVL44G4n6LV4cL5ZzIdyepOO
HIfbwdhLLd+Sstf34cdPjQ/x2E5OWbqFhXkoDUbLINuD7P8K1q3VIa/w3zjDMqb4amqdm/fmmgRh
bFVhM0CLDWQi6x59/C6I2ghaDEEi+kYKxO7yw3LwjYu9l/kVavYU/icbjcS+fgUCh+D/Zeyo+me6
OKKi1JaIyL3bE5UE647FKW+TtUt3unhEbGxeWX1sxCueLJ2xptuBCS+xthfDD2WM5QXfupaTASuq
L9KlEry27Y1dYX+Col/Uc+jab3q+rMetfRbYWNrGBIR0WfGVEr0bpmfZkW87rWRB0AOOgQEAgHRx
e1O4uSJZVbz6hRXmEeFGPaq8oRJJwR3AGvIRN00lkiPiMehaGapAWqc+VhuSpKbKjikWRIwqS0yN
lPzKz3cpZdn6WJLlMAal/lK40IjD9KHtZiKjGUDfnfAJARsTgMvC6f/tp/VWloDuzcnXnfOu37wV
yyDz8leTrWRVjriZVO1mzy986q2GJdnnq7g0/FjNeLvPL+UbWbD1QIe0mzCNFSbmgPJBXmNmsOfA
ZIzvn6qKUyr5MQFJGl268WHleosPqpzqC1uQFWfqJUsWqSyskdbxWSvdKtjuNeZ7TsGcfU6AeaxR
VyWhJUkDO1YE8IZWdaOa4nSsjlMmVcg4hA6CWM4BLVN2CjDgvf4MC+DE8QAAL/uIViFznleKUlD/
DSNydsZwQ54J5zscLWhc8ndJNdfUoCJeuPuYfwBV6ZKlxEOM3AJdz2X+9pesrDj/ISy4ynjJRcjD
eHfHCCGoPBW5ClAI+OzVKrji+Ps8pmUnLc4AzIJVNc9BNOJSZxn4vkn/SnQTBGCPkjkAgqRALZWV
03PMelyUEH8CWd/JxHbGfsVY3TVuAz282y3QUToexFm8+qNP/RELe/GAx6XYeJfao1WFyVt9aDTj
WZVFue0blUqW5auCE/7h9WIO4C8FdgS9uRGR7XScLCNgqMWQ1u+EfQSkFGBfQwDTC/6RpS0Wugav
O3oVDEfzYJRFPxmnnXOZBOh7ue0rfjuHAYmU3PP+06guO8pmr9fQHT7juN1TTZEUdt6ra8peR20q
Hj5W7/Rcc6ssIfBRAPl3OICrgkvb/JsykH7q7RuWcKlqckrHJcW9nU8G7HfZBy1Y3oFvoyTuXqOr
7tJtna1tDWBTVu57SJ7S7cacfthSs6g2DLtt5Pso2810FqyXQRI66qZeXyX2KVUIvzFVHMbOGUsi
4QJWKAOLLj5JsnNtjFTXm2lMrcWoi0Qdd8kNNIZNtcbHhX5bZBw+Lk04Ic3FVRSp2Ys/4oKQSpKN
ZTx6ITO/gMWpTeL8EiTgWIOm1hhFbLWsZphPwvvSyhL0C6rGNGWdQ9HgLsx4Ww/0hywpfSaiGuC7
sNmU+NDsDy+c9bPmmugtFCedb1/bfLfAvBC/X8jJ8ATcl5ekRMpwZbcko60ITrIzrqn+MfL5affC
XnKfjMZ0yDVAnvnEVivrfuWjJssv1KLNv0zNM+nmakTKRFcp7/2EQSnFAo8XASM/8f+8I2No6oIP
KUuRC9VFeLN2sNOQZxmLzd6Q3UZxK6fp2FSlG0fVQyID7x1HFstYE5JzyKtkB7n/z8W5ysa9LPcg
4xFownGf0l7XBbEY0yS0wdkercuP7YenkBkGioOxfYhEaUCLklLh+/QoA/0FHsyBEI9K92Ao+11x
Kh9m+AUq06KOyVoBslLH8Zx8gOmvbDhdk8ev9Y+/aADgQeg9egtC/StHO2begtBj9BUOk5XIxuM1
84eo66gATNnSmZ8JKE2j7OEUNcITaUm7Qz1KZszIDK84E7fBBqsKb0jQhm22HZkthawBbDPluhVT
R+SsHbaNAQqw1ynld1CWY6s7fxo/RWe2G/fC+syd2FjrWQI4O0Phq+JLvtME9NZXJ5Wm0Al0VtJm
SbDdRdgVO45vZmhB7vwfrPbrI6AuGJQNFpkAkx8kPVP0T4FWIlX6KsTS4607yQYu6cS0Be67d568
zTOQoXZKWYltz82+Xv16H74TP9iByB7nYCEYStj0mAN332FH+Q2R7yLHnF06IN+Gn93SOxHF8BFK
PoHBCwHUv3wseL63DYokigMYG+YkANMXqGPnnI37QsHnwp4Z1pmNchFS49eWjy8BsLO1JBptRK1H
/ij1Vg15/BHgZFnMrvRJyA+DKheA2VlVmVu1poRa2S5EZsdoej29C3GoSDpdTJ7wT3tffiIjyQ9O
lOop/BVwNwj1VeMz9LCEj6jsEO7nndY+jcLvP6gY34zj+4X3fI8F7J4uOk2mCGWOnPQh013mcSHG
KlzkWc9ICGYnJ0B2rFGeLlQUQQN8NrPh1DnLhL7ulRVZTXqsQF3ZU6TwI7OXfB5+eaPNlDbOF83h
GiXciK1rxmlzX1djH6zzGnypVzUpjlAuFSjiZBGnQa0yAqRzfNax3W7odFIqPGo0c2uQP9b3/jmn
1OE62mCyprsmd8ugwh69mlY6gNnBsh4PkfvRVkE94H14BtTGO1gGOprwRzyXdYXf/OX4hYi/XO5W
6aPHDJQ5obAzbJR7H6+qQEjgRBigfhVyvwad5ylovlPtFfBqFYzxOAhtctcOyor/oHo99zElKuKy
aCOYeVE2+tSljqPmqgDmOt9PV57wgSWNiYhw9PKAn3E5vVTpcOXyOB2WYhW0WOimqZdKTayIy5Wp
3fCthMTeaoREK5pMRse8W78rHRS14CM8odrxI2Qf3APSN96WckcosMgFkwEv6kOpbpJ/+cx+Jp0g
9bM78I38/BXUdOmH+yNn1FLhG2hHB5rRNxPUAnzQ8OVj6PFFx3NqpbQBodCvG/FYuYQERG9KOGXH
N1hi5penVtmCTDUK3Ybt8fJNkqEtQf6C19GqeNerD4+ehmpy6w1ercmqjT38M6pe+C2+RYW3Gp57
BgQdI3UBsp55oyj3t5YtpIIpRvgWHKHmpPwAy21A4xxTbIfF9A8IVrYa+X8QQiKoXjA9odLXRhYW
WnCL34qGTbs2hNNE0X3NoUcvuI0ZX1qQA3pldkabwt3c2u1xV1b83ZPRLVeRzRkjrUsML2P8oZOp
sxGgpHyaCZQeaFkjb7OAnZAjM84RdhgD03bznA+vRCCyeHzMWW3O16MqixODvD0tPWAgyuG8C3f9
tQBoYm4QQXoaWdNJ3uLSVarYFa1I1M6GBoexsXFMdm1J5FIXmwxq1lRBL0W2hjtOA3k+YGwCNNGc
3aP5/CpYdAKqfnxneZpWMnEYwB4TmYve9+R3AHgtcdC2hM4DTm42OBoNpTYslo2B+APHfZvQgTX/
Ha7MNIUbhJ2Gc846PB22qAuFdCkGHiF9Oo+GheWZyKuknD4ntna0VWassjg8viwnMLgB8ba36Yjq
HI5qDh1fKxSkkB1D0s8iVo7P4CB9NJ0cpg+b2qrGw8jy/6POQ37ixC1OPzPCGLzkGMDDgh9rsCnj
CQzLvVwYcYMPZ9jITLM0aGge8UDpWdNlRwFSRAeihPlGrZVaiPK04K+uN36mt1fTfbXjGx2TeTgq
2t4ONliflmyrhoQPhWXyVU5vBXlcySs4JMsUzDFjnoZJ1NvzTki91v8uVbTATVdUcdnz7Utjyh/G
UIo5dZ+z4NqaCMEagULLZu6YIqEkB9ypMTCnGX1YWAb6NutNDxADMPxK+PAhNxX8PvkCqvTgVMMH
hBmHjj8ot7lYe7M7JBG9LfSNfJnRJqm8Itbhk7mX+a39casjMR3z/W6pCzJVRN9WRmDLIMQRx4/y
wSGkhp+GoU/FbofMJ40f+o1HlOQJURDJLq69u6sdGhJ9t5xRtQ8op5wzljBO1zvyUnLspNEy3yAy
ltiF6XMoNuYKnKqeZiBtlw9cvvqVkQyyHZFjfxUHljXW+3OnUA9Y34I1Z+Bm3dKBoKdCwBivxknk
Sese6xKF2r2CClaO7zKDEY36JJic47Wf2cA+rBinn2sXg805uIiAGU4xS5OgRUhLIPOuPY1AgrEi
+4P0FhpEb6zxHTWwNQ2ribtx1L1j5TTYMKpRgQTR0pYuBq6cYsSuuyhl2OLFd3XMZ0YAJxrOEwCg
wh9JFZTMpt4e7w95wOUq+ohl2/URWuDi873Aw20soJHL20oZIHLMLyfqiAJ7vITCRblXKqbCgoTp
0q4uld9gGX80qVkZgYTYV9uKgiPh6x2JxX8fAByUknFYG84kqD1n4Q9HI1c+7Oxksz0suK3nouVr
hBoHaq2b2X86L64PRY25S7RGyklbmhYbZFLW5jv08dryQB9RCg6vvFw2shz1O2FPJAx5l4rmjUEO
bVDTLJvbHutlnCY4YR/R22+02nGEURbxRKK+Qxi1Eif0Mlq02l42FUfp6/kabmwQMRtoIKFnYhwu
2vcRNhOZE+FQ+Aq115QR5gyEUAvhCkba/izX41YHc6/peUxNH9ofhTj7/tpOsXoIH76xxeLFlS4t
HaNdohLYUDp14ZcKOjdGTi67AJTUvaUxPs55M+Bt8uOV9u254K2kfp/wzZ22FDN2UvWMsTizV4uy
2lQNbPnjSmRA/NS8SrnCnFQ+aJ9jyCUwwdxWWp++Aaf1v+38KEbkqs8hXv+/TWy9pnFhkeQEhG19
CBTVBrYmNm64qzp/KBiIlW2Y7H9ImkhGpDRnwu1t/+MrnhhmdQcxpIcTKahbJkfpoTomFnksW4fv
lJW7E0FX4/lrT5VHc8Z86/gbW7HRGfPrq00+cSFwvVs0l2HlPAfJfUJZByTvaASL7LXCXKxdoHV/
BErkY8ocoCyJvPOnCOel8b/sZx74cyk6L2hLcOTYRp3v2U8Au0Wui63GsF/lbbxFs7bseHXgcKFH
R0acI07X/I5RcuuYwwzAyzS4sZ53K/cfJK+Payf9pe/onslkN/kLWXoMFei9d+wqDQAN67QUt+n+
VSb02fVe7cNiQiYS7xqxLzpOI8Shs4l866mKM9SHoNfEdO7B2uH5ahrgtLnG8fDexeFUkZfElPcH
cx+vIXtJ/HzAlvIEDcINdDfROJ8IwBBJ/iny8sXk1bJbKPF2OSuCWGKTXvIqLQAZA0pyMHLlho5T
lZtH83rin97KXmieNPTievefjJZd6BSkEBeB4hg0uXmIZCsnWC9y5WrhnIKFRDQwXeRk58++tvUm
5lMzpo/bVsECjsGMAuO9Jb1pkQ8tjHtiqGP5sDCoJWQK1Mn3xbE8H28wbCaMuBm1JiajdYX8mkUh
VzJKycDaAumlur6B0OAspyeFBWrA2HovoK834c4IK3WdFVX06xohuLJ2ZTCGNTMVzd3YRb9Ezfi2
geBiF2Wg7+iyNqa2QvngDrbH0WYLEAOTcbdzOvmAriFIiF1kRWgvQ7N8/Hjo0PqhlPczvCCr3I7f
wBvgtKzUPfV0JEycQ6afrvAww0DAIYpT2Ap/ov5HLYwqAbTOfosqcqOBtykITqVOfFRDk4bk2ndA
s7PzM5G+atGm1JicjhBs8h70jwXrpvgvKFg0YiNDmn78uWhGNL6pfJthvK+AvrhxITmEAp1sA4pu
6jeTr/WPogne8KDf3icZEtkXS8wN+mbni9GJyeYevRlquc79xs9s2sHmeUXqzJljuztj8XED4Trh
zII+bAv+YuXFB378ZRnqBjvOFwm8tVB/Fkpf3LpmvAu4lADplBvkrcZFS/njugPz4gjhY+VdbDI8
ffNXfYs103m8drWq7HSmtvhZH7Ly4sK4GwLK8fAZZJ08IY63nZ1mY8OsBcdDF5zuXfrJ2ndMYrKg
UJsORRi85VOPaEo40Vf8/Cx/JEHQpiBa6F7gdDnSopCi7vuNSyJkQO5t6/GqI67B99FVDTiISTZX
urEN80V9G2ipga2bPe7JuhhBUMJR79rr+B+vbffByUZR5PF0jX+BaSry2YKA9WJ2/JGNHqqeySD+
b8aoh61Weo4So8ppOazIku+A56oJGDZexHyoUoHDaHxwdwcrJm6rzXDcUvu01zxt0pmU1YXqOzs8
/3tu01muaqtC6l2D/U8hVVmeicxQ64fCE7HNtjkxF6ixaX+Kc5JCzUBDgxiwk/zLQ9DKh1dfHIur
17fBq1R2LOfMGCs0RizAICEsAketxowS4Kl+RHznw624EmjHk3uX5sTY/xcDd5ToExd/z/0i/P7b
Xm8Sj07kVWChBzke9lfeNept7hmYtGQelmI3nVCdvJh+VwtKioOkSl4qkwjDvEeQU2XKxWyA5ciF
x38/tHI7K5BdiqIY3G86aVobaI9eVcFG+EHzMAy/Wo4s2DmotctERfR8k+kanIKJcIor7b39MOI+
JFEq3Or3uLXKaO3xyRfVI2tfrlor9WGCHEewoLDCXb7erEb7xKeGMPbNnxcIvv9ltTgSSjGlrAaK
xMxLGd1vrKqffGHpJszNQDKDi1vb/KruoUvNdR4XVqVutXdD61RInIM9gOjT5Vemm1czLf86UFY3
73q5MBc+YM71R6FdqciJqVFuTDs6J62J+eUs8ALVJsTjIx4NyNQgCMbDfnjjSax1EYouEz2W0pmG
D6l31qwCeJBib67xpStRFxJnqNwVZ5ySZU+LmMVbJTkivu879LsKPG9io2mVqDhjp7rXfLMU9ZPJ
1/0gZhWLEjaGPhu2TXinPRRLTtFLV4wkSxvJuO6W9JOLFYDVLyjTPcAvzmFiE4RP/YQLOMdWm8K5
mCaiRrcJNLyQOcM7DVYqs9+/1N6MoPEjkHOHyZOsUvzu2S/JiIsOj2IVfdrJcWulEwetXmlemsR3
Xws+25dWR1bFHoFR6HThkl8R4zs9tr2AmwDYG8ctQ5620q4uaSHE677WzCtXik3F2xajmOPfrGzZ
1GdNnFs7/ckGxlLNDpLIaIQgHsZiNIeMbCDMkoeRNgahZH1WBwX+kEUepsIi7F4BVFecEJeLc4wU
IGB+VRogFyh/nnEbdTqTFKHnpg3AkqEdC9ulYO3zOKkY/IzFO4qNQCyJAOycsZDYL5fvhBHojhz2
NHwgN68ypefJRl3iRimUkhh6QDhIPTtocQEkbn6CwqXT5vdtQr15ChdUYkSLYwo8fJ4a9ddjQspF
WPf1Q1Ic1oh7v8ktC5SxCs/Sjzjj/RsN9vSROS+h/IYMPYJ+431RWc5sTEnEaFsD3sNViFL9e9by
Ys07InVOUuG/Sqj/gUHM78DyHkjYTmgEIJamK6OrhzAzjirteGbJWVSYsXFeRi76Ya8PfHEAO+l/
q/dwrorHRwa6B3MAAqJrRqdSYqRfB+li5aESXacaX4WanabFtWD1om8692tqCg9MKV4nEeCm6a34
h8zo+rAEHUQUwV7+9AwIf4fC196kFIHby7PpRqZefaEQR170U+OMi8mF8i0M3YWJMcmVFtqnQo2N
sDpxfOnZ+mYA4sYkK/427p7UYBIaRbIWT18EhXzsu59OWmKeU1DVXZHtNGFcv2MW/DnxzOWZAtOf
041aYFruXG17oXvbhrIi2xcWRVoUS4xjPL4GCJbnYYGPobxRT4GlzIJcCkIraioFVLQZS+tJumBc
u2JFWCmPdsqL9oS/7R8FXryiSkou6S/EQFQdq1crfeft8LCG82dcnNoR57gFIoBhl7TbAjJeTGf/
mqObPe+0+tIcDHcOwXbz9FgsGfgqROCsKFZG1x+4QeEQvASlRcIuH29x3/B4wmesZSUjTX8/Cill
1OwMm5s7cYHr/TDWCH6rLY6UWRURBn0LVz1MVcV3kg8GkKBjDVIvK0MQOatdTINJIkVFS3M04SdV
PmmL2kc1dxprQ2HFw/gQKHxDszD6u8mXX9ITeZQUXekHgqSlt0K2l6IFD0IBGeajDOP8OzUQPMTs
6hJWtPrHu+f8wQeYC+XYJmXlbRi31MtBF0zyBU/rsT4SSoopPg0ZwWgGz3w5EqvxZhLzG5+aN+iK
F8vWq+GemkAsMN8ljV5pUusnAPnJAbrxI0CPjajd7hPhquvux4jrVIa0VcBWyQZS3ETIyplQHxDc
hfT4mUvaDPJKwJUI3sJniS/YmQztcHYSUcGCbHrJOuuzh50ipZKB/KeNVNWqx+muy6qQTZn3+WBC
erlV1Md35hFQ0WLmUHWHBoAIYjBFb+g3IxmR+qJmSbkcU9qltXZ55dibDtYl9y1PoCCKJko3YnV3
V+vyQt0AhHyeZ8o1e5H8H1ICE9K2Pmj8d9ankQY0iUbj2jD+ZBkvmwN0nObwU7i7tEA5YRqc6YCv
90Xnl8I8V4KQWhLz1h1YKmUtT2GEpf4UznBhDes2E+osnz5WoTcMh1SgEc777yFa4LqRh0RP794+
6Ifv92RZa96bIZ9oRynkkewdXrqbMA4o88viGOZGWLHaifnvcPRieHg5oI7blCz0kOT6JQGKwofG
JFmHsU4xn6xeq/j7MMXox+7YItGTiigSQYblvXUQiQRY5PB0Zm16oTs1xaqZvs6W/LIja4vVbd7q
MfLRXw6Becu6x8aW2QwUviG9Hf7Tk/qz9Ea3Cn9rPigzcSrZDRUEw4cDH6ltp6hBZyOnQN9O2ebS
73pfoOQHJlI8mRb99BiA1se8tQp7cGlL2OU1N1Cwc39WBXsSIUvQIzvi3uETNO+zSCWhQFsWjyuu
Yrj+hYIINwoR1NCxvNN81uJQev3h9Ae4OSoiFfini+hrCeYQ2PAje0NpKGspaEDJp3+Rs/Sbn5a9
RA9gfuVhVJlGywI7BQ+duZ4l6Okqt51Hbf6Sbdk0rjiOMFZc8AVbcePLDFtdFIJgX7fOw+WDTJND
1H5MPHT6rKiOyyopiJhFPicIbwh+vzNrtdppDQPkO2MBXQfz++V2MemxwzziY4CmBq2B6Bkm/pTL
+iMAuoeCHdY2+1Srae4EQmDoM4MPxbGRMtAiz/c4j2ubKWwHHyim72jS5ZN+qnP/au/Z7bG3izdq
3yg3uBTymIDRQb8hsRQUwwDEX3dpNmGEkVrlebmFoSwIvnVbQ95xY3HAHqxWGG2MLLaLNkqNJmrG
OtnxAL1918EkR369fl/SQBIesEf+PPqXSOpabhJoHSoyA9Of5TUVsGEpfXYcpY9nk9KB27eitHh9
dzIXcOEFSnDruSs6WBsiq2GAENWybJYwzTkXf+5tiQsmFdy6NVEG3qqrvHM8MtdmOFmgXEGi0fJG
Bua/BkSWdGgcGJYnv/KCQEBBtxvWGcefiRhdjr0mPYpagmXtCxA/Zw1c8Z2pGZO3y8qsZad0TWj4
jOUb0J0JRyYxKLqxWx/OyrxecRcFJCphOttir83xRQlvXy9dnI6OSKixzY/kRlE4whloBmuW56M/
JDOMfzHnnNvt2zmDPs6Hsg+xqZj039XrCNYLP9UpoHXtHj0gU4YTHkSOK500qW7BSJWVZmD/pFkU
odLqsZR628KkNhKwBcaKpWVfPvYDM/1hZw1jjm//blvioTHfn9H8+EJKflwt2XmaYXdTkTFOEVnm
1q+8xnWFj3K89KXYr6nzMEXCV4jcgsLKwHmAGFrKmVsgcXtOexk8wA/+ZVH9lmKYaC0wkmXJiJ8v
c/Q7jzR0GleyoKxwwVgcBlIww+vHFUdYi/jLxg6DKIy3bK9jD+jJ547PTY5H2LEIwgp2patsxe9F
4yLCPWl7FilGG+x8WzTiykcEZ+atoVwddUzavnEL/wr6ppUjnYkaAYgbBIa09U5xVuuLrsQ9iBYA
1YrwUtWNLcIhgMpyzi4pGIZzeAL+MTMf2BU+3bAL2thV/mXFzno72e0q2T12ptYhqVZcHrzSg6Td
9E1bOAEbzmHwsLW1uEnOi30tA/IBJvNXBePXMYBeDXuxrOgEoZqEzrWat3iI1/WkIVnqevINe2PN
zptPZ6plRq9LLGYJaIVxJA7V1uFGzJM+BzQhhhGNtrXDxwZAnK3kAuts39T/91i7s0W0CmRgx22C
KtbEjHEBj60QSrGfSjdYOXnK+OK+8GCloxeBjOu8JydAc/EhfMwm1FndeqaXaZjaj+yijjfGwOVa
7/sJBfbCKPEnqKOKLYGE16cbUC8bfzdQyt/S/HmT1mWoz6f/mmCP5VUAcUD1O/VGKHD3da39qCL/
RX65o07fuB3FAYstm/bNIMsAeOssR9hFvL/HRaBV/eArrbrIaekONtdRRGS5xEF2ebhJVVG6DAoE
bl3ob5MhT5D21eI2l3F+G5bo6zXwu1vHVdbq57OaEbrkZBjT3/h+TdD87O9bE0YkiSnTrWmNkrTQ
8/0snQ/Ruqg7nFooy3k4LZNA9r9PsinEg1t+G4uKCPhnmUQqat1hZWYLluAmlwlAMMibA5w2jdOF
2lQSofhzaaAqngL57oHNjWnGN+fekjgN1sOJplvFc2TyffxnLL6nk45732rKV9dmTV6+xgUlohDC
QqXtacYgUjLov40rKGSmWnFJh/U+R5za5DUebiTNwTbqdiyjX2lqFA8Yd8/oIS0aTnbpGX+zhtRZ
31Gb+MFz1nwEbXbeVaRJjZc1V7WyKyqQWdOdmX7pApaXsJsnN5ePBJrFJPQ20EupBMF1e/klEwOx
o91ImlTpt3syGhqXCo8yGJgXzU3JvWACJov+gX8T5QelPqNBl2i38wn3SR3fU3UWc7eTgbXPCWES
YDTAsbMqlA2TlPTLMl2C9yN+xbyDtc02n33n6n9bTKzaowVigob51OtOn9YKZkuQyHWjq1NAydVj
Gc2ewsqZ0+4cfglPZ0nxPEmNH1uMYskW5bx7sQMzYMFvHiTQ1RwWUn11O+bWQfBq3J7/i44AMT9/
sXySLAhXAaabbDPWnA6iQFCYByKe/FiQNg3Ur4hQ7Vs+2clu035LRSTolkOpCUVdZuxC//CiCdQg
C/Y0sgBhhMJDNgKaxbTsnECCvpU8vLdMQijT95EWMl1bCLavUR/vXDGCnr4aT3hoQgrc8kVGBz8T
jHp2lk/oQ4jjhqlAsyb1KgluM+2o3E+zUr/F5BxPlj91NgkntP4y58EvuqBBrfpyV/i+3oy0pnB2
dEYgEFejtbP+9a+Xo2C7i62l13WNf1XuoRyPrrGV2xWI6Yl1/tIPqWzaWbvIALK//lUvOC7gCeh1
kEPEoBiojV3MGQPnkFFniTGdpNoaBWJuGet3kKAVIu332lc4JTXeRwk/mdy0TLKnka6u744DaGg+
+RLMqqu1+LFm3vaj6RLIysWWzfRkqAAeF81hqMBbmVuHZ73CEyQ7SuKSa8zIUHaK2k91+xkQRCjc
5fZFIxriEBYAjrpaK1qcwu1q9Xgymxf18gtEep6AB6HMRX35UlRxtWlP+TAqwBtb3nlTUGxPX2Lf
jdwJGPC5EIyTNj8BezrsgFAMA+cMWhAdLes4Oidm13LzX/hXFOmm1pLlK+Upsf+a2N1s1Pvwm0xV
QtBDQr7bY0hOGRVG4wa1eKVC4dxRID0KaCitCs0Dd3ykTe9MVfcj165cD+L1zUnCMnC/BFaokcrw
W9UyGp87gwN3L4hOUIMPu4UVo048eAYyaQ2zuRtjN0Vt1mylKcjJ8/bovZa4Jpp/MGA244fvuHZl
Dr2KKlIfJCWB4eHk+wUKi0PXQZdYPU6w4onB2ZBRhPdZ7x6GoLCNvw/J2L6t9Rmo/hqOYUCLOsaZ
RxaMYGo7ZwlCJX7IX6+vnsA0xd4H9VuLULcolFgGTcYfvqesbixWCnncDEtXs4SDtBUrIijKD9Ee
TnBgd5dwQ+FDA4F0nSV+mXKQH1c3z0yBUgjfw7wDQBSvgl/hVMiMFsIEEXUImjhRrWFwDoCnXdhv
BoMGsMD6pfGVk0lhI/Rz6j7xxdBrMT6czeaEgsVaOd+FJECdSe815LCf1Ldl6BOoO+OHi4fc1qnK
oUzNzgJqlbbxBsN9OCY5212P9H9E7sca/y65q36nm/VdaJ8PBVmaenJ3HkX7322qpGysTjCpQIco
SfM9Qy7mPmPENtIphWr0pVprzWsUFd7LJ7Vp61bn5iO9gvloSZrVkDG/SJocwol9UR2wWiyeJvej
k55MNJnKDc7DQAGnADDu+DxiKg63LvYkWDnSb29Jb5IpiNQ9qdMSmF5R/n4ywfF19whgMLJw4e4s
WhrLgmPKiNRkWwzJoczuNUmcH/H7X7iQMr9ogUW4IY2/BUb9/ZP3yW9RjUu6s+F06zN9JKZ0N5fX
kN3KRZb/pj45Y8b//uPWacD246ku/HYVZpmwytqbN2VCVHq086Y0cnMJmK5A3ARLuS0VVy+TA1nG
qgioIT4KElEpuSsreaE6I4iqFU6mNUyDZUJKnuHuT7XJ+IGPgfMox0caG/a/Cg117cu0zR+wXIOx
8NLGj0yMU8w12WinP/sLbDJvC/hduJZCbkUq9Ee8Kiz9wOZrMQlfk97KPXxkuoNyLgG/0qH/XGzm
mapGk4R7SCYbA6ICs4CbgBlKKNGi6QUb1fu/JepsFbokJyn5e2qCj/hOW0yTcmg88ob/WKl8VMS6
FFbHvKyrRc9tNSLp9dOaOaNdoKmBkESgILnbvlC0lyYPjNL5uPAnCsxXoen2X5Mkjdt2fgk2RNUN
s/b+jdd9rlUkF+rgNH96DvgifST2xQ67wtgymCnMHaYywQq43ZrgGfLYLQ2DTZYyew702PVgOGQ0
8DckWB5NhCgL0Y5uCGB2Pz1u/HpsqNbHhZFoY3HEcAm9ksiirFWEgknYOPCL0iovv70VwdAvnWnx
moa1lDabA9VVW0qkqUCIucQpQyPw4yQGW8F5u2Xw505fev+EtljJbVtbuOLmctVczp0C5FEVSd7Z
65jCrU5460ZKOgsTAUm17vmXF4K+GkvclTxT7kAlYwNFuceUgA11Ks6AM+JDIrHeVx94TApwTNAQ
CV2kmohtiSY9PTmWs49w8jXV3f2Nmr/q2HRWITeJP4H8Y8zPoRTE6jKAkxTxGWzIuk/v3EaBJTm9
bLHaiXR7VlMWEm3GN01cBiUowkV/saqe9oPIYbFXplI7ort+BycisWprorxJSNVcVPZITMRt9jt+
RyheBxQxhCNJPiEb/OMZA1QCXNFZnpSXgIpB/Bg3EgX4X1+Mhk/g7EZFp86jsboNNe8T66awY+Zx
pqLibPIvGoutCM7QMQOLM9cOyXMvYvLBHpczpOpErfRcMyNSVQS1DpmYnwkbf6YS5c3YQKzO9qgk
/QsCPA9HE4ZifyXYZ9f0KwP2wne1xSpivGldkCBb7V/+x3kx4xVbmEHlZ4CAhDNHMz1Ow6d0igDQ
ZO/f6nryVsHbWoGf8oewy/FxIfasF4m5roXK3Uljka6CBmbPxobZcSamO9gDpJGmRV7xJIOt/5IB
K/6/E9eDBIM6IiyTdlTXAMbXzrn+wH4dPlTCCLqwUbqyzmp7IRamfWDoyrx3xwnWfR53b0shdi1i
hLKhI6eo/d7bL3tBUml58+TtmffZBuuDqoWN9ZPHvdW2oVxgs0lMgrV1ucabxp6sir5dRfluzy8t
BfRZYR5QrM+55TcdONhpdd02v1xzXQw9TkgeOstI9ehqoxETeUbFxEolYmQalVuMDaQELjJOfCIo
5/tBjxdaUAFWPKaorZpBc+DlbB/swY7MYClilJPLwm0JLN0ga9wSWsuzQyQ7Nkqcl8s8rnWV2dza
IvSPB5uqVhEHD2Mi3T6yk5+U5xiiPg0N30Finxwx9u3/Q5oRUz6fPUw/Gf0TXlr80lZor960dmfc
ignzWeRCgaP7EUkh9yuheXdX0R20QMqQHb7ruuVQiBypCiHsT2M2PnHBjex/BJkcC7XLQQ7Lrhtb
xJxCnZW4fRSQsmwL+MQ4a+bXzmT4kS3FKhl3ifTj0NerLyAfg3suhia58uOI7qCXI4iG4GEvGWVS
cW2JUV94F8oGxXkeYqhjA7l5Bsekakt4HINifGVQew8ww68R9HY3KH/u6VpESAx7Vv8G/lkYu1Ee
oRXDlz7HHMJ6kT03a5dWEz2m4XCtGHeFKGUuH3AKXtS4LAQ1VhW2DYpkVpOmJO062o3rKrp28F1W
rc6sS1AuwZyVmFxdxEPqCQq7lb2sSAbVhbYHEVyzxU4JoFnANp6J4Thu2DXPRfauGDEYczOF/8fh
maR/xrdRgPwRcBJXmlEBZZjinoVYJDtS+92WF3i9f68kgf0w4yQeZ6umP/Vf1KQes25+ja6uQJuY
Mc/PygHMv58bw/3mIHrBsVVWm+Uyfq/doUbIdTY+RhMraR9q3gJtU7/NHrQGZ8Xc8Mz4+Zxn1yGj
F7J1ZsES2TkebZY0p98BsVtMHy6Uu13x8mBjpeMhft05rWtgIMtTCOPzO9A9D8GANqRBtXLF52ZH
3qM8CFiPA8ncExiMBq+Cl5xTwu8Gyj1jgCfODM2dVa6O1Hp8urZrDfxUYQL4ypHf/pW4ATsTx4b1
czAQUgIZ8l6gHC2CscF3dy58BlwIONP1XjhLIybg94U6H6BalRX+ISDS/aekrrjczV6KlYaMZ/6w
qaDpAtNtbnzyHhNDUWALDWyQX6YeoTTGjmo5dfeW32EwdUoMl9aZ/nkLGgn7ut1YfC5/0dELmvFg
ynMkX0kosfobdA9J/Iqywz74a6b3q1giDS8Ja6VL+yWYS6wJntTApqq4q6emyX+JbV2hoFoq7qWC
8hA+a3Y05eZUyAahlIb36qY9dx1cEEZQMkprw57IsB4IcHj/F6xIOB1mP09hYAd74P+37JQpsCLC
aahHoPdtWSN0GniKITwcxO1aLlK9rAzkx3cG7v+JwXXquVdcaw78ptoMETBQvmSU4lX1pTbMchv7
ktuAQ1NU9GNg4s6WVSPGWRyDhQjkKc9Z/1czIwKyDDEhiiyfD1q4Yy2wlwVNUxiGzP+LPd2U9WiA
MsP4ngZstNgr6iOVx4A+n+W6585R3qBwoW+g1ILKqvw5iXo9BOT/qToLArCHZE2w+KEXJDRF744i
38vWT7/fYU+jzr367hnwrYw4ECHJBQeApF23luBLPz9oM87Tl7kF/ZXXlBx2DiL+s7RsH6zB+Yg4
L06VA6zXBMNXDriOf5DPTadv0Oiz3N7bJyJ2vyKQ1XavMpbqtCK71o/cxWHoQUU+W2f0ywQFdAUD
Dc4+HP0Bs6ZVvQh1ptEjvwlQi4TAT6uHFxGl3kODMt+rDW5piJOBZgNWMKuYKQ88kMRjjlqtCB88
keudx7Qqz+svLv6BFTCPA2LWnYvqjYMxeKBcKSkhVm10MhyGqFeWwiOeO8ieRQACYsUWTXBJ0RNE
/48YOc/JyISSus9maBc+GcVBjleyGkijHz96qT3HYCu40QaJJlSwZw3XIkMQQiPdr2/AkruJ5OAZ
nhYA8pRvdyI9CCujTPuA73kWtWFsQx1dxK+WzKO4fAkcq6BBEpQ+Ngt1/7cF53+8gPuYscMK+nrw
0ST+M/fc5m8oOBRKqDM7NCchvsVK14I6Oxm9glWyrs0Uj9NPFBBaKu+biwqhSa1O6NBLUMyveoP/
ZzWdKpZW0SQ41cy27sX92IWvrEQjGEusjkSAA9E0B6XJW0LCJfFrUybAYwEWlNOv0ghWYUG5L/us
M2MEzbItpOQIg9m9/rOEq4uxZd2Tr7dgkH2P4VoVCrv2mrqGh9nG2Bz4/AhI7y5ajhLxiJJDcqTR
HXcKiZqi+CdBJjPId12OsEl4L4dszUUH5c0SnwjnMndy1GFM3FVmMhGKgMYQhFou30fuDpr9Ts35
RW1gvtrMkIjVUWuzrr5tuvQcG3B/T5eKjwm+lUe37vIuReZ4mNnAwz122XouNGU7X0Em0CVdQzYv
aPg5HwrStTZ7FIrjCihGUU6ojF9lNvwpPKzB1sIph+huoJvX6Ndep6fQppADjFfxGaKXoVVccyX9
NfCv1MpVe6D43n7rBuc0flwTUyctRerlgQXsOrLzeWzKTUw1gGtMs+DvTUGmv9gvtUOZtflPxOCH
+6R5+1a/hG7vlk3Wbcu60mK+k254WTaOww4YJ7qADU6wmoREECdh6Ixh1caHbavuDMQOu1+uZK9x
IEauZexmBAdeG/QQYRellMqjlVoHZ4fW00/As74M1ynwLkLj6uojcNI9SdUv/E796gS3NBvFdibb
EnrYJZJ3/gDrLUHAOO60PY9YitG+3JEv9gtFWM4O1X8Vl0NhJevlIsKc1VPZ7GbTxR5Xpq8HMFFW
VJ0hpUGCpEhMAGUBxsQIw9nBHW+hd7PGs+ZZgg7WtWM1002LS9EGWrQdrHoOC2slaurZB+yuNIsi
PCazqtexq2VJURUjlWI4UwrmJ0bq/Y+ekMBdNrxYXWS5YhydoNqp92whPr31AumNaVSdbFkocQPg
MNJs4LYzTLRp+xdbKGUfWHMfpMTEMIYcbAzlkEMEtttUixG+O3peDFjS85/j8/XqdNUzmyEB1dea
RaaTyGHDOR9rxTalN7+zoI99T0ylMEMG/nt3m/iHK0l1g54d1p4DVmnX8CdV/vjlGu/fXtAnli/8
UqrfDmsLwpM2DohmV66xlSfXictiH6eymD7Ylrd+feCgh3bNNM63zNhlXmosfuuJBw4qneJGueAH
D4tLUmouS84eqdHz8okidgOVZ+EqCJC08/Gz3G/N+zJT/kWLRp2XfsvswAE354NMejwDm8f+65iJ
B3bLzuQ1eZ50+3ryNCxjgoax0DZL5V6upIKuMx0NevaNohpTD6MG0Z0CIUpNGAsUuX/X5O3Du0js
53GgupSsz5j7x8hh18/wXVkrwcLzetfZcu2mpz1Ek/kwPBMAuPZ1hqpFBqPdiI5L8Gtt8eGVhsVj
Lfx1rRO7qpOekpWwSdPEOK62TN+VA3B/micCR6CY1Wxuwt1GAVd8pS+ir7GmwMNOGO/4V0narOI8
7wJzDIRx4jzeNJ0ezCucRZnjYCE5b4gcFDLusgld4QsGCqpA3YH3GqMsYEoe3HM2xDgZCgivAyKN
mgz7RFQem5sDAw+IwH8JPf3HWre4JL6QO7I2CApxUlkkoexnp/pKCSWpqaMb/gfBCG8BR03Tn0nI
3o9ILbWRmpmQOaQpAaW2LrmvbGNSPcrt9jovn2hka9Hx7QKVdJ4IuHoIO10rJCrdF2/p09aKAo/F
uqtDmG2rurGY0VQNBS5HxLxPln/0BJ8FenLL09+djt7vwKv/q0N2a9kVgvz41Xmwa29udMeEclj6
YiOewDEa8aeQ+qzYGStCoIdcQ8OxZw7e0E8z5moiZqAfZkzq0XRfXAYKE3GnQl+O5RLFPisoFjR7
W36dhKBuRejEQFTxKOY/NHuSbmmpTuleCwk+Zg0BMqTwGCMA5n4L831xiRJN7PCT4qFHryUD6ORP
u4OseTQj+Xs7736g0FqWsS+F533ozyOY+DyVt473za3tF9+FJH5g3tEz0BuTP5JfEGiZ1yIE80Og
0ak1hPsnfo7sWX6ny4BpPyZYoZ8skxIAYVwBujPHPt5J2ee/N1UiNvzqBLCTGo5OBhCMo9C8cWkd
WDfppSM/0vD3rXKQPD59U4ficmZ5KfI7OTh3cDhKhKGbBEt/AAIH07Ki+7oh5b80puAPqbNNZ1B8
JIJYKuJTrzcAYsbW2/0aj8ReN/i+S89jfA+2d9TjdlSAl1f57Gx+sN9bRINfoCtspDK96iiq2+mv
0SP9RqOL/JRb4Ylh6gjKOrYRhLdfM5jhJaKThu5oPPkp2DMDXvDko4JlTkhI+XZDV6YJs90krQ68
/3FSDOxK92DdwaJ0THRZ08hoikM3Zs3Foc81YxKmc9RoaOhz3DbVGNwmWvvFw8zFV5wc0pnNAjpR
gU/3rdwfngw65IaitMTfZF1JkL57uS7U3YaSlgI/AKSqHkbGdP8V416TQ1G+aCXwS3p+tAWBLXFW
THGH8GVbJdpBmyIH5s0EaMnZUYemOI4psolSQCoVNOWliTZpyI3xgJswCq3W7dWWQBi+QZNWW4P7
H884YuO8C55QAPeGGCGgwm18G1MXm+Osx3lk2dXSzmKsMp5YyyyvEyKeQHMrTl748elXrgQVdxf/
CCdIHdFk93YNQDDZObLEZtS1Wj88u3HC6obdf+e2WRF7POJBxjY+YJCMCqdBen5FwaSQRIThRlDd
4blRHi95VHIltNhZlAW0Wj8DNsYTpTQAXESgPuYBJPjhB4RWvH9A1BtEiIdq35eF3tFV+ZjxdGLA
Z21cWyv3XIotVP3kqFN8erTDc2FLt1rIUXcmyh2dhXsZz61BIvrUeaDvRGgPRJh1/wFFHQaUILL2
aepPrZqGEv/1cDqHVqZQ3I01mykXfRf6nzp6TzyohmKUCD7szi9NjNEcIiEwZOOeC2HBQdCMRzFf
0Xyi/uoJxH7VzrslrxFmbdp2h3Yqohii2KD1S7FtKvTWywsJcEcbKDjUzwQ83iepOa2YR6wFcb6c
hRIcEVPwIJxetn1mexjui8TCTKHk0nSrqoUqyoDOC9TNigk7m06XXYVuxo0GLwARdlp2anGv+uh2
Y64YUWPDsepOmfmMdaRpQwVR1GDuePZ2+VD0epW07S/elgXyZIuw62aG0zYPaSZ8PNppklOxO3Ke
KqGl6jEO2y3EYfhhdT59aRMWGBplFNJC6Sga00Sl4fu1g+yb/VZFKUge5VAIu2TlbyXB8FhmviUI
uOxY4M+3FXEOAiPeB2k6jsdPy09ogECrcQ660t27U5xPgA5KYh6mwZr7nYk+lyRL2bzPNYAph+bf
FKqcSjdVdaap1C7O5Hu/P5qg7Ezpl1lag2Q8SBmR3qq8X/5kF9BSTsZ1Lv21CW6x860iVq1wXLsU
LWu12/BWS0ybtJmo6+pNSecRWHXHxDM7mCi+SFK/yEvxafnz1ND/ZaI5ICkFCml0+lcYXmjy9atN
84zH6soqyFq6tjoTw5W6NObPAXRZ9nqx6cFp1Qdvfo6tWMDH1x2VIJZEJf53M5snNx7THHRSWpFn
8XwYbiJ6Sh0ThrNonbIa9369iEpNlsbJGhwi3lIzUdzN4ncqLGLonAtMWu4UGO7BUI3LQK+ODXgA
qG/NQzlCDXLGZrNqpNk+yxm6oY0pgHs5OXiHu7bh6a2XHIXuYZkRey/BxEDhK5nSKUfdhPVGcGyO
/EUl+D+eQJv6SMZG/qA/jKx6TwOUL82JEUk7O+lhufkIpbqwNuQwb3UjCGcoGmLFmeHttghlQV3C
cxERGeP8tQ/z4azpV5j8Kse20KoD0XtJNj8vUmC5AiO6dze3WyFHX/Kt6y2d/P+LcRmO1sHV3uqP
ZAhK3QCiQbu2ha2/Z4ok2btl4y5Wl8ORNcdijDJHVGEvEoavfKYhNB0hxaluyNh/WKv+YCi7ivkh
xhxZyuO0mZyDE2ogko1n4JfAB8h9X/R3EdMKgGxOxdDeY1EypMhTAVbyBNjEKmUCNvcqNPtTvAwC
2eucifpNrtSFH+O9pPNIA4WwevscyAbZ9EGP3v40EPci+UJalv+XAW1AbhTwPy8a9Gws4Nx/LUe/
ZJyj3AgY4PTQppdtylJ8cKYl6LTRR/p9VX3dyFbtddt4GTeAXAtcE/BT+BGjY54pmZR0w8pnl94J
sQMPKQQXk3WAIbllBbikOTrTHAEMTHvPy7SjtUNvdU+AHJoNT+xJxLIksIUqn+UNWSjOpHORFvVL
MVFKOHdm3q/zGUAuKyrQdfCDTpGeUSVAoPad6DoTbcbj9iHR+zbvteExBV6dfUwzJsB+XAyimoxB
bilMrsaQ1mNVx4rtzzOdk+gyGFfZBxPE84doy/AUDkDyBA401S1xCvhxatQgHvdcLCySyjaj3mOO
Bu8SuwlbQtWts6dDr7kC8BnK7fFFhySCGIqaPXp3/RkOgDNLx/jz52llIKUiKD/Cihxhj5izw9Wm
S8eADnq04ZQ80ZewgIj031cXS8+udyaY5O4V/+WALqenPOTP7TmQNLE6FidGmoxwakWS8Ud/IO4I
pMf5xncygOb6kTRPboy+O1RuZFo5X6sXBO4oFdWFFt3zLwckZRdemOQOezTaphMqk2aBRBzWecvr
oKa6IeQ7z0SjdAjn1e08M+FRid78BZRcW8Upj9VbCldXRbcAsaOZ7hG3NWx2ZP6yP8E7Xe8DqHr8
Vh+u70BqjOEYj0v9ZPMJ0PomanFftsAv26fDRAQgU7HS3nbcsBC8LtcgZQcMkOqAdta1/2p6Kmne
BjNgssDJfywBEN/PXfG4JxRk9mzqDC6PQLygDT2mwpHSV2/oP9lLo5dC2tqfF2wStR2dTylsoNd1
7R8YTf+Pt5di1UKkoNqj2RdfEGJKJOvNDBHJ7Il4Y7+G45euejdReEvZqcBTZzXhr8lYSqYYOs1M
6lSHWVNeE+YKw2Zea62pKSDip9zUOndqNHQRtml/1zUvd24/LUX7DQB0cH8orTRRz4VYV1i9SoDE
bgU2qLK25IAq74r+xAi69w5LoSqxtPvw0vS4thHgNcH1QX76HcXkc+iy6OGpeuiT4X42uriueUC6
m9/qGchgkWEA4uIgwJq1MtpWeNbSHR5n5vfPYfe+4Pg3G3s404nLkRnTraiyFjDiQxOHKQz1nz2r
3nPhZkzfdW4pjue3GEB1zpXvctcBlGwEMO6fPQnlLJXVpYPIW4nWGF7KsQZVmPxFLUGnavsnJWgP
tVISbKnSMznctQNpP2Yjmvf6U0LPF9V43lW0ffCNhDi5CCUvj4Ji8vdbknUQaeKJ7ioxz+HZkLKX
JfSB9EsslmtwFvw/I/U2ODmt+xxvNtBAIvAdRwNuNHDM+26/LE4gSDd8ayVAK+eyNo/mfBppw92e
vruC5ASrpOZ2vFtxGbVXEjAWZIsDN4pt4jwSuudTK7cyRuwD3kXcDslNCgatB43+aRrqWfg6BwYq
/jhtg2snr3JFRIg0RTyE12fOJY9mFVPlgsGWN0XF6nm2jt04CKPgCGM2qhqb1/p48q1Bj33iw+kH
JKBwb9VSwvSbBgt90Ymp46r8WKId2S3SJj4KnXHLjoyer0irkCouVKZjLhEYUkTT7L6FwFtgF2+6
AXUb9gGQX3nxnexXTsC6KF4hw/HOp/RwI9g+GEfIS7dqbR3NYjVgJ5k9o1sWueupi68uvmNmNAgS
cSVsab6xcqXPIn6rXFBrcSKvbNqrEl2T+hFYkhmYDYjeeLfVLC4lem8yuF8IabsGhxnuF0odzb21
Nxd8aS0IOqZNw6ZSdwNjmeyCje/JbWiixgL0HyS0iK48xt6Q6dfOB9OrITn2JenG8un14dHHJABn
WE5RFEF9gS9CQysrjDDLZMBX3eFIRgWL6Z/0Ei3YV2v/x/4S0xFMZ5AOV8ALzIgsGV+a2SOQYLT3
F+GvhiIWnmvK/krrpjWsYRfsYjzkm65XauZ3ps09aGR2KHyV2s5EZTCkDY53mfngdTdeP1VRHtIY
/HschGUBGSlsVmNXr5O7x/62CZxWNzH22naxGfQB2oOn7DyYZPlC/J1ckNiH04RKp4o4tIEGi6Mp
90bkrpF0KKXqVaiX6zlMpU15L8KI5PrHVI2cNWXNUrP4NFsD9qvgID57Wo0jZCGEb/wOR1N2BSxS
0viT/a8v4rFhc85JjuYCE7+pTezJn3xjaqLW6/Gy+IBSQqe5AZXJlI8pzlxmhkC1p+FEhKzdnmaY
YCJeUwR6v/TH5sApxywmAxG20t24OUT3AVJjLuomc/L7EC9X3Jy2FcCRrsJOr4XXgymFWwYeDJmG
9bJcRz2a7/qNV5R3A0iYAaCeTnTHygzQG571Z2VqrCub7NJFAidSYwgiawlB5WkVYR6MQZdiS+wt
u3nnJ2ie5VPQS1JB7dDSEDeLcHlGZu4WuYKBf13pS2IHJjE0NJLcy7VJ3p85gcKTwm7+lzOhEkJI
CnW5jVlV/bBiLApzQRL8BVEtB4Ohwf6/Pz7PB7Ze7vlALOC8uLebVY0y8g7YVpZ1L00qtikCPDNT
lTcqmIPY3KwlGsTg0VfO2+UusqrvdqZbOthFuBxuXaHq30NAso55kXtTEMJqz3vQrZhqBfqoW/Vn
r90Vjkj90kuU3D7yvgjy4nebr8Z5sDDZ14KRchIodCU2wx0S4tnGb8Fac4goPM8fQQoCgtUlBy+q
0Liq9dDJB+kW/l5kRT4TQ3/rfrgUyb4PoBxc0s+F+YNX5alr0Tm47yi3KPB7wqmTcaSnguzhrcSD
jKgLITOopzsHbS6tBrD9xPgDivTS+EwsZGOU9ZVash6nqQIIKq3K+9VhZctmbfhzaqThloUywCOj
85sERvGmZVGx2h4+nL5IMNA6g1biKNNgyHCzBr1KMZiDOJ6TX3YjTx5h6uQWAXkXdkObRXQwLHXA
OryPYro2zYrhI5Dku/zQHJ0Vo2vZw6H+Ghd6fzJjMn+BvavcTr6YZWsrehWCJGIE32NWoB93CYXr
BQEqt7/PgbfN8t9ykA/UXFzKCUkURtymFglfph5KIxBU1tka5O76wPN52y1fXEyjz23IDC5Un0cL
Ue96cUVWqGVBZwNAL9QhEJV5rjK+arizLqReBRN3hOjFZ6RY8C7ncS4hZRmlab1uoYp5gRnkVube
eC8PE/xMSfI7kGTmpoI//QD0RAoVnGvxB5TYCyFg+++c3bGF6pvhznrLS/hCdDBBweJjrl2lkgEY
V87uQrrdD80bX03EMcsD8b4tjOfHUE5R16zOWE2p1zyvkZ/T/uymizRXvVqUwLT9E3UuWMf/YLE0
ZXKJeZc37GchbKoL+1HKP1062JYqBhWpy+BEWZKUzc8Z67DKLQi/uywYLXBFUnpLndX9FREAZoTy
EU8igzq3Vi/o0OF7rm9engRD/VSjMCI7fsnF/yPAsRvXRGtY3LxhqkNzLWgw5u8+s0gUiAg8KX9d
HIV5uJNsLzTsOpswtk2ApOfy0xgl/BpcDlQ5pVBy3hHhC/G2f/qizUruuoJa57KxInEi3rrByRYn
zbkh6Wf3DDc/qkkQ1/wal66m+S/l1wgySd84UA/sLPhradHHAhetuMicaFA/AkqYbiFa8G03/nDV
cbx+F2unq/R74Unytguu7X33Q4KLSZNkzzw5B6N6HFT10nRJAO7xYT1k2XSmDH/XWeiTYJkFH0GR
B0ly1hbXNVOi+bQezo6dvQCzLjFKOb0SuAHCvDBaS8NXAhrbaWGQDq7lU3Y/s/OXugz5xzik/fIo
ns6+JqNWHMZG1dv9i6/0UIb/9K9OY1vfBbL96T0nIftOxbkM2GtwDq/au32zU6TvYwT/pMBRYkiz
oiya6HnvpFJdfim13BqRQVm3bTLtZMsoikiGtXL+wuq3iINDNTIc7BM3vpQLq4Z1ckQzG1kN6oGW
J6xBJdTxVlDF9LJkDLVSrjedVLRmgCYPnArZYYkmaYsu0EYggADsJj5tCTH0gfVhy9vT3DA7ITbL
Iw/1UnebArD9FPwNr3xntSEpomDTBnpjrYg9Mx65/x5IIF7bwktWkG7iiKY4NVaM7TZbBSD0kVwh
l969hJpjzxlX8w6ubd2rEMCfGVrodYEBD/eJQzOsIwzBOIrm8DGfTPdYLhavJNkpU1hthZ/XRBip
xOkHAgtcGUZH+CqGloAhB+mOjx4zMy488pajtfjoTkZM4wA9rFfpTjHoToD5U5dpxSmdQAIXD0r2
EKezJ6ECJIDTTdQQfRylGAuEYIMsp0f/z8doUjKIRJ+mgRncrnKqXEezbAS/MImGjB7z/zj7ZC8C
pzo4+dR1Rrj5lzyPzLXdAm8GZ2sLK8uVjPnMXb/AUqVyk8xciw3Btj5Gh0SOWFB+Hs+AYk5WRREf
MkdSQTozIi56zuXDpPynC0VqmOFCZgpRS22wwobzrmfm6KPKMdle4kLwrw01sNTY16lsEk33kzs0
voFoyShYffE/MQ1DnLxtm8hhHDuk+k9nYIItL6Tg7/+ls1X9j87pu/P2EPqatdg4lFKNGTizgo5s
o9qQH/0yHFPJ20AUsprfmgmLETU3BQ/NFjhyl5msKof6Gu2wuPnpfnIvb3NWmdczX48lZ9KZkAHB
+h47ffkuGaIYveZI1sdkGhbjkBOsZg4R3FC4kOs13ItagTjqUw0aeDeVHJaHmHB4nhGxpvyAobnA
hLe5G4Nbx0pGM6VmSebaU+CSXHBtZm+n1DKcyQ/g+YuJzq7bUOLPq0hw4e3N7xuaE8LurM1Wls/o
moOKy34PisjeqvQyQkVrpiQP4Twidbum/onFlO6kHGuyWoaKFDpUH6Bd4SYDvmGvwmJIeelhzAjV
nRQr/iG70c74FSqj9as2CFJuwdgHaCkR9FSgPFdlkqrXi3P/jZIiDa+sKscXRJXpEXNTOQ2nG7cu
dGp1jNbLnfnXJDJpgOlE5SoAbq09H8HocszY40IGYTwy0UoCpNziAdSctOmXlIBj0c/kNQWsyocq
SrVos8cEWD03nDFJ8BnC+49xHlIgEcDMax5kzCGp6r6OeGXnhRopWvjIew5Tnt/qk6w2A/+KfTjO
VuUr4GtGjGW9gwvudVXaTlKB59ASQ0qGopjQjKpW2PZfvo2p3uIFVgjWSmsT2vXIUumih5YTXZka
gT0NZY/dlnarBJQsB+X6+hx4hN/+NOPlpsFMqY9OBOX74zlz8f9VEqkZo82LBahlCotfbOU+Gnbw
ww9BBWyli8Af/pbafV6MX1K8XHPYAG8Xjia9LBn9de7410wqUddPe5lCTOBh1AKCZwjQc3tZ3PzC
XDJBk8rAVMq5Asfou+b1ZtIBltVnULGsRv/ZlT4GUONnlNj8uRGCbTNKMdCoUi+ZI5JpVrnCNtyO
Xvhmgsz8U7pcQlJbkeYYTHrXn5U3BUfJqGHhTH9RISyVr5PE5aA43CiuO2aByzCawP+clxMe8R/H
iqUXHJ9tGB/oYZxElokyItyLS207HcSUkKYAB/FS6hs+SEXYd67QE8Gk//rtrQXbq5BS+TnIoWRH
5KlIgEr/yS/syS+oJZq5T5hT9cffOoSmmAfHujfboO0qUMupBiobqtG2H2cp4NlfOstKZ4tKjWVO
nU4Yw5KpoGnjMcv2WG79HQFlKdawupxqVn/+54hCtvxMbFftpeB4wbez6DSUs8uEsDswhWjJ2PJ9
rTjGEIIUu9hZT31IsUIRAuHmSsPGp1sPCNYksowEYUuWTx5dVx/IbcpGXnGtpgkg9WjdbUG+W9RZ
GXup+r/4qTi8Kd7cd0kS984tx+WrKoAFxaiqGw/4cSkA4Pm8xEqrYCc7lZ1EK2+K1/FHjC8IsQqs
Xg8JQ8zcTOhuILut4yXMeDFHPbJopJUjat2VhIFX33eUDpsQNn2Nssw21x8B9J+eSBSvqVHMiiLl
smt3H4qZHVxNvCDY3tRcubzVe8FBkUtKYowEfHQS2hkOD97eEQoy7q3lmVkdv4boSHrh3wzX2oil
BvDnIr/tQT33RCQE+98R92If5jdJpz+97VEH5hnMnRZQJYrvToe6PJ6hadArCtH2y+WTTwkg6pRZ
FNTWqBoerB259WeHR5pO5nvkHi4VwHCxPN7YYv+JYm4p2zcLKYnkYA0BGVV6tZdvLV0dgXm/1vpa
KfWbwubmv5KZIa12Qx7by30t/qzdc5nKy+D+jtMzkVDl/tYqk+YZvliUJpQDILKaQvZ6cTQg3ddf
ETp9tgAR/6RnAdeuW2melUYR87XS48BaP/JgDbizY/jIfCW0DxfsER0EQlqXEMtc2aktwfzm3wdw
4D5fMZ8L+aB1D0RLzLinSDbk3FUDfybBmfY41pchGKhSC4GgBVGP0kiaHFGSSXN4jBov+cQnSUku
SL+RmM/PiPDnoFG/1ujk4o7g6KRKZrWrYJHNOv/VKvBgFbeS9A4nlW+vMQ1mDap5bVME61pC1F4/
qLuyDF4kLkA47Ks3FOed4rvIAFHA0yAAp6FWpsVz0Tj+gRla+h1Na3A+6qZiZdqpmLJ6/ovSmJxw
J5AM/KthIPO6R+cUJUcFea/fBcXElzDpITo2h8DEX1mFsLM7FRruTEpDbR6RoO2ZU/RHSKVyZ/hA
c4+3zC0rMaG3YUDIDP2WxN2qHGVmEp8t13nq1HuWfsVy7iIp19kO9Dgn/ZuJ4wWCoaHTNR7zUsfh
vnwmTJPvKSK2Ml2q3ZoiN7c6sEi+KupYmywgawdaeR0M5X9oeADP/d4FtQ4X5GV6QrRZWk+vMRqJ
l2Fteq2ceaQ7vaDEHPWN33m0lAYcD21XifEypzKQUD7LDB9f3l3IOlXBENPvLpZkMWl681p8kdV4
7wnCizikuxlCKHJs1d0wGLzLDyeHzFTNN+NUjq2gkjfD1yJ6+HOtUatdJlGd9wIHqpCYIiFyHqJl
NDvBQF18JzwDeA0h5VXnFoD96uLHix07e7rbmjvD0tDdePo1V262q8Li2vxOnDJc77xlwo/jW9lc
uXG6XnI8aOKLYCUcbp7+qWUBGVJkPLlGW+0hNqeS/lJqZ2t19r1mnV6sONJYG5/e2D9VQFo2TTjn
yqzG0VY7C1WnibZ4Lc0cxl2Zg+LnkEHTAYjPiAiNbM7D+LTz6fR7g40PIi2WYjQvh4ep/YsFquvd
pT0zHvn3eCcYF5Kdh2YItdremhmvBeUSpEYN61x5P+MmXZGpT5EXPxg78OBSifN2OhCAmqdBuseB
LN6zaHjlGNV5sTgGSxuQfJEjYilhPaBlmCu/bP/Pla7zXa4veTLJPVdrobYkH6LfrqgDsBStzrQf
IS1RSV6f7KCr9BWMvyAELe4bGPXwcqGkk1Dd1/Aa5T3nb4lM9aov6t2GAge3B/p7F0IJPMhjeoGP
iFW6RX7sSi2z8G8IYCph9JwDOeF3Goliyu4hV0NAESrszpweSf5p3y3IjOPNKdJLYm+X8m4XYhcJ
AVFGoLjl7WvUxjjNZq8jHahhkvLVmVB2fVSO1oGiXud+6u9XqGo3fLTgcMXm7ffVfZCo1xBzhQti
PEtwdyjxEbtQwmvrbVeV7iCE3CMwnApzYB09wmkF5gIrNfLcV1uc2WDPBRdhFDh413YJdv26EkK3
NAz9XH5LVNZ9P8WOP9Xn+yQuJmi5SJwUYByUuz7k48+YBNNUDhD1p52kmLVZMBMSaqIU/XfnFZGP
+4VVssCojlzna+qPYQbG8283NtazRO6Ka7DJrU0U131pTgMcle5fUJrIPSmlqPzzgRZUjXMUnIJI
TFKqfjrqRxr0IaUGLKcbR0Z2yR0smndC9YJ3h7oCyneUH+H/qK4Gixpkq9pMi4J6ojfA9kFRhGuU
Oz6qTQGsVY6kCuZ0ZjJU43Dm/nenEnpmf/dEwlqLRABlSRaxu40LwjZeBcIARHHcSA1UtByJzm56
S4MyINPp3XmIQh9yyG6wnnYaYXk3ULLV1q76Zn44Qsiv+i462qc08QkU4l3Akm/32ywznTTgCRSp
NO01kkNab2qYkYLqXWkz/N6sj1bdEXEMc8l7tgup9+SNnyrbZ10lWMpYLul/JLDrIWXsRUD2VqKT
aZv+Mngnl4dp+6pWnvHiqfeilRXY/eBIQchCrM4wV5nZADxrdC4yl/KIswMswLMIfLCS2NEnhFbG
yvucjkUPoXJBn0uQxDUimjXI4lS8tyGs1v11GG0D8bCoDeejQ5G5oX4T2nDviBCy/MZkagM7g1tZ
/B2tc+rf1wI29/4CMF7mmvrG2TqqWrhscr6Mk50kapc0+Ed6r6gQcNPoC/rQ267RteAmvgde78Ol
WEQcN210hBQmH48ZlQswHARnkd4L3J1QcL2vwgdGxku6eg64tZKhWOcqlVFTi/B09NYK890ac0Ii
MerSUbC7XqvVQ5MTBWnqCwMAkuBjMoKwY0RBISMHX7L3mf03nQ5bNReSLLmWnixUGteTsmWuqsGS
v5aFCP7w4u/Z+bUbpca3O8yRvbBUWDCQk1BxRU+OKc8IR8aPiCxRm3z3E0Ac02Yj7WyOZ9VSahSW
wuAR/Q0rEbDduRyPX4J/nLmMSCty+Ijg5Pj2BTGbx4y/rvvx4+NSYjkWQPR4ODcznyHcdch1AU+c
vqjdo5tz0FzevNksHeHTiXYInZAGJfFJ1QYTWB3d6rjUveq4LnrXKuwaZGRSN3CzAW4j03b5eNdI
J+yafTvrHZZE3f8edHo+Jgu6AANz/CYFUcCqeDNHXbDT4KWToTWdRCQal0JyRwvBGp44scS9iR6Z
MsXIEPgS1mSyOzuFVGJUBCfHYE0B+8L8etIPYP/MOJETHZkR03tOJd83GRbbmpvTnp3UmeI3dUhe
+vuZotP4WQpxUrdLGNCuLuHMVsQjA6y/frS51bFnQk+EGJRIJo/vvl2ec5RghBTiF1RLCnpxwl0F
z0XmpZ0I1kfOIbkGm3HQCMvkTkYvfzKkW4phtUqNCZF7d+ROrhccjaAcCKfp3qYhq2ma4D66uV2e
yzNEpGw0sNc7/HXpozWVVfqWZ6pqeL3oYRYqGjffE6wMcYLsuiQpkkQSA/NN+muOHcxwfIGkvS33
fCdi56+i7nwkPQz/4uiHE017JPMbj42ByJY3lTbSVCCxcz7ngYV+/FC2ypc+Wb0+xxc0jMbEWj1x
35XAkPMGNkfIqb4M38I0ok5h8arqK5DCI6IsZLF5lalffB9A47gEFxgJAKaC6JgiwWo1b4XW6hcv
U/T6QrZ0Gdzk2Du3UIKZDYpmM+iaDRnWd2AAeIis/CPGdyCmXe1n6JbyFqgHFHonE42kNc2gSkXe
ksTlZuFuLd0NIv+Xc/MvcAfkRFTskq0lWbSIdtngjrd7TIcEZqQHLqdV5/a41cYr7cWmZZssQa7i
/IJ6eaXUPxS93g7J2eosrWzzx9VNg1Bjy+DpWf/ws9UvpPu+Cwu6UuQv3LqP1JUEXZROJwCTms2z
eOJZfVztCUOJNZ5ZqMKbnAixqlXJ8gKvrcbdqMdbFXhS30Boj88OL2kf8QpYvNNXY2bXNlbD5Gbm
Zdgtw5ir8qp1zqWtwNlEjWQTgayGA6kPRgmmLi/YtJQK6j48LFOKa4RSSvNDeUBtOEMQk6wVc8uD
KuEAAR97Fq0FXDziNb5EgCmsthqra2vs0CV9QBSF0BaQJPPY6ETqFzhpxvnD3yDASWw/946h+68G
Ty8aRVSyWh60WwFgBqtmsPKe0C1Mg4jgBZ672DYgTDzxx74JW00cNL4tJaM+7QVvMJaJTNV+Ptrz
nduperdJqspeGYdqKb2MwqCk8lnoTyai5lj+C9gimvra6uVOllP+muIFCVwMVjKXOaW7hfZho7GN
kybkHAB56RzrTOZX6p0UJ/Cf3fbmX1DRuj73sX7/Ij2IAHQ/nr0eL/efEGdIicFZgfEQS6deISPb
sB/aQVK6kyQZzDknncDrLEyPEjLk8f8rmB5SfIIpkIZJ+AT1KHkO2S+KP1pRdmz4ELARWSkCjdP5
+WZkOgcKh1zN2DQiYe2htfMcq7F50fHj/RB83gnBsZznu46Je4H4D6Z7pSDSF0Ujp59FmuK0tVqf
brTJ1BvtZZLtnHwk7AGjD+PoENwoaZFK5xowRE8BArNtFsEOdenxmNmJ8bCKq9ju4z58gyJXuhrE
PUohW5+FUBJoCfR0lN11h64Wbsozw/8Qh30QntyZEheX9klwqotJ2eDjgfmR2yfpoBOyMwD3JAvK
r6atIiWNv9OPSfAp+rAS4UZyRY4mvziehjS4TgmtFjVGZi6Nheou0ePHlxAauTZ7Osy4LUTYn8Bm
zpbodHxhkIvonxO2auQRXOt35uewZcfbDdCqajUun20hfsLnpL9NZafQYVyydOvZz+TYH6yW9mB1
m2eGTKj709cqlV4tNsV/iDBbAOhNd7pLm6hNKRyXOemeSDSkakLPDXQuEs29ipTMRzWuDTS3mdVC
w1OpPqIsH2B2V2iejIZ/e70K9Py84QdOgiWWh4wo4AF0LI/xME7xKEu83Q2meAP6R8zreSuxUuo4
/52rlaMp2K59WuslQ6DG9Dmss2znfS415HmhTaLTk+psQxXju0s2PB2A7Ha7UJQ2gb5WbMaGKBgs
7KUaJhwGz/HGUQTZlMqDZe84aaUHa0Q3jK73QGiMQPqn3lCCqlc+bHahzyYrHnvfqeppvnXxwnNc
UMsC2149fau/iSmPEuq+IaHUlJxkJdqp+++T/uy+PU02MRE3dK/LrGecYTIVyhfJGsSYAElOZWuw
qJRA58uDfbvKrbD+BcUmjV3Awwe5dkh3qnS40dpTXFuT1b5yevUwY7cHl8wbxDfPeQwb7Jk3hz0P
05GjbZo6AV0gaJn+3wk38iJVdE+r03RIU0mvMrhctlXlICZWlelZlowiNkU03v/PMji4JWczhkxF
JPt2Z5k9qcfjf/EGn+ev9U8UCfJfwJJ6Da/UdI184C1ZIxnndFDySkXG1ZTYrkHq5KRegK5y5B0u
m72j1k0GFPEDUSrJYArb9ulcNc1MYHWwS8UtwRnKJ4xhWVIV9UlcE/t3xYlfq8KRoWjZXJX4+vei
n4h/QazQjxTPR/Xrv902DpXWl8b3MbgX7N2JYZ4+PatVdiVA5he0pJ5FlT4+T84PrNWoecWuH+b3
hXuLByySxwqPnSWMaEhJKDVl3OAL2zKhr9oXVPYPUuJ93AOs/Oc4bs0G1PlJ+bwhAv9xlaFUoN8A
v4SrPfn9qbJiOvbi9iTPPRaldEBi6tOV7SAU93WyjmdLl7E71uXefUPfjyBd8NMUiXK9pvYLTGpn
5x4aLlQhf+OAmxBMcs89FXEPcuM6iQq4gA89TqhYRZ/gBjc0nPACYZ6Z8OgyBzkMcykcX0r10t+s
eZJyT712j3nJTaO3c19yDd5K3bsn2rOvSrTEgM4VeckNcPYaM+Mo7rxOfQ4auzBD1OK67oOtW/Pt
gmjduvSam6fu2OxKt3p9KfO4F28qOKqhAru9XF3bxWbRevcev9VTQ8d13KKgeOX444KplMRW/EQr
NLBGY5XBM/waWXsQ76ValP/CHD1CakERpyc+XHDP7y1JpfkKGx40lyvb0zQA7uu9DHIQeIMZ8CQV
86t06jpGFBRxBYlosllmECcgi54VTmuDu9e9By+dDrUiuMCv/xW/s8cYlfOVpKjTg9Y+dZOuAuvk
sbvRH2sOyg3g8ubl9OqZLZ89JyRpKjIttY1bv4cg/oF63Fv53Om9/aXr3AEhFpP+PvV1T/tj6i+h
jT01QYybd0gq9ZVp9qFtVhRIZpYmA1Ca4q3X3UBOCoYsemW25ejY3qNsBNbD3V9fGBWju+UTnJeL
KYs+r/Q4qgIyqL5YuZNoqlGef8PJ8qh0XoXUSuEzMowKPfiJhJ2iaKCwbWvAHVCdGZvmvjOn5WWc
EzhgiTpGtKgRq2K2p7bbbzfXh+Uf5OZAsHG0eU9crDYoEURmrHJ2g2B8fgiBhD89xnnv+uxbPrW7
Bs+kUWkdiY6NO9gKEKSUnlzzeKNgAIVy79OVNOcFZuujotIj20xKdLI8Zj+ui8JBwo6gwwyAb5VV
lfA72tbKhg6t5S79NtswzCHUR0dguz5U60t+jJnnNmLQT4bIPAy/RHhouzf/ZP0WIgfVeomK2HDO
8isf1C/A3d/yo0tKKFQMe8j+7XaINOnVYZaUyitO3soGa3G0jPkQ1mPXcBvPV3s+SxDFu8eBNIKJ
DpEK29JOcgS7xz0BDhAiOQ4sed66c+s+t9/ofD52g2Slnn040blEq3XEDaAnaJm5vQXYMGD7mlZ6
zVKWtAQOhyxE27UHM5xXbQKq9ts3D75ag8+ttEcybDlEgO5D89Sb3M9Y7qUvcZRZ3Sb+CcKq0MLO
dmcWDldLJbyfsHjVXVj0EW7ibRJOeEeNQRakNZCtWcxYU+8slmCXwB4+ZUJNI2KzFE6BUI8ar3bt
KSsnXu4HFZRhaqpWXfpILLNtP9Mzmsn62X20q4uOZgYgDNmseSNpfN6ysBoCeJJFzN60+OPo1dnR
JFSMVeuFCjct6pWfgn6vuDhT2YgJKbwg76jATZftLyqrvQqrZiq9BF6D0pTbv0tFM3SmsqUb5z+G
S5jJmRQJQaXjuBgcUiCsMxSyTip+JtIS94P96XnnGOW0b8jw595a7vxATcRzFYoTvuKznvMLINbx
HOaPua+Akl9RPW8Z3FqoYbFjLHfHjMjqP2VQScF75ZCI1Gjx0SRZw50Jm1+s+mvfRGb1sETqUQrf
sEmUp9qJXSJPkE8UL8936XveAeYleo7vczYw3jrIVW/x2ZTRt8O6M4V9nBx2z2DuyoGh1PJTn32J
Gu5mbKt9G1zGGj/gg21CzVO1AYDqIKmasIp05n1n1VB4/FsooT5Lcapkk/9qiuYO5CCYuc+/Krwx
jBrGnlELpk201lUKuYrko+PEjbKQy8A+jUOkEOgSdyP/s5iO2Qrppg02obsZqGX7w2R3sxNe579f
VEz4IzyLXB/TydmAMfMaZEmsFLU+OaCTm6McZuF0A3yjzD5h5cFHA/2+YdINE8HddHT+gyORf5pc
q4JichOFeNg4htdl/xeo3HllIxUu6QNOgglHp9Y6UDaIYQWmiM3UPweECihXFXyUHuG65W52HOTF
DynpP3lmrDul4rnKiy5Odga/zWWvo9GPItb8PWIHM9DHdsbWBEJGiBRjWghpACnhK25cmZkc0GVg
l8vj1n62uwm6eJ4zj0jqs357QhD4xsdF86LH/DFlRYW4DGlSh3duYRPLwBr4efo5vkwlbBsxnRuU
tj6Ndim2u4m97aBOh1OpQUEY4oP5F18jnAHu1LL9XTpw81jO3SkSwdCeY/UDnczchBLFF62pEF5R
HwH2clqrIManl7r24Aq44ikfjdvFZaeOXSavigcX9etWetWBn616Xf+VbI0Yhj53gmQdFAwukfZJ
wVy8+ovCA7uislkCcMAAh58snb2CLMjU9ZPJNZ92vcn5hjiCcM1WstDP0sTVN9jDkfL8fVI3gWec
Ex45lhUc1r7U4GsmXi/fpCuNhZ8s82qiov2glIblXAAAxoUoiCLe2bDoSC7WufJfvJm9w12jjmxh
ca5RT+YQNk0FMoJ7B+EDnzFT9JAdZFAo0h7q5DB/UyJdHxv6HX95bi+961HWDFqVabMUSo/XFo8k
n6NSbvJQF3DPhPQuBWbrpusrq0At/CWLInYCFI8crQlqxcTL8tgdQwenc92E/EtlwObqw2dep0Xi
3+asgKn3ABNnjDlbj4Ft83UYSPrzLYzBuyv3SZLLddSqgLtx5ZxAhXB6wBH0kIjITuDa/qTIuGaP
2xA89/gkRmu9xvUNxjyZ68guIwvxYzvsQ7FhWWMcACUTnniMwnH1Y79gnQJ9SsyuLanLdBiPEX8M
8Rig6/uvQcWTico/AKYDRkdITfrCbcgnVtsrtnjob1X0jDhu0RKJyEIjAZYsqH6TqU4r/TxuP1zZ
NYJ9pqQJwNyxzMhfDkpr/s9t+A6vELJNlrba7eqDEcoJQaDSuyBdl9isU5nLpYtBrGapoR6uQoqS
LbbSOvbyRfONbOE11DiB3m2WZnA37FVQHEH4va0RWSXQyLlL11qY8pv+TIyRg+oA5vR2zndBm1x7
5MKdgFRWQHA9DRWz6ZVEYkGLwA0eBZ5uWQOT+vgEoDvjK7KZeVz6x8hYdtqxkKJY80MmH/cQJqUL
suCCK6It7iHGPr75e3+3JZhJI6GqfRJ5K+cXGVV1kjIJyd8OE6vZsnGV8ot1HT1V8ppr+5BYHqek
r8PCIyC2lOmOA1dBKBGxpnoP9INyzRIS/FK3r12d4YzK+Cpzzlc7Tmor3qVxCNJnWtriIjNWsCSp
6IRiUxpB2Ho1InfhV84SvnKlfJbmGer0rJy6llJsrkn3CRjynya9S9aF/CHcF1TDDfF8FSHjj+zU
QjZ1mUsMD0f6lupBUINoMh4l3ZwwlswyG+m/wjUgxa+sAwC4cE0lyqsOJwyh5RS9dK6+mGo6LKUA
roQLA5PwbQpUdV3X5QXJoQotxw5hzo9yOlKSiikg9q33UEKlFsULfd5Ex379Zc8KY8XFazj0CAwe
l1mdIs7EzBL6A2vdaY9Mc2VW6EIlCsVTuxSc2s9iYyncai51RUVXI9RoGOLU2/TE4NzkiXwOj3Wi
qBQSjcFsN3X8VlJhkUaBzTyA1Ix3ZldAtx8VAiGBPLWqrIDCHFsWFjmBjl+Tp8oF7pMLLoqe6uTi
yyrVIYCeGJ2v3Oi9+l8MiIJv1Ui7ADLx3HO2eb0j9o5JjyyLqa1tLAZke5lwqbd+StO/d7XkArKr
MVE5KZp+Nbl9wsniHGTgmHd4jXTYmSRDODWWWwg6GRNLgX9iApraBa6KcJEQI9HGLRv0swUgsymR
i5vuvmNaqBAvasCzlEd5iX8XNbI3di4Q3deAwnPuuaxq/kiU2oqxrBWE2DWONMDhCXvbHDX6AAoT
oBZOITx13JTAtoYhvgkevrBGxKr1IcUXJF/MQX73o1G61hMG51kzssyTM2D3SrL5A1DhtQnJPMku
ooPezEqXsZVIykTWOfJQrgNXAKBrKZx2EJkbekhnd6Fa3rrTofh59ucPecbTZ1BnDITX1D20x9jP
6ZRk+Oh8eMLWkg4sCHfB58IktoinsBT1DVywY4I6p87ektX2r/0m9FCkvdECnk8vYoeGMwJt9gYN
/j2pFd4Z0LuH5VinzNM5VZNCckVKwucxrVPJ+PZVqJ5fld+N4dFQN+L85GOwhbLQ1jBEoZBNTM4V
oB9B3PkhGBAfMcQkMDTW1UUTVg+fcUyEPFNlbjwpfe1vlXrX33zX8xrkZzrdbNOAxIvmrGZ0bkB3
UlcN2PFQsJAjVAFUwpPCwVm+WsBtwmCzCMdFgp5MqWY5nwVXTuTqHtky6Vf+zJQfWFnZhFwAOszN
Qq1Dm+Gd0QWAgOb3mMGxiD7fNsIw/EH49Qkaedl3MHzpQEKsGRrBAfJNrrxqMx7ZCcj4JYx1fbZi
KFVHGkLWxa4WhMTZUZCJkCyb1GI74biYb8iprKZz54wFWU5jDkyMpk3QBMXXkZVL7PqvkpScG/Pl
XbMKhL+Mnf/DzfBxGyx2SgB60i3miWdsDRga1ujQDCzLe2NTeTAO2lJWPVIPHP6v9K9fAQzZngSv
4gVOV+qAgMqpgI5/tnmtjMAkZP8DmIyLW3STjYHe/hka8Soht5S/rYeSwwcDfINoH5CnQOny0p82
mYJbMdexusS+tjEXtNYRGDDBGCRPE2BL9+BWY+WV/QTRGfqso0WQ9tsYCemLYh2UO6w3Ha9fpPMF
/P7J6Plrh332w5F9xbqXjHIt9F5X5SuPsTwjvfQSY2nSLzRjvvB3GjwPXg3l+Fj0KqofDv6Gb1Qr
TeGHlSjQvrOnwgy0qXE0ZyvKUa1C/2Scw9oPYpffy+I8LLulurZ8KqH7R7gwGJqdUOOxQ6nIJ3Rt
DZZCW8pYH4ct3SlNMo8ol17RWaLPa0HnmPaxoxr9bGBg+M/aQiSToFtw9BmfzAFhmEpY277nUjg3
6B/hvK/RsIaZqtW8JxY8cy1efm4lMZ6U50z4A+WOlhUoyEbxIUFzO8/9tp0RvhTLPI958WVphpgp
sD9J1vUcBrsJFI3h68AX4/A1M5wVetpjOIwxekd3N3PKN98R6mYUpmThg/f7Aa2teDe2o39Yv/fM
sUJaqn9cBTcQb1uVvQHMaP00X/FfX9vNVH5NMs8Im+p6kBRFHSKz+70f/5FYalJ5jpDj/QZuPAWL
1X+2ofDPaSOz5MfheUeVfXhIu0Dt/Ic+G5gTf4mNhUpea8KxGXSnnA0HYN1VwMA55A4cGM59cY1J
R+wEO1GUycaA1DH6NiW4oV2UvBN0IBv47UV+VlvPmQpWaWnwTnhCOLClV8KCWPK5vO5YsNKeoD8S
f04ZBVGb7ofNhqx4YmbnrZBVoqTj3ttk1zFxj5Y9EOh2y5AgiPCNd8KotOXeYE807mbRh1x3u5TL
ebMcaOGiqeJGPEuxt+NyGyV4se9B4K7Bh7rWrvgFRh7VdQB65jtLm5dCh/bKdtH6dU6upYiZ4pQN
DCmvfNOZb7shWceMQZqhENerf+pSxrwE+CJqPT5DyzIJVFQ3PfW6y1cadMLlf2Y1N5mXR/lHFfgY
CQCltmPheIUam8CAFcJrfTL41u8TdCEfsDFzD4i6PtfZIAHhlesILUPHMEStDb5AryLpowQRj8xz
EHg2Zhvk88MPRsJDxyMqdZ6lzXeaOq7e0gbUZqk9VIxjejHspFsL5NcjjpSEpCq5DTfv6g3Jursr
aSgL2ZOGK7NmYK4tuna9ni7Dl6Z3u8vpQndossUI2dTFEHqhJ2bWexN62tdNNxf4/ex1hY8Od1LR
rX+vZx3ETTRzIIZ0gkFmPwRXTF8/HFQEn9+i/1nlNsnXLO1wACuAG0rUqEfbWqQQ58WR+UnDnUIc
5N49ehHiMbQpGIY05QzpPxN1BA2WsXgrBNeGssKmC7Xy7y14AxTwqEYQ4VuSvrVMClbuLDTJlS7K
nrbxVW4zuKfLgYiAPe0y3ZwdPE587PlLAgnRKLzwi22ahqlhEpxxkvUf8qL0vmKJbtJAYYWlMyHU
XZYliyvTntE0UFc8ott/Pka6OOUCHOobB0A1MFxYjhlYXlN/OuKkJJBn7kXgP1mH7f61xCNdNVrP
8u+jM/AfYz5dNHBkCR1uTyClYC7W2vWxPSpyhCIa0zBYqSCy+yqXasE4n0XJ3UsKaIJeKGkc242R
0RO2ylodLwHPd0f15YFUXq+Zdj0PN3iIcGQa7yDchrq+CiAqwC34Jc7+ECS07Zx5Q4PQAvf/2wVx
/gFQ0uEwnLqwUHzKwMsJYBRssh54BQMjeEqXOhg/UVSISDMPpKybpLrnRT62PadBsIOM6ZFdkRRv
gEZhGFknqWypHQB9V8l0DBPGaM3XikolnEgJ4aqWB9xjhGI/FsgHhLHZ0hSefd5dFOBRgyNYczzL
l8OtyNP941aasOeB4HVZ+tPgh9jjVX3MECCtsNnkQpWRLY6l+acm2QG+l0AQP6rH8dehR1NgWWHz
XTtXZv0bRwQw9v5UUBakBjLhoveTkc5I0ZE8Z5hz89ILX/CHKkzmtJ5KqVU/0yL+QnQJmy1m8k8g
NvQ1BcitGU1uBqz/VBNA2+GOh1XFlwE4lMY+w3O/T/FbqNUdSJJk6SkAC8VZtnzrhlnPNc4TgYhv
QLo3JQSaPDMAHmqhqF3GO94GDo/ZeSQb/ckZjJR9pKx+0EwxDkcO3NcB7M06J/DpCcVa/9506iQY
jXy9DUBX23d9IYp7QcYWVsvgk7aNRJgW8mJv+i13COcIkcPsXfMvXDVux5E4RPUINKpQccOSlaH7
MReplQURZ5rgERVKe5CPSMP60FYExiC9AUSLcstY+VO2Cem6Q1sczeH08PQwzYo/A88Zm1Jkr1ba
8IvtsU8m1+Ma0i8X+ZHXpqOaeQgNIplC68mIv8hLs8+Bfmb+r+CrP7LCl/w/qy/M1hneRhAkSwJ8
uO8cJMXScUtP/6nqcuNj3wAA0YdD+6JjwEN923KqoQteCnVr9F0GCIoVju5HHU7hzI0r9xBHibfJ
y82XSGaKgeBlSbCv2ahfD/tOdUMDsMVZjaouo3bbjosBrRzWj1gcqdug4ffURW4ztMwNGowCE+0q
fbc2kggOuKeetD5zgWxOZPSuSTTMU4zrsPh3UuPi3XQpitsUK2r6dxD04dTXJUwkOxREZHzOP6bs
6jLY4zEkjKAHx3/RyEq4UZ0xSPR/b4VjD34dHpHz6c+9JESoDV8Jd7eIxGKQg/C2TTIrFmLm8MWE
5KohhnhJDS11D+QEIhmNuO+whUWP4K2wDwADsDMxEA//3uLLq6btiv/WZgI56RVIzF6/n8UuJCqn
qwmGBVtwNmmPaCaTu2Dy+7DbOZnn07ZOmziDSQI3RmDx//G8da0pP7iSb+ML+yCQO3cBgmeKpLvB
8Zi7Buo39nkny/I0iDE/0CBBL2IduRsAFas1BnCKLKJWxzhioPC5umqnvWej3xqlLw2+K2+cUNUu
cU55/kHWtyOt12ZGZbe9kukptR9Eswx7mWkLtekCSF4xS+NkViWfYpqTYXOpFyaTC/0E8XK25odr
we2A0tm8AOzxKuNbouuYqJwSZ2AhdhNdhWuIWzY09LabJwR00edoEELFmzg8PlylWzBDiJjIdzaW
zOkbZql5yDHwQknyLeV+IMoxGXp9ELkmUi1LF/sX68okro/GLD0LLYg+8V0gVkz4Jjq7j2vgzxqA
AN3MAaSV78cRwXSvvNRv2m8Pos4Fax5cxUwLrpWDewQZ6j++kwglLfFncFQ3SaQPcZATlWMD8SeH
YD05fPMDzg8kFw3YST4uIdc2mBXvPrUfDBH7QBY7p/iYAI8i6Thq64yDaI+cq98ZXkMeLjxAmp+r
0121QGVQ8TLljqiZOQcGWJRBWLM1+mMAtup09L/R2BPZud/qKbsTSOv4ViuHf+aVtEkNqzvBWIuA
BwA5bDDvx12Jr+Wu122dk2TkAl4k61wgfvErJ7S0r+T8zKgMoN2uqVePJ+BBtzMWV+HtyhrsUJ5U
0WgxQK5vuKRFku/XSJFFpznd78cbDIeS5jbMwM5K0awOHseDOgesSjBrr135iEsK1/SlKUTPuwOG
wA937nh0EofR3YFRfJijRyN5ay4E4a5N7c063UsG00iTeTlmNwFXdPcVSN5b2q+dfSw56w6zTYAq
EwD+cUnZZOHjb8yMmdwovbtiJHgzt6nkEuS4FpK1EIAJ7tKEraMSGABwEsRMvCZ47205aq/yIfBZ
NT3mM7akQcC+m3n1LimX6o4/QJXjh5+WhWHVBEzJ37HBrWei3hh0gyk7mYLtatGNLrG8LAPKTvMS
0c31wv2AuFG0ZEBKGddP348cEyYj1yBu2cXbzsd/wCXpqv5WJgBIwyVnAIb2r5k6fFfg699v4Y1s
JEm2xgQm4Fe5WGE/YxV7L/jZsP7jgnii27VEQnvyVc6vxTC+qrQv+BZyTf/mdLpkdEwu6v7cSJe1
5BXFWC2Uo3bapzRd86w01n8qR89zD73RvdpYHEHsKk98DUR8Frz+bghZh3Fvo91DIeJqk23fVdjW
IY3ntWoODD0YvyUUOh2ldQRvBQoUQ3th+8Kzr6t/hSQnvRfxY0lHKAbHBRgUdY97C61tlywCRudg
yke77he7cFet/4tcwYixsUEppf4+uY2SricakaiBum2BC/JIEZVig709W1fdKek8Cu27e1bmzRjl
btBb8P5E8L8PrNbAiM3lBjNGXVbLwH2eO+ww3ayWnDffIH8F36UrtetXGpBw+PfA7W+Or1vuDH6v
s5OA+bfZXZGaIBpnEbKx/JJ7w+6ldkykIAdvqjD2++VVrMLRnC/2eztO1jbfoW4TUFbCekWLOzgd
TLpmDbY5yU8Z3TV7Eq2CXDwXa+diS1fV4G9D1EhaTxCFCY9AX8lY1DOdyJ5QFLnrsv1siqDFZ97d
jovW7s19mpuG0tQHrXTV1BFPCnoSZpb8XhqPI53YnNyuy/gF3SKDX7arCfNGEChWvBopx//kYmJW
EKwl3B/3vY2sNpDxvZbf9uByM5V7n3HSjdHKDQhVZF+zlPLYK4AR6+gAY9R7zMFKxizpWegGv3xz
9r/uyxY4/l0Z2EmGNvS7YzuDvfJN/X7vJqQ2kUSfmLJIUuajLnjRG6pX9gJR+bu0VCUVAKy7whjA
JIkgvxtIIHshuFmvv1jf4OJSLQDDu+TVetxJfAlp8ESAeokxjzkNoG7bKGLHzg2hsUlTdap2YGrz
vGvP4HBjuSDA3VB6IznlfmK1i4rhejnqSZof9J2sQ9X/EMvpsOlQaHPx4UiJ7LzvGx7icayYWPCx
Hz4F8SEtDWvUs5z4hjWsR3hOosT0VOu/qQzwmT2Y8ZGL9IFV+bgBK/nUvaBCdLsG29C/xBCg7lkA
q+PrfS3W/3rOaESsfOgTa+Kzn6BBL/Gf8SD/uyD6AY3bnlGmTV2iwL/TfAPjzdP5AOV3f6ULMpyl
PpFGMnKAXswXZBEX7snt5WoQtWPCWWxq857YbpkvGNdMeGgahfGPbWLMFaos6FDX3/wJlbI7febD
quqKG2JLA6giwETPjZmVkj3dkuGsg3SRY7pbt9NMgFrW2TjSa/a+B2dTXlF8gkNpaavoLQ3/H1MP
K3PlqHgKcuovmiW7SHaEFHGgxe3+grBOEOA/g5zWf0KLUYWYpCyxFcYiosRXPisxTd7xFZyUpma0
mjE5rLkOwSs0XSI5YyE56trkEocaa6wrFKV+aCLPDNmZ7k+mVRxaF7vUAreYd6aGRbL/Ry0zsH+o
kzIfe60MXlobVpCUAy5r6EKDOUaW8GgvF4hUPiG4/CkIiY+9X8A5XXf4ECYJEY8TfGAmyyuBuww4
BuMN3Pf4T4NMgfDZTJRQxa1AQtnLPOaY+7GyLMAPBizjiH1tCB3mxIhUAyWqs0d4JZPBhyF1ESiS
LZ1Z8BOZuKXFHRJCFvapXsoPycy0/EwEjEufyGRRRpmFcxXmPcahW6Km/0a6112GNeb6cWdXYPQx
1lic0OT3i/1C2E3OhPbRvv+pl4HRP5lvj4Ffj+xKoOyKJBPzSB6Ll9Ksk7FwJ+MKeRqUDkKd2ZjW
KJEp+JufbpovBbz7k74uE6oGBgKRHXY+opWoZLfzxhI5crAoc8WszBs7qVHMCjT8Ti6GgJlNQM3C
51CndyFPNqZ2kFqvenjCg3sMMWZvwXsFp28+YWr8tKKHSYG8i+fjKzgeyNv45kogxg77cR7GKyoz
Uh8JLHLvburTWCk2gFIl5x4VSnhRMcmsye4AHriGVLNNXKRYfXnSX/BkXqsqhGORGXBS1jINFU9U
HpxsCZ4GdSDQzTzUpg80EgtNpD4/YBtejph9Qc10h+IObC0Imw6NUGnVQkZszbjDT8r3oiaLWdWl
rsFPgTd9DJX0l6W+NJ2+XpjsWLbTzaZDq5ey3tyNFnXmLk5RcSKuTqHKiNqokhgcyYlH7Wa7q8TC
7S8/DLB7zkusbMb7joaz7suJ5ch5UL3h+w81zHnIhzxDMQKVB/cJtINQeHWQLyxVDfVO6m2mZkLl
SvqnwLl5Lzj7ha/414EZQXhxi8yW3UfN9L6IK692UL9OrmIB9mNOXgoQ+E3sgARLbIQF1a8nt/St
GZdLMi3z2aOWXiTcJn0fq+kyCby6J6xoggIaUPdCc2HyqzsY/aU9nU3TKF08lxSrSVJhMat9PVpK
RHvqflzV+uUOKARCUU3RvzcyCROKVDLxnjr+C7dCMjSte12kxU0paDeE5HzLJ09eNwFEYnFFr/QN
rG/SDezI9p13+JOcSigcnc56rsWRtdTBVkoxQyEwYZfe9PjHRspUn4TQr+McBtJMgFvZVKB+uHr9
pRw3TeVkH/c/NVZfkJpVYjk/n3XXsG6zA0c7N2WgZi2NKl5wQtxwsP5jIn0jhRkKF7f3iO9nm+gF
ujTJ3PI/fOHMhxw7kDbnloO6SWTy3ahfH5C4GkBRJ545qlfSkWTk8g+3Bqm704smWBVCIuR4m5NC
gR8RgenUrfYPiWF2sph8zacqBaHR+0sh1TEmyeyBF/XuJvXDmoWRJ+JafX5eBXkeB7JafJket8wj
Uh7q2JYFNB5b+VzikmjPk+WfjIOFHdfFvoV4dZ+r55Tc3lJR+m6Vmv+aOZ8rgu/rngwvYfDM+PrZ
EBjpoq1Q2bfKs3CopR+lzVJZffpqlG61YLyNlvstlbQbQTl5471xG14otbfDJaRsYOBdc5d2hUP7
6KUZ7ZEx1FZsYkkz7A3FDAJzz4i7TYTJsXEkdRNeLtdVkBENr6xLn5YainLse4V/Sg7a0nASB/f3
6F+XUfgmlAvM1NsLdj58wxSyetoC28XRluGzmF0DTPKndRvI3VOYFr+pi25SLjj19IydFWsZcg02
mvknWdkGHN9pPMM/GFH+vmb5/UljielUXb+RlRA3fpzLqjJIFiqi5MqxGsBYVBQ7iMwFf2CuWGgJ
H3EKi68yLq5D5cssEhmYG+iV/dPQaBOlUAx/ANytQpukfDkM3DmEiDhQiaKouBA70MqkMQ/xVh1e
xqvZpClBHd3UlEJSvlkdJ/86Kwa3LZ4oxzrMehI3w2VFr/oAuOjMdKRgIella38XaLjZX33UsNdH
XPFtIi0fhfXdQwLgkFRelwMfEXCKuWf2uj2d8Yim/tqi/qRHyMcgsWbg6WCJgYM5Sh8TmCwDeZgq
m6fAHWa+dYu9oY7QuSxwYBvV4HRu1nDoJV4fyFZ/smpoMpLvTxrPc6IBAGd7sZyw+AEz5F1GBPxH
x07XPTum9DmPkVVf+wE71rXo8tH3KANnn0tOd/0P5NCKB+SYbv8QeuvXJbR+sceWgvt/312UL2SH
jioZv42uLASa5dKGbqO2F/BA7hWVttsIun1kHEZDfulWovIi3Kx6FWQjDneGT03J4hyciqbNwlt5
K99tszjHGE+Wdi04kWmD1P/8Z03ke/cqjYTZIO8TRgxuUICJCOQaPblnMIUZWImT51R1muo1zNmm
iRsPTPlPxqEwooAYJLG029vKtFsfj2uXujxwlpSHa/zhZhDtmIHhq1G7zkSqbbgACw02hnjXgfyR
EqtC41+ftRykdIP+tMz49MPGnpxUqt7Qk0aC6CYqR/ybhGVMbx1UlaKdNrC0h9JJp9YXBAxJ/Dxa
6mvsVInuR8xKAoSRi2d2UQr+vIKd8pdyM3fmYRTTaPTh3EsqY6vXcIJt9FXyhUY8wgyQk5VX8nlH
0Om3v8zWVjrAgE2roL65oZcKHE4xfzYLC45CJTgucL7gaj9BuU6Yc6dphwhCUQT2rofb3TcmtMIi
+ayehg3lfNoZ2slVNm+ipN8mA8TKBRFU74DrFUSyRyzXmmTz6lKXyrrKcIhgBCj5cGHevoEcxbDu
IICt7rMXkBgDkCniq2ZpxTd65Mebf5hnH6I9LcaIxA6GNPjWknu6WzrhI+oVySlllXFIgXz8fpgq
1QL3r1s+P8YqcKVN7DQkQOg+GKa83UIVPMytll1aGqaqGKmnaH321LJqHQ1cV+x5Oc9eVkBrfvEa
rIWYWwEEW82lsG0i1norUv7ACj3aXEswfOrxARKAwffDuFR9yBxKle4uw6d9+o2jjcY+ROUzoakr
B8dib6Tm4LeIe69TJK12lLbEIvMGN8qErHcaWFffGp/5trILifaVjeRspqesf2/ErIxEmAXFw6Yr
D5U6BtR/cV8V6pDbBPpPrnEhWmGyG+EufJwHWRib42V6u//BJ0l8PRkdATvSbfhPXL8FCIisSoaE
PyyofEURIWvHnErfIGML4BpsxbGSvIesDxh+m5YtT6mUz+YZEyq8YsMBBAmGY+nkGvQnvACTHrj6
EBsiaZ/M1qDu0+mhjYoG+ZgdtzBiDjsIcH/3Nvf/MEOcRRN/JvGbYX6OZ20Y3RPYLAmjSJtL3ka1
TFAFZXYVOJ+RHRN9wofffha4Y+lsRvBW/vn6zQEWuM6eYzQg69BkGX3zzIjWB7MQGEmJgBl5P1ov
sxD1U+p3+8/XWZGMrhRKOi+n02XBIpiEaLmsZrIThUGX2wCxrAH3gwOQKWJlmmeGz1RTWAxIBsr6
jl2QOjFexoBPhR1ciNb/rQ2UjgKZ7qrC7Zfx48+RoFrCvFLHpAJ7nznbM4wf+CRGSOsxML5xWwZn
9Hvuz2Ue2tc6SzyetVsubk5qiiaCcOI5Acf+sEZEksFOzLnuHudnFv1o6diVOfp2vOkhu0HUB4RZ
lzEAK0k0ukNDlutapKeF975hSLp/TZd4Zyz9zDHGztQINaU+vCgVISvk5njC+aAzAfFeSvVufK8Z
Q6KEuTP45vp72b8ae3E5zgkn7SKFX/1VY7Z8McFTJZTqQuoSO9Asy1bBK6/EKqkLpFCMlGelgUQ+
1HR7lGj50sryTV4t7Kw35vpFSgzb3hruSNKdLrR9gOg0J5PRLskGLk2cuJ0HghgnBJKC7XKyPIox
5vpYJD9JJD2cZStynBw+xVQnrAFDi7tYHdWkb5dSI9JAKLsUR+rr/etA17jAnIhOz+8iMUwPobKH
qFRIh8nKnkP1yBFqvhu6Yuu/f5XmZBJwvZYO9FMK0NrDda9UwCxzW4H+LASL1aDmXia4/BfF5dNC
IeezDmGKbd0bTsMAcSr7HgJZBNAnr9Mjjtt8EK4B6365jHbmPPWTfB/uG0OTJ/Z4Rfps9BWPPXIc
oPfmJ7X0ka6gssrz5Jg/o49micmSWXvYD8dRmXRN1X//EzQtJI6WkgEqE1uR39uB57TW87iB5zLV
eH5nSnYoRVTDlXozpJE5ULB2LdKkEPoFdV8DyPu+ZnnBCQRSeLo7EGKan5i1Yc41dnYdtU86lfF6
n0V7/XZ/SCKFUPhvtwHQIjhzzVyisy8b1n9aQQwELUGNqJb9DV3tBI0YAETVAgZSLvFljM98nBUW
n6iD7lCyokCCgjp4/N+GySEeyUbv4rafh732q1WV3CGQjaHMP1lH3tSPFRuEvIIB51zGx7QUb228
osUwUoCGRDcCU05H/O96KgbCK1xM+UZEGugAnqhPe0BVjGyD9dpbOko/aI732m83Aa0Wen3s7az6
7Tyk+wlDjRTPsn3TD7qO3Kq4lWOrMhrrjF0jPbMP9T737uYvnsds/eztG86zN+ilugur+TNs88Yb
JKWUtmtY+ZguXaolxolRrUUdqinKZ+J528ouA6ZsLSgUEb1Tgmh6R32++/5RTINdu3cYJ7XSMiD0
0q8KaXkb+9E+YvIWN1k18vVIQ/+YgGUhccolSZaY28OvuKYkJsPeUESjMjKpsKnN8F+XYEc1VUlm
0zL8vGTIhBVC9ReWeL83aggSxg+IisRQSCzT3XxKKKyPJpzATsPst2sUjW8bYOJJsHKllyOyGDN9
cEsSxJ+pwK7rJMai7mt8SnKwAGOAcn1c3xbAV+wQRW1xep3q2TrapSSlBZ+crZbvT7VToYRHXus9
KIO9RT+4Uydg5Te3+qaTF3OR13RbaldvWxIjKxXSI+jFSgTEscT5oV5jFhwUi7YLXCZSJ0tz+vLo
/nKVdG4bQs2KI/egE/RvY9LM+z/gWUaiDC2FHagPgOtHwNEF508raxWSM35kqm+QZ91yX8xsLSNa
ru+KZ+7xRbTcZaBJW9lWbZnjBKETTteuRqH0wbKAPLhAj7eH7SgHDsLoc61ARc9ij+S9jSJK8/rg
rY4zWMVaP6jdv8zfjTn4O+5OjYyBBZtaede67kVW+khz4ChvilUP4E5bh6wKP9QQehF89TwSZkEl
icTUXGvRCBamAz4ilI67FuL0J97m2bzqbblWtTacQPi872pktiiWihBBEsCzeSWljwf36PbvA7V0
nRAhmF+2wjGundWUysE4RveVDVjV4IFX36XGImcdNVWF40/dlacuBWJAN6bp6QCUlpl5y4nD6l8P
kFCuwed+uSKAy7yUXjungcPRduHxNGg23lC6X6M1472E1557vWeYmLcJLpK+NJ/EwFsQEc/tPltw
BnmF87Yui2HRGO+ZhD+iAB1pSRIweHtw9xvfrjAgkVJGcF2tdrXPCP/zkIaR1q16703h+7218FKm
CmCRODapsJHafVmZyRRiQ3g6YwPqvgczfFdVpmXpMIQYBxLPROkTvTtsb+VABSaFv5zBQ9gzaKGB
s90aAeCjEnlv63QvBLOTMk66Xf0FGHNg9WrnBtPStX4c6PAlpX2b6oIzNNzOoZYh1MibxlJ3lM/b
Kith99UiPZOh3swtqwe17wYu0EsWIWIPOVwn80MBnGHk6mLI34JQyJm31cWBDm6THRDQPeNk4sb4
EpAXX+W5mWvXF35ufl7FP/8dfOkn+ywz6xHseZdxCXleb5z4VLIoNa4zsKMH0MANApHUAjSUwzDK
/74DkYWUTh0M6yUjroiJ/od2xyiK6BqqedUY5TOP3uXJW/bGE96wEQhStBYLdE/BVeMKl70YCRZT
L//b5tDlxeAFwETzCeKemVNu2jEC9z+UUxjGIEs+NXQ/XQEnONL9+GC3CQ45S/Y4A4HS5UJUShzN
BQ8KSZt89+oTFD2o7siBJutXC2Dcyndkzu5d+qgV7ZOvUSL1tKA1bGkaCMEjz4WfVvpOlxlf45h1
fsruXFv3hs85Lyms5bfzQde8UuKBeU0XJSZhN49L4akiMc1XWBbgj6Wxcgx8nQv2l5Es5MRjoxwG
Vh5x6dSeP+BCCdb0W6zW/6g9Zzm0JOqaFcoJsbdFDlefeuhf6eMyALJrptu9AiuSAULXgXB3Wu/q
JIkSnozlne0mfo3aJmwGdQXDJ/cfg+42lYYdF1TzxiZeFipyZil0asRN4xzymyL2Li8DIii0mYDt
SMw+uH0eGpSXZCa4LUETqBOUImdaLFjHD9TCfbbIbJ6Wxu8dsi4f6PsuHXgpOa+m56qBODx86e6/
3AiDZ7mIYYXQ+vUV7Z//EcpqLhXueM+pMw7365QTjBjndSwigFJBWCN/YccTZtuiJtMUnRqKhSbd
cQZyPz7a5XNah8XemnTgg+PklU/WCqgZXu4p8lX8BX0G8GMLbb5l9vbx25R4zFjH7dbP3GGb9mWv
4iPGHQ8SBzNLo3t9VW3v2CGIZbs4mHBh/9tCGOxu5j7TOBX5OhtMLloDUncL0k5jDa+BRhQRZU1z
WQEMp6zo/ZO4extHfnshCJAH4Mds6Sx637zishgZxvj2+jKlCZlvq9vd/zmVOt142ldFh1n1XVCi
A3Ye/qREnREghv9YgkyHYkjHDwxrVmzGr+n9VJgfe+zj/Z2XzN30huoDUwEHlB/A0VgpuyBjgxft
Ls3TrDxj2p7qgnV25vLQjHqc/c/h5JZPvfuzm9tYDPq9hw1n9KoT0Q/RSWFy5rNfzJf9VctjB+qK
cifEIyaPsyeY2rH7oO6+a/Iq7jRP/YbICTz/BSZOQjduu0aywNY0mbfnDdG16nLWCAh3NwBPDVOt
xhlqjA6894uNUMbnH3yFkAlz32mPs5wtO4/fI/iICQ61MIXLyiq1Ec/DpkcXB/mYZMw9gCIgmjvG
CPRn4GOstjGfFAnc88RC3mhN/q8yrSjw7MajrYbHtLxbFHuxFsb1sZE4f/5+WoP2wFseMk4IcAuB
GObIs0idtv3o8TXmw/l4YByTulcjJpXC5M27Mvd6j4piHpqiaKxiPEzuIo5R/IH9n5K2EW4h5OZn
oXgA6iKlNwdg8NkecAn9kNGFv5fCyJoJLtTZ8Mf/Ia/EPi3938PbvQJ15A8sKAkjOnPry7AjFztp
eVSbJFtaotxAvX3hGgwGeIdG/wNj7Dqzny5kErfNb7/9zm2aPMVSa5rEf+xlb5EXiuLKyC1MMRfq
+DO4jP93E3OeOLisv0OfhBP7jseQh1xCOd7SVMUN0eZrch7paYZHtMTOmJCBiL7+7aa9HU0jCpkO
zlXkLeR71DV41A9KE9efGwJ7EOl+gC8/VuEK80wgk+RtrhxdjqeNZC8hdRD2IDCovOFNUCLKWxQq
pnzqYSw/aiNDBNyYwapcpi+ioVp0mwWKyjD0N7BFopHSOnrpy0JUYibyYQI2WEoIW2dw+IPMf7wC
Yfz7IdXfrq5IG4eHpZHfMnHquRWI2a7/tpC08hOcgV7UOQKPWoKJlXxyiTuYP3r/goAbVip8T7+c
SfOAhna0cz52tWVlJNmycL4HujI9nC4VcGnU+6od6vOK2swVSkGwH26fbru1gr+JG3iFDNr/H4yM
0aImIus3rrpkD2yW7BRSz+LtZLwVjjc0qaHD91KtnOOvRPyCqIVkj6MG4HlhDh2kRqlXXZ47vO07
YYJOzHZ+IbVcreVoDWvuNlnUeXk01QqyOElXLTSWv86BYQs6CWtgdm96Rfw9Axm8zuBoc5cal0Vx
HsLQ1ljVSSqpxrZsPfuS7wE622VT2enr3dE7tOb2iRo7XqyFGyhRSKD+DIbX+HwfFZky1bH8wNds
p5Lo7JxWDSf6jzVPOiattByOjqVYS3ZHXilWQXxnHUqEkQoqdnX4WOpZn/+pcfmMv1DrUyDb0EGq
Fdhg5mXCIjIdHUHvLJtwu6Ljn3YzdyEwIShhtln4WLSOI34QhO1q/FXNMyiNQekS3b5mXKdGQakC
d5wUALk8D/NiStWbhpGjhqkuVKXEIUf0vwXwfGDWQ506P+EmEa8/TksnQjXRtU+1a7S/k17FB9Ol
0FgS8v2TDjWBT/YyGQy+HmPNdcZRQ9M1EcB/uq9fm5l0RHGuPHoENhuaoZ00FN32pkfX2xUDUGoZ
lFSUoFqkKEj/XVs0bZI4zANdvfZ+/AD8lUJvgJ1nsqEQO2Rjdwxo1e7kieTeWL0KlUEu8vt0rfHT
COcUi4vAO22znPfv5v3zOyE0KtwHEEaJCjWXXIHI7tVEh8P4MzkdmZ//w5fyAoXLOZ3ZNEHAxYBa
/SL5R9qXd6+Y5wl5nPOxcXg1tcZYND7nwrIsX+ZYcqVY9sWyXwNjqWYLveCkUMoiq0RKkcS0ZxCe
CfHPO2Ju/MaL5V2mSDax4WFmzg0Jj0nN6ZU6wR58k4kzpHpIwEp99Mo453uMO616ZPcMj1KfkBmr
ssaJ0Ty/rKfhCUoM3+UvCuGeClJo1RYxBnAPtk+ch4dR6x+aAGwhsURg7HC/xUkjOnaDoXXlKSpw
LLfv1DDuumbsIb2JlhUdYl+fAR7WL9Wyi2pTEVwKDW0MuqGKkcrUnc8x24vtTHNJiQcEvrsnY1mM
7QDs/XxyQe2IXWAvssn4P+nCRIebHFhh1LKVwXtI22GTiIl30Nb7Kl9lIixEtGYrRDun6s2yVHmt
vvDL6mFNma89B0eroF3Yvb5jHjuV/HJs00EFHkPrhPfHI1pxF8mzIQA8woLcEs8Rt/AMcFx4c57a
O4Mqwnia21EvP26RygCbun9Jq1pibScSncOwzyhisjRqQxnFLzCsxLhc6INdX0DgeWMmjqry98jn
5Cs6QOeBeXBbS0CeOwL5HRRQ684WPL+JhDLLycrUjWf/91rk4rVjGABSQ5JG+99oyLavccUbUz7K
pbFEkf8PM8wKAInxrVLNHSnkphaypEKoX9mgUWfaL2KztoEv0+fpwZV/U+JX0ZcmVskQl7mqaNYi
eMq8E+839lgh7VdjYIB/kEUoRVI1rXBdIvQbMZcjHy6y6UQMMfyockeZWIKmtMnfosVJYtD+T28f
42wdhV00qM4TeZ+RFtyfy7YZW7UTLoBjYifjoiblQw7/dftivTov3qeTkipV+nKLiXehTweiQVNa
Ba7BYO9tLC17vm1U8VhLKeXryi37PGejdT5vP/uUkOi7IOWGutK9O7sqjIIVkYGk8Xvs2vIZq96Y
9ANM11sk5e+jte+DlXlFPU5SVmMBsWiq0Fh+i4EX/aLnmAiNHEYN1T/NfY30N1IVrKM5nmlqdCWJ
IBhnOJ9svGkaxY6fM9eeVOROdZolzALvVOAzsFutvGa/upb/5VgIRzyjCUNvzsJkXQGHiHacNIxA
hqs2AMGfb3tVGg0A5c2Is1XNNF0GuJnDsCCaA4+DQSDoCtdhv2IiFpVh2M4gPwHcRxQRCV46c4Bc
AhW01nY46mkTanO5zdEUSCVSJgrwGh2MB6Jqko24F9jf6IfbyssVNl+YIFrIKuFL99SjgtyNCaLb
ro+K2lKdnPjvZeG/9ywjTM8EQM+v4X6pESGMsxrLW/Tgq6WbY4nMPfKYAwulK0gX43yzCmODYLt0
5hIRZR9Nk41zVjkeK9JGLc00RfIm7jJm2yLMT1TXE+kCew+tocoaoSDvAwPJWA0B1fr2+vR1OyFW
cIekhCiHa+99K78ljQw8TMeOnygtprmAC+kHCNgivARbHrdwFnyHezqOIhcK0WjDZN1dcc/d6O7j
rvZsZ8tdoZdTXrhEOh/SoI7NziPFeH7NhpPx7hZILM4GFxDk9qTMA/sAxC9EUzmjlFR8g1qxWomV
/Cv/gEQzMf7cRzMHLqk/10i/8magynYBQBi7qFs7P4SSjhIwZf3eMIuHItMZEARVc+TkNWQ1uSud
vL29cEjGTdZmNFzl2BqPGl9W4LoX422hPRJk0lsh0m7NlJeA48KiGEfyYFYY4WXafgtmUJ2Id5AE
BDm8UqLikO6faH31YxQD8Zj83J0xa2z/aCfkmVZiQe2XqKA7BVS16LYzTxRHqMWeDBU9xPn7INL2
ykHKBJ9YbDVoy9Fy4ip15deeBQrVXNYVkEDRXLYduxgJij4LFHltNFqX457cI5xG+5nzzrnyCes1
Am8N7PLf8GSX9taKYEEkRugzy4qcUnwiMhXcMYNCk/ey3Za1b6qTiYgHATr+StHWWTIRrakgxp2D
GpDTPsRkgm9ADEtC98rE7dUBnqYaVvB5VozrmrvbLW6woNR2ViEq3b3bDqmpuRVxMvqA3L0pXw3h
5cPUFwynpPttF3zvCZOuMwhOdjBOONzYrKZQq+UEWf/vXxETVFqMzy7mX+WHaKQSeAIcJ455lNtA
TlHg6M/xj0DBmp3X9FwrjSghG3zuVOhEw0D/7i3vr0nUSA0wC2TovUoaGGwvSEI6HfY/xwB9iKCY
v9Fs2nEFQ5OX6qeEJ8zZuU0mMJxt3/kUzkA1aazKxa3u6o4OBRtsDAblz0IlGLxEPiv4BasbyVWX
fuZRr1xaw90ajNDbd0DjMc8I5sH+cad//phGSksehEN3QdOb77XQdE6vRVqacZ5Vz3J5tlsogxHa
crAl9etsCRrTpbtH5Qh2rOReDsdE58/tCDAWDpv4r0AJ9JaoSO1iY94FgWn7feaMCQLira7+qq0V
iZweIpM5IYp27VvfEk/L9a38R5QBl36MhAHTT5wEm3eyCM7p1noi0CkoZHBYcTE91eX1NSiQed02
4wsWsbFsbulXdQEHtFHa2bITABbaC4XDG7uqmDYqHYH7zlQm3EJVIiP6ixzhO11qdNon98LVf4vb
A+KB5TJqf2rXS9DsELejX2z3JI8Ibb/sYRE7LcR2kVrMvNRVKvUmcvSRUgW2XdWEgI5WbspWsuQ/
lddwCTx+htVm0vVTRuYKhv9XrZQNRaZ8zsGtMGqQYIObbiS/sJp3xbDTTP//PZSjJEEZDRDPLajl
akY81EoN0nq6Fhe47cxDGQg4+PUB9m8Sv15t8Mqv9T1o75vAdTSmXhvMMcFxZFtwOy73S1Dd6k3r
iGg3c7DfD6TLzwuEPhepgq/ZmeyxufmQjSmrFDps4Opg9S9STQ8sipxOasM1qfq9vUuIPDHYCLkH
zR3CJyYkkmgQfaAJXzKvKZ5bQ2XlXGxWWt9ctHCyBt1iu8jA+LfNQhgcNpxBov5p8QWDoIFcsRHf
JJ8oFnjmeu5C3ViypCoRbC7tegjxsfrpnywZyRs3Gxe5WcHuL7brVX6otb6CmLl+vq9eu1UY1gUv
4KjPtngMFoNM3mQnMzU0ds0guAJSPNrNa5xfL0/A22Af6EYTEBkET4pBXtjFAhFbyAkPTe5k7kWG
Wc+04GODz/tc0TTN++9jEFerlHaLM3pNG/WYU2zajgh6dxt3tbsviNOdzFY6uERoFlUAMTBAf6M4
Yx/pBzIdaPHpD5xc3FecG41IVKtNGLaPjaF0NwmTofMI7Aee8VQYJw2DX6WlqIEPVo2hKhnO2flG
XZVK6AfMjjX/e3h2a0kc92dwjSwhdvFmvmRa+8BkE0KO4prrspk5vJUDGcNvOlge7trwn96BwbZ5
ncq/0g7BD5W1h2zQ0gApg01Yw3VoTlIkG57ZFHXNbP5Rj40Fc83Dp/pEXwvRnZ2tR1F9f+pm02Tw
DGDsa3FbyWsGy8B7ObhTnLVXP2PyRLtGlKxcbDmLqxk/LfQdjl+94H8LxDse0r6xvWwyL1sGR+an
dnBHztCW1nZSvi3ICSlaXr9JYzb3LseKXD0XJt6gOMMDaPhvmF4SrjRSI3I53Ax8PvjoTsLNVPnx
D4Sc62MR4Rd61RQoRH2+jptcI3qIAcuFogCoqU5KC5Y2xn9uXArn1BieaYmD+fRBK/r7RpIUOLEk
vNhJY/vzW3dmQNK7sNWEMx66ykrp8BbAEmz+47/WkV7+7Y6sLsQldRiwODjqWvAMock84hQ62f+d
tnLyD6Oo9kU0b5CvgKO7ZPuCCXJJuPfN6m7TlR0EH8BwG4g4+m4V91ZNojUBCFozFNcpKOr8Gjj/
+jJmcER1LhIec9l9WoLsB4IV8m9l6+xRsz+24OLpnUFmQp990to+vEd1/594Wa+o263TNMlJ79hE
3uM5YyLSh4gyuQKxq6xfkBXC3OYHNV3TMoDNV6fLaFv60FOL1vPh0uKu5C0jNBKlICkHFD2BxSn3
UZVfpZE40E8CnFR5GaxpMLnYDGnvG6LCteVPnZ9+kLJR2Vj40dodvvkC+58+xUmWMOfB7Sxu82al
AcFASvSkBUqOtMM6N8QyQgf5M8dhtmKfxB8o8FVFu2FuVbH3z/WgaIH117zeY8wcV3xF/AmYKUmG
7+Kkz42M0IMrmnCnKD20XNBYR+vuncf78KxwmSjIVt7qE4lMrGZew0V3LAOf2Jc4lzD2C09uk9Ly
fMMZvu6tbg1rvIQqOQLj1ledr4n7m5W68ST8/a9oM6uzNZQlIbFkQiR0fkqwDg9NHRkG4gIJLuUq
g+8BC4gwr+nOxu/e2Qn231nqeD0icphZZZFSZTO3B2uGOd6N3PeV2oevlv6s3qn+QuSfGbqXfrYj
rvDhNRLBjyQn0Cj2I6x+u8RJtYTTr1fD9Ox86+U6OrVYI3GvTCOKrEUZ/S7CixX5pVITx088g8ug
tzVf/rSb2BmCzeM9Bvc4F9fE42Gml2h/Vj3KgNOqj3xttuKJ5JMG0nKzCRk5ZBcfpBQVQEHUCuPq
Ql6272R4Wi8EDC/Sze/3aTwHK8jH2SsZRf9g7kFaYrUd+Wo+6fSXCFN3O2n6dSm9o/Iq30KWzce6
DMvfSiz3Wq+uGsPmz6X8TZvqnsRI7YSWcIibrPcIrGgNbRsNgr3KSMuTdePQn/IZB4NdU5fIYMD3
3Cno+Ix55/iH9ePAk1H/o3w+0pHbHsf0w9QVSuIPhrWqXhagvvWfcVSZgCJeyKqAcXHFdL+unSI+
iOV6XYC2PK653//BWb9j2JN4tl69mdJEmuypMZOC3/JUekOhtZW1uUUfvEAfo5krzIDl46MMqXxp
gpDJUgmBMFz4bmx+RSyLyNmjXZV5/sZSyOPz8FufzU1bor8Q83pcZG3d5Wt29GAiFJMiIQXB+B8W
pV/AD4ykaNeyWJ/0MRpmBfn+QbfD0xddPDmQ5SlMzMF7TlvtoD2xHnGJM0iCcyxb/eKxJnNhoCfY
C8AK7KeGFQobyju22g3sgN+/XUODt4PHuH4yB3LtLRMFkxoDqNOQ6NsRb9lglH6ljx9ohEKzTDiF
6bcWtkQguc6bKMKhprrH/Fvl6LmkQCrv46Oc2PFZLsbCd7vQbcOy/Fwa1L27CPZAhtRBSeDPyoFt
65ACz9huceTjKscex9feWYF+lVoPOmqLx4HgtN38klArVyGNm5k8Y6+XR4AlR5AOxtl9P/9mCyIz
oKnKvqsW5LspKoJnkpx/b5Pf3ox2T3MWMdRY9vKzVffIUvNsDVC1zYz9jSArMGN7IPz/iuxcE+do
EbQeVtSXxcKKNVxyMRvurnGz6EXWHcskm8OJdBRRuQXCCiLEcCjm/l00RCA6dnIsyX9QyX+ly/V2
dWzW4gJnZ13uiGRuq1yFF8QrKN6C+fxv/Rnaa/9Vozn+sCkdVumWWuUUBySvXIBds+wze6SNaYnk
6sXzRt6/9TMamt1rclnl5NlIF/Xx7zVk4pbEGccjBlJO1CJBoPRtkJmjBVWmxiBAKNIc5406LY0z
Iid84PBItNSGsNHAD1V7rj+PFMDqDt06JsfPsanJW7/j5bOgk+zNjBM5qDJKr/HEk6Myiv81AsiP
/Ah+cHgJ2jzMWu4icoKFBrqLcy5mbPTZGTsaNsRwFCmdyoAwQKrpIJ8iOo9LFDAHF2cx/ewSpcv2
MZUg0W5jueTRQXGl4FJ0v6Uk33UhWTasKpPnCUxNfY+MSYUuTLD7hT6+pbX6HOE2P+hXOup27+N9
Loc2QAVCEMqhh0VhNxlWBO6GvcRw4X5jjOMWrLfGB0I8yrEg6NYSLs4QbSlHJRoXC1qNVKG3VrJC
8fwg23RkRbLutzeYXVheErrRRXN2XYJCUrwDCX5kbok0kiqK1xo3wvz+FE8I8Pu/New+FgRGdF3p
FjjkJsjARuu4zD/Vr9e0b1OC/1Zy8jE5hdkDE/Izeo7KhI17mO0N7QtRs1j858tBEFr96O28NYP4
tadC8tjiZTXKG6aa8Q9Xlp80g8L41tfiYiUpSTqJzSYR2RR+JDYY2rqzVg16l6YyxajjA4YbfUOI
3Cj5yg7v/i9EiltZSerB7xazB1IUR01Hpu1B5QkMShajl6PZxD0ugNK02VpG4+4jT1OIIv5WyhlS
zpl5wRYZrvW+jR2avR+H9R5kMDjdIslzu0IBz1+CLWz9hbgD6mTsuYrSNAxHxP+iykHGnSChKsV2
L2gku68cDaZORVKTId109UMN61otPYHIVc2kz0zfW9ie1xEE29b9aMUSNLTFAXZ3YiOq7Ebq0zmm
IFgJZ0vslNtEANInUEkkUFna3f76fJ0bFLiUWLkWW4VUXZ8TbPzC4ktadMO43067SemAIdalh9Pf
unvTToB0UbhJhcIpkCBsLpA6QfgT6oZvu5Fb0gNJLgmr6QmzPDCcj8h1AMxb9bp9qdk1RYKSzsKo
eneT64xUYFk5FfDRTKA4Eh9R8m2/b/iHOXx5rXLf81m8MI0/ttgcohJTnHaUFdHPmQSUpKbBXiIW
VGTFts+KpT/YqBxREYVgquNjIHkaOohOXpwP29avgoA7NCPzKlpsOYoNA/G5jICM25KBxQ8oygRd
gSbVtyl4DLh9cmpBP6cPV1oCyGFrQ3vuFpi3FfwrBT4U4QUH2ac+V/bTDyLAedL90Ue69xD+JA5f
zzB35gf7BqdY/2oMSsCLGYpyAaHwqRHkP3TgMcWUbYiKxTO8lgw9rlsM0RruYfn01bSxv1NoPv15
bTbF7UDbVOfNCxdUUjMmUi3juanN50U63YFCKell21DL4/f7tzTWn+aepP8o6VJjrjxPffHB1P4a
atNX+7OB8StIqJp1zXbpOQxiaruzP94cEUxXkefdi6+zMGcqzklzmDP9YvidmDetFMnlK5cVo3/e
Eb9GLfqKexTGY6K1ySN+U44Y3xBL2jOxpTQYEQIQav5R/BaQNT7fsULlN4zSoJklyFiEQ++8NakS
oRWat/B2K1W722Ebz7cGgnpO44Qf0X/zlNn5yTCYYQPY9oCj1OTMOZ4FecDNH0AuLRsg83iJQhOA
IOiV8+ZjRLQjFxIYR9c9ChMvfo3griSEjbcJsNvBA/0HMx6iAdHsWv9cvE5ffKNWhFWs/XwIJw5t
km29FNxQsFY9uicZfZe+gDMwuwvWgW+DJWyCdDpLFfS112TKTpKtZDWf9KIUtILy36pPT1yU87iX
0I+JZ0lka46KFdODKCV+ICUk0nkwm5p4CPFWL8USsMZh0M4ywJiSApP7JAUyPhg1zVWnaDLui+fj
YqmFDf1sa6p2455cF9gQeWubKlsBGPXwl8SPamO8OB46NcySrfNhGCQX+XbFEjfpwi/DWYyGAxJk
5VTl1w1EsspfjREPtfhxPW81iqM0iiHtk6L0nAqRWKVOKVm4LfBmAhji/GeuYNLA3tUdkLaF2wF9
kJC9w162fmf09sy4xdosZqimBtR90qvo5AxrIgYQDw3pLqULv1n7VbINlamkODZec8zKVxROaiR7
RWjEU+SWpPSbywRgYH3/HbcyYvOq9T+b/ZRNY7Itt9bDR5w8pN2Ku7aMdFwu2GJLKFvRhAFKIFsi
SVy4qLtAAUtWkiJEXc/t2GCvTDxCnW7w6MYBSjmCEgfy4OssDvPRKKczRki3RZeZco8uUAJ6GWPQ
2NX+hXdUoK/kNmMx3rMhgJ0ZE4ZlZ5HTDYkTU4npXb5Ua4JDDRJrvuh62vNKO8yN7uPMlWG+v7yQ
75tgwzf9ze6y43yLCYHnZBlUcdY/jTCHEVfiZP/GeCCI0UV9AiCF9lHKca3v0JXjay2eeneUmUhT
nK3kPsn5RsVrKzNIw5QdlUTVtX8ek5f+GSmiygMI9jHyMPlhJdkaYjjtLPJQS/fwPAqJMQzCeXQ+
wiKVIvosKfuCha8uy7dgIwunnSKuWsjS8EJer8922KvVqxySCgguUzRPQ46Bq0ntICKSRRZXBW08
3hy9Vus7AWea7cmJLtgbH1hx3FfjoC6btPp9uztAqLMEJfWf4ILMUewZCWBeoMduxZHzpC8TixFR
/F5WEfeWdaDFLjQjMb5NOvPrfWd1cUsXowVPSCVfbC2rzRJF0ShZsE/cOU4heIgwVO33nLDmqsdD
1bmtHx+bfhiGbd60v5uhvlW91LW6jSbkBPRUmL6Hn4by8LmbILYtjzPEcXgYkLKwaj0WXhzHoKJe
wrHoKfB8g1Zkrw2Uegp8N+KD2DRqbdXL4mH8X29KsP/WsZssDVRDFSzPsAPcLB69F9RCjhKmqLc0
oTdIrgXTLpSYLy7B4tCTxdzv7bT/3DgwioggxEHyNElBO15PTP6HZ3PxnixDbSUcoiD0TVdHnzl0
1zG7/47f+dnPpODgnB4SiToZQWSks+kdCBcpY37iwfIX7uCH4owEuoG1mm66NqZ5yosK0WdsQ6+X
fJk0oFstPi4ClnTxmTlHdsmATokjAFQ62xkZZ3J4Uxn4d9jIEvShFsyN46axdhNc7fvHa6iaaS1l
zxS+LvbMc7/vNgrffYwvwp48y9DV+4HY27abeDWUnikZ+gKYrnDIDvRfwbAAK2HP9MWVyipmSjgp
fflmF1sMnRuEegLlI3oNr3YQqBToTCszJ2a7/mkOx1pQSa9Eu7EIXGrtw+5qvc/gbafUTvqNb4sU
sR6LUktPB/XsQ1u9ztUjCJ9bo7M5j/cfsClQPaU1QUD5kqgGwOYJJJynB93/ZOjS9dLrQo7b13vL
3Y9lu+WqJks8hFDIZzo0Nrqe3Z59pp7/NETETndO4ijZJR72r+8KRvfpj3Ow/jbLDqrwn90YhZPI
jXocIOi1ovie+VXHU7SI01PzHck6ebf7PmEHUap6q0k/z0jVyduJ4a80dmllw8VQwP+e7wyGh15N
xPlp8pbXvh009vHk2UjBgNnJQtq+rPyYi+A8N8i45EosdQSG8nxNVvpHLUHtUBrnBuBkOpvgxxmr
oJCjRD+FI4dGtLIdt1qgBNaNd5pggGv1ahLBvKwJw/BFDU9mKofpLwW3QygEAX6XK+h6iWwJAbCn
zQyjGwj1SgiSRa6fH7pjFec2kj3nx9q2vxsw+G2xO63A5ClGSX8XgADTXcE+c6wvIdpCObS/qQp5
5GMFMokAxumxb6bILwsWQSoQgOimhChUFWNu9RxcjRQWSEoSlOXwt+DUcgxFBPT1sg2tRG4h9eOV
lG9k8OKCcNg+CAaOLof9tTOozVBRdYcbdSNOJg44/P68N31j6usJ0TU0XHG00b/rcoRyJlyBntR/
/oUpvH5vk/6IXU1UxVHdYrvnbsU7HULAlEJeackIHZ7BacmiXzKeZwBUSgoFVtB5UmzjAghuXVQh
ksfqqdO/k6GfPtOdAfuRfhycoYsEIhhptLT6MM/TqM5n0wG7fbt94VmFyDH3dsJlU+SOf5TGfI9c
0SNcjLD/5qP03lSUhxU3bB8bTOGA4sWWBwYtyrzvl3zNarN0NZO+QxbBP9ocO3qBdnRSMhf32nqW
jgIa9q+9kyYpQ8rPJjuER8GaD57yD+K4+j7JQPeVm6WA/l9eEZU5+SPso9BqLJ8j093UaDhu7z+J
0NjhkzBDE8YFuRQDuwBil0d8TWT5Wu0BAQJ1w4cckqPrYtL17hT6+aCjsQgsoWks4NzXUea5kI1b
H8tZXJ2jjHGNly/TCVvweCb2aS5IX0ZbJ5dVUOOEeRbXJfUzjntP8NMUIQGm2LWuVxBdfvElMYl8
QE65yUSmdwMVEusY5huyZztSvvmDB04GlTFVwdwoOHpZ+281Fj9St8+FH7nOCM52QczNxs1eDCoB
yuBNqFbB9btiQmTf5v/deXKOQPTYvQW4vbooWMY4mAPoDQpLd076QUv3wJ5KZbSD2wrgf4F1goSC
SYZ7QJbOcO0dBv64ZjtmBWDCWPS6o/oKdKbBYXwx034Nti575qtjOivWbdInzCJI38QL2IRC93Zn
Qp3WwfRNCQYOOcLS6irRABJLEwVodPhD3uuWi6Ij60z9u7M9GtATq4mJW2tRLILWKn0wzKCftJVQ
dCWmkvYGTBI+Uz05+2M98SVRBO1cOW7/wNfbKiSr3w7vB/9laaQEGoY7+4Ztut9+OAwU/A+WCIzt
fv5gnBdbdESCax5GZOsE61YU4cVCOCjpKgqVdgD5eckS5aewkyaxfCPxXHbfjweVDlqhiK4q5FTR
XZyjBN4FL8oy9BVjz0j+q2SLQMyCRPVwCcw0BWwzBdl6XkHF/Qxdd3YHn1wQjp7c7iZzK3jOCxTW
ehpzQk/blQR/MehWdU3PHZV8o795O/oBylWDj2pXHvlPAg/yIBUCTGpf+ruAejBimEEhWc2C7SKR
zTrrB1UZ6+ZAOlCQEuFRQrqJlSF46xi6gt2JxFKw55Ng0t+om4Hk8Gtb5HlJQ7MCSQNxoQBXW73D
Oy7aMJUtOotGBFsRPIdsj9rSjKzzN4n5MjmdXzVAfNIQk330NEPK2+g4c7T8r8oHtL76JGWqLicQ
rd5iOVcVqzwKxdMyDN7+/pj6w7ZoyajAe161d5yAPsQrPdpdxhCSRQDe5+5zntPYTCqo+upwArOk
d42/YlrgOcaJMiG5KxmCgPCHqBYLeF0//X0Shirt7emZLRdBb6OBP2jMRlkIkoZESsaRJcj2e+I4
pUKSYJ5kKLCUTHHZ+9MZry5Yn00+Zgurq1iaZbgEVjoQWh/AmEM2mOOQP96XJoZJb2hwzpFcL+Qv
JyLtmKCKAcUlw/+QbbIlZW8WIg7pBd07+I+bb2bTh9A66Psgh+253wGgBKBEjfGM90oqfQs8dYJo
z/4sRY/s+/xNXYao0QtNFOc0tMiHNRBQLivhzcRvxu7w1J/om6Vc+iAYGoktKQ4cMZN8VeZMTjHo
3hy3iyaQUC39c6VCBA/7bAUVr5+o29kKuuJNW6q8gahcRbBuP7m4I5LYPwhvRq2HZFBm7pmmmT0V
pNX3WSR0YnRvW/V++HKJ37AHnQtbY+0aD2KTA4Ku6t9/yW8MBaXiUuEUdGKF1112cxvEz/UoyJUL
MTxFy7x+LJYrj3ByUtvBeg+q9LhCIBZOFQ41wPb+xIfXGaUN70glzgAHnmqLpiEhnCwbArGMpL1n
818FsB4hmAWVC8AgmDg6KIU6ll7FlQ+bynY7aLEMZhVI6f/y+v3g7/niTkJ0PF3say7yjc0AFT+V
eMAMukURuY64aNSHfq3hPTFOUgB1C229FqDJuD9sPxs6MrLaTJXIYgwIYCXlSEaYgs9Bz8mhwYxg
Vggh9dIqYRdVBE1JHUe8Jv0w4XfV9RENMxXZ4SniSzbCA5S2T+5sJO0+u8aBC2TTsp2PeLrIiOyn
YrRhZ/xO7zS5inQRBTM2N8ssYf3E6afZTR04RTuYgtD6minbVn3CVI+VUUNp54ls+pTP9Ul8SHxv
PQRqhhz9Hmu0wJalYtJFJDPWMg//j361i8L/IuacKoFlk7Q8URWo/Y1aoZd7kK7fwdASdjjHBoCL
sLfZZlk+8BjaVpMd1QcqlbQ2KQbXRhiDtIHrYBVC5YZuexo8SgCYVO1Z8Lfv9YR/1GrG9qMRR+WC
t6sgzeF5rIqhY7mrb6fpGDdZ6H0CEhpDH+ckdl4AR0u7A2aNo3K+nnHjDc0TVgjzfLFK+UIoVD+u
s0TxV5J6tJBY3l1clbhhev1xDk/MB3DLeNBi4ACz36M4xjKedZTsG89mvEKyQR2L2D3Yufred5+6
2qm+3z6qGZTGHrp1Kf60edbdLqSTsiwUAN07Wzm1JNrs/SEi+eFmNUmYdv1p2eorQthBf9aVZFyv
j3sNollGZby6vtjojsuIE9raaRLQ0RHn5M+2JycHDGXH0GEQK9dsPwGTqt3e5kOfqdeRK6YG4sNT
tVSuFQ8JaTBULkXqGfbUWehK6Ng00ishK5ezCHoTtDdOG0HK0YDxtrDiGMI9p3OVToeeToJdZPiY
KMAL3phkaYACwyVeTUd7e7C8KJ1RGyPcyR8gqUkCjVqZdnbboeBTl9Dp1K546+i/YlZ/fC127Xd4
hxwUhOVcYrkubn996DNzpxlFOPuu5r8XhEwFxtUxYFgIMVrpwlGHjI2S6WvlJ22FpQJLir6rvvoa
n5SGpK1RxB9c3CV412Gzm66qzHqeeUUppakImbzoJ743Qakz+j2mIaQNPg6GWpVtbbtOPNwk6axT
YetEgzVyq/H2bBzpLfYM7IPeQNBlmypeM5r4Wwv4dqfG61uFSMzB0+4sZdV2LwclslnxJQIPdkNe
3gaP+an6esqeI58VhpV7OhYbMAHT2mIJgQJtJ73KvUa8txtcpWx8v3lVcVC9MGCnzR6LT+TGEeIS
+VgvMWjPUjtL9Len4PKXudo4khWiyU+1VEsaNqrtmONVyWeEd4u4DhGRQMOF2ubsxOD6mc3Pss/k
p+8enkbTXloNC4060MqEjA1aEJ0/fRx6O+vUewj3ahfwlEOrQXRohV3zA4s1ADGTnIpWu8kaSltp
K7XRqrQEd1Rvc384VRRfW/2S/NjVHtIJ237ZuvekWqWrcH34O6Zl3o5PXivzvamo3jxY1SUMQcds
ZMxWOvpe6R/H31b5PvhHRVrZzQgV4f9isrM/QL2oh/V+C7kZ/EX1pTX520LAk3ETuJrxSyA7iKnt
0Cv6D7xZH+fQ4968Lc2CZqgJuwiTZo3BLROODq/AiiqTvzUgzeqaDRt4937ronWhKU0KK7A8lNgH
jXuWQBUjQFO7a/3zsRoA2ngYu3OhMoI7+/olxs7I+RIbVjDw8uOkJZr1/N5MbVyID2YxIaQgsz2W
FkHq8LFq7ipJV1E5Syl6Yj/LWzn8BqPV4jLQqNJTcEOxDEHP3IvGcqTpZ9pfEHkY8Yt0cNx0+yx0
0o6SehmB6gnIw4XK3FLizbjD9fsH6vwwo0UeyTy2Agv/90Vu5ub3PHNQcTZlYdFtY6WnGgMnY5/J
f6jDNT09YSHLjsp0glkzgerg27dDY5c7SpkV1E00ed5TbTKOfCNQ3O9VqiFSw07PSkBG2e7F6F0p
1xjFbIXzCGO1TB7cAvfYov1dMYu6VpzTet8llqUpQyz7TmcxQyXr7mkgLGU+Umdp65CHBfoz1hFK
FfxnT80DWz/V7WKuoGBS44rHedGhDrB6nFLR7iQd4xr163XNzkxhZeTLxsrj2OGCeS9MK73N8DxA
CrsNTzhnDL/kB7b8EZSNSVVU6+sCwoFxvoGWICjJvSseOjIw8WLP1CwjDuijYAK/rvZN6Qss2X5U
rZla4ur5PnLiYQV8DCcsXzAZIIHXfW0HYmlpgb49bbv+85j9+Xh4aGkN2tt06hSxV+OK0Pw2faVm
Vk0NwOYk70i9H1Oka5FTeBUbtfsMzzs1jMtKK1uii6osifNbkO4M4SBM6FVXbQ2Tp5x9RrScmicM
roM8ZS6yW9R84ARxw9LkN5oqED3cwHt3rPkKo+/ZUarHqkkAM8o9M6f6286FhCq0OLzlodfc7NFZ
fJ7Ki93SDFwjLHK61S95wTULu/LzgfuVP80ruBKzQLZ7TtqptwcDL9PfN0uzVizjTSXhg1DrJeTs
F95sbKvFG1BXR2V1Z9b9ektgrV9Yim1Ay1HFdKueEw0HPw91SR3DXLQPTSjqwvv5K/u2Y8fxV/kx
g7g6jJuR+3KqMZLjgRTu1Pvedvm16TKlaHWKyYUhcryy4e6g2IwoIZRRzWDW7mX+aUesJ8EZq7xg
O6pLMaDWqavKEciRKd/EYlP2p0552i7W0LOv0w1OcJJuEIXwrwzcbhxOwfy6ztypoyG7PNEAe6fo
+GocDCJMhWfZr4VjZ7wUHPwTCe0fp7YRTZmdRkIet5alM0qWC+lD5K/tJcXAtKZBzvaD0iBoXgn1
uZ2QrKkG7YVdhGVaN+xs9Ig2Yr0jtK4KIuAMmVyvFHRiZjiTn55NUzesUEEI2yMw78gtj91F7+Ie
Wyi5Naw5YsCGDuAkquXI18774xkeo/iK+8pvNTRQAbxySmyazO+BTqouYV+5Kwqfel71O25/cQTN
nAu+7rt5+0t0ZnIz+pi/OfAUj8/lDpdkSSZWH+oY01S23DUzeV+D9E1aPROHGlmadvZTjtVZErib
L+UD6vYyaHqcNu/Z05lIcexjm3PwaOtV8u5FccIr+sBLfd4aqs/Jp/qzKPxh8MIbvbmFXPwsgAU0
z5cMIzsKP3yJXtRbo43/emZvaH+emsYDDB+EHKK4gcmAbI0RVvEfRH2aUb814Q+oBAo+TUCJdLEt
86EE613MzwWxZT2yiMsUM2pDJJF5Iz0IqP0+qgII2A1fzJJaNQUK3IPrNKt6y4CANqVQ9f5NPDZk
YgzcZwTmGgfkMfiQ+AWLwPmLZjAfjlwdA5ZmQ+AO1R7kND9QWPo9yzcXPRmdscg+xJFAn05Q6K9a
H+HG9sHo0m6Xh78lnFYVTfny9sA12+mBVcTq2jt++m4gzWsoQYWqRMJ/wEOFJmYSIJgXEgQeNei0
OgULqXHAV5hi0+0cSBIZQ9PRqqKLTh9BD0b1WNGFicpf96UVNU7NVJy7cviDGhogwRvQNXfo+PgC
1zaIT2hpFJwvVYc6ZVolWHlP5fulZHQ1xT0MjJg+iyGniXtor9VgIDQrJjt5uDjKGjGROWvb5aBj
tMymggwmqdm85gtUE75yVuxiw0NlyNbbRj/xYWc2HY9GR2KLy2HXV1pP7fA9nKb/YC09mVzltf6m
cSGG7Udsj0yOjettwIXRAK7EGNCH0ZcYWDsMkk41V6F6roKJ02gTbLN+se0hJDW1HAP18+XuyxtI
Gz18T1QJuRYuMkF3OS4sB+bNmatP3cITjDwLgEZH68KNqhFF3QFaUvzc9IxQfbB/zOcQrSXDzVLa
uxA03Pmh22zSin3f88J0Roecx91/WEma6PpurkFzgPQFMpHhVC4MWhYUA/5PWUhUK9704MMex7sW
DnZ+swjaZwLF9fiMA+QycRdquSE04zcopLLR+uNm41rMz8cJfgVF65HInH2hyg6SvswuKbnD6aEy
id2bXixnKzTyOt/KBHgVVC8T9kLywaBdUoVarjK8Vq1gxN5WgIyWoWT/ppkXFbVFj6AC+OfX502X
nnUtaBLDFuE+AELhoD3Oy+dd/ijZcE9VfwHl3YqgDf9Ia4nP2wy3z3029Ytzf1loVdj1auK33HJH
Ze4CU/vf29YnEItocqG3MhYg6q7zPhJE2culnDdUf6BUFmAago8pQL+ZrUpJZbjECg0dKOtUtq+5
FSJnLc0u8qL52zGDL5lzvczl2Y3KSr5nqegFeGUJyzdeElNaxPsGGlK/AzJEgvMIBfyUpUIyp7I+
xOmohciTIPogt2PZtKSdFdLHWalgSZyFMM/fDfZefcXXeDioV6rhAqVoxXfo2FbpGgzLvOmW4iP3
4yiIUHccuGaXtwZcL5fTA2bUs+OqRm3j7FsS/93PQBP6CtFEiqqg7tDwI0qmB3PGI+LOrMYYU7yq
AV/yKwkMYWRu87PgO100NFEAUy6U4iNVP2g0oKy0bS2rnP5Ve0Em/1ZWvGfu2/vpb7MDQo+Jg/69
tbBvE2yv+FwV/PKfkOlBiW0N2sV20ZTF9Dak8AHImhz1mU2Mk9ryqsVhVrH1CUwiTflqqWZELRj4
iigDwN8MEljRp5pw1tWYbIcSda4pAnwOBEgYCpWp+p6RvaN9ii+tXIo0u23WdiOJqv9d4qPE1DjU
Hvm+xSeS09cDJE06YOXd7ZH04sgR+oXXPVC5K6+1u17KO9SV+YSqx3PseWYCF2gMiEcnLI8SY1gT
9sOa7BZzL/YHMw93JjuGroRuGqd6NUwuxmfsuXtEHYa68nID7hV9ZoKJsv8VM9y5pkIxUzoLQgGo
mlijDzWfar2KO0KE0uRw6x9k1ew4cB08nKGt5aIe4hGYhxccL1pw7f84voeH58H6hmGAzzbR8ZJh
BwgoOnly7z8e67ZXxtbuJr6HEs3pmPCh3tnPUOIMzfBETpjTi1HHyGXOVhxRDxVr107g0uO0KZZN
9ke+SuRSa3o2gchhBIbEaUDpN+mnsBRhK8aTWM1Rpzmz8UGIjhLjqSrUah1e1FCYqb7qxTBNXXkM
LsbDKeUf8kskH+nNBFp3huS89KrOP9VW0CGo3cuitJ++FGb4F1QGymudI4QcWjm6xSV2zJxv4LqL
EKm/xsviFPy4ZdYIauMxq5g/BmOzrSAjtb1KLIpw8XBbaS+2pZYPyBM3aRR8l9/9y8EMizCmhJbq
A2+DluKxi8kaTcKKvIq+GiL5OL0dXmLSAU685kLTiHGfG3cPZgTvhVjNBmfXakQ7UVK2ZCK1kuW3
nWCfQmn5tFgJ2ohLwaRH3DktJ8q0R3Ii8JW6/UyEEB1sWQQw2Ln0VG33GqLq4oeQww7FXU/h3wL3
1PuooiyWl/69+izO78trsU68KXNJyjjnaAhn1Kc+SEpiSOEJFfO+1voh1z8q/5mCoY7eZ0esT8lH
XXcrkAuVwBAE0lS0L0XRUME2Koh/vdPncSQ2aXeOVkiR6tvSw1jUEd/30B80lSkyOL+YrBTPN1Gl
ul+/kEBfLYYUwDWZIvtCvG3E2U6ZOcIft6IaEjKw2nRG3tFks0JiRP3V3lSn3gNZmAMFzOY1pF2J
sl7oYNOl7BELxZhrEvNVpjDSB0yAluaW7XygGlDim6gGqGAVKhEmHdGSN1mzt6WiSUBI1psE09Vo
2sC4bNvSBGaaDe9xsQ+mQg0Lmy1EckR9uilfrf0Rlj5cgGUf9HwBqP8Pn2W5L2YACm4xKTQItB6v
mtyI14g+D6Eb5AvFa8aYg1raLyWvC68t/o57taTBW2yZMZye62VOn3fKtW60h6j/xd4eLuO1JSak
1EGwOW+mxIrKKGezVnDIQqTg43PRfFL2uoUJ9uph3BekW2U6Z+aP5MHNUkjMkiEtq+ZCCErMCohu
fm4M8J1mvsrrAOWP5eQZqVebSasbW6I/pbyPBbYef7ZyBRQe4WOdL5iptRJYQ86Zee5aTYre5/Ld
e5rAgz8wDqB42rjbj4mNTOnF8aOkOMh7XobyMVaN2L+/7r8cPBRw7ifKa9k5x3bJaHXFUXJ3oBuV
YCcEQtChsLB3/KxqqjhfVAzTXPGO34VMUiqibf+dRDxO8BBRVqwpCdVNRURB9AOYbPSQeY2TtD83
z095PbaEaYQryTtocntD3WIW31v3eJ+9VlnhoJOCYszTpdzJ1p7lk097xUZtD30+5kujKbCUZknj
Her8JZy2Ots8FRC/rR2048XR1tqbMe3kzLVxn6/FIfqPPHvPsHxJbAfcSk1CewtPApkymXwQxYZy
YRHfBCOFOWUYWW/iEvqSF22I0DR2atlVF/xl3cMF1EcXwZXJBFAUqv5jvTAce6uThPilONNHYDka
VcfmX7FBlTJ2BBmZ40XcvN2d+ntU8LhjchZynieyPG+9o00Rbqac2+rrvhhqoF5LAlJrEJAX9Os4
Q0JZ9oB1xZijoPvYZCD0bQcABemdWcOwewE4pV2vh9u1aG2CMrLx/RR3nSWu99HvAkirqPXw4S8e
NiqnEMTmEcGUQ+0T0xXoPnGnjtCk67khGsM24qx6x9LV0vRS2bYUolO5nFMnA//hAg/DtL+vL3sq
q5Dnwm6PqH0XLoYecb/UUyzeefl8AGbQy3ETD92zEysVXTSmeUMRjr09aKS8OKvLrF3s3OMUBSyS
PRiya8L5sRibT1tFVgBGUAb9g4XQQ1f0DykRgJV5WEHmZMVttu3q6gI1f1dUBJ1Lvqk7f219Tkes
zwcWfFhwhkBwKgWCFuN0f7gzqHeCfz7ucCD1GkccLQ30PcNFz7Fx3xqYkXwn72EUlQPBgW/vJZaW
hBM3jC407XfSfk0tKrIQlgXmTyqlAX12s9QQFuvyODard9GsN/x8qPGQ/w7XPVLwu1RlZ2mjlyLj
Qc4lFU+1qYvKhHAo07O04fdTifUb950ZQx6ABJ/1sxhRM2zBWc8ypd6TvPThaBAHXyx89/db92QM
w1gKMNLC20nWQhx3VtdAvN32GTfyQizI+Ec7vmwhnVl9QjOwr710uVbc/gLeOGAvMWLlRJrb1U9C
hlEA5A6zT5/sNbv8SeVHuhA40gjkJv5rUmXbNRxtseYZie/d2JWRoDibYP8dsu87NCYlDLCUnWmn
5ANcSU38Fecdk5RO5snbxGUa2pJfi5yVzilAwwkJdJONYRjcZ6+pBG0t6klEcpl5vlxi8u+fbobJ
CUTYXC7OMX3qrRVwTcoWeUfxQyX5goh4B42bQe9R1po1JngOgTNCbbLJi/4e+MABOWndeOl6SrPp
GEyBaGurAqEPA+rnWglSopztHLGNAr9zwTQUuJEx8NEGJUOpNehGJXaUEkx1Ra35770afLGbmlIs
uI4X1KUWWzTDEzFw2OlDNwYyX1Uyx6TxDxbLl28QoXuDgkkRnS4WAA+/UKlKma9KQr4VD9ucT/mh
O+rsDx3zyVoiaNK9P58+VpLrZ/UzwF582qpGunMkH3EHIDsAf3MwRr9pzcoxFbhIK7rJRpAxDY0G
I5LKmpeksCTlbZtisrx/bB8F8chbepQ4FMPh/1DZ46iKMGIQJLp8HJdYxkOrWLwA4RAylMurxPx/
9BhinxRcyRTJR4VB0JPOAOErG5EtSPcmsHKZ1FKGNsCwFogsKLEd0SRApr2wSzEOww5kU3j1INWY
op7v5fMuSbRdOQhsY4ANvXzsLx9V2C/tetCpp7vmWrHKy+kHzKemNPvTdhqzhIv75jYxlilsTrP/
ontdO/CFu6EKlPzx2KZ5GYYrDVimdRf6w6v5UNOr9cXPtnZza+Ym4A+gWBY+PxIgPBLIz4D0/o1g
YRMMya1AuegLGF3PqSuc6gxrQDwGXPdCU66LJv5VTV6P0HMkPZi8k8CNUHthk+8jc4U1r8sX/jwR
028mmQzzEhyQpEaeugy7SN6f0r1D1sGSF+cDkYZTEzp1i6vRx8d0iVPlhCwGgDEGLUio57pk6e+S
VdTyAR5HjT4YospR8aklzjY7MJ06Tm3a7q+dC8SyhgcUeiYsi1LjiHc3zoyX5Uzrdl9HHJZDeMi8
190kXu1D5KA9tHqJBEo9S1CYT/VWUowxXoNiVSMgvdeZNw8n2bxjkGbAE+fWaRsTWX2DGD9qDyjf
UDMA9723fpCUHTZCqxmlX9TCwBaVpWo2UVj3WH9RJ+Gg+pRG4o0hBEtYkWqmvtBxaoqfyWa4QSvM
q2noE9h0aivuDBexqqZ/P9bR6bmHw1DflxI+su/d6FOXqx5f4nXOOGLyrRLMX+y6eajYJ96+DdvP
tOahPoUNUk/Dh474cPO51aKMVELYs70rGNL4rm1jM3WuRmzkAtjh1dCMCH98EErgDujhxL2LqFXJ
tBf7IjKwiIYBD417Cph+nPWlifcwH10AxjxRmus5slx8DP0Q4yibP36/pbIJ0MSGfWJXWLJQOsaM
we+xf2ZfRkaKQRAVB7s7rQpDAFEzDpCBH7/lHiKw2w1MhzlOn9XQTZYWN5o8zYl/7tM8ObBiqvsx
mwR5h4Qk4QU43elGXpCJdGdrRQmq4mmu8/BBPaKi/lO1dl0wl/TaCkGRBXDxQkU2RD3pMYamfxN5
PklUHbQtc1qba4K6Qj4Wbi4jf+oT3XPsThAc1D4GaeXUkT7vVHPOmap+d70wS1nNw/yioumrTcrh
Et3gE+NKnAPnULt4kQKEs63OB8fCpZDH1XofkZco+U+4i3ZnRdP5w8ClI5cQ5g5VCFXkvgyKimA+
U6WD5Pg3Z+/f+ezsRzY8qBPf4OieebiLht6m6PzVr0DJnJDV5Kp9yKgWEJQAVAQohy4FHAKNuo0P
fdv7QoPh3+IujtWMbbAC6oW19zi8mpbC3UQ/hPNckzqCKOJMKwF3F2jQv0l/KlS0kZBesv3GyFgu
i1+r8V/0D1+D0x9c1JlPXHpiC4lJIClEKXphJpd3I3d95VpK5S9oMP6jQa8X84AF06gKLMcgcK8P
QDD6mJL4xqPDZRKJdF46tXXyIzmMDHaN48P6VyRvbXwa2w71t0IN7wXFDQEXe8wbN3GqIGL0c6nz
waBngbFIUlDOymULUnCREekmFSDBVZPLe7Drru1Duy39mvE+ZU6OMxffyI27lEVMABtfhdOAC8o4
SVIhdYf7B6uv2jwoVBFN59X6fd66nF9wGTXfNIq/272PInP7desehrLiHgHX+tA/Oopx51V3+Fsk
lEq+YsVMPAoE2G9dqtc559jdYJAKiiXIZuMWYejxkEecxN7THHwMiBUSXGVHWZa9yeLAmnVp7pLn
caFtbe0mCWRxDAuHAGHYYd8X/waD6TpSywG2Cis9mgYEmgP/h34mWHQJtOOHNPkTYtqTMzJ+i28O
bodMvFd3MtYXt1hMUvgP2H7XJenCB4jr36AEtlBBmz+V66gm1qvyCp6BZeemTzzD/O6lLqjwOb+5
WHPTizHMD6f/fQiHpc4kbYIQrKbWunhiWzXzeAVaP5etV6OCf7+1eJFWXGLAJRZnTmk+NWM+SWx/
f8MLRuGZK3O0Pqo940xhxFYdGLtiOK+Vy65VGyZdaUHl+OIj/mxKNcwPvzThqWYeHISAFxzftUOt
7c3HSs1R3/zDxfYnArtCa/WYBPx6VSr9Ry4V4qBrCyqU6/xmoFvan0Nhgf1+F98rdAsNCkce6rPY
3rGQc1Zsb/sFq6wyhbRg09nxK9JGyXKcW7IxyMdlEe6lwFxzqA9qWPEYSbHqsKBikFFyDY1kLI1l
inBK6H2/eb5wK7ClXkA2GCAxcZZJvCbCFMCBCBl/wn++YJRWEAWFfNTHJHvixS6JhkCAl99yUXdi
Ah1aqA+EcHBE/vetcjIeLoK/8pJa/6dIR25Zd9I6DzO7SYBu2m/C6yOk89mPaQIe6REsaG1lgi1X
bieV8iRq6EOJqN1hxbJR/cPbGDR4bgf6n1yhUpAI+nNzZEgKdkLmQi7TQWWLInHEgcJaXnOjIJHa
DoGlWcdBwDk1LyQwyOzb09TOup57pC1auuNm3gRST1UgVdKKyXraG1F7A7P75XhFAPEbdTTaFhVC
gbvkuNie8Xnj7cDyvfGWelgdXvl3k1suENNuX7YcZZp8I52dbPYFuxtbLSisc0Ix7G384eLqFuFo
if8u2XtzHzzmOu0xrXHhT4OhY57KmH+zDiEGGawcG78PobLZBlp95V/j2Hv7Of6gUqlBOyf8KBcq
pBeEEvoSPPo7wz5XYsUOd/yd5NElc/f6+ETCQUHqnlQ2eaUhG0UicIpW6qovb9fY7JbMbifuVYZA
uQr24v4Ys8sFG0VB9W3nejzdWTfkBy1B/53ZUDbsw4ffiNa4drIb2du3uA3QPAh4WJir+M2wmSVR
SkqSBVIVGqltwoO96E4bA8pqMAiMEEFE+Sr/qGmwNcsZf6qJUs2xvhicvkkdT0PsuQl05pXjKdMt
bgpx1kZVnsRlYJpnUrc8KBq5eFbJkYIBrGfypQR1kieCPtFG+2MHS/8ai7zHmorFC3cFjFQqVOoU
7VMsccCMO86DOdvYqBSA6IMiJd2ZtIYF6Qk688Xb8TKEwMfmbSTcyTI3boyV6kKc6bvZcU9DgM8E
Vm5wkcj7Ack7RJXHiT+ZvLZ4Gqrv7bK0NspbBQK58V7nmqHbibgskdS2eReiBIF9mw8hZTLt4CB/
YN+DsCT+A3WFnVJBBjLcp8kf72FIuJjuow8zurc0922lbfX5SY513GdmVyMridPE7w0i23jgqXWE
xJZANzz/txJ69rW4qDf+prpwolS6qMoD81YGnMmBBL/pwcMR15UJGymPOthwqCuEzCpJJTXYEFkD
2lJj7+vNcxE7G3Ezsw8zMrXmG8p6KfntTlQ75iQXvlam2BQ3BZIPCOWOO32fv1Bxz/FV2bAl2LYy
K0t+XqaQNCPhbCfrv9jZToeDphYY0ZSJLhaB0CAWQzmdkxT5LU8TAcTiRIxrwOZH6EQi5Actk6C6
l7sDQhjqc+YAElX/coGHS0WStqSmhHbjpfuIKDb88XZnG0ClMRolrapXhJDs3xrP1i62mDLJNq0s
mZMTp8Veo4Zhs90StH1ylXETXGCd5UhsO5ft/c4dM6U9gKfIX7Ner3nMKIykcSSv/fWJ8tG3oiPz
ucAnXfTI27Ie7fGOJDitC+rbhdSPHSiVxNVyAf63BsmQvP0yc6nHL9DHmKkb2ovhqmTANF/hG2qL
8u7ptvmfbe63ws2cVtWQ/pwEGixlmo8zPktBBx/jHxnk1DAFdFRaB0RbP4PkC3umICr1SssP2Gyj
Bz/lOqLQYQYPJD9YFcPkUKSPmnoX8aAu68yH3zN1BCv4k13iVHgh4QwqIiaOrOjhji71fBL9nggq
rJtkgaWhizJKv7BBJUv5qXkZx8r+ZQZs0SDPhd15PDsZYgYPtX6Kg8HCIJogcZKjSiXFVHVhxCEI
VUsLVAGdujbCXRGtDt1RQXn9G1NZd8NwTB9FA3kFTDyrpXlWSoxsO3I4k6LyG7h5N2jC4cehhmFm
kL+PvPmplmd/ZtfhKZtz6RXlqp63CynJ6xqD/Rt7cYDhWmHAKg1j+UHPqGwyzvWOuD9Fb9iAO6d4
WIfedEUOqoF5u6ccPneXXy+on0pZXS/UNBz/Z6tD/d7Hs9A8s33FfiGSPwvsy+hvO1CfSFF7tha1
O8EYN5h7kC/YpN65xrA33ez0L6D7GMw28Mndu+fz5f4Jy7eBQbYXgHOB6fQp7w28+VbHvqzAXdGt
UGuZKiwpa/L2GAzdtsv/cV3nJT2X4AKM7MVTw56ssVkSW7Q8dZg3taCKGlGo0/VHohvMBhS6zlU7
yppcH3uiBHjyQYcHt5tTiWRP9HnZdRMApFY9i7MDWzUbgQAom0sbPLbX4xqwI1Z5EnXFHNi8nAcj
/GWSD4B+ysbVY+QOG3gurdHPvKLNseu7KFMkStxOBz/jC1x3Kg3B7uher6Vp5BI4FQXLC+KhOeob
+/t7HQv2Yle+kBnqQAyuT7MchDp1209bQvG5nut5b7qAEGRVasRdoo7vMUkGWPyPwTqyUL0mjtK5
aNTyrrBXBdNr+csevh4uh6de9UNsFbA9ZXPSJytvLJREvpD7POzG38hEE9A/lVMwMHWZAK8zFqC8
qAFNR5HHxCySSZQuMvHEhJv14n/4YmFi0O8SLIAe8PomWW42+S25cT2Ql6lrgn6UzdMXTSA697Ak
eNzKE60VCtPMZe3LYT0RVQmHYThh9j6DoyQnj4O9cAOBH6OmcXufPxS90od6+4Zyz1MmJ662TLvU
fGbfma+SiAWNMicZCWMpqqan4IeY0Lfa6SM/qtMpVAQyGyjPcvZLsXa97iK5Xef6bf6BcQuwvHOj
hkWVtjb2JT8Tz/842PU5e1jz6xLlAF7+IPiyuPJ06R5BZfU4tV+C7NN9lISeT5MyG2n2v/Buj/Rk
wfEsdhV/L6GExr5HTnkPMGab3D7zdfQfPXmwXmfd7JaQiWqyllR0ELj0xE0+Qun3iS+oFxqSXgX6
9OBnHvQob03/zefcvrDJQFE4g26CMCDsnjmteq91hv+rS+SvWWKDvl0BzMYCJdBOrOB9I1f4ramv
dkD0fmE4CqG2mLJfk+1CEoFj4PJ+W8RUc4QwOjraos2VEUv15Dys9udCQ7LZZ/CCiMg8Qtl8ejQ1
TKIFw05E3cLWk6IIo758zqrjh7EtyztZE6cfAmgY9J4qKXLg7ukQEJyWHBfqjqeinMPhYd6XGf7B
lrxk1VbG6di5RmLR8SwL1zRnvMUsybh12tEFre0/XUy3MEAHByRtsCJfNinCruWJ+09ZRFUAEh/V
x8OlYkud1uZZVotCLsc2kaWmhRwtaoEXxDLwMjwmiiXJ7Hro8drUVQfrZly5Nqz+li3XpeOyCRQq
zxfp0axHt9hBUcdZ5+WdWthhSGGaz+r2gYz8Q+1fBEII0YPGchEhT2qq6hldrzH9byXcSbxraYXf
mKlC1b74yfFi9OG16jCOoIPeYOcb7Xle0nO9jfAXUo6RJi85ssD1i8hbXVdAEGV+UUxpZz4oSTcO
2DZ/kqcehwp7bWy/KV58VXNs94ywU6q3OnOjwN2YwEEdk1ol9ZoMeUYefis+eoBkEHaej+v9CdCr
VDYn1ElnSxMaBRKHPOmqnACIVsx5qufRSH2Y6qYls7yCegOvYqe20Sd1LNthHYqQKIbD7e1V4dmf
TpZy2wsMv8uE+byBoTN9raVebJMGIJ1F+2QYst0d2vT0INMgRcm4uLZsBjmTuV27O1/vpmwcBOQ4
3WDY/Dc5IXLQHIYa14UYdPQafLWlwQwO6R3rJGMjyPozP8fQIyECH5IUmOH3dstwIxM6K7mrUpyB
om3CoW1HOv/sH06lmYKN4tCOsXJu+U6ecMxEqMQjrtQrdj2Y1+55gKzs/4f8sOkF7w8y3gmjpqM7
D7dUVp+97jQaZ4XzEykdkRM0m8q5ksi+CaHu68kgBLXyvmQNgayTOYJRxZCHgm7u50eJi5XSBzRz
JTLjwyMNkkGtFgKlq0eMu+3RgvBV1/mkduwMIs0uvifVSa3yX0Uy/nGyUPx3FvgX4CS7vptzFIWW
UOu0SAz1YzI9BCI/tHrXNkRf2SMyYr9Iz2BGxeyHYjBKJS1BYYofR0HgNp2BX1C/5IcaUiVFhMuU
5foXhN9j0qf2llYXQTYGc5teibsdhkWbTvDLdPQwUwQ3IjLFTSTMa2Vyadv2oJ/WP+invbO8keZY
MHaizA4QMOYOw+AvM/hUmP7kdlQCj0ymsn0aEvPtSMlbCHUShLF9+QyOVZ7NInSEyh/+c74goCx9
Zq3xbFu7m4/gEPRrDvc9mUwsz2gH3jU1GnZ5kcWaTu7rF9ToStr9YZ+lU6nkhXbmU53DS7uXgds1
5jhGdJE1xUVwauD4cpQFOJrkcJeo2o2kwhsjqVQ6X1+pUSHWFAsDY/TnLCgU20s8gX+p/q80WuMf
kVGmfmOPVG8f9Ids2dcU3RkwVUtBtMdZVwM1q6BtNMTLRHPI/GZHc93rHyFpzNztYysjWTMfrOi/
ZIAx5Wpjb1mQsWvAwT2uvOZOxh+PDD702q8l7Nd2mrmcTaSg/gBSV8oMG7NVlUdWbyHilXehX82Z
2s4XHawN6CQXRWXDH/ml1wNHD64KF4yGKvpLn1g/7glkHoGn71kKwx5Lbdst6a9+Bt95UN4xBJEx
Txny8V9vLPfJpss4MM9CZTUBa3ucxiVo0ep6Nyi+OGjiL9LUuHSfJn/yTmHzQn/D11UYhjDMtJmX
3ZfRjbUXmoQ/7A9N0m74pDypSSinIVOFVcqdk7xhlk513ooKtSTZJSCo0fFPsZayhnU0YYU7uCuJ
qMNpReh6xzj0QRvXXeDAl1s3J2nwrk3UxHV26VfksdmVAZdX7YZUKCOB1MHpds0V7Ack18Rf6/ME
bP0b1NqpKLwDRteFlsqwM4DFL0/7Tr/tDtELsxJYe1++l0haJCLNDqGVDE4Q9t5oqXQqz3sQPJ2v
gAwpN8bYBiCuzywTnWrvAnrwAjAvBNLBzIh6St0TmjCc1Wj53Oo6K+YiZiFffLfhBV14NBmmVMCJ
4tYJ3AZ9unDTljUiY2VYZh+qxijcqJdDouFzER0YE6aKk63sBxBhBeyREFdcqgad2IyAqnKCp6oJ
ZHcv5h7eSQzkhUIUL7a46t01oJVoDBHaclkv6O7JgR342xWtgwAsN+401Kjr7jMkUJbHsyaNGigN
u/Kx7OmDW5+IjxEC/x1N8AKaMmLWnBrnAhQNgt2xwguwZo0fCiT2+pBe668QS9Ih0t147PnzUSeq
cp7zrMprfVeyURF/1Uq81BNCJQgfTXrL8v9JPi40XqVgEYlsyGZmwPNyv/veS5soVzli+4FjLbi8
5g+tOFXrfUWYwlIv8hqOro1Srnry230pat7PPKAltdxQik3EIr0fKltdbin/E5aJIz2zV6LfcDFT
7oW18HbUV8TBkhPSfuEdMMsuOp3XscTiKmOe0KS34H26LM+Z/CtmvnxgJ75BDfWEWcRj40ftS880
6VLPlRK78IaOMkug9ULWvtuv6uitOnZaQe3oO/jZNbaQl35l5nbiWXF92J1xdZpHqAL4krwo0ejj
TsSzNrL1R7RewX8I4gy22Aee4Xo1QdVpfeNN7rrgGMlIWDTmK74BPW2u/GVNDE8jUESjMDp/cWAm
RYNYvei/2NRqYldjG3dm5sdds6t8AasDN3pq0YP9cLxcJljkEeFhTUG2KBPJnKe52I+I3rfabOMy
9jlzc+wRCjj3Tt9G8w488PK/XcyE4VXKV2QXXbo9ertdvpOvuwR1joZkJ32GUTpXW5XYNBV7S4AU
bGboj/RmVOFz9Mf1yDQt8A55KzwIEufvyKyOt1nt2uvsx9buTV09aecDrnCTujbpaHtPjIx1UUd5
R5KIsg5EcxhPURAz+rdhrF4ouZ0VvdEFkAHtw+rcpNFgt+ZhUF0CExEsmIqF0BbD8Oq/iRPNUSHf
+CuRTf7o8PMDOYhI1vgTAhePmkMLLp3J0ToXJWpqFNVYzJOUVqwIrWYM2s4qFnw2CqudJ+AWQhvw
M3YR0Ofr0df7GbFyjopibrnwR0vaSCJ0i+QIbZ/XWUEbw/2QZrTnP48Ofe5FqoVKGW14HaR07tOl
z7W8qBPu1Gc93jpq+QwNJ9PeSJdvO1a/rqBxgBGNYNCPnCnqBNp6qB7WBLyYUsLukaglll8SRS/4
9cHZoyO7fp0JevgNHTfhzPq8RSlSQbqoLQfIhVs+eXvSVE1PL9N1KlzNShWkrQMAsH9EMxAPH4Ry
rBUICBzhNBGC0gLZqqWWM56q6KUMYDHnFbvnUkpottvZ5niQJt8sPNb/oCINGYVuQG3zVFhHK+lG
ptZJIYqe9BRVpGTkyD/PY7bfMrqAPGi7ygpg5+F6v3NB7k8jK1iVF/X3aEPM98e8PGJBzJD8UiHp
/g2FqdG40zwboS6GVYTx5h+O3krHWKaUmj2lGW+h6q4N/yhJvVOLSlKJDvtB2O8rOA5lT+N/IzEN
ENxg+2o8TVxbqr1Jc498HWjeAzu/rFZ9w1oa90zi2jy246nHlwCRq35lPm2auK0L1AhbYuAZ3+0t
97rl/aVLMn2JkYoINSNQXzIeKue7do3KeuOm9I0KxGh3YFxIqBtTpNYWyMVzYCpBbcNGc/WmsnA5
dL3OU1jcUKQJe6RrmDvOJamQ63H/DpO7nPAtDRE61PriMGrOwnpG0Z140vLSAfYj8hlLYeDt3zrS
rgBN1X8WqWUoX5t9g8RrelD2eVP+Epkkedjx0vcMMhbEdTNVPgh9ezNhkR8VVLRRyQUyDyUQcopB
QXlVBsL+Te0UKyqB4mdbay2LbgQtVh/SUponyf/TFsj2V56S8fKmb+QuqM4GRoSLNcN3UwM8Cff3
J0SfECUehDE77ed6eduS7KzZFdtJiDWlYz2aiefMpQ0cg0aKJ2nCG/oxyXoQK4Ym81I65sZqdvDO
91pdRSMi9FaG6L8lK8h9it/FMS5Y08JIj1UR7QPchdixu4QmUOoLvy5x7Rb3cWJHcSV+T4XczanN
DbWialhlNuKDMi9HHEz8K/6Ljc2UtWRSX4zuEcHVgDGvCRvWUQg4ULnnH6cofV6CtgmW1QMJy6Ux
jS0SyHs2+dlwqPZX9DXx1noU9TEIueJifKmXCAvIF4drrAvajKmE8sGMtOSlEqdZTpEVqjQY/kV2
Y+NK2dyfsuPmkvbmHvqNBIAs4sP9GOHitAt7/s48dGPjwZOxPYo1edz/vtOArYxSYlnhjAzr9pnc
mLQ0s5iCMoywbnuyDNAIk/Qtx+mtb2yvkrzbgy0aiYIxREXYiQx5e/1zABiQEIaYBw0yVQnVK/CD
yurhz1BZ0g3RZ++5S6jLcien6C2uN0ROU8KgAPgdxDp/UqdLg206tdeEK9EloArDVxSebjwTv6o/
abmS/syNHe7yA7pYwcLIyRflEEA9VljFHEMwG91/bUrbqJ3UTW+OwoZnut72GKzUaERrj1ESxQNr
T8rGY87tApnY105BRbMxV4YHhmyrx9x0lveT9X2lqT72bJsSeLiwRKDrZ1Pr7ee+GArWpsLF137B
1PwuvA3sS5JfcBeomRA63K79G4+K/JnolbVMlwrE6udhZ7EXVngqyuhXTRFIq0Foh+0slocPk0kF
Ex0YLDgg7rYkYkBmc2ELm/jA+CCCcH4gYVIaK8gcpXE3/xxEwyB7XIWZKA8755e6uwBoV6C8/JDa
dxS1hmEg0WgJ/LCw9ANtZps2l/U7VpyJXv0s91lvOfo40aXUTIlTlVdEs01WmdG7bWc3w1YfmxB8
4jxUC67tXzN6bUrlGAAb0sXKlKMCsDu/UmRzTNWahs/UsPSgqFuHA37iuZ8F3GUf6CaTfmZy3FHJ
gx15zOlQEFAsvNyNtMRBJ1V9kaH5UInOidVuZbd+sZF3u59nCJT22k9rbmsLqXyRHAu2x6a4elrG
CDhp9upVLD5Fmjn5w89z0svq0aZwQ2DOKrQ8F9+d1U5EQ3hMeVBtaRt+LMR6R0t5KUvOKjPs2RL0
osBtHxgOlD9lpIjXWHDSK/jGoMYJ64QT+0R5HOE+G8pmeUDTnm6zkPKb79/RZtdqV2bCtoPC3G45
tT6WaMtWikY0jr9vI3arUqWlaDW38NW6eIoI+JWlgk/Au63kyQfFJxRsLnBbFMrblRfAuV54l9IN
KsJOsgsg/WPe0vqNV5LMIk2euEpKk8XRjSrmDuRR7diOfbyOKjPi1AHXj+tKBytyyEFWeesc92WY
2QeBeC/HozCGpAya54S6PtTVvjR0fC0LMHEYlcFVCNg/1yhkgn+UZ8KNx0BlyQOiBJxrKmi2JAa+
G3LRLd8LWRDL6PKBnQFPRUp6ZJEPXxd3SbdTp5O2ghsgLFPm2eiw4t5A28pUuYtcn9mYBvrylSb9
4IMm8K37b/gxGcRzcufKti4zXqMCCcnF83jt++lRJgAQTRGAjuA7TkxZfrzOWUHhUSFDJk+K8HJY
6R+a6ZM3Vimyw3ulPrkyNL3GNlmnRkSqeqbywdyrLfWdfwaVMT9kcywTEVuEwmCDR/4F909rOmBb
APVP+z7F+JJ7AYGo+MKsPxwKhxNBzAKpNr3TWIFRSnbN6ht9a38UmGe3zlxWy8UuJMttqoG1cG6r
ZVMcfLkPuL0f1wFbK6kXD5p//8gHYloIbpP2LTz2zHoFVT1ma1lpA5CzzRJ9Ia1HlwbIBNCtFIwd
OeoQ/xRLZVEjihQJi9awl+rJ136EdY1PuBPgsOl3Lo+j8ps1s+A9l45U+CwazgJteRbn9qLCAny9
QhjJW1ZAwjgV8dQaxH/nLGyWCLZhgpaz9rWUUZVSoCABb7NMsFKiEkHqCw4KOw8EzUGzgofg8AZt
rMtvEgWQhx8k8hdTw49u+sLvsKjVxI3ktW/8aC2oC3E1WLjSltasZxReXkGiP7IOzLIDDE9k2qya
R1hOY54T5UXtVwhab5Biygh6+IMBTNLt15VBM7XqMcwxFuuQVk/nL0tvL6Q6bL7VnNkhDDa5GSVQ
G3oeOyCqKD65BDK14F3ajmzVVp9kUj+YsdEYQ03LJtRig+dHvqGR9XcyYX1kSr55reEcNd2k5MIu
mFsqRBHQP+vYVqu3WRzxPevrYt15GpEMQdDsRBOgBIk6IsAXvkpCsn4w/1E7Rpk7ob3vPh50sOea
hKRDdHs1mAOJYytcjKCxpr+JrVybVuoBfH+g/RAAFYhLQWZWB3lCjjJaWeWJ4fgdW0Nj1FCT3fdY
qMa8Giayj42zIy7PiL5l9ntGoeIqLBL8lu05a3Uq14ub4OTqMsb6gu3K0HyVMjqkb2Qcj7juFp3h
2Y8G+dsKZmbugLJ4DtJyIZ7rTbU/hxhmXlGUf9iwWyTdhrJtYAA+SGIb5EaoAhB2slV7uHUeRKXD
aSQxFtWPyX2zym1DaRaXDybhhRFtnCijdgfQt5rGntYzNlS78dsKLwwh2srgHkmNbP6pYRRsNUBM
DRdQtIfNVmdIQLb2duKv30ka/2d6aejNG43UN8+YFZavtnp8+4zSAT1LrieJjv2z4dgx4s6cMUfS
Lht43GFIupK1s7koTDMZ6neNZ22wd8WnUNZ2icwxhp9UbwE0UuhOMRApiW3zQCVOYzWvL6+DCPnX
4mQ5mMJ3uw0y3pTy9HWG9dxubD+cJeutIuKyx9XmtCK/wwGEeT6ohAYAqPT5dHjAmDsGMKEUrMdG
E+bOEgD+1uNja6ESZG6RGmJj2eu9edE7GWKIZFOxMvucsdnvr+WOOZtsOZxZr4+eLJZCzq0T3Wwt
E+a6Q98PzRmPX/m+dcBz+hVTWPWGwTBPfhM4EEoWq3ZCSC5UBbORlZdPQWuSGLeNkJzwjVkBLACs
yGIRK63KdF61GtaQxiFSeQzfzmCWhto2kXUSTFjx1T8NWbroShrXKoWidGIdlL2SYsDQ6+Y9R7i9
XujKCY2bAobiHQ6tSH+xwUzo+Botmk/N3RYxdkT0WPh1srYp3VZd4F12AVuvbYxJ8hXgjBsFuzr1
genrZvTAz+eehyEwcyLkhh6k6rPtPnuw3fQsor1X7RK948S2RvGn/2xxNUXLhPo1NJyNzRdbmn3C
k5l/WvDfX/pqn9opWWmzmXMbuy6dxMZGy0X1YP/yKZhZWu4tHMa8Eue+6N90BH4qlppSboIBYAgd
YM479R7oy37oKPbz0WFwnwa0YiwGRmoU0ML6saSw+rfI3smWaUjQVsd3M97nLS94D+c+O4zV6Nlj
uO8FHJiT+dQak1JC3fOTCRHraaFm2N9l/H4kqy+tBtHBX38blkVnQTyO6/UJkujhRznKgZ6eFkrT
4vUGa8XfWAgnQuoyNXUTYZvq7F++YeSkrzwQYMQGVQFHFlA31mdb7BEL24RYVPrN4cAfVlLbt8Zi
w32hu9anbV15gOrPMXUQSUEqgRpJd0/NDAAvBEXQI2rZRwPkXrGWw4gg/kVhAyeqEhqJ+COJlR6h
xCfELtVvHA1xFXCECK/xqxSG0e1rvgezHQ18wdc51BErWz21ztH6vLb2+7ijnuNySnQ5AiuaBy8b
3Ebq63oDJOmqFU1wcc928WluRjY8wKJGXwgqeyMyQOBOf0IlFIK4KamVwA/cuhokcZM0zx1kdJjS
CEgoVkG8ZAUQCCtFl6NE37IuAphtNjZWlScig7BfFF4D/KZr4G1tFbKwpAI9zwPrKjhjHUMeFFSU
RceKhPs624zNaSosB6oFaMYz9kuspN8nE4iU2JbCFkeoiJ7b6tA+7o888MKC4MJ3yBT5g2ZnzY/7
LwcGBrktdzgyzjfrAswitKqHxVbbxrnLiVZ9aNZIc5H5vuW/3cuN3wM3nyhQljuy5QiMDTK7jtgu
g02ShwEebb1WxrZlFCN/tlSAH6uWm0x68cQEsFvNrsCZ61etL21OcHcz2ucC0a20JvQpQb4vR+/i
5su2DmD4pbZ1FFPkEAzmUDiEgmKTksfms7kzW7u9UicaEEf3HSwDWjWl8xIapHRLz4mNiVc+ufDu
RqoNP2g+tu590RsPEyvC7RQLhB7cZb/Lm/2cW6LNynGxgnef+lY19jEbqU6jc4sculBemTWb8lQg
y+Ho6eFopu1Kpvn1ij6eNGpBZC9+EMFzn0QYOTkjFKwkOJaUt/uVxwUVo75HtDuH+//lJ7pd2rKF
EiCflVGu/flGkkJUZeIdPbO7lZM+HuBBopdr6S4uBCkOy49v7pReiVidS/HZy6Cw9iTEAncFwXw8
qYyYSxRM1fmuuN1S/m0+b47JkQW3K6XQurX1ayuzUdZA5MxtuBTLQQQDnJ8/jVvHykieD+SPgRv6
fu2pRt3/UophdUcM9N4UuDeTsFz6IIiou2Zt4UXsaSY5HCWLXZE5noFkPSEMHwiklX/etODVO1Ju
O/rjb6vJ1KROPpVeZlxyRJkpkH4wqsxwC6et4wgEXLM0Gnwte4iPo3hE/BcVfNUob8NHIje4qWhN
jJCEU3qK8Nvvp8kLLgnEz86b1lBYSZ8yOujDCxxQwvHyrfjIfLd/wsNqYDPoDyKjLaEgart+p6aq
8rSFWepXynfcmCfbNL9Ws5VbIQwShOy3VniBUobRoYhyHhzXnzodhs5W3YF7L3+iVpbFwJbxaklR
HmN3Z3cvPtoMzr7TI32lHI8JUZQUcRPC893yYqh72+QpfJy/p5f2D/Vj0p/JjDZ6mdut33zdbLo+
C7+ldIjuD8NYrevaMwCZwhiaAVIAhI1zU6rQ+yg4/YncxaiV1iFJWWPxdss61gyuPUn6Ld25NCsN
Tg90ATg4zLxtNB9CU7MUi0uAw2CK8fH7SkxUR6A9qrXOcu20GjfofuKt2ICDJrfzqkf6bk77oQZ/
d+yHrRM7AtZc0xHpJN5i3oQJv3nk9/1+B1WNPAjWMhjO+8PSUmlmEyUIBp4iajg0CfnzmcfVjtKn
oX44s6nKBLxZm0iQV86n+TcP/QA8pBX/5oNAuwUY6T6z6xGUxzJbVpA07YnI4hL7o87YXrS0B8DK
T7VUrelJ0phvUCL8fFQk1rUdEC7SHakKlLMY520SmXFlaUf7yxHL7JEBPUhCktQmW1tSWgFZE660
JK5QRxhxKAba1roxVGZBeHBJecoiqUCnVQlDdgE4PwzkgtYnCY4lDUKi95IAreUZFqNPkwi/hr0D
olFLFjRiMGjAk7eY3TbyXckxzi2lR7QTcGKQhpKbf+NSr13QgJgu9KJTGkEKRSyhIRvnqJGqLvq4
dmy9OrP9qRkVbgWvd5jJvuuG966uCuoigsXghohCXV0CYS6i7K6X1qVjUf5rLVFIIGPXztyquFwv
ekYFQvC/XD+JgTBtt5nwGzWEOpF9Q2XoYuT3/hFlgT6vr08w6X9JekClqxcO6oDdllDOP0C2cPeq
knl5l9TTFK5miupj4w0gL0z+3ZbNBmFMtJVGheNXYPU/WvsTBcZZDG//X90tkfKTIVqOTkinMNjZ
fdWt0CrtKXBPMGzrygo5xKd4S65UobJylBMRSgaUp7rVDjAggIF/KbO9nGTI+CYP4Tmf5ku7MkPh
w3J8nvTvXzrLa07kEI2YhyxBEI5YSu0YXhp444Prxs87n5RMhur/xY57hTYbaMWMI8mIZdLaaKB6
Gek6TXyWqFnid6DDoSmpcCfb5JdIBsQF7i0K/X5IcsVEgnBQjqN815F0S2nYp4zw5Guc9rIAMzlS
LUVXAUApyp7jWsr1f2JwBCUxjU/BfMwd0zwESli4RUHx1FqMBdIZnCzpHSTbLCKxoU7Q/pfFMgos
algUQls6PrvGgH56xmR4wF0gu7OVqVQoLYaBBOacbpVJr6lZhYvS1eQYYq3FMxnrogc8DVtnTn89
KxKEqZ4krh14KrKHA9bG0ZzqdnG8Y5ugIO2HLtqlhcQLq9RsRyl+ZRlTSjv8wgzvCj6Y0uiHkwcB
OuP1szzWH5s7AszBGZ9Bx5lEsuF3nahATOddz9ejIG0vpXVJX5Cr35nVqIOlnlzH5trraYf/xQ2O
hT0RKCRz0GivN2GtVu7ppNRNp/cV9kIKPBjK5CvdQPYe+4ixLFyjg/6Ho4nVm9FGlTaJ3guBJd1s
cOUaMpqEZaIdxHrWaAHLdwCHtI00Bj2UT0c9tFsE1TdGXHHDpDoLNuWFwa52J1on8aWDe0Z6zST5
90fZ5DLDF4L+GDcFiE4BuuTZ60nxNwlQahjqYzeU+8q1ifKSvuczHQTbD6GNAy1qGugWbkA9nCEp
eaRzHwh5jw50PF3PMIaMs33I8UJ0aIJjcTJfOy63obzSb+o5k1k43hw8IrWqV7S4H2VHpzLja/ZD
mBT6sgQkeZwAcvaVLagJxkP9It3BffXCrVSHplKRqzn5AqB8XRitlQy4/xYg3f1tCwQTHypX+KXQ
PV1s7P9httUawPkDOYUbwaOwPfroONKJcv+9O+cWyGSkJqbol+NKmqUL+0j0qElWuBjiQvcQv7qf
QZQRZcGdnBt+MC/osItIIhTwDNLDRAGgn+19rBR9JbOb+z19OVj6yZWfsCstMn4OfMceScvbibRP
hIWLWRs7/wivfdTy4Y+malg7AlJo0jJ8uD4gkKCMuKjQkNhNvfQpzH/ANXylzhWu+AojpU9aDK23
4nWRC58cgH2o/FKChttjqSE5LEX0Szhotzz4QUHdBZ9IqySJ5DLv0jXMW9HU7XzW8nT3YNkQHSeW
sE3vum5y2f2+88WbFUIYbMtgmjhfBF2SLSFZG8foITSKOyhr9ORvU/XkVpBxWU19HCFbr6rlScJD
aaR0j/Ai3Nzx4d98qnEz/LE+HdgZXXV34FQ3yKOpifFyeyDCOw+uo3OsKvI2am/Tv0R70epYGbCL
3SxNLtD3XvpENcuyOumLDqXLNIPfS4SPzx9mvLGs2eKByXxorLoC685a+AhtiXzqtEf1XS5xt9LP
cMJWY5uFCcRZvLTopvTvqQkGcsJBbDGSpvd+jwF5vXuOXAHQQ1HURrfVqqK8NOKkZ3iro1RCYvWQ
MFotDVoeWEZkfs7KmVdhExSKNYUU/YIEyN87BPHMcuX6+Wt1BQgMOQiS8ItInEQmnHNNssvCxHPj
5JfTZd3Bz/CxQC9gsxgVnYlL788kIMwQ7gm5qPh2EUgFvumpDsRWawMYCQK7DFHzswXlzQJ40TSn
XU3hGBi2bOdAqVLcyCHNQ6yJeC25lPjdK3M9jg3Hu6H3dF0bp+ULMi2NepfSUp50MWDYWpg816A9
mTecTHkTx64P9oaC4pkVMW1wsrD6+bIvkePG/kmoZhoRhPyvuEidMdi81lo3D4hM1ZNwv5FpAxSg
cBIRQoMyE4iKTkgwgcdcUiKL+RbuLqMqvYlnQiDkWVCdfrrDG2Xf6s91UqUieDsTx2kbfuQwssIi
Vz0bx+4ty2gvcKZ58isGe/xsm7a2G4n+Oi01BWkc3onjqzS/GN/yZBOX6TO+GMiNganBmioL/XyH
BN+h3ELVgV1L2FMyLt8mIxbtks6aWbDkREhIxZbOZDK5l5q3ePI9fizv1+8WvLXiRBTVC8K/v4G7
rfY68oueTqt5XOAq9Vhtc8dNtf+k0roXtl1gzBQxzcqe2hHgbD7bgwJRsnUKcEVc7KlmiALlR/IQ
uxM0Mognx9xnqDw3hFupa4okG/NuEfQZdgOO9kXU0oJFkHyHEVAx6vznKEKjZWaMvoPaQm4vo03m
Hw0/fXL3smPR/ker2H2kfa9hs7AQa8X5wEoHJxsIkgp1lAYXJ06maZ+aH2dgEpFvPbvQmOheFBpE
/6vgqC9oeYxUYPIYHrHI0rjOv4rjBe9gMBL447AuNCPcrZeISUtaC2T3TodlFni5cO6Tb+ZTca4t
rl1yHj18VEfEpqISGfcPg9n41+znuKcWPWg/cYNfaNzLq6tsDx343Ji0tav1gLZcx9hGHB74kbO3
lvK2YgULz8eZRDL4r9CzcUT1yZyl128XlZdxlurb4ViMck5UQX+/8VF6I3sk2jFYohvQ8yiPv0GT
dDjge1xED1U5exvEhsZkbc+JjeaQIe3+Pp6dDKHHDFUpXh2p7kAAFG7lbiygZh1hlOGVA5aUFSLs
E1YNjvZ0eIUuSmb8+bKgyKkwg3Ge1cRGWJSqo9XdS1Zm3fV2SzS7PDBN6Lx50PueBVz5pXlujGYl
yP4SW8jrMCTTA6rhFAKpZngZ00Y+6BtRYo5MIqzt+r2S3YbmS4wm4BaumDiH2pZ0pYGdk8C5Zarc
XEamopJUITr8uYPkdLaWKyq08SZj+2Fbs8sMHKcIC5DreUqZBMP19jWKsiF6dHT+qUaW/q2bsM8w
Ey04XBtAlPh9YMN6+7+hoOszUOXJDkZsmr8wJbPyycgkYUzEZeWO4l/LyLLNR528zQ7+Qu3Ogb6D
OmpjFDqiZKbBUTO2ZFNwIYfHi6eLRvXhCawW/ljxrQcgrLke8OyYDfYqh/CHFKSVoNBYxBqGe4IT
3Ozb8pSIKZhQY5eD5LFXONXstBlBmMDzvVG3eVaEsKYVQeFx6dHnL8eeKb3CEyxIp7nMiyBUWC4e
VhBJme0zBUMZAgSzvTG03RI3zXUmNtbqA+6rwtyfhSpdGIWWbwRQ6prd7n5icFdzDl7q629WbWaM
Ms1eZDbasqyfe9QDRmJNyriEoN8TalNmKTffKAO5knxuDb4giy/QFpjcnB8CVhYXkdp8CWHn8A4w
eTJ0bpttgPrY+Bm+7S8efUPk+WToJG10conWnv1MfW6St4PNOkTcJtiq51rS56kfHyOkgcBgKMtV
+15HKnVHqDhFmiO7dPRdqgrsWqgqUB0TMRzXMSq11qcB31ZE1b28rWZQ+u+myZwQrAI5CMYfqgB1
AJffiNLt9xpPYqcU2RWhiTKzKu9/mr4HW6TEv2iWnh3j7RuTBGUvAGk1EBpOUukMlWmE6cXqG5Ct
yzhjPu8AHHgiEIu44nG96IPzhzxAK9POveMWibBLv3UeUB9ib8ZN/rxKARaJYtpNvget52SinsXt
OTEdJ4JmSqdIQa3YBuaZEGYZs5vdnaDUMfDhD3wrgj9oFKV3gyeh8n/VrkvV9cmoitrZp9/i+Y0a
eHt+KBHxWmuRR4xgnriaBqBUp6kOkrqIubwUedGBo6mtgvSCQopU1wxzUv/edpyRg0aBXSvii6Uo
u8ieBN+fbMhYxLGrDJfQfDMd/NIOMLOyBgxvJbtYnHKPVyQtTohFznwfBxghL2hws5/J5CnAx5qL
82bAXoLrvc08MnO89q4UZUBLKqrSfLuZxa8VJ++EKjikV99wSsin6O6qBGiUOQq8unjzrvKHhi5j
Q3aszbsyjIuCexinqw2R3oOmqVgiAuQfvoC0kACy1MpJm1lvMwfKPIboDd001Pdp5OMz81r5jrJL
ngDv6UtmrGmLjwb+FUP9y3Pr4eeEY/uXOaiOUb8ONr0PZ739M6PfT75ufea5mFwY1F/w7U5RdNLT
txwPb/Kvhp9lqooum74pt9m2AwZ2/+4omqsDnkO9PEPmW+kHUEcKxeICdBf9KsoJmHjFCTkqywIn
xoOpfEeb/bQutsc7tH38MSzkwbukjVuFaUS1DKNwcQrt+X6IUf0XlnmKlAQ7YlOqO/TY4jZj+Y2w
MuLO5xtteCwOkgcFJFC3f4mz0eTEZIQrE4uocBnluCs0UOyPUe4+9GZZ0rujGiwQatECZfuX7rrn
FLrLUYkBYgfqNMAD+dqzcBAFPwxwKYduE9qG2GOXm8vNa459XqnEYJ87RrJKIq+ZwrS6/1LuXOnm
vrJOgU5ZNW4KuCHIkKZ0wj4JOBVYeBXsoAdt3pMYzo/d2yG3B3C9f6xzKzEF3MBNndIiw8FLVmVZ
6Q8BrwpGhy3u/gA+kl6zqfynpmyyVg8S9T8DyqsH10nbwdBJiSDAvopNhHY9E5frrW3+VdqpvIJE
QGMomj10pjxTCnTVQ+PdKUxFCj6LiN0enMgdH5R/9pr75aEX3ie4CnxqvVcIEFr311Thvn2FUBgI
vjOlX75OyCEcbDECF5GyIZLHnv6qK+/pUVstTR3f6LVGkWWbaubAxWQCyRQ65bPrhnc/LHHwWYgH
BGhgHRku3RRXMHIWj7XUnnUIbsueho9qNPHYHpusgFjUvdxQ3fvm1tYnzGmdX0wfsDcfItKGaq62
a/1qSqtyUx/sFto7xLufTrXgAyNDwqW/BEaSJCewkivNHqivMSjYdU41inNYngEGuU+5n3WF/Rlc
cA/FLWJ0AyvBiTQCF12vi6WHF/D3D9SIu/wrrnszJBwFQ5/tt3rm60lEjX0vmwX0wQxrqDBNyCVC
CrGwqRFYvAqeSeoW9aiteJMhtUTnydctmT2WypLnE1FzDlL5iXvW+yBE9dujwYD1lWZXHP7AEIJm
EK/BGmkUSMO0G3hIovC/Ov396UMOdDDt/YOst0ynNYM7tsNyAhcbacscmYTtAJixNmUDc7X6Ck2P
rT3EVdWvgA4EuWaHZswJsz2UNEw5ywveFXaiySlFgkCJfX4+ZXJBG0Qh9N/QLI8ZWUS4PALUeHmK
crnt/1nx5QtE+t/+Y10Dt+AIBz0CzQbKRDkqbRL3Np39XRBh4Nj8Ry0drq+olVqosOD2LhLc7QTV
g5NozxiAioDf/SR2IHVmhogh7FaOd7j7zvpcI8C7bY31ozZKxea+gapQrqNrTc408vzKQqK6bw0j
YZ8CR14vImvswfOguPHNyIRUUoauYp8Z4j6OVbgIcdFn+Pcqb0C9bCrtSu4oEB9mJgKknhV5olpP
yg6umzsUbqHqTwP21u0kwD++7cAA5KIUkz2R7u6kBUII+rAVj12xWhorC5WTBoNbt0hqDzZe/tIQ
tnFwlvTpoX8cpbgy/VtiNrHU6vfLwLGz3PRPnkfpOiftBw2m7ZFljwza4zzfZW3YpDBGWuxxWFzu
bNcLyU0UxcWucBf864EDyjnPy3zW/OFeHYB+nOB8C68TxSdXxG0mnq2Od8fIOrh38yXNOd6krkJB
kPizF1hFpdRXnjvTCKxxFKC0MaeusHZkLRx1+np3xieKzel3dM9hJt+pyVm9Bx8hGjUdErXd9dgD
3hwx2bFogUe8YG5JD1b6wUMSe+yLKBZWjgq94WLuymatDX7I3H3enW+pP0sYQWZ1lw3mMT0iSg5S
7Jc83xafmi/1pt0UoUztNjGKtloHyMOvaeATv1niV05hAwk4JtQTEwDRzoPpDjHirIFBcf/swXXz
C1rWbAWyYQRrIZtLqiWT72II10LmojzC2Vi+aE0itQywsunxch+ypkTenGQcW4OgifTAXUz34urm
6R0FPr2PmTIeQ511XE7Y8PafHVedTxGHQJbwXygqZmmITrRjwFOQw92/K/AdSAfo+qRVZ2YvlkvO
TnAf8FVKGz3OiOhXnPwZcFE0koXmg2jzBk1TlxwzqPAMfyDTo3tj79jL6npTe6KqXNTAVAMDut6V
67gSJ8nINfKnnJTmHUtxFQCZ3eV1f/7PqEkqWyK07SaCmSYAFFmnS7/0M8UqAL/VSL3Wq8Mibrxr
OyfzVPYrRRmvjdoyBZFCPW85SJ1lIEKllzD02DZW9s5qoeL6bwm54vSEhYF8QIFrXAjcTAof8wCz
CQtRz+yFTfBNfwBV9Nlpwiglo85zjX0CIIKlYUJL1cjFeaVXtB2Ir2RJ2jFoUjqpiBgtrDxJpsj4
9XSYe/ANlfWDa3BIJ+7k9STS5Ea6AcP0/Po/rxteOPFNuGgPlpSishWyniTcz3NrEPlEBzGaYJuC
U68jd0ygKxFJD8PE2/pPcKo6wLDwitD4p4xkiEVmwXC8UCFzTZ7URo2sKeaEhq9MxsAEajbmHT/3
UODmvZ6GtyY7QayQTzS6jthdmuaFJN42VMTR7bWU2TBPKp6iWt4ezSvtzS0zT5kDfcfSVr+Qt4eI
zBBMhspOni265VNDPKgx99tUNE89xvRK4/wVM2psxt6vKir+la2zPVUVE13N4sXX+zX6UypApJCF
/Hb7+BlBDE+bvdadimVpBzKtDY/iP13cWumaitsJjxd7NGXmw44dwxuhmdcRkgxhqbB7l/hmU7Rf
YSHHIDIhPy4tHVa21aWo8ZGYU+sQB5D3b3ASBo8BpYhr+dDR3P0gR0HTMU0AFDnLRDFFxAH5xCKu
aXwUmcG1SBJ+VjklcvUkDAP+KQE2DM0O+U9WD3RUKq4LvlDQH5y98xl3b8NADch7JfyIOJXIBELB
pWqV9kv48TiuYTw1rtOC9U82X+tHh9woh7nDV9PzS2QDnJvlxPxteBHFBXVxUUFmdMLBUqV7C6gI
bOQTHSBRZRWeK9Hqd0b87r55AQC2B4BIwfbhRVOiCm84QPe7zqHZ3Jime+xptBb7yo+KbuTDZCNJ
I+I2AiSApkUYf1EIHwUBjPQBjS3z2JtltAbK3bqwA7Ye2eaE5DcOJqRYhTEWzu+Q232OPuZ2kwgc
KwfrhaaUfoV8g9Azu8dbF2jUMuAnDuDPFcBPjQFUn5Te+hSpXS5YvS5+jRYwFxApONtS0M1RHWsC
/MpiG7VvVftAa56LtXcgYqvnTBAvNybhGiw7em6PAqLnStflO1xIkN2gjdMXxWuQttR0MxRdp9xj
E+fI4nXLCfdMpkNeLZfA6rSAM88K79kpkKW0vIB45bf1CnnaFC/3p+i4jE8qqBzam1wUZQUdxCl/
gshAla4098aSmtLLSVCchr0sc/3fbumIesA34VbkgoM+CMAEI+bKvdxS6KZ6jHT88IfneIyDL1Y+
4di3Z/5CtCsXMo4ZR/d91WLtAPXX3G3cs8DI+GwUIoamLz4yJhsJMsSJ/9zpW9TmPxUabkh7iYdO
jVkozlboRHznML4up+QvMYVfFsulhWqAVIkTi2oVRD1CVncQcdSceCHX36a/Q5xsggDX3bwZz69H
esKHEkUQe1V3umv9bFITYaUl+6IK0A2UDWARB+yTK2dC2+koI9uGr3S61BVeD+xvd13RGT+tpdpA
pP2M0kRvR9bMVdbQwiXlIyc8uKoydIv6riqx3JJ7h5O7BupTwL2z0BvRHJp0F6wQceJxqxnmAe1x
P2ppwPZAXvmDjJKBOYDmJaIY7XxHXaDDeDhLgX9yFHfF/WXxY5paRP0EIfe4p111EKzXZItKEI98
yS/m0mJymnXJ7bDGfXWYmZdrJixypBZ78l3mGQTZFsgbkq7Moea0aZxOWkqdeMNbpVHuV3PBHXn6
pbH+q9MYnqknFchbIPt16t53dKK3vChTbKI7Xy8mBiTxIiWI8XoWWu/y4wt80lCT+KhO3J2geTOL
NfUyormZxOwBhQo3Niw6uE/qtcHRa7hakSyYTlyMxF3pyYOOwJaOBXtFGfRm5jgxU2bPPnZ1pKKw
Geb5mX2BM1F/+x6ZfE18QcSpkX+EP9BjFGjvBHjvSCJ0LHuJUEgJNeFpQypayyv+Tnk6CHOeTuzZ
S30o5XTZOuQVF5mE8HweA/lYZaVqq0OuSRu0Lon9BuGkouLhBPgVWtP0r/eAeT354YL0c7O2dquU
Dbp1FdZSZD+y5lCHfhiLfu1fID9pon9D9UOlrFmrW+06GMtrlndO17aAybXSvKrGAg/JGIrdFE76
9x4sVPGKQzxy51AIJbByf7eMDvQzXVFxrjgbhdvuuQrgctNiBKXxLK8ioTJ9g0PkXxPLlG95e28t
WOCAEoElsUMMUHdrFZ/kFTKHpZEMHeQ8ox9TLbMTzEYDziN3kUon2kGn94AUqmyqKjdkZbAJeTFl
z6GmI/ZGAWYRlxlnsXjJkyW1c/uDu3exdl8qtPCCHnW9TbjM1zH7x8r/y1qHdsawxAXgo/SmC99K
maqpNqCo2Pz9gtdYEdoKYdweQyf7ksA/ffQB3xpLWxx+WBtq4REzVTfYMQNK5tBCtaV0DWZ6n5VJ
jIxEAmtR5UuC2BVXAte9VC6pjVPi2PdqWSE//dHNe2VyBScxkYwVppO3lJbjy657KGpHsP36Zx2K
m/yjyeLA4ChfBf6l5tEcrrOTLGvdNsOjP1+25sv14/GM5IoOaGluYqhacOUlMzNJIRTF9fX4L37b
9rwDTU6Iw7M6zMYjDITDHU7jqZNeadgnv9y7d5rPSIVq1yZRdDKzQgIG1LNoRDt17wsEYHpXusvx
Ruzu/tcjC5eB+GPo+D+FASZtobVhVG7C1oqRNWKwOVK0N6YrLf1b8LC1YsH2TzAR1zqXqoGDWI04
TAT8lqZZGwpFw6If1qYEcWLMKxpx64In/LS05TqLpQHp7Gbcd/aKU6/mdaN6hN2CIq920mUv5rMm
BVlGc9op+u8ELVDF8ECaUxhllMzTigsrGBSgtuKoUnRzdm6CVZVE1z3zDx1Pr4/kF9JKGyHWpixi
GPzlfoKlFdbRi5ejNMJmK8CwIvyxEplcxERg1ndVPXjxL6vGZM2//npavVWko//oSEE7whUWiVvh
T960c9Eqixcdh1/gr0v5WGK2hJl+QFxB3MnE7FYNyckX6PvDCWcZTgyCRdidusgQ27hL3vYVwCTZ
vKjfJlgtegI10vp8TJNTqbWAd/jFX1UeuBZtSuHQgJ6q2KtgGG711eLWOFXPQjk0lSIolfZ6ywi5
s3BI6jXumB53/1ZClYaGKM9zn9DQk8mJnGPgfBDmm+/+CEoyw3+ybfO1fVDDWpZWfLdmx2tp8pap
NjFsNfsVQQrtPzm+aWJ+c46rhIaVTZYeUsh6eBdoJn4JA5Nd1v4CFqCXTI3oWKKFqBkQr2HWyHwl
y9wZ8dpW2e4biTW1dk1uzZaJ6h51DYIJCkJVm9+4yoOJxEN08Eg7fczTyaKYuLo90uC/N5l+mEMS
feugW+7+vGNYQFj1cDZrzbqjq3Ne2me2uOFAgQO0vOzgpi46JfW/BQbUtlt9ku2XC0MeuRcg2avC
i2ilMcbYSB1Q1f47sr2vtGVQsIJlKdbiMC2ZP3TLtbhcuomOe/HYrqRhc20nzJtJks8cMcemHSgr
6iPz3LVYMTasNP2b9pR5c0Kh4gG0aByHeEoI85Ypa0Qi0SBdqY5zSKkPev89xZsCbjt05ZoR635y
6yltJ8UE8slcHHLSevd0ah+sux4TN4oOSG30sXCk2SGKOb75m/kAKzjWDoGSvQE6eQopr4y5C3H7
T0otMK2LVaMes68/aaEwa9if+n9WbUdF3PRLqmgZX2YDSgJJCumjiAo9olLKIPSj0tF8bTvhHRhs
97OQbaz8XveYAZ2z5He6L/tyAjgc+uviSBKZo5BGI5Zt3jHLGrYpuiwgNlirZ7BXPKWSgDuQAIGf
KikF9CTwEa0A20E1w2wRVUij0O/s6HLbvTszjDV4XDgWqBpyt+HHYJyKqVUtd/zsmR2Fc7a2EI2T
onIlzY3bkRCRjUPiU0eXGcc54BdyWvSSPeTuGfy5fEJu8AepAQa0jtSRXc0PSqw4BCgetlwFduwU
1uvhjOMAwghg6j6fhQzelXnXDGk8Vgt4GiXGgQXKFuJCC6V+18QrihOs8nrnBw2y18/lkPGXevHJ
vHO6LDanddmYEsorchcYSwUmQuglxGj2xw+O/vQKPpIlKGVmV+PzxBPePhnZb8wz5N7I+y6xnNe7
akfUlx8d22so7Jbbbmocg76zfOi0zBaww1VZfjdtd/1F0usJQvk9iq/5zC6z2yzcAvRxjKRwuZLR
jJPb/SGPT7QM4ZmAcOl/R9EzuEeHIMhflNM7Gcw44AeNwTvwKeCEkGiR8jRTZnZQHY5R5SRpVMkM
vOzaihk9iyVmOMFIBBERSxRQYfgL3ebDMaZfX/oX5lgT3B6/N19pHkULHh89IXw02P6Ju3iZct3T
F95D8/qUbe+scyBXo0Y+xekGCjIvUqNR4mokPXD4cIKvllldWNieY7cn59Iz+igfUiHZEfXvr3gE
tS77Zc/p4dwrK+r9Dkim23HT6dL5EAcBhqnGEE1HLi+MJVNNhYD3ogzQwS2jVuGEgcSlfiyMZ9Q8
AgtSs/ySLgTOz96TqWmGB2qot/ulbObsUxXzLeMbpP8sCVB+PpIqRpLw70vWtuM4wETaG7EgIgFj
rwl0wNfANJPxV0IubSWYK/t0RPO3SfrvRQ2Mv8YrPl5C1HX2IEXMvw1M8hY+AktYM1JJpYBfMkjF
f1dchPtNcWjRfJP9OTOdAmkUud+7/sZr5ckXI0fdobr9ppzQgcOFzRM/x2rjClUZWAyKZvBBTgtt
LCapV/DKzNz08HP9TL0vjCJFZE8No0r2J/Rbocf8EbavyHRUgUHTur99dHICOIhIXB6WZzJ7qiQj
eC7yiFGuc5vP8y03UMXqMAkLPyaiNAv8SNIF6u1TOy3enTM/SEC+Eb22Omqr8qqdcqPstgjUrVch
wfn25+JJabEUDLqtdZ0rxeWEAmcVYJ8z2S4YbY87AtJRLltAQkNCuy/RNG6DA3nAsq52ptcZlwek
WGmj+7UWx1+F1B0awEJjj4qcnu3IHCqIkSfjHNjoJXrQ1xqPAjUMjdNi3Zk01vHeIaN6gKheDXgQ
zUp8+yTp9ZkoYliDlvpsOpJC0Gkz2iwUOGYH7lAV9szqNJBwR4uby8VpU/+xyrNwSFns+OZZ9L8l
AojlyZUnkUYbvBImo2/G7ynIDe1XjrZ9cHt0TYwTAR2pMHZS8U56uggmLjiinohVtrLWYLlYYhZc
IQSyIgctVSpycRh+E7TjNSInmPf6IsujgAEyAudBHBUXQ0nus79Kg9dpsW9DAGPDvEa+Yh/uKuQQ
N0E8bSqtqBskzemLxGZCRhS2QkG8MepZN+wU1jrskxeeANGqSCUO7hB9gE3RhvfplWqIVpBDoqfN
b9vwZLGE/TVhQox6Qkri2StK1AjYIB+3M1m8bf1UmnEHM+ei3J0wlMnbsGQ5rRlQIjj+dHnu6YOD
xbt1cJMPCV2aynT30RNlRjvYAAX/MI4dvoN69yuWput5Gjp3XOvuqqnDc8EEiolOcwli/Cg4VBSz
LBzaCIYt6sQIoFHSuJbJKXRrTqrhf3+4X1PbI+F3m6w4BSNiGJKpROofibIN3O7WywxR4jIt7p3u
Cz6RVAVpAmchFe8wtsOniWGiXEXu/AMP8B7BkoPW8V0N1KhyitnF1JuEPWqV2gqq6ctwah+UPl51
hMKMUNVUvXLKExgclQSfCGPkj5F6FFamfIYVp2WDrRj4lWMHU7Ce7+1nt0p5HL36hjBfo/eqqa0O
YBFKFxH8g+5yzLyhYDDA+9CAEgBnjTu84a5PF62plRq4EK+aQoJIeT0heqxoG3/qpDjXXK+A7Q9D
Hm2PKAvSNC9e3lG8ERgTSI++0XuRUEnv1Nec+V9cq+eCuCtdestQ65klBinHpOQ//P5B03JSKR9S
BMYqn9t70K7dG1tEpCmP1KxT+e1wPrH1b5NwqP3bNAVOrYf/i5CJX3wNGZxAiCH7BsD4p8+NX0kp
DE9w4ev1lQIvzWbszxXby9eNS7iNtubNOgjskeqyv8XgrmbpvZ7Qw8NxImOiIHabbWDqgEoDKLox
NRkiq6qHhTn+kGFlmYcrqVlVarnO2K8HA5ezRaDTJGSu4Iajsnu82gt7Y/AGU9QcQ8MOtT6QbeKX
eBfHGPjh6uSHMu7hPkcdOgQneRSd7JTKCyACx8Hxl+7plz+LtyBTCZAPgB+BAbK+GHh6URd/MmXh
/8lPfENDboC98/AowmlRZwN/wiQA9vb+6GC2N7Em+4fsURfarlF5LbWQAxVyTWxgNwKlXpyYO/8+
jf5Nwl0byWiWuCuJjFURKIEl8Pv9reFzjzQSSA/PAiDdxiQwS4bDXGjt0bYDOoZTKDVoz+FFypOK
8yEvVSVoMtfZx5g4EetfiYFIi4yg6hqBLvZP/AHduy7TDsfoNg7LPo5Gi0jGHJXKnObLucQw1eY0
gnFtroXRW2UbGPDgh45L3b0OMxbKJMl4/Tg4CPOC0DAYxopAnX44YsVccMBJMt5ZSrzdUME31htt
g0EKhfTnUjTjc7DzYSB0wbo9BKUC3XHLX4hRfgcv+yPZ/FKgKnCO99pJ6DFyJcI/6w57foLpRveA
vdRACxBuuZ04YAr+UR/s7zYM0UD+TcbvGE/2KIn1ZWRoOi2LgJKgo5FR22sG1EzZmBt4HrrzroqJ
gHG5pxaZ+UfG5TAAElx73vFOIXsmSYiiIll8j9bv68QN1exZDLoRY+VzuUp3Jtndju8Yev/J8rEw
mKXeKo8p9pRKQwNANSE1uz7bjEwTBplYq/OQgkpkGhxRC6UzyWShsFScH1rFTYEQDG/3kyncKhlb
hCwH4LdtAQD3/sf0rJaOC/VvypALbp5upD+e1g7TgOojUOVT7rkc3mB9L7YpwmJ3o7njrNnniX2i
daE7rcG/D2lbTpHGWVcAIrtT//Xy4Sro/6o6b1Ag8+RwrC3k/8lRBFD+84xil1wTpbeTpI3x5l+R
bQMqKM8uc6vc2qX10HSvs7tmxPZimOkfvubMoMvALBdgMRJLTo7mM/8s1hiZ33nAoL/zxMUTfURs
18TZWWwdB6/BFrjDyoCLbzYaHGRfKORQzCIGugoayYZW8M1uFwJH4p+d0Y85eBX12p4oLv6tU3FD
4eV2Pkdi/ydY6N40H7tgEhLsxawlv0aTkAUdGKE3/nCwtMqsI31/ji2AEc1atq7+dMRH2HzKs4+m
5g441XqP/803iA2qJsmFV6YmW0t/F7ZnxEBw8tKDZpIZxDAaOSK3AgO+ST8QiTjx6P+bq79yeIgJ
S/soCDd3hSqB0TTZajyU2DO90uokKvTlhQO+ln/Uz4ufMWphMSijEmmKmmIIF9oXgmhVi7o9X+6n
yWw41a0QR+H0pDx3D36p6W+G+uvrsKAzxHR2GiVTnGu+x1BIZH9KlWG+QWGMwNaCjN+BULyDw81n
OAjdiqpdxFrfUCMKH1DnN6GabuWfs0Dv1MauJAmw50Zf+GF8iZrZ316IqsNc6G2i2Pp8pzQcLcZM
zwABfQHCIyb8cZmURohMRU57X1JflX9VcHaRSBbmjVGH8PpFcnGBei2/zUm2zQKJhgtEIvxNEXbT
BmeLXd56uyK51fQhgBSeKlsm5MzaSm/yIMaU0P3nX47wcF7NJReUYnvOdMPh2yv51jA+49yOr29Q
9HI6dx3Gzz/0vjjTv0TiOzyfXk8H3Mo9pVlGPkm37ESgZ1Hr1FGesPIGS7YqaHmo2b7IQDgHHoBc
MAbbA3+CvoOpqAOuQtKHWc7rxsZLSlOsQpaEVAeC7OKW+Ifb850RWShNV/2rkbchFtHNmKI+UGR8
O/IqTnNKofumO148rkl8eo2RUEG2ptacNH+h7CkYH/16owY/7bsDBI13qRt2W77glACcPOMw/ZWX
ULHZI1nvUjmc/gJimYMNwxgJjEWg+JgoI/DzJRbQnLQqW2eKkY6aMCxXrIlq3ZZPwlywwbji0Pu9
NoHvmPdv9cKcYJAOyntMjnwZw4fijoZluidbFVjAXkaD9iDpUYEAiHtKTrp/CSe/1Pi/+12YJUkJ
Bb8ni7c67qz0VDtLMq2e83wFXE5ZILtVo+ACmezZiJiw3cxIJuodf46Io50U6pMb2hAd/Ryn9dI2
Xeo6GeI5OesJqrF08eAlyX0pcgL1/pJWNA0x5VFuyCDIPBSNsL1oAVPsv+pw2iTm7OvHs40wDk0a
+ogI61CXiDdmUM61wvXeKVIT39GWRPbe9UG/FlKYT0tHXwph0iU5AzDLp8ly8i8ZlBWyfEIXX27t
IrfrPTzlT01Rrq0TBNopps6ce4EdnWbdC2AJRrlFNjLtWkdcDZqNFVBv4vj3q4OzBnoi69SGgxM0
N4Xf0vJw/+qP2bl0DatYJUTKwo60Rg1T9qddkgtjGhJmHDaEzn87GrAeavlV3tlS6+KZ09ITUn2V
1b2sNow/XczgZAIyJ3sAG3iVUCJLG5ETxyNt2W5mJBewAbyOeWHstsp00wW02C1tOprPRmYt3IkN
LKopJflIAbRhYnWfzjZlDn2N+ixVs2LE3e3lH3yq5RCJiX8gwQORFF7uZUpEjp2VdHqIWtrZ3Tps
ByV4YuLAWumxxRKoHCpsepIl5cn+IJapDVal/6qhn5ufC04oCNm3wSf/UdzNISxS0Wml31odjMC1
K107Zt7fpXB7ShTKcGpXOqbG8dNPNM3l+Sn/L3rvnYeExYX9SZNXc2K0W3vj0blqddw99SiuNdJQ
AazupdPzQiDNOFhkm6VWCKXDvP/W/pzu4cyO+4a7NDqEnUKJ7EUz287ZjxRwO6LiC5c1V9TtqrVx
Xw8J/xdGQNTIxhSjvlXVProItHScQkxMlgFJLd99AV44WYRzs2QG0f/5vW4V37Pj2SZlAYWYXlhP
v9x/sovd12tDKzI1pT14lh6vAP590YgT2AH7hWo2hkVOUouBKyNVywh8y8zWxcojSo9p2eR7epD0
4oyD3XeKB4ElD7zZNX+uil6RvvmQ/++9Iwzf6aqFs8ju5OegrRjOxlLAkanmsWrYPDizf8NfL8T3
KqD0X3D2s7LvzxthXjlLGoR6R7KscnxOiUs7i419eSAkO1xcDXN4gRAuB9KPxPTLdkCQth0YDkYJ
dXkbdUxyGq7yUQO+0oQ2YRO5m23pUFmqYUA5dorcurRe8HDsFCbIXm+ghl9vmEL+5+iaHPENiDKl
44sCxqQpxDRx/t4rMWTNeUVPEIkflkmEAX0nxXpWnuTJ1IdyyyNHI4SHWtg4CjKWb79d6OBei3Zp
7mWPyDT4yeerViP+jU0vavt8EXYQ9ANu5n7/J5diOinDeifpS5RrLEVh7urxUa7gsB0/OFwlF5eg
ZUoCJUhvaNFuwHFN/bG3zKxMGcs6DB66/92lUpSiobzD+ZzShxiidZ0HqvskKgAkwIlO0MzaK3wi
CETsVSkKg2ZCChOt+Tmg7Mruzy1vIY59UMqZoOh0ZLA+R3DK72563QX60rU3VuoFJny9c2zdbd2q
n/QF6Xhuad736hkXUX1TjSTG5WTjpEUlNRxD7eme5NeSHMvlTIbL8fbJGaTiNDyvtc8cKa/bcveX
/CPscYsT+H0xVr+K3Gio7x8nXAp9Luy15Du5RPHmiscmKpiTCUEiWVIy6eNQZiu2myiibEG11+rh
SzK3c/rH4Qv29IaU/L47KtjQhFgiPtzKJOZSNmO+KQ8tPIK9iNlV1a8GakBgP+4XKAhgtnDfSMeD
NzLJsFh5xmxqjMG+brJH9cbUyqNLqlISrOt2CJj4uz992D9V18yaz7Q6EgffCdbWQ2CSsgxvSV1u
N5seuZMcnIy/wJ3r+RUNiLL7qAkcpzmKZKRZYuZPtbW8dvEMpYQOiV2k+AEdU9G77UnutF6fzJTI
L1bThxITWRSsQj48hRBaotOyCSWo7FUPbx392NoWmM0yCwwCMw4CX3bq181TFAJ+H7JbgONoNTGO
EovgXPHx93uBb0xd4x4MJI5TIJpb0uGG3pCRHyAYfoX61NWX5FYTvHlS//WzPBOI5/GYT45rCO4I
o+JexKBRZ8Z3Oouw21qCXRkiozIUVBwPQqfch7yqNzPYPU4251yLWLoNpTsL3XjK+eId/aXAXFom
DmlsW89Ubn5MNiFjORmqNLfCCekDAiCVhoOEVptbRB95bfLEht7qT0iq4ty3fkyZ+FzG7RKrXdg0
nzV1JrUpwL4SJPz9MvXohqw7qmhZiot+f0/D11iFre23OQPRHwXiEug8YWpQ7+WIezf7xBJBShV7
ZOEurE91tEnw7UcPblY0LOVcO89xbZNZX8Zm83kSRmomjwDBRJgUtx/FMkFok8KrXQTYQwAXfbbs
jvscn6ystoDg7OqF/g33qnoquMR+FM7gW0OfSAa/KyWawby00biTE9J//4E26QqyvfqFEtYuugfN
9526bW/ya+0snzd5mUJz/Oht66ZdznOmy3Ozdotr+XLEhuy/34sjE205CicuZ2VlIfgZez+iTXNT
zS1YQww/1wWXS3o6wr0fePRnTXbO/2wIMFRHBDZuzaBnfB8Ca9BCgx8ohZM1r2bqD+XpeLAFrIWa
+G1HWJQlPwucbHA1U9yCSkDLv5gMLKSw4Cuk72DtDE0XAENE7XXBVQn8sJevEIamV2938GCxsPXr
dBdP7bl9MLW8uuULidgAMcfxclybVSfrx90Q1wNotOcjP8HsLNJ8prRRCbZ+8rhkVifyWtU/jgGp
XbSn6FPq6xoMzEyRPBFdfBDkng1Yqzu6Bu3IohqTUQq1REHNFrL0N1u+85ZuA0KmROTY4tvHvTGU
pNKXRZwEBWf9AS9LvSIqO4NSXeCaKvhCiR+FsQjX5qjx5CN/+Gj5pvB1s+c4FyP52eNJWpmRz5D6
CY1H9RKxIUkaCRblNiOe05IFueyjSfz8Q44bweEfNPdrifGUq9fLjJJ6SrGstJP/HY1iqngWKnHu
Z/IoT74EKd4yvrguBopH5gK5UwubdJJBcWvRwLEh8M0V11gIExD0rPSGPMY+Ze8I+dri6AyXt1Kd
ieQAEHhB3lH0xif2kd8vxiCVSAve/8krP4QZSBTH8qrEmzvO7UjKYDyZIVk2ncTO/J3JLF5ewgGH
rjo+NOAHswMVvyRPZtPhaUnaQz6Mv9fJ9iMQqKomEaT4pjC0aDnkgZxYqYW4Yv7hFoAICjKCX7DG
fYBuBDoXwaWMAINCQv/mRdsi5SAWAQT61GAYyd6lMvI2zHDeLzON59Tlu6tRVlPncSKFUgcRPCuZ
2eU6b08zf7MKBK1wp51f3/k4UD0OP3UBr8fp7GI1tWid75BFXmcVKAifYFWuXYzBPc2g2R+hkowH
ftcToZ9EOS45PKE9p2HoNdgv1lDMU3JIPxucKBiW5MMkL687NS5B76yl8nK57KkVd4sAMenM2f+L
BUto1j+azz6z/JY+XEIZCPwlBVvLh7pyQA5UIMyvvagSCbesnX7FnOt/ReF9JQYYMT97h0d38iqd
pdbbdhJh90FlwrEY/pue0qlS7ivBuUPkLoXjY7wdFzw+nEkHPnd9rx04PK/KFl9POFlQcAFzXBHk
zWW6IaZtPkLvtIWnAGKVhTHeys6e5NiwGkFv9hBlvdLXckTLoc61n4cvGaseciuMRSyd4HR3b88V
yAtOzKCIJO8g5tF5MMjOSu5ZoYK7I0roDSY6VCkIdwUvZc9etyAQSzEunIdcWTJsgBaz/1cxqRt2
I7nmFlMg9S7G/OGoSKwc8wiBjGym6uQ1rENdrc0iL9f8Ka7x5S/ecT+g6eyttf2Su2Lhtel295U7
uGRTkZUsiDeN7us6Lo3hQnx5vVuuuUSPypjR+8QOYIns205nTEAcGqB/kMjrxO1RVV6sBtPZUoN7
hdoXDUNTrJAsHsylLhGfYb9NbXWEhM/n7V3TkUbvX8EU0BccMncDOLzayh0avZz7raogNc3QvhfV
hYMbBN6VskOl1iYSDckVFXE83vOHHk66PQjHADhRfH5RhTC0URJ9z8vtZgqnn3bxFRRqW1qTi7E4
FCqI+dZF7kWFzzTgkeKeOSFi0PwkavGZZZkpSLkN5s/DftujzeGgEArNMe95J8mxra31pXcYPO0J
DGLy99gdACM7WyzgOiavbaVTKmtTeJkykcIrA+7Ku477R2IY8gjV9zVD6k85K7r8w8FZf/2gNDh6
zw0GbHA17RUlZrHya/SddYwgV+wNNjJGwL14iHtQfQusXdvs3TERNXVLOr3eStgmDUew0phpXJvl
C/B88IT4juxaPlcsT/MFqpsiHV/+1Jw070eg6HkaXLC3ZKyhcoWgThC4Kh8ZlHxLoqCAXZTaqIvQ
h7Hd/R1b5gaIUBFxHMcdZ3K1Crbk0gw7gZZzHW2xmxwwB5eW/gBs51T4L87G3TNppuf+uV+f0dv7
mG7Z2ojaao2oj0vELAo2KqSizW1fjf5SCFmPB1e9tiO2/gUb8CgMAbhaHdGAjhNQg0E7fHTgWHTF
j3GrAKU5PbFWR0Dar91ntiv9KSiN740De1oI6knAncGUDXXKhIQCoVmDK7v4HyeFeklhSEUuufwx
OQ/V+UOrybxTUBPfUiEhXK1W5wC2zaZO7s5WVLtn4Nl22KbhDHNLTfUVi33Q8rASmAmaYBheQD2E
Dz/GePdo0wffBUVacdgAsK3N4s4n1tEmgZJf0QBfqC30lakgsSuJdzpO8ZSa1h9HvFQeXnKr8Bp1
/T5OFwwy79RTAW2Q2RRrd+AunwTkWWvdyNABG+RS1JRKgdIoP6xfIzDaX5RVt0xikpr91g8E1Kdf
wHPrWTK8izwGLENMOEuwySCty/ih9Ku7IyYqlOqalcRG31sEGxbsb/AzRsztPQVOG01ouVtuX95h
h7SH9EX2rg4jrBs8Fc240BGYQI5T+x/i69NHy0cqtOLrH7Jc3YrxaFsbsu0a9Vgb3tHb1DjSSXfS
RFFIEpMfP7hJj1ug/fwVlm5nTQcTIY2exudfq/QyaJJdxb8gabEUcRUadMx+k8N2Rv5jjlFtjYuf
T14m37+RAZTzJT4QuQX0P26nqqfishhcnLuseagH7ispBVNyI32hX8/1QjIEnMire4fcd1y0o+1M
FwxAxxiOE3HBMmePx4WNtHuxlR6xSmudkXb79Fd4x3J+p7l/CShPE8s/4ZUpjtqgj07K4oNmTk0Z
p7IX4eyqNAdG81lAV61zXr589q/8bFkRT6eq1TL4Oyyg300AVWK7O8Xe+c+x8mrtNT2Uyl2QlANp
+/oc/5clZqEc7h9mr1tQthn1BzytMUajNusLs99HICoFilL7iv1gAf0Ebw3+DdbeRmjMTPfB0H6V
ImTqP4l+HMnUy6tzXJZbperUZL/07IV6/1k704xzVWu3KlBlYkic+B7GXZUq6ynJ4O+6ofESE6HJ
77aZAlsgJRPUTsjjE5wuWaID+nadwRcaZJMn9+43kv+v908j4VvwvwiQX18XPVE8XnlikMvow+gP
UeQAil4zT0vn7086WwtRlsBdj6sxY7aLbdAKHTI2Hu8v4erxDU+Xx4mBNaxnJUBbMH93Q2V76kvd
hm8S0TZiAAqZEp6CFyJW50mYxKQvgOoLtx8TiLSCDZRx3n4pS5uiUnepb/Zst+SpJHC5yz1JAvjQ
fBA8tNCSp/QpCjhOQp0jEbwHsXhqHdU4g1dripAX8kct9lRqb/r5wcbGagFyXvgzm9mVJbBtiPMs
Wo/cNMl3lf4HvCjD+MWCIZWkSLTOS6TyDobUYgByVgU0Q/VSdelu1cDXBWFxTA9MUWLNp186GHjC
lVUSvnqvD/JeLYMpij9gUV8EDAGxlJ8wxym/H+YCxUcvg7IVdOQ8rmDgr2tvUhKHPOgUIfCkF1af
uD8lqfpPRxKYWePnxzJFsFNdTqCRz8q2Fg5mDOHZF5Wkdw+jqccigTF/0Vxmyv57QjJFxjC2LiR0
om4BFzow3qX8TloDQH0AXHZFMcIVfRyKFO31D2Df4F/ZvsnxnrgP+la450uzc23tMa5wUSJQZ2CH
IP1F135yThxxvBHkfLtFfLqwP1UuP1i2817xPlS2hem9+V+FUWSdjHUdbzwz1MutN7PYCPfG1m09
LUg2vq3tjY+iqE0nsAxiK5lK807Ww4cf36sOGI2weXMl7S5DeGTCF9b9kHFWqOZFQSocYp0pYTej
Wzahqlba7kqvICblk6YT5o7Jq2qWcSo6Y/HFG5QvV5Bs8sGEyPREaRDmSNDopzm0QSNpFRl0MS4D
X72iRd/7X92FioJLTxVEI/vwt5oQ9GpkfND8HsuuTyXheV43dhW/1CMpMlzYSVSDKvxmZMDCn+De
CaAK9Pi0svCOUPt9gSMTBd4e523fukWwFZtGh6ilnOPln/mXLQ5nQ+9EYu/+sGxOLp3NEcuNTMwg
OA2kpyeIDwLIEwIyJD9weNS8R3PXBaze4QfhmLym9hDmcBCvNa2tr0oxQvfsfy+V/QeUKxXC6uBH
BlXnAxIGARUSg3v55OnouYc73OXySmTK02SI2CpIzcwJa6hkA3MYOhxVBuIatmLweg6vpP2zbK/4
+VkR0K9pkMxzFG58NhC9Dd6gbOU/Bc6XmcRoUu8QMJMlGqdEabNJcMdoyExkAhqR6dVGhI7Ge6It
vHZsZ9U4ohlEuHfe9/aq4v7Szc4teEOo/QAtGG56HoQL+xNVJ9K1Z2rgx+XTawHMfreB/1pwnjvz
8SDX9GKsT8huOhC4uINVt1ubGO5CDleOE0ley6mfM9vu9J4aIi6JB7NCV/QKq7QN1G5hji6vBug3
VAb7szZqHbWRYQYSkf/ZVG2etyQogRLX63oWZTDEO05Wc20zKZspt4U7S519RiQfMniWfieWoi+o
XveEKhDmCVCk+8jfgAat00E2ZkelQkguyqJTCNM+LwEyrkgqMpQPfYeEpTAITXF2Y/r5a7JNWcn+
LHX1plcs9yaJEclTH4kaVbtx/DH3/DYygS1ZSaFxSCvM1K9P++BQY+JOxddreHkE4XNxZLLmMJzt
WjbrLnVZF9gIMjfu8ah+CgYXgKakX5YU7dsykZ3ixplpocWZciyFTuOfxhLFudtZdlGzLk9WAEN3
wkAwhAFmflLWMVpvMtub/ow7TfNYKsdHispoOP6bgfeNdhQ/sfZsY9agUDsOT+jOvcpIZDs2cBJW
qArh5lvYqytww0kQLQW7rfPR3ipP04r832u00BtpTuyDblty2V9eeIF4d9njf7dnqx00f7kcj7yH
lIuDe9eivSZ+NX+yErX8iL0lD95o517WqJ8HSl22NPDZatPUnofJg0AbbgNf7i2pmqJqgf+Eatge
gSn19tEMG8SDXrzC0qRb8xtfVOCHpSZ6zD9LHRnij1yUDA00R0Ug1kOUDQSPlJ6Y5rngMxzJavzm
tb1MqQOxvlBw5iq6i3MMNI40Il0McZIUYZ3+MCdIXAobWTCKu/eXIT+pT//vq3Ta+jjBG/SbOvvt
xZUZJ/MOhJz1PHIvml0sGD6CPN8J+o8wSzB1F0Aqe6vxzGEhAmufi20Bd95q/m2xfZ/atJ/EIpYf
5mK6xBy+00SIqlo/FSGnIVKDBWCqktVCZsm8NH5UoPiK1Knmp94Ov/LR8jorHqH6Lnv3gmkAGBWz
Myjng9SD2lU7O/S5dGZrzvGR3mlJ/6jxu6kyRCPzScA58o3I/nOgtLogsO7CqqKIaIn7RJlRGJyY
PpgjAAnYYLKdalPzZFZsc1VfMXM7KEeL774bsMF5+dhqNb2mS2jD7O9WmrwxSyvwZoUj2jvaUvqY
9w7i8Kr90unlgyJ+0aL7KnSjksGACd76x8i+7CoAiKUfay5xarMOJJkOWjBR9JMjgR0xQSEEwpnm
ITSEzUjbr3kO3ZE4vQP3ECp44Vyb/r205lEvv3UjcHh+w7ugRuMUtkFTUshTGJhN7PIGxrL+y1mz
5OV6osQ259causWznELV0peucU+445cH5XaiJw6wvr7Un5NdIqvuNs4iAbsjPh2EJ+nzIN/d6wEi
hFtk181Wbf9g3VBT0QU+/s1Qqge5LH8gjGmG2SqeBOPbwRDOfZe5cI0DfapPZ/ED8fujb02liDyP
yQ2p/Kd9Itd7+GMC4kHTjQMH9VDrMp/gbhIvh49eeoFoVogFH/QgVl6pQ00w+OL23FQ7pX71n0qa
/FKFCaNPOUj7gMaisos4o9HGe/KyfYuoVVMGVoRDk0ONLbAlrTILEEP52P6EsctdSmjphCnPO5Hc
UpAUL61Wveun2i5gL2/MDf510PM76mFGEpFMN2pHJyiweZ9lmmBuw+wYlwnV1cDIvNPhOfrIRwoz
3I9lb25kbI0UeUySPmZaXRVbWaETnszmJ68gQRG3McvCOKqOqr0JSMbP8ejgoBdaAtT9K5zHWZQ5
XwUcHSgjcVpa3t6l3XMs2zzzlMWeu2rROGakpbzuhvf/v7twprsThQKOf9T36T5ibAYe9KSdll1N
DzNsjs2yLwFa1fSBlxsf9zd9lxj4cVOX95BW7ioXIRibEUvhny+kLt8UARWbOhqHje8npXf3Rlsu
U9x2SzP3piyVFi9Psx2Bjn7gt8yVpNfb3ymXCSBtaTqMXFkZOq2D7sRqxNWFJw0trERrqxxlrz83
6BS+34+eRKpqZ4FvZMaCJ2BQ/d4LVvWkBgBQnBumKLRERcWfz0+C43zr+lVTG2pVLSB6KBxGyHlg
nAJa5b8Ln4j8APNj8uU/mKViqhL17j1deVT7DlPpTUH1zBJDOdgCgJML56ZnRML1eZNNluZl10Pg
dff+GaKgRtYPXT3P+QCE7RXbpSIoqlqC1Q7FHqXLGJDVXbG8sR0wNUqGedhdF2n28IKJPjROPjvE
AfSQX6XmDgVTEFbTl+aV7UBVAwZ4BLh4ZUIowyWNL720OWQ5sEtnfqh/gusjGZObM5YR8faHGwmB
x5E4WiI95y/FcxpC2IbH+DQFqyvjLfqQ+oRXqeXoqE+ljl5ZUfsEFXKyf2MI517CFcrcBAT5+6td
Ojh03N/MZBS+nKontnqoDW1bwHmcii6QhrGRLv0tNGlXR/dvX+bBAN95wDqHRaVxDHZrvC74vLqP
IBWAMOuwKdzoHcmJulR+lJPkR7EwpzD8acPrxdEHPViUCe2Rya3tVMl7aUXn/jZMfaFX62JXX3Wi
nIeHkOmZY/zbfysS7Oye8S4IKb3XnYjmq0SISZx2wfC5i3Q+PjnjlDpqMe6Z0dFpqFRfDXtrpWBh
SjjAEaKwPzqHrxUh+D+Qc9phZdmiP8C1JaQboKAAFv/zZ5Yuse35/dnaMI3VnMghQQ9Msbuli5FB
D2bYM8jxCYuxB0Q+6yyzT8R9qihQynz7Xfnz8bvZbo/ZW5PEaQfi4B54TVipJoz9fgF33CnwvwTe
IXBXLIfQiU+sN/f+RI9wcYPBjb8MJzji1UVeF/mAAs8BfpVFuoc7HOB/Ru1w74Y2Mp8ypeVskvH3
0hNluBNIbzIvCDNYnVnO19DHA/+3cpk8xfx9LyECknWNwb38c1Ot8vSa7u32BnjjbzrQQaa65trE
L2HN5zOKI7lzUUdYlaXctEnJSLQ6SYQ+zYtSsHLMYEdewJHbH/WQ+zBuOfoz8hJx86+23JUHoJCx
wDs5vEeg3BMQc0KtRJlsBpPO39Cc3ttYrf6Zl4C05mkfNodA2QLVFWvLDp4xv5tvpIqeBX3uyXv2
J2dplUvYC0cyUKvUoFTJCRmjJrNa9UCTNeBhswW2ad4pK6gCkHZRvzPeYhkX2P2S/Jpchgjqfdwx
LDfVR7S09P9U6oLkLNyNBS1JOyHqzFYayCl5q14wCD2KLGBRTa0Ua1iXGBfcZJlVUEJZSt24YTfT
AcHVt3x3x4u7Td7W7cA49/Nj+H7+BJt5ZbyRMVqZAyzt2gpwDAt3Hu2sdFrIkQSSgCUGZ19vn1Mh
uxWSIHbYVAL3B2HHTDIhOK3ta98yKnUfKPhMKPwbMIL8bfc1jKOA3VniqwQZ5okzcKZfuFt4Q1j8
mzOuQeG3FaHCs+gQ+2NW4eXTx+uZCQTd5OXXdweBihB0utI/Zv1+nopoELW3P7749FbSzQGrveSC
IvK/lGGFB0slaL4I2GpDZX+TGD1TT42kVj3y37He3Nc2tAZyKIdmTtVHra6ULKnfeH+jLyeqQ/58
Q8QrX1gqR0z4rGvkovI26Kag3dmR+zXF+tSuVP+DdRHczICTiE8ByU3LdcgQfFS43LeaeTDp1fyJ
+7RN7jhYktiWRIeVMaboChJMCUA29EwzTG+RqPD0Y5FfygWFxBdwIFVp++P+TdlirKQti3p+ajA0
IWi33COeaKe/c11Iep4n9dunzJkCuhi6I9ejOxR5ZDHUe1uuZwn5zKk/4pvH9CnJpMM8x7A+PNEP
jPsxFqlmmlhYrzZy6y6A+gGyUaVazg+TkXEXxAuy50UEWqE+2Zpt6MHlbUrxEjW9jGbXFaBJcA8C
kwrGGnyUuQUeUVT0PjJ8T9rGYfslPkkMyT466ImjcIBYLcFVConCR8627A/BWZqEcrIABTv9v9L7
veEXbiXBKGFIdDX8EjxP0B+kVTm2Z/ae1/ydCL//+Il95U6oQFsJjI/4HHRSgJEnY8UbeA0pa4g8
ymDVwzDOPFS14lixBy0xLSN235T7Wl24/Ecnisr5vr/dtqIDby9TrKsfX2cWDOaJWZiMioD5jLC+
UBQJ+OQ06ZtI+LXXAcWdeQPmG0HtvK+SS4320hUNvVrlf/10eXMsEcFEAjr9tpo4bEqTT6QZnQuP
oUta/M1z6VvPXm4Ml6iB8PaFddTy2laSy092wlD9xha7QSSY3WtHZSvEimUjMhI6K8J0B6JdPZ88
C0sYR5v147IpifleJU0UIsrkWRmE25DXKWbiDylg8FCpL6A0RhFzrEyBNCYn8BwWIHg0qAEyu7L3
Xk+v3ekQT+4FqFFYLC793sJyDX3rYnFFJSuq1PYJsrJm7FL3A8t+4y7U3gQoEJCoU+3VCMa+CMjs
G62DaidRprpyG+fHIAQ4yqVdBhV3kLbdpW+pAXwsyPXxMohKRoNHj0Bivj/ABpdYfkJdpcIlsdk4
o3q+28U7Z/AurUrVLSFaobtxcqQ5FkAkTaO7MSCeDVLR7DK1Gfj/F+8PiFylPhjxX51VmzmwJJZs
c3uAZOdJjIS1baB41qma6Heb0oF6Va+DKGYYcgigE0pobALLb4Uz3V2ZghuLoSG7KQMAS7ZRIXPN
BrCfNwbSsXg2W0drdJW5frtE0wRqLUDgrlsD00fQ5w8SLb5YB5YMfY/2o+Uulas1jjV96+tOyjCp
HKYtbaVI626aG01+k1anOgUKCR7pXo+om1F82s5oVDtbBdrTtVnnMQB8Hs7OVx9sjSAjfYpk6HMP
CW8lHlN2BeBngPRH/xmGJlWIs0MPuvdc9FPKt71cbm0YspAfloM2fPQw+bWo7/3Jyt88v8ot1W4v
MNwupxIXcZyq9a0rU9MTniESuD8XAicOwOxBFWU92N3BuuXZd2tuHJB95B/RNfOFHqTxndXxwFoU
JTUEFW342XDFj8O4IdnZS1cEN41NZpxdYJ7OqQzxHqkT61R9kafIB5WSoWfSij6NR6YATXF0CtNj
i9VaSgUxSZTcttT91eZ4stpMIzpcYYRtuhcQtfMV9Z4HSMZNBrf7CMYsit5WDmLwmfTJ+gaxCgCM
GhMtMFBSVvJbJeLUTVa9CCPhOQtLReMdg9+JBJrm4h1JlWt4gqgKxq57dkn7Yb8KXfIFCpr4wURh
g5Zb5TTNT6xp8zXQ4hSVtixDIsw02nOPOdvCc8EMB8w1ukhqPGq8STfjM8Vzls5TtIyx8E2WgIuc
GlNnk9XtJfMR4cnrPvUis1KEt/jBGNPIMWo3867meK/1WcwD2I1iiFCi0nTEtn27flxmS3h9bl6x
u0Bi75dOAe/5XkNf7VZAaKj/NkqacLSAmFGPHFszWuF4itgEWQT8BTIx9mIS5eP3jWCSA6QODlwL
a0Ph6plcKJmf4ukHyFthARrMzh3FMxydjBYrXvW0g3916gJROQr/VOZO7o/gup9eJn4OMmuvMSdk
KeIjxUqaluiTJ0gOb8FJepILG5BpsOfCPZHMbEmNt0ESkoROV2zabFIIQ/y0kYoYKnr0cy9mhpTu
vQiM9BDlpreA41OOR9cbpApel8Xct7rL7yOrm75q1zsedCdIQiQk33cLJaifxc6r1NSTXky+Xr5x
ws3D88EYxymdKgi8RAX64IW+yIgIqRVu+1O7eTRqjxxkXZN21j0pqaOpgGo+FKfNRRsA053ybPUc
DM2j/vdRr7rUGb90/RcAMHket2pzNKQmMd0dkFb2nWhfA5oqaFl9fMKRNmq96aX/VuWh9eRcC3jm
H3dzgTH1fUufnCA9a+RY6Zt5gQqpYhFLcNtfutC/9BQUuM9hK55wjEV+UrC6cHeK/pcBe5YXWF58
tP5Ki9TYOOjBMiX7B9QZGLgd8Ded3kZ1tVsPqy8WVD3TF4hFydZ6JswW6I6nQzWkFbUCIbwuUY5f
R93ov6W3G6WK7KMcFzSay+INymx4Z9s/QRJHUMzI05Y7BaizQMiOrY4HjfXyUT824FgxWP6Ykosz
pjCE8QGLfEgdfK3IVMiSqn0497ZO20qqQeImbaa2yNZpXKAz+uuykfV+sb9/8ptKoim59zeqjNNe
5oWhygLX/v2qoayiYygrWYzv5txKMtb682KDbDmFP+NYeIJFHHYBnaGJ7IRKtohCxn6q9w6rfErE
S0VqomRzy3q8cJCo3NgE2SLZ6Q1r/4mNmDuf0D1gQjFVkH0AY1Ia+X5x43aQr0PHwCpC619FXpVN
yXtSKmGh8uRY9ZV4nZSnKB1BAGIdgsIPXHfIvK/iw6WPMHWMmRElLeX+s+bzTECWXNJPvekevfkR
uFmnMIqMeioz95ybDqrFgup7P3Sq1ICF4ji6ez66Q+0GZBWUZCnPHG90AuUu9gaTr31fKFD8qX2e
b8bJPUgJae8PWMrOfbdJmChgrnx4kBPY0BQWQhC18bBoDOXw8ed2Jxlu6s0FjxeZn+LQSyXTQhfY
a1cJdqMo9O5X86lj9cNYY4oL0z7tQfHhpI3ABQF8uAastFZb+AAizw9DDBYNQkF5mTMgSHRBAq/b
QEl7mXxi0COgj3Wsgge3gDmK7HBUrQTWgb665L151kf2clBzhEBS+vx/n0lLlxKNOcFrTrUXk/aH
VsEZLlNLNpVUuf2nGWSBx2PRgbgERnvD6zhwuoX8wStYwmtWcbtZqm/5hq90Uu/ergEl09tj+Sde
oLr+sjim1p2UBudqLHPioO5GX4EUPToO5jd3sxgnt+A5bCYwvnLHsMPB3QgqJovokWo+rCq/XCHK
dzzFufAMC3csZCO0rQkv3y/7OXXvQtBE1wy+TPHt8tdsyuPfN/urqgVUJ5nqZxmosWs0l5woKS7X
yMhwtZ9FYkoi8j/kQUEhJOHGy87pCeGIOsWi59kj4SN+nQ7kbPVqMtRKNCZlonSb7gCeKwJFF0RT
patfA1WjUHBABwYTC8MJt9iwKCTaTSXhBtYoLpocnUU3oFQnkgU36JB+rlhE0XugFdTQebD+9FFz
OAZAaEMzWPaOLqaEdsnu8jYrBECFTt0J4ZIDdVbvTZ4W78KRWyy9WBl7eSjfPe9Dt/6wS6bcivcO
Z4A4R0APuFWPFXXnrU1ehdRhQATQrIzSqaJ2pInuwF8Nr41/6Pfn2dacpTk9IFNEg5SrteWt6han
Gxj6uYVWm/k28PqoeTawwDThJ/aH+KJZxtWOzN2iy8RJFMyFfO7jsIV5SIm7k95T4bWtJitZQyZb
qaKai/Bl+sYtnHhgN3TAsIkaIm78PC+//xM+xIb1+GWvLFPT3fmE+69jv2OqSi4+X9iVdrCgEyN8
TjEG18PuFCnV8XcJGzIM8EeIWRi3zfOvGPigcOKbckXPOtzV+paZ7DG4Iyl8GNraqo2zwwdqLWO2
LwbyoPP802bl9EkKiKPfpPmIGwj99JUYHfuCEde1WoZwfliNIvHFzMJdwltatsnDgd+kxQJt734G
NP5EOpojqtIHmnLh8M521tATWiiowR3F7rBnKxW0A6swzbtwz287lNg9Sry3/QyWWlP9aBHDa48r
m5nTwXtx7nrMVt6G09T+ymUES7Lwb9NBKhzsUlS57Z5eAs2U0OkJEg8F9wgw+ICnbmMYFMymjm6h
k/d478a3yD6Vf0a1DFIbF3aT3dv2UF97a20jRdYXD1if2EZ9g+S1PlTiFq85a1U7h4dF4dGmuw7i
cbTx1i5onIYMB6r8lfCykRiFOVG4RWUU0JrvquNCBW1fJRGny3xYp0nc0wq3gkry5plrAN0Yb340
bNx8SjxDne9rsBJQUU+jNTqLHZUjc9Mvv3WUOHIPxFRnwM9bfEM5IDbygUya/8cO57XGNgmEXe8S
s/dMRmr8qPZHxKtiad/G3714G12yR2QJaJzxPybUSLM47X7uc7WRVQ9JjyIEMAfHi7jOnMDUM4GL
MlCZ3JXK7bsq40vNoBmAC3Li0QkN2h9m/lMg0doFmjaH9DKHdBDCB3u+z3Jzaty29pFoUvGgnLWj
9OFghebGXP+2o0xUfNIAMRiOdpR9QiC71lCizjuGDOcFWeL/YDXnCT3UKj+13S67D4cCY15YBRmu
YT4m2olwxmYVpJnG+hbrhsNyY+RaySz0/8nSw/QhuX4hYlG9+Jfe8oLdZ9moxwv7zJmgJf1nW0V+
SodhulQvsk5Ns1W4G9EPKLXHzDAPcGilyQXfNFKPuS0ZyjfegcnKv8L+z4VuExqWEb8+G3PyHkn3
UC+RTSGujtDCF4FLxBC5deE+ytAnn9x6JiPrukz/bdWB/RbWoEHYvz0kuBLo8Fq4AO3+dvjpyAe5
yymGFZV4vIYTI+AXj+cJVH7kvru+OqUPkp2T4loczLqsB0piOSKnhgiAQaxIc4qh3xI86XN926Eg
y/eIxjXQdGeph3FNlzwkLdr/LbkfBI7w6wkM5xVvYXjPcdBdRotOtqP45nrp0qeIS0CP+upgnlve
E6NNXlzTeu3+nWjFAh0El1FpiHJkm2d0X/7k2+f522emtSO2dCvFs4/5GiTU3i116Rs/tjsTBb8X
p8Z0ZK4BHGzxnqf86BKnP0ix4i1vNQh/DGvzyizcesawmyhyTRB5/Od1QuXRdOqO5NxP4NMqDvNh
tOiI1iOMsTzz9hJrSQwWewtDzS1MFU5J5mcYJHRh7qmdRxBcCtqKVu/7TuqLtl3AfB39cKva2VZr
yH0+bfcVYxtFeIeYCfPiM5E156TK5w8ZY3PJ8xOEpzzCuUFP55IaGOUSVYXbsP2iAmXURfVcNJCU
sva0jUTuwfxfsAdDbFxb5dSc3Vf7WgcvWTYSBI+R1PLkujRSPYTdute7sYY35WQfA26uYf8H2QXZ
zhPtp6lBc8Z3WAGVcBSRo4TYGWgorHVZptYSoRDA0Gb61KAcFU0wr5TkQRBF8ej+gDt5RgsH18AL
Nd5UjQJsZqra6boCO2/YZNz6ZzrzLNqUmgWLLLKMoJJ/hbs6fBaJ+Ow5s1mDkNiHtHFlOzAWQ2ql
HiIGz+Az7ipwGQQYKXk4Wo9f/gllKav8CTbLUZ4Qad7KJ5eE1nzRKV3w1KhgXNbm6q2oDLMjl9KG
0P4HU3mdU0rWUc0c/QZIVEgUrOQmYa80ZEJpBZqpBls9m8DSBiyAQ9wqy362Qxm487AG6bUYG+Ut
PMPsWTWXl0BiMXfXpHr2DVZs4A3AT6q6xvB6LW4e8e+dNrU5Q1KA+gs5t1b4rVZmbI93827P9fh+
QQ9c2ehCFfcjwUuDiN+bB/edBhnNjtmTpblpc5gg5HK9GGdsw+tQRJfVnsf3trRCyM7LX5GTFj6L
rl3KPRStr56HbtBx7EPE0m+PvMqyLETieWckd6BxNbi7by/u17Ll7xo3mpAIcBaVJO08b6cB/LWA
FaICHSV0yb8vUYhpkekJn/B8WovSTCRMSnUsy059i+EPcapaVEKHbhp3JLSSYfez4Sk0BWWWEvLm
0s6afGMzRY30iL6lOFmGWwIfAxZDtvAuuOu66fHm5Y+P4XSRTATqowDBa8/4PY6qIa5cComzvegR
Eeo51qHRMuJoGdpdUsi6XXgcivBotmnC//3tfSgJTmv+CkRzvmjVkRqgZ8nBZ8syar3Q/nlC7Wwa
m02N5KToCAvpZfxxiVm0jPnRk0bSHEIUAMKn9pYFYLRQu/7XGzeGZJfYXOYeXs2zwxCkKh+1Qe5t
Gz3GtUq9zjM/WwgQ9xJZs7PkihhANRNsQgeF/1CsT9hpxWHDUHmY04cJ0Ia7tRUV48grE/7ATVMr
I55620gILrCvgau5fF/U5xOebZHKsMLAJP9lelJLA4wwnWALSU0XFc5MLRUOg3AKeHCj5bv3rqMF
wkGnklaHqfn3KYz5m6uGzsE9uyC4diMvCKGCBYCMVDsQ4gH8jF3JQHGmxjuWDVukPvkgKZpnSg5Q
QQJ8z4rCIsCHb1ubqLCsn5w8RUblTnBWyLZLWkFJZDoypIllecNB/lbVXSSG3MiARdUNMvagipup
O42Oa+hyUrS/ev8PKfQLiVaa+cAuRqgl/HUHJvyBwnpbso20sD/P/wwwHJJ2gZk+rzDHxbRSaTo3
KesdSRM9dObXX9sasjPTx0rvuIWclGjY2i39UPb11mFrVdasVna8THM2sg2yDrkJYr744fvLIijl
Ipddcmsrv/YuoJpl49hvQX46zth1YkZGpisB5l46hcLRVK8WJ9jxw+b6Mi2Hd484XiKnF0B7NG1r
RVEb68cESMMPknF1s4sRj+obrK15sGXWv0mCjlHCDd9wIfQmWGlO41HLzSIVI5FnVkJLsfTWEQqe
mAQ80MgkVrwggk05H1b2RxSa+U6NPzB9uIsgdCb/MXEGBMq+MzNvYyUU6GUScUS4QHUjZv4Mm/8K
8qSRxt3VQ4nLQCGpTSB0FsBS12HSguLjl2TCM5dMfN/a+1+dvhUMRwlQEwS4em3dBkjrJ6Ou0jj9
aRgRLX3BpZqgmhmK/LOC9/92fclFNXhrXH1j9wQIzEGpow18ferVtqXMq0aUgvQ4dxRWqy/XBnTK
ddZkQ/TY/qFpS6ll9Y5D3jB9P6MGbDb1wnsgjW0x0bcuVdfcNevrI1B0l7i6GpJ6aqg5urb4Ekq9
xWsfuzfigHm6sYl0XgyvTyfHFR+yVDnDE26RhKeu5tbN8tLqzBJBu71cIxwBGiJCnmXVZhWTiK+9
C4ch5jx1DzDHPiViaApfyV7ruHLtt1Nqw7Xs+g2YiaYxQ2+m7BBzTiOPlnfHAnE1AimJS7f7w9Ab
zSSbCnx/mExAhpApdWTfEFra0Wd05clD6x1bDNh0Kq6TPDs7evPzbhQQZaMk40/Hn6RWNpV039jN
tRhTNqX12792S4hA/ku4z54BB3EDFz3IlbsKZHq8Vlmp4Zo2iV2cw47wSkWybYp3d4eMzLT9fyBG
IZe2gXnRtEt8WAxIWIPW0SH7O5WJI7AbxQYiucnfHZTRbTsCuGahFqewdsHh+qtST9ooJr+3uqzH
VzMLR6T1jz0cdtd2gTFHvl6/tvQ9t1i2cn6mfWYyQpNVdZq+5+3dG61SZu7Nc4mrd64wavtAkmSO
vKDrFwbYhbVNZzO0iY4JHbpjKKeBAP/+NUwrpPUtztP8UI2Lko/giE/XbUA1kvmTkCJaiW7nz+xI
Inx27FL7skXSb/POQ/pgU4DlCoU/FBIdgZ1BF46+Ja00JgX3NOuYkIPf1i6SPGPt4C0iCFuPR2vp
5MVIBZKamxV7CSHP9nYC8HbtCX+sGeI5TVQCObXaqM+B/D9YmDG/hG/dnDhL2CLCH+mugABUSZM4
yn3CdL7CEUojlxAe0qGoynqygd8pAIIJ2bgwHXt7xwm+LBgTAAhJ3a7Haeuxl6XKkicrXbbVxnAU
KrdFlLT60hnkXXYu2FmLysp7q4siUqqbm1Ics66HFGKycnF+Mi+/EIxztoNP6O0qZF8E1bAg45pA
yJdoxrlnC/COVf1F/tXqhb4eygRvWVxrjVqxMH6vNpGTdyMpuZPs/l24JnmgdlVCD8t+n/VuKF/L
4AxAk5pAZal0qgH9n6HKGPemviUUG+w7buJmUCGcDFsuNiG184V/WcFvEkEDI67Qx2il+amQ/Bec
hkTccjWQXelzXb6FTqc4bgpEb3+U6737JyalSp7iBv7WMym5i3pfkozPUYodbL1815AgviEo/syl
3sOsHC0z8i0E8NqGUlR9U46s0tV1a4jYQ5TXFuYbDGDUwrqhXS/dgAemHQpt8IusPpcZgLpz1M0y
kI6dmuxdbnv9OlVc5Uks2ssVh2X+/QZf/kRuq+aAZCAAdqdxQsgHNMQ9f9XSHaAJ9MVhxXcO5SkA
4YAC0JHpbkxr1kI7E8Lbjd+uJvhVJRunojF9BYEwq99jQz9qse24oGvTeNhByBKGMS3HmvOI8cNm
5u6mUpBsDBL2n0Ogpab2E05JuC7oEJb7lhiJfUiy2+OjbuD4HpIxpMPFQ/bVfgBIn5ISCFiuhCBx
uE7eUfjtF6dm5UnNzjpmJY7nfwKmiLyQ5nGxEVv3P5aT2Dxk51n1cXqAi3KYAsMShg9eG6eYZNyw
WfyfcDkOx2Sx5eei8h54m91MBGOcNM014tKYJtFP6XsBJYBnPhK6MeXyT0SyqVttUo2ugrNfeSf2
yGot6dvsh1stoxhHJQ6YNk80zOhAbOBalXVX4HW7M4r6DkuC7qxWIPKFx+qGZp9+X8VcuLUknfrx
NtSmVyH4x9c6uX+ohSLc5Lt6evFalR09uDCITBTxkdomrI6DhvrjDKjRo9o0O4wyX5d+spXDDZjV
+CyVukaSHWMCosQB/w4MhlFND9LGRJz1JAuBnpwPvVbUTOKPDmSRBFts2iLf2xRlBvWZRMjvF66O
t4xlSSmDOH9LQLC7yb1nKNZQ9yOt9XTAvd0KS0RxVU9FRsPzA7CddP/nX+NcUvn3iaKR2pgsYk3J
Hvp7R3TqYLL8WqLZIxQAD/omOAs7yvNlKFkaDfc4P1i7xX41zwi8lbzsYxeVGL2OKfKPI78C1t4o
aY/PbcmFzEPiJnPgMaTajEBlWcuj6C5mYuv3xetND5/YK5zzNxbxfokQNG7VpTdRHall6I3Lv6X7
4r6+l29lOua4IOSnpGzehuKgvve6bpZQCe+STDBQsE2uXqVXRkbg0HyN/vhig385GWRrp3bOjViQ
pXb9V993/l99VdNWLdJKZ5UmpLEz9eq7PG85efxWPqEhhH9HvzzDoV+NOcvosS04Kx7doRj2z6g6
TRTO/LjLQxc7Vz1z/M+gvnyCCxKjFQ5gJyn+AzZUhkffEpOattIGoeUP79XA1dyzIdzetbbZ0SJL
rFev6om+FTG+kR2h3UHzeZLguzIN7aVA9Xwlg0tcEw+cWTet8PzWb/m1Sx2EBVVLOH3wNAurr3i7
huTD3gYjwgSsnV17KLgZQo9Q5XqfN4bzwrknO4O3r0Zyj3vD2hXJJFsJxYFi/1htNdF80qR2UJfx
m76A8aKERsM4ssEhCnMdhDISRLloZSBPa7RfwcTq1dldmjyVqUgIddeivlpYZw1RenSmdEABZBCw
qHaQfoTwLBUbGilLyq2zWOU66Gn2pj6zE84eyacKBzFw3NW8QNj4LhsZSceUBR0GfMV+6mMD9iyr
ucaKRfU7nDKGYPzbfRqUiD7HbDheZW6aKD1gEM7VVu40sZ26HzO6uO5FVRF6/qXZIwHSPN8wnPZv
D+y1556vRjOeyFPHJtdqX7hR+agaGjbRGi/s+2+laCxoW00zzyhwIA5Hzq5l+R2Myul3kMKBoOBl
Th0kDpFeqbe//3OTjEaCMvihPzEa+65dcdUTJsogtcteGOZq6CiyoBLJHLRYV3IfyQm7n1isk3Mh
ARd1xBPrwFnpXOP0Fpx3biI+oDw/Sbr5NBfpEg+ct23Z70x0MsyYtTZ++T7Zkym34I3CYTv8Z3YJ
Q/I6SornGAmdafQsC6U8a56FowZrNVLuGhTCm1brIc81ls+DmsBUwNF/gCpy3DNbrY7QYZnipYve
RHElL1Htrd7ggdq3QPQ1dc6Z6oCkzczac2MZ7IrJTQ8Tn+elGXPiIUK3aQ4tOaZ3NLKwAtLhUCB+
OIFQSiI06UwqFhfrtYq4Z3B0NrVxTCRrgzBT4YJO4DcOzpyCLODl0iJQyfXWY8ZYZyfgVNnwSwF3
5lAVzbd0SUilI4/WeS3ewW0UGlL4FAlyio+IC8qHYFTaFTKQNZTzmkNdbngh89NQzrP0qlUcrwZq
hfh+Re6AjgqU39FB10UtCqGKb6ZnHjB+Wq+Eaur3rxV95zZReE645uZcv0Fd65DJaS6h6T5+6Zoi
4e11j2u9WuFdB9/j8nwE/Jc5cvdO/3XIhST2HU3FTmZb8djqbk9qvbP55hrGiTwab74ZiLSXUSyo
4m9mpEqvBTbCzait3leIsNZcw1DqvuIqmvvEr1CgylBhVRMlnjbZfx0FqjcrO4bnF3p+AoQX4qt0
gEW37IKa9bA7XuVoUJl8FMYFDf5i6vL9fCY6fCn44+BTBMbDqTIq5uKsZatWXzLYRbs9Q18bQc/Q
odYYptQg3OBZPFN8Cji0RfFyugHZveGFzug10vBc+5yHddqc5unlJMoYr/ztGW6RLvtXrNAuBlCV
V6Vd/XWknjlR3Rfo8k06UMexE/iZX3rwZL3RpySujOhVz+ys1ZWiZlSEWRE7SJBCDdVWBOprWemq
SZhHg3BNMTDu425vSSb1N22cJSCCSKwVeAr0E/ICwozYofGHi2LMg0OnUdC4eyTXilf5mL0g+Qgh
j0+yLfHCqPcaGqmMCHIc5sXyWMtUBZjBNzGqiI3GdPW/LzNdU6mFAqhxICbv3pmmEOOqNumJokoJ
+AhUDGf6g9ifKTmas3vxEugmZFZR4/WHQShKzXx46lYLr8Lb0gN3Mbi1cKCCNM7wpWB7LW0eGG8M
errgp+ZrpL1HjXt+Cm1nscMjdDZb7BBdPelbZk1AFnaQT2IbxWFNILHAIlydRKqUN1T67KkKJGHZ
duFPetyj2qMRuIlW2YFL0GvYhDDnBYoau5m+gagFQAvxJA2Ac6WCIVqhJHecIFS3bSlRc98bbRKQ
w4sFJ8KB3n/CN5pq4FzdyA/LgRzFYRtku2REABmPzs15MrnuIaNEM6XKmoGENy/VS1pRnpS+aVNo
V8yrVqdhZFlhkYiTh/QHegln4YKI80dl4UJEL42KUN7TPkncDFU0hUwqutY3Lr35DsM96oyUWxBz
MB16x3WZ/tM37mZuD/1I+yqVlWOASlKaFmti+LUYYyCxgZMTAj9umBOStOEjjHgS4ZZg3FVc8RnF
XEVYYZnFwkqhRpfGtoQIg4GhY/Evm1XAEGMzUdZMGNCyurQ/gknoCmXxFFLOuPQ7TXZjjzMlFgDM
OoCu91Xm6Tzv2Vb/bwR29hiDtE3/jCWBkjEzgN7/OuEsMwN3CDdtOZ731VaV5VyY6LpxirZXAtz+
+dFBFgCQRExGy6emIHhX2lFsZxHPqTQoqiIN4XR9jAN+eK+9JvXnFbAwCW/Kt3knqc2sPNzHDR9d
PWxYfjae5a0A5J/cl/Z3jk7RBB9l/ao8dqBdem8+aU8fx/g2xOHzlmYOHKJqKys+oEg1r3TfjC1Z
KoAka2gbel8jM/Pxb3zAO4VxzOpd8w0zzXuFRikDowsIgGjQgWlZLWEWDIV5N4KXxoqf3JTKSqi9
0MpDgx3qVsu29rGKP10VSKqKCf0e7XAUZxkNTGLY4nib/VNSxT1jfha7BWLCtO6o67ikDGpSI9Fm
wwjdqizX0M1OEm4T7Uz0gLdE774dckWxVMCmh2cAxK1FRCLzGDzVaKPuL0OiKepzErYl1O+5ro6A
UqkqToHg/vN40BReJCV+aFXAvDkmUcBTZBSFBTygif5nd8vsz7onWx0+gvDD2Um78t3h+o94uRgG
iiCSAxkvBokgjasv8s/L7H4xKSukS6GbUxNlkRpwQcI838KO5zVjFrFgA5f2TlacSr1Q6f3ZaYUh
RdpGuZvT+zGfsFof7GYtmzXMfPpQrovmLA75oS0/4i7fw+05O6QFqNG/xfcfn9PUxJ15VjY5KlJI
vLhkJhXNUMdLp1kh1mt5na2W5HhAb2eLLseBMpQDw0/czkym5CG5tPM3gZYoB5MZEPLCMUa/H4n/
WSVW+SeRlYgQRtn9oRzzb38wjjaEDkKBWv0EtQk9bXhbDQEWu8+jLPKVYUHxijBV6Z0Z9N6Biu23
d7wyfUr9kA9mqpfMhNTzT7VcUyZ4ShYcsHDsZL2RhzvMTEZ/6qqwHb8wY8H93bo5RNe7VmpWR8EA
dnYqYwgKmGmfNuTVDskEV2kI5rDYY0Vb0XB3M4pNSuZ4LP8JtoRqSNJvtfMgMBTGBcnvVHVDapRV
LvIctsMIfmD+M61t23wcf5ssKO7QZx+Vr7UM0VGwTBY+8NwEz+fBBJzjwkMdT5PAierWZUGbfyvq
2Wh4shSf7ymDSEtoI9EoacMpjG3/kcvR85mbR8Bcxe6oxz5Z5rS6UUsCrQq1S3z3pMKaW6W4YxnI
qlc4+YElSJYsFuA0/4+eMOI2hBgNlFDX70Uq1pESEXnWDMOfqoKmMQ+fL7XyKBLyykUe5AFs3/RW
LxCSdXmdO+Lo0A/rHeIOnvatr/S2GhUjroa2cmdzP3uzMxGpf3Q5SYcX3QtYvvpqOpTEVIq9GKbo
iCcfBKzURwqdlNVSOh6GW/UdOrEgV/PpGNvtzG2Cd8apg5+E6Fqhy5TC+HBI2uykYjua2AN14NZK
lLein5wGGyLX6S20njGK4PROSXQqlwEyjC9yjCsvHsZIRzJm6cHLfMXNsxdaobDr9ORa1zsqMpnd
akjmwc/h3LBLWz+XL9vzV9AYgoaujbxKCSjhFayovkbCQwnZpYOgb8J6VeXeq+b8VcR2DUIlDTAE
2xKREEXv0+4aLxpH345MR1PP2FgGo3rtkdT2byhUXXDneCxPDYh4Qzsmnbtb0VpsZZ3ZA2ramcMY
OYFBUD+DWuAH1OVZsPbuwQDa63nZ1jlhQK07Z/yUPDGBOb5Y1nzlpUOPKCK5K/8FlkYSNMZypR7S
0PsXYjXnh4bBnGN2XIEElB0jTLtoq4DbnVLtjOXJH3Nc6xtUP4nGkHVldKGmhDdH3mbg/u3xhAI/
5fwMy9XzzCXE8CPOapc8J00uHTlSY4jViwsIOqZ7dnE/Byktric/VuHQoAYdZ9bysi2uitjKzFQS
TABQdSD444SAylTmM0o3G+w10yOqHB4rahcPjmov0HUTw8kRpwdqV95XDWWIMCXwqlkatjhaj9lT
f7hYPc7dMUUzOY3f8otk/RX9bEnNBeBqgH40vqo2MaejTUWOf9El3efAOBfw+ugq04VaWWb32A8Z
0y0XfGjnO+unB39wSFlsf9l7iU76PmGmnBa5tyvaHcAqxDnGNm8uTOSIHM9mkB7cAeorvECT8znz
+T0AJrxH89w+QJVXDGYoZ/pTwT7au/A/nFmM2tsTwpda2BfTBJxkzvMylWJbiiakcVR1ktCcVVDp
Tn960QL23+iRR+QkhkCPby0k9ssLow+xVpkym0VYwPMl1q+SXjnYhO6IRuiLKKVh3LehjrADMfqz
iwbIAHPzDRjeveefcwI/mF+ZuFlIvO4VQzDzdxrG/mItHs/hECrk5auxNKJ/0s2Z6qD0sFuljXQI
kycJrOx6AvqeWZ0BNQnLb6DJqtEkOFWXVWAwsWWOs04e2cG/gpNc+EUtrAdVg3Up/G4FYCxKsjfV
GqwNAB7abEb5pKHHXTPvLgwK8mr6FKbwjzJRkh0HoipeeP9CQ66Y+3NB72o3ft5P78OUVKO8X9PW
VAP6v0+1tPLhCZ1RGRnPSD6+NhmUXZz0ueBgbL9U5/PXbvsskkB0Hg8wv9gBA6Q6L19DXglDeyrL
+vhQK71m8quhAe7hAZFz8rYag3xG2w5bbV0gtThTz+0bhrdx6Y9/urKxye/qml9UMQhv5NByS7Xt
VssFSfZGbCtBLguFRwO6Bf+oCNYoAjEqVgMA96Kas6CQNh81WJRqNhN3Xn/HFJZxEIDwyGp0pWXM
PffwSKVttULU3+vozRjxoy+cOIqBYQkIvNXiiDSjcOJYmFufaRG5lOJlvm23VcKTwkRNVO18ntKi
JAt2s9Wdm/tFp4XRVN/MNXnwFtQS72oXT850g7+YIvMtJiK9rIINDmdxO1/WsdEXZAaG0nWdniMZ
9g0gKhsLZCaDFDk08cA++vomnkx81grhizhgc5Gy3wSgc5FHRI7QWtZ10wAq21ftJllostdwJybv
7vRCk9MkMKvy0XNVo78boFM5uSBr5+fAH+KwOCy4i9tlzQHT+lF+0m/CepCohoo3geYOT+qshnkw
Tle67FzilhHFLULBA7620zI2bXLozg8oy8wV9hNfJfL8nuhLj8czm3aPiwjPAaT6yY0PJqmb6ED0
hxQh15VVhmEfS8ALLN0Zwcdn/n+0X2QrBuUOf/1VOOjDJ0cG89Jrv7Pol/7TUMINH2IpyiyxSRTC
HKclyG9YG0PIEnrof/Exncz+M9yCPji78/SVIsSuY3Vwf6PTqILpQl81sedpiK/i2oH04VlYREIb
1HwIhOWJoNGFQsDy6RLswWj47i6Y9jNGyVsxGki+n+kf1/d/EwGJrZwXmw3Lmj/mD7MF627o7+p4
Y0EB+z/AhA30T69oIhS9xQqHKsOXL288R0FIAGM+1+Cibgaa1O8vu3qKvj13Af5FtFx48OB7+eQ4
68hbIww9tSroGHspaiQ91b1FOViwukF5cwldkhk1AQBa2Bq24h1Qtuww3ZFsgx4hzC1c+9kSsY/5
mHRqGVGYEiO3KbJwr/4g4ZTjvxjoE5dztx5TbWJHaejmEYEksgzJ2U/YRFDDe/D1Y1EfdiRQsrgX
b0Oj1Qu3SLq0d2zoYlXiL+4oWFiib3ZjNjhWGwbRvoUB/+lO1xExJLKiO6jxW1UAWISJRJBuVHDv
Ve6XqpIudsa5dgs4jMxNNgaWcADHyF6z/pXL3sS8Kln+wWqmv5tfyjiEGbXNtXoD98kKdR+1dc30
hRf2dHUb85Ux1HiGKGINoHS6s2tDp29HV8lq4UlTJX4yhC1vG4w+xV/LHAH0oMmDTA6GTpzdeL4Q
eo5gKZOmvyH96YyKEgYge3pqIJg2VKZ31GNjWimmo/ZByVg/qXK64SPVAUQMP7LcxS6DLuL9PrEe
C62nGu76hWG3RB1A3VcnQa6Wi4LIwYxX6OHdqZFeNcLjhW9K02WTBDJ0ivsv+zNZiXNWp5EQ/vJ0
N+qZjw04E19/sjAsKiTnLtTnuF/06N6475dpi+x54FkT8gpoetERTnTzu0dvYbXF0m9WJg7AnFlA
uciJOfA+LQh6ROpiZ/IF3nZTrYuB5Bd4thOMrqJFQvlpoSeVAAmmPxR4QxXlkAlz3GtZvOOx701P
uWDT/V5MCY3JcTo31dfYG6JQUk5KhKI+vkkZb2UnTwCSgrOhjAc3JP6llSnhMdPSEq9U16sr9UQq
kX+yxB+A3PpzFUhbfiaEmjxuyFlXQJC4gL+B2ffv4zunx7lna+Im1d42MRtN9hDeXd8EZePcPb6w
tHS+pWE0kPe7dLJARzct46u7tSfSDPB2teH9sm708GrHOTMQngIgKTO4w1tWnboAwo9WlMk5VW47
P8i3/cGClqovTHDNZf6QfIjjW3NyiYQv2DrEyUQK+mWnupUT0Jsle5983Ak559ShyuWvFU3m36xD
ixHTjXq9lwmz2O9Oa+klMqL42k++pI+KagMUF4uEQ5niVRsTZEmW+q1cBxFxyOCKpYZdVnCmZz9L
e1AeySXRc4bpV6S+SWm5CY21tUdYeU194LXxL8ITJKMRtiBxsTLTTf+qBMAI9qZxKgxh+bCMLXcZ
MwspGUvJVz2U+8SwBN6LCT3+BcSrEqhjWGg1Bv5h28iHLRqdWuGpKS4voUQN6eNU1+7FMinSqqOs
hdhubziZpDqPW5L2uNt4WUDz/Ygpr5Nexpp6LfEzNxJu9cqQQfuJdrdQ1Aog5vaYMKzQjvNfFXm6
enA53LbB3iI/wIrcp+Dy3UIne2fq+qWGg+JOKWqHx66KfAwQTro/icaeTk869SXNvdb3MVl/3atq
lXPLrBuL1Qg2dmuzuEUQoN4M9do/ZmVT+SDPks2RMUglXBp3RfancgtcxkB3oJu7rDJYL6QD3SrN
zl7wJNFEwPoj1LCFOUOrD6c7GOKnN2EPxdxyDH8jHrg/JfzWR/LH6Uiyv5ipZlRjoqu/q70qysoc
sgy1nPFsqee6a0TS9M8NMX+yOkNk7LNo6Y3AwQWUwj+1glw8heTTAu+0gUn3vXKZkyGaIPSVDLvp
E54UpOliZeN4io+HzldL/z78he9HP+/60nB17sGgGMdaLQhSIG1GKBJ+rIEGAjbEVvapuHerwzWE
8IkrqmnsodvMvKJv/cVyEldOrcQHhRw9PGp+qH74a/vOBdvLb0cH49rSxdKFWthZAud80EOKJFs4
cqHIJOm7D6zT9rlISo/ifdTtl5YbgbRgMq6ALDYJi/eIdEnM5++F7/VMZt2yzQQCnlBkVbxn5bSl
o98xId1o4yVEOXuhrtAT0lDiNGpuxD+nBgPvjrSifs8+hUOHxlMMEHBhft9b7MdfgGGjJtHguc4i
vcjaLGCS5XVw0Z3ddTx2Q8lKp6SDgMC7FwE4oayCH+svlk/zRZYD7WMvrchib1R7RK9YSIc1Fdb+
nhWkD67Q3OKRatWhGXeK3m4zw0GDOHu2tKE+JWlOdLT9P96h5GRUWeej1H4rzzLgQoyB9GYhC7Ek
Bpg+URcnwd+oTsA5DkuxwjYEY6JZBIVrFyjSGmNyJYhdv92yuaskQDakR8vStWcnHpe7yAhUTl7p
2Lt2NTNa0nqB5Ib/KF8eTHFmgXejR4V1upv8BG8J3Dox7Cs2xmv9vOo8az0/OqxwugWG7QyHbcpQ
Buvn666xm27TXUPZKfuXVgFjTurHr+U9g0L5ioxg3XoT9hzZ2pIx0YjKNoW88Mf650SstTrIY/AZ
9/lJXDSjI4OXUcqZCZrjam3tZilClO/kEviOxNF6WEXSpChRn6RMrHSoaUGtkZ1A5eX9wPpC3R5N
czMuo7XwJiXvpdaDMghRW3pQ5rh8jjNF4Z/Q4IM1amSWsSTIM1bMnhlEieYi9y87khtlQ5dKtoyw
N+78vyidK4DFqBz69SGlGSw2FhxkDhTLeF6aIESgpTHwkAQmhvU4y4u+1A+wZxNLuU9S5tq2O83N
vaejwHiqReH+RVGMRwtCNwyJvo98/Y5hs24dyW67PBKmY3BDQVWM58ryJjO6u3+NGbr/OLIVEH2l
LdOzaQaKgqNI0O3Th8gPC/4KzglUsmWPMoIyLc6RDSLxQjAznSYJtkMn+NrxjbDWiwYBgpBB73yp
Fi+qZnsJ/JPwmtuBiZBWmgHgkAqqlQFWMCR/4bpZ3NzH1vNyl+kW4k8nhml9Db0uLkeyP/Qyf8Zk
VzqwqUz8uX5rDjUjnMVlPkGr3TTRcf5Q0YliHLbAq6HjCSebIdNXY6rgUdht4NEVT6Ji/uTmzx+z
faR5+3H2CxTRcIEDP8PlBmuIikjr3gjGlwQVNu3I2EgTqHwRrvVNE9i60r8Li7+z4PyDc3RcPuUa
JBPg/N8gcMg8/yNmgpszKbEo0Pk+Tz76j6VV0qmWT4y3bQpiuxZPqTIc7yGTr/7qeDI0z8qsTZHR
JF46asod4pKyBG3FoQer6gOFIk5mzhBVjkhOoq1CjGOHw74/zSQIkio/LmiSne/Rsl0a/crQc/Qf
ca6DzLFZS5Cbe6waxD9A0slMTne4nP1u2siA4+ZeQDzQFoFqs5XUKVFUpKFl34HO/E1COTO3EkWH
AqPMRsVOlpSSxSJJOWlBdQIxFir8cjT7/FloCZGwg+mxaEGAwgCE8Cbjj60EY3e+HPpWDpk5m5TD
7XVBnbn8JsQt7WXJzlt3E7Cs+eI8pPlK/A5ZMLBYWKnSKCNF0ndB8K0BrWc5l2I7PPdPDtgck2V0
bLqs7oCC3AYiyNYEMIL7TgiezOjtj4vw4MZ2BM5RlKfGBMlmZJnbtLUSuJCZw84lBx1erPOS+ixb
nnztmEB2NF0l8lvERlToO5IGBeaWaXv5RvR92MKuNWTrebqXc4Ekh847850GUY7fiHn5vQ8zoFQ9
B9Op75s2eciKJpLiKgrq7v7xsZJWtcD7xg8HNLyg0GMO+hvStsi7E+ep5ILUynhBvT/BtF+YKi/j
k6MRtBzo7LxUwGCDvgEQAFqdCPgEwUqBxRXrukC0PTGKb+wYwmZUyHZBx5KDeIHdhb9x15MJi/wj
ErrXsBOji1goppT1JqGsekYnR6o3NW17bYSlsX0KA5Na74eT3iYJM0YNWns67n2jxF1jxPwVtziK
zbx6reFU4IvyigiJhvLAEEQ87iq29JfL5M433YlnQAjG8SogNVEbzdSXS7EfY5VP6sWMMuIXYZJK
EzoMF9t6vP+iyIGLF0ifUoJ7v7xtHN+OMUCS86B2UaKUw4auHdTpqMbWBkcRmLuK+qzuZVVmsKBd
9PZL7PS0j9nCVzbyrEwkZE3BLPSRfVUiaLuWUXUwrZimvIsxnLeonzIDed6pj1gPoScmjUFMj1ac
Z6VT9UIpap/GSJEsYVcYD4kaSGo6u8NVFeDDMl+rS1p3PELYr+boIfRZbV/bHmKLI7KrVoIRDk3x
vY+tyEkfFG72gRH8gouSh33L7ryIZj0cjU32B1yEk7tgmStKKzZYV54q3PB9FBk6xgMYe4D1Ihlc
Ai39jWj1mKfJe3vVK6NUcUVAF4YS4ZettoyZNXE9ab/xnXe7josjQS4DBsnq7FgLzS5vYRHsn9mg
LHA/PXd9sGFKOBa1YNycYn6a0ad4Nptrq2KfqBf1BqaLv9VykITC5Lu0dhbFIacZxtIZwyuGhF3M
ZRsSU0NF1tzUtoMnz4Mbiy/fjw1fyluLaaopzRlGTksJLfJGg9WVr2u1bnUVMDx9h0G/nOiKZiyT
sZCRm+KJxzZ61WR4UvvAGZHZ/sLWJ7TYhFWTeinRIZ4OmmbZ+pOxcSUr3tLP5wxB5XPBExdgBHO3
eFJ7bDDwM9MW2YjbB7gR3jcydO9gO1IvrIlDIwZciz3MNHNADqy2NxZz+qC+UJvkAmr7S7PWDIpt
0KZBau5h9MX90u+kr4oh3Z3LMvjr+oV7Su2opyoMTNoeKLqCHyI0oySKdA6VwmeQVugxGNqe8NE2
O1uIyQDZM7ZePpGNHcVnj+5YdKK9t7bugQGSNcqZOUB3lt4tfpz1VOVMItgA8kQ+ZpeG+DYMmDJF
PaTm/Ux2kRL5RPjfnKoxc0U7dwCcq8Lt3gz9+KtwXgRcRmaWf2OB3fzXy7BmMnltvyFbEUE3irpE
wAT14EXyNnbf1SIASKKsOVS6rA+RiEfJP+vJKbkkTmO2iXVKHbqukCvuKr49C9c/AjreXbLLVF3p
8VcWLiejugIJLw/WlWYoJnllS8W8E0egAKZMGnPMqatyUTLThHULr842nTuxdVCi8Zvlo0VtgA+k
+j08GQdmoMEhp/2G7mouHJDvPZNkV1lgyKHgUXWNRz6WSWEsqt9Q/CnYFrI+PUnlPUVkCyVReXSf
MaZTdugFRyYZqNIJs6ZsW5ZXHtwV00ekODUTaV1EhtDFLT69c0Jw/3+gueo0MoBxd142pIXtVi24
h2DNM4wrv+tjPfzEBchkftq34ptMSEp01D02iwFbMr8awpQSQLcQ81lJGSW1jrwr8Ecq8DU/WHWK
hYoxLIHUos8XbxxxpjQ7ihZoDN39ZG+gSVpvldR8DQ/p9JDeYhzQhIQi38Uwg7HM4NrVexaMuTLQ
/3JUY0Ch0p9MvXYC3JdB/K/eyYYVxsSkaxbcJ+Mdo/KC7cUMbUevq+XTEhaM5OP4CTn5dvSyGMpB
8P1PzaVdYlO+6Fe9mrgDdDeiX6j9sN4XM42vEXQuZ0qgRnuzu/dcs5PyKTWlLI3LjXJDzrMi2JRv
1PHZ5JHAVv6OfvxN4KmC4UEC0hrmqwZb0voULcJd7zNY63BF4fUMudhz0oFmLVG1EVmzdZziQOZf
uPkGPk9MBgmxO3pVGN7+sE8RiDErwJIjOYCpueSHPeCvM1XV3yhJnjUEV7wzZR2Paw/ApdXvcfRj
UgnlRUMW3NcEJLF/slcIEADgytajjLslgrgPyqVtXCOa4OiLPYUnWt2ghuATQoG/Zyo3ujC8sz42
VhMkiiIYeQyaoaoCMsj7yUtBLXbUJqFknu75pIgwV2AdmmAOfkV0DBJIY6sBhiHm87f9jRu0DrGX
A4KgbGj5U/5oXg0fBFPR396QJ6v4ZxMIjn1Uer1kMD2GuiTCkbFd66Q8gtYNL9d5gTmT6BNji/mn
eSAxiRq/9zULb/yOvXR5OnL2RTskL6+mig3RReN3wk5kw6SWG/zO0Dcyk7t2fDLEjOvhSFRKFyfH
hweSLOagvwUyGxLElJZLLUUFJq1p7DDJoFaN9sKCJBuhSMPWk3of2Yw+di5jgrShWVqtfvYyrpr8
T15ECGPwvjaEtLK7OsYqeDe0sSzk5skwHX7hGKvVWUZP6G/uCvqrJWAy4NPc1ih988Yy6MnNCJf9
ELyjTBe/G5s+T6Oy7230f8kSBwMngReAjrrM+0b0HCxamZS/8hPFOxJ/t0XdC7znByR3mGu3W0Ra
+Cz7JqKsDjbNyjytC0wIxNgQdtZuShhbQYMliY2fp6wUbpayaPjxJ/7K+jwUID90tgQi3iylUW/r
0QA9TQtRR11zOywAZmUa4j7oJeQEcwQdKyY/kx89KWtTeuNi4+yyZZYLfUIE+K+Ml8OUPhmP+eBZ
h/S6gUrg5ltw3JfIW6yHZnN9s1Fae2JN9ng9YRZOTzpW3uVAgbEZ/AqBf6CV/Zikt8XPtwFpaz8U
W9Gb3JQCNckEItM5f474EsdywolH2m0igcJ7lxMsIOnybAvD61N1WNA/XDxP+HblGT0Y0JUegt2a
H/HGeQMlq+X2jhdxs6mNCLqohAu28GmLxujIJJ04CTsdRr1mhVDx+HLfPdHDvQ7AbJMQi5jjfVPK
TDCH6swG1yAA8bjWKLbAbICZ5uYaeR3ZOx2bo7Ey4AzubH5MTAX3y+evRKE2UEtwfFWhnwX4snRH
AzknZCF7Nr3R/zkjXxGp7e2iIImEo5BCHRChAOsxPu7KzQ+lvlc5XvfUxu7h1VBImwO4fhRoVsi+
Uy+jQGWGZKnTsr4brWMs/A4vNq1MKAHZcMxaAdnCz7Y0CQmTauaMjLgDbKRV7fUNQJhvPhPZ/hKh
KLINEYApajAxvmpFN7wCQOIOt7YOzEHppgiRF84VxBslxGzKUfjBvMwDvNCZAIVjOQdmNOIjjLKP
0LKKJ/vhvI68Pa9TVlriN4G0wWBA06FLEThfgDgtMC2sd2nCQF2lS5dCmmtbTrc2YGBu8L76g8W9
JGv2BsPshY4FC11zbr/JQs1fMiURYo4ePwOBFXc58Acn0ycTxd3FOVaarPI6VXxNqNidcYJxdReF
5ZZC+uVGNyXANPnm6pG8wcd4tTMu5x0wU8c61IXSxegUZA0FaX3aLhZ/rHzz7Z5qmpEZPGs9p8Bb
FYbmbfFnGXdgf31EL2nu6FcAjAPywiZU0kbPq+nJNlsvWIeLY4MccIWcwi8dS51nmRQx7jGYSEBE
ZHzI3wZwtCzotXGSSQdJ3h1T1pY66c4x8Ezs3zRMnWaBm/NM6HcfwSfpkS89Nl8PmQxyYX4T40O7
q44pjOqu+1MSLNs0F0QJ1VHPHHiQRvd9sFjXezIU5z0TaRsC3fgwVCuOcMHskgnemAFivhZjn5uY
MXo8nG1bVIgOoq0GU/b4WJOhKYEA9Bm4A9Jzieo2SMLT4Kg1d5PPLT7Db25v+IF7RXJjC6jWfIjN
8b7Lycg2X/rdiu6CHvBuX3HX2s+DNBJloTEvvmfo8ufAl1SeLlUZQiYqXakqLqLdO8oPawzt3z/L
jwENk6LJmCdB8tlS1IPPCi41TjKUk0kiJSJbNbxTS2wUFtihvmyqBb4JhnpE19Zr2yc9U2550FuW
bf5FLdbcMY1AaL/+UxsVAv/fuxyIKHi9Bh2RleARRtVIgM2/ukl2UQSpeS/x73h1B25UBtGUN2T7
qtowCKXJk5Ob3thZyBcu/C2tnc7GXEHg7eJgCesLgHhM3Nv6CiFKOA5oMn9Uu9yUx7vKA8VCvWWn
4FXY/W4/ifnV5GU4gDzLZTgMG14TFQmQcs44aYSgQeB0gF9dtY80R/qkhW1/TIslfgwbz2GJWVWs
tFsOeyFU9O/u+3XKB9vD4JGju+++1gd+50KZXQhbZHJXzYhLL3l9GtD+tG8CHj8E5WqpyAsyajJa
79to633hUqUkliwiee4vXfEHq363KxcOJLhOaGFL9z6D40r2SDI61mLSuBIFsDCfeajaB41QFX0R
vgOWVwEjPUemRehB/82Xr8iY/V7Do/O2cILzbEdkAIjxwqSuZ9qwnHBZop53q3XxlB/8hEdntzgu
U7v2t7gCh82XOLNG8nTEU2QIBPu+pD+Ga1M77t3Jc4zIQCL1zAWRaSAk6bxFTGGMjNunvZtUzniI
eRUgl4RY9Rqy+jCAqp1DGEuk3RbT30W/T0fUnDa3WqLP9/AdBxSF6IU7q8/4zU1lML8uSGRneYmN
ZyGZnaorOgoFpsTDBWKP/XW3VCEn5903J44l1h3R8geVT2qNQOfkC/swXxeNb55djd3UhEqrMPdJ
o689j6enXs81kBPsZ36/Ydzu+IOAS+PfWsToHwGa7ReCrbKqJU3rTYacHCBKNBSIZW1tVBZomJV8
woSf/zVlrrZy2qLvLSh6u6EAyGENp0WXK5N862AOuiFu8BjZNefryuxI/gttty2QWlfcy9JPHlhX
uNmvmBj2D4ZpFkQZxOjladumjTJrVetKMg1mLmBNc6ZlBw6SoYSgNFY+fBBHUbo80lMtAQcl14k8
9eXrn8qctbktJERpRUrENalke+EmxB0fE8KWDjBsPE6vhmTVOFblM4wqTyXw5UGmwCZinpXzXmoQ
ylPATxdXbW/QIt7OHOZGGVCvUHRbBQBF7jMRVz1j71xiT5Y+iizdhMS4GLLEwG0In1mMIw0Mx1a6
8N6yzszNPoHQRIYhxa7UikCbYCcnXsfHZnQKSeeP+ECcjtxOEZIOsFVmUzSwWgYOjxo0KatSd6St
xCsPT4UJPC1U7yekX4xRdVuhGUdTZIU7/CL7y92bdZ4YiPBSrDLgjGuiimzA8L1hoDzAp8g65APd
ocvcN/zjph9CYoUY2eKVUbg75PQSNCSqELz7WZEeR4aDeTvzrJjTwnK/cIzeLRvf3fRsXcRW8kt+
SbrjJ8MDfhfciieu3/o2gqXXLC6eTzDDYMTUxGFItf07ENIeADHatGY4/4jNQT/gVHdCPAU+iZLe
UEjDpR4LiLPgl3uB9wNLLQYr5kDAMAc4u19eKG/2gLPTiSGV4ZxIZEjAUBfi0ZUONk3W6v3unGWm
olss8hBHPUFqTFt7PA1ASinjX0WxPvTnrqMorM1WBNkyIZBFCNzMkBUQQpTq2hbCSB3LNEvWHhh5
XjWcqmC5NzvwdSiNp2Zv/igyinA1Y4VDtx6v5nm14CkWFyLeTODxXvgaF20jrP7FMRR6EuHOlmJy
pqYnVJtfR3hpPn+dIeAMlOSRxLcAcDUixhjAqB2yMv+WhT70lUj8uDkauEOTitJiTt4zH8LLmHJu
frsUZy8B7Kc/xMw1ldHTKgCuXfKY0WEuLwMLtNiix/5Uju/rWa7p/0FaTNiNQ/qRh1baWVVVw9E+
qFUj7JSBfBXRq0/hwaSYQDcldgOTSZv/6E4Whs0/NoXubrYUdYlnFHOZQNiyxnvt5xLxLHZ6Lu4W
UZMayrYUdWQU9rnnZ1zVeVlkSWDX/v7J4Yd9Bw5UC5yb7eX4BRkdzFSPd9KpH5f4UXA3PJy0mXay
P9EhVgtJFfht41UVPUqKC9hdQmYLlvaPAJtUw2o2se3Q0ca9z+HbPMVTG+Tl8bN1RZPqL/JHNW1J
YMfvBDUJHp4xMeyh2PJni4jR8gW9PsdV7/+eCzYfI6EN4aPVPAA95LAYYvh54tW3wCshnjxMkFRE
S7zUbqUhPFFJXHlqp7vm+nsaaCO5TQ+M5uZPcAI7Zhvkzyg+liLxZvBrgLske54KmLq8df5OdPdD
T3oGcQQxCd8h0F80EOqkSgPRhFTsMHrRyJUfojp5f75vBeipLZk7k2y4V+qeh/iKjlE22YiAa1aA
kh4h4SRy6ld+goJefn2I2Qv0JEViasF2F+dRWY9qjutAR9u6ka5WTu4FfYY1KEszFjo3nvd5lNnA
RB9spSTaHnw9LDt1u4xjJL5dzw5bbhib3JRvdA46YRDhOjyDz3WdWwcpfJxrcdQPgT4JYAY8+1dy
HvaORoSSkUTuIaGcEXQeQuhzAIBufieSAqD/0FPDqlw+2uaeb/dE7SRAwmOGk6ZAot/9Q5kL3dIr
CNMJkxzXXnQ6+QVaYXw2WRq5igPRMsYTGND2+vEZe1iec1Ci4g8uLpedtokWsjgu5BY+GPao+XiI
a2Kalw+RH+uf6C9GMxEb2kI7kbvpJMMw6zTTPpiOrIrZ1xnukPefIAaNdH8BjPnj6kbgIPLycrdk
jnXi7bDxmelFWWnsj1XXdnnYIq8qeJPNMkX9Y4FTZUU2qx6JgXZGj9aDTEIeaG6kP9SxvfcvIBBS
9MsF31T3/VMDTF9VCGJZT3656OaafS0Uv0w4POddsDSp0OcK3pqoed+HkjqsJ0/L3yYnIk5qJITJ
QgTMJmVLpT8lq0C86imLHy8WqVes8KelITbDUrJEB/IZzclxPBpwUTQHb3IjxN2k4Kt0VPliDk5I
azUpIZVSbqiZpBvrmdVLBC6zQcE4nPNacCVrjb+Odq7PCmSQrKirH3U9Y8Wt9kUsdrdIQA8bnEO0
kvO31aJa7aeEsGwK7twyfr9e1Q1OnMgVch45nE/tQEpLMSUgzYd5qBlrfs/rOmhZ7JXIWz1UfB5n
haQnGop9xt5OlPfFUd+vLjZQ8QQjYSILnInuv0w/11UDqozB9LzyE+QEspYZOJHg1W625qU5A0ZM
j/qHq11OBtLaoWzNLFaEodRV84qWzyfNc2VHBnKuv0xo2D3SzjOhcHIyjgCTaBQwNbxJ1YC+e0Nm
3YKx3/dCZRoORlgzNNCm8CDJYO/qs2Hf2lZz2aZ8INxca6iR8jQ6+88dJ6dmwGJ660yxwPSb+DyW
k34Yl4WE52Kg1R/hHTRB1E2Inpu0CFv0BZAStX7WKiDwji5IuwSNMtI7qUAEL03MwQOLGz1sfg/V
IUTHud85cJaOe5wFBLTBeTXp5Po78c5DueqhRHHtpI9RRwF9nif2zwKJ4zhP69/30vex4zctIKiw
OpsKApdvoXlj5KkW8k0h62Bt/tpZ0pCHAUJIcSsrj1GtOJu4eHu0QzUO99I27vUyNLyQleAhw/e+
ALpokl7S/HwaivlHopmpNHvSehyzWN4WsTzAgu5uNUFkguduYX1BegpGtBbrlBSRCOcAU9rVTdNz
xqV0TztcGJU8frVHfUREAcK7TA2k6LDIFITMIqZvnPiBlGhKeG7tN5OpCFqyH4yK0V8sL3ubnvfV
RyMABEv3kl5cDTbc9CF2f9V4ZX5E5BAp7c/kbr2xbUuVvFahB6VXEDXCDvAZ0nS+LlNMMeoBWN6C
fg8h4dAWny+ZHNEAldDxHp7pmTIwf8seT7/bJ8orDlVwvDvnWlQ3s8q/s/KsFYFLRaud0H2c/B5c
cy/ip8sIPohHDxNtHV+quYw8e9eMnbnlMMuv2fE7+4CnPsfmm1GTea4SV5o9PNjlsaOHS9U3Zzlx
AE6PubqJan1Y/DDGd4l2U6efUQsBv4tnb5b1lfUTXuGLsaEZK0tUhu051RqTCU4hffNpaJlJa3KQ
XBJk9tn77zPdkImnZ4xYIiH5v/WtI1ns2NnZ8Z9hVbXXwW2bcyJ/tfE6SOR7+svH9lptQh5QbOrJ
TJYHsXDgyEzo2ieuyIL6EJjRMMiQZy74nWNdLS/AT8Bwgp5b8HDCin5Tu4eQHCD0pUtIxLOg2WMn
F3wSw/b/h7iDjBfFu9bQl1k1I75R4mID87AW8I+kAukHr93NU7M02kR2cIuJd6Rcp3C/BMcXw1Tl
ER++OFbC2g2YUr1GuRvhz0MWfLFmUmkWeIsGZxwk321YSGUqAGjN8NyozJyc2Yef4uFevnTZo1z2
fUDn520kH6/0Ecm7iz9qpBWMKuwcs5MOKbm4QoefkgeHKUF/FXuyKkevob5h1DQdBt9a3/xjHCo+
hOyteN1g6iT9JenGvd5TfF71wbOms3gL+c+uFS+roEjaXGQfX+TgCEG2H2XNE1xT3vq+HiBb0iS6
4MXv0u1AELsRtyBsvP+NiZ55+rT2b1IWFQQ0460hKvtbGFDxrwBSmthxl+U9m/+8usKT74EBeYvY
vQSZQD96xxPXj6encpDfqvrNXqMgXXVwAOIm8NJwPKZyJsI4gj6QgAWJnUeOROyGzejY4Gfb8gcD
g4EGsf6wEVgp8QcPdjX30a2AW4OjoexTJRIjw8mC5KHrF2si+W39B8p26ybI1gWW3n4cOdIko7v7
pdbwRi9rYlwgtONfn58PQaVJXs+a2n8AituUsfucXGjINbN8JLN6tu8oYwpGMbckeNxV3HsNZ2VY
Nv5gBikWazATPLGEJXJWIyJmOubMjugBXEHnvgkvmc91qi8igKVUrWSW2q9xyTqR4waDvt8qY8DA
iABu8RDS2YUVcuXPwlsq6OtghV59ZExcKihn/MqfmN8izeSyZnn+vE+R/vDsvbJcDF3Gpa2XzpD3
VDYaStJmUkLG4EQKWB7zdLfDloCK2MoHLsYKNLuoAnNuD807Gf1wCuq6UEqZbg+LxqIFW/KKSUFc
CFq9cZ915hXC3SozwrzP2rtOrKPxMPWUYN9VZj09CHz7ehjyD/XLDAbtr9xJT2mJT2dGUc1qgbX9
Zz0MYyCBtvIa02ac4+pr490NpHT4YNXZmIy2rDKs38Tyaj1CwjtZIr272imSNwm5v9UKQyxoz6te
geYkPnkSw3fwtDfCAf9q378pEUFQHZEPYVpRqo3q4rRsy5ioTSM7Dkq5sTvZSos7aV4GUtLY5CT5
NVApaZBAMeKzl/fepJA1SoqYc3DnBk7p6ZYXA7sKmJcqMxT2wy0NvXX2kXHIeZk4sMWU5QZ7fq4O
YqDBTz13nAzB3yO6ks3vm96kWn44AkPB4r7Op/zX3Lqjrl4Kq7QGbkfK/vK+EmnBkVR0/WrbCJXf
Jsh7tpqXi56Ue9HucMpSoqnFQpEK75KrSWBiZXUZRBbUZOXiSyUNG7MGxXKapBUkNtBFWhJ5yrFi
ZtQaWSAaBs3cX9xnuB0OzUtObTpbq0MkwTAoCVubsTA4+AT+ltu39cZLGSb2OJvRF3SYyCF4KwEZ
rEjeDsmsVY9KCFgshKluVN7lH9ZwfmDo9Ot5FGYOclOabnZIVxOIg1lwTO7lysgAl7PvlT4ZQGVA
b+ksc7oFx3Gt1SGgqR2wRmprLpVOXoEKb5F4A6/rIdRaoFegTj3xD9ctYAarsA0gZQ8eUtFx+oKv
pj/MiUzWJn2ebGIxyCZZ0ZpGe2e1IDfn04yvuMqVPWH26EMmynhv7jK8Q5tBvfXH27cCksXvIlEg
ZttrC/084VSNhKkP6U/RQiyjCrNpttbPkfTIOXkbVUESjY1GCgn11KXFD6vGQmZRcwjiGTp/i5tl
G4ggsjRIJdlweBTVMthFlf/wEKGynFhhq70brqxlsyRYbMeim2De2MIPvc9D4A77BTNBsl8Bg8zn
gJjaAyX8fMpIUVPeQ5fwM9CPHuvQzO3SBtBEG4xCvCAZValiGkG09G4wAz+hA9D2i6ARURQn0pF4
e8Hxn4XzSNLyjDQlp7fFVeDeOYDp4vgFL1dJTFGxAP03rt37Fw2U83JqCN4o+pUJD0Jtj2xoeRmg
hZEmzxEVLrS9nkkhByHDEfmVIWdwQltZY5USMTXsV5SkhGhWPDKsEvGKSEBLf7zyYQjyT6utHXIU
dHuiktzRY4w5ocBXgJrsApLxAXzDeakoze7O8CrfWOe46Qi0fIa29F+Yl2XPU1d0dfu9Cza6dOfy
HbtCGKdvWFBdRNianBn7VKEmdu3RbjReS19MqkCeyUXkes8UtfRyt//IVdvTd5Qefp9E7TkCK0cd
BmOuZ9Yn/tmliESK+Ec0RZP5SoNGKpTCuniWk3jJoeGE9yKb/dh/bi2p4unovsKiQCBlKtC01mlo
8NKzGEWOfjCKXK78iP4KwfVmqCl43JtNZkvqaNUwzQTGg27FZMdi3rzfClAFhPzgDITqJwSjLXsQ
VY8HlqNI8R22JUJiC0sDpRHpn0PETCOMCxM08ztQOMuxnW4U//NA/ptzNL1p87GDC+obMwU1pZx4
Fv3lm39fmnctFMvnUW/2AqFmNI71ubtfXUNuy+YJTLjYHoJvL8qqgzpHRukjcYPslZJ2nbdicIPY
uVx9gT+6e20FkIRk/tjS3YmdN9pec3fMMcIfI9KpKDP2EHJhx1w3K0l289eoLYYGQWE5nudLb8aq
1B0bQ45cLeGD+ZllTimWhQa0JBpde7uRh7Dl3tngF/i1HFWfSA1jHPskqw4Hra0GEgzMUEv3NK9V
9iwamzp1gYRsvbtERbOCOZzB/n4SJhixc77Gzoqvcoaqfzt2m22SC+GfQZta8yKPda1eJNZ7OYNU
MQf38ui/x+512KI8h2oD/OA8QWJp/vYf2TZhth55B/uzCFqXEdf27R7aXWAzYmfuxWCgiBtTRBKK
LP6xVvlrhArzcWDe/hvl285huopqIxnPfY9NOObRrlyRqIEomITT3gh6nBk457bG1AG5LUJFQ4Y7
tvvK5AteQxS+1ZcD062Qbb80aq8kOFvwfcx+s3IkuZPtKUbTrWiplT1fJkXiV6mtzEzHSbF1VWAt
L1cPbincgsKmp3s0CdhRu3+cQnQnwLaLkLEOeWthKEZKxZppsmWpNd1HNBXuDzB6QISDscgdE0N7
HMTCOFwZlP8A7nTNmNb0dQlwnFi4hbNl5jJz2UTNTH/TQ7JfNXMhJTlANFIjFa/TDE7s4YnHiRG5
09y6GvRluSuCFbJ/gozdU8wsrSa0R7ivclr+tCCsNxH+tx+4RKYc4anEax4mCd7TkqtNeDzA5tl6
JardgcT66AqfxgKgYU8Tea+YVwDGMiVO7DSu/87ycUHpd68jyETkZuajkjqTyB+eayno3oeriBek
LgNyQASQIp79k79rkp31m5iHJ7Oveylvx9FIMeXxuikH6j/y/wRiwRqK4BjqRoXXsgwJSLz5hkxM
RsIonoFpYX3zDeZmrVHU9Cw11uKWy+d5+/+ZFMguIdjrzJOtNc2myiJ5n58coe3w6oJdraVQbjfa
ps1TG0XUuxSMW6OTPDsD2vVToiJKKPNWfRDcwxkUlnZxiWS6nhaXwdYFOQ6G5Pnrv6S87VFZKwad
/F+wEiezU+aIMTkvyuYeHAB1dFGqFb21m97DtgKgd1xXFybOj+TluoMsxA7ezJVCbYIt/Y7qPbqN
gt/MDsbXjGD9h+O3XifwYPGrUjco9rrZwq1UnEmT1yvx/VzQapeldZ7juHWDRLKWYu3HEIg97gTr
ljSWtfNxOMJIbrRZKKjf/Z8r2fHatnn2h0UlUgx9Xy6BR1oodcUdKuhm6/BligCLDqhBW2eeeHGW
nNssoC/Ulk9Pv2Pwa8uf8zt7v31ciZvN8qVHbZ63/pyKGGjpWCw5vxgFfdg0/RcX35V/6i/uYUH0
MGpuRBcA9c6d3Q4FgrvagF15ha/3OE4IbbFkTinhhp/H4eRHoRUYDjGy0jz4MmtRjpg1MOtIgkV3
oKN2+cdZvhZq4j8eg5dIjYrH0BAKlSrdq4NFeph7I3bcASqR6u/v7tAP/RMUUV4B5CK/WU2FVCCV
qZpnlH3oppci2nldX69zc0Dhhd1V9JOBrl9SPV1S5S0Ys6yjcV4TgRsf+BojLA8ubVk+pK1rrZjn
1EITzZT7xBbdEyReDyMcJDUWzY6Y9+e8cD9cSpWsYh2hxTbXI33hX4EHiEn5HkRbiFlK2QaRCrxA
QxgJzeIIzR7JZpilUNRg+Ibg+ErT0xOXzjTn40BVghJe89pDbDGxekZqx48UqXJBnSysKuECkHiW
0xKyRpE+Quuf7SKHfhT2fUuXhzS5kQy5nN1XSgdAWYwMxl0/8KJ8jfI3s8PQr8Wy0kvGMfNKhqC4
aqEVJg4M3i3DbtUXrmS/jL0H6xz7Ai6S81iH1PBm3DYVMyyTBD7oyrSCs7bh64PWeY71W+rrNZ7i
CjnZaVu8c9FqOTgxrcuQtAOUZOUutqenw9SkXAbbOiQ7p/ZBh8awgU8ApTyH82a83nhHv6VYr3xA
ME7dHauG0wwlE9UkAn4yr23j+plb4XN3qdsKZTeKrjv+M5VzKQLke6zw7WwRzSH3TikP1gyVp5Bx
Oj+FM23+QfkKy34b6JdjGg3e4UNxSE6fB//uLxvxOxP2flx2S37Ramzoa/cmKdMnLqVITD0/PXs7
3ixNoDiSXmFQ23V9zufcFCy9red9nSETPmGPE5WbgfcoT+GbcIVg9CFADgFMk4Vt6GCK8QCdT/nj
l3tisdN5a5XCgR/07irMTP/+2RAj8kgkZ3QP4WM7OPnlyy/VKTH29L6SL/zW3VVzfnUTm41b1nmp
AnH76bTmn4/YfQ9rZq8ocXbwAD8BKS53cn6/t/e2NvsO/gyTKfPDJJ2v3YmNUUNS++oxHIm2IeFt
9R7WGbAcXlNxFNRfLyIBwB5O11e5VBd87P9uvCO/efDnYwlP9b8FIOMPtoBhIotPo5yzXsZrzBUa
6r/9dtECgGqQNq+goUgjmAATubiajjsr5gWIVuP8icKI4VDFcQ3Kj7X+lcHgF4+DOD4aPPhaZU+J
wu1MwzYQdhN9B58tTxwrUdUyvldN17gR/W8OAFvsKQ10JOO70/gb4qhAoqck89Ry17/gc7kAz7d2
w9WV8/9ahXapjYtIusx7EO24tOWFD+OdQtdHMgWl78K5N3jXAKRSjwiamoUs3CHhsE7BwhQmRE0A
C30CTLEYAUQ7zcZ8C7aJUXkYjB6M0z4BaJ4dVfi06Xv95HUfkOrlluWGtuqxoOAe9lRYHzoodu5D
O1D+4JLb8RAVhUYNGlZjYZO4mopR1WTsaVnfiJcgy5rp4kK73KRbnAW9hORGjy/9eQVwuYPcVNFw
EvUeN6uWwx2iry/hWmUrCrK+oTht6CXnSYE3/tiP5st+6Wmc0srJfE6j79oaFThjPzSakmOaQLvv
xY8WboIu/U3Iu8t/EUyfniLuQjykNmW4O96yE+UKfBYUyVsjxb1509txVfbKVeUhhwQLCwRXMeFM
uZlhus22yy9xHsmHCO9+tqFTPHlIEoK+eTg8icYsiP0nVyjd1qCdZPYPtYqFQBXZX/SsWkhfPJCu
FB29YmK0asTsvkVbOOAXHYzoB4r7x+hRMWfDGLusN/4PaHteJq2W1CKa6UDI2RiNbWorgGz3FftD
/xp6XOqvEIeQGKFr/JYs5uOxb1IDgY8NRDpvYm08yyMRAHgcOltWM2C5TBEt/ivYnPTpDtcHlqiQ
mP+Y/2Ouo2CYTptcB3TEIHJ4EUlGxEOsyS6rUmN8YCflo+l7T6CLROhZVQO5s23fYzCvMgyadFzQ
htTeuHjss3bXaZEjrxF9gdeJ8mUhmF/UqEhsjWImAHef5aeBalAusssC7lBbCjKsDwi1CNIlrggr
csM9/55dfqv8qjDtiNOhZK2VwLL60AJHE0LHAQC3JPYKUB9Ge2O86cIl1jcOGRgHT7dbABXQG/bO
s6nxJyBSCserSi5f9BDm/TAYhTgMlC8KNg+OUpn0mfzbk945qTndGPxWK6IyTrW7txc00pXlG1KN
exnt8M9JL30AWvDQe9q8kyRE0jMwxdYsB9K1fTIBLMBj/DUnew3BCsRLcpl3E2DgFUjkZbrFVZ8k
la+m3DmJb010fZjNKmCZlq+QABVch0E5ErOQ6ZwnZOzjnMJlbM+j8Y0mvSbaK7OQGUxPZXBXLtsq
0GCtPsyJIwFmScesMBr46vmifkI3g4CqxBkrnoaQtmTf3tRsSR8tDZj1w7j8Wm38X/xndOX2oNMP
gGqGVfiZ8cJonxiyeTbM/JOPXqean389D1bt/3RcmBJUB0YjFYNyfB4yestvD/89vdvrlfUJznxF
kJFNl4LkC4VYyYOQB0a4MG0uUNkpSAH5rJrMFwcmfGxnP9VnvLiwSmcHzsLss18ZDqQ/+xKGm9Oo
4wg3L1096KH5JHe35AFqpzma6hgnaS5GmtRK9qPfB14qpnDmD99y915Z1I+NfCQJnNL2QU9iofC+
gWcv8XuO+OUbsIaU/lRTGrWPTcnVNOXZNV46erWEQm6GYLVCw9M1nGGwNurfdxo4CBkGNUpQWM8c
crPeCQshvBkajxHH4zwV8B7+e9JstR2DVkhPhqY9oATVVulGTNNEkg6ZUUqBww64WgAQfctFeaAb
wza+xB1I1iB8iR9vSxcoFvqlXLS/Zp4EO2eRlEi4vs6G11b4C8OTem3j059Y3VrSEbwqQbWwKAAf
tlcJ429obiytXXeNFM+iQ6o7C3ImEW6KWwNF/MAe08wFtzMwRFuMD/fkQQ7qw+DmDVAKEFj/9LuW
u52qBR1NvodSGxRvle6X5annUat2dZH7+hZshEmh4b2nXE4V0ZKzC/QFgPiKTtgeC0n5YLgocXwd
ni0FJLVL7vW8QaL/7/oKtwY8Yl/I0GitEaW6umUkWuVunt0n0zpW3f2Rg5SaX6KCiIFCCZf6v9bF
SJxQevlnqNnvwuS7ERuH+SXQDed+3Gjg2No68SdSLSaDS+iuWMti4RAK86yVgiEvP1WeeHABAjUx
xqSLAizTwCcFRSuMMyCgdriNAWKVMgeDP4PQ/mrg7LIayhPCWJPSQ1VM0K3KSBzdwcJksDPI1HsS
1tJl2X4HpJwVzzDs8olPnZeCGvxUhHZzS3ULtbNYhamZGDDdcr0mw7Yvnc3cUvH1I+JC+cQiqKsg
xw82QZfxuOHcH7rQF3HVyLyONGKTffa48fqxEFyI8iZOQSnURK5OAaZ/usj2prrrJAsj6XpoTFmD
NJin5ibUzNwtmxfJTZ7HCVkJQcUHi5mjzQn9Cjd8nZ2tCAosOdh6ewJK9d9QbTN1R5cspeZnkImN
wH3h8VS9qMoiibQWfREvo1h1ASiCfzPj2TzuRo6ANEfMp8J97ZydcGXVviOITpjnuHQtFbl9TIdE
KduNyaW+EtBfA/8olUSYKUhRs+8ReSpAmS12V/6M38Ydeh4AexNgtxC5tR4uSwKnqB/cGyVMl0bS
TJFRQzwRs/C8ELYD1l2MR02UIw8BR54x+ww7q+0M5VitGWyHzoFUDIORVgfAo8CkVgLOMqGMpC3d
9LcaU9c8wzoOs1HKJnDOww1y9YdJXpmRvbpweRVt05d9zJHJ084LGZBoyYq5XqiWQjYVh1sbiAu1
Gem7REUmbEF9miqZ+qloDSz2OYVvrO9LhXc0bv2T8B8Ida44bFSFor7PGct4bnCeYIsGaJMutD1t
HshA/TFqFSI/DTFovTnCr2jQ9L9Vka4Im2fvsOdaJSFIh+28ri4ASYxbLkz0TnAQC5UhN2TOPkw7
lgrtyvw6z0nobwpjrkwUapAFqbOComAKtjlco959OMGhOphWjFP6npcGQ5tx448ZrgG5y8W2WKkJ
4W1StYLygvnTS2XTz/t0HYzZobW7/Fway6ku1iFcvqIW3VQNS4Zgmc3vi7xnJuhYsIbMpUCqcF8O
r2S8KvDKBNu4yDfzAsgB4/f9otWmZFsRRGnQKqq43E98wyHSROMMz49yhho2r/7niQknJDQROjtI
1qW75EUa1uENgQ/OQhVRsJ333SVOk3FrVo0E53K4v4tNazrDD7cKa9CsJNVtkMHMAvPe9PnK4SVM
SKCNrxeIl2AIchQNc07HDBs6CK4RDQ51YwT1qyVmQjCbJz1E3A170LFLWDzuv5IuYvJxFsqEZXrl
bH9HV5J/XzKtN+Fd6ISA2Q7lzp+GC4e7CRX2YxRTr4SgvaTv9ZgWWxbIhqB5Ax04u5O8a8RTsPax
LYKrBdYh3pJ5JQUn6PNaFs4ryc2lmtSb80reiM53uAhof0eOTkjWh3oSm9ACiPtHAWHhbovNqF79
auGIqo9SUueoE7X98l8CN6atAqTqyfBreN/Rqh4nZ2bAcez49VgYW81iFZw7A1I4NJGYxJMMZhBK
g+Bv2HPfL6+4Dtv+m1cmmULxVSLOzGgKHHLLCoE5qGFBz4H+adxQFdgmMpxIYaIVt4bFk0SioXXe
HR7nGmpUA65/wnvT9htLeIv3+hh18MnC1xO5F9hspN5bWKiUPIEjgv2DWXl/44dKMXXNVW0fFIyZ
+j+UXpHYzfrHAaW+IZXXLX9zryp3STPfib1rBH7uZbh6RNc7UfCgBIxJASbA/cmBQqf/znW46HBM
tVcZI6eYYVDJ8YSLZtgI450MmHlZL8RULkDWKinLeJE/RmNqzFhvITP0kmyXH7M4S1RzLLealPS8
QoMYkId+7qywYkUu93NoTk8VzwAaiqjSE0G+h43mrgP9wS0nxeDS2/BCMatj+62Kmv0aD+Ax2l0G
rRohnA4EXkmAcQBQSojQKxULL0uCgiLl8cTmn8B6argie9uAHimW9CzokiZbiwpm7JVrF2PCjCRr
At4JbA8f8sgPIigS7QL9PXsKaaTGxoUeggwlwkiSJ4L1IxYgzOTXktVLkL8lpFxgaJFSWR69xktR
DCbdnxkMiRpGuM/+amFpXPvNn2wKCDVsjn54wvvW10RDuBqgIJ6HBbA/qPv5UNqvLGGkJCTrixhO
5dBrAZxgVJvkkTniXUFT2GFnhzFI/MclNb6DCBwUnoAMrO+2E5+MyoatZLkD9UFd8Tja8Aie+lrX
e5qvHnO/bmBgkBBisx6GYR+vDuUZZ0HqG+aUk4IuQLObQcfnVlkd9bwDyGpbLCTqtNNDmgmp5OSO
3bCCL3jjVLJISU9dmLhCUEMF43xT1aeH1ejefyThkSDyT1TumWZ2WU/g9SlhJE60BnO2t5SAkCQB
/rguBVDdBgoeQBezOotDkIROl7zsu+GoiKVRZQ4GbXV4r/rU2yHWG4UaGcr/gaQ4Re2qf5kk+isq
62f3TaraZuORY/FniAG30nmDnzG3Uu4GQbXGtv8U9vq6CSwxZadtm5p286OKO54y890YoqOtrFKD
MUJOPNobBtIpr5qP7iMmlxeS1qt0Fy2HdjehYiVnhL1fhy7d9uZOyJTxtNIbZ/llQ/nbQ2cJOm6I
EBagYX3c9XqLPiBJd1Fn+iMhEk0CIlfMOTndtbAWdYBI/li3CZQK/+6Kb2pa9TcIxvoMwSnpwHn2
LlxswFVsaXudjc1e4VGhf5uHt5gIPm0hFPr/+EF4jiwd2hIJPcLfGivK0XCMNmqfDMur/TxSgLJf
q7atv8bHOGHFhBf1vmDTMJ/43yUDM0NDh5PZRVif0jj4Gztiwmif7MUCWBRZv2BYWc8i6ytUeTn/
RauJ6IpcWlWhE9sSKP7FkRrsoLbvV9X+yHiqjkidffF6M23fghXXHIDTEVoihLEIe58qr5iuHCZJ
NmdPY2vQ1EVyIII6p18Zi8PUzfxwOO1iXZOuMDDQDVaqGuUwiKGBjM0hsaip3uwQPdjACgDyUdMl
iobfaQqOJ3owLjnY90Av4dMZ+hst9Es+gPDrEx7j5QBYkSGncgl6l+7u//r4k1981jQUI2mqlL1S
SEdlUYr0quvedHODr8WgO0WWqVtS/q6REOizxIeqoNEftIlAwlTOBhwupUZ5BZnJK3U7WRXQ8K00
Aj5nEQb6SMHX4SyOHWZ7bBvNAvXvKh9E73cDNBCdzR8zZauIYuAJ09ldHg/80XWm/uL7Pv2m0i/Z
slcASMbO+QIswpYIXdiIEo1aeC+HbYvfluWGuw3rAz/2wa8DEX/gNULucKK3dL6+F6R89Z1p+1uH
coGktiWGDXQsJ5H3TDqsFimKKtcXEWQqQukSHEgjGFCGQyAfwrbCMq9Wvp5rMxd48yS8Cee1lwI3
Ahof6Zo+dTSzkpTW5IH2bjAx1oHqFBB2UWM01ErCSEaaf6/nfVv8pRbyLd+uz0ad4lPWwf90DPzT
i1CKi0mkEEJAhIvm0jFsX5hNQC1OjwJqZYq6thLiHdiTvaWJoXK3DJuz7yXjCTyfIh3/Kbrfv9ws
JhJBOqmge6bQrnbWqg79VGhRiD7WR28luy2p2ufNHl30yLLgJYCuNHiEU0tc4FIxiUmiKGHtZzIv
Jl0zxTDwW3lITS+JGCP/JRsCrAvnSgR3pmDYNdJGO4U8rXZbwoV20aEkR1aVWzelIoyb7Le84FR+
sE5b7dGx/oqfsJl9LbGwaYhErtXRrZp2fEJx4pi84MF2WqoI8yPgjWIzs0YaviEaCFzWxHW2RtdZ
/lh+ntzBjuJswOLjTY6xpDKhDThAKb363YWTSirf4Dz1p7Xoytx2gkVRM7qa/RCO2rsShPp7AFao
W5/TrzN3YYGHav/j9xZ2d4tV3noMDN2/RSrfYfQP+yeHn+gd2XdgIaB2IVVlTbpvpUuXTHfU7MWh
c2374CULVKR29EIgy2SIv/GZMcw0v/tvDxOfNtZ7pqe+UxYrKuWjvnUY2fMu5uRSvK8+hkEm4+Zg
N4No8nPvDt0Bd8kXZPAf00kITZT+UvcqJ9MThkadf2D9xIfQfTUiWlzeNS5Azy030je9Wx23PPwl
9gEKEvkw7fLacz/VZM0Sw3cxL1YbuyQbcv6JTwCWa/QC+/ETrv0uCETEpinsVt2CsDD3wvR7qAOq
SGeECWNdbRaZrJyWFx8oTD+BJFfo/y8wQ0mdv8BPlolnlM8KPziuLLJ+RgxYOIZZFQIpieWeovMR
EAGXSYmQaXBAQIikXHZ8NkuHRdNrIVJxi1CcvH71LZ5DfXX0sySIhEpfGW3pk2QIeF3s4MZ18VfG
TaX3xl9ndjTqOqtWdhOxh7Evdb90vdWLuFwzB6qrGyeJ4CqfMAWBFaF136eX6IfK1gD7ZgrwygE7
hr+Tos9WEt3Q5evnX/B4WaeD3no3jz91mXhR3LTOCyrt4qjC4IN4x7Ffgxb54HFWOS0rvTdLG+LP
p9cNsKb8/nYbyiRqyXBmdSZOCQVKEfVRVV4xfXq1564MGdZQxPLEZ9mOXWLXZKhGQzicsPAxglQx
sJhhyLIduKaOa8p95dSVSNuN35QjdxDqbYOvb/qF3/6g3bdbVoraedvMHyG/v4pMXiA/DkK5NZHF
/bhITX/rZtFZ5kda1g9UC85k49gihjYY74afnwMY7AzkF+07f5cENa0JgCYFq8c3WCqJGWsWWhi0
F88FfzShjMjWLA7d7KK3u7hwHw93Yfn9COR7Zs26hC37tTE5b903HoUAQKHFYA7X8OnE3FXnZGFm
BCrNvQzkM49Nx7r+Lvs4+NQNLaUi43vnloj8A6xngMQFodpAWo2QR9vN/dExVf/K1YRNamUOqveI
kZZ+UatSPWO05ucK9bT9U2SN5oEmqex/Ru1cVXV0vGVKRQ57yBKD6x8kqRgnCT1whsVz7lsuhZRp
mhYvihe9cs5+bcxVrmQCHTxsEjNxkxldcbR8ENnZvW1GIdsSGnMCQpEo1VxYd+J1fcDfMpvGn9UP
rZxMM1c/S0wHoyerwWygmgirglDHRJRf57ldtb+SQhzgKnrXum0uP5Nya/wos6YJhlrbndJsz3Is
Cdg0NqNwXL49BJaBa25TQLnXHbOOxAlGjyI/ivSrnkzBVMC3b7ynVk/PjTWYR7j4qbXzAM2EfuV2
VySSXGMRm1g1gDxhGo9LFzARqxiumgu8BdaOJP9NFhtlfqVV2Z81s1I14lgAb5plSmlzeZBeC71/
ATwb5+uiHYhB93PKaBuRIDaLicpavHBn+AuKA3J1wHOA9i577rv4S2TXScSAq3jqg+Z+b3F+i7Jm
Z5tmDh4r7xIeNQxyKVGLxLekaXv4kZ0uly7jK0aIb8kMEd8J4IEudz6yNFCpFfpABsVwsswJaoeC
8Sd20ho0yBZQLvZjwzIbIJE9Fqvh8SuSAGMOyZLII6CEoVFR31rNO/MygFnlexpo9QRWtTN5QQyS
BXMKhEAFUTLxT3rSpCTZweaek2o3GUATdP6VH9ed2jOousW1DAew4VhRZzgIvKe7dOoXWXL0jSAN
hS6bZBAnpLBDbURMvlYOQzcdJaR3NKNIMIoSyn/8o36WY7ykAHWdCAmmbPTd001zAZHOpBYNs48A
CFATjAxF79MnYUSCSxw/NenfPvNyzhxC+6rs2v4w3GthkjbagAWbsbVFF41YNc+P+EMwHYUDrwBn
wmUfWWsygoEe8rXr7mKu7Xk0+VNXc2RZz1r72MKqsCXz3mixxmgBQxHcPRliAr0+bnqvrrFvk7Rt
U0umRDSd4aF+ZCREiM2UWF9swU/ch8x5MQcIHBpQK5kns9SNRtMiwzc9jKcjSMxOwBZV286qDUFh
XmvcgIYdAQHYFuaTggX6Mj0CtNDQ1/00k+gyiWOAvr1l7Y11iMWvLavUJPlOlZNFsDr+al7zbREA
lT5+b5dq6QYtIS6aMx5Nj4uNIzn5hm5JX2L8xh4ICNrOdg1UPymdkgzoejOm2nEO5E/WclU1sVLl
APp3k8ypWoZ3F2vok4nv5f0Zi64ICrDf51dkuQCB/G7ecIABXhwhEVl29VidyBFukBaboJAT0nvO
jd6frJKMt0V/GqF1N0i5WIqLR8dqQdE6W5Yn0p7DNmNlT0KMybisrSa5ljiSNCBKyAsVZmiOPBYk
uvDkPInR9Yiy5HYn7Ytd9be7uc22FPAGOf38SIhF4Uisirc1oZiXil0gw18gydP+RYZfKujJM7ft
xRB24LK1mf8H3jnkeWCkKm2XX+kYp5QAk5uhN0rb46YGUjg56iNcFDCbOd2yoynlTkZi6KM/3Zzm
W9ddK3bLpEKng0tTTA0L69qOFAXgpZALg/0NmwrjLY5EF9EyuLVHqmcspedxu4wQ/LL3CHz0PfOq
dU++aoT+R/BwsJR+n4vGOQRoI8n4buUAO1xn0GqU1u2VRAAeSFRfDzpViY1nf63H34F74fdSZ8cT
UJ+aF6xavB44WeLJ32IxttArth2Sh/PrRkT1fkyrDiQwCVqRiFdUSX8xYkPSsJe6pNQ+oUCwtIHV
7WRIIvxRkWLe5FzG5bWoyyU3uIUdjhu5AEQQEkzYHWPIm5yQTt85tq0XUJFxazcK7+a2LUkkHcFq
VJKkgcl9M6F7m2v3boSsHeTQ8fGfepLsbpRxdKiLAzAv5rxAaKXVJxlcdXAkwVbF9vUZgi1N45i3
DKRN+Nw/zhOphr6LEqr9twmX2H7j4CHswTApcNqfnezW/BkXyF/QlXfSQoX6GqUtviH5KHyOFzjS
QI6wpKbrC9ldEIc6mFEzqiJw961CMYyQLc0i3QwOt0SQnAjjBOnknE7JiCE1yCsZRGa9vNKnbs6T
mngDMfljw1XpvHMIGvZ7giCDQgDFTtZPpk6O9U5JYHt5q1bBR1lYZSzFGv4RawbWgGnGFgPmx4td
UgcgIz7kARDfyvcr5ZiYFmgQ6/9Lld5RXkYK6Lf09PoUu/bM8282rgTmGMMT45h7e7PscbSkBana
ZQPkpJ94rgSMP2kn9xjttIfnZK2B3NygKzWPJKg4kOpPZX7ZIJus7u7yLFn4KSy8U1+or6xn7bIB
9xwyoXXbcc89nmWRANYjhJKXHoHaSsoF2XYUtlDauxdwyIUN/YMeODVG32YdHlvOxa5EOdoiObXo
OSKKLCx7eiBn6kKZTMfjdSTdgScvd920UX0yYpHBpTLOB+lTmjl3BhCQP6kXpvoq9G+cAzTg4NMK
ATq8WwM1S1Hk6oQ8GHyTu7pE0gfMkEeLIIkY5EsjDkMLmmn5upKtciBYUqzosKrnINPb7CxysVlA
9Yzg3rTW8TypUaffy6+ET/9v9ekUhBpbfTWBPHR1AyTWlJQxNfftSXalyhyudPn8e+6XBUweRnbx
DAjBQRalW6qK0B7rXxyA63w2qV6mS9/X9w7PlLi4FHmcISS3vl41RMWLh55PwVvoeq+rTIxzwvlJ
SN0g0dsKVD25v2vTfLG1TWZrOjN9/5LeqCoszYYU2JYcDDU1wUij8fkLkLafCNiluMVloRrlMclw
zUiiHX7dyYy7s87dQS3EeRfV3K6DtfAvyGqOpQENbBFx4vReKDXyVQsN3EBo0o0zFccuit9PMqlr
zqsEDzdI4k0T1Ic1WFvXuQZ/JOczmopzj1yQz4HX4Sdp6dIfsw8fdQ40yRaFfmiUYSWXa1b6+oj0
E15kdIMfZ0AYIP6UfEfyzs0hawn5NQOj0ATQaA5mUBUgQtRU8G9V/XJ/Y9UU/pkwgDLBr32ok+L1
1WDDy9GsbMFi+tm2lqx8yg1jw+e7FocKi28XH6aO1AKL43omaRTdrdyt4HRdznypbwToDyj6tCMI
6na++U2NQG2Af616DrDcvzkd5RVPfS4GlFTReYL2Da5s6N5aBqAC6asMb+w8mQ6bE882uUaGoqlu
9jIrlj+aHcO0s3Rj+71MRD3GYQUU1jXswm3oA8qCsDPYPO00ESos30bDm5JxK7BAKG2ypXKirDjW
q5aKm2iVfih40D2xRlfMIfnPDcu+tuJfux6kHTyiFe8rT3HgDxwm/9HczSHcFYymCzghrS4xi4w2
UkvG5fC7zvDoTOnJRu8s6Ves07wL08qJWjUoYL1LNmOjX8EDSjlkTL7oFw28P0o4j95Ho69FN4+W
RKL8i1iEBRD8+K1niXXA1Shu6FAKOyUYVchSDX7zEXuHvliq80OwgK9GCAWGSlxZQTZqwphq0l8M
MDKDTzPYycDnbs7O8NqxiXuS/+McV7mnvnVqZqqPFCkwGcRU0kQhxHJvojREGPslQWh9XJ4zLuhP
ub5gyGvyO6x5J8ynQ71rQ77P5ZytX5xqpMutE1yW1geDqkE63CZWKhs370jTsvChEcubW8wc3A86
ydSJu/MwaCqMHtBbT5cEq54ttwpyfe3oA6bS4Zy8S+Wl3LVk0p98dkRf6dOfiPYOoxfbPAUSHlwg
SGmcBRiOB19ZowEKM35fWpgRx7gw6wRWwUjjGEZszLDpPKL3QvTVhouGG8XtEUR3cW+2u3kzr1+R
04aZKp+xFrSFB0S1U7LxKplT+vkUQorrX3vdbMZ1cmdInW+iajUuUgChQUcrkqnMQHlNcvdtcqst
RgmXIqXcoy4HM1Q9Nksisc6fhOWlvNelN1w3xNUQkzCdntnRhUcs8w4sjT2isMmEKxCPdzrFpGuv
LtkiYj9/EB/17t20Rg3W4KNUsf+Jz6fF1gFcoFqP6K//UabHSPx3Uq0st1q7uFniGQr64HpOoRaW
PvfliStDietLpBoNGuIXOhLIJ4yHLbTBeCH9KDsnQ4hiWlnHFxQzQYwCmW7fjDVHkqHCFShG2qXn
/Mf37/+BToFkDwf9yF2peJExhGGdM0S8g24lIUA2I7qwrMuKdgPzMF/hMvKy0498VQmkVaC5XzVK
zxFe1HfBmvCasEmQbp8cy8W13RojfdFGOBE+qO4OXLkAJprQkLi5RmgxzbaIptlTk3DuFuYHrG/x
J0cg7u2+m8vX95y5fwkhsEN/N+7tG0RgdqmGcZskxiWpXv4dnXteg/fHrbINo7hAtKWIdQI2/e8Q
sbYcFk9jGka1LJ1b5bJmx5mzH6DdEysMpf5XkppqIqi7Az5TquMnxpmflWzSxwO0PXYiKR0CPGRB
XW5xb4shlfD9h3a6oKX5XN+q7wt1aZJ+5sFbvZSaPiXzKVp8KFSuk2Kd8pqZO2RpnN3PaY6pHRTr
1VjjaYlhrfiGmmHVS3dfg2ck4jpWe6pBF8QM5mxzBR8gSeAuhS5YvsZf037gOYkGI6MNQ7Zlye5E
y4NSyX5dEPl9QclQjAkrYztBkGHCTtLjQzfRmHm5IezhzD7a7CgWcHB5WIZpV7+XJjD7PlHkmiNj
MRBpXQW+9JJyuJcNRNrHI6k8bcjus43Fyiyn51Y1n5l215c4ozZrxzJx4UpJFhdOsN85QgEBoTuF
dCyCgS3urmtElKCnJfx5isrXBNO9Fsrigm/zO9RAROdv+f9EmrNcEF+XkfUjYbOMfdbf/aZdOLKB
Yr/kHp2NRvlAwdgQ6QDlI2grNBpo5SOZVqHCCHaKu3kdS/KBJcA0NPmv2gtc3aAwQgqunQw5n9Ic
jeMj8G7beZVP2yd2ZplLDTIPsU9WCBgwNs8O/d8JHO82+wMzj4KaYzYS3DsCLF/mcbgh5z3irnir
QdtA+FrLA3hki8fwrkwCU8la8Ikr0biRUNBQZonb4mVOBWPRzL6xRGVkLrlHT68Ipos/d+CgLHVV
IK+z4eovfL0rRYDEi2mUSmEwyKMPIDbpX8qdAWSc3kvNBjLSaJk95tOXGf3/9zSv3+Xwm1eB6wKt
aC1pF5DC7Uco7PL39fjxZ7OnDMhqzVLP1ub+VUMdLsziq0V1P/XVSPVyY4xMcfslj/QNt+rNiQfs
3o1oCgSfwLJtccjAPFquUvibv2mTjdcs+jElp3FoIZnTwtDjNm1PQcawipQMwOz3kXgamv0jqN1e
5oUo+Wt47HEodi9gXsoiZFWSWU33yYqHj7FNwYUKci5BoCCXjLBJLt3HOi0ZuT5KPvuD0K+VFwA0
ox18tcv4RKpNfEwTR8DBdq3qUSozOzPbtr48UA8jO3/58hAL2+2FwRw8V5yp+ZsF9ZS01EVmnN9I
J7ukaZBpzE04b/6YPzI7+sn7dhXjKfSIX5pAHo+mzPLdaQflUACKBeBq9K/EG/JvTBCRhErTBlm2
k4erIqwRBU4rNkKXb7IUtkPRKOjzgYlt5/EJmU9SO6FVVvgY7taPImdKCt6jbghvsrYlaTBUgXLa
kub8W+CGRaW9GOoZ1kBwZ0qPxWY/fiQ5pPlZvENTIp17m8Fckl9D2Zqx/RgW6SB+w1rHkzy9jEmD
BqoCzsjx5ANWMFla8zZOcqS6+0bK+oSjo9xsfvoOXtOvL406OHw5mz7SEcavMJfHEF6uurgEsnxS
ARt/tcXqvFuxDsisyEl71mz1bIaftrWWkJruS333xA4hEB0qa6hVzSsxnG0Bgy0DjTWqIaT6/UA8
0OgFQvaszs9wXGCmqraNbiueLR0UDN1ljnKuZLHKrF16ZQs2+4iIYIBrxgvuG6qpm9pVZrhca7pn
DtzBYQn7MrN0FM9RsekGMGI7sPkyIA7w+1uHDCYW8nvF5E3VbNkDL0NTQi68DZPNrGB/ioBaBwsI
sF0jUjconn7zdMC1CIKwPZI7vFGpIxLqenM5rdTE8vDMrhp+Adxyjfx5mdR4VlgBUCW9DapAqvNs
kjpSDGdh9YlnB0XnitmUxn1/L5S1TxFlgI2zuzWTdAv9RxtN57zZC/0BTbxrXTC0bzkik/Y/7t6F
/rpISGlht5IwbkQYjkvIW8ufRA7vcFNn877RPLTa9L8717t60J3czgJy1VUxbtimA4sr+hyX3fRp
WoZ4i3WL6hIDYK4gQ/R1LZ0AtDtApST3loMou5Jvw6QAIMtUAYf15qRt/Ql+ws/WbDu9jMConSUN
yTvCBaj8kSVOV9uLkRSw7WUBsAXzrXVOgBfT2XqFQCIHu7YnyAi8Le4RakAoLLaieG9LhR+SeaYQ
ZAgfxwiCVCcmQbqdPDpU63kuAhD/tKGeaQnu9i6Q5BOSYx0/cN1ciUVDBkExXg0v4vLyFtAkC3GE
Eka619mYqIghaY+ALtXavCZMzz58BGXQ1mmbSO9s5V9odeOn7kJZ6en6gjfu9hlWUmgTAlLq4v4S
sFlaBmAv0Fh0vG7KZWWdnHHKGpzIguoEGzh9/kKt5XCVsHGgvNrt1M2HybsiZ8LTIAmvdImSrYEu
W5kh7vPR7NEZBosk3VkIwQoOT76RSNEE55pbFhzIGHOl98xIowpLbqN8SqQq4CASPDjJBBXH+9zr
KTXvJIa83hnxPEJlPiQ+lv3jbwRBE7fjsA3iN0TyQ+30FzwARNz4dQeGqxcLqzOv/ItvjqVk6iw7
IDZr+WuJK078hJB8s6xx4a18gDvFxTJUsWUmiOcf5E+futJDGSHSdHq7DgC99+QqN/uJJBFBRXnF
Hz9r1sDT1rZIaJ80XRMFWgVCQJLbjwHj4xgEQJmsZ/5TQoqGl2Jq6F7sI2AwxN6XtceaGP374YjU
HQJCuAEEWAfU8xVkLnqfiutxkZJXGwaCF9YvUdRX2Vo+lhUxwF+7oUdMBx1wWkNS1OeRc6LRrN2r
Std+X7aHmYP12Te/FBzv8URc782IUDXlV1W2bgoIBIazpwNS9FTNBkp09BTQ/M1u4015Q/0wNWN0
aL3jGdV3FKqfDNjVPgKNzqYkcBH3/1kdtc/45JhuWGPtK3FqN8txjZ98lIIpSTBc5WvQ/4Dp1Iti
J1SGQtVZNL8X8Ny0vEF3jqrFr8VzH98zZLtou5m/Xzv02/24ra6uRMpE340zeSuitv8furmW1jOS
XlloKCZAJyyqYrvYtsO0nmfxfU9bhmDLSW0UW+tciDB4EgBSLnUPn8IpJV37hoiDRCTlZFfeWyj0
qTANneivgH3sy4N/+9IlfeIvJl8oQENdkB3NUBzblXRxxqekehcX+qVOAkHSNIwBYJ3KvCfke6Pn
k6tnszuZ+WSA7+U6wZ2ngW8kWbyMXA13QC/yM0eeQjT5OMYrZ2G8WWtHhotFhAaAYoV0Bz3HaL32
U0sptf61Cm9d6r07tor/p3STQ7gscIHAxf1I0wdU3F+d9+Q/X/QmL5oFMojfrVKnjG0KbuQscJV9
rL6AMYMSQWAyDNX5IQ2/MgQGsJ+W0U9WOj3XjIRL7U3K5Hx5qchPXqUNQZhGGgph/Fnm0V8J19Tj
Il8RmVDXGbvfFQfa3+eGCCo1+R7obXSJ7TwLCsTq9C2TUJOfJy01zaXywUrZG4hnFi3o9wJQ7M8d
Svzf3CoRxIj6EbNX+hLqRmF8emSVduYcJA8Q6QVYw7KSSu0iMgUtd/bKFBYMUR6glaMileYXVdDT
OT15Aey5KiLD75W+rgzjfZI2WtD3SttjuLj7F2Ut2KF48VQieLO12RNpNzo9qN2KOfpTeQWlpKbV
Zeei/lzlgRBrU32CJaTofazb2xkSNbde7cMCErQYpOd1H9nvRz7l1bBPOXXinc9CW+ub6Z13Tk9s
IM3Ev2tfhIuEEgLNzPy7gnzp/ZN70Tnw8wgRJNGE3riHDAEuZ41ZkY3OPjw+TisFS07NEW2AxlHi
wYR3sJ0e0XyXdxMdcT+2Td5LvYwCqNBqjOYYk5DocnsVeLksTBAV1HPxsXk5OgMRpilRl6UNXE9R
lLO4QP36d1IIPlhq4E27iKb3xGFe6zpox+rSZezJoJMN543yfhK474N+dyev/Js1x7gOHPOA1BOn
MwfZMwQYpRcYQrz6YfIYJ7RssHELgU6/VYmnfNWwz1NCrr1bMmhbNqf8IziShMeUysuGThtsQW4W
QiK3U4k9nWVQi+vtva+znZx2Hjl4FF9UIEkRBBoBr6eK51XjQbUf9mCzc2oCu0mV6UAOoaCDvFv1
uewdFJGKJVPtlb3tj7ln+mxwEwqB0MnfXLjpNA5mdndGdmbRAJWN7Ac3vIGEaKYSvnpZxkQ0mKOW
l72xuzFt11pSRH72wyxstW73fXBc//51yLCfi4K4oxdSqhnB6STxX2hHrvo6ePt39thDFjr25JIl
4BuIja94quQyxNcMhep+bRi/O/vNNEj68ms1WERyXXDkM4AgTnuOz26tftC7PZlD62rCxKoQvKJg
x7ORTYk/hPIif/wqLqfcMoYbdffFRZenQDa9eKXkorJ+7eiAgRaB2oC0jpvr2yvshpyu5Zlzuv7m
9IQHZhBhayXoULgVtobgFT6RTkaHDfsVAO+M4ABpbS8Xdl8wvtHSsThZTXENKE216XGn1J3ZKiKI
ENkeIznn0NAcpcbJH9UQZRg+QMg08VTDddE3UhpVkXuVRqEAMsosaoBNonwZPlhS90CiU5FdS5GK
yU+77ER6R8vmvvVY34mwDub8M38/90z35xs8kVUqBdftMhvn4uRPeuJNw0/VqQE37Ysls4c3jxg2
eKVNXoGI4EOQPkXV+j68tS14lNQtQ3cCdjl68XRiQtAW7MHuQ4MXiHr+Ah7wJhjxwvsLke8ZAj00
eIoal3uAPUXhczc4Fyl4GhZBZgTXxobQ4/+AoDYCay+2e8o24nnZnobeTuaDprnck+nD0LIYEAOE
PJNJ7UKybDgfckALaQXHLNkmhakM8B0EUATMVYaGNYibCtoq+hPUH5DWx+/+StjIlLUao1dgjWII
/kcsCv9VfgDWVahv+R1g+2NZ6Y+IYn/MMFO9uN8YCS0p/pf9yF2sJ967VDkUclZY52IBuNBSs4qy
wq33V4YjlrFwSivjHg7rvnnBX+1b9ZKg5UhQFub3TYcK7Ca7pt4nEvjLBtf+au9cvcXt8WgKUxWD
jqLHxZOXYVEGFD/wzW/mfrNtBpYWK5fa7OM9azqZKVUJ4ddLR8vOzuucNcoWD4FzS4ApexloKbCJ
NrpQFzeFlDeBJHmttpq27CScj8eWdSP/cq7UDjwZz/vvL603a8jgHuAEe7RA63+Dh4YA6NzMDWUL
08quor1lpAX1V8F0jPNEMrbxvXdcnq+ZJPRuaUVI4Rv+0Zw/xUk1qDNqa5s55orZ0O2KHUobpnyZ
4PPwYwbNe0uCEWc7WmVE+euKyR+3RYPd6vZMJjYZQ69MJyFlBEerT575fOhSTLkUIvU2UmHDro/F
ebNdTK9Jf0EwsQZZgwaIG53GqhP1wrVaeTC5wIBxWjNO0y3XKvoX2vsRJGmTvytGmMf2fFRtiXCo
tsnSXeKJY5MqU0Z9xAEc+akQHNSFmukvMJRL446t/HWaWUDGP92Wk8+JB7BTVWUzyxbao+fs0SXs
jpmOLHV0ZeurmK9yGVHOtYu7CUoqGNtsK/cTHV3KqjqXCgyu2K4UUcmQM8rnFAkaM7KynharOihm
Rw+gxbLDhQ8LppkOMX55O3+NcX9JJQn9CTpdHf+gAfA3W0XGxDkhf9W1L+EDhiWLuWqZV8N8suVo
98GgzzGA/YTgsSGaCRAywDEyy9xUMnQYvh/rOI8MKh5eJ2TNH5c0Ty+DN5PVZ9ul70CHveOYXip/
VrZ9ll0/3ZU7YLlVEmsnFrkiOAYx0h0S7sMm1cF4nfZtpNJTswIKw0WAuYYh5XFiN2EySVHNU+dR
AgM0ve0PC1n+W0MIED3alW2DlZZQZU58i9+QWBTIdYS6iVgzVy0iEwvk9+9wp7JvtiW+uNP+OEZY
Rue5+6Z6iZjrJf9CZut96R8FRjXH4cIltGXU4N9b7Lp/7Orrh74GozHnIsvkckbjV07Bii+jg24+
53E/ePgD9+Kkad1H2mXuyIYsjJd0Hnvr4t1HIlMfq4qpmxUbnazsHC2S0giwTBRGxzaHZkUKU1Yg
DssEegjTGyv3sTCG2x03D77OEUKFb9fHU6KSGHHhs5icJd1DAY+vH8w3omOm/2UTRh3LmsEqjHHS
mT/nqrONwHsijR2dqf/fvsuWvI9kga6u0gRV3MR9bk9ZAwgCiJRqKF7w2ellEkRJHPS3VUAJ0M+T
yC2MwNKxtNUNXWujvRLkybrl2sNdw4yyWummeBxdk2fyBIf9Bxv/lvtWfkinOA81ff/GElsAEzuR
G7NX8iu7t5M3dDkCYbXa+0TDUbLP9X0vVmmRaXY/epbd2BmKyB16uYNsjGpxUHXCMzaxrNoN+8dU
fKdQcw49+SIKkbZnu5Vc5nRI1NAT/sUihf9QZMsKq6yitWX38DWeZZyinMQa4RFQM6o4C863YK92
tA8c2mgfdKK6tRYTLnaRw67Mpom43MtKqTlxESZFWQrCCpzq1XAyu2D7OUU2MxxxImz49cAMaM24
gcGoIP64xKkxfl/EcutQ3yWkPdJea+t0jFacNUGHbARxWgEYmBt1m/Jl3loY21aronr/6QtfIfmR
XWTGUV4bIwr9M1Qeg0wRIGtRdMnJIPbQP71TqHDHg0TX3PKrgFk/yV5D/JfPWnpwEqjueX1IGsDX
fqAR43tiJoM/v1JQNE2KTKosyMJOZ6j2nu24LJokY0Cif9SRCyKhsDZ1NEWfAMFl4o1z6N6M5B9o
sNg4WBQE+ViMaTxDNsNzT8vFYCCezhNdhwhL5dgLwoBHY6tcZDt7QjnFnIAA51TROw2klQocR6yN
4cqbz98lVZ68hBvQz36tUnD/j6okDchxPlygqDySf7OAYoXcBZsO5fqb1i86nDRXH2ka0KIXV5Nv
ZnKf5aO4YjTkR2bNbWEH+r3KP95ShRIDi3t3sNNqzSSpNI5xotlIv1LerHFIruANdlFXbKHO/Kn9
4d1+LKErL/zsy9AGycH/qF6TFFrUkpDA5Iob/1nVb+oEI1WjLkdS2P2HbF2rfqz47xm/nkzzYTHb
cchVryHJ482+qmRZkhCkW9zDVeK0YXh/BQ8pHFB05nPJbiGRmtn7Y6el1z36Rh+XiniAQymh8JpX
FYK7YH+eJLZhR5E8AIr0XomoEoy/g7aPNYW9kDIrYiMI8/pqfo1FaMyDkpD6HJ1G2YTQdWdP47rM
K2etyPO8L8mjMwcIhGofFqHA9eVxCafSS77aROM0QFXHNvZ2xS5fx9z44fkMeJ12Jld0KMLIWg0s
tuvsN7VvZtcr6jiilK9k2gTzZlAzfYb8KNZJP0NTGj52k33zA+XTxr9z5Ch0TldD19WNrCHzLaCs
+QbqH3uSrb4i4Z13pUcmjY4mXHAXKGbH0+LCVOR38O3+1RjU4kcyZnsUlDPR0xKS+46cDkmQmji0
Byz9vDWDehkkeVJOwoHOUYptoV+03LefsMMoWlnZ6JasVlIhsdM20JzuoyIbt9Ijv69lMbHPCgpK
HjDZsQDUZ2UQTISkQK0fXyNZPxk5zUO7kUoPeaFYRZBTtj7yYIJT5yAR1YBAX0kGNw4ifzR0gv/J
Ok0z6LMgr5t2o3kuJ2De4z+aR0RNNnyqqQnrP+YlQiB/UUZZah4vgy9/SDqplpB8XKV3ZMYxZc8Z
5sjKAePOHYeJtz8giNTLKKjgWK2DuxStl1u0t+M2gFycm16OTn4YtI+O9W7L2STsqHoZpBfBYC3I
MicZhFWh4QewEkxrw4Spa/1Qfy6GxZYy8DGghvcNwCVg/YDg/5HfbOEXLYcDJrKyjcdvcrmBGqH3
AEV9/knH3iFQYRkdC377diCcuwTsNmuzUPki5Vl3odYrnESZomz6EFuoksu1okCwi6Q1O3lsnomj
6FIabPF4x4HvcCBatr6uBprrDDZpK6b3SKWa2e1bztvap8OiS2Ekf/G3nHJkg261w0dBkU0SPHvl
+XIhDEbGc37MG5v8gQyyOIlhgz+OlNgMcGtUuWPoKO7Pvn+iow2GIcPGcFPBpoPeNtkMQ6ZNuDnQ
g+dlMQAES4Gww7R6mjSiGmIKZyTKwuUv6TEQeVD+huV1ue9L/pGycflyj+xAdlmJSG6hRXwzjRht
SncKLLWOYDRU/JAbXcLmg1hK5p4521XDj83/jfi9uFX6Bvhs+7/WTC4OLbBiFzp6fN96qwIBFlnV
IrkBQhrIDhQe7Rulo/qUbrJQ0v4hAzUkWoSzUXrLhtOacR0HzpHD9jm6vi+0YfMPoi92H84ablFQ
CMr/b9TLe++fWq+j7HFOqKt4o/WRckI4YvVcGrKof4o9XnZXygRrhsDEfeo0jQfUi/xXzXWm5vKU
yawJCqQ+niKxusbI9khDLpNQm+0UsolNKzVEFYqbWQW7jnsGDnT196C7IftxU0n51OpxxI3bbH5T
l/YxGR85yHgJPhzFrCcpDKJJVYCNzuMgVTK9DcQNCmSp+3DSIyZUvTDBcFXKyAR/ZWC0s0CVGw4v
+S5UiVO46t63rAduk/Vnh/s/q9DZ87U3xjMvqUTWk7o4qqXh8fpZ1S0r7CTe38bT8KepFdfrp5+E
mUzwMQTU6D0F/1CpYBBJR9/bMFWSoQb3xACb9R5QZbMpIx1vFoJo9Way/f0cOnxaMHbCJMzFskG1
bdP274/1uKYzxzFg1aVSfnxOGIVsIleYy3sDInHoPLKDEo0TIgSH7O3TY33qYuvD3EI+ZE76GajG
I5BY421luetcywJYBzB0v/3cohofpHO6P2whbs9IL2AfwCuutrxD1yDATa7RHziTXlJq0vjo3bKL
Xpka1eItYFvHyXzakxFNGEFSqU47uOP8eEuKD42QyG7/PhzTRcZZPYu002PANnY3CPHqdsLloH6h
ae/tGdASOgee0XQGi6ifMsGB9KIjWm6ealGDmdS0eBaBck8/8CCca3AdDNgORFK5vJWyvRxflF9u
lCdAKM2CX4LK5UmlPsby/Vm3kDV1uRZ+MQviJey9zd6dy29scqm0GzM2JnefLwgkHn9rPBFvTsFV
fUCj+M8DUtDF52rQVd6SUFixF75S3cmA5mUzGSR5kVnfPlyF9uJuGmJeG5X+BviF9NX2ePc2mNdM
ytlTYMA4sSlbMqfo5+o95UWxMmNTFndpyojIDajrBHSIhalaX4V88qU8SMWsB9tAVuekSeq9sHuM
yScz7g/B92Oy0N6egVUXRcSEc/+T1HFlp+tIi3itEE2L4QutdPgzRhxrBBUn5/h3IoCsfzVuCwYw
7lw1dtdNYbUQwVP3hC8w1RbO+TOy1GC+CP3cmPd8Hg5mGG5UjkATY/6e7W98HXMwp74wSUOqPoY8
PSs/CdoOGFv8uYIt5NJZvtxekGGA13hyuxcs5xUcHG/yBMM+IyAcmH5U8UjYJO6bEE0L19YwXRNk
kkNOzne7zVp4q+Hy7NREwdH6RV2rhLhyjbs+2bw1etTrob9JPa643bwHD/xPv4asrUQLe2w6s43f
XscT57Q4OI+NhXXBys9PWsal/2vuXfThh4tZvGfFZQVMtRz65xItW6Bkao0vA9T0zyHvOgc9p+ky
0kczVU8PD043H+NBtbGVKFbAB9aU2FO2flOSMHXxljd0tME1gRB17U4gqM3layEjKUr7oM+5m5ut
BD6kTg0CgNNCNbiwgWNMzjl7oyKbHxgACrgJtcrALiVGZJ4vT4viM+TekaltCJSLpGULfDrGPI4F
RTJgjVool2daAyQERSpxutynozYw7t3QpogVxjvL77nbJ/zrALAvlH3eEDQFjLZFm4/zPigVdnoX
uzyCEqSK/8S5Aageicx1mz0ln6SPP24YC6JChmHRl9aodEoDuPO5Eed6QHnyznoMKpE5yimVwLZj
XMD7Igp9b//EAyNxvDBC6hFm631De23MPWhZWPdjVDWQz0RDxzF6MDHmY7y/dNy/z6JEE4WClYUF
BCyDLqoeUyWb0HAMgp4/NBCboG65c3NELJ5KIcW7SqSqiKzRliTv4r5328Y5QAV4xBBeoLReLAZj
7adrTXYH/DuWRx5BzL5aVDxa30jZZM+cVHG9714ddk+E/81AnMI9LBHpaXxH0mNmkmmQkOCvZcpq
Ly5qBmnY7vpOz/M+K+L6vx+FaCrdTRvlW7Hn4kLZJQxo6mDeNIMoy08O8e24wITNyu0p0aroZqvq
JKCOZSONO7u4NlpwzesiXaUtE0Sy79qkVmIp/C4I4/6kwOhclZ8W5wTeFKLjcwqUrvSPzADFc6Q4
1TnGtKXWslkBvvgQXEGDFbL6VMxIh0PStG2QmQ0x72AT/LVCD84Wznvk77KSWEsUQe8haxsnl0cI
fHULeXTzipQPhpO60jNuiABhmgKvLp3AUvOLmNX7dfwZWDrRcgTFsB3QcFX+QnXmBDyceYaZX19E
nFJ6sqy6eV+G89Kg4fmC2XwsZC/rTIE2vQm2deFuVMfHMBSxqA1PwPSE/7h727mYk8IlDn3vg9Xm
dKRuzpxDx4CzNDqsLwa+W5fTdK/Z3MnFer71+a2wY27UAcOOtTVUsDSV3CZPxsCXIaaGCdxKW+9C
l9vIY03YVbyvgurM11jrB+P1AACTLhtZs0Ts12okXI4Ned7Zx7cqg0CqDOyn5/Wdb2Uz8rtOUy70
ZwVXYvFXi3Ur5krAXTfD5N93/4BZtub7LyU92z+O2NnVQUpfHgWtEU/HDUzmgT7PPBx8kryxcZJ0
d62pynMAzrOUCdg8TezH/eEsonFlPSgJZXNCfcAd6FyF5nww3I4/LGWYSKexURtrBnsP0yhpAKD8
TRDWrqPWwgNG6NZXWV36N3qARnoKi0KJ6rR7SCux7tn4x9LnCA13Yjf+MoiiudfU5e26htgBIZF2
R6TbuEZqF12NOMXKbdw+LxDS8PodFgIALgV7k9hvJT8VpIPh6j9MsJTwyoAqy3Xs4VopZqSd9bzf
Wbdqgm7hpHK8XPYGtN+IKRkJQpQAnnw+8gBgjqiHu5aZAt79WZPJxPgJF7Xa1VFBoH39tzvw6Eae
GudlwbbWXfMW1G8L2/24V/CJs1gFdeh19c86Un24LavSDaZh3vGHj6kAuMuKZ6tM5rB/kls0f6EA
0ryFsqBp/iuvd+B3jFwB1jy3IYbeQA2rmvyAe50VUvVLf+9zxY+y5LggxldDmLXrmY3P57ekqxEu
/HPZ3UG93LLaRMNz0sOGMB/lMv1wLRYXPRRIr5/eDOUts5T+AKHgbOfBgMQaZLwbCVAuBgZZ3hNK
hsHfzB/OuMECR/WnFz8rcQ1MJHrvdkS4HT8hm4Vm740ZWPLwUgU1hH+ycNUFK+ecaN5qGEOT+Ro5
uacuj7tK0wpDAe7/St2MpxSUYF9qUfYaueKyeOkhvkKIygiRu9iFjyZa8IJUCgMu+e+m/8w7azmw
Vv5pBg3G4F3ybynkpPVMbSA3ll9zEsHAvnAG15ojAH8u1Dg8lNkTKPmT5RjHii+euzVUz2maQDws
DvrvZLV/w1EMY/auwjz5JECYGZLh+iNWv8O2PxZ6ARHeHlSofyJ4+DxkFzN7VS8kdV+zBRjeS7We
mIYRwbNwP//eIbfWYOqUU+254i+UMpvUrcDg8ZZQdK2I5N3AqPYOtYdtKW/IeXS5UKXzELMliFaD
pUgfYCxezosm43ow6Puep6XlfJAD93pl5wrDUJkzQceJDXJ99qW78ccBvSiMvbWl/Xf+nbl5S77n
Gbllwg/bhlAusX/LEbK2mS1zePwqZtJ3ruTCUNQ7fXhEKIOfru6jMN6Qh/NKEImYowGLgewqW2Zv
CVISIftpUkH4ySwlhKtIYeqWvscHIYSa2Z61Goht/7ktAWyirJD8hJ+se3RG4xS2hhJp8rL9426t
B5NVxSAYsCR+ZqB8MM4YvQxiwRhdB18idOyNwx7HpTjLzOvj9tKJztW0bb7iYqMur6iwLV57Boh9
P7ZySwAUkrVfuqJa0xefeyeHdDt3WBPY2IGX8PWAM2+526xOxwc8Hed2sQkojrMZwhVYHwczGMrm
UmEYFQlcdZGkKkxj8+CuWd3YmuhX+B9IY5bU+pXyxe5wfITnb13u/DvGYsbq6W0jHpDt6dtawNxp
vTDmBGqE+uhEubvHMeY+NV3OVnLNDkoywZeYRFLGOeat5KEeOuq8mLs5uAPnVcA+ZgbOK6uniuI8
hBYqBHZ2NHTif757OvVW4gObMEV1HOa/OkuWtSwyiepAPpJ5pcqdo0SUUYgrfzVAmvHj76WohtwT
xkuU1W3tP7h7B0TgUMZCU5JAM47WDPcQIRP/7bikexQ1D2XXFfIfl4pABXIsw4Mppu+U+jaOWy+S
JuJnpbkNd9iz8Mz1IzObKIwnFZNGPv3yKnHMRQsyZG4trbsv9gVddBRELrRovvF2Ce9GWLvS59pa
6wmzUeHiThmidPuasU7oCjz/wu1MNlg00lWZqE1vCe+jErHknPfA6lRQCqx6xZSjevE+qDu7Skla
Rp1RECh+JE0fQP2Za1YFKZJvJnAHftSWqRKp/FcSqZzkf9nySc4tjEudxQZhzN2FB1BuA6MQS0l1
0qHzUeW8TGcvHrt2dPeEHlh9ZZ1lvelKgL95N1DMkmbYyxfSILqqz9TZVJXZXT0KCTUyDFwO6rYD
J6RGT3NDNTaVdCSK0YAJ47z0zatriWHj1nG4ucVv3H0mWPr5TwXCZXUCEbAwNSco5xy/DRz8izKF
vJ8+LMQiVTniix1kTvAKsoB5msy1jC34gMzx3Nz/0Wjlg8D2Bm9HTGZUWtiu6rmubLR5l0/zHUiV
dd0culIPDDFJJoBUiCKMi362xBiOlv5bXujrStF6AFImjbJxBx5IDmyGWcholr+Afn+OBtxSIPyP
AhIupsfUvCYnJFWW9h4CEj/PvHkU2MErpogIGO2xy4SEqUiYI8+jkcaEl5hAM77GItlizBFJ5HcM
A/oIFWUqudwLpNlj9hRYEAYTiZkLYwiqN4vlGC8AkSd1Bw91tf76Wh6181it7NrbYmI8EceHg6uE
HycIOwN8F1YTDgjf5TxY/LedKy7MAag0NyZDWecMogmu/sOdnmrGEw3QnEo/kkiDKNXkJAum+ReZ
JdqPWuxTReK3Bi0LHwyEUKJ7xtqjhtUQQnKMmkxP2cNf4tbtfsxWEYZzFIRGXncXq3x/gJALamcY
qKrXuZgyt8ks9bUaefX6Bmv3B/wVUi55ijW0YklgaBBg6Afm/zeOiZoiWAEJcRSNGYUKmR/31+Ob
bNRGda44EyF2Rjhh85c1R3VkH0wAVW/ZRzIGPRwd7+XeAJNT+Fliq3WgRoLjqcvz/x+wFjq2hGPj
BHUlckctWP3PC1QSB9c/VQwIZdEAoevQ2WF6I/TYPmYdLAQVadZwTqt+6qkiR/UV/ove4CrLuoik
rIwhyXnFNgwCtpQ7aabKLG+LBNNZKP612NDTFKZJBuhRZg/j2nMsn7vweolQpk1Z+9B3soLo2avs
eIy8JBMqRd0IY645D9h9fIxWPoy4V4FQJ2jbufsb4S6Ia4HPqrbCRi3R+WiPi0VdcfAlibUFPqCI
oTX6MV+tzTSdC0u86FBi4O9gIpSPCaOiWUOYn+Jsn4Xn1tZMypPowv6wy2EZ7RpI5pWTUw6Q+ze8
FCNEkJQl5XGlcue5CgDEpqIenzR6PRU1CiCkxAPexJQoG3fBBxMi+jPIQj8d1/xjfBRtG83XsDVM
ZA+D4XvD1mzrdg2dFy+FhkYb91Vdjg/3iqUJ/yuOZqkuHoBc1BHCbUfT673fsi+1RDfdtFZVIxad
mqp5i/DtzMEqka5NKTLX3WLmsYy+kVjav8CFmz2fF/DzvlEnpQ2SulTb9vc7hLj+xqDMGdgMyQcH
5faU1X0zjWoZSkWaTyCWuBwUtKTRCgsg7FB3JqlV5XsK2yx3YyC1G0ZhDx0tsmTirQD4pckmVIze
Nc0mzlUGULD1YWWbb+iMD5pjUdBXCZCI0KLBuiAXyMIDXHiNgF/NFMwOgtgigao7eSL04pmfwBk1
Fx0BtX13Ml0Hgxs44eRNjMaXdwo7ZRGFXB0vTDwn81/JFSh49iM/q2lq85MTdwGzjKhrHzcoOZid
9cnscsrddE+QZbB9So4SNOb78UsKUB0xBSsY4u5rOIWY3M0xvieJeHejD17lL1S8lLgbMzI6ly6z
V2i7ZRjbQ1Z+YuFTGkMviCFNlmlEatckZFMTpjGBbWi43l3nKZStoHaetAhl9FSNz/Pc3rctbQvO
uOlh1o+wb+v7h/94PC0+Y2RZleH+vS7Bj9BdqIIIEFOTSB/AyHnNGoe2dCBw5GWjNjwEeMFx6u8g
GumsEqbgeUHA5vowPB2WFZ1k0J0FgBqZD29zxhUXg0erjjva4YJkjenvpYhbhCJYG2tqTdoKrpK7
I4SWdxo5aKUco0JwKKZvavXjCpY9WDBx2m/m1ubhKCyJqhZSCCbN9OygfUYAbx0Ei7/BXiOvDNvM
6191il9h6i6c3qHOFXZmyM4pycfLgkigNP6imkO12aB/UgZDJqFo1qGrKlzHjECbIPM6O6LVQbC+
YiQr8yyfcnlCQGoiZMYvKwTwrfmCCyChLsggOwNK2kHThCCcoWqZpK4Ty245YnfR7cWPjXm9yhZP
C8aOtVQGpsIGKZfbNczcRhaa4DH+MVfc/DPJ3XaHDytdNj03LuAF/9EaQkLc+UgT4iZBWFQ7mpjq
aMeFdr/d7wd/8CF8PjVPy5sYwzeH1xQIowpsikg2RL/8u3E9oMN1XBRYX+4zTpAZxLdUG45XScxn
md6UvYvMWRz2oOhQ9z0P56Dfmfw4SNjZ5f9z+xwrdnLyPbH6fueQpap9lkEmb18Kw8Rp1bkugSXn
0VzPmaqzEtX13/xuycjWxLyVcSQlFhKErP1tYTNB1BqJVtYS5Ik2cMTwOTt4KW8xddo+9NA3Tn0F
N68Ti0fh7FmIoKioelXyJy5A1Up35xj4XRIHVW0OcBgHSjq1GiIx/U4BVvrQsPJoelZTjcu4C5w0
Mjm2oli1/PWF6IhKkpz0yZ7B4tL5XKd2zjMbsVrYnlhrljBk3D9KKSD7mMfciDic/xzOSLuwwTHI
RFEN3pJOTkTj5ZXf9LHKnmBc3uaIr3wtmAND8GPR65EJBnWWE0gp7RoiLwIz8HBvoGgmFf6umgFB
GSedNwUl4NtjnT5L5ak/hBe4gxpCIN3+3gNP7F8y+zy2DcgOA5h6nESNPul5xYE5+gzLuami6lVT
f8Hz/swVxNimUSZL1Tt3XLNupls3cNEtQF2SWmc9ZH7KJLHhZSCYAATUy7h7HmBlJfaHg+VAIdec
WdTlKEWwrDJVrfS79OIUfq1lMbixsY9KItuu2Wh7j0UbxjyVnRbvwowq5ko1MK7nv2OgdfG67mim
NBrWGzzPIklSd/9utOd5KsWaNSnYpkwnkPzsoEFyfa8ctNmfRqeq41RMgvKWumv4Nf+4TXUsDQZ+
H2hfUgabMmjjpoT8LgaRnnGoiWgA2Z2+ZjPBEK+RNS1lgH0YETMRnpcRYv2Xg1gzNQEvJ5PWCyLa
QiwYLnubv8bfQsaaEO2U5tq7h+jT2BWsiSrXShsFslT82fWypi1rcd+0SK8e78aZl0g9KPhxKYzN
3ehGPqqrvkuJCk4T0y9FQaXCzEN3SD4naUDqOQp1xF/ZNrfoKYxMXqgNwFl8wqnqah+4WduyZiZP
bib/mc7zdTeIk6ZZU8ehnkm3afR+HdVLFBu4MHSkARrYfhjZLaJNLiofBou75VzdlTjlpuXfYgAn
uiWn8EDv0LPP575cURnNmlpVY4y8NKWOE4shve9kwxt/ez3VkCvpRK36gY1tC5Qpzd6T0h7TF0d6
pZlyhVVlnHgwGNvnur65Rqz4Q1S+y+4oIfpJbHyzXFO07Sm4Gn+SfKZuGJbHwDIZ4jTKWBYd7Bdr
VD2ul3EZdZaeUlANYBPYeZqRBYgtZ36B86ZTuDNun0WxxxfYP26T4zRer2gZxhB+pgmnhZg2d1AL
Y+I2Ez6KsOxLB3xwyOvHiTyleAG6oVgagJBPoIJLD8Sb3xSPC6aArrfAsJ5Etf6Fs5ySzV66GHEg
U1sRuRWmK6yZ1VWevnwhwmRs1ieffgek13yoYVTOw8YbtcLxUKeisR4kLQDBdlP3WGUu5xPtPa2A
y6c5UJs8S7vRWb7IOh/xap4vRXjFbXeSW/Xn0nInAh1aTszS+KVLosEbBZjnilN4fX+4ziDpTjds
jCszt00SxIZ58s7AnT1g9A/yg06h6tVn5wFkcW4PUXOphL9TG3bkt+TVjL84K4dM7clCHmhtHZ7x
pEjbVCPngIywX7vOv31Obmlq2T3XVX1SQUshbXenbSaYHJfyBmEjhtGfUjONA1Y/Tgcg1d0OLmGb
j4zNYUWb20A1e71wNYnGhZUBh2yW7N3zVJIIAPpolDxtF4RG01E6D8R+aqc64pZyG7nZ3AJaSclz
xJjY+mN+WwF0dJNOW+akr3A0otJyUvMlpXj5v5s6S7Mk9fKvZ5uFIEc8fzOi1BwB3lNsmcHWAsCp
Yk9Lh2ulT4CQGbYJd2P/1q/fNZz6rcuBe4BBD5wIvKHIxh2t8Y4m7XzPuq5pnP96ig8FitwpAOUd
crw9qSZcUGD2QBN/rH8YBRPlIz/FrjKHS3VJ39kqqGWqGwAbRs5gjBkWO1ZjBdP6CDewUrxfEA0q
dOVFbFwqGedBv2FzQjtcred6ups5/RqdeDfe3ThKyuZIGoXj84WMo5Beg+8TY7PZrqeHNkeUz6NV
lfp41YG172ETue87tYahTLHXxXToM3cOeZofJdeYCJEmG2UBH/hSzARA+pSEeTU75qoJC1fJa43P
C37lgL3ED5JgtN5yOR2dS46MHLCwAIKvycbBcn5uWkUcYalmQbSWFRaqCNQM1E4EMWPeAS3fTg/3
V01oPT1LKLOWU/aW0iTN+Nm54nJmRsFHF2LLcmpgcgg8GJdnqYr1meQGNuPGE7SaMtH7vPExsOje
I9zpiRWuhrltu0jQtO7ETRtgU1LISlHqgNyQbExtpLyglkpLk1/ZFOVUj5xVVN751Kkve8hQySGU
gpl4vnnPq2Qvz5jVPqsVNax/ILsESSHk6dWaAgGZy78d8FnzoAWd7ZN3EkUZGkAIduQR/kYoTROP
MLBP6d5rHqFqyxLm32FOc+of8rjRZZeKsccTsrHqsPYe+PjCLE3IxKtLIsBGdHXhYznu8BwVmrCo
WxuDUzRWhbdx/+1Hwu3K7xkfV3XAYlWYbijN6Ivq+U6cwro7CnGpXt0F5sWfHingm27aaCTc1RBD
oN10xwoSDPn6yUoy1lBaLzuyH2k8Q6LqbNK1U/EJVw7/5SMl0QqncyiNMlK/+LKC81OYR7IldrAu
fsBnnWWKjuc2Dd3iXCn0kvoXxZXmgDpZFM2qnrCXt+4Bl1qpO3B/AS4GgZHzFz9gtMe8jAM+3V6E
lnCXsXjPVd3r5+DO06JF6yoIQCEuW9CwJwTC7B3KHGrGyMkzpRwgvA4oDM8cjoYgxm5X4Yuye7XT
uz/p1i3MolE4p+1FsgTPaTsJ43ofJD4ti59PBAerWbxlG4OeJ0e8dFUz6i7mCxh2nF3kLy9sW+BX
PRRDFI9V0aLTRkRDBSHYsbKot7g5eZkubgJTMcJPVjIqHY+5MLWvaf5RoqL5xMtbykeN9d0k7IQx
57C0fEUlkm0Wqys2mwaoAxYaX+L1yLSwC9jlKZIMTjQ6AUonJl7POKYvQI+mmrIdbUV4HuCJgAFy
9yea9WzTjdHzW01o29QXyEJuNcIn81NL4AQ4k9YVIfz7CKW5TDsIDljlFsTCg5CEps/kiiX1VZ99
ANIjDbenbkB6phCS4dVDBqz/TZaQ1NHfz5Z3pGCXhlYGFEgmF3t2hNKJSJHVSsBWBxoDsOICh1nt
7gNL8asDDwxJ5WBK1aRs7gRpbCu+zVkgxk8X06Mo/5KYygywcqDqKcTeI+YgG12HJOOMog6nv/Gp
NyBu9clxeQHyOwC4mwoUxMQbhnVv9Kec9WFK0Q771CYocpG2cAviNZskZBt9Jd/6Kxdw3rOs765/
GKpnsnxFKuHGtDiDIUXQ10RlmG507fAnXLTTH9Zoyt8G/wtF0Hune9QIs3B+xC7zuBho1CHmXN9F
dI15wfslpAYOU3YacOKuqWMrWjPcC/OpFOk58UDm4Jcj3q47PuhqNSVo8SP/7nO9JCHG/6STKFTj
yxqYtapdj1Yc69KLStkWTVTdHfQcZnSJ5MXSGqhTA0IP0dHULzkCqGhtkk7Qx2f5Hqjrs2+wFnCd
sJORBu2SMfuZM7m43csu91d3+IUP1DoSuQuhXZ6tzXmkeTJ/rq9uGAiccxdGLA6fGjzFdGI033O3
EiSuj4IrUu5JH18uyEuomEDJ6BbmZRu+IllX9yt610UbFb9DDMvYUoNtSAhfWVlWzH2/ejvOTy7t
nhfccNMTixUh+PyZj638OCHN+O/179CiZxjmEV0dYZb0M3MBwqfYnScleSROTi1WnVegJn1VWzFn
GvoTpGFMaQEYXRfAjFLGz7Hnlv0N+FJjv5SfDrq5gorwvpYmnS6MbxMO8zgfCnzie2g6/TV8NDix
22WKfWIRRCNj3WjnYFEmPjpR7jfxn1GrDqqCPMvFdfYWsGyTJX+4jtCeIC9JKqeLX2rQNACI+/TH
fUZ+nxzdJBb7PneEniwljKF2pj6Sokdn22hQrkqZt6bzxcTzuviKiZ0ZTTflmiYkJhmgm5gxs6O8
gGtyORrcJSxNRa7BnIOwg+/Eca16jUf3LXa+ri8Pe3N41jENh2FdiB260ggttd6JUtFKpBvGChGr
jO1ZCm1E1yxDcaTalnFT5lKdUYymULclZinGIDh4ytd8u3/tbYyIFjTeg9W8O86LtKgMmS0k/rwI
xmu/2DPoPdPQUI0HoI0NGvvxlWfF2Tdk/HmpF+yoiymttaUBAlrFhHao7Px8/Z8hE0Lm80M5xmwS
4v8OJg3t2sNwJ0ohsNeRQcUpqGPZQ9PtZyMZkHKhsYw3bCM8B7NVLVdE/HJWPGyBM6tIFSRBsA0s
ULo85lPvRLsDa737m3OFS/EeSaZBuZ+jmiCsV4DlcYYqJ6sYJivdbDYPKYMrqmr+UEmyQVIjF03b
igftFX1zDiEYo2RKl9VaxviPuCw7aatRnT69INFKVXI4AAalItjc/DYvVKalbs1Cq4D/LgiWozqT
fFE3P5H/GjJRv81pxVIToIlDAUU578hR2y+6Ajor9AJbKNHlFccfHJT0pUQd8H2xKB0wJ32lxwZ1
PqTER5V641jBbNB2BMVUN+Rvx/C0JuxFUookibFMa5+jDDeKtohTIH6zaEbdGjay7sA7KKLgY1tC
15Ka8zVwju1BnyznIW96AIAOn+9oxvhnb5hZzfyFbyl5YORuM4yroEXoE6izmpSbacJl/MnVWsUr
vV0smLOMTrmAHLL5sevdE2eNFzCgeckv5qjffqssMtCRbwfevGocYgITYo+wQiKx1p1bUybuGgUy
0+eK2zx0nZflosGVK6b+Ldeuxyzaho2nkkxROmJYqvwpmjCxm6OQp3ahyjRCES8ApdlmfSvtD9Ts
qqR5WWxoGF/iQToouYmdDerFNbokJ9Dik6EfadANfLl9NzxVnRWqgU63VxurQGc3P3FFpLBFOwzC
t4TODr6gsvRGLN1igF3AAnN6M0y9MhXnxmdSIqYM1AkMVaWq1UPhhtlZ4ES1quZ7NXJh09TmNUQX
v+Gdb4+HP/qIOCH565N+qCLinDEcFnGrJnm5yq6aTU1Q/pF0ca7zV6QfJytrxFAetrRC40P5x6Xc
Iw0i8/52tBqW3ZIZvKWmCM7MCRfaU51q+2LI0U1nsj9bHOcXc9vI7EmCrZC6Tv9/b0RLVesicDxQ
bJ5iLl9yZwHadgjS8WNZ3rbgVB/HMe3vaU4Wtwux0wJcBzFFuZ9f1MTY6SNvJMLFgL50MtXZoHTd
n1E8R9YTZeb3bqZbBlrvd0hHB5SoA6E07IvPjOE9YXVfLOxXYL5Yw0+YOredMgXeiTG701gnPocD
+hh0I09/DkrloEHN7G7RW+IiJUtos3WOuUkDpizvL6DHLGxji3/oARQRzPOCKOYiQ67scOnoiuj5
10ZxwMctLbWRCA+8Z/dYHWJaU0UOb/koWlhmNCFbznqrz6l2LW1CWEo4DZV7uaQWyo51SAm+Gebu
E0Piz8gTCMQeX9grmjYZ+TCGjD0I3aWs4VxBqqvxhutm4SF91obBFlsFqdoj26JlNlPoYbaNGdDj
sWjGRFwNH2ff9tIXcI3zPCXjFK1lMid97hdqWLhWP90b99WnnRFEXXpgFCZUbOQiH1BfO2TUODB4
8UMfrgsdZ8fGpyZjkSskcMmiPuVmk00IbLUCwlqrcuFeOnBZoQiPeUJxtBsMhwQcx1JEJKJ6PHma
oEqrki2NWS4YN6BbT5HghtuaXALJVbJvyLZ1uVDU015oX1dC3vQxQnIjhQZe9mnomh5XbEI3aDbx
wrgLaxE1oGMdOyxoHH+tgA+iCwJL/Gfn67Z0T8Nmsg+C8AN1ZQ3WwyhUgiFCNERhwAHD4lJ5MPZO
DCE+MPfh/KqLBPT0+Ae5pAc7Hnt9kSOUAWf+tkoR7nGWZRW0zncrvYQ/dcaZas/e71HvZKlzIlzk
mhqK6JFDEzGSYch6DI7J//7BnQeJPok11ytM99su41492Xbk0/mATg39mcOSRD44gUoaJHzmZgO7
K4uoyJ3UUXTIjeAqwtJwy/bkv5+Cynct+sqmjb/DJ0o7+BCSFTTtZvyZRrGDARG+DczVUvHQfNOE
6ZIot4yBBOovB2XuuY0hCnQbclAJBpBnRm7GvjexccN9QGSJRIze+GgL8mdPUZWDHwlMKpxlUk6e
+qoCE+YF9uKyXOXotx4HKy7mVdPofMM/cSPwEDup8R/9/AaVYHXYuxQS3Lk8PZBzr65Kr+/83wvJ
mrNKnlWLKppp9Yjo3sFBuZW8+upJuf2cR0p+QVuQHOciSEhXdKMnR5sV6e+5r5nuESLTutRiJQuk
DftZo8F4YxBXZswENGYJ4BjhUfhilMJSDv43V20PUeitwTb4aA2OYYhf8RRR9R9t+yb7jTqLy7XL
vnP3h/h4lbvz8lH4wDFsBNAd4bXoZUwSKekVkFdggotB8EDr4p9VC0lp075tKC6+G4DkpH7Q3y47
WmckD2jSDPOzLx6yTuDtu1hrMk2Lpf4b84EanlljzsA66fwJoQHv6mdOqVcBLkESc4uR0UQiEU73
QL+Ughv4npS25C34jyWuUfUyFkwoO4BJyHP4+yW84O9Im1/pXyLN54tLmY0mwxyDEgdrQCnTVJ7N
0nJP82fHEY95ewa+eaSsprhfG9DyV803dLDia/shSJ3xwL4j3sAP5KEW4NVi88XUub/cHLVRyDZW
x48HQOcdMOuPCHtht8F6P11bj/E3K5iB+/5SZlIKT2/GpfG7Lu6u5cykmsxwB9+KNV2wghBXk83W
u3IzELiEnOjx7oA6/mSL+PXRyIDxu/FMgiCp/ukWTwsf+cwE3Jk2apowP1yKGRi/V+aLzFuhTRTx
lfYpRpE6lm1q7yFmPq1VRbg0PbdYSkLFnRvwdx6uM7V0DKDYw1VjULqWExjQYl75P/flN4WvJF7y
5E2cnwMt1J8XyJnsH9s/2JIV5glF6TeeN7fJnKAc/JSrobpNQjG/Chs8KzNgTZlv7H4AhwCqzEep
X3zE6PVsWaX3YqAoS+7xQw8Eay5FgLbNbJ5DwBpQWwJX89mulI/W/jWBBUO/PZb9PuTeGx4YbKT5
FdGjjSTxdc7mFciYQGhZSuA6nweOGt55utnKCC4txSHwInPNSddkCc/P4uuMvY+AVYXEI/5wvH2D
y84B96mmCc/RrkUQCMBzhyt5zgS5ABKcCi+sopd0WcU6hPhqUzfUQv3Ln8OFV7zafnumnon9cZ1A
GlcIS0PQ0kjQYCiAQByiy35Ld4MnKJQ8p48wKIgJZSHn4LptzAY5dT2BhUz4oByEAbOD7QKQdnWA
6UZA8itdOo2xGeYjwDCRNjzjvZGIdWa0i5O4jvX05tU52vu7OwRtKP3C2gc9vTOkT2roYZyVCwAS
uGw/i0iVRlPkXBY7KlckWaU/MC/2LUZopm1iwf/7dd2qMk28rpBsJNpsOGLi2Me04G4hl06ozz6e
nL9Vcn3rXObtuoPzUGIB6atR8o0rzoB3keeqvyH+sZ7jqIWa/UmEYKNydu9a8Io1qbb2NwKPVjOB
Ql+1jtP3jfTFgUNbFFNktTRdYU3tOr9wmRL57OVralCQnBrH2PKIPcpmzENSAItELG7l4iGvlEkG
roWS1v4W7x68Dh+UC1NiD4r4GBoPfPdoOLKra0xdzKOVpu66qljODlHOzwGRGm8c89ic9z6TwcXE
IMS5gvyjCy6GVvNIEB3C9wFTbPeq6UFQXexUsdKTyyQ1jGzQtLj719KG86iBYc5sFZT5NQnTGyg+
Js2h2A+tC+VAPHTEyTulWGoR2wWGcrSzbJuAc8FoMIyZtQq+Gh4T6NOnn2yPprYnVQux5Ybji+6s
+AHYZcPVI7ZTr14MRPnDqqHW+xZdWY+LpiRthtWtFaypxWTHVe25jH1FZl03y+xmAmrbYlDRCd+e
NZPc1dfPZbBzevhjBdwwD6et44aW9cwtptx/N8G/v3868l3oPKknQs2SuG51v2gmYu/6rkLx9kmI
dSbLf5xhjZZ50mJIXCxWamFy9YgcO1IbYxWvWkReGIT3Vl/a9mWYfDJbxpVtf7WWfUcfqPnfNv5q
pPcksfRNPOSrvXGGWmJoKqp36oTv3Mg+zK+nuZ2imnkPD/Lir2/zq1Ij5uycioHztDkTDs7hGcUl
QMDfThxpqq/vsEQxxum+7NYo66DQSf8ygdN3fiJRdoQ6q/X0LsKD6BL2cqpI352vnC+YDRdBjX9p
lJlFTvj/yTcYH14P8HxG9eLsU9MYqRwU0qxWATGVUkcoFITRhVgsYYD0tTCYL2oQVh5Rsg3fDIfS
V/CMc6id2LFW798UOB6il5qH66n53hXuCyza+1/bqU44rMJ7iX1pvCgh0Q3rwb3AIIFeef4SF1AB
SXIJ9YolQT6+Jxixb3fersaYLc7DoR2FlFNxQXkw1zo/YUxnxblc+j61oJYJeF1hjiCL6i2bzLph
YjM6BneeW/any5C3L63sAHTLlj1EqhMlTKKgGjvUzgT2UJ1Y6pxpRiK7gBQsX/3q4/9CTqzOorpA
yK4pEOflMoLQ6G1JxJcKpLtdCs1hUydFNDX0sx2hbK534wWlzcjc8yatk7Q1fIb+cc5bibLkYZC3
htc/DBDm70Q2WX0MrVEeWa/PFMvyo7idKTUfjxEIZJiBQEM+nMEwHAOSyRucX9UtbOA3dCn8zwzY
gVKai/lbbhgAerLhpL4ghctmoyGW7O2vfYxo86qhpLFk1lYoPV07VAPkNYfjRNfikEKSCJie3xhw
FIxn44J3R0xBSpJogmpTKPhet29rEHviK+GNg42KuxfZMSRaM89TKGzjswXTzdk5gEJwpoBVyrBV
2QVskcZrM8cJvF2dcfMbWH/wRPZT66KcnLogDgOcDcprd5TLLFMjuYdvtm3ZKY6XUP/Pk1VetEwf
xCOdIafFQyhPGhwzeAwTgMRfRVgNK/K0STZNY0wgnlyTIuiiW7jaWF0SeIMfwAF8q22TQC/yTiX0
/u08siiUD85z3+ug1+k9wQ0KyJKdWauL7rMalxK7v3SFf3yRxxp5qnXRoC9Hb33o69LYpzkm6+DP
V31bH/EwlSEl2HhLADuWafEMdrHCI1ebczV/EmI2+Tazc+5zMm8p+zhv8l6pzhlpxq4ISvETv/SB
p39SEs1NMALxKXHwUY8l3tyAOJ+ESoengw/1P6x55sZE1+2eTQJ4pR3G+wrdmKwg/xSre0v0WmaH
VZRd75Zs/56k01DOZCBxV6FTolmjvzS9skmY5fPf+2sk/rp+AIAGC1HhbC5i99r/WQSMeSwcc7Zo
GXoNvuLudmKmIUJ0reGvHL8t2Nadk6J3K+W7v/KX6jGAc4FMgKTNCzIC1OpwCDx6DfUA8ICvXzSB
Rc97YL6wV5xPvocXR13r0mokbKGSmkIM0cfNQQcw650Mh/C+7FEDVxzNJEXEHv/Hxa4Iw22t+IX7
Jx+PTEp+P6Ibrx7eAzhrBnWk9jjqX8WY99Q4lTWFpscr6aVfvyyJwrYz9DF/N1yG5vkxuTdRtQMC
yt3pB0UK4Are3vNReimlQqhJRQuK0n3GvijCvZ14n0U4Wf2MtDTFRDqPqRw5VNnxgj3UwOuio1Qc
jyWoT68SJSFPGLex6TOmYM0GBnszIamnWO5Uj6hdxGR8IUm2V/rY1TNB/S2EWvy7gdlCLw9QhpxH
EVAF4ZroHolHJth27g+SjQoKeYyZXJQ53TQfkE3EACRMtX/zSZIBKMJLDQh5XKbNIUlgcNHygrn/
0+lK5+NedTthtlgzKHT/qsMxjOE6UbhFm7g3WrzjdQtzBcpkuNcQSsXHxti5qbh7uwixwMOyBT/P
RWvYe4knM200hcmc3iWACqVPTNkiLuZGq67ukrO98q0hMGaqkTVY3Y/2Nzff5UFGhrzyJGU6A+AD
7M7Ka62zucQI72Irn/SrMBRxueAJckEOS/h2N17dZwqyAULt2Ylrf7KxMzJy5Cabzd6gWtI6PPly
FO6O12P3mIo8PmG4+AR3ZJlbdh3redSe202/k0VgMC9+KD+OCGxniQf0hQqWT6guafWS68sHRdPo
XhNBWVVJTByajktbjcxbtpAPA975jC6Yu2hs6fhQGyc/8clY4mMMgd12hPXL9hQ+KRQTG4VBhB4t
YU9+UyQa48z3VKe/434KVT/pFQzEMkELjxzWPmNnY0CZJWEWaM9qZ9KxTZzwZaSN/d74lh7CbE7F
NFk4sYRyVKu/yyu6DqlW8CoaFddzccrWoYs1HxWILt2UFaNYoU0OKfRyh2S7TX3i56ygN/+e/IVj
h24KIs0QbIgPZHFiuOaDLudFJZ7lUZgujlro570DzdfJRbNfZEny2GaXJkxzuidN34Kb+AT0X11N
ImJ3QVaa36yqb1H95+wTlu9DzVYhyngjtbLQ5hY3f7GL56sxAMz0leZlcT9akspWrJ2WdcKn83NW
xc6nVOOOCH1BxxPD43E93EC7/ehnWFpzm44J+cwQxXUTToHcHTiLdoBxdQw8w16V5CS58TQd/4+J
jaespLq3iTfczwrjRABj6340x/o/HLku+8llyCYJCwpUzWVHQ8mqPZayd8EFF08A0juBh3GL77eW
+eXz0pQyfrLjN7Xv7o28j8Gx9/JU9XMTYvZE43drewr1KX95Z9pKwmnLiBiiHVJ4kVC+/u/Wbmp4
H++jmSfNwggQvhZxFxq/dgRtyAUI9xOr64+2tn+9yMOm6BSwOSV9tAYPUQpyOSOomQtoNK1A74dh
eoQPCFYev5VuCeyuWiKiSEAIoZaY6UdwgJVRkntKk3ze4w3OguhibzQKwn4YdELKthGvE+CZ9alZ
Y4sVoF8d0GbkLqs6179IC6FneqLDk7ZiifLq4W0xarDHHcLBqogEK/RIb7jCM3lKJaK7Hp5ila78
7GulJrPhj+pq2B14JttAeAl/mpB861rQvOHfdZxZZZ2us3BbLM8mZqhYKWzLuvQQMCcknarXb176
bDaTaxSsf54/6eBnEOpFMFR0LkMROoj51IZmi7e9DEV3aoZRGDuL9nE0Siw07FB/OI7NeA/0prJ9
n6M5OrC0v/lWYx5MERCVgyUU98cuhPkrH9QoKfNw8lHUWNhUYFy3c355ielx2cYM8KMUMQl/s96M
1K3tovO2RAXfEyPkHflQKCqeen/dwj/Ug7jNruj2HsYNfGMN1qo3ARcGqQIVuG55lnN+gCTpGMp0
pI4Z3EFIld81P3f4pBhb7Kpc9jtfh/RKmrN+eA4daHwujEyTzESx+O3IMZVXHkGouy0dzxkAyvNy
f28hmY/SYvD8BQyCoQ2DAsqdgK52fllHwK70rzix03xx/jSy4dC57lraf0oKbwN9z8K98SMmP13k
U42+VDAlxpsvP53CG4XiN1fxwLwsNMBHokg983OjmASjzGMzjtXQ17URgGvbS3UYQ4sTcQeeWUYH
F3YxJ0j/X8YbzPdkRjXlRNQaoS/Eooa+2fu8DuQNDOoKXZQDcJ7k4+OnwJalDcazFJAVWtWUaq9s
jZELOoSLO09cE76n/Enhit0csER7XLxuzh64kCknEeGkxPK7GSX8n4ivFVhDmqPtCk+GLROQCjth
BMx7nvUNouriUiLFdO7oOn0y0lA2og0HQt3lihCIxg3tZUJovoQtmpIarG5n1BHfUSjCrJqoeASl
4AWobYBT/FJ4zTTRBVVjPf8jTRwxJsLTfWmxZI/nvCFHhyLssSuNv8/MwPqxhXhiHGAD+1/b1RPL
YTUrrYQORVatekECEMKVv9wcaVKNd9h9xLegY85B84rHfHSsudoObRX3Y3zjT/tVZuBUcnO+csaI
RpDJjJRFXWuWD7j/mgZ99zuwe2TuKkH2EB3iMiJR3pxr2B19JrApgwNEdR8dQNjt35ajwH1AxcJm
8jmd3sI0OzPmcwNC5mf0OlZRJmcTj/5qxp3iLGmSozBPzWMAd/h262H/ushjNtkAjzwrEsENP2YE
miH9vYBxUT2NR9Hlg/ODPAKwMkooA1BgHnHKlwAad4pbMK5xIdxkrI1F4WKmFZ6WE2D21H/6VZdm
djxme2cVnCoWgQoeCcMuGQVF69qHNVlqYyczzfICc5NQuiL4aipzvKPMnf1/Dst6GF/27ARelwFC
R9zSZ3KlAR2S+ypHFTW6ONOkFbNZ8DONRYHHc20DZzV0VQcVpDXZN49Xp8tdtOp1fSjScmhydPh+
dp3CehxUuX7NVmQCim/VsKKNvcDTSys2KcBxHjAlqFFQMd7ZsTV6jlesB6ClV4GLRG5RHaymcJl7
Fhs0qHJXqzL3/KUzO4JiEVS4ZauLFRooAR0/zcWx1y0PZARDRTVc9yEgUp7mdTFYMuLpOBhjvv6+
QP1juTz26WFwwqVsmuKRmq7Dk/J5qzEUV33MEKjmgKgFOXKhUQs8wOwCHHScMslJDJ53RHDUyFjV
iufIGXn5RNb8ggJYpj3BZUUBuy4kGOPo70RM0Mzqx1jWz+cXlSVHGocp51w12ObhoJTY/86CO2g3
UvIlCA2dziVW8Q0gHI23zbjZsmsODLsSfPa5URiTWWzwLcXifC337t89aS2Fde1KhJjgKpO6cdJt
C89lkCRsLO3/l8zm1nihrtnbgIKkhaZVEyyqV7wL0TdZ2YAb1WjS2XGixv0Xov+E69XQzIpfjK4W
6tLyicvxQocnNZwlVFZOEDxpsMtmJt8NVxUKgYw0GE4h0vo1ftiIkp5LshexsppT6oj4fQV6kN+n
955i/weTqsVWPWUjivx7B0PKa13YqVyYaauuhUEgLASzLSHXlLFMj8aI8mbde/HWPX7xKLIgpTDK
p5lCc3rhUjuiAT7DOtq/uU/IGOlOSnttc5KxPT/fQBvfYWyWFbN3X36U+bj0kNS7FE/JwuyIAu+e
980P3ZSXaiOH9jTrmITa/97m3WUUoeEiAb0WrjYZI/kwohCM0qjniNjeUMPT41TyEvXjm+zwD/9/
c02+YnYucTAQ1XZilCjB/COFS2iNVKPqupMNXq5EP+74O3pFa5P/WJErfuKUymFR9r5uukjHLE3k
JOnuGCcwxsED74jIqbY3jmVBWlZL1CdsyJSd78RM4TEvh5PmZ+tiBpH2fEBrPb742lW58IR2wPQz
yj5Qk+U1pMFGTlLEXXtknjvKN6iVPgjgjujgoFEN9B6ACDq6UIOGPG7qBwbxC9hGcF6dSSWz4Iob
EDX9Tijg7VXQQ0gKys1vusRrlCRn4Km0ZMZeugxCJrPhVDX10PA8ecUddZQoXe1OnyPdOtEz/Mjm
Hlep1Pd3kGrg1EwmcwNORDTS1tCwXdTRHsS3Etpxd2YPxMGemUhzwR98eCOPxM4+7O1O8Iv9266l
djsShktlui1WIjZuK2JDShu7g5fJ033/eqmpJGauBZPdohrDXihuHa5h7VsacrNPOYsFnhxoWpTY
1mKSZ8dnFxwFA+YkLEj1xvEOcYXWut6vyaiBFZsA46tzXDMTNlAkp/Y4I79V7s7rmlenMfezo+Zl
7nU+xYUkOfMYCpV/I0R6aPe9ind9fTa33fF8fGfzqlMRrOU00pFGHzIZ78u8FsUouXREj24sCjMl
HwOe1HhPQq91xTlK/hvGYEwiZoIpnB6gsEs6hwoZI04LgP4fv0RFUUlxwglX8EF09VPZIR+Uhsc+
4u8CAozWrKUdmygtD6kd2mliYIxdff+9a+xgSuhiwdbrAK+oBm79dT7C4Gk/JJT8prMDask/kJeg
acJWNNYtVp32pT+GqHm2yujFBube48AacxQFVMFxYuDf0mkYqvUXQqdiwSVnVD2RIatf9c8ryGKj
38E2r9+fyq+O/YbzNW6NwQiRqHo00S4HQGIfl8sE7LEGZy99yFc/mhlfWmxniOQ97SD7YsX7c9Z9
HOGmZgU/vRhigv0jVhhcHd9HRZKmsbYE9NwAGBVD4ARb9ccfBFlXRv/2Jh6Ck3RSrc7KTG+t7vh/
i4zpwjEQ4igCnbwo5WXDTKQD+RCL4dilWHOl4msQV1DWVtBhbYklNUJwYnQTyFgrpwYRDLzS4Ou6
ntilqobAN5vEKMgtnHo2kzOS/O1/7lKuGU8AWIWafmLGAxKaaOgahdnCSAUTqyyxyywLynFcFRyN
H7TYcfnThXty/f4pA9g+h+rLSjau6OYLWkqtTfqw3EZ5Nz+txb5ZlFHRRWyZ/8KhBoCe1N/1vhQU
KjuxfoqiG06SfsaxnaJjbEtcEWNVnFAB1PUIIae0n6h721WNriRYpT1KhIjPjdwL4xlwtGM9xDlf
uLmZvo5WknHeBlDa8JXdJijUXgu1tneiu1JYFepO6SEnSQ4v4HUy8OXEXEf9oYJV4FAbgPKnE6CS
CWzeJJNLvLT50bEaZ7+tXlAsRezZrjrV42O+faGheKXmysG/9QZ/q7IAqwO7fnWIp3GwMpGs92cH
OLjlY749STuKJggg+1sExWgsgQh8W9tFTnZun3eF+orcIsm+pgjw2I4bknX6gCtzKhfk6xSKdGpj
HKuCja/KwwIXrtOQ0FurbQisrxDXV+iSJfDBmmBLuEwFAJCQ5Y5xC+l/wylkriqWd0f51N5c8Qa/
LHTvyUMRkyzs19z/xHPZ17fa0PMZmSnJW3HCipEmY0oMJFEVKPaevJmhOqRiMkyoeQo/wAuVf1hd
KLUePtuWWjnqP1f4aEheaqYtNNgLmmk4kj6b00qocdKnrBW9+jRYGk6Eq7iEQ2vZp8W5mMGvJt6o
3YkHuiaC1HRYQt9yt6pq1L9tiV6ka+N9PGhL9RrUflK0fTfadxBDOpH8Rta+CWaK7Uj4pnahoJ6/
XUkoM87SVrcJGWHfksfPNLyoTX9bo7rg9tUMiIQ0Hm+BjwHH7gvYuNGapkstf77ZnSfXsrK3qL+S
637SNhmjT/ZhTwlB94KhOCzNI3XUJq4SOqbsLIOUxqNzjaFoTnhusbcxik0UzVzDkDVTv4ryCHCs
SNboDsiKNPlar/dpsb49tQHg06Ezagf3wkWAMuMbgFn5vujVKpnAW/JxUFjOPi0K1z6ZDI1zWE9x
UnQtE5phNQ2hWBc2hYPuUowbllk7J731o0j3knKT0jaWCq1ktyJvUUXJoi+TIMKKx7BFRdILDA5X
9SrUW8+HabuBlPNr/2OVSi4h/jYPrAZUiKc0yKXpsTKPwiB+XnH5K7HkJjl2M61gKX22hW7jeydV
cfbLNcmkjCzz+bwlNfwhjb5uDBY3YnJfzfOiImQBergnlfqOxLgx/Nl+A8LaVy56p9XsFXwSXGJ4
RV4WxeWQlE0Pal0+kl5gdbvKWcSB/jR6snSQNOf56zUdt99cjPyQVc+PBxZzK7lsQemNi+7zFDRJ
uEsZBDWqCa5V0Q7VLcd8PsLWqT7S7j4OFgj1GHeP9ydhckDkWq+Jct+RtnKiKC/CZONwWx1mTocq
dpOfJ2pi73OMiwcj400zzJ4TQkCQnmPzg1gFItfFy5PE9sCvU3mkeY0YCq+vH7quCIZ/4xDGtHjX
fLxsALiKKO8CPhTI+Ivz+rO715UqWVUke8acOoxuap/QCVEdLvmMjINVOA4BAqUDuur9q/BkxAlP
5vNFK4za+kLEW5iOvS+gJ7T0aIHjNYAxTCBwfyNwdR9V+K0l0Xjaw7AJVKKHnrA0yvzOkRZBpWMS
0g2GAinTiHD0XsPlfkS/9KZmEM/Ceh8Es3qlMGfgxsyqpEgG8J9PWzgiXL/0aIt+ax3jrxV8wEaA
ffbK2L8SD/ov4Ub3JFNqUqX0b++MzoCS9k+ZosPNWC3QKzlPyfwVYmFvfdylA/MHpueYBkUL1HiY
8LfwbKQcokRe5ykEUmtIfvq01QU/EYBZ47zmvIZE9eLukVjxuZQz728PmGHOCvTXBv8ZbvlPT6ob
hYfMWwGRYXWs14PnH6AxBUBp2HyQ1ZUelM4yiFeL+dZh17nR040JUvI0fcYbNFu8ox3QZRw747vX
2bdIOnHs8SErtV9YCL7AGv8Sl0KuRxkKQ1EVrxOmi+Z7JDiXH5mot/RrDTE2QBsAqmJWuYhYOjzf
ExG24XdEVD//KzcCahSf3hlxCRkLQXv4XhjPwDuDew00xT+He/xYvFmkGUlvQKKXIfFa8GytJkvH
M/FvFlLQ+dgmKAuT9p1G+BFPQaR62tGhacMOGJAD2/ysLemzpbnpt6aqEUw5miPuHDvU1SFIHnwH
7Mh5mhz57zSiBdXHAr7wvGBmt1TDKbnDDkivEMRSWl6uxmGqera+d+dQrcnHNy8wK715M5z+zLEN
9uowsqdPUdw9t+hCY4jhcXv1xBKgy2SCLoG+J69J5zO+I8yqCvvlihVH13Q2H+az0GCkADjgEpu9
ojP8FhXlp2cJnCwkF6NUwimJyDT0SQPZY2vKec0milljsqkED9W80FQLGssNQybUMrRNOr2xF8Me
VJCpIB13gVFe5NDAv96amDhna/o0Ett6wnDSqdczsqioaaq07vQeGrFjd7UUl91Bfs0DFGqu1VrM
5+isxLFGdo5BFNoB9xCrcKVTqkJw4eN6btLjbhmlCdVLM4ByN043xm8DwwhOghlKPjg/GvMwPUyb
YZ06wrY79KovYtmMdpq4OB5dF3eba9JkZyow5Hr7kpTQPPAoU8Aascyfs6+jnYwFTp3jhb41hIDP
6FkNHW+kGZnAS5SsV1/vbsdTEWfQUnN+ljgEh3sN/h+rDv+cbNdzouGW9HsNh9Dpu2VQwoXfVYn3
2Z2AihWHkP7pOdrm/ozVo5tEhZO0WAn8hwfLUm612Xk1RMloU2IJovkZsGaqNptY1D71Pd4KYEpA
whZtVV6Nq1POntn0UYaoKw+Y4U8YElNiiQOz+rqFxwM9koiTTxjsubUCSKtpu4hHUjcjM88ynKGo
v4GXcU5tFh3kIgiqY1Ih3G8Dmi9qPBjDGimHO2Uc/pTAq07yJMvx8cQyV/T7RvaQ3LM2O82FIROz
5lPgwZhwPwbKAWRdpx4UL8KPXgG7VajMZmFowiN5YRHeoiePSxto+ZS3ApCvzYGlBYHWM9w71J7c
1qvo9F4orCuLxyfa+/YvnTbOGtkxtnXxFwKyryvc+5jV0dFyNOe6PXpya3qRXwfeq0ti+eli8DhQ
TosZ/lLzsajWJS+JXiQJf1DUzBLY0LEY1n/Cvh2Kt8ENJe4QBcRtug3OHfsZZd7HGSHlt+ZT7z66
ChT9wV24HgoO+g4/qLVBrlnwcKI1PQ6fD28LOCRGene+qoWw7rBPtqIrIho582NN3NHgysUZKTpQ
hdNJZynt17Les+z+G4GfPVROSVbuGulRj8h4X9vtH86wDuqzJR7k1ROpOCY/SSS0jwswzf/LrgVW
8evM+pMtHyunJrkvYwH3bAAaxg5Dle6X5pu706HiTL6RBDO1B0vS6JS5LKTsTunKLjXxGyjdtG9W
o52gB9L0X+QZmiP5tD2mMnmvZXJJEMy2t0euaDxPGocIm44jGVWxlevJFz1GNO+OxE5rGeXMmGrf
1wgUMLD5OVsYnweGXbXUegC3vqineF+pU7XCo6NcjF7ZkUywwGHs8PfThYGd2RenKRtbW8GvIaPV
hDDsH2ogr16nn1SGFKJ9HugOiiUR4Hud2hmwZEWcy1rkX6OQweatEIlbxwg8aouNCBaMcK+peEzW
bZdZSPAdafMmY4mz6cDYlMKpQACdEwsI9/9EJ2MeDTznXFqw6oE7wduYkBOg6mWkDBvLAUu5EsaI
yxUc2jGasR224fYTXuZ7m7eEzKGEwdpMfT30xrsjS6BLyKyO76IIVzETrGiohv3obc6w0GlNNy2k
jX53rGfAkuN6rAaDUGCZRbT2STt/ALf+wgTeVZl8RkuWohJBIIRBxjWCvtrJ24/xdUeDfKj0IFJY
wMDaDF/MH9Sc7mYuVuxjhUZ9bKMW9dMFz4aenGpgswSiJd0qWhMl3o5pabzTtXhWDelbyaR/1f6y
eV62Sk9o8O8ycrUT89iBWiG8qiqSIBit1vzXri/pEO3dfUSNlxXdqyM622sGlIovYJz9ObNrTnIY
1RBVTN08/0MvwZFvHPvyKnFTK9Md4ix7az+KD2GyytBRV4NOT+FvG3pYtxB5bM36ISNlY09zEnTw
EtjQPkLBTh6lAT+Kl5pDLOmOks8QCI99gHyV+9dKhvqybXbp0Y4LcgjBHeqn+A4ZLNkoEIPcFYLB
eOv5bK4R+Dc9KDnv2E/OKkg6kOiQKopWFULR4IS8kUNNAzVJnh/KPXNowOU4SkXprn+X1CFmcO4e
6dPQFjvCgh4mB4Eu77VFIOjVkdRpiY2umZuzR7UA7hbypK5fqpMsCvCjbY8RehXkRi9Jr7kfkCtz
FDaSiF4YX6jmCT8H2XHVOT+WZimfmIlmxfp8SHS2JhF0swIg0XfJ8PHaiIO/+Uqwoa/AkLadLL7M
v+wTWUabdwj1H9BZzYp7ilU8d6AscJ7KeylwGX+g8JBykTapnVrONqV0gKBNcrJOwEmtg8Yu6xap
3W+WHC9q7dGgpNFrCI16SDhTix0aaSB52M9WO2H4pB17UgWcHRQ11Kus/d90DIV9rmu84IQsMUoZ
lFomu0gB3LjNw3IaXOo+953qzarQ352sZUGWFMj4btJaar76KO+tkbs/UTyT9MdXFwRbX8C/s3vL
yQ7J71Bv9ha9DMWEMDxDbOKXo4UhqDeJgjF+dANL03EWxfCrm0hYjpxo0MFeSIu/hts1/8Z2NYZ9
c88rfmZf6J0qNMcE4WeGKuNTBTV/wFrmY9FUgfiHqH/U1WyAiRX2O2ZveL9ffakka1aP1MBLhV+7
vxtvjSuzwxL/9e6ZG4o9SvVTyIV6jseua/E01Tv8fTQ0S16uKtXfodtk6CXCMqcHL5N4MKWvRQV4
afph58Sgl52/67+iMi89Few3CtthAzG321CRg5FpP73bwmindM58KWBJqsj4+PWBI0Mq4z+tE+xo
vUItxaDiQj8sKjVHVXXJ5VuyalgWWcyfMP7mIRqbMTen1y8unAo47aXtSY9rT3pi53Dwz7QebSG7
7+lYWEqXQFsTx3BEEjrcaEbofPHS4Dlc8QGSQqSX+VC6MRes4OxCjMOXUS6VBKtrbDaFZmaAi80S
3kudUot8CqX4IAyissi66qQF/0tUfs0QN9rFiks4oORA1quVtJ7CSGSC+J0P7ORZQqmJmcKW/I4g
zmr+cvxV1Pdb/KdkBhjpZzgIxz7dUF+/U8e7TbGXbdCXs2vjQew6JHcXQLnH5x4rYQoJZYF+Cebe
lwLUWw+aG6WQTwhoQGSzQJvBik+YRSz9n6h+tGyK7c4lKAGiDfuY2HdN2PULkm6DPpJexNdjz3sq
QfY5UdRj9Ic4vcaxFltpDem1uZ8ikNk9FUHWu21vuoIEquD+CAU+7XzAUW8ZlPksmc7IpY/2BYzR
wkQLu1ND34mvVNI/Y/EJ9vbFOqhV5byZj/RSvfKx1QPjRsnULd3L6GOlF51TwpfEm/oLwHBurylu
rxcMrHYY3cHInx0l8KUn3qzhz4Cu/73z+hbDbZk5K4JK3clVZADFQYRPlluiHj7eCgaOfGrgHPlb
WRDDMpmJVNwOObHaRjjRWdyRA3BqZezuqqicb8UC7qfAQQV8+DrsealSgCzH7J/cANg9TUpk4zbc
FwXOm/A3Xv9k9JWQQTYoMUengeCMVf0oULvi32QmC9zwomtztd54spsw8anWabF0ocwcjM340ykp
YPIHK/6y4A7P9vIzW6QPXqu6ScmGHQAAPA6eGXlYRp0dJofgC79+atJOEMe/JXlp+kIiVXkAAa+A
GWc65k+KlE6SAKF5GHGDFtuQptxxJf0sXqePeN/E2wbo8SCEIlf9XYPb00h+4+cII6lTc4PUMChR
eSDkiEzD/NMuikqIcXrj/iymRD515xm0suwzQz6i8S/g72tc2dcY7ck39OZhmLiBlBbUJbfp90xa
asBmMb+jpdtdUcNwfpUJoMK+QcukjkE+AcC955lp4zllQGUgSnIEKD3TMag3SBX/d2L1RR0xUcYu
DFbWZXRtGeddyrwVBCuxMcsFb34eR1i/yXccitoub8eR+DqzReVF+46t+8B3eS7TzYI65V5w2ESv
9IBJNO03Culd0Fdwj9ABQ6xorPtRX5nUGmiPXVXa8rn29YOqBflwv/LzhaGYUmx7+EjhRBVlAtTp
ePaaGMQ0NSLiSYiE79Xe5lEZ0YSFWMDB1zusePpoiqnlpF0avF5ulaQXVxxOaEu3BRaiDyEyuxv+
3NVaihQDF4+thf8i15EjIuZKSnDvRAmtqVcaOjthiZnQiRWYDa+n7q4C5dYOCe3DMwo+c5GmFd37
FRlm7abrbFM1OCheCv4CBK0okUDRSSFwSuoAvzvNiVyeobjJ0KB+9NRuPy32o8L+geJcL7hcUL7S
T9B9hTDCulfN3idNBCYogotFQqJzD3CsNFl4LOmmP465Yb4UpgnWnQljgC+XwEP0Re15HxCNm3Zk
mhV9OE/FOXzMVLjmSv3UDZwsH8q1YtJuTLqP9iOG/oNNb9qnFnpjPNPmSxSADy70Ed9z+2w3xtUR
vvVQFDTIqhhgPRkxqIhpLg9xYizGdPpVGwA8G6NA1z/MwywAWfHDQ0kXMiSRwBKYC6tu3j+u/GAt
uWaCQ9uQg+/qKtR2dwjkjawi6LDaHJBQoppe7P5FNTLMCm4bPgdVXDBJv84AsfEwxsglascHRCbq
bqyNuimsOocsCloNYptEt2Ha0VvRP3kGqtg6Wplvdiks21v//8iiqJtcPTIWGCKk0f6d2EKdw2nb
xiUBjIez8fTuWar5bI8koX3/3inzJdkns+ANnWQk9oOgxZBAlMXO+MRPblwiagoGSK6ia1yufG1/
UvWCcT+ff1mRvkW/jMhhRYiDlDwBts6l+/a0zYbDqhxoKFlQ/PSDNeMbOGeFRhVz/PIbR2ldTNYR
URRBd1hXXGwxV/gvZORgb6fXgvFvCgHXLBziCEasInPWADmRkOFxRLXfLBscIBQfdSVNb1WT+RQ6
RMaQopCbJ0qlewmyEMceggH/VJpT9McgG2jkFUwb08UC73mMJGBonyMcxC0HvH9WmmukhDZPVW2p
dWqsDuHuxoQMl3eEEazNkk63l3DIcFpHYdguVBUmmEb2R+CmFsT5HMixpMN0M3LWaF1AZO8PKMNH
XMYwkquMsYaoGnakA8FALN0rszybq6SjtLWOM2VyqtCEirCmOTvesa0RKgT5U/BPxZNTUpoV2TT3
oLYRHFnq//r6Rt50FXQi5gRqkzDyQoXZzzrZb9z9Exn3QZcH4S+LxrzBnjpcIsWPNg6vebiizWwq
h8Dr7Dsq63o2MfCJe3oy32ZQTVTsveCJkqGzzeOWPKF5S27H4OV1I2IAS/sv/4x4sBlgk61oTJyP
eOEqBpsvB07kUyf4s1/34p4qow566kGo61Ys+DPnO7YKcbJQZYnt8oHMGmHsl27C+rbfki42o9jp
bxUNyxK2o7cJpO8B/19E3J9yKNIE8zTjbCLomwF9MuFAWDfFxQD/035aZYBqakneICXnoD0pMZMo
nzTQsztpparfl1Sh1zcTllOrnGmvtdRDN5+axr1eunuiYOqGyTuQYsY/CrOZI/1n87UPYKvIZdCb
OdoyJa3553Gcy3V1jZ5XBoRTEFIEPIS8QFWrPw9PpqLsEUenbHCocJlJhW64CpPuqdbnVdgyqAx2
Wvw9N+wQ8qcEyuxBylEZ5juTUoW9xjeVwiKIH5keVyyWfKpY/CauFPq2jK3EzSvN8+9qwK015lRU
VaymBH0Z2N7HYGuMGWOuIQ6zi6nycXyx+xineoxwLd0okovOaXmvGgQM9sinG9a+byWzH797IL1s
bXMjkjaxOr6zLx6uguk/yyqHfrbfGOsR9VRIFKLt1tvkojpxbRNeyds2rCZA4mhllEC0Gc6WHxX6
xeWHxAu8b1nQtgEouM26LjW02s77+LBZzAKEWryMeni/9AkN1q7k9SDMMU4yLIOAA2vhQq31nuge
TOkW74CWpDvMlvnzl1bhesHkTaedvLPhCr0jCH0ZYPIlAbKQ38a3zT0q5fMS1I3UpAJCieyK1soh
S4VbJG7AOCJyEeoXmuh9dmeFUyYyJYRomAVCDq00OoPGqhKmkCb/U28R2DGBh0Rkym2M1k0GKWmu
7NjfILSQH4ox5DjmbMGWZqNDJwJ5pjWHFC37vNoa0n7RauVwzsHzs4x1bY487KonRL5onXYJg7lx
XL+G4cFjBd7HlQl5KAeYe8uvNdlz7Sxn5CQoaigT/6CTdfvkkcD+9QH+viHaDOEQbp2iu2l0DcFh
3CrV+NKBctedwXtwjEamE5jZKqvaMpx2p8HPP1EwNtzwVyazSbPZL0Pmm+T+vpLt0+RLUTz9dlp2
YoT6CC66ox8hMJx+OMHfT2kRtBNRfIvwXW2BlLIFrxWI5867ZFcAPUr4UR1jok5B5vi4TDXE1Q7A
5jVWVQIH2tC662Spsd9Vlz7TkDg81HuFnf3kxBF8glzjIYQUubX5ROptqIbjJxxjpt0GYd6xcrTY
I/7iaK+qhwyBVGij+OoMNH++LQz40FDcTorvqB+XFcKSj12zFDqmWKS8rczo4qqnNGJar5ZiNvAi
RKNrejRv8ha5GCkS6stPyV41pijB8K8P4HpBD9ayFr8xGyjYrMH9fi7VI/Hv0quAKUIp8upPctue
lKUHVQg6vwvRe303jFjfer11YYePaj6ojtOPxVNgs18+7TV7MxBDFRb1IHYfsJ9H24WOplH8xg8a
F2ZwhkMsfLRIquImKu+8WXhj6qkVIALppjGHw4sij+v4iphcCX4k5XhXtXKl1viWiNtJMqM+FRMm
11WntYhko3oo8C8b8AzeBDvb0BTzFD9IqFHAH8jchvePNwmPb15rdgQtogAnOSvSHIKQ0p7ABJA8
w2HoshzH+V5kBd3wJ87ohDAGHuLyYnbSsJAgJdd4XArAcbzctwp2ytyq83KyBJCUyduKRmuRKVZK
Z1Hgihfly7JT4Wip/elrnLoZ47P8CfkdS38nh7jiWcfeFdIwN/OZOjuV8/dTyU75rCjfutw9D8yO
7+55x1xxZibgBPd4D317OLSbJRs0vrV6PhHLJRsjPVL9sdl2PW7rQ56T9pj9TYnfLN4mUipmRfRV
5OY+05lB4Yg+SZjScZUff3SHbLtl9FDTzGN/oLcUuSEowcRdWQowG2Pp5JaFFH6jmY5b9TmZNfsE
6wmJOxbZA5KBqZ9Wm4ESwlqLSsW9QuJvoQuccmALRlnusZHzfQmGYQSZMmCl+kzgRmKCvYzkE/QY
8bQUQLlERiuXmuClkxvwGqoQBdXWOG+Gy8dj5cBW+yvVijb5Q1s44tor5PzWsvdEDiLs7nih7oDe
2rmElqxgF8OyyfGOa3ftX7L3ZPRv9HCi77XwMFSeM29pOyP0R8e5VeMmk+F0E4pK/a2Z1xQEp9xQ
6E2hDO8ETJ5hKx2Y/9YUlkzWZdA3d4Fn/Si6hlMd1q6iRXKW1+WdMZH6APbZjNMvHvGfkkeIdkWs
In6xpH7D6X+vzl4GTGI4id2Ju6ERsArEntQbJVsfVsS5u93/pLr6vzUbcEu1VDxwPPTaic6rYSJW
T86nFfL9MuFP9NOToNDJhYcHDWq+3rwPNIrA1rZvQnclIjlKU39qVGHbdy5qrIpchee5uhjTwJDo
G+frBpov/AhSgUVLofci2yRhB13TyuSamZ5n5u1cuiEHYnWlt4Y12RkHATB8abcOD3MVNiivxO37
DgMDFiW1Gfzlqt23mJMnC7LUUWCvHmNB2o9LRYWA9wtD5IdR1K1YwcyoW9zF+lgXjZi3GPhpRqpl
rKeUw7iMKzo3iDM3XznA5KozF4BC+KDCFfkPIDo2A2NenSY8CaJ13syRfFM+OTvyV3og1mgV4CXD
c+hQOPY41EUAyn+J4HYRQRuHVYhCq1dWRGN3pYYnj4VZKNwqMTVfNOP2ajSe2TuP5ocePUgT5AhD
QeZ12rhhvBlam5rQGCDmGuDG4UESdYUUbp/FacAK0Lsy5rVFaD6vo0jSEU9WHsqtQZI6FXHBwoZu
J8Ed4G3v54txpYohLGZCfl8L4z6D4pOFPozS4g8ezp0OV0upt0D6M+DI5Vqam9Hs/ZKv6HZDievN
05+qMcUqSUdk851O7R+9eYFiucfj7kirNW+dpIqxa4Gb6M9WV2AYns3zOvBKVDTgW0B/vlZUJzM5
no5pDeSUvTUgoHZqpBlJirCGJdvCwyOV9RRDgZ46DvgK0cIZtI60o7y7W44Z3BFiXL3YGL4sTDQO
3pys69p3nawapAUYmHzzX4LcSxVaHzOopsCXYWvfWibbiSJg2B2X1cVf6pPGtaUhjh9wKt+1x0//
TernCgS52jYJlGrveuINOWFCdBQ/tHFlJj2yP9u8GJHGaTpUZgjT0PW1TMQpM55gPkrP9NW3tGPX
RPmhdLWiTztDV8uZe3PJyBAr6sRGMl+yG32XGQZGvFWd0A7QrVvp5KOUR39mN+78km/UPXUsq/kg
Z5rLZZ+3IUi+ZeZ0NbtvKworfxWTwg+WYXEqZo+oTmUuweay7IjAKoPOF2y18H1iNnbA/aM/uRb3
Of5h7QJH7p4DM05scymlMGBIAr7nrllfwl9pVSxdAHqtQLNWunSj3vWQ89UoLeelag5UwxOEunr3
2dpt2WeCkdhwq5idRP8AMSf8LL9N1GgfKnksFSQOFSt880a2S/timR/drRblFNAuCVRDeANYPTIq
xOhVyYiYBv5lmGjP9h8JJ8PFl0ZLrNGYEOW1WIc4/8Lz6sguMgPKXSlI4X2nd2qe1nJuju99u+/1
rsNGW/fsxufZLXVs/O4j4f6yM1FHn5MSAefxFPwT10zxQ0nq6hdb//awINHM7oZPSi9RwLFORCS0
HIySD0atZSy2uUBClilqSKugT8M3ZZGE40/bd4r5RlEchVF/XRa91fELeEzRh95Y+cJZIdzBR6Hw
QLVpfmJNN2j8YeKA5G2tln3ZymH6Z6dS5v0NpL+YsBMBYwq4dEOub2qUMVuU0G7GOSrZRWYweFJF
1Nzgdts+LX3lJ8luZ3iVCF5upudLfTkOcgBAAThZFw6xi13k/J139XZr4sJXZSSlyi+ltFhPwNC5
ungu6VgdYLJijyG37UcAK7WWsYzUSO/zSiNphB0eOx4k6+7Fdz6obar7KDRbMpxFn/XYa6LS0Vbu
6LOb9u6agJjfIgmrelbSrRSxALJ/kfvrLmV+ey4vxR8sJ+iGxVUcpUnuhwiif74aka+bbMvyPxIV
smrdhD7avXD75dsuyfHBaiaZsJlQwUeo2DPtuh3dztRYJUdYDaeJ56ZO8IpwiyYjxazgYs9q00Fn
wnOkc+Eqk5XERRbL6jhmPA4l571BpBriuf0kinvc8oj6uzKaajweH0vCwYN+3QrUJ2lXD3l0DbTk
9YmoOwNFC8gZ4+0655BC8efoxvRVRr0dTBYuIgo1N6rjFT291s1mcoVejGg8/IZNzt7YYh8Sc+Em
pXt3haZoVwnpFeXnKIc3X8Dx1Qx7PuCc41Sqdo65Xn9YfJs88ob1PhXc0RXl/uTskATsz/H2SYeb
8VilozLEgIjjoC2Li+czdwg2/OvTJHt8h/DicYaAkcz8g6TB/tyt+TRrvt4ks9pQpIp5Owaeez/2
Dknat0SmY8iljTIiTMUrhZX2gEsWMBafVellqWMuDvaWNS0w3kbMBcd+Z9AZt9WKsEYJLHsFF4tG
PAETccRYUGLrmthaGVcqDujPhSpmTCRIcOsJpdxmoz3iBRx+cMeU56ZZuJcjl+LSCP0a/B1SqcVL
pYP8b/ix/VTTA8zIYheQVzMMfFno1MaM7Hx63VNL0+ocWStmahX3ktB6mcmeNZ6sSRsR6+qe9A3I
BAvE/BORbu2WfM6/4BAhM3K1NnpY4pjmGc81BsXteoM3nlSerjmYKjWNsT2qYqivNnREb0PdryQN
KmNJo3qnQCZoAZCWfd5pMuulEPtq5APRqX8Lq1ktYUSQAjZkOe83LaozvTRRyu315mxyCLOXbd8q
776LZelIMsnmT7x/Z4SF8RUqrJ7exEh72+94IpJ+Sz2Ao1RbkVYDRlr2jDVUD/jJuYU0yRabOo3C
lyBGoxD4fFuVLB92GRBn7QLDJe+T7MVaK/ZQAIw6P0t65RNrP8dHhHtxGydpoghFDvigaIDrYeBy
M9PJP1tNmgATbkQ5jR3SME4hTtAraR6Icalbyyl+juBzjYTC/ITpPTX/BSmKbhHCEic9DREft8Vo
W3VpfJaZw2TzZIpDsUzZk7KYp4R4QqAa5pxpVnNH98Lj2TDr6pn4tskdAgLohQY5UaeODluWTqtK
C0Cn7i9k9/9hW8nxSZJFy9nbwqR2I6+L26LGZEN4mOS+KVIy6SKjFyxHUXKXfm7Y3hHpp+C3BhFq
7zYFbm/2tbtBTGDu6A3RRWPKTOaMy2mKBBhi+Hwr3aOyj/uQkP/5XaIa/A/ZRSe2nwtSou4fUult
VbU07hHdpJ1ZfHauOgDowbw3w32U8EE0MFzrlj4F3LGrzTn2CBYUzqgM5zmhQhI8AMFOylCqGlk1
1KQCKjuR9/Rzk9zkpgRiYAK0u4uN1sozR0b1YUcb/EOfG/VMYZNIvvPMisxKe/0EgBPcgSY9Nsa9
gyfCCRd0dLIA+7LgVuYP/sUeLQTmFeiEhi8iMdzvYEzsSPo8SyouMdvZwKLOwJrrDR1O1Dp3c1RA
uLgfmcNWd8Zib2V1u8l5FZG9a/Ohlt7VKtgwFF8N2wD7SKiIOMf/K54CRsgo3LI3thbxGP5bUkR5
qMRLTkkILHiuFYvLDW3209IEEJnLqDmNqH1bAOXmTcChrTTEJmdTpsVp/AMLbOQ/LiwjF1gU1/TK
+RA4ZJrrKalmcb/rpcAxu1HPWnehfrGbXemgt1eAtwkdq8QLhvzOQGQNRpx0dZKeRpILTruj3lcT
LqWqq2xggjton01ODGhWtKzdq/ulsXmes6t9ArDNymOTkf3a2SbJ1n1zZnPTNvQhH4dbF21V6nOe
LJ8AqR9oF2M4X3Oiqtkc8eQEQsBd1fmQ9bS6vIsVpGsZLX9+L1PTl9R8PLmH3tANPRbqyqe2O6aQ
j2Ib+gWajgvtTJM1PmorO3DuazhjabPJIGT2V9kqZfUTcJz3W/a3EchhCo6T/0dPWbgyv6ZOwXlJ
evYN7lHPwkeOWdkAP1bEL2TyfpeEH/pJ1XaKhESOZ2DR2XpG7iCsAUvElLsfZmVcSSskpvg2+FEC
zn0AJ1tbrRJFt/QYImt504rzyZEEdaSFkGcq59wvaQ5Bw/8UpeS7Ny4NnbmAtoC6Qr4rl/0EN9qC
4yHI5J6NgEXEgvuDl3ozM8XSSb9zrptwYNF9mhqSgFJz4kr/0lNd8bMvhReQGHLv/8ZdEgr4Tgur
ZxZkQ2AdcZ/3/rosT/OaCCtGxiR8xZ0wNLxXWYWzr0Uu4CBVnEr4kXU4v/JX6m+4SFiKcqh/rSy/
Gz6ms25mYB75KY0lXkO2xQOSZBbsDPNgkTAWiFPzvKM5iudarcY9Rn6xM0a+Aldphww6P+D9OtuQ
2cLXwXNbPZ5FyKdJtHlwJt/B8FZwGM0wBzm4kPIcEg8cw4nR1fQ2aYn0oOJ4DXjjjt4RCEXARa2Z
iZy+1S8SDn3mfXTJ3AEKwnv7kGWit3wU1PMmOIblcQcXxCu2kC1/PAWb4iio3jyVgerTtjcr3Jck
HhaSWgQs3vWLDH4JkUfEyj3dR2gqrbA2JzKMEij9HnxPdZowfH9vQSE0MkkeRHn/ITR2j4K7e6LW
ctHnMjjPjmBkfFbMjc4kb/1uPC1NpjGauBK/JprMzFISIrcGyYL+kUEcoGXeGMsVQXypsRAjOCJF
SCiI3n2+YGOQ6XC/cRcnu4TY41HoQI3VQbiECmmR6jSiyBXozJ7wswpyqLC6KRvNChBj0Fw9/Ad8
KZCJ/IX83ydkN6Ssj1IHO45vEjSNYPyN2WbB+jbUKwQvSkelOate6jAry5JismIBdrSvuKfKEIHT
9oo6AvbOHHf0zmvpjmwOzzZND2GoRhBIAiN2MUEEvLXecnWT8qI5y6fc8Gav+yoEDteycKh/m+/p
aDpGiTmzVDPyhRMBTYIfks42lKdKGXIfF2p1/9Cyt6xmX9LknqE5WFc6eCSLGUMqCxi/6btIC0h0
lhu8H+UxR/381yU+g0VGy9cYkVNAWOpzEVF81ydqw794W9Fy7arhBydLLjgu7bng0t/k9ei50Do9
jXuqfjRpT/68gTn8sbJnK9eBifc0rLeGK5AcOzhf1zhq19QazjgdgYdZeqnD0dGXu93jGsLLArgM
HRoxwxCX43mlQ+eYRuW6tu0L6ORKHi2WThjfKs3J2iw7VwxQepsrQjiaq9+l+QCTlYbpAncPYPuP
UnnhuRLDpcELLpgOp9K2SNuw08XowTzAMl9u3uqZSun+TuJQZz0O7todPCKC7RaXGcDpnvvQIGZM
gjai2QwVryewgPm9YSMY/93ABpWu9nWytMqUSQgX3pPAeVL8HVKj9v4aJ+9KDKilNOW9hc+GZtik
X8ge623J/IWfR2I6TXZf7qMDEswfwV8n/4QafWoE5Iq5BqV6O9+ya8NAGuxAhl5m6br41fv59e+g
XKsKvU0xP4Fn2h2GobGZcmk8yye6qWEKyXe9lXPG1tpooxds2m8aX9ToKyb6jv1t9GcaB5W1l1OI
1vLrmYlCco+fRy2ZPpjSQKaMEWVQmD64EUdWkb1rELkJV71+UzH8aqmdgM/OnVraEgWE+1Vg5v5R
EE4Bo+C0Ej1RNIUcTQ/s6KCZpvrNdFg77Dw79Y/l/WVypYKXXnmezyAqsx1/VadczkNLSRxuEBUa
wjbRcwjcccFJ9jPd9kt+DAJcr9ovCyFYoApZtEAhZZ6opGPwuHOsVGcAtdStelWKvA5gIjJ4oqBa
ZuGnDIJBGR9tTvweK1ktH+v+9OVVvGT4fL+RR3Jh2286yPMI9xTanLAfKv/kgLWbSvrO03AR7h5m
vwtT34CqagZWfpmDAPlF9HR3m7XCy2hBSlhJm2Kzz/K6NuSWEV81y1wvimxmxpbtF8kuuP0rOt++
WeJpJGV+aS2ZR88vdR7OgQizjIEtMzHDCEBuRxTJmQ2ULqbX1X3XIGZwDbdQSS9eHd2d7bTQ38eZ
+fPwIpd3chTmjEDuKO3ucoEwtMrUHGTorJ7RK6ocxRhnm3qCvdJqvnzJe3I8rui7PYWoPLXuJ1Rc
aIeyOIC3TTVJDOoD9QUs520n+JZjh5rMgu5UVub4kUQxhkzzt9nkL+xUQOW77ETkZHbhjt1+MME2
pPXlsV8qMEsnUYl0eCaEh58sHJ+PcheYnpNVULJbeL1RfiIyMXoHhDAoe4Bo0aDyNDiBXS6g/x27
rVgavTPYeTGyJIdElALa4ugD2hM9Xt3ZiTYeRm9pGxa3E7MdO1C964zVJFT9QrIjE8trc/aZoj5u
tHPbxl2YWxNY9Sble1axd/8Dcv50njYc42LdAc161V+Ffvz7iwto4quLP2wEQtHn2JsIKWaSbOeF
ELR5HBcYtnHKkcRsJhDbCDgbf/yQQUFbc+swCrh4Z0upNnnObokC1DKMpty6xNMlXfwuSDGy1Nak
CeBdMwske77Qci7v74hDqPsJcODKw+o3YhGJ7mtwYk3uSJTksXQqf04Di2rwfVvCEIdY8l53scaq
GV/vbCIYdtIQQsrQUzqyy9oOlV1ElbYhMGMNrUToqIbD9cnBePdsFKQUnCk/YUsHIOdapC1gz4cT
+TSa0uyt09LtXxP12hBZhy6+0sX8qp9g+kp2JFKPWMAyUt1zSxl0TGDmsE8PR7IxbLeaCf2d2hdv
KPEGnyeAEIqNIAsDv3vbq2PJLoXNJQWR819lV//Qs+zpmdoJYW4STuhDy7qymMuIiKb8bCfwGpfD
DsVMlL2akl1P/poul02Eam1j9HkA3Ross7NmU7OE8ne4x+eHiPYq0Hh/D4tjr1kQL5jd8B4qer5P
0dbK56t5OWW41mTRj3PUmiT2dzGeQ/kF2xUGTPnv4vWisBdwrHc49ZNWFYIKr2FjejXOdGvgtAVp
fBeaZK+pfuJ4GxCH9GM8Q06x41wWWQQCoMU46M9Hi3X+wiJIK5ozAAnI6NqD3eKyY6Q+ytfpfwcU
D3Bq5KbW05lFROooEogL3x0UWfgjRFOqoZ6c1YmWWONp0mY/ciEF0/xQzd8BnEU0Qv5AhEcVk1na
6Sh5K/P/9vFmjNMc2EZaRvJN+tt4NhuBKLOy7kXbjaucy64GTZW18DODpg8pZtEf/5Q5cEGLsxYs
vUyP/x5cNU/xrqYGTjmO9F41wRTfk+lMcW/Weba6YHUKXS7/Wq8r9c/qstx8mPFtKYGG3myTrUOb
pMGSU5Fb1OS1Tvzfvnu7IAGpqbyRD+kJXARdJo21XAhCgnBVblfJivxAjcBAYp7F+CB9fLMbF8Ho
Nu04hzM771T6285GrdyNyidMkmgzj8oe3Z32xzdASI4DBF8rbYrZkTq64lnzNmz0tJiqFAE6LsZr
6P3JaKLhoHs+SajkQ0N1/99AgvN02fTayivFfIq3+AuN9R4NSLt14CnndMT7u1UyRl0n0gqS3ROo
zPXRMmbQDiyIWTyyPFGXMo52JL8X1Um2Ztgh+qADMPYNJwyBMDWHmqLyqzY7FIM18HDlHciYhxFt
eBHK7870JNjFpYrI5tAy0GHl/dZog9pOPjwJ8lHldjRS2cdbW9uYyJAsu8+gDGerHPX2lPmaiupK
M59HfvjnSbTr/vqxN5csSg/+y4Y9Ne3HLeR8olknh8cE9QQLRFuatPJmtA8Ep4FZgjtEoyVRBNfp
P9nzWNFRuSR43CcYlBD7Zb52W8tUmQEAgCqdgGymkJcyUxH7cp6KJOjfFXW6cIVULu3E7JRXqskj
fcIK0mYQFHh5gD9ciaWtNtdTNb3A1dpLy+i6eH+0n7AmJIVugZs6bK0Ho7wS61s9c0mKMcIml1Oj
3P6bMaz3GpZEKM8a3QRa7+m4IRJYlPa1RaWKiDVR3s7O46V9J0mXUet6qEeKFZZSghUAkXFpeWJd
5pl0Ith6tuu2selNWwi4bq8TwbWq7DR/ZASxQnhMBnjrSaJlnuuR/H1ycXczMll+IqHBozMsE9XQ
q58CQaltLJWYQ5l7bGL/DmL3KAGpI2gE1JI3g+tAAd4DFy0NaY0Tpgf/zyICHD61Vc9RVCGBpZnQ
ud072fIhlTehV8BA/SN6lmoa42pmri8AWW2mHT/jxgN2XJ/ut1ggzX07+w+64z5iDtqk08a1WWPy
KS76/2H72BnfNerOEFRBT1tikw2wUo5eKz+ZcfoZy44ifP+LdFt8spI+mLtwqTiiW+5D/OlxKi7R
PSvqt6Q0D1zyRkvv6RN7mtuLifoqYqjKflktLNqMoGZ0HXxKQCQHpJlBpkhFpCLrZLdMBOAsAjXg
2LzEwLurwOr4bPOzf347YTQtE/f128mJnRbRG9XUhMRbCqZjxk4hVCLhE79YbSDx+TXfMKcN/9K0
e4NFH/IBxgLVwXfkcbICAppXWwqTyVxGjGXTxEOt1dQdAz1+8ZujChqnM2xjE5u9HrXXJwS3wudK
aTmdO+xo1vBgJdBj2bpIfPIYIiIP5qYXhil8EjMz4Lca5a0D9veCgzRCO4ZUHeY2cWCnHjy2ErUT
SL6nzTuNs0uPvXqYwxQujNj6ACM2hQokOIT743VwRunM5tttf3TTYnlej6SlirsQL1XOxtFeje7r
3NNyS6yfvguKCmEYiJ/20zVEHfSdfdOJxZwf8vNyjceJpOsuR2VoeNDhor/sxKnf9baGUEb/1eLI
ikddiJ4ekUNjUwty+f/LM4AfkdDLDkMqb96X0dEf4Qc8ZN/TJ7hhYSo/d6BeFMH464s+tAqtKGJM
8iBxpdh8vt5xzjEUlAE7bXjwIu29kfwFaAaxJFR3a0HhUNiW20KEb7N41sZRzq14f1elqva2gzoD
xt3G2GROFlcURbOc9n9/iNlEEz+NCZhDzuEoWepRnHh0IaitKEvaAoYbKOAjd3wxIj5alhxWSkk1
5Mx4J4PpV1ZQ/0R/4Wplb7KkZJqw0Lccukobj93j9Dvj6PcQfBTIo29Mj40RqjAa15rEaLphVZxt
TQ+nrEN8N1bomXGOv3PI8Jd3lbUDT/tyyQJsVXPa4ddqD1RKsHd5KDafYxuXd+cpn4Vvnk55uuau
E+XcDrDbtduXFLMKcB7Z8l1HbWn82rZF3JYBxHPaqUJTyxRTWBNHP8MzqfnzNr94zG0a6SbxLbEQ
aayfJUo8+hQWckjhvAJepdGwLP594eJ1DKuPUqotZgZl180l4ve1GOgUBy7brx18VF1ChGB/qySa
xLdcXwxi/pKCKoXUyam7Rfqez30eLXFZ20bkapbrxQ+ds4rKZvS2WDuLMuPJw63KLvQ476tUlkvP
+gxhsJPXqfnrfoo/P8EDyNjPVDyaLJbGQLMh4Wxjv7vVv1KQAaqkzr+1QDKCv3FU4q+/1yErTzAH
99ZDrhu8HutXAY36GF7KMN3GX2SCFzgC1toRDoNs8T++RHeDk50u2i7AbtHELJSs9Yad7DPU2/H0
UDgCDR+/y2elyLbXWzytFf0EHGk1XJwBKkFdoCku9OxQy7ElaJvQK/zoS8x2wf4TMRgh3ciVCXRk
CYQUlBYZGEw5aJwWmOvBpYMFp8YKLMh1rpS17KJRTPc6Ry7gr+2uyF4+/2+iGM/iwCXyZ5nAxZ4A
rf+40dYNqp7ArrUY4/e2N8WGD4plPCxteQjE2xV0Fxc7VdasDaHJzewPYrBrzd4sBnpr8hbQv4bx
Ag4AIbU/eTKKtDSi9qpRPA/2MXlGEIxsKbLGraOBNeYa7y19Ycw3Ix/eSRJ9D9fJeZnFc2nOHRLF
aZtOAHFCZ/gDF2qF+6M/+w5VqngEo40EvCu+vKNCkvzwWwcxjewYVvCRnrGXULcGvjRnzPtKsd/h
abBhnaQ8IaQvH6HSq3hpQbsg/7Iz8jI8Ta3RO6GoJj1S3lhZfp5+Fqj9eVFHJ1wGcM7vdIhNfDU3
R+B+mpbGrH5t0nNlqora1kRLNUWcx9BsCTt9c8VG4V3wHPpC28Isn9TWo6ep3fVNYH+RSS91cCUB
xVIIeGGiAtzurYUBQgrspzz3QOAqXeUW4TbFV5DHZ8C9sq0v2W+gseYCnR61vmxo0MPXbWQywbCX
Vo2XoWuER4JAlrlvf864oEoKINUoQlBoD34TYh2l6gYDHj5lCt6siBiTxPyMoLJzLlFdRUsZquqe
hxb8G5gPFcnV71vhXGJ8ov0zXvbdDGCR3Kcv8/MFU1OER6WdDIQmJzUtSFkAYwUtdCITz4fO8591
+8sNaDQYfgmOe5tOjURjsW4z2U2ic0VCvwxgz93WRvz5jxhR3E8DsTpW/21B0eWorEBZWpkS2xzi
pqlJE+VhzaxdvKbKSbPnur8l5RKufOXZF96CLOp7aPPgh+D+3nbYVnkPQX4rtXLh583wr5jm2+1R
UlLwdi6qI8P1nyDbqQYCKZIhKWTD+L4KGdRlPjg57XRIO13rC6urafrhDnH6AOG/W9mb8K4i4KK+
baI71GDMvAsD79iC9FLDLQTYy1TlWyyl2rKOFnkevxSYgLk1JV8XxrHXcrrRNqn6cju5QQc7oh/0
QsntWFUUb3G6vp4b9ieqFYJ4+/ja+PVygZA6GNaP7jdU3+3PuwwZ/mlyVtWCHsYieYHW3NVI+JNa
rSl8iJEF1dpInqKHnZSBpXjTB2sZX0adlAHSS1FkzvIAqx7UK0U/Vllu0qAF/LU+ZEZD+IcHId+4
4+jZVrXcrBi0QhoWmVs6ZIAhYkCvnfeKgUR5OdIjuzR5n7wO7cv+KiBaXh2yQxhMgKcYt1FVsKWo
0zYiusIQislykAP+/HDeaZXsyhdRuiK+XGBgWQVGp+OQm6pgIVRuS343ybcATw2bv1XRa4PRVzjh
ROa81Mgd9rKbYPdCu6dt6P+BLFXTL7hirCXbvwhywRgif7G2gSa8/YsPYGK1E90+q3V0sXARVASn
JP6VtxoSNQT8n2S/AYdup+JJ3RrJCLcMrWFRNI6q71OTk//b6Fii6Y8lIAJf0wNDbsXpqEIC3D10
u2BTtm3N3o/IZmrF8kGVSpwB0zdXQYoBJ3fSMRFsju8p0Y0PG9JhaACI3X32Pnh5O4R3l0Ez+9/s
S+njvcTtTjoZKGx5SIcykhCTnTXXL79iM2CI0Z/X35XHsrL6hr3O0CR4Y+ICcGnSeRfY9FJ9lrS6
8no07yZng7qBhIgq6h78YyJEiiahRKheWrDflA8dEAgU862kdl1OZ5VNvwee54f35XtxmmWc8ygY
XxcA/pyHjecwUt6O+iKj3imgF7LjrlWIeyGJO5ET3vk0zE6bnrnMZe7akYqEKQvJFbRi0/acQDBd
BrLS506ytvoEtxC9rZ+VneBbX/6E1+WgDykmNp/FalI7t9eaWRPwN2p79IezkvfcwuAAOkP4MJOQ
sLqqPmrUvnX8pPYcX7RoME5oAT1UeVdkhF6ZHEon1XgUnsYiXJyBPx+f7doCtrrjdBo437osn+fe
uRROvIn5bQwE5IosJ5IJdnVdAysPuyY3MAkquqBgvTItN9iCWj2zzi0R/Qefq9crYMo4PrgLv8Sa
71yPkNKmejJy3terbnn1Qy9NBE+8btJp4U4kooDnrTKvsGfwiPp8KFZ4YDBuR1SDxWj8kui9We2d
PDAYbzVivsBKwIAcI2WVuVFKS9xvig0nHGRZNzy1eEpp/ME8O/ot0MaOk3tVFyZxN4TXtQEilvON
aWksqrAplxQNHo6B0IKEo+gjpYDEwLRB3V0hst5oO5qZDR8dG6gLP3Fqra+rSnswmQJwbR8mgLx6
8mgcIC6JVSfLVs/SLMNrvm6dkUbCPZ9xg2iFa/YlYTeIA0swWcnZgJOgg23duphzNiox43E2hC2j
Aifvm0mxyGIWZScCJqC+3R5BVgv8b7OCahoL+ybh/CpsF9qPA8VRRoz9/1s0hVgoC9jV68NfJnYZ
pwcgFx6vVcHx3l6LbM0VsJH7jysIfk5FDrl0Lwyr2Yun7nB3Z3lgpcW67yTQjOshHO2DeplYB8hf
YaIo0K2/m27ZZDhNU428aLxj4NHFnzym4Ew09qJGTM2b4+c2h10Lhllg5UJLmVhSzHXj07xKAg1m
WBZjPnwgf7d6FlEvBzgufxnT2GpJ9U21QrCRYzDxbQhDvX82lPNoMSWGsoN0WE8VsSypwtPL0tRR
dfkV0R9gfresLH/bL+o22Mk2gE0dv6DV9KosAmD/bGKuHWJ8Eg8L53n0WK0Zqv1555farD19FbB3
v4xebwE5fjFI4S7TImUdSouxnF76uFIPprB7qnXjb5XLIdTu+3Y6ikC86wHDEoUl33B3kiwCO6zD
XuMpA96K2YGPdiZyp30fNnt3C4mQi5IXdzoNG4FTel1flHEucLKELpnYosw8mMTQ8OlYrft/kZZc
JNM356AxKp7jKHtbCPtPObPT5npf5nE726pCjFND/DW972C0wQdHbAsTEe3+AK7ZnpQ0PGLt9zHK
v73QATjAYA2AlhUXpdquTS/M1BgTKCzxlZxbUjzDyIy3ZzUNRziKfanNfTOC90EYb19gjbDbL70s
5UAFY4kAx0zHrosr0TMiZoiAFlPSkpxF3gdmPSkQKpmxctiJGVLdYdUFLUPT1+Odrt9KMVujaqko
blYijJ/x1sBKV4swKXoElmXDIlGkInnaQzb0NpUvKFibNeKlD8DPYPui81OLUIMay7d8EOQVb2XG
ID6YbKTWC1v3ydyBBgxEsGJwQCeckmuavIfMRR83SlHvmknVfUY+W+bm99iW54Mofq2XpJ1iLLpw
XQzREECuHlgO0TCt0GHVirNJDcJUqIRRjuksj1Si1M0R/apmMyfqKfrZz6AaUwv2fa3l9+N3KNK5
SVJaodDkSTMIF4Flm7W46rDMxA44OUTUP22cH/nSh9mfYE4fIF/Tt2oO8hq03taohxdtpo+IJPG1
/eYhwMoRXbQxRRPWg/Fg9aawfDdlZ/+iHMZWF8UEziQbkG+VRatOltzoZLj6deaxcYNC/4pbCZSE
q7e7LgCZYeyEF/nNm9KLVywbJMhUR0sheAwnGWrgYApbFSHGo6cI2lRfkZHGnsm2HGBodbS7x/zs
W9BGUL2OyaY1F2gwrX57WytaSgy7T9C+12Exc9o3G9/6p2b1XYcTvdOAyGWg49pIdSnxfgWjrFPs
i/5TjMMozjT2cRvw+L32fP5sv0FrqqkBA+lFRXSN/K698w6j2Ow2FR47PFEKPfLlVNejui4Eva2b
/1nXVyFwFNKw9DVDltyuhMMPjYr3JSw9El8o28XIDUyghUxvWNgO8LM0NZsNDS1qGRGeXqs/m1Ez
g3jQjjJuinxz0Zyp5ZXAIcMMrKY4gObtoAaLNekzcn7guQsWsWVUh3HXHoa6VyPsb2ni3DS0nHBw
5d+PDVY4qr5rqQtU3JyNj/si45gbA/SdKwiHo+DeF10dTgVa3+zlLLkDYJywncN3tw2mK5mac1bK
f+MUEiKLOn3WZtMgk41TJ8D+XeLbdtCmyVPWC1iPv4Kh3d2Nj88y6oPpR186U5/nUHsTRAZOWFha
SG5ppHVQ4/0Yxe/4/XXXFKaSe8+/e/fZHtS7v2DvpSemDbVqL1GQ/TOYfi9wFhu9xN64eclnXY8I
A5uQWUgcxFOgZ/4Vo1rmdUhBbaZ6XWc1EIUKjRlDF3MocY9PlutcGibgqXv5DHZFYk9XCbCEcEj8
EUTGILAF1QT/gkr/1o3IZuskPghcAe/D6Oj8ogL7OTV3YvmA2Kz0rT2CEjwJ4mqtCWRYgG9SrOvg
T2oKwZESWoSydtYaivtlViDsmbqXbG5pPQ+cb3qkrW3o/PBfjSsDv1ibtu0DTKfH9W7tb+9A2z9p
qYjkeUEjcYHKXtwnNk8fhI5xBtAqaM8p7ZlzInKdVVgFg4nRdP5efWEJ/d8KO23T9GzxGF9lc7to
olH1AC3QB+f6apzmR1fCCqHjJ41F+Zn4NM4tLFr7pmY6h89p0QWqNDzc1pZ1vxFMLNmANRT6ZxDD
cdBbB83OEuTskgHOe+DMcwxJV+ouvt5I4gZWAJ9WAFfM71NQ32C+bdxpZzN03jlUJm6fPrD8ETfU
vn4+HFh8bSc5TuIUlc5FEldiZc/wQjaJJlInFdpOWYnQabvcCGtSbXmtH8ZUx6u4o0ukHxMb/Onf
KSNhPtRszNzQPMPO2o1zDxZc/e4fvRdSxX0h6PEQqB+hgKyHEwDgunEZTRSCsZCVH3sh2dpXIVnv
Rigi1VMD9Bb7LkqzuZHGACXDegYCJ30I8sa04ux6q0ybGXmy0+FkAJgQiFqPpdE2kxjMYp9ThBrb
ZuvT7EL2NLU31n2tyxgbT9+Y44pdgGfCx8NI68nrgS+Oxaci7W9qn1d7WPuv28cqhM9VeryjXCAv
LR16u4W02RwK0I4c3ne9+KPTgQrjce7fD/KZpEq7rcbKiyNHLat8RVPjEdiu/XuMuwI8SAhZTiQS
Q5Ldc4wwjSrb0S97jh1T9+Iws3yItUyHn5EiGCeUXSFJOaYWqLPTlU5VQoSCw7Umwoz/rZyAtcGC
FU7OUBGAXRhRolKcJ3JfhVUm1O4iElqA6JPl+YoMjLnTvjPqYlleArvwdbKbK5wN9xE3sc7Um55N
kcJhUI3rLSzHQFlTlRxDhenxdg3M7+pJwPlA+YEQMZIALnSu2XPeQPuw7n+andukTia6TFZogdd/
ngHR/IcpWKMAczhfQoqqpAaQvTwJQCRgcGWQtypO+AP9m32dJJPK37ayKmzC6Kr+A3i43y1rJp/q
QcKqi2ohwYkvsF+eLijm0M2xczHRS+aSE2LaHPXDwRGXWkctvaDRZ1AmxRnfZXBGSViI3gK8a9ky
VBVZOAC8RxKvSyq3Iv2ce9YILzK5rDV4yn9HhgFjY1kjbBN2FuHIgE71OvlGQmckXUTkaZonOoXc
kX409RVtK399V2Fk5OZwTwpEOXYU7dqHg5Z7PQ12YA/2P8wlQs5VjfSOi/oLwwgC7F8uWQGGTf3B
bnotdEO+iaQFA9gHvFld3Ihdpga64tGmKcJmqxwvNzsAZKd/NV8vHO3K8dMWVA9Q6JI4fuZcwmcz
+QqLA8sxyyTcP4NMG2rVeufBXXj2NsjPny19j+y9fxh4hDxn59Z5cvb8MqQ1nqwwY5ZiTyanKKd0
s+4Dyw2hkx+0a7qtZOspC6sjUc/BObUmrIyK6uDtl5pllVDSDHKGaBkIjN1gBR+lipRe4FzMTPbn
DbYIhUMGHBdQ5T0/yhxNvvp24dY5E3D2im/3zrtacbaHS24b80eABiYjrXlqUUeB6HuhEgefKaRG
xlwnMtJlYR55ZKZUVEJyov7s0Sbny4z9jieem3YSfXF7v49prmzqnzwnn5C4k30/xKa1nP7O6JC0
Zk/TIHd8E2J9nrWW5uw2QrTuUttfnPsGqBy2Vq0gxeEN/qVZ6CglvvUqfpWN1HMPli3AI0HnZUYi
Cyi7r0KYd2NsNJcmz3qaNj0qjHAjJZtvE67U24EZCofW0XMSVpxBJ9mbR8inqCeV1xp1NPzVOyrF
YvNPDYlQhNWxz3nTDoI07h6/i7m/FPMUbtyRb196w3ttQqAnytPXzbdDbHXpCYL7CIvbWO31Xz+U
tFGFu31wmtdEag+XZsGkhy9bT7kf/xQ+buFKGITMvQH1I9GYK16EJfQaFF1XracX+HTWZSn3tSY2
2l7JrMzF9Zhjrj57nhVZ836DWz94VYmbUUEgi9AeMDZB7IezIBUCfWYut0Z398TKSWbFpi6VvA68
dgF4gdpKxE5toztNns0SA13U86Zj/I4MQtmcnva3gxwmIupZDi24B6CMsajqsqaMzfXzVCNE0Kgp
q1AIp7eh5TNZhygXXGPHsBWBAETBfw3vT9iHfJjQTn/CBiFyaWk/HoOW6rEKe6oTgJyca9OR7Dp7
kBDR02mAYnov8nGpotJG+/FuyYbmB0W9TSMPJed9ys6j5UiZ37DrWPhucHffNryBiZ/L+++Gmdyh
ARENMzc2pU+zNgEy9E4cAL6rB7dQErmubtcjnCVccXYAP7n+S0cpwC0t5eG2c8sokaS62uQsShWe
jvMG6skuQBfvK6tWsjlHWjzrML3WX1ZTxl4yA7oJkI4zg/qmPnn6jRxj1E+0p4pE8nLsN+Ipkkge
60BmonvJX8cXqQtUY9EYD1vNPtEypNx8d5rs5YLuygICDmGa+fQZgeI6g3mor8Q0uER4lhidjSDV
c6e8f63ggwWmbm7RTm53Q2gVW8YWouhgPeJgpVKf7Ij1FKRbSMtc60+rWNoUjninv/G00cVGhLDR
KyUmeUBpi1UTDgHObFX0XLD3bSCpq61kxX2k3AUng0qhDq/RTxQ8X6yHjlsrL/r1xxTrM0ZB43xy
V2YWinKn1vDX479wifTil6UblwFS1SD3SAeuq6YaWwelB5cyF37p01Jhfrc844J+MFAV6zPvoBkN
itiPQYdd1pIJiNytpVly6fw8qxHPw/5AUwOCApq7R/ogqNBwYtQZvDMdqCMvv//MfknMJiKKMcKT
gW0+MEPQ1QBEH2ncGg1NMpft5ACQY8/l8evgymYXixvgOYYBwnIMLTbOU8TIcj9F/c+/izSqZ5ZA
2u647DfvVzcZmoz+EbsfdQX49P7DQMT4oxfEKdI0rImV6aXim8k3cn/iA3rIR+IH9zNkY06Tzy/a
ELcV94EfwndE4LQiyNT8fkAl0g/GTtrlpzfoC5QB1UyVoWTVg9Hb7Ld8RFs3cMsvgj+wWgctg4yv
IDVcWe4N3LgNu6nE16aLDkEnMT0puzFM+Q/f8hJmmewbwfz6SSFuVD3UPI3hjOL8/OvjrOGes3L7
bI5XPDd3qH3D1Up57/SMTQTMB+qlKJtrRj1guL2wKGkRqL8cdsDUP8k/48GhJNxif4XxWXrRDofc
D5JO49vCqt/DpL4I1EfSLqmbD8dyrQ5IpXzbXeYBfc0FK39kwdkzzPpqhJG7RMlPKEBUkP8wfFoi
f+BGHGCJpDCMfn6AQpghyMWh6KwLvEJJgSjhmfKdURSemrYJoAT43bTe3Rc+M9dqBb640b/BM6CX
0l+YWDLkoellRo4s4WuUR7tIB/WH8GSuFYJ+1+PmSc9ok2iRg5lRU5NJ/Emc65OHX5Idoo0L7T81
O3MNz00y56HvutP8W/GQgLm2SS+oSxWLWPpOK7lD4Y5/miUbi119zgstyZJfW/0IJTD21q8fYIfM
eTYLH6NuOgpM3DP4iL5ThEJSYdjU5jLYfDrRdXUvdd07/XTA7W7F920KdsmI3uWNIzo3sK5imHAH
FhDrQYfI4wNCUioYyfPFbquM2INaIjGTeQDaf8zSPdCEZ4NWdKgITSG2Z6YJ6dXz8xGCHglldyLw
cjCdYTWjrmwl3p7ELfE7pC6zwzt/946lNObr7dv5xILPPJgWYKm5OkbQo67RLACUQwAPFNa8KPAK
+099YAiURkVrlgeiZQZMDWMLoF1UvgexH9nC+X97ZljvsZi4GtcUQI2oHP0Jx9FavF6/dIGCYxcR
aviQnlews89rWPEr/VTrOFIR3HLufXjnxai1p7zYI22FoRzIMpKk+DOrFqhyv+8YDdYHeLcU6qMS
dUtQKpMUXDGtwPVaoJ5cAy+t3f3L/L8PN7xGfMYGvzNsHoCRkw7FwqwDSybPDwx63VBVLPEhY+3y
IorZuZxISP3O+1hsBw7FcVp7E+M6IW87F2EZrRnSY+QiiZ7B4U9EB5hMhjKlE8xAtgcZzVwqv0Oe
xjT1GJN0qmirZgM863syXBB16kr3X8ITzYErsv+v7lPjB1CM2S5dcJMVGSQaH5CS+JfToeyRSE3W
66YK6qoCwIBKaYZGqM5PaqF/lKs0bHBDImTc9ZyHvxbM85i+6YnT5uCMDvtYVnHqX1PrmLTM2D5C
swUzie3Kulqlt/lzkG9bDKEawTfrq10ecJQx5CZ9XdGSK7+kMxgU0sdDNeoBwh4ZihtRIJ5J/7vQ
PcAybjlhl8jhLm5zA8rlmmCe0CaNWxiz14M2GH3e3oaqP+OXuGHH5MeONhHjPQryjU758Hi0cDDL
If3JhRvOMw35yVKiNaVzZwX0sEyhSWcKtdzXxfpDGoxCliK3ZDOjDh2eYfJSUhHPFOZ9SPyVZnzi
BXeZQM8HBmu+HTP01o8u4XJ0OtPTt++zXEnREQoNez5mRDx7yimLiUKdbzmsP0sWUJ2L2gE3ss7T
iRhKHylkP7PwlNTmP5ol4vUAqJKqAXcqzYS6+sykaN/qPddu/JWekoOfC07hsq4BD2n4msJdGdjr
jGU9UqaVhkdDWD4TlD8naqhHSn7Vdo2r/yEEE9hGOsBm+uP8hs0DhdiXEeMnkc2zQo+LwO11Cj6v
LXrTVurIsBYjMIuOpjJaP12/FODb0BSdG3fxXSin2Al3GOKaMxke312YHE0KIt5zWZueJHhg4XVB
5ZzTKcA9HFI0jxGbCQ+5arvd/V4fqLXZ0ke08jEnKVcBoC0hXWPsEMTWyk6lrCo22VqFmulfLGYD
/aVXPVJpAW7xC9MoDSrQDQ9Csc3cnbOjHYpRsLMtgjlkswtymf+vlwMYT3dj8zSrWMA3DpCJTZSA
1Gt5AVZhfXY5iybJq3wYhUFJC45WYo76aAsekYlEeUpjy/t1ycvbKwEumA4CTcLISqVSiNSKL4EY
MwY8hJrf97Mb0MgTI3yrFu5WFYO6RbMr7J2/MqZBrnF9LJTe+swKONCLzcDIvIW+US3LKJ31H4yd
gITCbBS2p0wM39GxfrCma1laqm4kVUb5BCoUWx7WuqmtEEjE5TpvTdTw7evEa+J3uTRJZ/VPfzxV
uxXh2ToOE3F1AcC3SSkzoddlfkjpmmUcWmb+HW1ZD58gmSHrJhStG9shv6dQxGPp+khzIH0VwCvU
I1BcrWIfyxK9Ti/mXj6RPiq7h2hqqnIgjG/RJ5yHodSXdnQstO8EjxypFk2t0bIN9NrfZZHBiwy+
FrpIZkE3PGGI0C2HjjsQD/EBcoSjLvvWLWvnHoVnKNeL+XLJHJcDcDnBE4JE9uIz/wypqsvQdw7X
qwC6hAdqZK+X30gqbfCtSc4AqWMSPlT4/QOJd55ngryhLBQcmgF4rZpyaxfsA0zjZ+Sw5tqB/dCW
0NiJG9uslufDUjK9J2RLZPkt4fky7LLJhmM8mHSNMjNXrJQ8Zr7oIsEXsTP8Tg95Xl3txwHNtowl
qzQNjEaYIYP4oRpZI47pFwm2z65uvpk+uLhi/LcpUAduECjATqKswd2LqR0YqaUJLwDliJ20YxLX
m1GSDjck4Jy3Nmo2fGv+All19pCyulheqYFd/6hsg1tvlejEMdCQ7BtkbEJfiaSEamhYtnbhulcb
zbv+yWs6ikEg9CnfE5SR6phFOehUQDZkFHTrZPSNYd9I0E5czpPq7tFJ55v9YjsvJYf1fyuji7yM
pMORBzV/69Qs8q9wjNl5FUbvMP9guFpX/NhSDvYWuWlehslrJpuXmJJW/lSDKUn6WIUkqNGnBA7N
UkyledtsWXIKDcqEPu3/cBT5nTIPNmb8z/lVl7XrWrdk+mHuvpi4Npw3HFPjUde5w0BTS2bP6bRE
J+ZNeDVtxsE3/gkFLGL2OEnuTrQKuQB0mIxBe2M5K0OJoW4bWqb1vlqGxZ9phIh9Xg4GSrJoeg+I
ic+Yy41eTHEEk5dpZQXkIqbtywP8ebiWPzzlIiJ6Nc4hwuF481Sn1Dax2342tAYrixd9eXXMIjyZ
2e0ZeH8+bNUvxxCHNpeDynCB16fWoHALkgKE1yE0NgLe20kto23N8wFv1sgEZfG+l0utm7hqM+6u
tYMuvx7k9oWXOrpCGa9uDvt55Pprf/woP9RDNX6s77ubm6VWcuUO6d+pRxpoCw/JObqzXV0nYP01
koiUcbvdKz0RrJ6j5kv9r0ColD3uzGIMD7Gpv9VC3jRqrfD7TaGmzhHSHaTarwRNkW7kN2iQ9NzG
LSQzUyw4qgvUskPvxkaSE+yNCa3WnTD3VryKnqvo1u5gLJTZF2pSymGSF/heIs1IICf8HiO4A042
dfUyDx3V7JuckMvIw7ch7VQXweUhnW9CKU/LFhsxPMNdhfDvff7R//8cqxqw22L6wSy+7uxcX6w8
hByCbl51SFK4hf/m9mk61UDi4rx9jxqlYXf8dJ/uJXzX5TDWNEc8eDGdAoZPgfgu1QDHidKvULNZ
ozu/Y7cSkq5wTH1BRcJdbyKwAUcPsI1hX41gnQzVxksBztfqUL/kTLv4dLOP39A8GigH7h3Vd0KH
CrQkX7XUHP0FVDM5hPffL/lHsVgzVo28M9O+IIR70E2LkG91nJ9a3Udm6AXoN6R8ABzuW4jDKBuy
paeGI7GYPCMIyOyt0nlKBswAMM51BNtZSVxuBCA2sXWOYCuhI8de6GEgnEHPulGzryvBG6ebpti0
SU2OWXM772bJMYeP0swFU6FbDffWvVH/nyQxKMAEe2TlU5Q7AqeQyr2UjvyWTDogR4Bmg2096AvY
A5llKpkmDpjlf8g7h0AZ0c733lhgTwgry/nUEek2vf+KIujZyoapObSKyCBUh2V9Cbxw5CDi0Gvp
IqYTQEyBJe9vhBFbvNx6nlBFR/LlStS81r6WDTfV4tDf58efKBdMte3Ri4PO09I459JpLfinN4g3
xHcsU/4XE7rSFk6XknrPNDd/wux5CNSZO6g3JBqU0606k+zxxMAHEkZg+w3GlscJUIDpcaHbbSMI
wFeG//xKHnxVuwnvJx00SqutJHiSUSN+MGrbnLxOeQrntIQ9ub/5fnJ5Jf4D8a8Ln70c30QBI75O
93tXbHw1JBz1z5hhtEOpPbaK6FrUWex0LJ2uhs2d0tHmFm9J2L3J0XYMiQVE8McjQZTMdmqnJeqq
FDPr4mBSRh4c7ENq6KbSkbLgw3BiSn52DNneNiiA/01Zza4O4MV04/o2hKAnyp7kHr6QrZ5S8ZLo
sgEHHVE6t7yOLeK9ZD0kderLCwwpa9QB8p9qGwAjUyMl5IoGxK1ARBTpCmHHmpzhp6yrHb4Jb/Gm
gCIxGgmP8iz3WsLD0z9na2d1A/Kux1+CH4iBMFDJaT/0fbqJ5hH7AO3/laEmmyY6peKw5uGi81Nc
WJMVczFHAo31A7IZfsG42nimo3gmS76YeeI0GOVsU53ASmqUcHw13T08Sd4/d4KH4IR/QgPzbX2c
pejrQt5VNMz1EXKvfXYEH3h6bHZ8oo8O9j4bAJWtovlCCjzSjB68hlSn0Z84GoA5cncLAsSIY3Ch
hVZTA/dVM4K3Yuxu9KVcq+W3A8CMt2u1wOLQS+C3Skq3Erl8Vcn56jyGxFf151W8D5Rpg29RZ1UJ
rbpvwXzfSLsDSvga57N32+vY1nFpLpaiiWmLZFWWHStVhr6EqQFNXuC30JLW0O9oMg6q93FiLjGv
Ch/klGMftk0UC/O55nnA83FUGU48IdZH2hYBYmeKdmOfw969JVOztwTqnJJMDsueVHgwLgE4RDZZ
zZqL3SYtRnlJ2jJeL28iBLlkufb22L307kysJSzEA2VzVXeU1i+s6TCpCWg9ZyUy+TKV7g6LGvNd
0lpmIGd5u9M9WSeJv+H3jnKfjuH8WSVvkBbZcSVmlR2BXgOYJwYD/t1Oasm9ndyd7YjsSblf9HPn
FeRlirooVKluCnqH0mVdgLC6Pi5ufa5sOa75qAaSyxyEcjmWbw+d1/gMlziBgIoPyznZUsvLnsxh
faWL1hJYgnmg+nbftvXz+lp+GnsFZpJKq6Fq2qo/AO7jpSQzxJ+rDUROgi8PfgNtEwTl+DCg9wfm
5OGjeQi5caXJ6UOFBCC7L2/SqITi0UdC4VkIH2y4EDEfB9sHNWKxki7fGUncPXhTFqLdMmWL02cP
nR1EzBxxmQffdv4SeZUeUEglG5jrXzvQS2NXk+rKrBdglAg8SuddVis+E7vqG2gbDKZHar2BqQQz
65uEuDjBm0nl9ZSH9awDA++SmDxeDV5rvzr1xfPiGO2BZs4leXlK2DqYrvx4EjNl26EwEO1LcfV0
DTfjmmQRq/AoleTaP9WJExU4UTbPsus/Hdh/41onICWmXxIlpcBi4zy6M3rKrXZJRyEmUzQb9qKa
euaLVA9FnqKsXNkgJOrKkXx9lAJMmFxUlwCnpHjDlqDh9p5AjUJ4Ct7nBpFiuwNVYXAUTPqcnZx9
dtn1sInhFjhN4nzKKNxtylFueKsEr8pv4CAuJ6B/kP4exn6Dib5WtNmfzU5RB20r+Ltw1/U2vx2X
q0dtpIwHuFUoj+5+8vmwEC+W3S6GHgF3Olo5LQBh/llyRN1HRVuSSdmj6AvcwJa6eQQxwuxJ2w4E
w1ltntYMpCZt5Kq9Y4msu3j0ugoRJ8Es9cUTYWGvP73+mIpfJmPlnhEibFHtIstqw7Fp7VoOkO4z
ET/qOKoiddZ7v6VLa//OEYvgaxEcgYhM2KOAOGGfJo44ELuctjkLwqzyopgT/WbPVFjESCYmF3ld
jkF/6g3Lj9seQJkX8DXN+xmWXFUYT7Ef6R50kWGSq++9lohYZ0lzDY2+YaeDQ/DroueeGleJ/9yy
DbCzFBPWk+JqbwZK/coym3aAFxpcuSEsLhhwVTnwvK55Z5O69byU5N1UznqXvw/5qe76/dxo3VuZ
XWIETVrxDNvEmea+pONHj3AG+9y3GjVeOWU+Ne9AWyPq7+JQwHLsswDhyyMydrawtO8B1CseoqLE
4aoSPWpeIkrOsqwGl0hSY4Gt1nx0ZkosWTi7lYGciuIlL4k1LvW9uUdgg+q5GkGYGKrVhQPcisKU
c9pcw4bP7H3W6Jr1356qUosJGkEcKbzivbw+gc971Rp/Z0JGrKdIo7lyMxrb/kgcTIHd+mkJtaYp
kN4XwPM2I/3+hIeTgdEhoVbxUaJiTqIuWy714YwUkYjzdwjTqgkaGRqr5SjUDT9uYNFe4LABj1yF
EfRsUEUj+KOqTiQQmJQW005rPWGys/SZTIct20ujVsATm9HSSCmx4c1dqpTqJPBJZa12i0ctQq4I
0UtMis/d3ecpUigrGppoz0fb6QBzfd/oUjGk2wSaeWR+Sdilg4/plFXUC9bvT/v0Qy422au7xCZL
dDqX2n0JZHmDN9NHV9UryFycuIpAeXpmUXRWXwrrlfUCcEbWV7XkDMzpnTqSybBqs0qlLOYhikfM
d0aHW2lkZMarpHqjq6rSUGwxMB9GPGsXaBRYH/INO012U5eDj6LJ5ZJr5IOyKvR4SYyaAdhi59DE
JDjcCcosUkm5pM3+X9sy8IlaDZW84rRa11kt4Gy8BRTMsRFEtr+DSYiyA31+A9dA/f+tk+TTStTk
MsLSVjkHE0QIja+gKBSjT+V6wQyduLO4eF/LbCUL12zx4PEnon5PzZxGYJOrgtu8nIeOA4GdGsa/
zpvXoXYkn12UVvU44zud30jmaA/ISFS2zb911vFK0Ny01CajaLAeX+7I9MB69PHQEyREVHAt4Pmf
lRnlGDjeSy0bSLatTNChtkL28esCiiEeKK/XBKjj8aa1VfPjM+4SFC7bIsE4L7CfVFxYyPkso3MM
YzncTQhCwPfLr3sbzgaBPR43u3NU3VnYoIydX7n17b0v6I78C4isyZNjdcI6cOhwFtQ6WUVoVys0
BFGfwwHRWtdb7zxGUqr21qLomK800HD1ARRGTw6ySTCjCGqevD6N+WAi/kFNgFeyYQZ7GKAHuvJ3
ecQlKDqAjT0ckPjaEl61eoFbe73MNiSbi+EthR+94DG51jMZe/CDVnzkheacE9c46MDSc69L139r
9jd9yniZFv92Ve0FCXAymAeFUzWA8HASaveZw0wQr2hwZznC8jpZ6KKPJmM7mh9LbQMWfxQOWutj
dmUFjtA51p3fZ8mt7+tFAcF2nMKxSO0hJr35llWPLiv7wfshzpa6m2h2DPGYv+CuvKWatEH9bL02
rp9XVBeSHAZNC0wjjLw8OIGZKZpcc1h1DBfrpgqNTuFEt2KjGG+AosAiIUxvPNFcXL+PPg1WlaXp
EWjWyL8CRsCgtKULp/zRSdG+P/CXdpBeO2TksW1lm3Ro+uLGCNxPxfe4uP6enzTNQmvFYjKBsT1L
kqRsHJFvS5Ptsz+NBhDCV7O37aMZMSOf7rfUbhI9ON6OUeqiKueHo2jI8H3vKZy19yMCUEH3wH5X
XXyOPFNqe3xu7cvd+uac31oF7pvG0JDMVWTpkkXZnTe7vSs9J/KKIH9vKpRJterX2qsCcAExT0Ua
tBdtofzPEuAbJHmuGaFxuKZLOmztjtGf1XhOhbH3L2EbNdAFkr7QsZaHa1uioPXKkqY+oSqy2NQI
eCaMN3KiPgR3xHAPBYnuv1FN1ygTq9xFJ7Dwz+XPG43JSPlLB5lN9RCvQO2UsipHmk6pPQbDGveX
cu8eEZoGce0WxJVI8emSaa+Cmj4bVgdhzlF9cleLGNFigwrZsFpTlc3xE7643SNtSlNeDlFcF4LF
2boOMA8qkQfg9RUHxaUbT4F+/95Bh3/4VKtBYAVl7k/VlfCTpLs1t05aNoyO+FR57H18RRHdC+U+
piYSvaIGnOdYLbYqEzirUgEpFFbAnffIo++pGPCISr0TSC8WMplYYbLaRntlsz+eRLNqMh+qjlIb
VByN09Dh3RKa+ho+eU4lPjoi5S3oW2bkA+9+q70cboYNU8NjXT/HEQNaHW3DvM50CiVnsMTWmYRX
/08US4IvG10awfmz0h1EzSV7tD9HrVr4Vtr3EABqpIQQewNQZe9y4oaDTsK6ke4OlAupGVxtsKas
6OO+YQXJRbgBDoC/7KP06b7sE3bEyU9lzaM0sfLn2ablTBoVehIAq69WIHkPEkx026uCFd7VT4Zq
xpj8OcHwzwZhDongN70u5rww8GODcIsd1/2q0kdkSpt6hEvyi/eoxlfR2tIGRMONq+7OUIJFYLQ4
WHBc1ck645jispR222/bOCoPXP66GlriB3u/FGaxtS+PXZGAcDVTb+mBDCIrYXewtrGWlfuZ2v5q
40IEFC3KMVHb3zGxeTyJfXa5zPjQLDrdB4byxnjzmTVxfXaSYquyr5uwKBYXKRj0K2+5mkfDGVMd
gQrE40okHrKOyxVPAwKQNqlxy0aDvazqSOrB6GCxNDLh7K2ztYF4UoBTnYr1egms4c1aXGW5wDvL
nTwR0siC3MZHFUAez1/L3nOQAKjeDvOoZJXaHtdot3a/+EtMFCkkQ1Vvy91kWQ+HEOkkFiMvpS7N
heDKusa8u4TrQ15KUPC3oZFjzVcUTSMGA3SKjpYYpGaagZE3js1998F5nTCPZpMo9eMlN/pNHY8U
qF8zZROrQHNldEip5xRiy0tiVYf6CzR+um+jwWazRVFi5rAI7BH2ONjmIse+FaTJt4KiU1kWyoxG
9abQNQJ6+o9qT2E6VKbLrz64oNyidyfmyf0VwYdRidy8gr+U9o6rNwz51rPMAqtXE3WfSDfyYr40
5seK9kUBW96qO5vn3SeKE8ss3DeZbwzgzyxUxcSTNdiN+2d5g/X/ZhqC8sXdxjmTjQ0kwnPBaQlJ
3niHJmalNQ2ntYZe61Xqa0YJHk2NizMuG97gTj8nCeWiuwPIuijWehtIuNjiHLsWO4qqf5UzbvA+
mXRBcKTOjNj1QmwXbFNtOGCdyyrua2allCul7P1Hf4k8IgP3kXr3zKEvoQp23iNCHUmx6a1suaFZ
G3HxggLZ43rWAxnNNtAbZmwYJejke/CRbvBH22S61Am4vhs3Jk4FQnh6oKf/BcdfaaS2uEJlrvON
UZc5tBBalox57IK/8pNUhArJxZPs1VqfngSIvbb32Njij46UHwoXjsgPQfvLGQVkW8SEsoDdAcmG
3n+Jc3Jso5ImB2N/rJBTjgCZfCQ/uj5r/rbagu9+0yUN5rsHc4wr7wWfSQib+gITU4uuRBaPYAkg
3WFxH+O8Xs8VpX+B31mpC33ytUKG0n2QckqURR3iD4svnINrGvvzXhKY4o8NjXLeulKkbqJkyQEX
mukuSsgZ0BYv4yC0C/zoS+Tkn4ppyj69DxTOyQWebSvySa192hEHLDdGApcJr3IbLLq1/80rheRq
tl3xzomnn0iJTclWgC4CoCQ4SMNKFQTuR08G4NMAzDJjWsgoIjmCNHTyledrSt+fHKk+9dueychT
JIueiK+y/TPuE+bMGOoyUdfB0DSCNhu76Ne1rhAsnDH84gIaeCIECnY5FvrIHU2MiXoOFbioCQe0
JKIMEQcMhLhjkSpJnRNz+CeX7/PI/mLFDPiJX+kylxVcCujzgTxSYnnJ/ttSn0HWALJvt1D6IMgj
6SOeRP6h516PelJ+dNqjpZ8acrW9NkNyyeVfy75IWLqcI3kixlaZEraKD2dLcxjMWzplmKednJEk
MFzJwHPs7gJAnTbq5RzXP7j5597nGvx0t/oOH5ZOO8t/8h2dWO5icknx2OxmKrzlqFrK70RbhD/L
YONBvix1D9bNEEsBNB3mUmr2uWThSWdPGvS4wN4enO8PtyauweGjsJxEXNeivf1r139hGSUuJXQn
/O084JMh54D9ReyhYkxpzUyxKnQ5RjpVOFM92YFtqhrmxq6bfVC+wTrIWr9jNtjsyMiQxp+72BIz
kLgiKyezaXAgM534ILBKlBXZRei72gJ/oCzaDa4TcYIgN9AfUqgQOIlvblfb3/g1L/NmUFMm7eja
AKvFgR2ehDAFOVFiCGrxjBiBOCL2dLch3EWGn+gBdNiJRoqiTrHDjebsd0fslb3uqbDWvkjJo1tF
APA6mim/O5aKMr/jkO5Z0Dv9TqMhQDlHuxvPwZggHUx1xSqLso0UoYn5wH/2EI7UD20nATU4u8jR
mSYqrAemkCXv/v+qT7NA2v1ufeE5AlfbX+BT6rp4bvNJZH9jdlxWbcSBNmNH8LFZ0j4SXQev1L8k
sY19vDCVaa+gzOGG6X8XKzJyuiWoHy3JguLhAo+EZ9JOIe9CqSQdFiINBPNkYVK5hBiLDTtHjUAD
hcTdntZr1uFOquvOhnvrptXrh+XYAS8TxbGHwzFeDFboyiEBa5oAUgGfdisxAqOt0K/p8TddoZ1i
8PrGG5obXt8fI6WTTD5pJYAbfoRl3uHzFIztLZ1ye5EI/TYSGZNe99S4k4eHFe7qnmDSC/aH1VA0
TI816/5+n/uLaJnoDGa2VZQFVmvL528UL9N0fWddelfTApJ5GGgqPghh6fXdBM1HO6lqon5WNe8S
0WsyVFvROQC0Be4PRZLTSXCPChbZ51qML5jksmZUXTpUp39yQczlFR6yAmHMq1NF58POqHlW9AkU
LSD3YauqAqTz6pdvWc36v6iD1iBCljk0XjfqNsODAE+RP4poOHaAbqmEnqgkIMXFsIRR82kKup2q
4Rcn4D6P3Bk/Pgh5icnKENaDEo40tO1xRchEz2veNGsSjHic7d9DCPkD8sGRRUKyiDkWL/sxN0aU
mOnJCnP5LkjPBTd+BvpnVatMWza4k9npeNbZGHyyDrJgS0l+/UNVsbVlywQ2kqzkwe6Jnmovly3D
8jpzjqk5IqgOUdeex9h/ZhGoUDkv23aesbPw+OzR2sG4hRDyAWDDzPjpkFRqyH0tNXEAcv9tnJgh
6BJru7ycFDP6yKaaBXzNK6/cgvewXMA2pfndIf6Wh/FHU60NPh2wLZTcCUu5+WfgDsi2jL+21V3Z
9dEkRZLZ4ob/F5jtiqYv9v3rBtVYauMCzSjYdIvk4pwE79CKpdwhaj/DElQ5MS0PPtcGbixP/JVw
Lubb7vugDjkzkJSndCo2bD3meZLoyskxVu224OTaErg9cBPw16jOeeTCK2cx1ZTVlTMcv9xAo1zO
fpsZmUFP+rvXjFBRLm0zik3jEkRLeDNj5kE5kN0m7+J4Ifqmbx2Ma2d11EIG7vXIu14OyO7VDLAF
lYz+PdUqG6aDDkzFTk29ynnPV57s1HX8Hxa7Ua37LK6NkW2q+d7Rwm/SbPhZWvZXkbZhTFFmOayX
MZV/KexNa8PF8wl6Sai6s0xt6B1WxCj/z9mxYZQaFcWxZVIFkeeXSHdU8OR7n3CDhryt1PPKnefj
DR4ncELKosyeBgpwudAb1YmSVpJbdfRW/JXI6nm3o0eDII+IZTlP/Pzpg39ETB9Q3k5ipj2B6e5v
WKwMb7f0hEo/vfUjAsbkjJJB/UNPBXgK3uIuSaj8nehYYdz4b+vCUtR6VW9XTzcqjDBUBFmnglGl
smady4NjUP3nbmPGIj3lihj6yMVsms4jT4rjbgdUEDvW89n/7LzXdH92jS+6rXmtg2IHXPgePWll
CJDncd5EIQw3ybfJ5kigT2vPiY/bkOdFyu/k5EvoXeyd9bP1APLSouKJEFBZDhoVBPu5k7kWX05Z
VpdTSCLNzCsRvAYaprYApKsxLUl/H1w50l/EZ/+/ZxuIZtjpgVZRgoK5AYlR1+XB2AGckBCSv0Qe
2KaDeosVCaln734CXWPh0ioBimqYxpuTJGhhqLAEoXmN/e5jL6kXYi6ZE82JQWgQs+8PJEUhXLZ8
MrxkyDSWJF3JGGCvbWQrW15xWVnmFYkEGFnzw3IDf+TyvjjvymOaiytzhf9heAQOOQ7BG3IrdhBL
Eqqx0l/P4Y4ymmVFGJIoIoZb6plixIpE+FpzvRm/E/TRl/rnA8iuZz5klrAuWzufs2hkyZDKIw0f
u5JZZUWVhJViICEU9QHwJs21RgNfzAlB84JuY2EZIntS39EEr65NwbWzlzAJqSgWzkxQbkxg+NvB
NeMbIPcnPnbzmYgFBrU1OG+W292f7FLvpKLSjmUAn1K83Z5bIJPyhwdYEzxugdB4lM5SoJjd/4q/
/0EFV4IypFAthojwOgeW76q/RSfvzWhJhzdj2PGO1Suv2BUUO3a12JC2TvEnfCkyTho1hOVzZ2nE
O/96bYAqZGX0j252pjIudSNEtsagUXx6sYcBzY9ZfeK3zO7yGbVggtWh4i9KPMsfw4f6d0RRq5yv
SKygsLJz5OS3+AnkRo2rHYuEQjgC2r6GAy7LZ2XVcLtUGEmsb8myakjZYGv41uGmvHeeONGM1h2W
OPGIADvjpT3/TBMKSX5gKGbqgjLbYlfVJPQi2ngbFiJAN9Nfj9mZQ9LpCJYvrAf12Ec3rRS87Zch
wVK1lxrbsDg5lQmIctez+4sPsf9nbOLbC6P8Zpzg2cWFpTXw3+s/gBoUWRLuGI5gvVtp3gOhptgL
81LlKOaNblPciVo8zmJHnelWX9dmdkk2tJfz+zgYmd8nmAbM7TSRhRUlNh0VMFuGeHCyuWjl0uKR
qbwoCrQhyNI5h6Ws7de0xPqfe+lLa7XZjGpYet5oTxH7lT6nGcv7PkXDwhlfc5YK3ZluA960zK8T
ch2AWzPlA+VvoBZiNE1UGJy/FuVM5D1SCuLc6hBqQmTzhe9oEcT/Abk8E38+aLUH8Tn7yB4508eT
2ldIUZtTU+nz+YjuBhL20VpjadDlQlz5EAk7Ai3NgIY85Gf7PJWm8MCf0I6NiwesOjV0RG0kBua7
lm5LxfacS1Z3DVL0c+gTgMPO9GRkdTUCh0ynHxGyv+R6ggIq8QZJbvmavVzpD0oUtdd9PjfPxhau
GED+ANIaKCH+95BirXnj2yYzSu9nnZ/cm0Ir37co3oSQEHwM+4FGk8qgcCSF0Ba1ws/o15HHlcFy
aVr8f455qNhkAiPF5KeJdoaunbvle3PFO4k9M0uQV/TSawEL1Ky1d0tgZWBcaPCo6hjNWu1uasf7
+au/CAfY8+4R7rijcLaxeNeVfC3M0iCVCnSDNb+fG8QvQx3kwDWXy0Uif3P2U5VrejWYcZazI3xO
tt3n6/JJaiUiPN/oedWDpROzcoBch5A78BGENP0d34CmndSVuVCUf+0CR3G8kGZgzpZfy0oUXzYz
a107oLMIiKqqU3UkU1GxArK7thIyYjWaRo9vrLY/eDMmS7y51bklXtI9+BOi0JibcI674/amFPWl
7s994V0n/pb9PHo1rtLwV0JjJDIBlFZ9ejL/PriWaJzLB+Q9BnK2NlhZGKiTQtGOHJLCJ2N4KvNx
aZPc6UvGgoBZIDIM1AkqJ/5soYg9iiy5srkGHUbuMTwW29I6Ydo+5rljTr2DW7XNBxCKwCa41UXs
mBDn8TvRCW0/f4ZVQTiz6HoCcYJ2ONaXXdbv4OrxEFOfCLFiVBPHn8CecLqe5+4PYsApX04shw35
c12q6hE3g5qWI7Gi1caVMQaZU4ME12ZJUCeSpeNO6Mrk5D7ckeeo3mUD6/VuB0osS33U3xIpJXEA
3rwzYq5tM2QBoDmanSPnwK16cYQbXB1gzQNYgNGxA6q1Vk3aSjXI7HeIv/h//UKEMVZSFcDrg8Am
SwhzVFC/pzwWtd3m0gXk7QeG/TlSmSJ0mawwDlqFEQRKuU1ha5gMzQnYCHyX9jLnRF7VYMoJJvCI
fVgeULcUQUtNBCl1Q76fp+qA1uw0UECqnAm893BOtwXXcrnRHl5yF7YdWwAC+gOFvG3PSD+fW9a0
Nr563SvM9tU7b8eMhdZG0b5ikZutMy1NNZk7CXR/JzwrTpkNs2InO+GmmzSVuJukYH944uSU78Mj
7mCAeVIQXem9ldMfJkfbO+gGpfP3BvHK/BvF2mUjxwW4TG2i4NUgLj61QMr9KkTYzTjfia+lkJx4
8r4dkbfg0zN15wPC5wScUWOz/qW5QyDYiHX43fIqZxziKpPEH2mRRjKSNcmTgI0OcGCHoA3Zww/X
M9cyuGELA1zoy6oylQnPWINtKFwiv/OdxNEFcPdPkoJBdO9H89jTU7y7freJFVFtSZGuJn+OXXhA
8tn1Mp34rL8ySKt/8HUTkw6pqpn3/z1nCp6kBNM6KOwCoc8rQVglf7v5kmxuiA53qCMdhoXPqFO3
5Rcrhlk88eFcJE3fA6n31WCTxp8bf4ATwOouenF1EBQW8qfB+gf0tEFseA9KRnVyPx8PUVyieBXo
/ozE5L0HfRcHqBqB3Rm1fP5dmUsU2TvhyAGpreHS8JaZtgnMSaTM9VVqsDzS7eGhtHGyakiHdYIc
gcB2oZsif/WQYeH64J9A/8uvlyB3VvR0mWT8eAtvrNEehz9FGb8LLDBS+I9ZhVDJ0tUxGywGcbvC
gJHeGpS8UL4Gazi/6GT7VO7mGNED6QxoprSO+jaj3f7WGk8w7fBlXuXwFoN2ZC5K5meuYYRtqyq0
VfewNYHQJ0JKwHtLoqpQUH0rVNamoVzrsFnehuY5SE5LnG5XUyiLzVjlnDuvqOWkxsPfOQUbMTYu
OnrHIFJ4lym6xeZPHVTqmd6ncrA32HAUxY1RX8o89KuuEY3mwV9vHafEDXzD8VJnry7N3AcUoHig
2j0XAiM+z4i7zSQSxzY1NvGGQUnpp3DVhDgNBXA8PxJEILy4RtnLch7oVvZdBDujYtWa1HJyzE+P
QD/99Ulju0+fLb/6EkjkpZqfu7/cs98wZ9SM85Ga74BWaJDXZSy7JPn8Xdr2lw5tR79R17LMIS3A
+KS8kK8BK2ZBgemqOjLU7a6tGa1QuRVy8TYiZZJcNxOb514y0JQ1Eyp2wB2meIYmGeFN1s0XSHEq
jiRDEF3n63QRRHl9Rp7H+EYHOgqwAa42dRnocmrpiTOuGvG+UufnwjSw4hPVHT5VCNIdXKma7r1H
ZfLc0DEILr3FlUx/6umGTvfCVRpnI4xGc77RCf5kA7g5xVzDL2yh6Ww38oVY/vKeaN1TZbuzuh49
qQh/EMaIRu2B6ILRk8qi4TiHGbsSAJmIMDAANVDzPs9ssZmLM+f9zXLtNIhXB800nmGtDg0OTJmr
2Rh3Emzn5TnDi4wx4f1vK10xI0/ffiOoNJA533n17+q1imv++bvXpgpENW3ZYYt/GYBDG68T2ou5
BWDqLEotYItyr7WTF1a8u9ho2r/0xv4y2txn+sP/FVx+fQGt0aOCfvGEH37N298xRlrKn0aAS4VS
oCTblhqoh1QDB/uXSFwk/ucTzR5lhiSYPrjCasBhY5Fbe8yRwfSlagUI142/G63xiaft5GdG3vXR
sOM7T1CUf+VA55cNgQHk4yP7kOAiTTrkU9LPFapVnVsOM4vxBnBb2zcHZAc0r0acNnc4ONcypYKw
kdav644R6nUnquUqyfB2FiRDNi7eaV2GXy5PQb3aBubmpjgdbzW2OT6fOgBH38MCsYmQaRQ4pxre
JKOVRE9ZNgc3MBjWrzgeCPA++YrIBj0ksrV6Lli0sIAopAOO5eATzx+ikWbvcuZYSQRmy8Dh7Bw4
dhO9mrSyjI4Ohft/J1TfiB/wUCO6F9oTIYTtTZhdoPDMyJNfXXGAz9vP3cyIZsI6E6XW0nyuKc6C
z6ud2v054xlbLlt4qPH+eUKrIIIIUpoV0UC9XH+4TCmPVFRBDLdyzd+gTo1XFESYCpqMS9BxpbKy
5keoRQRH38r+5LbE6WzTryE6o91MJBs1caUf+1e8e8y7RlVKcA+OkRbsXEjO0D9rYpaztQyc8nwf
ep0urkpB1abh9WeyXddEh+aMOv2GaJ1YNPwiK3ex83G8Iuo+Ti42Ibt1e3YCgPAHSs2xOXqo8wfi
Z7xDH3xIfhx0KSP+WA5prdDbV5cYz91GqE4CtZOOsLFT5GUL4XwtG6GTS7VPF6xLuUWl4PvKqXTg
SIL5/+BrHmwwdgFVTJhAOP69BwTg48AmINAiFShVnRPi9/5eAV+HqJ6NmHEVSCBImGXNVAIX6HKv
vaeO/BIQR4xUdodFyDyrp3iTyYoyAqlK2XkuQBP1dKP24CwQiaczD3OP/gg7g7NOBJTvdYbY5AX7
YJ/QaLfc4U/DC9tFC6oYhoh9dWEjD7LQqAqj0QxU98vAeUPzf0N8A7uiDhE1PtSfwOr9tmqsHCpB
gf2dwlwBACgt0BEMRlwYBg/T9en3Qrm8RSl3AYxCKXHeKjb2Z20zEIXvXdNooFh42rS2YXhLDQie
5ddw7WeKHM9qDtNGthPnzvkIwVDlMrkTYi+1RPfN4gvfHbK1Xf/u3YchXeIQyBp9JdDpY1TKRFyh
6aXl7tp7bd97uvPLe2I5EVFlkdGoKbToumdFRDgUfcBR+bkM2huqXaBuCc2zKF+DVenxb4OunYIQ
ZFTi6diQ+Tx0Ap1h1v4ZmAZp1gMOGx9A0qqVfAAsDgAXMHIihEtYzPtCFnbjPJLQKWvuInjpUgx9
Rz91K2VZw27SRl91CuYSpJpxovJyJW+A1FSE2k0Mo1X6g+9fKHfAUPq6fDmL8rspXCBhEg1jImkN
opNOohG2n+76GAvOOZbo9kRYz1YmDxZUpdSMCrWtiyG1XTY0gfa4xsGc2QR/gFnQCtRsSo5xiwNI
o4U1Lg6Lf7pVZ+cebbFDdwxx6qmmDDJGnOK6ZSsziRP00rTYM9xn7SxXGTQkIgscmtS5VvwmwKwW
le2Fvyjea1nyxzDlqyvqtIUPcbuMiOxAVkQZKB33wuV91w/UMlpy0kjSpH+yifkJVFpId3kciSXN
j2MO0GgPXsnyka6Fd4kgLTgH9Y8DwHCKhHIgnz3SSQ5+QTyECwPv295Af/ld+zi8Tit+oOH1sGbM
tovI7FieEyS9aTIUR7d9sUKT7vCJsJqwUCku5zScaaZXiCnGT5+6yLnF0ntblRXunz+ia7lU2Qc9
IOgDMsGqjBu0RMPbjzpvcsGBf97O5w8lc6APMncE0UXfvB+uGB3mp+MeDUO8ptmU6FpxkLT87vOk
Oo7D6igIaUJBrGK0vc1NJSEi5Hgv986NIfuKAfcqJvL9NzcEtifLrrElMrHqbuyYwGxFq30/GT56
1sEbYnfMwnJhHq4IJPAgqMSxN9kPQx0M7qnLDXig6pM/iWhqKWpEv0QprkDgVLRlAwFVkmaCHVUM
Q0Ea1szi66aMHgFNjxxNo8pNK6BHOkZHybze7YtGVdpEvwpEcKIDSEywZ1qMWon7QCTxeZT5vP5p
ipUNUXOzmG/eBXfrR729UMhff1P6G8nUC8ddkLoC/UZyQFcgP1rhTwV0qHVVanMINQluUiisgpuI
NFios+XfP4JJaN80USaprIz8Av+XZ+rIHUjwPCSR1OzpPUybI7b6wWyLT/pn0jzgo5AuQnhYC8O2
MdtWTpuRTet4BaxnzrGt8voACCOYWo5Kj7xRSjJrsslk8oAZxwPyH/f+m9adqlutILo3QL9sT2c5
kjgfhDqZZnK08Be3Sw2A0Y9oB/WzNlW7sQszLHahbCkI4PYLw2yW1mC8y3DWnW/KGNvBnZOhvHMZ
ACMo5DmK+znvhie/8vbNzLDD77uPZPVVij6uKhq/02qj97bNO1tAizrap8W52j5z8XS2zE5uZlYk
rBrM/s8RO6oLEc+fCMP2k50lO81QlYyflhtnMrt1qmjA0c4cjdt4h5u/dNdLqYgT4Rvz0KMuJEzL
rEmCtvvXHoaKRQcRN5F9aHWqSP1yCt3EU4UVB1MqWSdbJvj9UDZ/6hv7DL2T1lpu/D//TKxfS+WI
cbG0whAgZdqBvmq+z1ylke7kXaMDHZavpAqXzUgvPR7r3dqYXDbwjU79PsHKaRkrkbXg44zjseKj
G/ImbRxDoBvJ5/iZ3+0ECnKaIErmHFnOsyC9DwBDbCOpb43MLU6vtVJ5QtGQ2moxmwiprhFhhLbW
7TwnsME63dpDLDMLh1gLzgVcwTMMN6XDPpaov9s0C5BFnhRIBj+WlTXE5FTcAnP7E7oRGQjKdW8L
UOgeCQz7t1eV1ZLkEy2qr15A2jpie9rR1STh32eugy02wPJVQfGqi5sbx0IXHUxSOVsd2P1mR2fE
GQ5lf37YUYXphAu0b/vpZ1CKFdTG8NUp6y5yi3fEIoYoRfeTu8R1GqLhQ0CvqttK61VXAAwKGusG
T75oHLw6vvycPLN9A12X+5FpxmSJtB+bhTjJxGqJkLqNAc2AAgk3RO2YIx//M02MNnX/ubHLOkIq
eSGp3myVx0igxlWRHr9rW95FrSHN2MOxCOCsenViHFC28RQE3VcxYhAiKxGYWR3NG5d62ca6tWrz
JMF6pvZ852WHJBw6uW1WhSulm1Ig9x6iAGWC60llkq53uSER0+M3PY9wuOioKwSbhu++qK2IAuEA
9E2cUSYJk9b6r7IaNtKHY1D2a6FW3y1pBujreDTg1cWOshJJ2hEgLEQUhsfiDoZbThxtB4zILHbp
iqdGtjuO5sxmDTVg8NSqyQw/x8C12uweDXxSVJJPT5IAuW/uFI+i7KslH1waHUqYniS8wR5aEeDO
ccyPdjBDlYgEFULyZZjS8NTDfoCa32TbJN75V4HCKFmxaPOSL/d5LRjGP0jW2KRmlAM5IcopkdXu
F/uC3sWQz1m9sxGUmGarQesNfNWtJlceBgRzasxXvbt+RdGP1GdcK3Oi+CjW75hnEu3XVlA2A2hc
5TV+b45hRVl9vEHToedB0BNmaUDGZ1wm6BGgPGi2Yv2URuHjlox49WKvvCliGrCycoh0iz8nfyNu
TxlLPG+EsDka+wpalqwrDUdAE8N4mPhhOFUDZlUDESrlhV4DLYyWEd1wwO35d5agnzun7F/4Z4lQ
NPc4NXiCc/jFDC8x0ymuCYCSgsXldbyggCv5OMxVgftIL+yBhNIFa2az+M/aCw16RCcGP0MD1s3L
dUN/vvu1CJoms643zbUx5dgVMCZjxfVAvbFqLla6NXHi/rgqEUJg5lZpvYOCqU6KYLsFaQMOey5i
elvUmYJL4jJUvD64tqh0AYrEAANS1Q/51c8EAbu7Z4Edw54QGTka3nusl2RO++3YMJvccCo3VRk5
S0GYevj5pj0PSz17pRXs7lgNqCvkLWnTCOemhSaR1gpFOZLfedLV1IopPraL7OBkp1S/Tlh2Jv8d
faVy9S/wZaGCacBxRa2vgL8GfkygdVPRswfz1F4PaTOS0epZDktV/4FRohEO1+38RpIN7zJS1GuK
/EzOSQf6FMW5hDmJJfPa9Tb/3I9DlasjGrkgTr6FDphFxhbk2Xk9WicY2bWGNUKpLenIjgGA2pzF
rQFvq8RFh7x+gRo8XeqFVUoCinzGsSOS8KXdPTje4eOFuNbUp8XzV2fZ6VIZes0kzyLu487IDURl
r8bHKqAOZULI+I++T+Tf4crytB1K7AXHctrh/fpjSGAbKuNsdzOQE5B4knubhXIdx9RUDEwR9Z4m
SlAr9Gxf4EmwlpGJI5B97tkghVkT076KWz2jWbhq1aWazaxHtuIEHLUDMWvOZ1ywoSuh2sfso6HM
gLL2Zjn7VmfTUstvxIjArqUF7ic20U52LH5pMRBtzt2GvdG3A9ew7npeijyyyK/s9c42a90ryQAS
C9RkG5JHFgeYY7qGEnj+gOvWFDzMxwakOiWhfl/oCbLF6s951k0l2nkrNqCp/KWbAu9rpsedEGLQ
52y+EmBpsUcMIncU/AruNv9jIcIL6mZQUxNBBLbYEU46Ff9+PIUexA+w8WfATaE36tApOPaFOy/R
6R4xKS5p09+e5nmFInAlHJtJoFvSS1Yd42eED43vLhg7mjR6GqggtZ5CDHCkKcv45Nz8s5nhosvH
b+n2uw2AzSH5AFWGGDwZEfjBX4k5nxFW1hR32UVNb5xaYA2VFI9iP8l6z6lD6pzTKJXpK7iBrnU+
t/8N+aWaHLzmplDDpHMZfMyzMmEPoEc7hExftPJWYpHlACXy+PKMZql29PlsLfgXSYytizNYIN9d
pDUz3sv6AT+E0xCx9VCAR8B/kgLUztcrWcxesQk+IVd3Ji7xdO9zdrqRkAXNSbKqlUaL/N61YMGp
g0b/m8NhkSANm1YJQ6qbso8HYj6tBUoZgvcpbqhFv+Rz7F9yzFG2ecoGkkVO2E5mIIp3xik/Sbn0
NZP0BUWKR/s+mLuIGPs4hIQrjlSyDXdh4K1GgwYdidqKyGQFcATTaL9YF3YgOQKEFAvaFj7sd3he
B27/5kcIxxEW+1x4nl+Kv1+kKSVQIhneoKlblOO+snq+GsrB1T4IAR3UMKHnQtQ9NQrhd7symhHD
l5EnaFEMFUy4LCj9LctHfQxAjcwiXyaY2UDTbcH0AuaMDg02rgsE7TFVSh41usj49rFsSLKy+ynh
E49l757mPmB6DAmhBSH9VTYvwKKTBBpjcZtZKMH9csf9qyAiuOVn1flQKRyM3hFvoYw5mZNxFi2b
48sPC8bwmIa45SUVLWL2bW5RdDngSBIVRo3X3FGtVKuPtq5k8+i1saAkXU2/qUGtB4qjRx/MMSbd
YtG9S5DpYtaRT9KEo5FrhAv/7gUlrUzlIqpOG+Tb6r5hQp0xnPf6JNXYSOYF3FhZoev57s3H5vvE
Vn85IQW5ROBkRipfTBJgfZ9l2kQt9AWCa+KHsEYVFjO+/RmKCKFI3cvbsXpzCVmCfi0i4SX5TSd9
HLIE8yW1VUXpYGdOQ4+6WnRgibLdNreAwngMgfGk872IsSl8ZqucKp2LCIFWkA95R0x5Y5susT+F
SqQKwfrYiu1OA+n59o2ZmJ+DLSI0Kp8GB544O95fZZzdCBwPDcaAzliEC1S3lXAtJYygcCXYjHjl
4MTfn42VncEZhEGebEeHWuUmpJVhot4evk7Le/OjSoXlC9ppeMquL7k6CkCD7hvMCgWKSU96IgF9
XB6FVHvw5goqtYd1jje0dCRbLsR6OyOGg7Clg4MeB7z6nxKdUQq42R1gudIRXGkdeWIz2BgmevSV
0/VjHMF4Bq/lzEZ0jFMD6DQAlA9u/NQT6GdKlISo6/odGY33W73oob8hnT3nI53dMxBBpaquNqqB
SKHdXoq8njXJ5fpv+udSJU6GUVMbwcaZBmTEumyggHxbmiuppZirn/dh/zeN1NFKnhZfwy7YKPS8
yYkEJ/1vlJ32w6WwSBhd3Di10t0ycbFguYKTZTGAop2jFmnQxqln4g7HqzilXtcObTiKcHUJ75aJ
BEjcFcu6QKs+CV0mypyThJQZ8eO/YSvXsoSDsSGP5+6cFv5oYeGMzkzPgwGWQWvxJkpb00IdGTVZ
vkdc612fm7JfdNLBnOPYikyXo9U9hQ90KGPd4nEGTwq/KsXrRmSAxGt84UwEdTVWgTo8PjlZCDjF
XoSjbVm6yGhRBS0RV0GBce5rGs0/99OQOXqt+TIQCvOsH+PYi/2TV2uFSqjnbhtlzD5NRnftd0DZ
TGCzNGb4k03yIYqoPEf0ii04k1fiykunR5LHihRs54viB3Duq1OXBholCQiu/z4xBZhsy1o49TY7
zTaGUnRKB6UpURr7GVOOy3nOvnUeM2XQa+XJfUeuvWEpdVdSipdsjtAxf+3jq55QigzqB4gECu2A
/Z95C0X6o21kB6qmn1FUe1ALNNn287BwOKUC8xGXS9gYj28ikhsSQZg5A2I1PZ/aEWCutqhBixaq
C3YLUvx7Z6ADMXGBhuatAn79uBPJcYJIiy781VoZGEnshPUBVjRLd2knyb5EJV8JLE6f821CrsLN
BAvOQXk69BKu9oOSUzPVfhC5sB/xQQNAdJZ+UEfdrAhXhoS/kS79DcwVWLHSL64MdQ7B25ZHFk1r
defFWt3V6tuAAduHvMoK2aUMiQ/EWuG/hh95OXkDRrjzxvkPWy6kt5lWarFMPoLy4wf09qgCWlNb
SPEVeoOIkcdKeGty1Y1PyAEV5xVyEV+NVQMc4G+sTwMhjTSHDzqO+UtRo51DK5XtAY92n5zBwbn1
1X+XF9LeSB9W0w4+po0sPjYCMqKJKhqqePjpXrfnTWn6Dnr2ontcvokyWyYuLVsFHQVO2IMKsuK7
qw84GFxGMXymo9FwG/LA03wXSa62uWoY/+WnpPjQDIKSoVFbxL3OsYI2C/hZxshiw+Fb3xFhS/Pe
yVypZKAVxAVli1zfJaHHqmotwsmmjrRJ/32p/tu+tP9BHF/8fUfnDT1IwSr4L99SP2YxAgLFUH07
gDA3o3/TFGJ2dhjZ1EH3VicNyZCmVmOctgVZqLaWDtHDTSLIw3Bj5pxkDL6hZXVeTH3zVoIqK5yi
aL/AQCHLlZHBfWS+be4l7nyoFRMv19Q/6IoB/QpLiwFwRisJHSsI6y3byP+Ye5KEBI0oS/dZFL1p
nVmRBWQF9aQjmb51dRCtEHUkw1njJw5bZYt/oLPpqTuTaFS2GSEb7mWV5TkZHCpDpbh/E7le7qpZ
EEJ4KQggi7r9vP5VA2oOsgoo/Bd/tDU1OPu/mJ8k1Mu1i2Zqw/bn9J6GPEgkOZCCCMNVM6x1w20I
kwLmD4vRB/uMhpO0SfKsebszislIq65+SdSVCvjvwm+H7H1SBmwLhXVCNOHkutcId2dziQ3bnOiM
EsziDfhStCwB4qc8ipIR8zOqOV+tNR6sO9NfbH56SfpPKVVVeRNeBXs+QN0dyKir3kA1uo8UOa3U
a1nN+h49hZd/05R72JpbTStrc0j0Quzt9nSVER1UoVV5gv5V92GNqOEYM9D1PTOoA7AXb00PeqbH
Tl5wtWs7FZMVzSLvlR/Mp2/YwNqM6yriE3tY0kUQuEW3eHXBoJ8sCmhHKnsKMD2pGLBJfe1milUv
+GGWuOiSwbLJaKhJR3awP0J86J8rLIO1cqTX9sxrdMSSEd7fRKvgm/9ba2qJ6g/YOLyyrmAUx7oU
QjpArovWfR01n6GOk2GVlEOlUQni4/v+rMFPEeFkmXSEfm3R+2r/+3LwxHioXLkK2m0tLpo4OxqT
HsCn3pjJ+RK4oX83/TyZXNhb0b84r42kfrdyxqMErTmagvgd9deeRBm2HII4xOgZc0UL/hAIjHhR
VKFChtpIL0+A/nAhBWIsZmdBBvLpeSzX78UFK3z6RTo78JCW99+EXOdjhHZfLdKn7D1nNYst1ZWE
BcmRpdf47SPCTyJvIvSzMkKauZZl9YYGHPJ/ou3R9fa+R6GYLP8nF0WIp39f6BnLDpLhDf5MP9YW
oWpT4gtLhgyNEH+1MtqcTPKm2r9DBDrFyJI8K0C8c2rSzpkM5JQGJrJfUtJbiRqfd45aZKlSxwcX
RMg3Lm1ZD+VegiQp2ZqVDykD9cuKcnNWlWozBrsQ0XzPuW9Fh6QYG1YCsI83lO9Jg/aykSM7qE4d
sH4UUST3Cak6ueyJ7I+uOjK+Gy2YzPBFDl8uTJLP8Gt6VeP06WLsqAKJj+Fam4XBpeu0fu3ZcgzQ
fQVuxfUoJpBr2egA9RVw4JGDbxJS+myFctNzoFF0uma4pBeI4dl82hwMO8bttuMClRTGOnEaRaiA
ETaG0tGLFz/XPvFeBFVZS2M5qu0zdoPgQx4n20muf+yG0uF7VppRFTUT+AOjOoWRnEsZumrpCd0M
vVlcHyYE9RHDcCtD3MCzYFypInOnCJlieFCB+vravo6oHD3K5MsnperQIe4RjIVE5q1toSROsEQP
c4idlPRGQJTwzMzWHlKwLqoBkG4fhs+x4+EagKcHpkizLiNrtQ2CSeOCEvGDp7KvrwZm7wg/oLu+
w0Mu2/6wJniQRNwXMh4nAL6mEzbrhwal4tv+Qw5rlq0KfzC8/oGJD+jeK72xf+vXp6/KU8z+wbhg
YVQCED7PhEC6B1mqFdyw0rUJ20MhvCwaALBbLMzbcgdGm1/kYie/qUzgeEnfOvNl2tmcd3+yiMnM
X3xlwla9/W7krJ5ZM+2hKyXOnlMWDvoE2t+iA0mypp8jjyGfhZ3QaY6cC4rLqi797juoaasEnbMW
1kzNmG+4hEMN6zFRe91xyIdAZpK3UskEO9uw/JWYhKvCw57DcEjUMBIcDoPvNkgfgLwm6xfcJVes
1UB91+7NYnW+00HJGKTb1T8ijtwlL0pV3x3VFDkyh3IefMO3ESujy6kVXMvmjNCiJEKhEor5iJQv
UaXLQwVf2TrpPAcukmSIRaEhlcPC6RqEGctFPMSoJ2qU0Q8u2Rnc7RJqMrCj1IrcweUa0Lj5mstU
7AcIq5T3WmrrTW4k74VWMzVqUvUYCClEXuYSCLS9trUdPhdgC1Kx2pqZFOI+qZa1OPJnT/eDZDfS
k54+JHqPMSzfzhuMrIB48BEnJL2HDtxlzb1te5ZRbZmXCgy/SBQ5qRTjy+NnLZHvFtr9SBkAoGrO
M3NDi5tdWszEqjqxIRX2eLki/2FcwkcmZmwyZiJZniGyzwhqyADIBH8ysHbH822cV9FemaZ/6XjW
+awBmd8qrKDOd6SOChs0EC1vtJHF0qjdOU/G2F+VyKuZhPzzIXP2NgY3ez4TydrK/k29GJK5Ra/d
9oWxxBngHNSwij4gE/UEK+NWov3kxR0sImFuw66PE4zE1wCwVy08v+82kYNnuV08dbJrLH6xG5oy
DF1N0z+FAr00258vq8ddeIHu8I9+aBYTQ176wvosuxJmvO33/m4GbIteyfHB5VRr6kYi2yL39tJz
t3P5VN3es7wYr6yHdW0mADRmB8BDxrdj0VLDCMWxbmxMvde+C2KCR0v/5x8gJ7P5u9EFSz0OYp4I
uo/Srg38/et5796l8cYl+T0zs8rQE9TRbYHIL64m/M/99cJTDzqEByirvpgqWafqTUNkEcyY7+7p
mzy0BPlAZBs1th087vcYMMvhODtychqP4pkpU6t56RmbHz5QcQHcECBdYf8YelI74mIVYOJshhOJ
xqtsLevjcktVFqmF8AOxmpO1f4nY/8WE9PGyoUurWOB4o/kxLn5hm+09VOVUjjS/lDwxvHgIHFYt
Uttj4r0t9ETETO/rY2Y6kd4QVswAHPXKBTLcVCXEFuC7gyNTMDbIkExff8O/+Ccbz2GBvWQjZjBp
CkOGFxE4eJ7N+TC2mCfPYagD/g6RjsczMtvzwg19dvXx8xCuEeUXRD05EkjAyJhVmCdv3IuDjSp2
KYpYPUwO8gDLka5L7iIAB1RNMZXCM+gaXHux5xeXqAxn5J6FZOoqAhbTqUBV5zu281IKwcB3WyXM
fb4YL5YCKg88ak1T59yfxbjfZk26yym1NDdilEsTp3gn6LKMhuH0/e//d6WNmIegyp7IDva9z2S7
XLEDvMlhDDdfeCyTDVQ2MldbSrZled+fY64KvlV3p4aJJqdZunP/6OKKH++ne19n+RJJV0N4a7eP
wLSC4CHLTDXjAZYAqh73bhwYCK5e+o3587zIQsu9liCjW71jKL4XoiEUxIhNTXsngD+1HFde1JN7
DY4Ge6xkXL0KdocBeWIbe7vsHySknCiVHmvWRTeDZrIf7mEoG4tyQa281hz5kNDL6pLOTo8o3QMY
6r29wrQixt9nR+fsF1/sGoq/FEiIVsqFuYxclTeQX3cGNE6Hme6ts7aaP1g/wZ/9eLW710Yv+9pS
FTft7f0p1dkbVmI6Zss8xguqF2D3/ebFo+gpqHkFIqKuOz7DkXGl/fsUANJcqgd8M6dUkp8tCNkf
zlk7UXvgVRut3SxpKSz9f44Jm8FrOkJhtprVfIkD0K9N2HObbARUG8OwT8/9N7q6Bf6DdHgsZQJi
R8fYQu7fxNji5qdQtv80UfwkTgla4SubycSe4cVbslSkb3hUWI/MCluREos15K44Px65DyKN1/rI
rvnPXcNoStVD/ZRhP0TrbTw1IA/cI1aUHthled4NZjkXZMc3HJeXYYwix6mR1GAiac43R/NZdelE
kdqiwN1QSagLCPUR6NNUJPAbhyGps39BB5qNQSfORlh5bQYl+w9WUMXK/oQnBjOSNZt9dcPbt4oa
iNhrROgQg9cxEs2wu8EvVcTb+aBT+JuTljpM8FCGWnTDsrEmdKSrN75CPPQ3Tyz9r2B9YWTq/NQn
tqvZh7LW2C1fQ1dwAgo0osVd+rTWqZXcyI2Qyp9N13PMK54+JtqTEy7wonkfq8YiD3TNHLMn3d0A
A+/+mi1BZWdhxalWqWh6ZgIqm52y8ScoOwSFBdktNTWUFxnOCg/+UcBOqgSJVo0lRMoi0DIjj5Mg
wHwgWnB1vwtZrNp0Ai4qF9tD3RaB3k1ikLYWJph+qPlxTd3dsMgqDtce0tujUELPlfu47jDHB4KD
6oKpxWs9J/97zAy6rYBoHgvdZ20XmD/W5hbN9UbTGzndfvJxOzR+R9kbgPF1Iq55wahcbjY/8Hdv
t1nXJwF8lfGpLbKlroxXJIa3+LBvnGIPNR112Glc6N5LXVINkfJgsB9glQndXvvYqqNwdpwDzUTO
UoFnmLdmwuSCFbfsJrRwPvEEd9ItuCmVRm/3xBU//iQX2O27Jih5kIfW5GmlNg/urBdlcbJPiXrF
IOfZZ0ZyGtd9ghp3tWYhQvhsJlavJ7fWZNaiAVGNc5PYGrKfixrHwBQ9BklLLJ1+WMwijgjJJChj
LsXc6/8Y6ZXIZln7tjgqtjcBQNbiXpr/7F9W9+rBNK/odVkV2LzsNeGZ86dUBk6iFyTyduV4gLsk
f7owsKOHPbM3NMUNRZ20WHIErvHwS+/BRVtGD/kfqdzGu8uTuXDEbP9caeC6z1dzM2P0RO6Hnink
Q3fcX1G6igmFwLfxj4cWbqjoi6JfLTSwjJzrwUygMJQ94iVeQwLLcqk690XCRtz01FYXona979TY
52Lrr3efmou7ykLoxngBUHwEqTFZ3yXyGOGEtqUeF0S3Oh79u49yRK26SEsqobj4dkF8eEPtojEg
W5tnpKldjE3U47tIei8Eqms77F1gL4/RrrCKusEE4q8VxPf+yKu0HdB+8qXN/zXlM9jhhjGi9SF4
7Qt1db+aSohe8DUWMBEwEDkyjNAneMmp9is0qft78VcSotme8M7+h1MS32NF8PUaWzjVg5IMgu0y
2CB8ktXOy56ztXARlmY1GTbW2IFteScC3RxrvIgJlOa0NvUNc2uORtzq8fXIiqIc00/S1t3Tp/cB
gqOETijweyXO5cM7ihDLvAKbNCuE5LuE9VqexB1XyMl4bHhWPKMf14HJsQaA8XzCPPVM9BxOFrgU
7QBqy7d11ruzP82FWLCUHaCmtH8LdOtvuM9o0HKQ0WICUMoKfP7R4zVsf3CDH9Ijw/zDygIBLO89
dVkeGvmQ+YyAhP++7fLhzAVrdyI9SylmbVtzW9p50WUelPz82UfXorHNXc2gbyzfNvVJ3nzIvkse
VpJHEABDmGL7TbNaxq9Vi/GRdRltPJOYKyRsy1p20qiv2fdmBVgqARI4KFp/emZ8xp+ozH63QnUP
wDu58J3Fq8e6tIR5P543hxbFwQnMxujJ5hCxOqos7jBtcAKNrzXMK8btHQoN9M4HjiviCMAIotf5
iooJePsWNtI9A2JoiGf4gUPdqx3AZDaYyE7zSuo0oyfd+oXka6g3/e9v8Xtp69EA6oHoyOpV9TEV
/nLr/tb1BxqTH6nc2yIB2YqIXl8/16/AxtPGMltZwOH9YOlMYq3niedbYu0DUydZo0reQ6VHmqzN
Pn70z2e0MhueAq5TkyODKmDkjREVWRN/uLGi8nhWT8C6SB9bbiQtPiNAf/L93SYGLzJGUpJi2lm8
lYlHC3giNGkebDEydxsA/2JChBn62NkaDnIZT6retZCyqLX+zBXm2PqlS4DfTZYPdM54RrYurkwQ
eTuqGmRcEPjhJkz6BPq6D1mOQaO72VPdPgndFq4C0Xm6FWVrL5PoCLyOmTxI479Tq446b2hcSaPu
ICN8g+baM97l+8YYFXu8+ZQLvnNynQWXAkJ7Ze5MdSumr9/9N7BjhHCCJgts4lX9oYyANAcHJaDd
Hu0Z/FDeBNlAlmjLivDmzsvmTa09+Jqug68VJ04mrRKvytCg0RgS2IQhUkzN7ELDxOmsAPyV4F0Y
nH8ajYlyY7u03+bbJv6blcicpFXt3e6uIKtr5Eihw/xAp5bnEoFnkj4ZSOD6bQGuMcR/SpZpmdTG
L8aB6QHWxEamDYnCJko5pa/mCqK8EQTdJbyQlISXqQj31GmeuVCyInF0fs+vJs8xK5LHiivbEctq
QsN92fGxzT1QEUlRnF9S5J3/30OkcJNwVDTFW+ZvldC9qmMtDnMdRh1WTajsjfFzMuzrrQavtV3s
ZiXgh3CpmUgcZYRiEQykEq8JYI8RtqT3rJMd+34cUTl1Yg3K9yxPCyuckKgKsBW0WOOm8pwhTHMg
F2YmtomRnTFZPGWIkQ1nZi4fGjicgACnmiqANm9cYUqYblXDPocdavkw5m0nzumMdf4pXFtBMDdS
dfDlVg3VeyZZ7KM1ha2oXcc5tHDlK6BR0NrBXJVmY1wAonjWo7POZ7GPI99MPsG1buqsZDiLZ2BO
eTG4R0f6ZrXGiXeaEtpLMYaLYZ2REEm0H190uxXgmeb9hKI92bpgZFMmpNYb2FAanImBpOCT+Mt9
0TXFQeZqSJ/VaLcoijm771DXeLl7qLijhjoW4I+qHpiiwVdd7xe1BXZ36Uo1yyzQlMCp92qNV7nj
JDKT4GRmQteOCX30S6+5W5U50IGdo9QS1kiWdP3DoLKC6QywM1BDcBQgI4Xutg5CqBrA20irGM4c
XmopY5AYEPcb647Rtnx83XoeD+hR5GOMgQHXvGxrgDsxMt1LF42VgctfW+39KQgyEFcWzUqy4GNL
H3nPEQn3JUBU33GbEimsHx4qSIEEeQI7bf8mRiU6d0fzgQhlmK7fARVm0fReeMUlHMofm8gKwfc+
vvYcMm0K6O4vdyAMuugtei6lFpyy31KhgYIhnqrzXyo46ZpXpY51OxuinEIXfuTrl/Cw4Pf4fKC0
3kWq+4Aq9G8484m+le+YpR/kSjnf3rpcGnsebORCkGls6eto0sPqbxi7eAarmms9BmFrOkDUl+2O
OsIZaSCqUMbxHXmkRTjBRTiLx2gEpn7aiyAB44LmfnV3BHt/YLJ8juUG5gpLVBNhHN0pgfOSXUNX
MLKXIAHqk0b70R74bIKnQKA8RIDndgn2DOMj9/A8E6yRiVBwpwPy2vWTVwEk3lrVF0gnBzsl8NiY
/NhjfYZ92dvSfkThhLfIzg45I2hwXOLhV03er678O5tkPM5U0A4p0TBQve0h3AReQ7r94kvT4u67
Um5ruQgT2X/BWoa3AHC3bmfbfrseCuWCdYxW6R8vQ1K+sLxavwFyCDmOg/pW9Twdx3d6GsrcUE+6
3iPP49noiAr2NUMqGWVlrSDjD7A5JGW46owZt04z4f7RKmRqWDeCe0OVxqaC86Dh9bMsNovfh67a
6VP2Zvnl/EjfrSVbq9FbZsZu3bjuJhT6x/Ghda3uGiwMdiyrtH3S8cvGXo8SU8UGof8T4lciPRpm
0YfOaZ60i5odz+H+azD7NaaQR7rz5pPzMN6MbXH0ksiZRB3aZcAw3iAUWvI3NimvOU+0EvMaTSzK
+bsSl2RD3y9MNGIfNozY02Ex4YJPinPfc1hhSpCJgMF7hY8mpQI9DjL96EdzuN4ej+03Oe2cmDPj
bN+syMrQ2C5nQcU9RtxArbNbgY8rKEQNsNnHhjtXb1vXZnf65w24yK2N8WHM1MfoTc51aOhtKWSg
qJ7W8I7yhVZ6N/onkNjeSuqSK9n142KfYxP5ugtMxfVGU95TABlcXtzij8ix0Z6O5QyrKTBFrQH/
frsPE7kQVkW9eH4S+gmtrKmj53Pnopq1zAWICj3c91WNBRcxXUZvVEjeo+K6DBOdiOl+yo/5wuwG
4VRthJ69ijH/OSoOnPHKZZsmHf1Qh4RNGSeSoXsssO5/1OrtE1+yZf7Xa6e9cvkigz9qsiCKZLdi
iwxE7LmNp2NnpTeuYej9WZVgSNL4Jx5zmt5RNnBr0vYE3hQ8FtU7poq0LCkK3jGWmxgqHHDj0fQb
16OICVLT4BQXZ0/Vt7Q73sLsgVVpFC5tMVdMoABaRKKtpdzmvNLDoHO/1U9sxgv7mQ2wTnskGhSB
UEFeQV5b5Eng0MtDUcP6atc7OdjOlIKax3Yn3H4fGoE6Xfv/BAIVLMECFKSmj6vtpQeZ1BVqFqJ9
7miwBEQ0i+HfhZ8WZCWideNZ0r9lhiXrRslIbAfNK+5LtkSgkxQVslloFdLN332K5cKhPXBROd7R
+YYERpaZHbxHVGDReFDIl8STHgH5JEj958Acwx59kKQAsMFo/O7g6Ti8Cg8/s58zfb3e3YE/A5Zp
8FePdIYUebf2CbW9dQgPPswQXR7drCykM1cRsixJa15bcZia05BVreNkolO+Og8TMLDlOmUj5ggO
RfWBdsiXFsGMs/GCD8PV/+Ql5+u5u8uFsfqT57futh5jdtjeprxotQbqAmwvK15bkTaqG21ducZk
ZP7R3fqmcpv0t71G9BrphnZFnamT92infOF2OyXFqUQrL20sWVGG4kpFiA9QS28iGpuHGRwWEiL/
PeXxh6/UTFQL44XOY6+n6D1jS+TyKrW1SziSHuW9p9LQeEB8BdER8MvXXqUKTQA7Hkyvu6+lfMLJ
v/Clh5hr0347zIt6ttWbOiIotPKwYloQe/dRX5GqVdFOpDxOpmf3Vu9J0XcbYVXJkMO3+GItQ7ZV
Vu8yJzfXZhYjmnAgPqv2uGVJ5Y5SXI6fBm3/GARsGoSJkJvojMA4UDA0aiCHBfJGyKz0+S/9YlZu
JKIqW/w8aPdBVirttuXXMZM9pB5AaF0nLvP2BtnUDxhj8pnRboZ3xrRmOtzHph9U57Mmgxpn14AX
xOsPC8/GTVMGSanapLsd8Cw9ppGQszBFDESV7RJUidhBhlU91fnksC0p6D2A2/STf57AW+oJ3Nld
CwUuNLUkPXLxTlg1OohQIPkf+fprBv6uXYLxmVBWFKAmeu0dw8y7WDzpEE/kzddOprsQs87mrxN2
dr/DQ1oNkY313ChXPked1LVSxcIc8CQKOF3kcCPp/OMlV/s/ITAQ8t/MXT5mLqwc7fArtbA85boh
uFkaCISRagzLj4uah2XjZXkZx33rZmprZ9iNn58IwTVJ7u55sZbIrCyBWGokbGMYInYa4Zyy4DRJ
tWzgjUTW2hrtIL/8CVJ8HYmk00ll0BxxEsO8b4oSKb9NnBGRyeeCnHQ35ujOzjQgf8bmiBsHAR+r
pQIJ0JiBHw6lsHmMS1Y7iZuxsRcheXjflihCDZLb4kDsvHeTqDrRyjX9Ak7umzIEWV8ShNvC4VoQ
u4qJEb+sOocjEHdMSNMvVb4CFcPRBf5mlKs9GM74kE6PfWy7Pk+6A95jxPl4geWfTJBatfXmgsxo
9zRRYPKK2Wb+z3lus64y7BWoSNLQ3YxDaFeQ7E5rqRIM9ziK9n5UfFJbwb6QAVRZmxWzCEnTWLtE
iX4mOJUbln/ym05NjHOejQKOekDxx+JtwO8NoWYWQZvtMUEYvoKhc3gdt9e5fAaUhL28DieVZ6Jj
d2SeiIKGX4NS/maS5zSKomRhdRc7DDdH05Ls8g72d66B9DmbtbHEhe4BOv666hgfGca53zhPo6Ez
F/6I612zY/25KgHAKIEU8SXk0WhTKIg1u+cfYzrx16Ra1mvA9Ul6i20yHBzMurKVwOHcEdryLKlG
FEppUO5JoT5y98Im5R/D2c5keq3wILUYxU4FOubP2/v8EeJOFqzkgtJLlLCg0N5zLE8x1jBVVIVA
OE5hqbaTsErTexT05r3OguhQEgztiSy92XNR6JTjmWSqt0UTr8tOI7Ca/cjuGPOVYNqugYOXCs0U
3GQj9kyd7aSAYwVLlOPGIW7oe7kdAX/Tq/vO8Oo2eUTVrEZj+YCVV3af4lyd3KdIqKE6jN6xCq2/
EctdYdTahf9yrkvK/QGuS2JLFS5jA5yDeusrFRjoNmvG1WfOcQsSVpW/QcoTbztrUkpMhc0TIjgu
ffgqd9bqNPzHcxV/XWAg3FH+L5TNZQqY6a2SNjXI8TCTlGs+lghMkGFMIaE0Ue30Ycl8hmC0tIzV
Lf3aaL+9lzsOfs41PcUb9vJXhXe9zW/DErOtwnU7aDbyn0K8NxasX4O2uamtDSMp49ZOgwgSprJ8
JNh6+zrwJVf+nYot23ykUpdQYqFnQwE2e+L6gXSgHJuvWQJIMIHr46w8tzsN7MewnVPsXpWjvdnC
QADFsBVSIL6ILrBi9dP/AhAcARn3xDr0OVyDoRb8Hfv5i2Mjvo6FVxS58mfuKYgPrWq1+0QTk6o7
YUNLN8rSI6i7PJkVm7YawNFeWvyCqr4c/drQ0G/gx9a/LycEOVZ1efdHKia4YJxD/F9A3irsQwAh
A/QPz1UASI9ozh2Rdng0TnTsK95FGmioogwMJnzKFYAicXW/KBQIdSOQKTJ0KKFZFUzWXiinoDAe
onBYjKsIRGpgYmqPpCNmJCC6gc/YKmwt44IV7zWVaamqrqfxDtOUWWQURI0pLDa+NRc5qeF024hN
9xxLYq6I9pJFVhVEVoTjb+lOjhf/Url6mf9x5UWN4RFixKc5quGFQrr2VHdZTDNhsJaHgsMS1zc5
4mThpGHx27+W85e2jaJBmGUQDjU9L46VnqiQYj4WshASujJb4NrPSN2ItPJl4scHFj7sNVqALrw3
2JfPUOvwUXpvn9kXf1Prh2W783RpenjUMs9p9ZJ0tnPDvBI73fs26gzFBtPZs6zSwp0QOQ17VZat
oDANUW0uqRgGO/enDkKpFAzFnSarfd09IuZCj96YY9B/zaE7cjiJGFQlLj8twjUqF7mBln3QLYYe
nXNMIAEn9QXAkXPbq5a/Rd3Ma266VzANtL050SDFIKodsxoUlyVbKYso23p7JAMkNsikjqNwz9Xa
eZfm6DgYOMPKsHhuhiyLMxJBF+V7sp8BUQS2/9oF4kmn8nB05Wvh3JFDJrd9Ow0w6JTomrso9k1H
jmBkzRO2PHX6PnpJ2E0cTMtoVCX9kAHCJZDlrJui8YSBoEohy42yh2rQaW6DzOqu7J2ZpP7MTH0Z
xrMoCtnGAI1jYRBAOzkiplBPukwauphpauoU6gmJSyYg8L6UQzkMDVyh2kg0CusfpXCeqTS5nkfE
+kkrXfe6tqB8z5O1khy6qt98RJwZDN9/dHKoeW+SKaHj0ZOixjYQu+23YIBSB/s/gqR3o5r/SkhW
XcUgDEciFbziga6lQMFSqtOxIzLK99ZF0GIPSyKKw3Qq27tWuBA4vJeYl1Fp/t+N92iom/fxPa6M
TGar4lubpaMMsZwO4XuG7IN3g3P+4EgQ2i5duQxleKRso1Ek8k9IQo8+HvikYlmNuhAErJtag1n+
00E+qWsytas+gq0l7sUxp071mDOa7bmPKGtq79fCjeaMDF3if0P2/zWIy7ax9n0O2Wt26A/7YonB
k0AmcM35qTA/yNBRK8uCPONj6SPvVaQIzrhtUG994GrKkr70nsub4vfWqXKxKQNHRrMRbuh6vKqR
uOd/nlKVT+UzqLg3Fs6Stumjh+A2asDvJ2ZwHH0Vko1pFQWJo7PZQ1dGzIL/hJYp/aE69gh0eXCT
meuSLc2LEwRgRKMmeqATSP4XVO60KGDQayga2JJJFyKs4tNybETETb5Y/yiBpzDQ/aWWUGdqXq55
OLtsO93raKkn4eH14gM4le8OHHXDXSlpsTKlOxsP/GAJsHlaRAQN+zA0sayw39Gu6g8582bILtIR
aFN1iHv4AXC0bXWNRlh6pIeJUqpK/5num1eN1DwEEorIXNqtnuRahFBGPsgN/ccDwvpF0aI2jV9D
WmSJmwg6I3A4Z6zzHIOUzPNj4yUuKfyrbGKMI0mG6gIya8gX9DcVHW5biyv60V4NGrKjDW+O9x98
wQ5qXLnLhlsm4Wng/2z+ZzyYM39IHg4ZAunPj1aES4s6VCi59z67Uoi9tGwGMpTncYcpRsYAFLca
QQv43axzdffck8MFJl+RW9uUA3riBXxEWHnb59ilOfWSNjAIJMqy0fb7mTAAgBzDpUanAGNEE+gO
BHksAw6M6LZS5nlihBN5+38e5Xv6/zWOYP18nKoctzle7xU+zu4CXoye3ZEPvNdCFbjH1EZiN5Cf
dCjx+pTvStNur/J1VQwW+tvpkp03rF2R4a6BCgOAAEfskPUsUPcO+78j3pJvspaBGt3Q+gzn8Arb
NYpQCC0q+2RhfDTNf2pRKlHC+5wd8xX+hnr01rANalzx00GmAISZ3ikRhqrbQhUicMDCJJ7Ufqma
3uS5CBMaHeFkNo8M84s5ZgH/BoMrd+UnmcY8PRmuY7mMgDeb05tzfNDZLngiypLjL/t+i671W8+S
NJErlO3Y/RPozIubODjSzRiAZ3f1cqxGTUoO+i4PEN9odD68nNsPsY3UhE18Y5KyCAgantOqaPM/
JAtErfmWMURFFnkaHEdeBd9KQMJz1NG5KFmLbB66uEc3nnWPN1pFnaodZPslJHH/wtH1UKXOHKjg
6ZO17RrXNDdwTwQIIJb06sO/hXlBfBXEvbkcKBgF1JOlNHELcw1a3pf1BDDwLQiTxwgKjXov9vby
Y6sepC1CqG1rWhV1TAQDgzgXqh6UFs4JVz/spVJ9bI77rBPWYbUSvJZwSF6tBr1XX0OeV+zmz3Dh
5FPX8U/wyvpIamyQprxTpjT+PvMiTauBiODpRSURO1SDxJuq4ePxOHBJhUDTbZ1NozYwBmsrg70V
nGwJI3NKpeLAuRqxu2ZNPNig0Vk2vsX0eipvzGLINnbvR/PF/SysFyZTGrU3EU1JH4WkaEu6Ye/7
JZ1kbYhiV+mNqsPG+1TYGQ0jHtd7chpTSlglwZsDIougeNRb/Cv4QnSx2JiBRd2OzFjzIkWiNXau
HWUVaCcsr90lkmbCTF/eWBysHWpdoJqOBzNqtFcdGxkqpGwXxY3e12bSkESDLdgv0ObgDboxX8WN
OoDfQ+fCuOw+xjIl1JLJ1wRib2uFy02tcw8gxgjzZ+7v5GOyQaYySYnzNSShl4IbFam1QeG1BFlf
4a265s2oBiyyhhXtaplLTnhHgs9UV76eB+Shs8EJ+qmDhwBUdOFafgr5qdr8DJrblKwYkA/mKzr7
PVRBSiiDTD9IuvXRgeqXzB0e3sW+fX3VRwD5uSpvRrd516jr1P4sWw8hxQd2ty7FEuTuD7vPJjD1
yKoK/OfrD8WazFAwYNJNznnWF579Cx0jZragKeWZHrcehjT90+i+Vr5j7XCwlUf5ui3jHbAF3rug
K16jOeJq/mDWZvYXCno8astlpSj6n7TGY2AdXlO1406FXwmPTnL1ZwRWYJq/snBhn08D2kfPgvy9
pbNNdgNa2q2cbC+CJcgv7WXwxYS6DYtZDsOFThd1pkHGruBCbwK6aeaa1ARtmJOCTmrY8koXDUhx
qIlTcu3eX1XZTKk8zmoYVA0sgoJHJWXQe3GHp1MnL0HJLwqOxT4TfYqVD5QBVMgh3t+pUN/Ysnv3
lECT16W6oHLhe1jlQFbNDC3dtmloO0SIkNCGrVxxz394qVCmCt8ueFRtgDdqHJZvOQjJSbRhIkKu
HvL5XhBImHy1uMsNQbvzDp898zqbgAZ+wIK2aqpZG1xyWKBXw+/VxqXok73P915JvUvzDPEppVjq
9JLXDbvFQij89mtAhSaJilE+7pmzBhPRxHIAaPB6u14EmUWvA9ruuCYg2Ukbg9j1CzPqRHfTIoMw
EaxCdRkGmXmND25UiekkiQlKuHEs/xZBKZp24O7JibtezrkJYxtyBpEWVVz7xYEOPC8pgvWgeOAd
S9e3f6Px59spqb9yFZIA4bnV/CihmCZFG1CTc0nLoJZwhxOnmTeH9MhbBvjHF4qtntDZFaOjTXb6
USqwA0wu65UYmc6D79/9temfdHQC6hTsDCdTAai+r8w6HSqN5MuWBzf3V3WbTKQ6UVL5bk6bnb5v
IFZZKDOHyF3okRQTgccFrPPeYZJBZcVpS+yVjuf3pch9TGvGXbsHVdDttAM9Xl9VS7wOzEaHVPIv
yH86YcK0NGNqVQUE3s+BpGL72rObBoN5RFKm41iJ5K4Pg9d5mpkEa9+XoUKMa6xAHm1v7fwgZeP5
5tmxXuw++58ts2Oe5A92vtQpfsGUsrDc3ioqYXAd9+EqxFVZPmDkEFgaHPguDnU/Klm/VsTZEf+x
4jwIFrS8z0BHFwhxdQ0C/xcjVUxgme3y9W5El2V+5V748Z4SlB3hzqghqkYS3T78cViZw4Ati+Pg
IkKg2d5JjEHen0REgj+ZnDTGvh9VWYdeb6IAHp1xrxYS+1PbtdclsoRviHkI99jTRDz17OL0vGTy
cNXrYsCvSZhe7Fzlzk88pRC4yKm7LHwAFvsJjVcbfM5TF9wMof0rBlXhMz6hUL5UHSgytWShoDff
gr2trVaWKVYyiCWn24v7spZKuJA8f5oQwvnGlXRRBOztgYQJLpqz+L2GYBMQMUGhz8jmdL1YIpJp
zv38e1LaKCVr5yjwmQyG5KM/MrNDloiHC2NZ2mMBfnO9vgeiQe1M4Qs98Ksa8lCrq3pbx+UODe+C
Xonv69eWSu/S9QFOHaptYTGzkicrCOmL+KEQMYcV2TTNf9fe583fQnjrl45PuKH3tpKxECiB6mg/
+Qx6px+hR8sP5xnj33WeYHsGJBVZzbkJNvCeC5rDRrFB62IRqnCl8jknYP8m5l7PyvRVPd5SsJXu
I+SwaKPpXXxbX5BIA5qhwMC80fDnRIQvG3uTBF/veCuzDKDT4Id785R5V+f/WuTazdZokhQ0M/Gj
QLCB8w9BlxwVAlyvuCvqywmv3cl7IBHePQ1q8TdXlaBWctrRa23X/FyRuqcEvUFE4qsuUbErcO6x
mMyXUW7vonjHJ8F3ou2BVT6BtOC+ZBmbQjtLkBsNAU8nR6W+TeXwMRbhq4g0aCYWAaSKGo7j37jh
GM0vOQ1GqOIm+gCfa8PU+/jMMhQaD1qC0Vp2VNXQeePvZhDSvr9YXEfRdJHdI9CqWewB6dVF3IAv
z/Qp3/17PBEioaVLy9YHApwny19d46Rkl/2ll5feaQbkrhSZ3mAcWCqtQ/2riyJS7szM3tbxJQCS
D7UCoXOvsx9b/EGXVvfOviJLQfxYiusgFrhag7znNgzpFIOPt44rGJsktWgIP1jpszmwXpYbbCil
GraoI9Nir25RolCSKV4JnQoXTEHa9wuAO7YTZW12Bgj1QuOsRjFF38R44Sb5l1nLfNDGbc93ygLk
SjqRiNdyE4Astu4XBXBvBcKddw1z+G3nQFK9pi9hr09U4T8SQs1ryKDH8hUMaxW6MnWj0xbrG3iH
3WfpTXphOlmDc+jp61EQ7TdvcQnmKiOMbDTTNlZSW7HmeLahOtb0zRk6N/FDdoHmPMRSehpNFBS3
W2O/D73QjAmRKb76W5rhPTPRz4nOV30KqDibIOEV8Mf88zwF0YsfDg9PfDngmSxSdqi9loNzwvQx
KqZIJDMQqwFvipX7V29TUg09eP6FupQDy0trRPQK9ZznSX1qIfBRByiKgIRnEuhdhfrdYJQ2yC1x
6++ZbM8J9oso84/tX9B1K4tcVPrZiF1Kgl54DIpWI83VolhkSmw+Ma94kumK6Ngq+exGxGoMY1uV
RIc47DgQVgInaMzMSKP7wdN0ep75xHa/sR1PFjhTUUcpC+Td/hrRP+eQh/q6z4Kpq2p0ADJlONWB
RnV7YxubDcX2A1JmkOxa5pf33Gk2B99F2puKRJkc1jMXf1omf0ahRzKbVXtzGvGY236qMKkuzudT
VWpsMsHLdS1dxMr3ZPS4nyAVA38duc5da8Hy2T1Lq0SLxBOdFBcqW7psDtUDMqdaW+vKW8fTRHQk
RMtE2ZhHENCP1sd7RGDVZPFNcPFoJm/xp9ehqgE+LfUsqpM1Ls+PuINY+Ne8hp3Vk4CtSfk2Gb7s
csjgqPplqa0VSrTkg9P5eE4i4tsSKT4K0ubzEKTJa+WsAQlQ3R/iP4jKElNOXaqkPrQOwef79Why
FQRJTZeZv2KqR+ZUJgdaPYm92jSFpORmsRQruMY222SaR8GijWU7ryzu8yJdwZly2Ko4OTky1YNA
dFtRiBiFnjKkAyC0pJ0JvrKFHgR+knce4GDk9O6lEXCdR2w7Twxx+3QT5LH8k1aQwXXq//Rwb9sf
xNHyp3FtbRGCkFhgqpQpRn6G5YBLG/y2CNEGvtetd+3eM8ofy+zpVqHHnJHOol8BFNf9Xxcw/xh1
GHml0teid0HM1GWCkhvO4p6mT7aMp7h8CmZF3U04gVBV+AV9Ak+3wlWCp5JMMMnbrtSPYBewI9DH
qdJe8h9zeIZxp8K8Ufx+x+N4Mov+TrX+mrYnI/Uv6BDGnL3+462yNvah4FHOvG09cpsmJThrsGSm
q7HFWqq5bIPlyenar/EP27GXVv2x/aCeeQfj5BQSfak7CuXeRAw36xEco8yAB3RC5cKzwepD+K9B
MrX10uZ0nBBFdqX9r9NGXNobSkpYoAvwW0CaeGMnW7oCsyqvZFwkdW5asLcJ51l4yCPpIYfLRG0U
xoEaAVkDm47TmdZ7kuIHcssSTjv1syWzfRUhJrhe6YmZtEuOfjisltJTd8cym1TCB4X1uUecF681
qgW89OWO2DWIJjn03PjGQ5r2eKlQFyT+sqN23mjrWJS2Il577MM2k1elG78648xcjUBbiQTCXIGQ
Uewxi1lJ/ZTHS+C3eqXnPRhkEkYl//Wd/qNASgC7FTVTTof467I8+btO0g5MJea7NfAVUOm2YfSP
tEEzSr7ZlQm7DZrwF/On+h4L8rjBr4VMzeMre9uFPhrl7hYlbx+ijd0TTwv6KFyOuhWt4Qqc6N6L
wmLAuqyoIUmPcDGjdjVR2HNrI322/fs7l5i92mn4WjQqbRbZ+aqn4uYeRkQeqvJXNehB0BXRPC4a
Bq/6WmGGmBDsgil4r9a2IT9OBcyY96sDTjHdvySBsR8QOT/oEu8tCW5zsUgavUYu72WZxK4I7M8Y
sGjSnaPHyjJygh828FtjyCw+cHc3eFX6eckhXvYnienhezWQFLPcOyDrIM5t5Zs7wub8dnfN+eMF
pDPRoClm1r5EiC25MumhKoDJU23LL16Ci9vHUGAh3gOSKwFmKvjAkFcF4HnC1AhjyLgOXD4CqdzC
kSpEc5BKMsVNn4jDAx0ZwsbeZRpkZuxpY2bK0MkNjYQcQAsxF2OeiQhSbDFayH97dEbONsX0SWfe
D9iKAj1goWqEwgo3RDCKDNTvmcWgX388RJj7S+CKZZJM2K5dA5V4J5XSxZ8csl1vJSXh6VQVTM3A
TjSZw28SJjOoBiklNUzFOU+C+ADR9nW7qcA0I+Rle+PTCm3gk1upMY48RJW3WV6vfL8W4yyzFOo7
AfyxeuIDT8D8A9ggHhNfV2yZHgefODI2NP8Q/mKkPKBhn1VlTS7dAgSt3XC688tzPTTPh3tco8oe
tjYbu+Tg1U4TAOIo7O+tDe+5hdACk+2Ln6hzhJpRja6ooGr5g8aXMrBB3fGBmbLas6AkS2mRiFV+
QQ9SI+Nq1dJxgQkvhhDmCIHYQcSkYLoIPg78dh5Bqh7IxjelomeuLu8TxBYQLrwjQueuPHkflrIc
HTUlzQpD+YNH05y/5TZLwDq2733E6dMr2ZSWFRJsTZkUD9YLdCv79yFOz+oQpCGjOvky936bxeIu
XT2cVKpSnUDJYX55FLaAtFjvEd1KLQ55a0HKcee9l3aXCbTyaxUCuC1f1i6+JgPKvUC7Sok+Z7Fk
DMNP+Vn9LFk2sMlliLcQ1GGzTvDM+ADxmVCD0MyFQPPyuSulaypfdTVSAzusA/A9GrqLSiHh5yvt
bObwFBh8oiK9zekP7U71WIHvoD1+v8OnpUu13Ef6J837ckTHHMN+zrZuVdTnaVKA7w7L8jeM13pG
IYLmR3n4z6sLmh5QRpWA/3uRle7z5KXcjB2xrd1GukwB5FM4kxlpOerUfR3nJ3S29pzzYaCKGk+r
FiNoMFlk4iBRdgQMSq5Q/ux/UmFmkQPUVg9MiCPglEzGQJE47WKIgYKzZqVHVJ9Gnwp/eNwUzw+Q
o/Zljf1Iupgz819SzPbcbcbXEvmrjXrIyj/znX7Q37h2pcD2IQNowwkW3FgmJN7X/d07ewsDWwTr
fyROhFU60KN1/LUQD/6SHRp5+dLXoV03XHAnoXAsfKhCU5IweC41/wXkQMMRK80P/8hEwKgvloCt
hTfsF8EbBmsw75VyHMY//bMiJofiwnwu0OTNJvYSDwalofIdzqtCsW2VWacZCrKrwrS0Acc3QBX4
xAyDYImobgvoydwN9Tfu5Xt69FpnItycOy3nxPFs+5VV0xv93ToTv+dYNIInpP5rw5gu/yNCf8Pj
OISiXxlWP1iaWdwyyzY1mfEORBO7JOX8mK7ouIGZ909k5jwH9jayzxYToFwGPbBQ+yo5j+kmhVWp
RB81Ousi8S0CWZDszncBq5ZIDXHH6mkstX9WCNTdT6iZ/opCn5jbF06b8eorVeHG7ahVvL5+AkKr
pRqYsiuSM40VoJywbV+DT1Q+Oh+owyMn8L7spwXzu/4aBuXMuF/N0IVDQxikmaym8t/FVMhvIJxe
xDlw9bSlx9bIE6WFlp+5ZofRmoPZkc02Ks2OIpYSRDTP0vWMESEYehtxXaflLOIRYRJWTzJRFSfu
MbZ0ga/MmWXpytv5P35b3Q1vrtRLWuWLa0r5NxRq3pFRqb0DoCiGbDfv0qw3ix4illXHJkOd6vfl
gSe/bRP3fjapbtsL10A4KeUN6Ql7WrKuQ/yuuxWTjuc0pZ8VimTNh5fEkJDSNdlzr5NaOQHtV+Nk
z7ltoqpjXZtqeOfbVBBTZshysN9mjedW0XScQpuponhDlk2hHZECUYJQAmP3D8KcSMAK2U7TcT+g
SbZPxKbvYtCOLoXYbZEy0heqy0QiHBldtuULwVui03BKeHTgP562DTGqkegHfg2VoFY9NIviR7MM
ORVvpRKwdXnJ5fNUuzRmPIfVO97vgEiFdnxgxqO7K6x7w+frrtcH5WEnEAmSxZ72xK8qVqTcw0nr
SAfro8DPg5WbyTK0eEcCq1RFyxi2t2YxIlh7AKwt5N1PZzgFqlvVv4QjXWgkVUwqM2pj2aW64Lfx
ZccGjsTytCztn1Wu1TWqb7QFO2XwJqbz3DXsE43Gb94fHDjwsKlm00hHxFqzn9FpA/SQZQGarfpt
6PMe23UDbMZNRjNeqQFpYjuqv15S2mp3stSUzDd0XssQA7seSEt7fsWUJamNa9L03qRRJfcGTvfV
J143xBNFNztdsRNhpJTWW3ttenYXdLJ9HdFc0oRYEg5atzPycbSw17mRE63m8zlqL9QlEQzwhkVp
CGdkwK3p5TlXWz8OC7PXMLCOlVvadka7xILU588nBBNWnStHTzOhiQSdYW4cDgdC9kgrFxC6mcS0
wmXHPvG2QCZuQ0+7E1eL2kFJCsXyEGCVMjYkz0J1ITlyk8I3YX50ySS2wVXR7g8d8nhqK9vPM/Y6
dZkDrscDXEDO775HSPnB9G5r526NnRDwzk9pNUom6+yAjwqm1ktgYv/3fhTtqC6wsCKEuHFHPOA5
mRdJbXeUqYEsbqqLRCh2chPD2ZA9Ob1O0WuW283XoTC1c8KxPDU80pHKESz0tzTCu8Ba4tkzZWso
u1fdIP4pY2C+RfwgNgWvMRWevG/irlpeieqH62NoXS7lsUv0u30l0nutSIYXwDaLkVRymtrxIUJK
7oc/Psu+EWavDrmYvvzR1oYfL9sJoPU7fQFiy1GobkD0DNx6Zx0AcyDsCuzBP+ULIx9DqvzGVLoK
Ech4sTBGgAkzHeJ91z0REv8FJueRiWEaE5NcCy6hhaCiiZ7oiTNLP2eJex5fxrm4XqHxy+TuPx5+
DdvqF0Mcp+V0jI5XPvKhZJUE5ovOVPkK9895idmd09J/Rj/XwnFNLu+//4aMU7si+gQL3GUfJwpJ
qtbaDLjsuIrKXmC3EPWu51BZNM3A7/EY0kz9VR151BklfDUeBx558DmELy0RVvuSk3eRvhhZA1dQ
aCeGSEBr2+yWSs+EefEpLK7pJ4b0MxCc/JCO8vP6oXb9bpUkwEdoWLoKDTZKw5NmxNVGlmmw1orU
sk0wGq05obqCxRyJr5A2Inyh1jfpbIR0z5fYUpt+EOsDkejlDZIur/f0YsSP3lyrtUoQS78PcPgO
0LMG8/9Ex0Ck5Dt+y/Ao51zUPqRlhF+8tW4InAWmINl7rEQoatIh8yfcdoKdRS+eu/bANOo+HBgY
kLy/G0JpPSJXJ19nQtAIy1DaPDz2YKnjfwC9loXEzp088eurDgjo+Tsm4XZoE71Y1mgKfsoTxHIa
DWS5Ulnq86fwe9WjRrXw1Qpet8g5livn+9WA7mbDu+bK4VKwLeJyDPhrXxaFVVXzdfocNOKKh3bB
qgPpqnJoqj3PV7drrN0veTZz5yz5B5jnEPu4VGrFazJ+TnzjpzHqP/u3Furm6EOyWt80zhQNsWX2
Z+YP4x96id/d81urVbTVZ2e7ble95Cr5GIJ9ECy3mJ5bPYAoVsYPf5/c/RdvuNf2QubJIXPUG+as
79curmKBD3vpVIlbcs235Eo7fK9UszrQ5YuAQtDGbj6Rl90UP5TtodGlHhluB1cGIWl7aQmrOe7g
4+7FIM+ogZmMum8Q4jTDO9ffQBuiVhvG97hVTUafx3XFh2H4tPlHycT8Yq9T/J5PVAa8gXXmTeEl
9zCAFXVQqJNkqh1Yu0Fjek7/H9N/8IenfvyvB7UEKcS7+JuIylGtnoiLWBwAsW6LIRvM3RJzrkGJ
f8KecNKOEhts/sha6/XKj9qoNFcPl9szhNtaHyb+DrldGU86mw6P6GGD9PZ/hQ/KiMBeY7SEkJvg
/siHvbwpgdhubKiMeP4M0bQNz+PmuU7DFRipM13mT0q4qG1Lne8wrbNHSjxeFn1MfOAbPdjcUTIg
6GxUHVb1aCd7j5wvx/Vva8he5VJ9+y4I3F6O6/iCrtaMw1PY6eClYERBcpxoC+WLo8VmrK6s3HUD
nrG7rA2OivzCdV/VCsNGIGt9HO9lm25LHQifUe3dT91WFepSUrQSNC+VXJH7JIQcq/UQODuShbzA
6usE8pqOWw98I0eAN07Fa1ijQsZq3/jSVbGTyiAh0e05/g2UNJFE8gv8wvq6JVV50y5iqm/AQ+Xi
+zPXtMziF8jd54Xx0srNpkP5ArqZpy3zsG2A3WiYbjm4PDy7lujIBGJ5lnr8E9GSaINXXMGnBHNQ
sc+YGyy2nyyGLU+2DzDNB4wfqt+YHHnwjEAQ97g8rHWq/Zd5G4trZOXRQa0p0akOocnGrPBMGBxR
JDKyrWd4ImUZs/RIydL2wV29UlW1yDk/4cnpKU+ltv2YiJ+87LBadf9hb33gyBsDCrjewy5myDaV
XsXgPRFn3btMSIWwH3OFTN+GrqkhZCUCtn9ZW1MQcgxobPipBIjr7PZTz1wDVnWTnucBhiNv5h4C
vnKSdwjYYbWJGWrszEERf+8PbSGaU447cIOgIyeYzL6xAXk1abGaVrwaSUIoGklvOqDqSvrNliqZ
m4DvCCUyhkf5ENZwCa6D2g2FC1Se56E12l72tu5HJLLdIMFJqEa/9vrzX7FU1VDKfDkMee4PO3ZQ
53LfxdS5RN3b4r11fg+1jK2DX9G25wwmseZSJ0W5Rd8RhwrvORCudyBiOOlWVaylUv3E9aupFC89
QwIIS9F7C9rrT23/UPToDqeK2h2Ot0DEnJdfU6VJ9IWMt0g3878DF/C7EUPi6t7xg4IHCZsvXzDq
MbFINHVHeOif56Q2hGOY5Glcbpac8TCDJXEgZhpeSb01DZlz+015UobdzCJC62verDKMt4xEUor/
NTegd2+u8rMt5Ye1wWRwT1LMn1ijz3dtHMYH4QSSDeR4HqOgfnlXsgFYopITpMSeNhQffX9n0L09
71EFAm7BriHrsqKI0byGczaIuSO/z7/TSbT1llXVnFt7zYiNiR2BPDXgF/fttANsZSICPwGOI/7y
aIr8eb3Xscc9aVc20HQuix7FA4gHramS+NRxsD03je0hoVsKNz4jZo78cZllUBmMsVV7KMS1SACN
po7IB9GHa9VR+m/NNTAZcnct0D7fXaUu48mNKO/O7Rzb45NBCoomjCC0zhvE7qKrRBxPqIE66twf
jrsMHJq6ayKeXO35+9goWPCoBSAM18YyDpFw2nRL7axMApMSQnlJrSE3sbIpwtamIv7CH1VWSPQX
iPBx5s8x5cbSkhx0fJ96uhisbCpybY/XC1jra2JtHAjUERFVfXOf5SE0dgGAYT1eAJzpvMUZbzlD
318ZENLTAijld01UwCoLX2SOMcvkooIQbcLOLTKQcsEZHIiStG8AO6sYb0GSQnnaZpTWzdQjvhQn
sMQP1CvwvA/XjqspqVhzLxUToCS29F0hdAunH3NtT1V+KRjUyLQgw7pEi3W6wSJe4p73SlBdRmBZ
EbqUP8Bs7yx3lTqb/SUxZ34R5uq0fW63BilrsUjljhJrtXrkJlzVihcSNDzL78zxawaq2uRPNKhR
kD/B3o7HnuCG6gMkfRy00TYI0lWteHAIvRPRhKC5HTtVVD6Safe7ULqdYk5h9739JM0o+1IyzQzJ
na6El4OkIgWpE9JkIVMXHkJQqFjBnfPitK3dlxQT5PJPLPtQ5EGnz7E0FVjuIuhKwjzWo/rN40Yv
hKIs/Llfc9KDe8f5qMTbeehZeCBNIAPIioFETLIIH0rfeGm0FBfYRSswrcD85hdpfL/RMYjucobD
kz5yMGsnT+0YLaQzS9dcSqnti3/0L5eLQwVJbhbr6W6ymrw3+XTTpq/db2yBSweie0SmYM+GgoEG
CqYoplCv2bFCE3UlhAtNSOpYyulMLqKTUbECWlWjf/gnvJ1KjqluJibbdcp4OPe9EdKjqMZtIwSx
E+321ZAYLfXhL6yLMrdBh2IdNHArR1J+vWNQCkoJ7C/6RkCvIH8IKpwRhFskWa3CCWzLtlmOOFzM
oPdABGrNgS0qG5GI55p/UUknzSU816URiJuu8aPzWmKfqetCx5szU27a8PMtB5y4wrKON7XNvJGN
is6tDNoovQimVNagNK5JAHkcbCmh86IZMoXM89fnf6FYnjG74bY2T42VAfidefNSPveYCOesNhu7
nYe454i9o63rC2b37yr4/bj9HxQnL+Nh7FMi6a7l3c+ivm8zZH2OHKit2mmyrq4yuBpeAXKNUfBu
yWqVZ8DXi9iUQNEzbh5khuPBnaZNhn9+rme5Yq3PFwfOsXo17wfrVkpkrtUPIt0MRSBDeR9EgFHC
BW+UjoLJUnJ3+lIk70wGgi1Cu07cfF4UdQamS+D8aYCDyj8nZqe25oHFnLASgS52a9pTQ8eDsDbM
8b2mnodRJSpwRClXXDd0w2GbKukhoaL1XW8KHDglbP3j4uT8TZY2z37FJUH6Zug2F942VaFAVcbq
aIv/ROp2u89oNAHp2aE8pEvSSkkr/gP7igFKrGcaE2legr9V4Hht6uVlA9rRiw68eYkcFvZB9iOD
bq++1CYOi2In58mc9gya27T7rbmVDNFOPkbmyXIt1Nt3z+Bm9UUFwIM2hukEpwza+jgqVfOBcT+Q
FjN2MxoZ1+vjvP/hUV3seLMxDPIeLLirkUwXuALasEb/A2sStH0IDWFrtGgzZNJtcNjPji7p1YZR
JRA7Kty8wLVa86kjc3EGCYq0PsvrRlE3D+7PWnlo09zhAsS1MG7EyhZQjuXgZQrq9OiAtB0cW1N+
YKxHLgT1G9dpC5H9BXTF6jWnC+jWstuF8254VXYulx94c+VQqEVzjXW8ttmzxrkdZjJ6hgy79UvS
KXXEtkulNnCnPkXD3xkbGONXzY1Trb2bkH27Bdkto0JgFHolGFU5dWokHpF8CND83pi32iG29zuf
UjBiRRM6AUlFQu3f8Fyyqm7mQ9mqw0U9K4hSDvPgUDvDHMXNhABITg5GXD36+ZFcB/j1bcsgzQpO
mKGVflmAmNJD4FoiDzSuBkL+b89he1DtBfyXC8oLWPDHD9qcsuZOEN9lX7o3CwYFeVQtrlP44/o3
CSS5BlOdR/TivB9BW6mZb1wBzjhR4aih3vJTSuBgc+VRJu65A63Fba473397nuBqrXBck3cbcZbr
gwaIPiPPoSponEZ2XW40QFDGegCWL2eTCipy1UoWuuKO3CBct3UhEarKnIVMThobmN8lxmgoLqwu
FvcV+1mx1+fsDSwz+uu28zsH93zZyJs4G1Wc4Baj+QOH6TK8hewMotiA474mb8K/OY5N5Qm3BwbJ
kWnvgkdVRzmmduJfFdwwv80iVhD6RVVyXkMAZtKI5mI+zAdkutfZNL0gijgvrP0w1y3ZnWBGl82l
q72DWy7bgQzNbIdlK3DKz4md6VHc72bzuTtYv8GKYVdocQLsGaJ4l04f9AdwnrjYo2qQWlC4mR7T
p86sjX2govbZLq30dUuxbxIZfpGR0A0VPjGHCgr2oEcVcv+KmCVBI60kwlkOl3RFTvYCNKxDlPD7
RxdbxhycfSqwXtR7PzfZORRW0QR93znoggVUgHO5/FXPxc4XYykF2meiJvrfWkD40LvoHeHcfea0
lSxR+/1z8BtGvGwuKoXwPnZVWs7vTikBtp0WzV8P09agkGmJlr+a21It8vrGZ6RpXU1m3SGpTjmn
Jg2MQCBQEB/rWv4bVFKoBkGXnhWtIUCcClmK69c6HivWO2XnSeviNyJor3n4/CGgHwL/VrXxSVME
nOqtsnTV5E5Wgs+3tAHRoxHghKwZy/ghQNjcSS04C+W56MWBfHEdofV7+p7JxMlDXY4O4f5O0Jb+
Lz4RQGENMcC3/PX8yWti0sHFb1TX4zYhnpScCvZYz3/HhdhwgnpTeoE20PkdzjrBONl8yBprutK3
VcYRdpBrAyfZes4UEX3VYKBIWesLUgnWNIWWvK1XL7LE7vMdK2dWyuhZLeLJ1xREK6CdSqYpon7O
MXLLODJw9SijLRhtK3ex6HGJpiAjGmDPSIKQwJFfyuFAW+ur3vEb//uEH8uYw3K6Uqk2+tvOjrii
llekfQZ0a3uaHAizVJdrX3LKs2Jm86T/ghrc+Z5TUVFjpnbCNRhX5tdkMNmcDcvScJTByNL0+xsS
7xxr1skqsiSzo0ES6sJpZOpq15xjRWjT42LQKYvvl89FRAs3xHrlhglUnMxzTc8G6Q96Z3oQcsZi
6mapefumRFzI9ncuTG5lIpe4AQskIKAllXIjKfAoD+MsL6FB+2w3274XwUaoR+m4qjjk1zbEm+FB
CmMDR6CpAsOnIBKsr42YLP5oe64PgPkc5jRimVM5vnb6IOUT/akSOKF1RB1MWK9VcNKcPyI+Z3Nm
ypw0E5dtobmKARKIskjVUmN6xO4DjFV9oZ8x4jekvtKuEx5Qt8PHqcBW4zQG253IR3xZbSfzEk0E
B9uaFlqZb9N8E7cCTU3G8wYnL5x1v6KsHLwuEtjWX9AUohphsUPjxkG9YgG3a9uaRmy1dNghbWRl
5VZEFzoey+LuLD26n0EOWHIRYNvdaDsqzYiUzlNy/49ZNFeopE74dRrW5hpHg0JyFsceKvISAiIW
rKXXj8GphXlVXAwFchqn+uauVBQ6d71LrtouPRZvNTiUB2PhMxcYcAAc1PUihavAiC5EVhQIPmqb
XpmcLbGiPRyngX7zK/DwwPc+A0ZFNirWktKiuaHlg/RfYbmpBG/a+6HUfXQmuY5tthds14iB/CPq
vrqZGduwCdhCDSeF+ZrvfnlLOO5JfsLc8lrAZzI1ZB1jc9y72YACSu/33P/PY1w8QmNmEK8u60b+
dEyUiE0aMr+UESuMuDLcb6P2NuFUt4c3ez4pdBPxU1DHkPvRpzlTfIlkYojmESG/vT1ROtQyxJom
JlY3KHRWChGNNh4msys5FTWc/LHculiiF15SRI5M9JUPdZTKCEV1DagLZNAPlmptqdc+tGhtIj0q
CvVTG8DMftxzxMN2yW1+IuHkd8CVnpRcnHr0kA2JcYwZK2xvItPg39UBQ2I/IJSLgJSS7Wi8NCzv
OlWeTgyU6G/zULXB3fghPungOcd2Yytiy9R2uqaf9XzTjN6VewGY2iOn4v5ytt01gZtZZxka5Fmv
vNbAT/yLgcTpehFf7dO3P+Hdc9OY6iUh2PsWCmd1PT6l9FBFN/Kk6ZRcpRTj7lNQmb5bvli8PZG0
7ldtIRLYZYzxazvvbcnTOOmmzoyyWxDbnjbm+Wba+7jl1ho5qWwKJVv59iHGTxePCfHJVFoDFcQT
dK5LHO3pdAmrCc8MEWMlUSeakhqnTSbB1u7Meank+I9E59WIeORiGyyo2m9Q3hXBEfM7ndlZp5YB
w/VS77mT7Uji7JtagUIt2dtHpiKfbivaD6ifLwJVbK3Bp8lALPT2L13ODNEWgnvcRVGwWTV/x3Ic
rbPMCLLIw2/MwOMiMJqd2UGWTS1sFw8RyrAAZzi7orRteEICOjNMtIS4SUvGYyq13nTsl6uWxVVI
a7ZU6A8ywxOhdVTusblxK9sitSNDZVbYDnqV7DoRhM0sxZkSSNiKSaLA0PH/g6GDvwABMPgK3lv5
NtsZEDJvBbSIsLLXsAD478whacGcsr0/mhsxqwKjlk4EUoWGvJMNA9NdBMj4N7opc7AccUxn3zHP
YN5l7DxfZ0WeeceL/g1Rm2QLqxCiTVGfnKq+pGP/7xOyWPQNcKn7j152yruPBVe79i/Q62nb6u23
VXHuqDXDnHxqQ+A2Pu/mHTeKivzenBI7garj8z8jqaHxPlpDmgQr43/dUee0Wv766e2KpTzbMZz/
xj7v5pAZ7gNrOob6oTB4x7qHGqvoqvfwgHlpODbchu04ZSujdjDwRw8NpiAuoW1v57HSJaYafdw4
KA6qvoWjToigCz3R+rWZC6RGjoU+jE+ecaADQ8LhADNc1m74ELLZBwLgUV4Vau2+g1kvL+Oz5/Jd
UeBUapii4cVlblfJvII19fk1ZlYJfL8sPU4UR+l9X97xRJHkvgkf6XEhh3zUyUaMi7tDkmBwc4hv
Au1BNf+7ijebt+/10QuOxGxWAW+Qu20hozsharrNY2Thr53BjBGnE6fqOjKxgqLwQ9nCFRw67N2K
J8ie+mJs1EJMDvpAfuGRApQTpsmPRvPzCgqkkm9vCx5knABGuMjHiEZVoGs7+oqQ9QRjX+wtpVxu
j1HjU6MFqxEhYH6mAP17SuwsHORy+Qezd9LH4kXF6JErN349pvq4hP5cJnMoJQvjY14uvgIwQIxO
mvfDJA9+cKt2BRXckcMdGYEkPKCTTAzFQfuel0SSRoLhg/hetsd32bcPGBdxDuJtiYhCPUIQt5Df
WyeuJpTwpCejoyJawtf/niDXf++oVhC9S5isiPeQdTOWFPd/SVVYM1TtlGHq2M5FkPt508XG63nh
9i6BLrcQc51QuLJuwuw319Pd8dC2aiD08tyl4iwJiEUUg2oSI9pGgrnXwVBSV0R1t5fFvKWhmrGP
r0cl9mBNeSLBN78IJWUV1ZgOqjiaIpzhjSRAl1CqVdy0ekB0fY7JooSo1gzmrxbM6CtczF6wDmp1
BVq99fkgSgBs0AJ9fCHGNboHU9h5xbZe1q1Ao4EfFRIi/342I3VRjYRkdc1NkxweBEPn0MPPPvdU
LqrL1YjYEOK1gFrQmbjo+6DiY+9GuWWFQeajABK54yUa9xlhdFo+wJHj+vptdvJUUY+8MVjPT+ek
Z4f0QTYuB5AE6L09f4A98+sx4kGFAPFz0e3ZGUCSn7td+47DDXc70MARuCukCHoE7LWo3ZvfBB+D
IL5KeTPdN8hwDduveev0WbtTxlcMvILyHrTM8E12grvKWiPai6+ttbODTT6aiwUb/wVeSdXGVeJV
fvHlh/ertp6/bWH/PtYBW1kIiYVsnRN0knIEPk4Yhio26zu/FXogkslZ7o5a7VuTdET5jSLnJah2
O0FDkMxMc+k60HfTClBj8l3XAuIwQRTefpQcelO8W+XglWtffuk5EtYAoPbbT5qqrv+L1IPbTp4N
SJ2AqQzabfxJ8X8P6rk20wvsF3JVey3Kh47fdXod1IODd+FchngNAzwJqzYA5CD9atUgqfBe4l8D
AzuO/W6NIMPq95C5Dxc+3qn5aNdoe1Q24QNJCoafNyuU8xErOl6Uy5beLpf6/HbheNfrrXlAerjJ
n+n3bPGEvXQayTDCKKR8EQUNkD4k3qNP0MM6qKhkvueVBZd09PKbY9FJ1t9KFxpAzlZmpXYsv4Hr
z5IWJFe65MM+qkmuI+EaZzYMVBMn7dOPLqgxuDgJNaJaW8ynPoCJcrU9129zh//5f77qEnwHXCBW
sglKr8Ncbj5cbOUlskPvjg8kd+k4Xxjeuq2y/daxJ0LMYInSY1Cxj3o0hDhmjafGAkyq2Dx/X+xy
7JzU6Qhvfxaycr0dIYwFXPxL+98yZFxCzTwhmNH5k7uipgK1mNjzBKJ+6JJX17UTvCG4Iha4yvkT
jA5Z4wA5FDLPAJXFdQPt6bnxVM5EWbkwpBLP2QZSpNrL0amRLALa95G8TOsQn1X2jpTeygdEIH+f
ubxtLLr+62HMG5VRpcuINvKgGK2VPatZPjNUVBCLFEEwSntR0Li2scFodrKxvQwjwrmPoOXKmzDn
SMA44N2kDb2qt7ZSxj5T4CQnrOnLXu7EMRNDhYRY/02le+XVWwnBVTL5QR8wR1mM/KYFP+5PQDiK
C1z8SwJIfCOg4pXGGBLyOqDN6g+Zao9pPRPSH8wxiGknMNtu50v3RytEDC3jBMd6GVcCqAgRe1nK
JNlOsuWfiWE4Pz0Bqc77nvIV/GDx88zUnKahj5Wogs9xFkldWDHCRVWdPItUV09MzpucpHRJG0oy
D4t3+CEa+0Q6Vc0xhlGnPx3q2GcxUnKRokSNkBRp9LUN81XhYtF2bTVNN8WWPuj3Ybtsnf+G3IkO
xmvKTBMF3VEWFPMeZpNBdCatRUTlQ4a7u8Q6d5nfl3e1wzd72/3fRltRQzogi0jJXAK1WEqCOiio
2nev19N0aAF/oNrwf5dL4ibQ171pscaM6QktsD9tfJETl0HsALE17ETIhlvPViu+fx6h2zHMIQZ7
ly8/A5jHGMYs/ps4m/s+bFGgvzGahbJXOEYyBJtwFNR67f/4HKZxNd58Zm9N8/thsXpRx7WS0Bij
ogman5Sa9TkE1Y1HpF/5EBisTCXLUvHeV2yrLi4HCrRum882hkgwshgzY8Nt36wdpGWUMUjxonep
oNGq9hQUCYg47g7yIqZcjz6Es1g4HDvVcfPLjXZEpkVReCSqcmOdd/nqBGoluKpBPh50tLEIjb2S
QEVSymsvLggPmw7TLQ33QQpbZmkl+RVxlKScf23Z6AutiiEUd5YJinAPAiKXSmVWbGjiVloSgtNI
WxqUvaw9o8nkeOq4y4mcXY0E27CTMWqw2iKuFWGXUoxG6GX/Awg8h4hZi/OmoFzpjzPsmXJlmoL/
KwPeby6Q2pqRRhwTNXNeLCOXNK5Ezwylsnkwfzw/PK/0GCXdLi+oKLa8A0Uvmc4CB2CCwYJYBcKr
jWK8DjbA8eDUG4TBPAwHLT6hCv7RnMp2ObgOR8Xo7fs+9OEY4Hk9GntjpdAulyFhbnDQobQZ41+/
6WECMfL6WtQtrcZDUV4KChdkce7pD9fVHAJX7LlvpObaubWQinuxJ92/SeTU33KQTrZHvE1J0sIo
9Nzd7Qxd+LJYFiT29KeWBkY0wGtpJjLVm8MEbxFgpD8W9M3aXmgsS1LRhk2BJm9i/jhnW9Dswwmj
gqqVQvsYlK6htsdqK3/oKAWF8oUmwqYVsW5SUtp/qRwO8cZceyvJkQkrR+Q4G8q61783gLKeKZsb
rH8v7mdtVohC8oPUaB7w9upXv64xDDYwcXOOpCb7uSDefBux+/SIeyEssTkEC3mXjKgl2+x33Y/B
IPW4w/v2TCuEMJTZD/EDlOLSKwx94Emfl2uHpUJxK9GlEjxZOVfYHCu7HvhnOucGzONtpDbt3KOx
DM6nhVwj7cQdNPkMV6Pvxo3ZNOXEMJdeYSaIdC9TDL8X344mc+kpI8guTmWrd/wwvR0whFEq89ru
sn2dRpMaL49Z4QjtyXWlJuLCUtoIbU8x0EOGric8+l4Ntfr9lKrd4DN6e16jILwu12TzXYqiv80y
rTBnB6BG9hyNHHcpz3K0vL/2EbPQiUPRAtKiBVTN4TOu+yAp8ugZedQUk4nb4piA1OcUpWw7iunT
Jsu6xIOYQXWYqV6teNU82RN60WZFQd9bTiM/sgEic5T6q9TAlh0ZU9/csgLsDJF+4U0RQmijxlzY
Gt8rlOOGs15KJcJdzwv4PAp3voESB8hr24QfmVUBO3CjRu5T9AwmYcTwFH1Lj/gJLEBHHy1Mh9lg
f19YJumfXhVU+KnIot52lkHX15V+pbuKRQyytC/JoHAljEF1y7ICbrqrGB8d5C1iAvFXmUUD029e
IcgjhnTppP6tDseOJE8jTfGITkqQpHk5pQTOw5x03dGgmuFls5lORixj+WWe+zAzro/MQmzafWpz
AJPXgOfi4pYGYxO8PpM1jEh+/BjAOWjVKde209y1OsvzoMoMkNtqP27RQkuXcpQrSEM+owrjoDg0
9SxdvTfpFObpTyanRmwylwlYtRyG4oUa81GMMjeNvzcjevrSPZFdHm8UQMDsaDkn1EFD+MgxmbaE
UD8M9kcjArR4cWaShI9bxIkUl+Da+SnhV3yy1vn6uGGxtEGur3hdzf5wAy7L7U1jw+j94GRBBhKg
/YHoYKY0DQKjBs2lw6WLyjue59i86K7UPejX3DmEWaw28jfCHCiYaLcFa6ABInD8mcfq9VJLgrIj
nfFnS5yt+65Th3ij2nDKW14trMbaqNB7sHf24r4O6qmIRqWfMzDI+OCiCGPoVBLR3NfGRqRvdu5g
gCioAkIlfamMBc0Pdu1G55D1b5y2F7Tx5K4mHrbIN25U36QTOfcGE5EeKMX+9cTvV3cU1FI5lkKM
VT6iFsu64UL2GDwWD18XncZvcl9ke7dL2TGF9FKzkOP7CcESgtFKwzwrJmFARUMSyYdBNVgg4pRT
mFvTxlKFs0L+gBN6TGf39S2GZZEBElLto+zrQ6thZFZoET66i+8KM+tPFK2rA5hIQJ4rBqgh0hc+
88iwWkwyfRD943rs7ItjvBo9dsX4QhwbA2uuec9fzk9B7vGXa8MvNTTFNLQgFnAD1r3Mo2G48ym0
3PRQ1wGyT04Dzuf9juwDqL+JwE0lVuQ+CAQPw+LRrAPVsF/t2DkHRw9h7pe7fAMhlmSD6w7rTjUZ
4QhIRY7gcxdtNoyR9EjTKFkH4xjtNUCkv0dwNh6cfDmOl0T1qsgeDf/eoBHewUXIUUOetpAAhsL2
QFT+Xq2XIRpFhD8dSMyyAZxmVwnZrjvKAxA5bTjPPytg7xR5vfbVfJQmwjEGjxYwSqRfgGsTBHym
kMX2IxdKnKwq94oCOoo/CIFiKknNGksq7Bgh5+q8u54KWBPd4JN4ORA5025+sWnDApXepICrVuwt
8lslPWZkT3Myz+IPwKIDwEapZ3AqtRMfyqX7ImPl0Fde4LEn1xTNpzkPjWGcZdg5iDPntlHozrMY
koqWK3REZjju4R5tPkWa2yhI0xMyom+IJKx8dgYbj3CotFKmHV4aaGmhgt0axXZegr/kYQjOzS4D
IsC0ck6fL+HZHtlxWzo0UXMdV+YS1zNMm2a9l+P1KNavXJCdI9Lq8A3CgTc5nOQS03yN8TAcrKqE
uhBCsbji21SfS+WqJ266RdqUfjno5+L15WrVIrpn8VcK9+uQU8ifh6o7bX+TUMUg5+9nG2R3YBXw
9uQFRNspOnhPcwu4KFXsoP3/lQSGOuosPAOZ+nUC0DdvyHSKd1hPwhT1pfyvISBI/SEM3zZDO7B6
vv8EkHTgj0jtKghoQogNmqTs1JeP2vcV3af6lajEOnglJmcB0vMHdIlc/t9hfQJBgCRr5fqNzU7e
I8ShDvEfda3LlPUI3VD50DvN2ITONtp96LWHdojcr9wrCGLGcbT0afvTd857tcM6ybDs7T0ON162
8SVeQRujEOzWyyFp77hDW/p1YU1lZTPv58W0x4SdULX5r04KX4iHcWPxMTjGreHeEaqpwTQ5s/jR
DN4Yy5TwQGv77OJ0Mf4DUb8QXV19t1mz78gBkhRxY+w2oiuJaei6R+G4ftC0UlZ1N0b0/4h/l3Pl
nwrO7cznvFgAlX07uqUTRvukrzqC4NkuVCpVmqWJ2x7/ovnBQJPd4d8yvKqZSX5sNd7pUrZBPuQ1
yloYTPiZ82yMqyVOdWll+Yn6RDsEnvDwkKg1FyM7VDdLBst3oVNLHLoSBt2gRGELUOE1TNmcbMZp
wY5l0zO7RRQgEHGBxdGVyaOcUruPfdnHtKdC0NltzrIW7T3+B15HTDwU2m0wmBvR2RUKfJoCp80+
EHWwcTCcQqZWyNae0zGTCrnWKGioT5sHTv/0WUnehqWVMWVblFUA2XYC3C8KnFvciKbYQt7deito
YqTAmhuwkjNz3XRxpmBK4kRRPN6qZQBhT6vvV9Cwg6WulZTqp6BBCDuXSOXg9uPL75PhnVwCqeYT
6Lr+MCXLuXMBnUj8Zt4978UsciLaAAslUmo8WqLOwu8WJkjKhszDi7LefL/eVwTg6hf84rwEyREI
M0GqE8YPitrRYNW/KZUXtrU9WlLm5u3szZ0BmyxxykP3QDftKRTqde1ZQ0iIJpB+Sgo2WhnPS7Lh
k2w9ZfxdvH9VzTuJhgEHZt8emMmhvhHTEkCjiOrvwVn09SlDKEkDN7Ucq921++qoI16MCvURoejF
kbu+Ze3tXguRYo516Hfnxkbet7LUpSWa7S4rouUe/pMQ99mCtGVOtwIlaQc0QFIa1y5vrx+ge5fK
tWZo3ESTslaXYpM8C4XsiMPp6aaBCO2UISQq3gPM4GIvNpaLo7A3p2bmhBpjr/q2OZjLBEF4EbiU
Z/T4OIH8AP+l2JzzHrUcwwguvej710OjyXgMagIZmUv4I/zOh96kz6fn3eb4DO8Ro88AnLKPAhz2
Ue+qZ6JSbfGAt1TilY3hhf1hyFzsg5hajpQSv6uJ09QToupwEUIVFWuic1Uc8T0K8+kdAJBkd1N3
OlPntfVb/qkr7+OOcitukZ0Bzwq+HGqHCvtnPt4NGjXqe0K5mhGaEtxv8SfF3ySP6RUJKYiwjJ1U
lMzh/pnAoLgfrB1CsCJ55WuCmTE0N4+RrcEDmmjAmLRyYmRrxrb6c8gkNd6G9Kz1F9XMqK3oPYFB
NRHl+XRIKfBiDtlE+mBhr8MdIbPOsGQQhWUXV1L/AHzQA7l7Pa5/Ls0NnzdZBUsEqHyUjNWDJzNW
d1mpEm+APVZvlFIlCOLFZIgg779rsYhfGOrYnbhHqxGkNec2lg0VTMb9sLZ+/bHHwJosqg3z2sq2
zS5NMkFffK1KsKJPFlW4ECioSY+gDMb6dY9LZ2Z9T86VyxRbKb8Yf+LSTAC/fEEhxlJGbLGo2LdV
RUBcwMDUVGZSYd4AfdMzpC0JTNvAWnh6UJ1fwdX+nD3kfUGEMZ30B7FpCagXIijNGgX1dMemalbc
wYSHsYMvs+/FVihB/pjhBcUkIcnRTAgsZEe3fzf9HYz5wR/SlZOFJFW9acu6nWRyoWqjf11Xri/A
QjnTv14Q95YfH0Lt6eKuJyZ+iXpnDjocbYg0inuC7cvbWe2imvdKtcCRiCFu6NXshmTrOVaI5eWH
V316bjhFcS21RgEvDkEa6mmXJyeF2dS1RvGx1m81rwRzKCuDNTEO/5RisNb7O3SjSOc9aprpx288
iHzEBHK26ufGLE+8S7HuUV4M+zHOABHMUJ2lE8tZ1DICZbmSmRckRk/6v0ipn4cQNKHV9bq4uK+x
9+wc6uxNwlaR1fSExeXh9S3d5lu6dy/Zsiu+K6QyceXqIy8M5CW54yzcJgSes9ptlDgJh1XrEM0R
9rV33XhSL6SBfVrOrZ0m1n+yKl3LSXiwNj0OW/+tnmh0GSEXhWB6s8breQT4/Mmk68egET2sIUei
ZCFnaMMhXK3Mm2IQvX9bOhKUl7tENp2oyfrXoKUlnzdv2D/Dph9NFKTh0VcSq+sTNgT4s7Vsybyv
4DskkubHCRf4kUpX44PJtXvWWFXMCOhlpDnq73lYu23XKbLL7e9Au06aQGw9chKsYEDpHd5d4NaT
LF4Z03N3MjY4c/SybvCkPbffwbbg8sn6fW37EYVe48pBdrtmhUsABsyk8b2FDG9SdQO78ZcJqq5p
fpXq4K4XASh/dzR3qUA1XaowkJJ5iqONxgGkU1nlSPJc/c8xwkxK3UZt30PVE459ccCpV37t63AJ
3tkFjcMdJ+neIAiFseCOdWk5wbj9CQ7+N7lt7vJZOfTU7BYVhWZRrEcaBqXKe3Z97Foi1c6jfjzT
tNfTsU5jjKUyExfGl7Zp131A8otfZK7ANmcj3cQDiYExfSI0wqGAh7utWoj/EVbaoqyyxIswrIdl
22ialjVDMHMV0ljVpR5uU3yh7AgbOUHTtVltvoEe5CVLyCRb/xEiCI8VPU3RcK3gtNGvC/J8gsDD
T9NGMLYrHlXLg6p327XgT28rJ7uaoVnCWb+NpSebCQ4aMtTDRx6vfwvVkouh8dJ9asA/Dx0CF0Mw
ox0ng7YR2u4qewjda1Uy1M1zicm+uajGMmJ2XXz5DwSo+AhruBJSffnudruX57TsF1NV2w3mNQv1
CaLEtAQmAccwN1kttjmKFf/OhxLrXy+aKy31i4MpIphy209tlH5alyL2FB/5cnknTF2yP5hbm6/P
xh0BUsOvzpTrNJZ5FdrQPXk3Q0VEH6dzsg4P3/oP+Sz7gdws96B7XXT3YZIqjhZWVKPZ4T1bfvhF
8gEuF6rQYwPr3XCiUkPs2Oqm6x+mjxpupS3qupwDhqkW2XyoIkUrbcDKaR1ibF2Xi8TAt3Zc+2dA
VKEQGK77zKLp9C6eiWAB2a/5WN5JIE2gMmse57SxhJgTzVt/Ov9xjSxbpaUouSNdQsXY05gzF5zT
g4g9uPjQIhgpeQ1ITPbji7mlUm4mUiJcxEbreuB/Pzr/U5A9ckkpvRRaP4WqmIC240zFFl+aAxkF
uhJotNl84Lk9+Y/KGIbNDjnJa27fmYtfznIuvoAMUJn4W3KF4NloXHCnL3RcM3yWe453r608kXVU
SUssQWfyc4Hb6OwwkPP/n/0pAw77a2I+8ZgW1JwWPDAARAzQ2DwrXbEhdFj+AAt28kxf/eKpM+Lq
nenIT4icWv7xlkTj6Rk5xJ11XaM9FY3z+RG7ifuXB1WYimMNHXplOu/FoxQnWcdZpZM8qSVeQXxu
yVD/ZvcbUFe4L3yrnW4YSWwYKgr8sD8pyhJ8mx68LxL8vSh2Kh/n4Oo+JN/c+mQndyL1BDYBOgxX
W15ryKUNPXUX5ve+i78DUquA8XCrY5ETA46EWg0/Ayojwb9RcSpq6cohjSlFYV/zhdNpfarWwqMr
Ywm6cRd6Dwosk9Ghx92KIKS9GL//JcNhDJlF1aCJyU2d3JVz5qAkgSoXbdbcsLrxwuhN7Kas2NuP
UJOP7ePWiMQTsHispmdCBfv51F0CHByuOoxP5B/IjqcCpEjKVttQ2MUMi00dLi0TxGSuDepQnkS5
PX+VQcN8bBvCbUN9Q80rWDbg58jNKYGY+ZJRxzNEsMoKIuDF9l7qqMB2HLvgp4Z7/9+9VhH+VDZJ
gsqb19EXzj47qHzJ/jYYhsd7tckYWEjqgajfmtsgWq822KzXxGtkZ3S8VgsD9RgwnJEMl/3puWtp
o20NWuh97bmVZM7oRB0TGGs6nLV0cAJsdSI4TiaDvexUGPCi6n71MGidO95HmPyzDizVjwcCi0tl
4WYLOL+Dj0n6+OsQbxEUUg7HoE7HunI4tceDrwiye8789ZuD4Pr+yxlfILIoay6miU/1dk8X2onH
Pljgifa8a+rgEUJyuRmSr0FcFbzP3teLO6cPBzZ+2nEoCjLCefSVW94vbmIz3NdxfMusbTfs927B
evaBUfCF6GRN8jznxm0iMciSAXHvwEsWhI8HPUFnVRXw118j15J0HtRvw0UhackOKqcvDXsHsvOb
j8It5sUtERLB3su1/lwX8JWw2PHtrGa4p4QFGkG1uoLCnf4zI6O6FUXhuYbYovc3qAFznBLtLQrI
0NBP1MWHcuqLeOWcbG0+NzLy8ErcWfO98EQ44D1BfRfNQndxe5GgliI1hPoPm8mfUy/x18MXfHGE
86NckZ7Xbe1CKtOHq3KoMRrVy59cKgJ7Cnrax/l9pD3LE4xL98PH/XBSo1kiXqSNDkiZeJO9q0ds
dPC6/h2yspV5d5eLW57FvQ0cLhN2Kz4t5pyUZtwAuJhbMw0Be+ybXL2KzlXObF0iQp54BNex9FtZ
8KhE3IjTocBQ7s47icgALMxB+fdf4a98bEY94/5vO2nS8nybcWk3Aq27vU1RhKDJFpy92Kp8+QF4
skkXXKdA7TMQE5/+9MmTLEOEWvfOYT3Dgk55McGh1G16q6FifLvd1WGSGU+6k36OVZ8OeAiunt6R
sVO11nYxnuUbYLEYRYwewcvGuA1jm+gatPB5Gnlyt9J0NAS0KsLQkw+/22ihW9TWHmKW1gO6QWRb
PvfTYOJLZHTLJchwLUYXMWEht6AaoCTWRU6yHrd6qdNyMagmpP0v8vUzfj/TMSY53NZOXwYiOUZc
VYViLBgtQXMXz0mYU2AL3xzdzpjJmz40P+VjK6b2mo6Xlmcv2nnctIwkSSSQ+Q3zPt1dtvF3Zb3t
WW97jbn7W9lkY1W28dWcKQLL3cYm5yRxtS9mLm6YIJZzW1X+X5YdlvlR6Yd66FsKF/N/pe4SvFYn
8lh2U8wlDkO1z1VHt5a9936E4z3ZSHfTYJV7ylzi5cS1NKwoVCmafTDVgrHWpGsFAHcwfl0PIhVt
7Yl6AyHmD6fnvqaRNAoWqBs/pXltb8CQPATGqb9e3ZP2ICUYvsKmK+EFdFMGSNLb58grLnqKZShB
FcUi7V6wJmpWBpf2LXqG1De8kulRjJ9x/DpuMA+swJi2PjrrBlcxLkvCbGHM4i9aocFS9mVaLeAP
sgNRrxNhRz98Y4JWClS2zhVWzejrXlcDQEMoF3U+24xHs88XKKVFbA7hs40IW9iXJs9P5F47xJg5
YAVJiLRs8P230S/YE5vf/EPetEoHwLNtuXPcWevc2YrvBCd0ifQruJHD47xdPuJV6LB4LCofU1rR
AFmDkDWB958zleeHhGhQ6aIXChIONA6XOCv5xnCIo9kifxxgBTxY4buXkaTjk95rVgtFl54hSr4k
Ez6HqzT3UIa5IJMaUnN74a5GFMea+jqB85HY2o8epr6JX8iSc0AqUya70G46Q4qr9KIqWUV4zK3B
aIqH+IpCeedJLcCxu3IqR8ux5yCi3up6UysWHbFggQENO74ECdZ4SPmHJqgYNK3GtF4nnkR/N8Gq
jrE66C3Uaur5jBthKa53dvACZ88Zr7WCyJg433ZhZ6kB67V27V5w2SsRTHltgP807CEmyz4Q8W4D
HyTKAjk886H5PqvjEuqoD/nP7GXgE175RH8o+A20wOOEwl74znpjoNjFqy5bPf39cSGsmf7KAkc3
QHoMD4ed4P/yFDJGvrXDXwWJB+kAkGBClBDlm2Ugqhfh+YogVmoP+vDK8T5Bi8AaMQxkfXwOJegT
/VtmqhuRY0Ko08wksY/LxbhWnj5SCAEzdooo8MCkWkhG4F9S29AaYVUB8FqxMxyQsWQ+J01Z0PmU
PAaQnyJ9vHRzfgX7B3wLNfbpppzGTn+SY/mxrj6NxyrCBuJQs33km+TcEoZfLp0STrA21nld/94v
SdaTgrK58W9CQ0hhAEPRkxhzvdr98qETqnM2k4IZZrTmLarZMg/dOC3Hk+Q33aSJHqeZLtb6fApf
H2MGwInzDK2bfdT2NHMhJKkDhQzvcRicVgIVM1W++ZRBtVa4JOy/Rfp1bTb1gYpAXqsSdISXeW/u
kkuemZAl6n3Jcwmzt3fDOXlKCLq/pGnSyZsJyKfs4Wj0tEl4ITATRCJqB1StdZRvUN+tXlg1cQmb
P++LvkoZiEgwpGBU0/FgCNeX0qmpHs02NaweqTfLeDrmOkdK7Y0HhWLRglf0v4dMpcrYTXgPu8w1
4WJ54Dou8TKNMbPFGtkhyfUguY4cJfB6gccgK7GiBl51CQj1ZCx4oafQCIV9+PNHrFArdpsz/gB2
3s148pNfa5hACfD8HK5YX83q43y+Bh+sOOZix5mtwSSJUAQl7D2ezytLJy4oI5s509d7g2xBzD3k
D1aHYR4ASY5k/+fu3xXfj1LA7a/mTAulAy/u8xgHMa5XclrZOwewNDIv3EehRngSlTwnUvSwuh1e
8uUVnweRI422tihl9FuZc2uXkrTwhGxwhOEvIWnNqiwa0vLnr2sP25gxMGt4EGShTmne8PV8dm40
6/A7G/VYFCc76DjEfhPlHNLs9F45IPB9gRYz69HiHenU0MBKAkrbpgk5okctVjB2mS9eDrYPTDXZ
heVziF+fH9pXuhLLj4GiVpw9LIT729Z/4WLlm6h22zDbRMzn0ceKtgqGqbNqIFe2BdBf3FbnSEZw
IbkOtw8ootC4rMCqXCNnm2JGt61YA/EyB0hmn5zVz7Nx56EorX+U6ElM6AOWReQKR/fIDPiDP7st
gkddn3WtjYDqTN7vpimA1inX/2SVzqzg3hCZM2WhZGY5v5AVT7WYxV2M5jqsNVEdVeRDLhR34Pje
fCO8y+ISxlz79kbDh8kPnHpNX/K6ntD2krysyBtvWWTgcJmFk9SJ1o8SKMAqJqlJKCnfqwKOtv3m
uUH5SMhbhf547c/YMLy2vTHGmpLbVeNFZqxbEgZmVcZhh2RVHtrfE8xCokDMIKy9ivcPmeKoofqn
yNEHuKkL2AIVHYlHM+0V09mjPXvKZ6QWDegAzgdI2JiD6E5xV6IKrrTqT8vVTa9TFSVy2iObMJyV
S16tFDDc8sBRbVQ4S5IqDjozvq97ae2HF/d2eQuILYQAYhBqj5wovixvTS2ffbQYR6zNmJ9+I0pp
MNFxGJIb4sXGZ26sF/Ox3UgNNPWgJe2zb3Noi5PGbAgV0HHMjj2dmgWWyimg6p8pR4OvyK6LW2Pr
UDGeuG+fa1aJKHVOWAY3t5p/1ZecfYsABaXS02ompnVPjP4Qk0ZaaIa1YFK7++v89mRyi2oRjer5
R61ICckefXtVL5XvM9NcBFBQcuB7tw7m/67MS12AJLo5IBWt/3pD3y2sBNP/yl1Ab1zUGEOgj6o0
nwqkj4sfwSq7Z3sIpHL/lsy5cNGix0wkkm5qf9rv2FcyF0YtC0tsXZ26RoiA7/8fwhdGXkq8nUct
7Ezn4Fw52quE3OymlLlIgGX6JQufGl7OoROIRShgsavS1Jm0xAZt5ShTb2etUQn63WNHYKsdZdUK
KunTgpppHvEDR5uHrBvBP/9WyzBbMI4Lqfd4DX7xlvgtrlzJwvL2JBrBQFFvIeVhkkPPyVD7yC43
w687PHTCDybbC20A9zvDNLRwLnW6NnKIdvqfcAi1IbHdwnQzsAJHnOVRqgicSiUD5ixGC8HcpD5R
LtFxLul/y0EG0UEnq0QvM/+ttzVd0ULb5EUdKejILtcxuVABRoHci7zCRqVg/xbjrRMNow5b+d8Z
DN6VQxE7oOsgxz7u0aIvGwU0e4rVcGr5hTz2ZI6fqvIlBgj0E971+eR+7KTRdYAcXmsBToIQXEdc
gERVtcFYVZomBdrGJe2kasg1veTDH3f80lvjFvQM8O0UP0/7Cg6Y7e8RRcX10U9M7W+IPrjJL3Wo
qdUKUQOLNlqD6jjn/JI8vBFm/32Pjnzkb9oHnB7bGgRto59B/sZQfp4LRdunvdPGds8hlaCGUo3U
PGVVaOGnfQ5KuCquBqqMOVKxscNcfWk1gCGrzZdQl+YXoMxcj+NNKEGmpwah3LP9+L+Yxz08EA5I
Ihwl4PllatgKjY+23/dcR6Okt6ystHU4CrvMnF7wsS0/nDlvBvHXVCRcqI4mD6q/tBw0RvH03fS8
4ZbYF2GOnQllmzhLP7hHJ0y/FXLtxlm4PRaIHb9gvRPyEXMUjSAgEXUx8WasYP1tR3Sf4T0y+N+C
lo18ugjrzo0dQmv97x2FTioKcKqbjEEgRJn1wGyIS7vNSrxG+a7UeJB++yJL07ZgkWR74VUN7zKT
OuocYbBRVlPmEoaH1i9usTubhplPpTc94NhFfrePCbR4m1YJstDsJvczvw+3L4ynZsyOtwB/QK9a
BD/9yaM26G4omWL0qR9RBitBZzhECrOfPpMIGx+LOkQZC6Dkje/rYueKwFlxwLqLazM6fPuHrloi
rdX87PyKVKFq8JWdZQQMzAJh8yfScjvAhnTImYMs7u8SXu+G1w/s6NyjMCmk99h51f3sos1UgT6n
4MeCUv9uXsbdvMuDb0stORjBC54Qp9ho4ilnwPJ6CYYKFHxdJwYuJzHoQEsCjbXYXWofmwfrZ1Li
eWnjZ453GTJ8dvUwExkgkjN1zL4a0BoPbrz6cR6JDh2z6HW9cXaUWzSGCynjLa/FfBLtkF3sVykH
+TBnP7QpgE4++trEneVHYbZTGfYcWUVvXp7hm2vk3a7NqvM9m3hKV7pVq9U4xJi3I6Gp/UgTakfS
scaajHUMEYI5yslfR0rXBAkdvtr0XWYwo3fTG8eIe77wLHqv3zjF5MgeHf4mlKHwV13rxB/sbgC6
b+epQ4XuWlA/KRuHrYiLiSI2EuqD1EqIbzv544BFjJdBNBAUPczZylG6S5xhyckd8QUkMjRdDRGT
KD0vexk67d/KTvecQzSBOY+Rs8V2T9w43GM6ELZkFkl5ikdTHUtztSBual9uvAXErvJmakccLCCQ
zm+LmC0/HztQVN97RarJHYs/I9kdBzCtZ5YcIO7RP01MuWfY+gzDKTwbiVqzWI8SZT7vSXFk9oLf
CWOpXDMTdW9LkRLr8ZZspFn0OepHMpnZ0lI3Hvv+0Ha51IHvl67FFwWP3HyLVlmv2KEbKN/0a/6/
kV/PdRfmN97jeuUa4+N0/yi/0DlnZ5B22uqzi49D1/LWrSnxNPz+qwAozkTVOhK00QbkJKsGzRYo
KhIFwKYQg7LL71WJqCp8ircbbXdkc41OYbJPDSjUrwz5QkWovzEBFgCfyimLhmwG9tu/2POwrBAM
Lv7Aoc3HCBjYoIzV7BmhmGokVqO0JQ7zL9YmrWg03OPAS3iHh4JheeC17+pmvKJ3P5Ft6mUf0smP
TMPCBz6YrwiBsWvUAnoT8wxTuGVElGMBEpIgGRty1A1GtmfMbLinSvb8YYeyRnZbODpWSkDcUqT+
ssxaleHrIJtWuqrK1DtaAymxfAqoxLhDosooOlgmqCkD1eDDxy/TXv4VcVIOje4uqJL7n8HapYE5
M3XYbv+7VWWQiqjXcfhiLjqFR+yrBe3imGbPHJapXrsJZugjEfKKEYYiPpfOr78eatKtJ9KYadlq
ZEw7xE7y6c3JkU+lLo4XLWcZKqf8PzQGjjFof3yOXMok55KBv5HJrmEgubmHAFZSxxVG8EYrmkMt
Z1ZMqXemPpwUEix2Q+5dGw/UILRDl7/9gL+shJJ+L5D963kSg+ME7O5+APOtua6M/iHbQC7pWl+9
LW88rH0bUtSTkD8acorhp7bZ7uLKK9nwT9ANeC9AsiA4UxXSSxQqDS1mVpg5VZHJjICuqW+Oj79h
PCNh6wGID0SA+kwwfJkprCvPbTdT8vGtMZs9Kw0wkDLlTZRGsl/BTTbyjJg3607ReDeXRExv6oxW
wl6R9IP+fivuVFynDfZlBOV+CNBuiLOHJUQQHhDtme1cA2NRn+FAxe276wtCtBW8LQhJDgGk+W0Q
dVWk+ZE/9LWcv07Q/VgziZLhXGAeLK9MByJguMx6Vb2yYdvKV90iyE68Jx0ouN6ireGf3/Fn3aOY
BAa191DetbJ3Y1MZLXVbkRLc7Jz0TVshvyjXglF4R5p6PXdRR3U9PXVddzP7TObM8a7Qv047/b8/
qY9FmFqBp/1WD2H+p6U+x8993+CeYW+aax5T3kWQiOHvM8vti/ft1NBmBOaSy0zQ+d2CvwQExFEp
AZgVwbNBBYGXzoXvBk2PpHQAqpvgRJwqhpKVymSqQaM2+kIv1V70SFCAaVz4pZLxzuXFqpTaKINK
IH7vZ1PDBU0n80Tf52KX1buP5rxARejNONQiputt9GhHhTYZJP1OBsZi86I7LMjhls90pmClZ4gb
9V1aF8P07wkFWEyZ1MDd6FYSQMtKlIsx/yLVQQaxpiIpxUIiL2HzLxbsA8VmyOeYXsBZVJcCxkT5
zhxeMLH2haKlbwjq+uH46E2j2aHeBX6hnNFplU/lVE1/0TTu7ov825jHMr9TEo3rg35mEEF2tMNY
Hqgy/feEvKNiL8eyyTRSavK7RL7KSMbZkUlo5NtKk5FQK6YxPI7lgvft2EE2Z8TgMCySfy/RArcY
Jy3loC6Nd2xy4qtg5HPWkzFhX7UoxYvJNPKfX77l9UFM0jnXzp75ZobCMLB8fqZFmTTGLBvPOSsU
F8oZJEyMkuWVOXYNZm6m2JuCxRfjW0HSvGlaNH3FroIgUiE1Q5VIaDXVJVamr8wMKSvlkXOJr890
QzKwo13jVMXv5/E+OiJarxucnDFSqStg+H55PFU33GTTiI6kn8PW44vyVQmbrriaj+C7R9RHrkCp
S6xpHQ5Z6Pk0KTIoXcwOYTwCgw6HmhSw4kFAt8jmFCXUa96k90XM5BSH0o8c/GdR9XNVZ2fPD6iA
4+rkI3SwExyDIv1i6L2EcfIZpy43u6UQUOFsTacwHuBiDT13s/jqNkAsiv7UvigGtTVSqUjtCkY5
IAn9MMu4eMETVjTicsyrEAOojjKiZ0N/2CaDRRGRGeYfWLaUsMH5tm0Qmw7HuoM9fF+R/EP/LYNz
NBhOLw4bSxW8KiSIq5IdYfbjtNRW4/GgIZJFGnb7++3N7Nte3/lvWiYMRf5wJMI7A9QuR5bCWbSr
QiRLTon11GpwENF5tSzHNjXL131X+K1rINrNszCTPEgWctV+HBqeEeT4d6qMXvneTcUIHz6KmVyU
xh8UMJsbhrFfoANhEMtWB+a+aNBY2QlXbNr/fkz9fSZBJ+7e57EO9NFcfzdRggjyofNJfK+xgnCz
RF9HKb0pv+ZGNNwjzLVSX6RvFroHffDrE7EO4pA4CNB2aiibE8gFLMcb0l1ukDr5NktZqoBdM1A/
rudpIQD5JXgBtkLxa4cn11/4ep4eJG45CjRF0hrr9BkyVXzKK8m87A7ExOSTs41RHYgdtd6KtouV
YYbo9IdGg5BhYRfc3+E08niFroM3RTXZE6BGMMQg6EPpQUQI9lTfJkRFTLMa5EuHuXR9xaS7jRQN
AKDadO3fTIZ50OfDx2dHiPJUQiX8Cb5m6Q73a1aKZgKQB0/GImaz28v/Jzoov1If0RsHtmrK/nNv
TlTqZpmIkgz1VhcSinEOgJUOJCUKcfJBViPyQeRDK7MkR04TQOpDaYK66bszHk19KHHGVkG+iq4+
4OG0XSalll4WACVhcy7Tw8GspoCXRMu1FVWdvz/eJ6ZoRFWYTHfN51x2OApy8ERElpNHTDDDPzQv
TcMSLDGoB2H77NzWinriGCQUautckmT32nbtVYYjVQMxYYkGjUXtKzZjf0w6K6etHpbxg056B2Gu
YckiEVnMe87z37nKouKv88phEDh8+TZX3FrPDHErGUwjHKy+szpojWk8x6LdBuT9+WmOjz27GxKu
Jo3Ui9eMum48zB25b7BVHRtwkS7pnhnwxjK23H8VaM4yVX8So1PAgmpgKrskjBTg9P0BS7iZliSR
SW0uYr1LFbmz6tW1Qp2NtSfdmsO+v2SDt5nw3GI3nXxRFTaqI++bDX20BKayRM95XCUHXMyQ5HTM
cSBhV0lcpbURcNnESlmCAIqY/fwx1ans4b+tUg7k34/CRNBMMWCA8R6a90Tso84AGFJEzX1k9Qgd
Nf69/w7aA7X2cWQ12ebDMcgkqYli/gvlOenZJXsr6ZunPI9MecwXnDV0q+XES76RBNlPZ7Uez3nj
gIRE+QmxkWa3kCv1dJLiiCaSNi7KDuQl0XlyowbMh3HSJvdAqpXS5hfQUdpaVoyrGZBXWXX5rliC
wyG05/i9Q6H3OhKrIOLxRbeZTgZ4110TUFJuMCXXdHeErS2+bGzUpPPbOLv8OM73vyNQ4Vp4FSna
Ih9dr94gvWeJ5c4Mc1DvSmyYiqWqvVCqnsfVTk+y+G8cAaSSdXHkVOo9t4/X6SbosWTOHb0w7vhp
A37oQMT1m+Q1UGz8N8j+iOU+sdj5evP+ETBxWRzRjvj0UzOIciPP0dlAXzIPy9o9OIW5Z5MiOk4c
jDQlO9p2qisnE2IIEaZHCttfq+aQOB199iuiXjpJSggt8bipXwrybccScK9E9YOOjz/Mz4ffxpeY
8odLgITNzEqSHBZLpMhbsQJN79IdGZ+Qv2Dq4mGtoGVWm0kXVtQRhJcytmfPzQlmgMH4slEkJCYy
lnr0sf/G1s3KTTicmDneZPwXVSMxhN2sgdqiUcdem6JR9zHm0LaOvYQqxtvQvuE2kXHc3xa0UZKA
noHQ4vKlP0gf7ccS60j0iA6QFWrgek4wXu+sptsngb/YYTrcMk6QNB57tHyadPthO5HLdthu2SfJ
RbksGPRuh8SayuHeZwVzpy7c6GMVq7yVk9zzNvmBTj9+QM8v8YDbNNhRtNf34hzXjsZ2zdjoedvd
YWyMQ+puXaPaAmB1JI2bts+LDHDH+NGpdtcGQRCtcLubqPqKSfF7Z0L9TOLD7/Dyc2KiPIuQ1ulr
CBZ4UTGzIUkuMYONAV9/J5hvwUBoWSK4kdF2WacVFiDASML2jubC+9gFs1db3cLxYX6BY4XH+L+N
yWQCf/0oa+HfPEOnhQDEs3aT3k+hI3cqilhefCkGzQVBzhPx6M8ZVd6HT7ZAU/ocvpwav9GFGp75
KdEdqa5jGdOdIdMno4FEKkSVzOzvwy/CfevFVKFyQ+0mr5ThstWmfJFnhaM5UrW8bkgisdksLC7d
EVyuFzcHq1i37cgkvxf9Si15UGkvUPLT9z7JqcpIkFX9iwrayB9swb6CAni4h5QmSu3LspkDHYTq
7DbCf7iS6bqAfLXwMNVjIINuR7Pr32S+UMvbKf5GZnUa3DS9pNuN7kJKn8pbCAnzdr5QXh1gW7iB
S6c8jtIaCOPLirsfzllOCZxilFvVMPYYGvpoTGu71oMxVzywMBE5BaK7Qb3Rhg1lrDED9XDVJV6Y
SQgqsO1hYqxn7v1czq/VOM4Tzw50dIyTwJSvv4c8xwjDzDKoOs0qcBvpYTcJRdzhuop/QiRv6UAW
Q13jUHOOcrmP4NweBoxIrxXDhvGChK1FdtR3498lDmARbQ0VUWgzVMG4w7lVzh801s9x+lsOzLd7
7ltj22oCDIL0Uh1CsaBYgTbZUjzvGHeiYJJfX+zqF45zWEb/BRrGi6T97Qm3EFl9J+G3sIb+EIfj
7F79INs8JHqtO+mbDraX4Aktor5uymZ1VduWTsltqLExxNMvngCfANIhrHBfQB8/LpWEfyTVhtxJ
Q7zoRa8pzTsfDlIQO2vs3h+ZQLPArSukO6CoajR65DCNaEIxZwx87c2MS4IokDu0UiA6llM3Khvn
xQ/p/HH5LDfLsSB1qf7coJCc2jAgic+soxqPPIIlCGJnAk4ZjgUf70G+aHPvjVbD8ihfxpxw6yLi
IsTw3bKq97sLb6/hwDu1pSgNmMafTBfhqpV4aHrtAtVUh4+tTludHEt90Vg145ffHNfV+c6EWe7q
UxFQpdwyX1m+eYg1cncUzpgj6M9DgiczZU1LZYO9cjnQFGmQfpIbE2B/cwtwqJcH/S8v4osbjfMd
rrZE3SKHgY75d1pelmBczh/0S2kOssjVhK5BJdJzw8xWfRIvhNpMs7/Slny+M9qroiRP36ahcAFD
n4Lq0DwPdrOqzeuHhrlSJSoy+aSIs32EEpFsocMTA2NankFaC81C8JKulC3OAU1gSJq7sygqVinv
KY7jAe34vzp86VvbiYQ9fZOEuEehe7+WzvkozPt3fvpohbP+Y4xY5Irm5u/N8+r6kIvKvdY/Ix5o
DbDCmgkLNH5KY4AznlAQAQAEu0euPh1SxRIGKRn8cx0PbB8N4DVpzmHwJ/83nrQTuC7wWc1jPNYo
NO2Yv0UKxcTGCK4eqjax2uiFcQN+SNj6BQAmqqnwzqNYvhmeblRGVWZrDfTICz9G3kgXob5z3UUX
kUP9XyVB4ZUX4ZcGSb99GtJPt/abGOogpuzcYjFo8+0rPbvypk8wmezY9t9ZZoD29zNOAbqgyUu1
r6/u76ZY6UPqiyUpQMParcFotJMyy89Z7YSI5fWCFjGcC54BtIn0v9ku7fC24WQ+W44lWp9vY1Co
qS33PJjsQihuoD1/4+rXVZHydjTdcZBYKs3snXodqALhWNC5XrA9YBe7OOgReTkd4onAtIK04B6X
Ei99SO05prftTHEAx6Tpbbw4KbImpptGT9F7lNG6zf5Z/zHnmQKkOm0jO23GFH2NkLVtbDx6PLFa
yC2FFNz+jOXHmK1feFo0/UQET6hvA6XLpYcgtn9b/LMk+bkcU2gF6wCrJkXfxWKKJsuyQjr7SMhh
p77tgNR0zbqsCSniR34xcH8S3/AFJARuA1NDebIguanpPogY+qYma7DHrcFouJ3FmGceCjdeGwxZ
ckJREmLX5gKhRfZBXNRMlDhP8HhDwOh1461jMoY0ojEeeK13up0iHT0L9LTE8YlB6HicbCoJpEjq
DVXuZCERm8lriNAINZOdN9f2GKGYkhnJ//plTWCb1UZyRbww3h0ODVC9JAC4xaBBhRZzg3+0cMZI
sYuWj7Bu6wmf/CnLUrYp28wty/aDNXiums28r6y659q0YDYHskeu94XspSKsdYqqF7NWHxVLUscg
xXWT5BSHr4mLTZEGe3yyWXlpUlcdV0D9CaC+DzpIx0uQS4FqID5TXaZzm9Zf+pqbuat4hxUO+eIL
eCS/cl8xTErqDfkZlCYB8+Kb7Uqnh5vdEvBOeeUvq+UYecR/MCF+AswXrn7ot1S0Wdg+NWmmw2+n
dYOgzymtgA6OzUb5FtLS0Wm/JQWJxgkMXXHTCg1pEm/xTBFw9mUfqIv3ntW+ii+2WQNwmlse/Zk+
jzv/05BFhtK29VaumjeZWoHpr+98fh1UpFDbzS1XhOF5FXc64Jb8TN/CgCqztwwJce/hRPkuTx12
ldzBkN/jz6t2OVlIAvAjV+UnB9QyU1RaBEoRJPtNUCDBi3BbZWOAs9mNNJHkyf6rrfZOln3eU7UF
/l3x7nip3lEYou9e5JMxJ28b1047lm2mKiCDQUKX7E8cThh4vtmsd8OVxI1x5TdTFlJuZ36VeY6H
HRBWzTjGychEnQgHSEf9zr0Fc4PxHi78jmocuaxcc44NRZhxIaAaD+A47V1fnWO3Jj0zOWTKC8fL
jay9Csuj6K3lc8cqBzfX5AViKgRD7F7RJP0JwOGrFTtnVRJSbwaEX9lqkmXCbVKk7vAB7kHJeiR5
1OjQJ0+V88mx+AK7sBh5SubGvv7DOc/LynQ5bs8QgEi22p7JomdGTk+EmiSwwWixMkd/qzBKF82E
xjRwxWTvLQOPqumOOABQwuE9OnzI06ydUP1SLeb4Euf07ycASAB6Io2IHD+3i/ur0+IFD7njx7Xm
OlFQUYXzgTE3jbXkM4tuHvheaDim2CtpJp7TIWRSEV6O4GPq/hzxekBerN9ZW1vn6IOtAeHN88/j
shAZpoPj4V9rr2RT9SROmbFekEVNhIMkQ19R7X8CSjI/0kZyqAhdhITLtEgHw34ON21HS1S4zXvy
Ta8v1+z/2razwr0WxXDCdIxdGn6W3Y7he9zmpRfhooDtMC549F1qQtVeWr6BiKsn6PzqxE0pWqum
torV5J5W+lLmUYl5TtLTydcDXtj7yxBbcpEkaRiFyoL5knigF+3BMUxBev8qtQf4uXYfhv2E9H24
pfqrEu7NhDjBc/oPE4ydA5oeeDJZYYWMlaB+7gZOhIzMijS5ij0Sy894Knpgcag6hv2QJvufpj7j
Zz6mIGBd75j/3oCFyMhLsmUzjq2/rKEolthXutWY6ca8qoH07KcnhTpfFQeVWlM70iMDRwh9A9Qe
YJw6pn1FJ66Bbi9Pg7U3t+1S3fW9AuN2TwvvIQmY1kXArVTsbrZv3xn7lZ+Xbkh7hR39gEh3umnz
X75s5hxpmmRzN/J0L4Cu0FdK6CnJI6iz4CZuoY68Ya6KqwUSXG2yCQp+thrL9pXAzac4xF2Y/+49
fsscw3BZuDPq+J8+KNHqEmvc40vVXAMU1PsPJDVie9rTcnWy+ZWGUixaQgzPp8jYfW/uqjroN5+/
6mHHSCX+n+E95UTM7TWJovI2KJU5us/P4sPGGuWr8ELuuArrPvqriQ7HjvRQymtYZ5m+aw+h91hK
/T9KMZuHeUprYW2fKBEc1V6aNYFX8NqEKyimqrH6yTIazw8cJExx7qP37KLsvyGHiwBiCdzsvOsw
V0krKoLfaihUNCSaG/+1+xW2fYOoOuCm1tg88di7aP8YzcxxRRtYOdLW3d6rvtOY6bHmxTBadpPG
5tonA3a4QHil6g7YT0Beg4KjwNQ5qiHJNVQ2B7sjsKkYYDaF1IwACwpTurMcuWVw1va4IldhGQij
PbBJJk9tty2ijWh0PHLOMkQtlNnUkpD78PdlEnzwmbCCnSsXN3abtPxtNdlpBkLVtEPm3JP3Pl/k
4WVEgMFj2iE2SCZp4BB7i6Zzz0NzFmMoYr/HjwjUkz7F9EAVgS5Sl4pBO5gmBsGxiLjfdBRGC0zw
tIeoze+DYmF4hkywy2NpwnGq4N9a7s5basx9l6kmYsRaCXbTMm/SQZEV4Dogta/TWyi1tjWyMn0H
gNjSI5SvepffXd0w9GJPioZdn3/vGWlUsUqjUpTeMF+1ZCGTznuBYz8tMiI4fgE8f7JLMYj5O7+z
ttUtOjB8b1x5rQcEEiife9s+asiBkB/D9s1rqwUavJJtiSpXHHIItxarEn3o1ej9sPxxqlxbhB93
bOJ4JA4NKWHeRygT3jFbwXlss1myEFh7CjIS4/apUiRAauv1Ks0KGC9WagUsq4znzFHF0vn8/nnf
PeyYIzgMVTqIwdf3atict0h5X9Slw+B/QPs4Oow56+Fq8GGZfsK6xaB/nkHybEUvJfaKoicDsL1W
KTcUVED7eTTw++EqFrgPa0pZpH9DbImTrfGKaxmFGtLUXG8Qjx6Hgxlkuv8yGnucrGeRMNA81wa9
waYdjP/ENecMgaoHQsmDiGSXoXOPAGIn+RLQBjBWHIuiswK6PTH/1Ici6+J6oJZlS+PEEzOExYFy
mlHUoYxDv2dnLTAhF0bFpQePDumXOzqconDj8NX62QNCRGkXD75UIcaakU01Rugv91dk5ARY1rAx
OT9tnU6OZzT/3bW+/o+nPTL4mYVjNIxoR3pb8QktVQoi5UR6pyEc/5WIjAtXgUJkcH7KbF0c3sso
4nXzBP3WEcnsTLKgLi50+yxqniQhIfe1MVQvtPwKJJaOiISTD1pHu/HWi3yw1YE/fVqZ3giZWTKm
ozrBuqGSECFvxveDLgEyEqW/UiTZ0hvlx7dcvY3xS8KAaK2psiH7vnpFc6TLwmq/0NINmy85Xxhv
V0lX4bGej/c4RISVw7z+Py8Wg/t/RPrxO76AwIPEMrVOfr20xdSvUPz+cO3kBiEsCLOrzSoRwi3w
5TeduTh0Oj41yJsamU/+HexCwjrWiZY2laTI78Mypgu1n9Ws+54VS/EB+NRWCHhCxzoJbkfBQ0EO
+dh98OnJKCrvmVkRRF4xttaI8iZNV1igoBMshSoQjjauaeobOp+UQ0mOSC3RMihxH9s/odNwXlEM
ZNFXIpz5KAx30NK94U+t1C6LrsKSJ+Y6Gs92oFsgvM0VFWqG06wDeS5ezNGA4+HzrMj+3zd5B+Yi
JMvVBTNj2mpLnprSQJuIZeU5GW75iwXmEGhCMazOFPSC5Kn6eoQDkUeJkJQ83GkeUtlox2NHH8nn
d+J6iGMgLyvomJZw9hLnWNcXNAMhIYHnUiU4jKeb8GkggFmnKmFR8dfTc+r1pfvLDp/tQ8XIB4AD
m+8ZASF25x9ZJDz0n7VeB89CyhKaXPqe0DRLhyydfTSnP3RXkD2g4sIavvtVyHCEzmTvise2GO1B
2dvKaKtZXLrGkiuaEi5nfvvlbWFpBrHUgwjB/5BiLVsyVi5t6RIjMbaOXufik4AElf1AgijMdCh+
ONENWNVwSXuhRvbIv2ju25W5O3SLYHhT4jsRUV84jzpCvjIg8xwwVNgn91PuvTT5oY90nJgIkioG
tVrq9Xq//hmCbdhNpnCikQOapWu9TpgVkRRkWx7pAgJsG9s8OMGzPD2OmebeMa87HTj90bW77X+p
veDSTm4OTZycrFv/vKyFuoz3lZ1yh9KL3Z8Y+I6ZdfqaDRyB2tqUxTUmZzQtOyWKYEdd2WPsaM4o
Of0pHcmQews/ExZvnRVLuJnovAA6YsBwzvxuqPYQo1zDKFsirnFibT5Ll7jQ4WbFdPyVrE2PZQFl
H+NI5v595SXAuvMmXJ7cHImS8tsNY+n6dcjyVK7sg0A1974xkRgyTwRK/lPQsjExgQXO4kl2X/1/
Kw1QAv5LwdMuXycZrqAhK2W2MqaFkn5xddRGGWoudJtwQLnK0TULhU424gTZgqB5a9UiOX7dB3V4
GHTFjykviEAvbCBBaluF0DXQg1oiRCO9H3WUjUqLTYZsDkUbF9gqpDlHBMeL+NlFNUj0e/jgjbhT
smbc6e65sukAjAWpBJyzEUhtKrE+hh7OQh4oKUBZEv4upa2Z3TR+0PU+3f6xnxW5f4TTSBMJ7bxE
uk8qvVO5gLLItpRivN3Mm13W9/rx81fYQ/OpLXuWc/6FosAhbveBIkdpKzggpun4GsaIq2Ow0bGC
wsIjl/pLpOnTSUKN9owTl332L0Ru6473LAV0ukQ3AyVa7jz7QWwspomuaRCFE/JrnWBMR2gLtaGs
1hS5ERBRJ1C8/UCKELH41Xi/diKfwwRXSakFonT2CF9jIU80PEwq4tdN0Wei3uUaFXlw5yyQRNn6
eYpNZhD1QvtTW7ahJ6pOJ30cQH4EQUMC0HmVLfGXpmHxJuH76qiDQmxG0td48Rk+Sgmy8xL1iT8W
FbZV14vH1Om8yvbq2upd+pR9Y/d/RfDu6lX6dQ7ULwL+YRtZLqABM2d7kIyOEsGrebBQ1ZctWOu/
FZUHgBtY4r+HjzXhhqCYtsA5dpyBWRTNNXj0/YDKiqZUZpLg7/WAo4S9ey1gn5eKP3Va44YEN4iw
Nh3QZNLX8gfPMWRXv5RWp9AW8M0npnOWUaNoIOV4BksTC79SfzqVrvWN5ouxDoQVGbzcv0qPzXGL
P4O2X3v4ETjEFoOom5/3QvXY266MKXsnDjYQN3fuLYw93wohSlBg6B6QMC3h0E3WIsbBaMLYVwXN
Yu3Aay3du/Zb2hwffQIfhjFacuxAAX9a/1jkkhXdkgB0EHXJqsuKiF8Mzc61W5N8QsO1WfjZjkGr
2Llv6xdXKq8LDwFRAVayO0RyOFBdaevUE3xRUpNAsUNudIorTdpw8Vc4wEaAlntbgnC69cj9sefP
tpFy+HrKtITl865dqgKOqh2RL8UU2qRk/s8+n33bV5x1uXdjTzpeT5JkwhAPh64S5fiYboa9KW35
JJhc29an464WBMxBo6jTOE5YVF+b94Gp3EOdGLJCqhVvSfSE5wlKzniQ1XgbF4NM7yCgg2kbANu1
fiF61Ooq9T45B6ttqRH8jHKIb3mHc3vABw/rhfEk6NdHvN+ldpYpYWtcybLHoVA8aT8uPP5u53ew
8f2WWIFgTROFtNkDVqo3WqOKDmQni670I07aSeTL+ZpBmdrlffkNDCEuUc2EFXOviEecU2ajIhzB
6ZIBGMbzOZbVVicqyPoUt+NZcYFn55CVSueFee1k65Ruj8fA+aOMfkl614LNJlyPBmV6WxnWnM6b
lg/cJ/xoe4ocQRI2ZdtIX6qa7bgUrWlHkgZitZ/H3Lh8D0TH9dC6vkfgxY1g/cGxC67Jki6xAz49
zW8YcmMt40O7wlPT93RVo/YgrgeU8+uV3iIrR9G1+9E8L244+mCO7BsJRKLJTF+tguFZetFFHN2g
rpdkBMZ1YuF9EFnP1PgGE0fg7qwy26u0PZfEQruI5MGTxWNzsFN7qoy6fZ58mPuhLLterfIhvi8v
f9ZJx5m+iIDlQP+xZ1Z5xYZqBMc/GhriLU/W8lXz6OLtxzeuiuo9da9yXmI3qQIqcNR4HaQf1LY9
k/uoShwyQwh6ky5IQEQ1M3XIygZdWGF2njjcaoSAwjeOODvAqEq51obzteNPF8Wgw+Zj4H1D6BLu
wLulfNa8MAWhJNh1HxTuXHqq7ZzU5jjhOfv4iUD+HZcrRFSEALHjGZWgHpVvPaLxlisdwo8PFnxw
XtxSuqM4HsYm/eQ0xvXA7L/GmzqpVlueRPRbFOIDWAdgGLx2VqfAqvu+3eqYNoLadNdHYxOO2Opq
rMl2XUzRk1Q5IsWZMQoJ8mU5Yuu0Pjns3ligHGNlIvY29TMbW6QmF4KCbK9jK9hoLdMwZywZ/01P
wgClgwotWWYHYc7O2zZTn0a2byRzIspHLw84a2Qxrjm6Ch9XrD/+YKEQTT0sm5uv0J+zXVBr1/h0
DlJDVEpmMTC0IyGHPb29hWjqsNRnMHOFyMtBNxfaUYfI0/71t8aDYTumbv78KUvGFInTn+9LGHPl
yj9FVY7CWi2KIgeGODC2ZSNolpSOYx/edpg3pp2J2rKj1xO8jDZdCKVDwZSVu6UMC1CacjQyXes9
wN270mtJAOcaYwUEZO9wi5YYvIP7nzgFiBOJR/j0QxOEHHBnHzKFAh5HW7OwB0Q/FIvW8OtjQP3S
9RXl5GJDbePf8kJDnyrS8McCWfglLeWjtO1dRH0Puzr58V0bpy5H+emepA1CM836/ZZdREcg5+7N
9jbEq3NRvsCjuPb+jr80mps5CkBXSHb+3n3hlarvPDkn7nCJAKzTl4mUFCBfxTAqC9VpVNwDZmXa
yTUGZSAoMP21LD5d2PlPlXwiEZBtmhnwogTTM+lHoPUVZm9YzLIDCAR4UWfntpFfB3hN0LmhPjww
B04v/dom/KXpiiB2WUU9nQ9GuhlVrn7he7xoYzDH+O4KydUQd4eXUWUB/VuZvXycejwlbxm32Kud
xShh4sOJ15RRdbVC+dMjcNYMUiXXcy5l5o16xqzyo22n/ZS14zgMexIziPSsCQUBPgqNWA6qjmAt
43C0roYayRWTXPR4JiNkt5h7p9m1+C44Ak9XV/ANenLrIHQ+KRMbTE9czUaBxYOpdOI064coA92b
SvXaWjDVUcg+PbLr2kNRiW0q7mP3jIrvOUck6LKXBrgqTp5EDf2+UeU7IDnA1qMFfRUUQ3sXQLGD
X6hoZl1K4ZY5Enu72Iqi2KcbC+4Kow/pdpUoIzOuN9iMAy0/IJFZdNaRxChwl0o8UhVRUlOqsdqJ
YliFaoDCxvUTyMgP6tvS2TETsQ9eKh0xDw7fhvFTpHH+NGYMjYyTjJhwQVjlrQ1psmyYft2PHUfl
P5Ssi94+7ONs2E/uFry20u8pTR2OBtEJEP8oho+LBjXVIXsMibwtmkv+6t/kQwEpwBKiJcNdipma
/2wZsc+DjWRfR7jm46hO+kK0ScLbPv75nZcizytacaHRBWxJZq6z7Me44t6ryC68arRVXnNtKx21
I7CyWgwD8+INVswT/ZTd6s1gLAsahbwUZXLT40EpH7fvakzVC2L30iQhFaJt68NnfdXJL7Q8pXzO
wYOl3fvla/cNkNHUhu49RdZRt9eHxq8kDr4ICd1cn+PUAcH92uJsCghvR4bWllc9CduIB+VxMAip
vyf7R5wmG//Vo8Zfck/87jGSfiRNE53kHxxC++zYG5JTLL4X0E/dIDkaXLJppgkz/p57DVaNka+Z
30YRHHTarKuLg+RxLTGEOXQ/mBOp5KULEmPztZH7w7J9Dc7oN+u4p3FvqtkzwV2bbiW1tvZw8mkF
pNg6t66CPsrxeOJGYGQ/ZNafk/K1VYQdfnKT/avd4KWei970Ef1OKkUJh/lPsWgXCuuwdCo0GT4p
ijHbCVf7fWbWWHMkasKBc31O/ybcLI3Q2pwjA1G5dDbYyi27dDnHUuDPtw19+DeRrLhq/4fkv29R
VFXPwburJl4BVl1Zi1GpLKgDqxagcNt7EQ7RRX1Xi6yfyaSQ9ZCryxvkXfVS8KvfBO1AGQ/+Dmxc
oknOYPaEIe2mcl8q2CsEd92twaCwh0eg2a9cSvwZUsC34HDALy/9fUzfKt8WWqOx3yXgnfdj7JD6
EIU0Gc14uYH4T2HVm7UtamWGZWOZV8rDwALK19Mm9tbYXPrZftUSj/vOCgzgiVg3QGtySXnw9u6S
YdqvdR0T6haqjaq706zcSGeQUruB6VZYRhbEpbWRzmlzrY5FsPWVL3gBlwj0SNTi6Ws1eHTbBjFF
Kyf5GAsze5XIjUS2RXV3zJU+TlyJ2iBrxZdvTp33MeW04trRNayZu4afs3JUC0GYHFiaBJOW1IkP
FMvRTxUjYaMb7R0PTqUidxw2AoMNqGcO5i2diXuFc8g8cIHkCNKbysc7VEJQOikO5mr76J0u0/gN
uBjM339v7LEyAlwerJnLRgbgsRPIacwYAMDuxhedqVBJlKnfgjMSwfCqTULEKd1kLr4RcaJGk4NP
cOXreoMHfaYuG/YeIw5xHLgur1fWLvZdHhO7nkMpExNN4PBp+0E7xnCbf/97VTrloqES9uFJDBzd
TL1nDKyrA5ZK3okXLrdoqrUHL5Rlya+T2lBoYh46YbJ3narpzKcGMYKCFhjWAcXqIZonQP2yChgD
Fe2qBDxDO67biy0wTqxDOQpGfzUJ0E3FlHhaRkfnHQPbrThA3TBJ/G2FKeCu1H24aRt2jjcQsMYl
GqGA1Th4hua9sNkYXMruwq8e1WSRqHbH8tb8c1Qrx976mFLcXuehbBqtNquK+mdgZ3rfT4nOwZuF
4VlAi2XqJd9h/ADfX87iIYCN1/bC7yjDeCzhKPvRA82gwj0GYQmo8tso8gxEw0JvVoJPsMeQlTN1
n5Bsv8CeCcKYemjI+HJFcjpWQQI2cP1Nj1WRzRW04y5/5mgODXHFL8pLXRMD7KYEA2t0VE3/fL2d
1nEoen69LY79uVoCbR7Ln2knmWhL+dz6TQ6OBM/g7K0nUPQb1Xl4h6OUTIYR5H1PBz+Js68RHO0L
+5B/W74xcJA9ccQwhsM3KAuGvC4DlHrl8nkR5ZF+YlzdsI9G5aDBsx8P65Qrm9FYQ1J4Kvppyxuu
IH+Ud1uQxR+kECEaM8Md0oTHLfAbY/sq1EVOAUQQHdD7rsNhZYQRuLzgn7OAcNdD3mN5S7VC5oVa
N3Tp26qJt7eU8HRIEGFNjMXAagpXDDMeWbqCN47N38ExeQDJe4jgmcVd2Zgv6+ZmkkFm/fJdy2Tf
cdxuOsi8nb3vGVRliTf/jDbyH4cbboUVCUFyMv0NPNk8xO1jDCfU2cfD4kmRTh3Ik4Lf7q+krVfY
NTlrR1/8vukKMIGo9vOsD+7I3n6Op2rmJ9Sp/nT6TRGE1nxyT07a99V7ZeT8Vqy02qh/ugo6b99x
w/YD6+7E0rC7nEbEAWxfA7/SCdsRmXx/5lt8hVAgA64WP/Oj5tYCYT0AIMpxgb8ez+uozy63B69w
2lGDFvdyfQITiRJOovTg4D5EWpRxin7khCxErHmEkHMngy/c48gTr/WMb1BV6HS2zgEdqqO35xSv
mCAXscY7o7WRMd6EZcN9vlxICLxrjxDYxHbjVLIz3Upbfn+ORjV2mpH5imHbkl0WKQ5cs3BzKi/K
i7VSV3lsGUJcjbJ7tR3wCbEMSxhkBfj+xT2aTi9X+VqbL8Z9xb71z01QZ1JmuHh18NoeagEYbLvt
psuDgW/kyi+7PFJkdDVLUeOjcicVLg3sWlc2AUQ5RSB7GWz79o31sumR5ou7Kny08GCiAP/Q64mk
pdycTFEIlfnqf9MCx2Hjz2mhKA3UKPMMDdWj+HgZDw84/X1bYl2SZw56C9nJ096q2z8U10sM9G2Y
J3eUEhIVe9I60Z/zvvzTlYf9J+1tshFh6Qy+wcX4Av4CJ34BfO5/ZuYWqBh5FNm2sK7rhkZZCkok
rJDPfyH9dJ5Lg72hoEm1mEA0ASVrvnIuDjL8c2VbkXzccxYNuzFiVVFAox10tuzm637yEt+UacyZ
ibARCvVDSevaDq8gjvVYwdstdyiC0xgzhGglDUvQirnZ98HkwRTvp4zQjeFdAhK28BhTOpWm7fuS
X79tm+RK0vVjhb6q/qPYZUAp2Ers02E2jHGS5tExKKBCMPPVDdevenVMkz+0sXkQgayoM04EZ4PQ
OQdGKSfrm53iaV2XyWPdvRmVXnQr8xeduA8X2DcGILlLvEfkeOPTu/P163dLx0g/9Oz1JaQt7JUU
g23lIASW3Mgu0mmDcnmcMKbWpBwWscEQ280vdtIAkBntCquPpB7Q7SuYP0/dX0I18+I9Jl6QtBDU
txJEcwkP96AIrudVfUwxP9GOHR1jA62g5Y6COoIZuZQuMyddSth7WVIe1UHbe1IHkEVeeQ5dZZI3
k26WE8D7UYZ3XQvSv8AEaxgq+ksdXFtryHSRw+TSBei8bZv166WwIcMUJxyck21wOZ//AjePHGzQ
bgBfQDsdgUTW+HTd+keyRqfNu0blefSwZvV7d3B6khFGCJaBd2ssv7oV5H8UA/ENW9K6DM/StNrl
08RgsCjXJ0MjP0RMU7X2b//EfjvdnraQVKVzWzW6JAmOOkF52H5HzkPO1eoOphpkVGsnlGYIoX/V
aKTl7L/I7sFcdr0uRFar0ge6Fztx/bV20wgwbLka43/swxveko/MU596F5pWdgHpWJLKC9Wzwlfa
zVaWh0ZYkvpe3OWjEGxiswYxKPy9cfZ1/EqngD15coM8w7k2bi3wkjUm/S7gU1BRUyeWJLo5oFAm
p1PaW97Tk3WwDHjvZNDLaRr6T+pnVBe18+444jUioxIXg+1PYMs+2uESpe39Hxc4mLud/OG2Q/wk
jESY7DV20GBd73ghrs9A1GPJbLyrKm2PYr1Ms8c3v8PrpO/RPZRfLIqRYylkp1+8HP/H/yNindtQ
AimnUXozkV62mNgCf3OP+ta1uE7IGf2NVp7ojrhffP7TUobhoGBZQncNS9HodOA64C0rJXMTsKu7
FCson6tZN33Xn8zv8gwjh51SyecjFjoUWDwsl2THQqlr6aYA6OtVn7pS+2v4yT0EkhHxjYtu1Esj
Rw4998hKGhlmdZXhb0z+lYHG/GZIZP/aQuF64iVLznt/MzN+iWsncVvPY470OAQmPYgVgPBcfkd9
vffAzvbaY6NlOMJLbEY8jkAZavj502uF7y5lVWXuH4oX8FZFKDQxs6yXoYNwZUbMmM3wpLT1cl5N
uzv/mRMOUTBnQUOLlH7FvLErfuGWrpsR9ZOtk9kT+wgMsqRQxpB5m47y7/fWLAUljtnMto/h5ktX
L0GwYOZ2P+VdRlKW9Gf1+OciInco0Nz9ubKuChmZWTHxnLEHrTqbs3DnjpMeczj8eyffD/eJ6HH2
CTHlW8zd/k2ZFiQQ7BAIKUhNDDIkDq1RX4YLy3iHzCkszmhI+IUXZ3hNY+7U2oig7y9QG7Y7oski
y00j43eXXC5utorxEv2oC//ym3ZlziieoXc1IwVzzANWLxDjZUmrHm2lu4gFYZ7XI8xItyCnrUES
rp7BzjcoiXdaE963FbACOGbh8Eu3JlzJ0pnm8mbd3QwfKdP/WQUivetVKxlV2POU7zvLIIRM3Gzq
Tq4rKr66lSJo+7ZPKStmEQGKxyj6r0m5u9QFN8T6CR5VmO6teo+YhsbvjjDmosnGKAWUbQcXLaZm
0oo0a0xqEA+vB4Dt0IosjeH64wkvx64lbrpUwbBZZLTwNGsYH/uxGg2TZvqOCAXy62/mVg7OBv7J
ZCgnV6+rwKl9prd5f66fkf9FOT7V8dJ3v9FSZzO7fNPJXaQdEYoIqwn9neCMoAhzHgqhXlRi9WKT
BDxXpKVz+5q6V9OLF/GcAZUd6s8TSZWO9nw9KOiK9d3oxiGLkszzSMDgTpgjQ2HnX0EZtrMJmDH/
t/zw8y+kYShmMI4IqASQy5QjfXTMylzo8nR4GIe3yiZ9aKHuzTF0S53eOxuuluRj/gxGcTM6snod
GsQqdzcH6pTDOoYIF2dokn8SkT7iDmFDsgtiUJR3ly51WWtmc1g5SbOUg7S/6AjHhBBipbiuQtmL
MUw1CZieJ+tIypiJ7i+INcLK65Mv0WTktdLUBb+68jZ5mNCDF8QkLfnzDD+l9LL+5HZXagzd2QIP
WpmGuKq7CE84WASBXh2HdVHug916On0nYTNDPc+zuzPvSI60ZLyiWvqkioZB6GUw20W5WvKJzh7+
KD5YLt4R6FZgZxCccbCXqH9b+Kb5ICWnsP3G1TA9ovyyr2lESuCld2Aih/hb0zVkApV2W9Hr6xT5
auqFQMWWoVwlK1aD1y2v/6SS44JVVG7xHHjCpaLD3r/QlNg0kLz/aehSd9slPnFGNFtsQIaWPTpM
ZsvWenEWyiGuwq/lACa556jBjTCoietpn6lNHhx3+0ojIoF1B4ccLZQ4dNyqcHXPSyGrcekZJjwL
SEF6bEfBrB0RuVFANVeCm0G2oZn/pV/LcV8mxi9IeEddF26yO6/BwW6CtE+38anc5/+O24IDp3am
ZrGw3aIxgQmaWN603XioWh9kj7po0Z0hBonwjgYi5+s/HqeehAFGGbJxw0vlgFQv7WijrzgIL/KI
ctWNpY44NL7lyP6ZDeqTC16Dwup5FeUOrrWkp4HeVG7EkgCrOzwcX1e1Ggibghzrli1fDV54pb23
RMUrZ75lkQYgk1xQi1fknwWkZNeiOYJKsGkIK4TLDm5VjAsCDGSahblFB4uMLtcmXn8TsuHcvYGJ
CFRa3WrlJau/l3QFVDBDwnh+PleesZCW8/D9k8fLgJTvQohZxk+qcaeHljv+uVxZDt0qOvu79fNF
ZVSz+Ro16WDOl2nhSlqIocYMP5N5s5prPDDPzmoo64AK7hgce6WAWBBLgtqNGLQEZAQszHyuQnLg
J4YW7acIM8JU1e9pgbMoLbBfrKojVLriMHS+qWiHy/ItguI1sGLhw3z8LjoP2fMcDNSdau1p5RTF
/lPpc3ism6vWM6Pj0kyPxFqimCIJUys9WrpM7v8VnybaTaQPZtTj8Pff39vLDP2t3ufoxl8o3mmU
Hi55nyRZe1Q+JXn2fc447Rufvio+rnm+J1WNVyYNuqqn90dFrVOdZFijNgw7lWrEsmPVgWVCEtQn
nnUQKrUk4a1b1PSwPGoB0y+nn5hK3Kp5ni8p/qbww0SaWFkbJQL6eT9LPlKQ2LvO6MBNYSR8Berx
qlhxM/TmDF1lVz+L1iuk62uQg38PWslod5/nUxvq/jyllJ7QspAlv7r3i1tWOhdjuAU12FC+Brh0
+CwbxmS38tKACpF0yue7vkaRaoTX+pokvFQ10q48plZQwaDHEoTMRkEFS7K2MbIXm4k2aFX9nOnD
hawXQpwvc4ky2ZdLBEzhFLbjEQqskbsXI2xWccAOPl2TZ2lhVKME/GqjDlNuP9mbOBjndScF2Lb3
+SjY9moe/dlU8jtGWDYJqjN/2AySBziodrOmps5GROtJVgOOEp8QRgHNTyUBp3v743TGLsp8J+ew
0rncA2RHcXBD8ip5F4odCF+PjffzNypELdzvFNlgwAdYCr+sIffGX55hUVOQulzJ0lVlsnbXJQIE
4qRy1eCN/aJHUV2YdLrreUT/vRBQmTxAMLOMtjd66ZEbv0zOaJ57ORLnjM3oGpvyus7UFEa40wd0
oFuyekw8Hkmgk/LbZFFNSfalbprhfVKs77SDB6XyLKwoRonjWg+TAtbRT/YBUMDHzVDH69hKfYc8
TWSJXkpBLFkcW/+bsqMkYvHgwaOwUCd9HFQSXxQ/OvAsGerE9VW4wjgDZ29JBIa4XADqzul1CEWB
r4+MFUEm/dTD/V9hUUqmM5KZJ7COufbyQBpiKJEzW9mNglHC/LRshV0NUSgCz+GZRVcM0gMbTI/f
vhZztCnvIeQQH7KsuEDQdAP35gwqr2tEKkNNrpV9eGbMgdPI0r95pLexJOatmdFDV3EBIFGRL9xt
0dpRM+93sBkIQFOoqtfzzxnvJGA8Gy+VFHi5MJuCn9WstTN3tTOtKBuff3/A4UoeWwnq+6XvSI1p
WZqpBvQfZVCtkgEE9PRoGEIf35xWqBRAhTtDn7033Y8BvCOOKvCvd8OHS1TUN1da+QbEq2/pphoA
ST1mi0+wPEt4GRWS0eYYUL0bYZYEhgE2xVF4VeA3tDoRkRqB/8Awd80QfsWCSypAzX1835cx55gz
03C7iyXv4//6zuoh08E/Um+/495xqu3bY33mpmMA5rN3imamocWFt2ijzUEJRbfMphhTU4MbnWla
T5Ywh2j3l1FuALi2aCmXE7P8uRR1Tm02LL7t/3giU8J5xKoCqd30597Y92ImPpw54eLHsbcFk8Tf
jFHXHIYmBiJ0Mo6jtq74bvsMcV7yby2Dv59q4rUqUEIEAn8RcUKsaLHDoIAlZ7+XS554R3JAI+nZ
D8UP67ztr0pIPd3P50toRdT6+2XrBzdIgPwwWHYNlu/jCzjYz50FyK+6nMvQkD2i1bMgaH8V10Jh
adcWWC2CB+bM5G9wQwuBou2lisUphayzmBCs3RpaZp+RhcOHVUH2852MlwAThEpVBGgXC1jt1rSj
4vsnhiP/f+0NHGEK4McLFYs/EXc4tKAnoCM8xoN1A8mZ1hA538JStD9zimxKCI4SxoQDAGD8IQOE
42vM20rKsrHWoBw2MbwMIV3kQCdCz4F94c6X3Xxzjuvb3TqvyxSL7qAz56EjWuuRWN5hIoB9Uncx
zbIJ5qt6j2eS5h/pCTwPn7QmmXVSgmFEnBC3OvG68Tq86DQwufh0OAz/MU/LNxEb7nFh8KiOGqJO
b00+2DqdgA98qamZT/TCeAS5ZvKt9YvLruylqf9ay0b1kE/1ANCKli0Cjy3rJHJ96PyHljG+Uju5
I+RnSrvD2I1wRSas3emRF3qBU8QgAtSgsnq1Optkf+dvU71uG0G1TcFkJW/Ig7b/HpFhNCW3lwrF
St4pZiKaEM68G9K7RwNw8iuIwRU7HbTmTRHh0W9XIRlMlJ9b8B430LjMO36MfK0HG++kL9dq6Lmr
NfgQ6NpKntk4q41g1IhomOvBRhZxQKMV6SthslB2nPgbqrWPDgPwKj+3/P39Vd1novgV8AtTl8bt
KV0Y1YtOWpBGpFumx0hVJ5Y/nsiLMOY80cHd1sXChQ7l0GyTq/lRgecmR5+2GwlS21wHMF0EsV9a
/1igWHE6EJ+G8A8G3dBv5cZXcw5DU+54trmHaCASYSC/LWib4zQseVMOwpwDFiy3b4rQQiYdpI2l
yGuOM1Onm+aZ0Czx3gHbvalvd53s/FhxnBaqIucPZ86ALVdN2+cw2vPCEs1PrKn88oRDrQZJra5a
69ROTXceGpYaq3+y+cvR4SvEluUo07GslpiWKxMnYIawo9zBK8hPwXO2pdH/xxz+CVrfgzUazUlf
dqcjHEnaVHvo7grf9K4vcz+/5M+6+TdaUe6/lmRQzU1Bfnc2SGqeeOtWG5mb2iwb5m16yyU8TPqw
D1Stt0y2pRrmmk9+8ilNq3sSr5V63T0wfe9solsQ2vNVszvIegnbBvtyUro6tgkGUJO2It0yFAnR
AzmVP6/Lnbybv/5JAloN1YCmG4p02p9IIsq1m/yYlQJ3FL+wuvuduAN3uWFrh9dykzANK+lZ1ZAe
xEhxfZDxNRJo5cv5BAVGZ6KJFU0MU18q7XrjQfy2O+qsAIPtZ2iSxvDC31VVEXZhtTeWFVPQcODz
kwSJFKVHqRL0iKaprGWjS01DM5LoGRkaxWJZ0OgWfamv8JbGXryIZH1WybQwVsdSP3tTRxGElNHx
DWpbesO7j1rY/5C7FgkRXxCjxlTXAExEL6mTIDhstnSQR0QIoG2I0vPmOhfmMRlGnKLcT/i/GTwO
+GdEfL9lVducL5CdE8s1CBu27nOhwkClaYzGJOCevKI0z5po3hryEPS28Cfn//OAIfPfKKernBRm
c0QmThPK4vwoSCLTGauGBNahCwbY1b6NDM94y+8zr5XyOAFnGYx2Cdd2KpdXgGX/MYhrq9ZyquC2
pA13RasAk6bTs1RNlu8GVfpWCOCeeYbXKRlGJQT/I6BogKnc8iRPPi1GmDR/pY8tqJ1pWYUkZkNz
deJs6Q2z0ocFxqxbioyk6LsKauDmLjYcrUyKrkSdMw2MgEiXOJfIVba1cVKKJ9O45LeWFKz9xFGK
stpDa2JfrzH8ZWZkDutyDocwt41SFKVxx4qK0ezV+DYY5EWKfCBtf2xyO+Bi+fgztML0pFFn/ZQf
1FiSkqHh4TZo1lgQjV386x1DsYoooIIroJQ6rcPZhpABn9tqUY/rvaJrqHoNhQQET+Kf1SsiK4qV
xYjrYGh81Jt4rOK0jp5dIgzPy8eIdOo9DKgjTWzz1x+mv/2R0yGHIb8Dq/KG2prVIEkFTJ8YBYz8
8A9V+8k9UU0375Ja4J/waUtKoqYfJW8VT6cRyS/nxxJ0m1EKQ88H0hJ63pIjXGNEnDvrGeul7yur
06qrgf21BU4v/aYTiuzoq+7uRjBYGTfTzHhzF1Bnz0PhPJIuNyX8xpDf09Jya914o120cihqerTu
Vk7mMKUo1q37oHH9D/UmwW5Sla9A4zCEicf9PKVA+n/F2wEGV9cUnvcROkJMxxJmDxQqLPdUWIo8
aQxjcncb/rsNlGFIjTmEgRbI1gQrUy8eBSVQMlqZ3TYJyfpK1dtDsTaWhUa2udrrKCs/zXzKEuZQ
QgBHH+clBRocL+76DOYV4IfJFMDfnFG28HHn+J5Bu97JQe8RM8F5tXsbTDMppBG5aAhdFwirkUxF
DT/8QDER9U1/nSLMaafBZD8rI5duhznzjE/KHL5Y6jkHaYrMy+eySRNmtHrXi0oopvke0ZYqFzvV
HkCd4WFYEnPvq9QH44/CFkQaE2tP8KXFJlpcrDpUjPUy3pUUttwGhe+YfOcQ/NLIKLtg9ZT5HGEC
owoK5wIgUlyEi+8fE3UsHIMff+QeAnUcjSPm++ZWwADLmLbeNZRhM+RFGlhE3uSRhEto5VGX/dq2
/MQ7tcXYtt3ApN/nYCsZH2g/e7FmjUmIziBkByrdO4mG6922jJfsef+xCxoO2PCL7rhPgVMNICZS
xEt4g8ggmf1mFSkmrfHhQPrkZiqh6KlFaDumJfDosbHLTfNpPSqLSx3c2YORdDFO+LyxN/G3KRSK
6N/W5vHUm5r/06g4BxPe+A6cx6oJx3tIJ0JBwckjrMsxsHxh5UUqel1v1mem5QfK1say5jXRoAnR
QcvraSpOW3mKHRJGa2U+cSse4ZaTTOUPab5Z5kvVvfwVtZS43gO4AEs4eBVbrLLqF8udPEzklqNu
ceOdRiNBKPi7OR6ZQb/UrfqFEn7+++5YYiBkwkfuvnfXMrK2IeP4lGLLg9AskR5AK5wIDsi4HcR0
cW0GoeEppSOe80TALgDfhLngZMAANu2Q/XUXaQRpH+7TOyL6shspzVYQIfZmdTKleWlGSMeL6rAd
wdJOYufpx5siBOuiD7pstiZ24MhJtX+JhX1/BnSg031gzyXu9e3cW3ugBsBX9+Bh0ZAtxrxxjjtt
TdGrVGRPWjq4kxtgBJGEAydUyCLzbrYw/M4dPo0jRda0T+A89qcrW/u2sAxk/+gpPDsEU50ptnT4
jl6Rw8xviXLsdcwCG84WibgVEg2exxwVchIxzzvatrL3ew9yWSEZzMPKUSfPQce3PhzxSYRj6jbf
lajSEGM09rkM6LT+/W8QlrBcdM/OakSqdb0QKyPgJ+a0JraJeY2Q/0KZ48CZIu9q6uLhq4BGYpk3
24ZQLkLpAziS+9Hi+BPJNv0sJC3MgPupsxVT5vfeSQvz6kWw0LSOwvEtkeIcUky50tQ/l+mGA40C
0EmxGNqV0XBx14WlpBtHGOgFrZ3pX5Qzi33f3yyc8NYhPQeCbeWWXqJcJw2FOEtW/2lCOMIT9bBY
Vrf2XwGPCwqVsF/A4CPej4l8yYG4cW93HtWBe0EGRVRANTvgfrRwmMPmbLWZSCGnjeyTMNVH+65m
cdW7Dd79wDsoLOlWQB6jrVEZOn68aXDSOZuUVFSRyhkZqrWZfOyJRakhSkjHoGLOUSjH2eNx11+g
ChYR/PFPw9dfUAGoav1pQKc0HsPxS/lQesumTr4uCMEg87sQ/a7CRuoHQsZcs4MhyzhRgJk6RiC0
NsUVVPcf93dLYr6nAp7WjW8X3ekQdLIHnRONf8MP/QvBLfcanwltxlfdlkUGwRZSkVCXGOkzj9Jc
6Gg4b72cn+AtkIdJbtiXlT8NcPVaH7zLHqrulNsQTRN1cw/oNFvj2sDBZAZ+fUuj19KCcX3x1p2p
mmcFbjLehs1WhBRdTfvUpXqyKqHBsFM+TP5aq/Zku1qE0pXT6ulcueiZj/gdwIS00AwJ869tQPvf
eqRiEGuO4sN4MK04tWOPyasAWJsyvZmNptFa0skXuBu3IDkK+sovLtRgISbC0+DfhDjr96CitOn7
1ImBoUZb98mOhz5H8RfMfCCo0imq40NTZv7MTsBuR8+EZ0OhqywOyeoTw1oH/aKSnsfaUL7652Qp
MaAyOsCO9+BROZLJRS1VRbUi6BO3xPlygb3hync0QgGxdudReZAzpQk103Btm32bjTzeXAUVQM14
0Ms9ktLayiCLFZGZatFXJtNng8Dc69qNykBhCOixXIbMANtFDhlEts+qJBE1B2+zcF+E8Xsb1AwH
WdDq1gh+WFKVpxCPiWNHgEZrwaf527/eP6EyQy4BVrNBMkJHotbLx8Pkfbr5Sf7i/x29fN1NAsjY
csNCrz1rRhz32dqPYioertFnRnYv372WTgvIoVkJDmE7odvTfTLtZ6ZL2CuKSwdBwwfGZHY3MnW7
viiOoSiQ6dsM86405GTdOfbTQFmi+rTRTxey1HYhbNyVKApYWv/GAAXtykKE/RZv8h4Z3lOHpIiZ
eIhZmKDuaCkPmwP3lJ1cqCwrOKRRLeGBv3ue7ukhniYqXfyfDIt/HLt9TBKA4kkmsGWInInrR4+8
4MAVEKzcKGbkznImq3QzeZRWpWxzP+AHKkCYExJq6Xs/fvMb7RBDMXvQjiuUfYNHI+lz5uO5wAIT
6sdYchHpG6qAkhtPPgTUfGNi4DD6i284QaRV4DO6Nk+eWuv/bVQgv47VRUfrxFzFrASwLTyURMhk
4ggArmyjR0KUpDHn9v0nXj8FNlpGmYWrKH5mEyiqjSWk/nuJR+doBvULVYIZjCpiN8mSzEY5dAHd
oaplTIi/ZClEq91GI6xoowoLJSm7araG2jhdwJVkuCBkImsJIuzPQdDk3VfiQkL1Pn4OArrvQEK2
OHAcmvtVhyN3Nke0E1xIBavo2u//QbF+gfkDHHKxFHFXDJG89JszPN97JuKL5/ywTariEAoq6mov
hrkgd0u6qFzLYXdk9nGu3i7j6Wr/PDbw1cp2/nFDAmdmVXAO6Nxm0jBVJfbNtmKBMB0FnOFunSCF
P5+x5Xsf/W46e6FFE1TQ/X6KXy3hJBMx2bGtB8bMO1xpHKxpx2h078cTaT0fSewHO2R+H0g+XRCK
gWCm7xC68yJP9SxBMNVxJQGfAnyUAviOg9Sx50/tGLgyE9kV+aUP3ufVAvGR8Aw81cvGegMWB/A8
uoR6JcwxWa3Ru33dAB9n7qygY+EdbBl1HXSoVCqgpLxG7MXPTr/5ohJS6Yu1eW7IgcqAedvLB/Iz
lqJAyGj+okkY1aAWk5/EuM9j2rXkbOzj3e1QQaApyQD8pYpFfijBioOU3NC6yW2GpZXcSd/zBZDD
ZQ2IufTHEaX0K1HqJKuCoTZoCofnUWb+KZfFkoyC/yjRyRlxi/m5N+JQh3AO234yFqArOAvmTeR1
fHvj0PpwBFxyLJp5d4Xm/xy68fIcfVeM/tbbJXzq0LNw+GzuW/+/FwG7ZmNjGAcEuBGjGpZ3ivsD
TAyegIyZ+VIWRzrKQP59ofg3TbyLE3B8zFynZF/7OFZVJueGdcLmxXHcUZVcp/CU0YKuSdjlsR2S
/7aQwUut6roTwh4+Gff4ZoKAlPBMugHyqlWDxlL+ZSLDGPOJ57YOjykLH+uaTPXKuii9wBLofXiM
uZiwOcv6abZyrM7abYgxqRw5Cino6c2ZKfLKG7R6fTWsvxXGhEjZqTe4e5J/9OAaTpEz+3jQMeC+
8gKh/2HuWcv0Cy4CILAzfyaNN9bpzcMSIPdb+PjlML7imZ4rvM6QesVYN3p2yWJYBXmytkWmJe/L
OL5UYBNbCIhy6HMah0Opt4hKWEf0ui56untCU/tbtVQVTbtOSr2MVeV1VXcdGbH7u7jRgfbmmTaS
lP/lm1vMsoLqJK/dtVC5YXBCBM2XMt76YF4mMNqR3n8JDsHYNPU1MZCrmTTaiG9FAXaf7ul9lIYu
KVN6wiCHZOosnhkqBLY0YwHrrL3PJaOa8hFcRmAulodpvs/PlIRyB31cA4ijH/8AFEbDFkMK/XKW
XkB10ps8s37e35c9H3ZdUug/rngecpANjBfv4Dzctci9CbA9QJTq+72L46xkWppDaJY2I2uCQ3C+
7gQa1eqZRo8MR8W79GG0B3YwwbbMC24k/iZonil9g1ikvQdvK4q0TJRHBoOwLsdr+ZTwufALhKAW
84Jjlwjb8Hw5odNQEzsESII6mX4HUsQBJhJEb8+iWBprExswFTHuPoraXRCKlCLV/KIx4FzKFd7A
qW4pjDg9K7yTH0uE1594ABfpqmlScax9SMY7iou7E31ffJZimBnJsi3dvtIPvrfDojfve0+HmDy2
xtfN5ks88p25EgXZtYX6zFC+MWhtsfVOXho7Y3EsvYskdZf2RDKC60M2juAqa/mkAM1Jxmig2iC5
9LAAtLQfyC3uNY5rTRFin7bc/C5vdAITtMpA9bDzsJ625LxlSAT5LAau0gxq6D2WVLIT1LRA/+2c
HaOC0PzhnnWLJpeEk7Si/Qu3TzcNtlhD/dEjeN4F0imcnaV25wSc8NtaOTc/EeflEXqH5h5tA5G5
Guj+A/2cCvxq9qM2GwA/eGgEoqBcE1BFOQb0c1VOe7B37L4oy+cYnBQZ5SG/ALWddnv16hALIlqW
1ATxM9a6xK33fhV8z8YgQmRcirJnZSNEXj0NghW/Gl/rMREvYCFagZpdSR/P1w8UrnSn1LeFmK36
kJIAe/Ymcy+4plZu9evdX9Ck7DdbRqiGxWMFn1BY6n7QTygoR/643yyPFVu/g8DAnZxtN6OszH6Z
/CzZzdPY72Z6+vCngIQ787lfM+TnTias2Pr50O+pQX+kFI2FZPImqOUh4+J+gYnANyzrV4gtn54G
LnNWBeAz+1NCasCIqf0S0RG4RPa1QjshXKR/aMvkzr6NEgYzl/6ZVRmwD6lR7AkFiFpHkQdp9RW4
IVpPhDkcjTHyWmxNBnCEUZQzSlAg/oto336mVBocp6QrJo3wgC4QTFOm1DVhDermBgM7zS6P2sNQ
63Mq5hfAAmovk3PqQvQb48a1ZQ42Db7TeN3Q2PpaAXhJ6WgMdAFPtl2BZVCPU0D23hst25AyWg9l
mkD9km1BA/ckuBPvK8CslAgbqlstzGuO3M0N1VlMO28fRuCrnbjCzZXfCGhLSzJFNRdO41jQ/G4P
47fN9YeEViwycHMDYV95q6ctCtjFJuqV1f+Mq1PtUWVioVNjn1Cbos4QbtqnjvbMhLqgb5qCXUNB
Z0i/54bEN0LsNqNxl8oN0Lk8j+qjqsLBoCFFWD58XEBqggcs0tOWO3ajyPyxP9JlnOqkd+LzX0ys
rhp+E8WfqA2goQAPscAP3ABKs8tepJq3g8yyZTQxeEEUHBI6xQ1fgHkpH5VhtWH3FxoEeBWyzR57
0Hl+8sxS/O8JJ998i0525tT13Kxo+ZzzyP4cS1/L9wYlDmOvyIXR1reEMvfIEgijXqQK35hW75vX
KV/MkwMgK0YieavqH8TbeyYhvZJ+U5ovS/2fg4FUYpJ9/jiHVMXAGiRhh9ZgH1TJ5He13wyLtjHK
soqnjyoZu6M5xFucQvisituA7bZnTwYbMJ3dZ7KRRGPh/LHAKOmL4oqb7D3NHrunz0LLvETj66jk
2+bL6Qyu511CLJZc9TOQtsFaO/76EU5prlmOyGHqIW/bJo5UZATGrkwoxW96OIgNKx6p+WP1+6Dh
KnlZq4z6hat6s/lYPbH7euzp115vAijw4+bnupM7RwbZ3uGw7AFPvn1tjvxEveVfdYjOxmaGe8lK
IqOm1M9jimGNKWbMyGyGNvRJQDIVKKVD/mCrbYZUm+I6SxZ5/mUDV3qq5e0139mhcm3hU8jI340D
MG6zqlkg/ilbEry2DL13WynQWXWiDYxSe9p0BLyCp8vCprFt3Fz4gfxLDD1nzq+VVy5KbyU5vXmW
1iboWNMt/4alxhnFafskIru4oTizvjODORL1RqP20XBAIDAFhkAPwfVgxo8pw36qsBcDp/ZqnZLp
mVfSQs9ETfFz7nhqiFV/Kae77WqavOlQNrftg56I1L/IsG2kW1w30OcLvhI7ogCLhxS9V4y0elzM
/2J/VhubVGOEerJ402BDdJhEtyhcZWGHl1DStP0iDHtdU1hNAfOrULAUKNYyj0tDQdbRPqX3MEYy
wVTck+O+/LKZjew64KfMslk9LohkZa8gKN3nwrDuuq6IM07ZHZXOHkN0AEpJBNTAYH84ML/TZOea
pfyMqgMHU3njBJwvOYGMhsFURmzclQRks5biAff0Fnyq6gSrthiO2taz+ObA/99MV/IsmBVLT5O6
XzTE7iVXEXE88eKbv9b/0gZeKrHrbjaM1EqUXdB79NQnrzsRb6ZGkEldxR1zwyjRO3Rcqzs6MezL
iNjEwKuAZX6xSlAW5Lz72ZWwS04hrMUVJoQ5bdXp8+3dLHOw8zzRTNje/r34AzRMTRgOiRf4CBIH
T7F6FAAJvea3Ne13CoO2ubQDosTWt8FD7JNVyfpdgkyYDQ+WysV4adfc8XerEDTBATppfEGgpC0T
rtf0hUrcoHrIMYoerFUj06ylSA3D/x6Vmyw0iKpS658ZgR7KW2Y5xeqQGk4OGhnNL5dr04oblnKD
xzwjNBIItpUo7BZoM2o1lLZcMKTzh5ZHk6cq39GE4NTb2e7BxQ9SCnB97aDaTCrCusjM9S3IR9Y1
I3ulqFWDhghpkyUKGCjmr6YIEjagDcEF5mCCBoExjeRplbfse2iDcak5fgJ0HyfHeYRse6fYMnwX
KCqhBFAJoAIZJ1AA/555T8OQ38cDLGgFHM5HeCiZdToRyYlYHrRqASlhqybJlUtqQ8DADdQ6ERH4
yc0uGolwocpfsUI2XfuT4jaoiuASUgAGBQd6vb3d/Rx2vOuRZDB9XX8+W0vV8VjI1aF2km6IgE+u
io7oTQWtfWHUzn0jeLpDpsZZA1DaY+GMIhE2bPueX2yvtuygY4a5yl3O/PD2L4lwkHKIr/dLH5tg
k7ugD2Xbp5tFYfwg2NhEpWPPjWXHhwhlkHngEtw+q2A1NrV/PYcWzTJoNDjrHzmRFtKJeFB3DAp5
Od0Zh0TJekVoMbXy0idorooRUM1lttSHS7gknl1NeSoTLoIraTl6xE0QgIt66qr8rzLn2w9Njra6
hBnTI7OzLJjE8SMMizZTHuVQOZQyQAgbSY5uV6Q5OsiRxDnYvNXHE7akXoRTM32LbwLzYo8HpFoA
DdcU7n8bMt043rjg2UIGgsacd/kfmYEbtd+tvXnTyVfOyQoo/4B0gHisrgHw0ftaXZX7iufchZsq
7R4t/E1pXuxgvpUTNJnPKZToTq9uVh6ZeReQrVfvdBGhtekN6VwhxiOHZeHjwMxbAZj9i4uNp5hd
1rx8qP/YbY1zdomBbcmIhBxXnwbx8td77KNr+rltjkY9ahtyqp3IgNg2gZy9YidpW1sMaaMf5qZe
RgZRRi9yiYdU3a+QcL8XWkE4qLjUBz/bFeODInGiER1xSDOHB1BfMkC+HF1CW1fulB87pidmcyWp
UPPIgIuvRAYzo3WWv4gN8pplpgJBAC0YZE1u0Bz/PNw6QA1ZdhppaA7g5bA/Ig9YKKPZmHHVT74o
+Q2VsbsMTPJJC4Xmx6tv0HcqGRTyV5agA8Fc3Mza1Gy5jDPvXkyEgJTnlJT2mpgLBaLOh1ratFE2
F4X9QUJ1hMw1a+7anptn0hCNfZAMnkHovJONlu0Jl7wY1JteLhMIvtZ4ggGhoaL+We7UOrst/E2g
QruA62sgscyHlcgzRq6tsMi55/ERGcCPKmpluANHMwoqpyBTmumWBpunxcAq2PlnlZxklHFtNZHf
kYpt53TqT+QvQQr0k6Dg5yAKX01mDgEtWRK//UdUYLz8P+A6VuKW62hSe4QX56cD+Cy7XpOJghAh
sebREXJy4WvXpv+SFZ+rASGcAXEOWLvwpDvBwLG+3YcEZjI/VuVEQ4Jp5ryqnxVbP71rLqLeXOlY
Tzp83gZD6qMNatc9fxDcF84+F72bd/Fa7+3f1ZL/psXY3NtyjqkjXj84d3aa345qIyzQrLzDJs3o
v7TjUtsPN0WPVUPbcWCTPHGhLVoNU3bUs8PudNRZpQLAEqy8WiJ7CyGrWadFjbhgxLW4u7Ajw2gF
B5llkIbkVu5F1rLp0NS64hp8IPU5D1mzT+ohJ0HerNkvavpc6/2/Zv2tFmE7NlLHQelRXA7IncVx
HPo2bhFZp3Gx1ubtylGIfexVaj7F8xrD3k6G7fmahTZt3lIS+XpSAPnrjUFPv3lwoqIaG2jLbu2W
cAqvjQOykm0RgY1HCTq8N4HJ+1fnlv7XU25XNRXqUS4+WfBKKYUc4H8vErF8fVEm6R/PDoM0EgHq
s+RjEE5tuSeoEtFf2Q1rehg5HMMNcKHA2sRMdGK9+nge4X4sak1ApJ8DzyfLJgEzfQ5EoOOqFLZ1
o6Uw3pN9R9AMkCKoyVhkCQwq+UhQHrz7RglabdJTZN8zHR7ePWC/wOjhZslRj8QX3G/kxid8lLuF
N0ikIhSMaib+OXNA9soLF67qYrV/LSM5I6dectzY340Sxxo9ic/6IiukoW0KSbb6Ka83axr7er4F
Xzt1wKQ3CXJY+c0XnGPToIncn/aPUr7OA7y+H4Ba1X1vpWPPtnWCfMn0mi3lgLOYgnLXtHQK0Rda
HUd10DLE0wODLCoGQByh87oTSlivGASfvqwX4WZyEFwJMQls8IYRcEDR4qQyNV1UukCiPyM1RWlN
Fi80ZPVB8kNnfgGAx2Hg7HSYohY6en9l5SUWcnX5U0DeQNodPDKH6S+CnmSQQKnO/JP5ZGhzMFq6
eyWILEnYd5QmIpelcOjutCdIdaUTck81OK0E+ZjdTUqu9k5rCE6wgySMfz7fdEZfEJhSkT55P1mR
EQ0lBwROcN2Gc6DOhjl6fyL77jTlYS5ubc/PUQcTaVqnEKKzp7TmOFGMhRBtogyYawzQy/mjAfUz
VzRZ9TV8jp6OCZwYLnpi8f4vYT+lSv4H4Fxz+WP3XS+MdGbT1ukkWfxpEFlmNrLz0fORoKvXbF2a
WP3kb11uhpC8AkR9qgLr3bkwSpSEcvnhrTOS3Gp5zp3cswl80GJQRC35W0vXzvny4ArzEtfa8dG9
Gzk9gUCWbVIg/yn6Qe/fxhawfL0Gb6fj2gwZUhlqw4uGcbHwgLUoWjBxxG1mTFcSCnIlbx4ijNRb
7f/5H8RgMa1pkVwGnRooRo5GAAu1+bBHmktxWmlLJWcOABxYsaqiuKAjXJsUvCzjiL9K2UFNPokH
MkcjewpIQspK/U1etDoWIDEaTw3BV3Yn+fNDN6QnIjjwGZAV9It6kHHpuFu0fc1sRjXPDm03DsE/
aV8X4T68mnv6ONUk6Has+Zq98KMz5IhFJIkZZx+Og+ko6vmjyN/yMo9KTS/TgCtTzouX8VijDy7V
/3/qQ7UbjmNkHhxjq38x82VZinfV/Y/84HYgPk38F7A3rcNotkJHRI2voeu78Fy+0vhG9UgkIEwp
o0b2kUx7O947PjHJeHn7uQlRr49sGow2fXSl0ODUzLBZf0+a5Vn2HtyxXA8ELounNsZ1i75WvBgO
nT3FTDCbjfgAI7/wTDVHdlvCH1ZwX4VMu+Oe4hRbw/4yOZT0BpqFFyXtJahXXjt14wHHWI1GOL4M
YSf+VGXKbGIrTnwOjdhYNclvIGxZupY49h7lbT0HPrzUA0Z9moeQyQQjryAjEvH4NyKS5U6bR6ag
JPUzkU7DQl9KjbDpHG73HbvmZYUyu4/xaxu8L34eoMOEUZnqiJwxskbAFpTqM2iAwpDoUpBaB3Wa
8m8BDTmFL6/C8An+gy4/ftu1Dih+HOq6oraOrgkau9sNKh4BZncCpe38VXjxUW/xtwICfIPRk/r5
LKVcgIp2JHRwDIxhgag6vUxUAE8A6syhqDmHCeCQFdz9fJWqRhfpDhNTRPHV8iHayhrf0HDCWBJF
JkleygJK7BtYsGI6bK9HHpiFpucOKRgIs5s8aF533oZmqL2VH94q5sEhhWXvOTaxi6Czf/ZOSGnJ
5VsGBLN2J7yUmY3ii9qq/7KEwR3FmwmN7B51EMB7M6TI+Ui+msJJjlJo3FTcWkt2+9v5FHani8iF
c8QS6VrFPQku3oddI9UjXpiEuMvH/mA6S/rmTQrVidf96j/DxyphNnoqnIW2WGMTkGXrXWPC4zCJ
G1JL/m6LJ0vVkbi34hKdz/QKWM722We6C9pAY9XVF9KUHOg7Fqh45ADnAw+xYCMQJEUaU8OAjxY0
g6GhjUDL9Nxc6+2DI2HHqdaKUkik9c58qP4yVL5FISCmIPlaxjIuf1n6Nm6cgJNTDC8EX49/B8r2
REOgpT50fauKG+eK3gtf9w4dv1QLJ/GT8G77NkNewlPFM4eVHnTjqnADEtUXFaPkSLziyixoGzoE
vwvnJpTnIr1fcEHoxnnwUDKCTDVa3n6N9JbKF1cmx0qlRQ3b2g44ue6kbjKXQah4JJINBT9jlQgi
OPOTmCCezNImltohWjh9PqJQz4hNAsDM1byD9uHKGbtkYPWfmIv2F/+1b7xz6TC10YlyGfTVmJTw
BD0ByOCPFRI5eQ+hBx62hb77ri5g5FUXuEdqdoekCITIz4WkitubR6b8DDq6mvznmzYGJH5VJQee
0hpuLhZkoupoOkBXHSv21bIfEGog04Y/b8EUL9tMS9jdI0I1+TnhYnNXBKSilezWQxQqmJoa1G1W
qtis+SmVGKLwJd0u8PhsPt/qUP159PirkmcULbwch4TP7I/1NrcFC9GBbzKEDGYEPUDAS9qix9D0
KsX4GBXmNV1qY3VhEIy4l6oJBUeY16BRtU+56lDSnoJXV7ZrzJaaBeSyxDMa0ybGMISRIVPFOgwB
zqfdViZsTaaY1JF7ElElMLo91ncT2J8LvZmj+AsQovTZqsoKFP18+96C+X93jPGTGgqoVMqDdorc
ifapOVqxnNlOFsV7eJEstdNi6+xuJv0rAOt7qa0g48S7D47yFxuGSlpvcYQYS/0SpkqHNQv1Nm5A
7ehrfiaONGvVfLbQ4kx4M9UOG7sU+sY7oCwHeY2Xtk+KgIzIapKgmtf4iSoP4db/oIcZWPqRpXeg
LImZhxVsE2KSysUCU87MN5/IFoXVy4+p26uW2x/jbPuXE9coUpBCCT6yWmgmcgzIJYyTUePybLQy
WN1hGtEdolo0guKaFPm2VoS55mdsRfItRTkp+SrhMNEDQfBfiQriyxZFC66a3X2LSpqJEfVJzLzr
7aqCVfB8uHzfTI42NJv+oKJFZ5vIX8bITpvjJvpXDxOpL3rUWUtHB5dLa6u4h2N98+8EBgfDJC+R
YGgGN5mbFvOFuSro7Ha1qQ3Zk7cerBWThOIlFyP4cxz/ogGw7oAZ7TOqZlNL9GkwEZjyUxmQqIkX
1p/DnCcL/iksOkdxZf4ZC/Uo25fJ84tgAs+A5mYRjvmUws7AJUPMJJMR1Y/a+L+AKx3yIOmROOWJ
Sg7Pm2ixnGgbUYfQ6j1yOz6wEofKKFKtNjVd1q8fl+P3HTen6RWTvrMKDZPFAsx+5zhVVWNoPweg
olX+bO6unJU/WxIm+owRpmDkljxY3xBUvOFhqxerMA8Oano78ysGy+ss1nhoAQTf94FXfUYVrnNg
mQHhZjhUr5U1+j7KX1c6AvYQfeGvMVBr+K+sKK2uTU57+NIPpZzbbmPx/g5tTagItrkyf84zR+RI
mos9j0u8Qxar2RXpgwyjRbsXKv0YDyLl/mr0QGsFcZEBnROziWtQvQUpen2rwshuelhwRwQg7xtd
rjgCaBU/T3Adh7d2XKXhIdky0sFnTG1X0Rjrd9r2qUwPebdQMIZGaXBdbu80l3EHnFdjg8pOjnP2
HTvf+vpC9Z2wnuxvvoyqtRV87L1YHonVntlRWcCjmNu6tWWzdT1//Nvr2xerSfW/LVclMapqgriu
mqVOrdtCeAuLFQwzQf1BoZSv9wi6vLJAMLn4TOTh3+h8087U1OoWsLbZPjfLoEPKPJX0GRJnP4X+
qdLYPpfe5Mn6YBU2JAoBCLWoK9PPXTvNviIZNAIh+1eRfrQ3bnAToLwIyXZ+ezHr5cl/t2/Lsv6d
KQUdVOkSGcGxvnUcMHPi/s2VXeE5UhisHX2yMWjXul7+NBC605ab92u8X7RqiROfAmQoBwZRRBx9
oiypYKjCFvg20rBO1otsNillLL5wwNEVwLT381iXx8bga9t9yzWzWQ2sAJTiQzfbFKVgrgZ5ewMY
7E+kTf0BKEeUkwqKEhPCe+jGh8ab9ESd0xapbBV9RA+o2TVzP524N1r/prlgApHqeqqYXBUlkrPX
ozIxCSCvIfzBa23Bg7AFbyX/PiuSgalVa1fb4TtJtk+Sbgsn+Nrg8jaTU30UNVGmqiuPK1Vf0BSC
/8KQ6br2Y0SqWLjX0bWyVXBhWlNEmaTtUErmXRXcpTJz3LHEOlQI5z7zAN9Es59Zl20iud6LkUC5
EccQFXyPMIq5o7zk5HbSx3UwCcAmPG+uy7P86sD7qrKaApBLXs0p7ATl5wXpAEr066w/AO+FlHM+
u9rg5h2WPwnXAFb9l9IS1dPI14V1dDIj7CV4HA/qpi6pkb10O/dLY+QdAxko4hJIufRKToOvJX7b
oPp5QvaBRukIhlBLmwDZYdfmw5426L29yaavfM30PaDBA0v1HgBJtJGleShxIHEDvQ3u4ycI1gdV
zQQ0+2S4vuXv67I+kXccvxzMNxxqC6HXX+KRWzBwPaP+37BLe3a8vG2Wo5vNyIeig8Ys+LcBdeF3
QH7eJSHlVJRV8JNqmkPbySeJFwP0Zos8p+J2FYRzkcKNSFv+hjDAEZQu5MVh1Gb/wU5HCNbepHFK
TQUriq9WV2wAyyiJBplBsOxTijGweE1SWYANEJq40o6AJ5ROI242krB4g2B59CznpV3OSm4zjPL9
Q1HIK6jeSC02uLZA5IgUFv9R2Bz+KZrnA9uLFKiWZezyJQlEK+MoF6iE2l6NCQTU1cJJG++d6gKQ
X21dLAIcGYwbbwf7EDr/9KaVoHVZ+90J89WT7umE0JFofvR5FjwJyKd+2JzG86qF7B3jfoWvpict
OFmRUF4oVGSBB0Tqk3kWalqJA8ZA+24Ksf3WAM9YpUz4XqaokOC5RUioVDxpddlpSWKiVni+tj+e
rYKA8g5tyZ9OR5+gQKW04X+C2oAdH3NPn1/F9VBjTRZikIj0Fs2Be6MGICsYXi9TrREmKxcCkhLC
QTCqleUJEpUaVVKXCFxh1Hs6v3EW8OSx4kjRe/I+8+ZdSnBcgcizWceGEBfoCRLYAefsoqnHmewg
gPbjp3YfsVROSReXb35m2tuRII3/IuPw5zqdALrfMX4OBnj2h0P/X3YddShtFfwRJec/mHGey3Mg
EoS3IYsOu7jGFXeQorrroCWGgCmguJct4K2IJQDY9Gz+EfkMRAdWW1r19t/FFVuh52f01kFnzTy0
m6ybRESV+ePmFOB/KE0YIlO8MYEcZZOu+1AgHpz/v3w8xUC+V9rixvMi4vUmUvZMBM+qbjj5IENU
3ybyTgXa1lAuWdUsGazSlVhRVyv5E2jySszppYBthyrDoISkqKo4TwhjQu/RkDO+GFXoMOp04s2M
kISkksgGBRTwi/1b/zRoKezRuLcbjxnHgEQuWx3pVDxzMffyz1/ICsbXfzt0ujIiK/Ma6oDjHE0m
VcOTlPy8UahN5Y/CyGdt2TNjZ1GMQL/l1sh6vr7KrEZMhpo0yZMezLliHSeOUZNTrohXkk9weqLR
rHjKD5VArEHjKL1SswTz95OlFIbDETeeSxY4btu10anKANp2xyw9q0hLGTBtgfU1yUdsqVwJO9zP
2A/Q2UllT9PcCMIFiixvR2tpxuwh81DQBoQ9GakTwO+9i4OqrBp/MpOnVQHZbbLHIEJ/IE+ABzky
GMFVcZezAXrj7Hz7tKVF1pdQn2fA17Dlkwp8qaujfueui2T2upUiydq3uIBLKlsYx0TIqC7Sigee
F0ACMLyfsbyFV4LeTnqWvIEM3EB2RE0ENnx+wJcJEu9g8oNYXrTMQpUGnNAQTiaa3wNF2kQI76x7
6WznM1gQuABwJkXtutrRtIE9vtLJbdwTdVCyTIOI7KV/2EOEIGHOmHFNsloiPiXRSvwcnkL8QTbQ
pqCFlJq9l//lCNmDBmvZIEdm1yOxp8vs168G/AM1uosDZpwQ5elYxLiCuypNPu+ZZF2xK6n39kE0
TLE1Sfmc9U/+Hs8Xaii73B87HwvnaLnm6SsAwnjsa6xdvAFBX7YIDvtYxScQRtf3VtIib1+exsj+
XjZD3VypT3mUrQWzrOCTpKWZlevMJkV6qdMiufJISQxtcr9NnfZIpujXfB31rfZFv9Y/WLHS6OpP
NVcVzrntFfeXrV2NtQEzDtv+AOBpERYZUJ9ToL9+mXiI85+1/OlC8k1myfhKAUmT4TxRYEWNhs7y
FR/6GBzO1P+X2AhXjYvq7OMjlqJc18+MrxxoP7CCozTZzbv8FQsR2nRVJ0dBpIzx5rzyfLTPkt21
kfLwN+nmLHg022gtKFT49p7o0WTJN14K3OooN6Jox/RkeKDs/OycON5NOhxGAUh66NdZWCcI2+jV
yQEvH3w6eR1buU2/SccpglXWBSuqUcLRZ6XLRNUQKk/34xiLo/yoRdxWfEHwSbvUeHnOOzBoNIoP
8O7vq1QWyhUgYMtrP7jE90NKw6fZmct9CCRueqko6wooWnKrQp6R48xI2qKEMzLpNniWSIVZ/Xs5
x3JDYilXaGId9dFznc9rvLeMpRmvKAoWpNU0JPaqQVuUNHmQ8MqZ7cQnZ4ZymqqaTUvOjdI+CDYD
SQwfkHz+cepBaKe7vuZy1udfTnLGRwJfYVuD5o/NndiFT5Sj+e9oA6OY7SNpojPYmtjLhaxm/PCU
pmblPwtW5EzF0Owbg2jH4cKYeUWM2h5bZHah0tY+3QfzJQazlNcOTwwSWkEAp6jthu7LTeT8W5JC
/Ejqy7xubQdesfQG6S9m50XCfqjv0/qpmqurkwjuhvGBwppvkVTtqydAMidzt4xh4w0eLqEIQV0O
qCPr2r0BHISY0Vws4ovRbwnase/D1tl8wM2Y3nWgrmKeGSR/Jfv6K3H81ag3S1sRikP0WvQWgqDL
wN0Y+ZeFsiit04gOUm1ikaIREHkRZT/46gjIfD2PjqUBySLz8242Qv3xgKUOr23SHz1qnfwBml9X
JMKsVqlb2VCHSysSd6XZybXjKtftis0Qv/jKZxEy2mCTaB61k8KUHGo42QlDwS1eo5SXb3izg+J/
95Vjmxiweywkot2clmreXaJWdlj5J2lbdLNKY2ET+JX9Y0jXk/+4uUkilLFov8SHgzBOjqmMmsJ6
DL80Na38klM3Z3mEiM8k2vPUot4Sn9vCiXrqsPuqStl8zoEkbxho91S2o97A2H1Kyj+svOpXOj5y
yJUBguSPJkPkm7YG66kXnIOpu9egjhqwuH5HHCqvFfpfIKmQwYfhrXvRSUOoWqoz6AoQZgz9zJet
WjlWUjxjfvs9/1zVKiBKVUa1AVk0Mffeo4kYuR+OxtkdZ43HsnAfcI9olQnmH/JC6QPVdOdEwOjD
APCrdRShUdJYA4sGJ+wv/+MC6p1Xoy+vvUP8KEqL/6RT8B21BitJz29sIm5kRfuTbplMkOCA/Zf7
PY9Ad4fZweLeMd4J3P4HmOX0MTIdtp4wKoR7PdJ3GW444nDjSUNfKmzpDIgT/TMuGjsbzdSCayS5
beFcb8Ow+hq1qiPPYRwbHjtt7vIYEWsXdztLNNPdzpYyUlVHUoAX5X+4i9Bcmc1+MCjr4DmOHyqp
uBbESMvudbThx08JRNSwRwzkcgzf8+9NqE1tSOzox1UbsXNP/Cwp+vbrjHJNPRw2i8JrZjVwk1yK
/sSHr4rO12bAcjnswuwMWPBxLI6Ba+3fryrc0YvqG7Tu74vPItJJ8kmePtyQ7Lsa8GQ0jkQAWiUL
QU8SJWEfU0xWTR/MzXci1f+kMa0ZmkcwplDo71QsFLoJCKKKDreeL/9kR2PpbU8+e106mMo0uF8M
HTgUObyA2G3HoBnkZoUZ636J28stg5LCeZcy1+n5MlyatwRn/oDbKlCZ5rgJGoZzwy/TBLjqEjP8
V++w9/e6uzMMfWtiyUJQocsiWVJlWAUm4qJp/WIjPMydTpgLLtz2gbpFUc2NlkptVCtypwi+ZjCQ
YxzhBWCPjAg1/1V+e93f7yEmhft4G4NK7Y94fzWCBts3w1LmqfUI7I0acYK7SNa3Lh0SilSUHPUg
trkpVD8Zii+uZotaqyZDFuzkJG72XOKocDLuHFNb9v5jxyiOAVsdGrNlPa/szFkzK4gagnetFmKh
1bqKAqQB1EOfh9vCx6HAsW8Z/CRyPZUKQ+WkS26ahLO6MgJ5BPPYAIuba1dvDAzPauci0SgjX1Cq
9CuLKjHhPgTqwaX1Wz82V6iQOXahG2TZWGrE1yFodV2RfYPvf2XouUcqLS84JbEiMIi2MytGHO/G
YR78jNME9CSVSEEHLsgkhbOAuMDy4aS4nPizP6hROV5sz6mJS09ZzwlbfjESUIJP7Igd73iVkdj2
CzwX5CZGUvoiWG8VjbHt6gafJ+p10VdVEWr4+JNHuwa8sEOeC745tGeNg0b4amzLs0aTmJR2p2da
ngUZEk4i3S0tEw/AvOqsBOA10w+OfUQuX62/30q+3PBRJzkodfJdr3ZYLfkpb+JA38wiUU7RPi/+
IIabXNxzTToEJ0iyEEM8uxrcIHIN5IKXkNh5n8ESlymQ6W64Qbf5oyQitHDSVweWYR/L/hchCwdA
Ub92lz+NH74tFrlcxl7xUnm/4VGkuKE2dkGlO3R96nhnpJrdInQY76/oRHNyX0hlLZ8FwkLD18cf
EPYsK1lvqOdV3D0rE/8ZuJL9/IjXy4hyPo3w1ScT+9oIKSJMZGt1oLO41GspyeUNnB6kHwTc2tjh
j/EHujEnKIcEPC9LIKj5he/IyJb4JAcfBaHRVlNqwsyYlNjW+iAE48lJv6TKWQwR6vSKxc56xhpG
SCd0KUqkXMssWvn/W4SZzP8UiS9+osXxc9Nc4rTCoDPjqXpf18nYfFng0hM+uHWAdwYM2aqRzS28
gX8TAzFf7O1tOGYf3IdMGRtjJT3F/Jz1VFSr1RszjQ4+vJooY0R45DkthMY7MBFd65nMtlxQeMj4
cSyoCZmay6lzXWxHrAqA1PtNgVOvjrHhOhfq/wQCaoFbnp4SaOmvLOAx1R0Py7gqHli+WfF+Hvfa
AejvFryNdP+z/k+ShPWRZU6i2xSxGMBvU5ARzyjRTAm+uTE3RrfIrYOqXnxj2u2Ji9xpr8Z/NeoS
37N6rFnnZlpneBZBPsxNBk6p+R9NiR8PM9lTDg53rQvUJE/rIqL48u0TZqZuWw8o2JEHZzRyQ3wD
nNPgvYIlSTWxXcSuIdeW/0tZFNciP280Rf0gycO+PZVoDAtRiwxGFXC6otAV2VTHrs1qbABz7REA
G15SkYUis6i4zfYQh+YkPloXPjyYeRDLvr3A/KWQypPZMFTLr1wNJdCqa83YyRdHxai9Vakni4mX
dXPxRyRsTwG/rGiwHQjveYzVc/7n9PV6vEMgKc2Rg8pWniqToviL9BbOgK0ocKruCoMrqMXUKh4Q
yO1bGq7sPU1NK1vDYhPSzGGs8QFZiT22FCsRhHN/S/eww5dzzeHH8Nz9glR2fQMIaHuHM5HP5kN1
m/eUk6PV7gsJflT0ZJRhvzpVmKousN2L2IczhZLjhQ451ayTwrPztkcdTn9r1kU4bgTu+Mrq9DSL
twnkxAP3NPrTxN6LbES6UcmXgNlTmBEArbEALmvLbiiAI/1shd33JbgK/nksBxa1doLWadQ8Mo/4
QjwyAQbOvZKEMO3KVbVc8GT95vXZJxx7z3fb3qNgVHP8XmnxSEgCdLb3LGpCuP5va0t69t18KSuE
9eszsS67a++8ceMpXbfxh/rjrH7RXJFxOZlTbdn6ju/+uPSnia7FRmbHg/078AfzAPFmOMzei1dT
8t6KgR3fJaf792U8ZOotksPlLqtKBVun8f6gmxu7AGt+prAh430np+8kVyZpTCKvOYZpLt3/LDEu
LPMCbssx7ICRgTKM8Qn0bJZunfOHPl80CxyXaR62kZdvV/DqqUkc03imhzy6nqknPWFFsRJnfP01
9lyM8K+MLmOsQgLBJJYvmCb1jfJJM+S0hycVXOsOVJXbNCOsoqappPXXQBCDKeuxHTldTsUUvZzM
3v2kjSDApq1fK95qDOa19ZSAxQW+Y8gxIYwfK1Xn/lrQq5kGap8oZs70d5w3eh9QAYWCBEV9BYu3
IcWx4Wbo7/csNywVLKIidMqJlPv7+6b/mwJVHYIz4fxyqc2C2ubEsTRCjqdoVQ11IvSmjb4wZEVu
eN5DxRub+BybInZ9KZqI7Hkh9qZ4owtpk+K8TFiEriN3F9GYCUEL70XJzudT5e1v97GnXNDTbYWg
E8E8ICucK2aUlWeWt7WJDQnHAVdrHxTLFpVWkXLdHkPRkNK/qR9AX4CuX/iPKZo5jt+eZj87eaNr
+rrWRHy65HNEcwUEF9q7gCc2MVKiIlMEgrC5zaGxhC6kAZIc4zf1amoWqS/e6iH48ZMVqMdv63fK
R6hL4h5L3DwpOv0jKVsGYQwD8EF/HFxL8IQ414DcNe7/3UR6y+U/eEvijrRMh7mLpW5SktraL3bp
GAwo/1YtvtIR095sa0pNjkF3O7EHn+aeNsgFot/4ZBOlFspJ8bbZLAcRp1ga0uHh7SvoxikR9YN3
KweXt3Zto5t04LheHQRI4+6/C6x3aUcpoc42EJ6mGlNli72mjv/zUyPQvFHWeOqGoA1bHQZdRCl9
bD27I0XSMPnG7XZloCiRphfaEAki1TTHUXHcZEzA3AvIyE11aq6kQW/7sVyTYG5I8LDcURoAnDBo
XJPWxD/mEcipcHR7gwxvqK4Ehs9t8Xzdl6nsVtLOG8swvzRXmrrIZLHI6CBO3xnk2NfpdANliDMG
j5h7wqEzsOiVd/RC9XO1+ZvoJ14kAvYBVNvM/nyAMtjGCY0R7AtKU0LIOVF8MIK4vRrE3ydGVCqP
IdDBMlTEXjzpFMIH6fxoZ2ljUmzsHHbTxKlB3B0nGA9tSzE1xrvXOB3ng53ovTZh+zajkhYeaOc0
fHmebN3IA0lDkOCnr6Y/cjv+t0E1c/cxblPlD/W/SKLja8Q2xogKQodSCiAjwCwLoRiKwozoTZ0o
k2xl/XL/iwS604SbGxa9TY76wvWvx1pIeY9/Bg4HFRgZBptgwOwPScsIKix6/W/YGu6bz5Rv7BRA
dc79Ur8OW64iqLHNDguKfu3j9cghf3ksZ3jgY1krFRkIrDC0j71fK7oRn29KhNYjiy2uratQwXZp
ip85Q1VHIERA3T1dvKTUTA2i1UGyW4T0ayJ4wuWJnwDDNnKVSTr26NSDIhiBBmPycyBB+oMhq4A5
bxgz5Cda07Qy/EzwUhczPONhiP1ZctYYBcn+V3UagnFvoZxA/8jBafvEZHzvAzukHx/tO3k8wCEQ
oXylK9fOhUtJU2Cv8FE133Zozi2q7WDeIPz/KOb+NRpYb8amffyt80LnkQursQpQmpVrUyXirBr2
cvXN5Aj/lkrk10ERjwBDBYo9z7SWS75HcLZfh3r9THmbQ+wr/YhcknS7zj2SZNVOWHt8ER4NLNmb
ASFkrH4dDhD83WlmnwVI2eHm6BNWkD+pvreXluYoEWb946GyVO1h+aJl5JA3oFufr2LL936YWzWP
J3AxabLUZS3zGhojZoeRgX2sdRFj8frYSw/W4aWOP51oUOW6KvOsAAIgzqQMx7HqRYaWjdW8ffWF
4fo6p+Y/4RO4b07y8HvjwdZmjcTbYeJ4QA+CF3TRC/Z05C3/VFMY5qig0vsPSeLn/csyevih7Z6Z
TefcHy+gJTGCYTw4XLhkEzm2Mia89MAt3kBk7XjoqbE0GG/EjqwJRDSlP5bb88XLkEWHvVuCU16V
gUC9mbZPgVfwhRltoXMQ97vSNQPiZb9m7L6Em4l8LOmewDqHrePF73OXmu1RQyHj/HBQeIdMgSou
efwNDsZKdJSxT+3vLWMnSZ8s9c4bfejFZoDshB1WgSy03AwEgagmOb4Zfy9YLUnTs+3C7ygQ4D+M
4pgJkPhv1LUgNUT07yx+P9RBPfsWEnzxh788HKkE3jJv0Ywjj0GiG4m/NSKg42uowgFEs4l4/Wm9
foPCsSeyllt2Zi9N3tDBvA/tFV8MwI3kMSwl5KV9lVoWcLXia8Dp1bFM9h7Dohki4c1FEOVS/Hrr
cupn/PVJEH8mrs5sEkMY/ADjr3qUP6Sou9ZdWY3AaFGcRx2PdLnW0G5t72uZzhAK9CXMA3WLthnm
a2TxrJOsEs9bOlTm02vJ8Xag2WOH1qfR+l1z+1/Ddq39ey2BJ+9YMENO1f9DRtswTbC+R5yEepl5
OqJ762C56d6/qQCT8PD/lWDqNKmPrfrQPKGLCqEBK7gSdu2cQss/Y8ftpLBIjASA1aAa9/RaBYu9
ZcosCr4rSDnyjyxONg/Fm9y44LDXQC+wTeXJXjzvNUsBK08JD3hBVgFLbsONHM/7nhXc8s0XJmfJ
uN4YGEOtei4zNV+1WIAAKad0TP8XXWEGf0N+iIPjl+f8rkY887+My4nIRg3vixOtWV6D1e6QwYmJ
dmTJzZv7jKGnHCn+Sq913273DKqf3VWZR/eVEqLwEuDz7MD5LW9x1nEq6lIBMzAHU/ezLv/C+c5f
h+utvw+5csTtKi2kHCCFo5zINre2pQL5AgUICT8T31+UBSRGQwWWwgOEuMi+ReWz8IVy//i98Mhq
J2UCqkXgy4YVi8FiEGpHvKvyx4qScAKaPgwdJc8xPuP3wrI1cmJz0mDWCBuQ/RZcNNyy+Y+Z59pn
gxCFS3JFfHkYywKsYPO+djwhd9N7jJtZecjLfTN0P27phNWW5Zp/rNGZ8Gemd+TPWfjMP/aZ1vb0
suYcyvjumScOGCTu2YNqAmRb5pYyXQ+QWklWtJRyOjN/5fvnOYPxYyQf9dxgPKkzXjysPJEIazbc
IEwXAfJDn2AGVg7DlGmfECgMbp//ndKgFdxDlKvdKttU9Kg0U96AAGsQW/WqDPPpUl9MM1XwLCFb
us0UgJVn9D0/pAH9+AYCRT/ogO4+fM1XwsXkgnap8yTxjkLRuX2M/dsH1WLH7g1kLEVQpzm1NuW8
KxQ7lfou65YCrh8jFVDdqPGfOw4Bxe6/A2QGBf+POVHH62uBAdPzeLFbsZr/GqyOXYZQeBnnwj3G
6P9iRFqdHhQuTYMXZM4auXqKMgtxtiLRwMywKpBqsznZ7nAYIfDfJDGcMsC6iXKyd+2intAItLYp
ECLc6/OetJpQQJMD+Z17jcBvfKPVNrYW+pZl9DoM5vyVkQYVjJfK2OmmZl3Cd7NnZ44XlQjq8ISn
+0Tx3goKyN1YuCtB9RpdveoXYeuGk+f87TVDfm7bjjdvs/sWlZuHPsuJbxJYjW4iZwIrbUSjD2B3
+gES+EBOdlWMKKmsQlQJwsDkUUs5IMatJTy89YmhNhQLwu4/O3OHsvUFln42XZCa4Jr4kTk6lQRo
tlvf9VZoHN0+AK1uBPBkYFBjWeQTbY0dp8w1kL1WXWusuu45T9Ff58P6RnCFb2vXfk4kUsmPYIh7
3+t4F/RiWwie9fLFzndqZDsvyWGsLoAtI4Ddksb5xng1rvFWqq8ic+NgIwG+MlRZveh1YVvIFRF8
tL39FL5MbMyqk+b1B/tMnDBZjggaLHcrFaGRgvkG03XdceyAICplJvAcCSdiCkAWaN1FIY52+tH6
QHd2+ULCRrzdgGBbkTQEzhJHUZvvYztfgZPSGiZ3+ESjMgYfJ4FyEbktv/BKOfTQUc9HyYCQ/SzY
8KFe2r2EpT2EoE7HVyZnaoVShMQkc40zl150Ga02s2ICLNcAiQW2HPpYNJvJ5B7rGzFnSLPsnJsr
NnbUHza3zckctQRrHt3zpz9OKYpP7Xxs9kNIVRzMYecrJprMi6jbN43VVwJbRUJ4dCY1OzV9HCX/
I/GOJTjIxbZiC88gXjcVW+L321GprwK4M/v5lkKAIqq6J0g44mQtt21a+gYXCHgN3cGSDHeufsEX
wbM1hXdI7m3ltVHPFixn2CEVci3R8uEWBMxpJl0yMUlDfh99msLYfTtwigAABe4jtW0zmkwN5Mge
Y8dBjtvg1ClogLQ/LBAlqisUpdpZYN0KQ0aD02ErxnOZXMbEH7yuQCd4rI5Mu0+n6oQ7+aowidpW
bGRGqXYbGNrHcZs55kYJwFk1aW9j5tZiPkwvrwZunFoAmcZ5lEl8pu8swVoprjkU148/z90NOcJg
qXqbuyFUqVG7Y6qPf7v3Ow3sfYRv7N01ChYLrkbdy0gsQQAy2kU0B3NveAtEeWx7Vrd1BBJuArdO
8uLGYWmBJ39IuEqPtc8T18M5eErEvki7cHKFUbd2kbMsthgBpvM6Io4k7D9PjtevI3z1v7SApEdp
DP3coqbbj8O+QMWtzVDxBR9yYR3VqjqXnqy84AzhFIKDOqVkx9UYAqUfGgTc5yH1esNWGaXfCeZP
6gcr3WfIusO9fEXh09Qsw7kvI0mpiS9HkiIXPOoD0783NiXPDtwZTzSz6eVcUDU95ccyHQP/xIk8
hW2auQjPuHQt5SxBeqnHlYF0qeU7UyT7ofq2xgpHrCk2wbv3iKa3A8HIuDgeO4eZGd9a/fHN/VPT
HWk2LxIXHyKUDbjE65oE5Csd5p0/t99Ho4qLEVQ5/SW0wnaWYRwp0oFaGAtRIrxRqv6obd8b2n11
PNxmGbK3Vc5+RTwQH6WknKi3LiCfcrs75lKKfBaz1RqSBWOosX00cH1Ehpd3OLYphqSm7UrZygQd
w0El003rgAowQu4P0JFxbnUOTGm7GzjE2sQKSCe9J+o/71H0dLQo/bfFnt1pKEdZitLvGosyxxTK
/nRm6azByb7o9ZJAHdR/caNM8qeNlca8GR3jsnCD41NW8dafaWxYdYY25gwG3tGwTH1DaYv16ws6
Ip5Gl80SyP8ngAmLehGmFjFymb76sT1NzYwi+o7SrDQr6kIn087u81M1wJIfRKbyMwSzkAWqB4ka
A6aZBLV1rkU7Bx3QnstC3o4kQ4LfegHWO90PRta/bDQds4mAB7nK+Eu4fgeA2ymE2MIluMeD1YBW
Sh0G7tJDkpUi121EX1ud7oypuoaPPF61+yPIPqWj1O1z39SgijShIvEOc9BN46yMkPeZKS5cVyHD
0hg44deNFDRl35xlH9BozRn5bavrphj2kphjRXfqpO7DKCHdHaO3HylNmJkQOdhli6LR0CCGN8FR
DKfBS4kBrnEOszTwxVLCGCilBbY2VvoZ8Z+tgnzKaw8I90L6mFzBpwTA/tPWOO/DJXBCNcnpZ4JC
hv/RwsOwpjUnnrVcv2cN6RG/U4EocPuwcsoLiZo3dGHSivH9/6CaMm0WfzgFBnuOd7oYtqpH/h8N
YX04QOivMAHELfHKAaa2kAGs08rXT9PWrNMLJTBljFlB6D7mdlMMhnTQ5ikp+EPiM9WRy+OAefSA
WgeeYhj5k/8FLiHz5P5Xi7ZBZED0KJhkupqOSao8WAropJiHs0fm1IR4QtD8nNibtHyxXiadEhtx
xJKBwMSTQ1uUEb5Q570UsIVOQeKBoUETUh0QANwG9mu486ZuSIeQhjyZOpfB7QN8ocR+Cz2mlT0p
9c/fzpRfYal8e+g8uNJSpGTWf1WiUgpGeOaPZjkXtUJS8QEQMV6q0vk8igfNac6vQseBJrkxs1ft
GK3Fwd5e+PLjpIHqTHt3WVm/JoGdHTZvr3+4SScJLjTAfxPX59tOYV+4V9M3p5HNvdhVXCnGRoQC
7B1NKAAFID8BgR48IroF5KBS30AB2YsR4WiGy/f6i2HPyo/uHA8lkbNWQ/Id4WO4PMhXCZOccgTQ
2ITCaNNbdZ5cso+QnZP5in3NMtAvsJX6MWendXPrPO3qCLYQzfGs1nLwO2ezTu+CMJIGxbUkoO9V
cRwnw6vho5b90f/Ps/yNv1xDyERn8Sd5luH//e80sqGgkwZjnMis3hFUp+nUwLIJJmllNQPKwpph
9hIiYZX+SeEjDWXjcR8t097mMnypdJAjEtil3Kvqk2P/VtzTQjj/A9Y09+Pd1Coenzef7A2tJitN
kKA/MPb/MEsge+Rw183SuciMyP5acC2iGlx8wK0T8npvuHgfBc/1Rt9f+Y2jJGNsDqEefAXpCHn1
46BJ4/3cUx6+CoF/cbQn6KzPA8TYXEDuTNUJ5Szeueppo78PhwQ09iFcj5Rascv2ZsqI2unubjJN
QFrYmzBkB1p9yRC2Uf1gvVxz68yVSEHZBAKOtqi79WqCI4puPiWz3iiYSZE+JENzx2u29KnrLzqf
KP1N3M/H/iSjky5C/UXAxQMSS3U/nsAS99XzVGf9vRHs1V5SQF8AAK0M+vYt4zShjtTJijNQCGwD
H2S/Z2iKZyQuf1EWZS8dacbTs9apMVP9Ub+XCUzoThQ44isTmjD5xiV2GjEuGU+NAxcCRcPLoL4L
oVgK4O3auxiDiiuVjZrOQT7V/sIVF9+/8uELp2JPPLpm+lxrM1sd5MEro0JpXLdpUbh4ij8bYRVq
/QXPCahlrneAw474cgC+aECHR3SiMdoP5LujCTNH4aqpNJNSQ7b4YqbzZsmguQLQkVrMqBfDB1Rv
MICMphvClek0fVGpzsNfH1sYRuP1wkxLHk3A9lCOI8IJPTRbp/Wdy8uLhFaPjKzyLtSGCQnHgJXX
Zqj77fVt4zU8YgeD8lfJoZCC1CQO7b1JeGi4kmEe7tdvbURNWK/xL0eaUL7X9yZZoT8OGZRMk7z5
MVGAcDrm91HkiW9setE7z3Bzd4No7YMhERls1BVBzq3SXdMhUM9NrGPSs9B2YKlNDCb3uEAAoyhF
36Um59BhaylcutjW76iVFLvx1JIQ0WS7bbblFCaSawNF5Qzb1ntl5jryibNi16Zoie8KRN7XGZe5
bLS6PZQaIKRixYs3TmYR+KwCAOhzuMkJLi/F2NSZrQbzlUT3j3IxCSR4e0jajdStGgnqD6E4bliv
wort5USeAGbsKQXslqEs9iK8rR+9eD43hEC6xWc0yNVzFilKiLaj46aHQDGN9EqF2/acCbPmWphN
HcbZRly0ZyBTJURDsP3MvhU67YAUmfR+pgRKZrJLm2PnijcpVonJZrxQTA1dWZxMfMruO7mzj7Mo
SJ/SSuAV4P4lau+Q4isuL60iRbczlez2nxcxTX1LFwKve4rJO/hbrQzt9iZ+ZoYadwvVr+S77Oln
JKOZIFMQfsdPMt3fvCIFpSdZ+Y7gtjlfHlPiVkBpUoDOPqgb8an86cDuZiS15Bv8wGSXBVMQpM6h
Sr9qWLonN4/oxHAJx4SUcpQBUQPF29kA0KQLn2q7odn06+0ly0UgTvnvu7hY2bLr4EbUfZ1f4PsC
wY07schk/XVQfa1Ct1qK9dLGOviORbTrYwMt2EWK8DfGJEVpizrsCNOP40HZ6oMxNFBd4T95Dh9y
/VTcN8TW7bH0v2W971AR7U3sEqNc3lGyHEnCKW7N0cfSMtIydZK9L4zQQsnLSTlf+SnBASE4K0va
1geoa3dJWCr9Wji2/WE77jgo/ilVRWlZhdetXH/9CyvmouobalXHwELtjNvz4atVm2rfi6HGr0q/
9NS29MEhMtmVeMXQfSQzaogTVlGXkD5xzFkkDxrANI8kzc9ovWryhrt4zAu3wV5xCtxEqcYr9H8+
TbvgZlSgfNzbDLihwvVjNmCoYEXPZ6IXxvzgG9W1UFZ05IEuFi/GYCwKB5K22S9my1kXN4fgLNzL
y1T3s8XtSS52diFU13XfUekjKSd7I1xkdedvN1y0sgZcrVV3iw/AxmSaFC6qFxFegA71cvdfpuJQ
0q2+NN9rgtKGLShLTEov2FPGQBB+qShQOjllYX3u0Ba6Y+i7RkP5pChk8PIPtkXUi/pOrosWe/bO
MexMUUIo46pElkY34nsnPz4QuKvVGEumjQ8lUtS1dEhsmjvEEuPG0fd+zWy4ULgm17/JV4pcb6sP
yet3UYoCXi/Hif2K6VPNfKUYJ+7RFr+5+M1tYfTJqcvmeSbbo7MUSZJDAgW0qLEeOHQkbrb+gzAW
eRXyIlEA1nGwWocsNqlxd72SnyvaNEKtpxZsRx+S7DciqFrpG1rttsIyy0zGySohyxKr+psikyoh
DTTF/95fdjQfou9BLwqsZlLFP20hS4AszcxNp4s34pZVuPMMKA013xkXckwMw47HccgadLEqw2Hb
70ea1wSnOQr28REhShWqct3Ga9RUUfO6Vcdd7jqrcA6TXRsrI5kLfk8l/ZUETsNu6sCjG+axJCnN
8hEAsWUSiu1y9O9rVnhNc2s/oSMmjwP4X1UhcfS87AmHPC+IzWj1l8CvWyOqgR3c/5YPzy2bt0QL
U5LLVBJ4mpoNKCPhM9nDE+pisHIQw8bmbxSCp0vjH1CmsuYuEH9wP/CdaK331Scomsvae5KQFktE
7YtLc3bngKSkzh/nM1/p30OMMuuwI7OP5LV6oN/yPduXXqejetuLTPGtHIgToaSCJJwUIALQ+I9w
oa4gYfqzF8dvqUA7mINrtalE7Anx3pjm4RIKPo5JMtUssXqp8L3bg0KuN1TsWj9eLQMhphwECKiS
oSVN9iMPOrsmLxJ8ZX86vawsP3DQwN/4Xo0Yrw6PZ12FyX3Uct6+hapy93k3ME5X38GE4lpp/QFt
blJF/vuGaXQd2cJXTwxCBj/EuOKpY92Diu/0l5xe12xHyyG+JzYaJQxlUx/HhrAI1TwqOPAb/FxC
E17YYUu34oAwrLD3wmdBm0tffxTTPwiJ5u9gF+5Rbt+2J9JZO+hGUR+PsPSHsgwhAR5lP61cE9LN
GWsMDP6jXys3+SLdspAld64vJj/lUBaRYRltGeIu5m+L62abLI3JQa120iDuF76JdX6PL6dJGk1m
/9B+sXwNphcNAB2MxCf1Gr4UtehmAOi3492OVJKzRbVXGhvNGXdmFnhqyia9N1b3xrQiWVlZNSs7
AlDkJ9C9ASAmp7zHcSdFmFUy6Jx41gJM1xspmWR+FYQNwGh6jZGqAiz6E9wREEtEZ+x/NX5iq/di
V3Dn1zUu1FFzwF+u8NxEs+noGaF9vmzaeB1XHpO0QlNqnZhJX4UAWuFOprUMrzEwLXe9C3VrSfQA
bToHEoy27ynBbpF+JI2yemQ53bEimIA+mu79w6wF4ZnkbS+yOQR38pO1AI05i5T1kUj1wEXHn2lG
TdqgVoKQqSVNTQPzMG8DOeDitgliaL08Rqk4Hg3sbsRMkTN0vTvol5qtxYY9AXox5qfEgX+nwtaa
dHcXdWQzIME2oHRoiat892Cq29GbGK4sMvfXpqRKf3m5ky4wMZSGV9VYctUJBQZHBQ6By+XnZAgM
C1p2Jlh9aXr8xs8lzVLubGYlgWBPHF5UmMq4/WO4GTYi8R9Pu1aF3yflL3aCHeu5Jd6B0ldoiImb
6e/94RiOFUu3IlndXbEbq/TyC9fiPw13Fsc3VACzaX0lFqQCgd3Nsnek8Sgd8s3MkH+eFzSf6KDq
GY//zeGwMAcocRfDTDscpjoB3HBnyE7ADyGwCE78ksttzS20y5oueotsz+JtG3mVN2ooisysl/5y
g9Su4+dWQkMMGifs2T1hrptaYN/xAm5z3e8fKUoxasK2OGayphdhSJlNVscDP/wXIx/j6MgedXdu
eEUGkFmmE0VJnYAglS/Y9Fea+uxJbyWRiPkorSst2yO3Pq201i4B12lgPeuizi4Z3myOIiabZrfA
mRvAmyT8lvEeDVjQ3x+Be9SYNcd56IzPB75OZWQJ+ACcrS2BIXr3MCcxXAQ2VBW1QbCsufN6tmKl
N2gdvOeTCX+ve66MEU6QHzL+Dxb2OlAn1vadLs3gkgE0uGYU3TAHnAenK088ehS0mhoQwlfhS8FS
DcXB6Ntioucp/CZNQDmyWJEIbvoyi7XEUe3yD+5VABR0qNROnkP0BZeTG8R60QxLQdli4R/DCZPs
JpQ7Kzw8fvLDOWAY5ft93IRxwIAyS6N7VV0+bEaKkQw+6imS9JDn4zLJ+Y3Jn1517z8WDrHTMK2q
6n+/A3qAUPHXv2Ukr3uKHj33FLc+BYI3j/oF6ZOrwh6Ywx6E8jh9nbytBPTW19zlmq249iDhMmC5
v6VicZCujxz/jV/0xbl0ez8+miZize42YBgMWnXNhbeviEueQb85QbmfetRYsojudm4nv2iICD/6
NBID5RQe+3JQpVbHUIpO6BphQllVbTMC5V5/817/SpY+TsHdBwPnbTKrfP7oCFoP92nq807e+sbV
pKzUFfYvWL/NKyeKEWpxhpeeMCq/N9COpdEvQaku8Qg+ZKBdVTCQqVBxoppOeRVZcTLHH9aWuqww
hB3SjPWTpyXeh6rmY20tsDIvRxXjggqKk5Ela/OIyN+LRjUk8ZMEXycFZR39/H6a+kspjTJfGjNA
PdIdw5mcBw7WebTUZHcj2zxXd8XwFshzxErYRsYn7UwbFV0HM3W/eSeXd7dPajG0KsftqsUwtfmE
0Zdvcrbob15yYEInPsdME+EHDO41JObxUfVx2isgBMWJUPwvBOqzb8qEE1x2bY9d7HUJTgUQO6iY
uHoDmmLBfpNddC5Zx7EAC9cww7CaEs2m3f7I+jrp1KVzsbH0F+0UxK8koNCh4afHUe7g1jUdT/jR
bWBQwgbnia2mVdWZa3T6oL8IK52OVRUUZufLGVgZa0RwptWaryz9Azcuw2SwSKMApvtmC8u5yqO/
YJk7N7n0yqUKsWgu8ozTIql8H2diPjNCkIdkC5jhupkCUrQBqPSGCh0SO9UZLnsSwgN997xRLXMi
tkRx26xHn3TCC/7c+hh2mYrkwrej9sQxs6rMi6ywyZ5myl38Nsv7evFpMfJk9lt/UfUl7nie3vDH
HkSBvajlVehk+Ts0g4ayNmwlSB2DXPRjpfIeUZjg6jQFGAewLIJ53dAJU3vBgFdNXoNWZCc9m2qk
R8IKVWW3Xy5ehF7J0coawYsmuS7KxdJigsmWKSB+RwwqnHRcNjSbbF3mBIQoZCrnUpuuH3zKEenD
k+u/MvDCAoqqKY3XNqJUhImKws+BVIEkOKVoYVfo9D1lgBpPyRTGcsxaUVT36QSNrBBJWnw8Eyjx
iUk6ugWwz1a6BL/29penGXK2HBJ6izolra61BcN2y7lu6/r6c/yjW2XjbPfg6X6C+34Zx8VLuhlW
B0up5GNs2HaNqk5DemxDkMlpQyCh6IrZ4VfSDvLFEGaG80LycUa75iWNqnkFf24t4jIbqgj7DAVI
IEnaZ0pQV6gUfDdJOvZPxMup8YEeVUe7vliUSI3mMzHZusZGD1I5t3BiJppx5sJ9xTq9xO9t8MsS
yNZlRE/ePvxuiDxg5ncBzfAhNKKcgAaDBUYjVxOwIxQ9maAVKEdLQYnrF83Br76plVONuI+r08am
lX4AEiYkgrAx9sBxmjEJVvw6/JiIgV69T59T14OXW0YZ6z5SExms9SKXTj8DIaID2Qxn7V/0/ZMD
qzhDJT6LRUVMksFvspoAsrsWQftgHbL3y3DpkE/HeZMWl5/RtXUUJfaEyVlsOIhFANecWlszjt+r
772G1T57jY3qxqQuj1CYcUA1pq1t3u6jKgGeTSmklYX/A8peFQVXnXkxuMahUMXy1X9C2YLW99qt
R9STyg1HFTlTq1VRWNycDLmp00VHxO8f8uGxhnym278saqqfCXzFcGYgfGWVm8ZeeqTHz7y3/A1k
PJ41vW0YOj3/3MD4s3yBbsESAYvzikSwcddM5VuvX4VyzjrUsezOTV+TJQZavoYyxF5X8GYm4jCd
3gGItPgV4UBnaycvY1XO/t5LRTEug/bUT8iSRczVzDOBUY9pLh8DFepqPq2wtc+ONT7Rc+GFwF40
sIW276TvZIE9tqWOYKCq7bUN1Fe9GfoKabs4h/VOwR7xPOQm5EnOTU8zJjt9717h67P3Pk4qdOtq
URh/aAoWVcWKVbYh7WgnDvzTTfu8GNCPJvhqDUQRhO9PH5KrRdTG8AwdVZLTAd4SpkqFTPn7461R
I+ZOOSQyXvSObxmyMJjsDENprL1QNfAuTh9l0Z8pOeMtPJ6v6ubPVpiUu0l7XzheDNWdwn9wo0zF
cJDzFI0x0/XfIFCM4NE2cQQxou+3NAVLx5GpJZZqGMaqU0gcUffR7BaG6DceMI0H2sredOrSyyp9
JEwf8g9MBjQ48/rCKnim3Cbcxg8DawgvANMjNOylORGZ16MvBU2QYrCRCp0/frl89odYPplMtSCc
iIvLvbEBG963PiCqCntoB7WdTdfJYslsCBZib6rcQoiezjb4yRffWOCepNGRo27GtgZGzWftYOde
sYUKBJfqC04j134kJKcBQmszIOim8Kq2l98JzJWSwQf82vUrNSgbpvJO+FNDnyfjZgP/SSlJ2T+D
kpLjFGtrod2TXzED8M/Lu92LcZsN4wMRjZXBdNdDWCm3gSH/+KwGLA39baR6rFCDOgmCTYq4xc/E
qG2KG0yyVgGzVDSWdBqRenKq3sOxQSoxAaoGg6h/Ggegk6QISIoSlAhs8N96cXaCxJ6poSX0ba8E
ytIUO7FcMMU3xcYbyEsV355yhSqNHQ+PZKQaIK5oSO9TERJB9NpC1d2Gk0xC0Ftd+qvDnSntEmH8
XNHbSzMwBBun+MldZ7TcASb3Be83hwX9NtGaUCNJCHb3zgiTF2Mkg7ExWpFPhywQ+2cOAJUuvy9F
NR3UD8s39HQKMSLewDc5ijLzXN/fVtVzTz6Orscxl4LUopXgUhLegbPGI0aNOhGVi/u71OL32l1r
prbqoZc0M1tsqeL8pbc1VT2j10hz1K3r0wjQLAzK0bpnbUsCPwCKCs+3bj4e/w6W+RuSxrcUSnAQ
r22QzltdIxhvJQJPnt5OxQte7TjDhOYOGHwwxpGxvT1bFMzoFT4G0GqfpowF/5qEvCzwpy98x3fR
5HcTB64YW/RyHcJ9je1PzHLzZ7X81m/Y9bEBCOC23U4LG+trbCzWX+bxtNxFkukx865HyFYg5Gny
XhM1RSeUhUVUsGOSwEZzYTihVgOniJBJD0SAk6+i35Gc3PN5KvkX+EwtwT9ym1N2+G4HqgbBtnv2
zLF1C3Zqsnq5wLvLRkTnVTNQRpSD/b5ydP2+C855LUkne4vv1I6mGVgX2KZ8ipnjTAgBOjhpnNxg
p2OWP2okJV7omlOEzVG8FQ1aE0fq8PbfogGt63O4bOqcItM8DOk2pZ6CXm5CHm1S/5ohiRc1tZDw
H2EYL3LfZ52lyVr2D5sxxuTXBx8khSzc8mRBPkwyFmX9TO0n+ibNBu6medJg/tWBWxmZHn6Fc3CQ
naOQAuUz45S1b4cOicBHhLLR5xEKvTlPQuonuIO1u/L6FqSghtnlYdL4iI2MKxlHk45PtIM169ud
/vLIfi54kx9vQVHfToxXqjGRLsGzCPGLMHazQDFOtnrD7kHtAGgyZBGINGfBDF8fJDY3NKMzd9No
vELxPvQae8PZZyPEqSBSSCvJyOmuE702NX/igzX+MUoBHxOCKB3i/2wMu/opgBjY8AL/68dPLEW2
vNlDSqZVjMLMp9DH+eRV+fT5swDW/Ovzurn4bp3AoqoufylP12Mld4Q5mX9Yg692el7/BsEjxkzS
aQ0fcHnNo5Fr3R4LxzF2DifFtdra1vlDy6e9yaJIlISKl2Ddlf3J2C6dI6UGIUFpTDbJAE/Hmt4+
eHm7ZjUwVGRFYdD4lYDx/ezkEAbTOdXibvchUuLeaduL0qe5GRIWix+y/aeUCSPuiVeFduWGyYlw
tsaJpqM87yaEG59QH4W9sQA17AkWZ+yG8DHeejKin3m+z46LlOqw9Y/0eGHHoxn6i51rl8dvnvr6
gjsoPLModqoH9y/2H88U2kijZiuhQvItTevKuROAhuwoSinlsbQ82XYP0Pv7U7oeyKx2kZz358dl
2DHRQSywuiAmtXI7nsnJnPQkyBlUaXU/ARucFRIRCriF258I+Ex8GwlXnhjF0YYd5cWBDtqHMI+L
/SBUKMYVHeUsZ57/+KeXIghNEgFQoXTq/lllj1Y93eJh7hhB3dANstXgn9+hpHrKNguqGJGe6ZC3
awaefwcKKBRRuphvdSfLcZExio+7DObZbV+1wBGoGwhwHXbJWkkOQjq5mF2EquvmsCTd2a4vmbZT
2tsnPbReavBs3NCcoKVMEWPoeRmMVaEbxoJG+5YV9NrN1PY8c0/GVVJGQ6sR+m2rHG3VcBfYAvBU
ZVJslkEAzIpUAkcAZ1i6RGhp5Hi5FABvvZsZXyY5F1n9hs/dLJD/94AXZAmkMqyLHEBm0WhGERRL
mkbhHzCOy5QclBYs1gCUU461O9g0Cxm0qWNfsfZwWBHRZalI48iOLTVPm0AMDVgE235RXP1kmIWt
qT9hNVkVN3S5w4QRETL3tpmJb2n12QgjUuQ/+NVqTH/1C6WgNq3JW0zq1w+qLrdqiU5UJWUJV94t
5FZUVWSLXTaSmbxO3HjsRXMPfbL0jPl6LaGUkjS6F5X0gPMzKH1UBlqjXiwxOk7wK3JeTK/wkXai
TTQrNXtq4DAXgrpnPAfALUdDAewFE88r96MGNxDKPvIyeVPHr4yR2qK9AW8LuBjPyEIGtbOKkWZH
1Brw0tWwrlhIg+46re49WgqRBiYRQ2bCxRZzLxVxh3sj7cN3d/+6CrtMct2IOmvYKTJdRg1w+M4a
p6S4D9ORlTtltU0Xq2zFTZ8g2+iqYS2bMKkGV0GYVsats8ZQ8v2uzw8bNk6LRfRmqgQObLKxR0XG
FFnEj2ZDVPb3y4VSpc6YR2VFm7EOIeiMh1sPRAcFxT10gp0E2P/SOBvfAcsmMzTHBMOfru18ZJPK
lLXdEDqMG6Px4RoFb7blHQdi1MlRfc6TWUFgt9oUsBKIlueWP/bb6WvAzK8aSpiYKpK38dR/gbfn
iiY/jZ0VsV8kL2wg6IPMIuwrKBa3+57XmKaHkhHZ1l2+2PRhMZwS9JIgRpiyWR4nfPXCOg4uJifl
4lIcoawEK679RpQhf3KRKA11XzUo5DUiD8+papxsW7Nf/rccP43uiOqT5iEJjPljmwLvVlWJXn5i
ebWRFv64ISj9/AKJvknA1LpT0bpNS5OPNyjhDt1WlCkMrhDbEQpjzjvaVsmgM0JQScc1JFEdbetF
e07ZEzE9v7j1QH9pqnB+1ye1P+4fSvpadQXoiAUOLColcYyINVRA8j/XyJcEJJoM/P538ZbW7vdo
xW3vBmd3cwtEcIieIA3LQnNp+x3b5EBpcRg4TahE0BqdFz7euyGJPzIRHAEqbpONHWCONilwMK8V
3YXj72wRbMhx0aRTX96Z3SD15Te5BHQLmOieAiQFiP3k9OcZMULckBwMOKrxmSfGSPFvuWTjw71i
mNrtoqSormj93PnfR5FVIsEsysfe9OfNejQ2v7t2x9nGBjIh89zgUVy9/GXV7cK98vhPMpqJQv0y
yAdrGkkbjz3LYl36e09YPJMsSo+NfL1V1blztTmM7axR/NJSSsX7cwYduqG+P4DRMjybCRMq/l9/
rQ6e2y7LYLHxCgK6LxjCZCjn5vXmBa3pCTqhe85sUpDf7CfkQWu1F7dw3BWddc2LSgH0wQWB6TWk
ygyITuGErQiqyQitqeFjz2xq+AJzK9ZqJBFP3Vs4nLqSkOfl7j7NuLZ14hTrJmRYPE032WP8Dlj5
V5sp94PGBbRWCZ+13J3IPQ3HQC3PyvyODREc1Ox6lpjOPIyXBEZG37Uss6MkL0e+7nLHmcbMpPLC
JeHDNFTEb1s2VuGskd9v9kFmF03MgUWZCSVdMjYqoHnvKf1CGfNJMKdmaYitrH9YQVJLwYXLqnAx
F1FJ2lSAetnZbXicW/0YdE/oOCJ7Ytwztq6oqTN9vl/AgvenWVdFCaB6phoHyxO8AKX9uyOwP0Ir
4dsKhWaUTawO5agvF9OlTG/f+4a//XptaGJePX7Q0fAZC0KOrK9vYRmF9p4agDJ7qjRXPJmo/wUE
/HlwyBYTb81GozrpLE9O/r4J7AyH35NnGVeZZJDrWMfvkOPE5DGt0dtE34BZ8j2pouj5sixj7JOh
pdhlOKwHOk0njnkKbRzunD+KBbiyZ0ij6dPWFpws6OTuPEMY2cmP349LcjrlGNaZLMv9y3BMOSOJ
VmRddF/KY8PWuZd+TMcVaUlI6bO+9f8BmVqKi+H8/sQyXKfIwwxubfHDSDmkip4qqbFAXsT1Bve6
XOURvPD+AZjppM7XL9XUwOoTgl97buLOdQTBtk/1DhoQZE1sPgK+p0h9MhB7XEZtOkB5p+LjCAqH
l10VByoa5+xW+m3gONj/6jta0W9kvYvbsTbvyerAvpTYr5c+I+cwyMCbm8HbaG/IcQhunJb+Ofu8
spo9kqEEAJPQt5Jy6R4fkdw0EAvYRBcGbx6Ts84YpV3M+kp+jzaPrDyrzaH4znYhYubjyUvhJo/N
GVSFGGumsby+s9VEKQnNWyXprHW1zmSz3Kj10bFu4R68bHKYfq8isF9yrfqO0d9IRtOoILMz6wdk
SWYVvBkIrBCprPNZVU5xiTtYbUx07FBwD0ZnoDi2CGKEfCP/EEnB4DfTPHf0DKXaN/FHqWFcBCZU
fLkIVJ/EcBKkTeEhDFqC7Zf0FI8VpamI0o0PazyOmZlIgnSe6K3T4rXCz3gfFoChZ9pLx0f7jGDE
I8w+iYJzrMgzzrYskrrhi0oXSxh+qY3IThgld69WtwuqPnyYM6bY4y+zQWC2VbFXtjTcxKnJF5Jw
GuCWnPQ+Tb6p/r44XV5Xz7SO6XNqS6vIiGReCL6GpF9iAOPQwA0ZpnPfwBr6bMXELiyTXUtLh0yt
K7NKQUxM/fnaFmuugkEJx1//EsVWcYFo0XZQ7iFHr+i+ISTfe+wrfK3F30zWhZE9o4ssGfjyBnhO
CxVIoLIedNGhMl64zl1oLjbkhbYF/YPSrYPtVrmN4jQa8LRTZfBfL/Huo7MCW6RDoTUusajnJdW5
MD49P02jLecx0nQPm0EF6i5A50/MRc0vYBKiYn2AgNj2co0lBBn57EGWMqhrGXLIenPRB6gtiZmN
Vrw1cz9NxfS5yhEv6+3rIsrK0M4rIj+Oh0v/oZPcaA5m1ifAEfmJ8hEcu+yTB+eBG8OW8kb2gP9G
nEd9qX6CnKIqJOLxO9W0zhJL4z+Z7xfQN2WL6t5yHd3u7uda2AyVpWiempcwUVAyZ6NG7Qp9V6NK
l6sccOc9YlIPX0I2VRBHlJE8CJXh4Yi4EqreVkzsMBRR1YZALAZe/fnCp8TiKg1yuVVfqIcZGvh1
F4ZGqZA4gvsIHPckV3aYYYuLRSjR9ST7KM+k8+YdwSQKrAiBftrZeExFjalp5Mno5rd1UDYflNJi
fqPtzdHAA1mfr3CyxCVdVhYuj3n/dXIbVXDNo3e0MCOB6Va9cf4p4lGEoxISKoXWjbkNWixezqzM
nkpncxTmwG8q1sAKb0mggZSbzLt7dD0LZVvTxTDVI20wXnCk6NRHCyhh2YDov4GWohHlkj/sSrHe
36/+c4SJVwXSmymwlgUhY6HnZmohFmihhcS9HqvA5NslhpqKZcKZp4YSiAYL3qrADcPJnKJt6wTE
Zf6nocbuFgicaPUgNJY0QJBHnjT8jYUbvSE5dgZlSXrYxS9T3Ai4W/i+IcL4xMaXo8GzbPKNUVQ+
0Xd9AxyXbz3ZfqP7jWbWd05yeKPJ1AEkFD6fSyG2CWVRf6/EN+DFYOBPAMkKx7XPfheq3plw+C/0
/HzEsGs6PfrvufkHjHXBs+j4RBYVrXDr6fGy2aAZ0GYhCbUlwyIPqw+0wfDtsPOHhY6Z0C9tb64L
q17UGtsF7S3gXkX5W0SgizltNEvN5xqIxEaRpbJhax7Fhnssn4cDdxy4BXytWeWa/yim6pdFXEF6
Dojww6saD92vHyYQZdPsZdfOSBwMHfRTbW2/fnvASyYwg82tT8AKMqlf2DaAKtNCI9kJNiNAc3jm
exgxBn0KclQoqBQyWJ3strOHl/OhNzAfhy9AQD1ivDOsPwZ4Uob3AByNxJHcyVNo4K5AP+vqBwdJ
j4Ac5LT567MlrIXljTcQWB1KFRU9HW6YvzDndUp6gg1MGmyv7rQmcEQvOwKWNyuGlKAu43lDBNXN
JlQKDtC1W9cnm2BP6pWGN2fTtCK8gyl89mXIUBtiy40yDm8CG5Q4BM5/y8E9Y0a/dSBc9mp0HIOl
GRDaMREfwIxKRBXwZlTVQSiIChaOcVGeRDaGK13wMu6KqKhVeyOMe7hH5/1Z/7LrKdl60ZkH0idZ
gkxF8E3O8X6wr0chArrJJyF39S54eiiRI2lb3CAjuh5LKIxCwaxEldAxuuR4Rqog0o6TaBwv41Uy
oCOf1G+PA7HxA6KOoX8KrMvFWP5Et/7tWnN1tXu2v2G9P6KcMSl/ZnVL5Ni2517GKMVuT6yk1gZn
H59gdZ0RJlieBQNKVTnyjSzqTNrd/3ZDyk8L0MsUnzzQCMNo67A8+vUbvrKE9fySiF12pxCZwsgE
u7ty1BVyLYQJfAx2EhBWqeEc8cd4JsSRVRbz01HZTGmuqp4dXXy6eDeDIRYZJvOCrg2Bewgpr8kN
1KDLdyHdCZDqRVSiFTtPgujVXySnaVt5/W4cpVMjoposswzBViRl2tvb61hM4p/HIMhJiG94CDOM
gphJW/z41zVyXGG299jRs1Ix2vpdTflhbfWDc38QsHsDEQn+bgVdqb9WdyU5Sv2lQjRqvUkb2ThV
3A4JHhB/wv+Dj66ye8RgtDNIkoG5DGYYvjqSVs8td9fQpZzcsLZeeaY6PX1oDvBeFtpOHMXIXgfR
8L3JyefVJVkyhO85SUsGVwcgggpvoEt0rHH/iLHct7tvZlXFLq6E/i63PvkpzcvxJwSdO13QWwtH
Y4/0VSeeT08N8HUgRc40tneDxma9Q5lbHrQMD6591Q31ZE3CEEuoEZiwIGEsuP7sD2g6XL1LQZXI
FK67oVhDU+KdX7Dr/4Jx0vOTloM+CyVZy3BuUeRgDeqMw1V52qEAZsf4OVa4JsOqIawLsby+78Zk
9YqKwq0JZktIDGOvNktyOvMA80atuL40reiVNy0FzutAb7VGcSYjEeoJe66N7g/JkUqHll9zkneg
GrUPg8tQuEritw3fducZfWc/SMxPBzmgG6Gb6Phjpa/ZlaIiHOgQLIsUm4NvYdOWyM0/nMBJtWbM
2WNQdJRoGESN7jxn6ws2OIhvLfN8wd3qOm9K5aDLuAVCXT6DikzgtmbJhwFxwBtsT7z4DMH21iT4
0L0YKwGjIonYpgosRrW0FXfKz2AvckbRXAKAk+YS/UmWu4pmPqMXCVAGq65x2I3ndpS7PN8Ch6dT
8SpK2G8ouaIkLSBH2yWj0eYO0kK6BBniSxXqIkX7vpyQ3CUzvXn9Qjvmlk310rky28VI5L73qwoU
8h/jIRimwiF6zUPxi7SGg0LRkCpE1xSVgQoZ33xQ0MGnV0KmMkH8kRZ5mKJ/cFDoB1rOnB3ahhXb
dIIXkqzHH/IPWS1Sp2sMrDsiRM05iwqfRHUNecmosPdyX5AfQkZ0K6AcqZuSPfEzYES+QPHXmRRw
hKKor/hEnnH1BhOvuqv99bYnc4kPk1g0AO8gp1YjHJTryeJn+PsqBDoN0jUmyapTV+8c1cVdbQcO
GoIIb41eSWb+FpxAPdMAAQqbbcF+sV3pAjKdu0GfqWj73SOB3ek5uTFoZjZUri0kTDkJlkX6YtMp
BiXFBgvSY2Wbem5WLsiYObFcZtvXgDcd0qa5kgsDInRPdzK3uc7KYamy6g+KttvBL1fbNthRdjaS
SE2F++kPqDaXoUU5wum0BHtgZqSUT0gNkU27V3vj7KOinZ/JYh0Yikgeh0b2jDSjnVyhrBcXlmSO
NxVSBO5vo1898rePeMUELI05ubhc2Ypg+Hf49mNAYtS+Zu3ZYgcngLEIdSifWjZug4agu8IokO0J
Rvh8kj1OupnbwejOj5GZOAmKK1z1DBx3o5+euOOeiVUDtL2iqnzAXKy2NBohHat5pyJpUsjfLtCz
C5Kv3enZ/K1xhe0oqlXE+AoP2yLF3Tz1eQfMNRaEiTK5NJM8cp1cqqhXcmpcONJJL9aRRFh2LT1q
CWkpIgbQ4jiyAP4kmbpu1qqjAPeF1YSfKFLswK0ul8uk7U8xRDJ9AIt86tK7ciUpxO14tqRKZWwx
6MLIlbeqiGpw+x9vcnVYnGEIdqoF21qt9ibqPy7F4rYywykBG+ibpxwKLpFS1Nhd2U+7yT7AK4r8
z770UpIXzxqqQrsiT8Ub+bg34CWXC2mA5b0OWbrDa2tCs800WDy+t+EXQgsZgZdaCPblA/HG6Mka
Lm6rWzmqcLCli+q8A3oFks0DNssE3PqMOXoGDPIYnhmBoTDx7HoQ37kEiifxhbgja/NuKxFfyAep
haoDkVHot3TG67n3XLdH5goLtqDGbcPGOZHe2jYYJpolx/J317bUwkjpfCd3BcBYYJIt8KEn0ya+
FQF/mQJo+LVKJxb+opL3UXYNrg3xf6iHTOM68w1xDAr9shOwNsLXb+sQqADjgxF9jucFxTex9k0c
Fn8C03UkZE5jt/Tch1gKfVyAYfTE7J68JJjpciLrH2NjZyjGkKKeoYSBk7tyGNSKN3esBsNnA0I9
LmK57rpVq+Pd6FPvpePANQMXvNSRM6CglUm8o85XGgBJ+qT2WOyIqD68SvdbHWmCWtRW9pZOlM7p
0KcyR03kQQi03/IRGcyoGCb6moy++Y2tODHwEBi7/ufRBJzFW6iLwMR+t3Pmto0wq1JL6hoK6YLg
kYNG0xn9vKcwpdHS1BpwEtFYO7WL2VyHgHt+FMmMnzbpZXuYyz9cTux3gJHhxwJyVsblS148fuIq
jWAGAhmiWApxMgwwzXctrlLVpJ1sro1kZLjosj6KFJt0aYhm5uwgE3mDTP3kGZ2+uhthgvl/zj8L
jPAYAUog4lFtSfMWrdw81Zsj6/xWKp15smMVPVBZXoFe4szd/zb7pHPHFEAZLCwCWiJqFNW6ODpt
jmrXuxoYjly0u9Mv/qv5IJwVCcmDstKv8n5jKRaxYVdGf3kkGbrTGexGzx9SXCEdB7yb+TFWEoTR
4iRn8odZC8F1VYayYQ+Cl82Cxy7Kk+8IiMb1pE8il4pzwsgmpT6UgQaVt8uND99DMJ4wyKOV0tFQ
l7G/5OK1+7B6NYbKDLHwH919u9RtorKDR+pUodStuIDIrnRjP/5gd35qpJ0HBK/kY0CdrGziIf8R
kJeKlQFzdcy/l9kOVPtQAEbXItyMOrx7gaoRMg/IQXXNZ+/MgFWA7CV26sxHSnDzmb7W3YO5YO1s
AwYUEb4oB3fMqOeJ4Bf6n/AxLy8PNhDoDjvAHrKccKytGBL9Fg0tq2yxgKhGVEx4lZgCNj+tIoSZ
5y/upRtpkDhwoXtUzym5FfS5B6w2jpEZICKlmU7H41DHfjY0SuOz3lmU5X2+kbWGiUFoD5iFvdgD
1DQ1vMbGACJVu3TbEo3xGaJ3D7VfKw5gSRJLfJLn2BzTGCZ7ABsBvrfAn+5NaJdMOHlk6qhFV2IF
5en86EABsNEOFNzt/SzK7pgbRZ9iJY7ZUQeGxSw1NPJRV7XjR6fV6OQzPVUEaQ1bUSaiHONFf7sP
2wkoN6El57qM9YZYlMV5xkUqXhbAs9dowYbnrMH3Lryf8Qblwo+7t0tCXsRIj5QiJt+gpjfLDZJ1
0BtJndJU19CJZCaEuEsvbWfV9PbtO7V3ym57/wmRdLR350ysfRmPseZwpqDNmIM9oL3D8Z3QcvwL
AUmfe8Hv61+qGL6A7CaAI+DObJVcG2eVhy2tvWz/63Jaqagi1PWoX8o1EMZKVd/gmvOIa7WcdPbS
CfyZD3YQxKYC6LOwYVCPQLuZp6/L+sao0A73WCwwATBggq4F0F74+h2JpS4wk5CddxYoc8QM8MCN
CdPnWv89Ken/NZUTvmn9xbJlmZc5vKORC7c8kopRVmjdbI3bYl5y1MqsI9VuPPCaqaQZ5TTzXXIv
Cjtpw8+A5WR3AMooQJkKMJLs6HzDsgYA5dVPDGpXoSkhTMG4Cnr3fhJqzWMm2NcKo24U3oSWHuad
HgL4oaoeJCwjZNZ7GlHw+kXgmEtGlYdbrYMrig8I/1UQGURxp3XksBOXxArMIXHyzd2/9d6J6AxS
Q7ZM+x7GMeC44bAbaiD3fjwmt+E9EggY0Bw6MUSeIYjaC/CGJDcNXJBAFThesHPJkGR4AeigMS0l
H7IGeSSVR8HRUMzxm7pzozx29ZMBw6gqGFn9zRB9vFb2pqzHwDpzBpLInseQ2jU+45LwIqXXxayg
Qkoh4UKn5rm1TWC5uh5vqzi4r5YnyZv+sUbUydEd2gVADZc/s90xL2fSVB0P9Cb6tP0/CJTlgKhI
k1NbfxXWGPAeE0pMxNKzPoZVJBQ4hTAQCGn5j8TNdQzpshX05dhVHGmG4Cx85DtOY8pCqGKLcc46
xS2Hlf2+mznif4Cr0iTYCl+C+y/rmVSeYsH+UuLiYvyC1C0me3gqplGst0gJ+XlNPKrxbs/8JjyX
eXngc7Le28WweBK4PoXzC9p7JKSt2JMon7sm5ZVMX/bPrhOX8gvqdZW9ap2ulbfOHNrInE48SMrj
Cwtcu1dkRrM7diaYwlNYAhZ5235VrBcSX4Vw9MmQxfJC+fD1qV6vTe8JEovIJGtG8fg8S0BzpHH/
EoZCApxD0ZOnQAPRW8+ORRKavK2igzQnXaoB+5HX88oZ1sH45rlVGREfx2msmqYB8iJ5R/1KR50L
i2wDqVHAAErDvOkAgjPcdHL7jOapP9cYNJyKdl0ePA7Crd/UJfqaCHUjGfG6F7D1433h9lyHNRqm
4gVFVjFPai3xnvox8/ySiwgUnCVPB86DSaWdQV8XDptbMqCziSakXKclLMs1P8zbW5Hh2Dt76HQA
xLmYwUU8tPi32nFVgWUG+Lc+MPXQyAZkAE1T99W+D/cMW7yLDvORjTntDlsdhQVJaJReHstabhXx
x8382g7mrrOXC7M4wgUQvKMrWLfJwgAkikOkX/giLigkcxItZK/INYjuvJh7/cfORdgJZogn6F+e
BPLqaTOBFUY9CPWwzV+I9b0+xFq7YLm3o9kI6GMAjoXzOXsAKesulLJLQCySwYe435V0qQ1ybb0p
oTgD8sOS1+tw+XBuLX+lvuOOV2xRgc1Q1/uYst6Q2SuH/klNzO2BdD5mHOXaG1mGPZ4hjhMW60Uu
YCyMe4akbhdX+dYGraNOWTNHBIcaD5EXvNaoVolQOv4jtZVLq8fAXD+f8gz7+4mozQrhwt2lYsbd
EemQigOGODXTxJgxWsSZu9NY+bL59XiIoBv/j+Z/j6C4ScDoChFtBEN6RemgJbqeZD0YG5jAK4dW
eeTVVIPerzZ3HfItw7bpsrhRznii3D+prSTNTB2Il3anNfa1na5aUUo9dtObJuS9NMdAnXX564AU
IPlebhzhs9gYG1zALJIKL3EeCCMTh5CeOjNc36hdMyFBkXpRoujMi+e7frnkha7e5lVqXERH1D8T
tPq5OOw+fVQaf2XF4aUV7Q3TSOqLW+jlJx6mZRSl1KkeFsmTFABhy7mwWxaxh2n9UI1ZjbyNVgER
oahqXRaPWdJztZg4yRm5rxapy3qFJTArH64C7cM71VtjxhA23ouf6+h6xh2LPp9QTcMc3f4UeYC6
r7ws50zMkSg0Ogmxkh/JH4xC1o/UsFLCJipc5T+CEvhhuCUUMwvLMyiDQYZvyK9qHgGbatfliGqA
bwI2BHCoLHevZ2cCNhfl4122Zy+gJHrFWP8X60lyT4car41LYf6KLftV3K+CyMnYA9RXpyAj/D9A
HgNdXkO2u8GAhUMMdHLAVCiCgtSWzm3Copg9e8+qfGvVT80bHC6HBU7mACGIyqwHwmi0fRKGdMuy
7QQ5lIWYykGxF3hOvlXD8OjvqFek0tL6Vr/ZjgXpXvBCk7zYH6ilImF1Z7kI2ZLGWU/J4LgUagh6
CeAGMAdNwx0S6VAugI4c0QZclQq4Yw00suVKZmb7Zg0roAoaWB00MiY1NIUUIDYZaDNRMqC7zJ/c
3hsqbYOxi+cp/AJSRlyKAeOFUKMIDnhzl0MHUBlmsu7PMMwf1+hADWWMbxgB0jI0Fpy5HkCJMroJ
Xi9jh1fIjbDJ3mEcletomj9TSZ8WpfKy+bda5J7pT1RXfYZxwdRxicV7B3VqcQUlTw7MwS4imFQI
x5Cvwt9YbGJu0fC4EJ2azLWsd8UQGHyQHP6zLQs6QIEd2AQw2G/L5Eoa8+8DnDjkNZDid1yBfP9u
JCEm5ypqbYA6A2FP9cehzPmzvTFXghaCtp2aBxjmTPRRVjQdpjOtz1dUQ5fsW9N+po9s5VAceYDj
tFL5i2rXiOGr4GIK3mOzRFfD/UF7PQ4HIWA5xgI2hmoMNegZHBbA7VVKAcJBb6OJ2fmJmykylP9G
GQgsO42cPEsvx6u5UiSFJ+EYN5ehAHySBJxD2pth4+AgOo+lGUAuGYuBUxX0dM/S4lQvbcRIi6Ad
973lcCLsJryxZB8wwBR1Vjlc0eufQ0HNZPLSDNtJX6uFHJy2I1FhfGEw5Ioygd8/V+HKFbDLUZ41
UnF07XLv7ggQk0EyVDNVTkC0l74au2ej/+86nU1jWk45ih4SBVL5uaen51iT2XSZKQ5UZUZWepQm
RZv7qDih1lG13nY6q2LT1mHezAiOwNC4u6S3E59MVBszWbJY1kAByuRWO/WQ+kw8d3Wu3qx1EIzD
5/4Zj4LaYw/Jb9P/JiTBZm4r5SLrEDKB3b9x+Ip0qI544CmluZL+mFg9OFumHqtwPxxj8D+XkAql
HEjp2TQLLktDar09uqKEkXIvkKq9XW72Sn+CerUwgW9ERoAHe2JUlYGplBVGtxNCyFrk0raZEdaz
yi6UjPv3ZZVo+PKQJZvmvPy2vU7s3PpCYLFhTDFkZTOivaC/plUYI7uefw5qu4k9hxlZcdYPg/a+
XYdrQYjBGjxRiO/CfmbAj5NvGQzDefKM8HXtw2cfV8GyRapmHV0A/p/TEtEZZrXjL44v3Ig8Bd6m
M3FdlY5IK7s27jCBWStF2cYRh/86kfiglw4JPU6/GzRfhxkCHqnqVZeWqhNOHSHc7ZctPxVZOhD2
FJXLj1ixq3wdFVWDvsbww8M+5F4sWi3LE+Qw0feU8P5Zl04Tp/iaEViwJF2WajIeaZ8slit/JAI8
1XGSelRDf1cDY/j0DtEExgFSGLMOfCrLfVb03Lz4j6iCkJPf6Gn1ouGnxLg0C4VS4lCzEgxlpdW3
LHhcR8O+DLMGjD/XXrILEPrPGnS932ZKeA/4Vu401eXt+VJUs1rSSxxTyM4jlU4hxBTRxPlRHlqO
uYHnqkNKtWXklwlCDjqXOWPzDVgRHBJdpBBjw48NFboreO/06YvnzFj9t6tKxjI3mDAwcJilbflP
dUIhvuyN0AAyI7AZ7Iia6+RLVbID18UvS0kWJO85dwthLz3ihl0b9tM6ZMjx8xE3iP/s5UGXoMS8
yELXpcwL/5cTDCy6NH4miHCXTXrw8FWhNU/jASGnDnShz0vKfqk0AdrCxB37SPixnk+qQ2hiTK1s
eLe2Lt6mR9wlXmoK7XoDYCIlBOaMonOoiZ7ETN+knvKIKz3n/WqA0Re9kJFr0onkyQu6/8EjwKxF
jpJUwdoXkJ/M9gPLaQFwNfxNGsyzyxHSAcwjcUspc9koDGu9Y5wqxQDr9+j51nbSgOJ1kcqbne1V
lO2lYVxrWn09wEyVAs8f2XPibT3BjcrqdIRlIwClkSWebzNGfrxeH8erblxTRZeObnUgYsIamo4v
euaZ8mc7HCyWzkupcWV895sVpnjNKTi8q8Y6biSQ2566xphbZjm0SbWSnuMQQOnIrns0hqObfgfw
SZEHtNdBYKmlbAbLmZF6EGJSLIcSQnRykUlzDyECHfL9DV8jvmuYtdW9nN+GF7ZyFtQqPKvrCyJv
BS+vlVsUlGI2KKKDOW+XgQ3gWV7N4VKjP03mHcb1TfFj68u1Ryz311PUP5WTZk/jPdqxn7Kin7aT
VNWjhH2KUXwmI8rfUTpQgXXlNbblangSiXjIG+pzxGmPSL0Z4nF43w/CnI0E92hjYEIVVp0/7BGe
j/VE2DHxRzI1zDkeVnJRvy2HAnHj6bu6+p87JIn6ulO1qdDaul9JBVwdE8Y+qthwM1NcXFjUd0W+
BQ0LmrJ1y266Z44y5Qhh84taxGTH6mo+sMLH4Kv5IuN0YFEeH7amYgkTFSTEodrfO6p65kbQ9FHw
1XP6mbgTJ8seZBDD1RKYGrblGmIJQPwke9vQVDp6HHUDLWIcM5gb4vq9uH39L0CFruW3qtIug0Vb
yllnPOMqi1UevG0nLZcR2hoc8KJkRZFNeq5P3Rw/jBRZg3vbzPP278+R+DQ13C1XIVN71xCqc4L8
jeLDhJ6s0pMcpOA3aVlZxLe5LsXJ/6JA0nYDy5M9mq8JAz4cVPjw/SH3IDQXOqzTIMPjYu4gmH2/
X/DfnEAcRxZRzNLLrnzBKLrsx9JjJjwB8DelxClnKJ/lLpsi1PQ/48CO4izPQXsPG3ydUvm1/+eM
OOU4PLdGnUsCexs4iDxORhnn7eZZPvdowOkEPRy2moi1HTqgqgNS74mZgZLB4l3jSiJe8Reo3VpY
y0q36y6DaqzkqEwsdauEdv0EoYI3aZV5cHGzwUqWEBghUqZPiMsydWPJxEfo1eekkFESqH0sniU2
fWyxGZB6bs4mb4WGbpUrUsOnwZC0XlZ/NSN7U2q+Ds9wMxcCHz5+6ea74az+e0vsRipDqo+v9HN6
277SndSJ+0GKTEbQ3BCFl8kH5oPp3xtdy06p5xw4Bh/rFjaSpN5M3wUlMnNQvS4IIeEgW3x9md1P
OUrkeCHMT64WcatxECqZkyDSf2jncOm0YL4uhjUhJloMb2Xqvvp/QL9VC59vVK8uPqPDcjog04pz
Q6dkPJNfHaYyoK4w6UQZaLaaJoiwjpTstLQ7eSNo25lYgCUy7SM650bN2vnIPHPiJ6aghJR8+827
Nhw3bz6MnjNnZ3lbtrMiimInOtyELhKO4QwIFbwSW7eznepxxh3RPkczNp2i0kaA0dCGUPwQOuwX
0hevTVRsjxAKbLtXe5+071mYJsNqlxd6UH7NgsHIVArv5uhiZCgz2ZICnIGkVwGECQaVOIT7Aj7d
8HmSkCwoj8FxMnaH32SfBCJ6o9dbS10ojha0c3sGjbcnB1WK0z5bB7dljUk6J4lU2qBYrRR0N8Wp
luDOlFcR3x0qtlYTlp51JdaZ4kJBXUDEf4FKYmK9VroYwUtDIW2FOqvcrOU03hBf5fEVPvbWLbe4
WJ+wDvML+VFQjHpnUfSQNqUDThh8t0jOq4nBnvfuRcMJRYj8qUcWScaJXBgQ3Cvr6j1QDpaMJVHc
i/gqFaev20xXYg3TyYN++BJBR9s1sF9MzPG4SNRDEiUDte7K3Ek5A9RNkkY/J8m0Oz6dSm8GQJns
brkm0kE50HKXMhe5/oDU3LpQh1zRsnDV64mVWUjFYIfsHWW9KcnbP7mBm0c83y7Jly1OR2eFx1HE
RknEjiRlrOplUVQh5LueDGfFwaNJ3ApqajtCy4v0s63/rAwDZbl3HsHQqWy/16UH3qdjH+DrAWnZ
F004l8/oYQRU9/HbzxO3P+5EHDMTCPel4RJaMHgEIwE4s6XASTMXev8NkT0VITV+sb0qZzlcBcNO
rduwh7NVj/AebuOFlUBNAtbGlKMrtF15n94ja+/ro5YGPtgXp6HBdAmBRoct5/OcE2mNXG3YhLRl
daTOL5f2PDbw3L/DBvdhEhSCuVNIYVNaC/Z71pHZR0k0K48iwXDKcuLSziNTCLqam1xN86q8PTCU
2ugVijlmO4yajP8/aow4RUNb1bNoxoGfmLZe9CpzEhrJlhbEOLJRZhxrf9QKPSuyX0oqMXMhhlFn
qCCOPHxMzCErHhIBkNZpTdcmXTRdj8vsQavr+2vKlvfqOJCEYuqcWuuOb4yqm9GaYZQc7PX19n4Y
KPt/WXpj9srFJhdqtJUujjNxQYJPkqw1veqXNxtPdRzC+88eymnNeXS8lxt7ozh82543m9h6O1sm
/yeDARdSuDORkvAg94F/6TyOT4bemVqk+rLcBQDxjn3oXdlo04I2v9gnVm8R1oOC2zOlKs+hf/7n
9nrvSfJKvht6HXlhCr7WZLaRrQ0vg0k72tXxSoYljQWTzZ2s25XsWnwJVlg0EpWvsVA3h1fx6OyL
e8pworttk4yf+3gTDxSMo51Fb3UgW+aFXcrPxb64jvsdRShgdd69l2u3hb76rYv5DNAlWLH5dVjW
Zk2rNdBSdSQZ2ln1kH3TOSDjeaq4+B2x3MoL+fdqYkOdstI+F/aznyTeAHkmywyb3qyq6O+nW4/c
rcG0oIxnaTcoGv6t+GKBBbbQFksJQOeS+k5LZ0pqQImAkJI/6h1SrEGBhNhUv/vgAgPc7D8dCjjU
74+E9jEFWjKHDqrE3D1EAeXoLrFGK2cxEHneWiMKnhZEkOtSm3MBzBOCPnIOcW++qpah0xYvS0gh
rSAzowbBCVKFUPj4R5OYC9y/8SfUWQh47OOVjfAuhArJPgmo/0TWViPRhGFr7ZGREBMbK03C6SRJ
8C5hXNB3xD5MsxD24buUsdDDwP3Rnddr6HWnI8Ux8XjIHuUgq2PNqBihlFqcaYdZ8gVjw2TS31+W
uRGJRU+ajMBO/rD3VlAqCdJXHRlx0Emi5UJvuH0t8hH32Nu4kN9mFdFGl6SdbMyiRJE0wVBb+7b/
QnfMeda3MR6dM7JdmOKWp7gIF9Jkc+SL1pcYhgHlaYrabK64hZuai/9gqFkAp8FapKKTdEuq7vln
8CFhORKs7YwQPrSzMIEk4kOGgU0gFAigOVM4JlK8vg6LjiiR4YEG+m3P5NgCcUUjpGOolyNL0U54
VhKPd+nPHy0diWzYQmCJSleUBfLV9zJlLNT9nwCZDGi9FGmMD5POyOL6IBprK7ocIcdH2I7/lf6I
xMKk7jP5HCkzW9m0TxSX6CDsIJMvP6jm8qsj7aUUZFHG/GH3ugKDF2bX0P+BRXGQUq1HjZsMFXt7
SG9zbVjI9OzeXgIPTfO23Mj8cnRRi0qLc22f2zhWwIBduINKgiO74hXZj8eX9SEPekOPfgfgSymN
+eFE/xSqlMnhpRciJBEZYG0be8+rpyarJOp19cwP0L+qIcUvTU8D4Vndo2Tt80NVyFbNTIKkm40q
ej0y/jE5n/byluO3Lj4CPQLe1ixk51po/8/a0tJC1ZAh0QGi2UW5gN2wV4VF8VjCK6kEMRq1+p4d
yLpF2TWCN2q9vI0n0Q7c7iuXt98Oe4tb4KSJ/aU0HQlMJlHabwEJcOzjZ2hWSirrUObw6B0LwzXq
aqpCdYeVe/PafL423rb66e437g8yVBKbTMtNW8rsebLX0jcxfojSfrzgkdKeZphwTRakvdGs8cI8
doH04tzH0SbvxqtnFzDUKSNsYqDvRvfut8UyBMCHEobgairLTUsptErjiSM2UBvw50ryvynxorub
6JTMMCf3fZrfP1xQ5/Qm9e4MnLnQ+WMn/rEnG+OjwgUSKRB9tu5Gdt3V3ODX6rd4EKu9IVyUGEws
d8Lv4hEvR1ROp2irekHChzLf7dkougbdnvnm8FdzlyHOihbpF8UlPbEPE5giVKRyO7U9LoWdKBJK
yi202OLaLrWAAp7vAmw3ynT8yPSbKp3vG7MSawA8VhOMamlPCoH+zsJXFybAGQpWkR/LdhBhe41F
R7jp2qZ9byt9S/voGU+eNthws78yh309F86zi/UJu+TE1cNjiz1cSgA1Ym3uXRJv0EQu9K5a3oad
4bmO4jc6eR+mvHNVSN+WA7mCpz5EsaGgS+5JgMxzDjiZk4ZrLBiNlyfr6l7QOAUrXpRjbX5mn7W+
f8rOIH8q6le+DzVosD7K+6UGmDhBkresCVxAM69BWSy5soildPeGSnkk7wn7Nee2YKAr0ulJ3Rs9
phgPSd5qgOFxtzRXX4BlaWjypWyh6RYxIw7+PWk0f5tzHBcW6z/7XO/YXJShKe+ppwj0LGRvrTUP
68m9GNPxwPWtiqdnFDxscobuTWWTso63yTIRPXhqSDdlXebYrpZpocMQ5BrWc2fTakYkzv38RSlW
rD2ptH8zJKL8KSQzUbwUkcbEWe3oHjcbcFAyfhOORRNn4ejrpM/7ERZBD8+axMcVj13rdRYHBk5Y
7r9j9V4iLWBnEdkaay+N6vhqh13DWYVmOUkftu01hS327IfPxewXaps5OTaAvUChSzoI3+WVxQkK
7u9L1/ybiMY1eEtURJdavl8oA2EXPpnqU69YfIVUPFhUwXgV+mtee6GVID6Sek+4ikE9uLzL7xFR
huAWtFKM0Pr/ksquzKSUEFiL+CsQjGr+E9bMcUI+Mi7DP7g7vdWuDMEiQsHSXKP7/KWL4/sK67Ic
6pPbEIDGXePo0KbiI5e+rZrpDV/CHn+rbddORx6QoHsHGJMrd9MNXgO98uILGC53uZ7M15j5AqkI
KbjR8m0wJWoSkssr1h9WAcnB5K4Gy7gfnlpMkvIWpY0jszVf7SmmnU6kZcsjldt7KZlrwphLKooO
q3BSvo5jQzZo9TI3FTDKho8q/dA/5hye9nUYqflr+YJ0tU9Ld+YFrBIdcG4rPB0mGZQ4Ud31ZIzm
4d8qcN15FiJhzZVmPUkgWYDOBIw/gcLncKH0sDoz2ZsnBAdu8zpcJPi666Bcr9Nnl4UP/lwzX+Do
bUVpH+5wKkZZXBfe36mfNwetC/GnNhrTCF9mL+GEQ0IIN862zXl7bXhvX4QB8LfeDnAQIZGyu3ZA
0o0jLY3O421gm3oJlMWZRbA9gRT5TEgDGUK3B0pUsiBIJBYXqEhOJe8hKjWkWUa2w7FRTUtx9R0M
IkJM3Fkqo0ZP2QFGlEUEpJ+L62uAm5/LvMjyZAPj0JmwMAfsJTPUzJgedDWeGJw4GBT9ibR2NL65
hMQQXkMkR224BPjEFnGE6fG7ToTUxfl5cF4P45QTMJl49oMP0/ZW0dBXD97vWrsNwXJmcKM4mWDj
Re/beBrvLmVEWbyaht2zblTvZdWbf2gkkcHQf5HE9UqvuN8o1IsmlHfh5MCn/TTLCkExvGifyNFH
WHJlFxzReq8ncRJkcxShskKIAq5uGFwfyXp60HHiaIH1YC9GtJ8HCMEU2yjuZ1+snyrng9HRBuv+
KG/QBYyGdq3mg+ArsD5rYhNq0EkTmVeuAXX307xGHQT2I/lxBjnvktQCJz9pXVjMXdjMIaiP+6Bg
Hochc/vz2dqsx0GSigO46W5kFqtNKRuKj+s2qn0dpmWcfkqKt3SPOsGdyERvcoiYGQD1kAV/Eamx
FyiHjzW/+wqlUkqED/lhg733yQxSrwLWJNiE6QVbWi4leXegOOfg81dgVmd5d9WTmkvYZ+xY7P8t
WFPvZVBDvh7mAd3hNQ55HwNWZ+/MKFVKQV6Fi1x9gzNPq7r0x38cKFHjPPad6SdvcbGyGnTptV/R
Ajc5NMQlqovYnijg0V/J5uztnaC7G1sA+hF3mF4wG8G0Yn96OTYsmrL2kZd4Xf+X0Skvtcw9l4wQ
XLH+q81gDu02/mVsZYUiwjp3rnFTIyQPVtknsiyBKz/cp2cRLQRIuGJxpLBQ1V5wYYRedJ9/wB6K
7bKx5qq3IHWkvXHwG5JyNcOtA8HEUVbWi90n/SCnckXTK7OGOsqcyQ4Ah2zzhYvmuRZZmaBFPmef
qwwgXVIAx4chD+Sq2CYhBsO4ytzGutObBcuFW4+bc83X0lFSGMKLCiuTSNDrFeHBLxDYqBSfG7MO
v3cQ300s5R0hhylI6ZPDWs+qm2Ioh3o2xIH2C3OXztOg+5hlfQr2R45DkgOihc+ki9kYIK0+v9DS
VgD+NXk0R7yLHh+G84tvw4E5KN5pTrCzaWOIG1b91tX32jR92o1GMv9Pq7/eRSc+hnZp4hBvSQ1N
2x77U1OiuFU7tpa0piAABy+EaaGKfs2AqzAs1GPPMc2164zTuQyUH036HawEslkPNYOjvOLzzg5T
l1MjNlY/U2Ubcdt5W7x3AYk8YfKJ1QPvW6DQrzE1hYM/OE2y9/0JcD/D2mAY84qoBRduSUdGTPPZ
SI5zdRGQuqHj8w0IunFc20j8EsAWa+WVTwMxy3PRYu4WmrkD7N+982iMIBqzQ2LafhgnBCwFwNaK
aYfTQMJ6STBLVmI+WgM6CIOdiM0Vu34+tOImWAm09rOi8SS+40hR2+lI/y9elCLlOTGgCk7r/JIp
rbO/H+/AjG2KDDIkFGO47m0y4JxNAcJJ4/+LKEfkSQ4xcaVxXrosNSDiDQxrU7lN8as3ORSB/B7G
ZGMwZ2trVEs01QsOJZ55p1f+12nurqDCn4d38mYan+dv4oL7Wri4uoHSRumjFQP7LtFkKixejklv
Y7QXUUzRd3u7CLMKRUfMH/Dx3O3vb5vAxr5wItcsMw1+T7IZR7sXtfO2Iyf45KaFoykUdz+yp7ej
ug27XhvUQn7cJV8vpV4/U0WKjKqtY9GQ5WSmVH+syUtH9XNy9IPp7vbbr5rLAWfVJwb9RpS0j1jS
njyropYYgxuYRRc76A0c90ozQvdw6zaExaoMLf02MrDW5n6zwr5iSHxBGqWwlK7XUAg/NL8edpDw
ZRuDE1xnyfDZMQZ8ihTkL76kj1z9BNwttiMojfH3/PVUIlGaZJGOxdV9fVXzV8r0X7MqTwJk7/7y
e3B2QufiGJVwWjTtxnYMa7DxzhdveSbfML4/7yQqNKwicbHj2HGK3H/xFbgXUnfzCQhzguQ+CMnR
R9PPi7GxYv9XUnIR5oHEYfwe9eFQDkPwjiCFXfN+avu+znoVdkOmaJVkYn9KJm1R/PBVV+dNpklJ
IyS8lWfQhPPFvXKTzRya9meOyHRy+dgtP+qUGvq6Nd9wzCy2WlMXeIrk9dYqTHjSRiEBA8QZvpG8
jQmNYkRlnRuucQrpuCkG/rX4c1tUdGGlEYYc8t7zQ0wbvouFUtO7hmVYRXxna2IOo9kSD7wbQ/jA
aEGhF1cQzsHWoSjWlxhT3chWfHjtdnEABdh3fQ17y+IVZhvmEhpCg/3nrmbJqapjQx5cYha5R+ot
P3k+z6qjNwBoL9r9PXj8E+ilBjZm8pmB5TakSRq520CsDLqlNqeusvaDI0YckvCM4HQWBiZhrj0Y
JVbVraC2dVNYgL+ucFjIlntRWewFjrrZY27bQYoOFq9i5Ne73ToGGpbDwuANK9uXR+DR74ktVLO+
+IzT4eZDQZ80mjGYi1f/v/C6MI1AxFSPgVqIMEzSRBtZObC1rIX9CNR11sTTL5lqPTlT4ppFNiLb
MK0ycf+XGszkDmHnwmYKiW1RolY68jLKb/4NwpinyyOSubLqEhO7kJ8npK+VXw/GEDlJ3io28e+i
lx36/4cwKJUyPegB666efzCZGnckO8WpTVYNJntrR1jZjCeiFTzzqO/m0rfek1tmO2WCgOFOBBPk
+CouP0J4Y759sP4qIi5NXJIm13mDmHGlSdSS0qcKPG0YdAdIrtBDJN+MRE3zbPAd3UL/EmjI2CYF
MEmv+3lSUG/NEjF10ZTxTx75pHT0LQsHQc9sWEMHhxUEw47UPOXVAwY7/idjmDqfWAg/CbU9rnmM
I40yLh9sxomsg06EH0cH2vT8MHb4WWjNkT9BAG45mVWKd7KPbVLbeHRim2nJqA/izTecLPlTh2J0
Zj/Z27FKITXBLQlKzrFAXJ5mfJTy4t8GVXG1XGZwI6HoiB9t+x3iVk2EoB9oJTvQ5nkDZVaCudqN
TAzy7AHQHrGuNo1gp7fcrWx4LyLo0svhZchlc1lKZoaFBExhMy99/3oZrLYhBt1ewlt4zkXIRKz2
P4/2JPNg4O7FmP908XkQkmUTQkNmXNwwH/iD4qpELXM3Wo0+aff4BX5lBs+B0i53vUQ8mcMKv8og
nQ+UvMqv8GWSEtFMS3PvWZeYU/eCphE88lyAYJ04/CrFP+01yZSHWaTRT++L7138uMXxoQ9KRdhv
J+sYOg9UVdkhZeWDqYNEdT9u9LBJTfDXtw7rmmDcuxE+0NweClu4BuMBsnqxeGKOEjTuExC1fKLK
UAhEBF/Afb/NMh61Z9+zYA4XENuan7FtegrjdxMN7ZZ15s3SdHCrMnEqNDSUDpwut3eO+POeLTLw
22bhWAGQrk9o9cMACVCiZGc40GgZ00E3fc7EQVgWtkipGhR4agDt3IDXvm51QwzH/ktHGUMEp3rM
SLlS+ij0ZdZGyfnjZxOsUjFSpBkn0hPOI7mtn+VN44YEz9fP3DiRTbNbUznrXvtiQZIHL1uvCdA9
VfMNiO0xiobQrzxOL54NkY+bkhW7NhaBXkKaJ2rwkW9/B7FkGIR8BqhTxUdAv8OqRs+uyXmO6gyF
CpG7ny2SU0XG1TAlYO6PpdC3JFG4he8dlQHVbh7dTlydX5M5NMQNHE0+zSGWIvpznlv9owU0GWkI
1koHFDTngSIEXkH5ubnZ3PC0rx62fMxpiUk/ixXyf7ulAmbNAmkRyu1Fm+O2q+kvmiZKlL9cyf0w
simHxD5ducxLMC79B4nKeZwJfjZlcnreAYA7RgAY8oYtdGapo/3ilfRjbRbODrptGL76iXaa9kF3
LNo8o4hZg9yakOgVJKE7YHm1Ovqc0a/3l3KMlezCLT69+v73u4bSn1l/15ThMjTlE1vPiPO2y3E/
JnsKtFnqm1cuhk66dngcKTTbUDbRmpOU/TrqctIRtTc/kTbU/tLSf3eT7lP5X3ocuEl3XuXaQzFK
/uhGR98Y1GkfY56Qp94fm1kRmHY4k6+lWngJrpFC4QkfHD13NFSaTPgJCDHLXypMtJGI+5RYN7k8
iCrAA8kwj4XNIYFHbcA9vrILTltRlj4OMXu7lmNkwWauNRBBXw1Ts7s1TSRSPvjaUkWzTab7yNTx
koJ3V0ORHs5EQ6NvAMZoAtFjdtHoLMjpZJ9zoLvNFdz+mMI/daWeOwyxfckJj4hnkjzqafJZCJyv
KXQJfKMZ5LcG9B459ehcnfvuCjB0wtUIoyUvieGIKXJjtNqE0j6g5v/YbjlYEuHItXWlC0WuwL5T
Mx2vKPBiR3uD4Ax/AlyHg13j7n49wLcA2Zmvq57PJo08MhHJPfNCMRSdTIUoNcmPBzKFdb2ekuJI
cK61jLY2PxxBPPbydK4u318aRxBgh/EfJKwCIsXPBnXbBRPglkV2rkXfG+MjDppotIuP+012Tn5V
BK5hcubzQ8xP4ykoihO9YuEcmr2oLKnQi/D2ZVU6ayphQgbspjJV/QrS9+N4kBuGJDwF6tkLjrhK
NBJHjVO8r+Ki7tnxWa58xCXZDLlqXiyj2s7aNv8iatPvjFKuY7sC27+Y/tm6+EhA2Mem6mAL8/Ul
yqIEKmCAnoQb4pMFPiQ6fyLHmVuhy4JSdTNJu9lK2eJyxrLkhU5+RKZvpN+2UeIRG1fIt3vV9SfG
W3BKFUXAL5vay5HTPqxQzd0fTrs+mLHvAiFPLt11vK9EmHzihFz4A31zBeqdmxtREdRTj7wyzCel
Tu9OsoOwkkIgxp5kwkhA0jhKQmSlaafbP+iQXv07USN9g4EyYbVcgj9AhW/yrx0f6ukzK2lPib7A
y4KdBI0AN49nu6nKom+qaJGcfalIoq7xaZCFEBxjqsguJb5P0tNeEUzt7nWaYN+UmYe+TNTMFuB+
MIBmzICYytKuNWe/MYNAS3CFPOiaRCo/pmi8CPYyN3qQxQKXaabs/G8lV3ncw6Qj2ykjyOPCfgSJ
joCVdR+pQmm27XJlCR++H4wURNtRX2UX1a9+/CcyIE4n3ptVudJ8W0k0BvTx5zgSsY8dymm1zCZz
SnQxhLaDbfW6LOzw/7o086yT9lAtOg07hT0XdhVRXv3h/5RgkpJfJfM6lsEBl37itXta7BX7FYNy
UEYqIrrKG9NrJeAWk3WfOvc4ORNm9gvvlYavDtyXyeb5q+R5kyG487aKEUE7rVSRBh0GClJXfFQL
VKNVLVe1wOdK4fIf/8+pIEdc9vjxdEk3Lm32B22pSLht1P7Ja0G4K8YrFo8FXR9F1CFyy0eg7nOP
aAdTWSDzyEMD5qoMa5mKY8wNKE7tU0MM9G4gfnzrKmp9/ngbBbjehT/B4bIPnQOlxhBsxeD9H23Z
JRcFcjClwyqwDIAtWSQLvTFwZ5lkXCheiN7IRVqvJr6JW7+ULVMklx9QN/C/iwEvyVSLDPI6tG9k
4PsHUG7arescf4mB/Ct8jNVnQ8GauS1u7f00rrB4fXfUGY64obUhLKHAlmbIvH50T0P0ZFA7HbY3
i7HLiHJcejbxttDwkjoBL5LPUgqgqbD1ohE+GxHGZwKcMIiwI+MiUGDpLn+BoHgnrKHyC2z8ec5A
+sYuFswMrvRoDFYDPxUoyc8jOl+TOxHzy4LD0rDjGmGYYYeOKGRMJGWP3dj4I0OHAY7C5QvD7g7v
9drofU+JKQv/BgnLxyrV+G9ivcdkybmxQin/cWAr187cl7hbNwhkHKG1WdGL/SkZ86XzuldBJG7c
5GvKUYtY0QdnahyA20D4hVUXNSv2JXpCRCbWhP2c1VUI+FeY7BJfdKKOKqICem4BSQQwx+jMHXe2
HMh25D/qB3ppycTz2XZI86h3ZWbdg0I6vNpxI8OFqrevAmnj5qfRzWyBmcsakBskfAjEXopkGQHL
0bVP/awdFFnwZafhcD5vIPrzvMBY7PjNLgQDKlWyOjsTXZBJ9KuT8/WsfZfgMjbpKwWV8jLQIjkt
UujRPazFL68psBcp7Szbj/if8Ya5kRhKtV+2+lNDzLcqLqIE6RLBnDJaiXituQV0oC7pbJ56fIdZ
m18sG0enxtEzYXmoOqnA1xJwYWV9VT5fR+ggAlmopqoXUftbI+jfvp0uAbslrn1N2LuuOkX0iP1W
2SHte5xuJxhkZGBiKs3ZJlGGvcI9STy3O8KBOeWIxwNmELajSxjSoGIvg850iknC4ThoXKagdxTA
yjGTHsOh5epIya0ipVUVIzBs29/9o4WxIksW8M41inJwITX2dn1R3ltsiBgrd1vNAcjEvgk44JJY
TJ6mu9hKlB4HBs2JbJwXVdFmt2vx7yYTC7uToS1MAuAfPln7V49lk2IMGqroo4w8hk9AVc+ICZNf
esqtlesPUHiMuHEscoh/v+PyXezw0KMUm/bNyeWtd067N+osOr44vwpsRY0ccLBH/0sXlCPiP23M
lQmvcDnKNUP5mJpFnmiwSngjiCvSREewsCE3y5h3Ok6Gz/2n4h3CkOtx4ivipwNtz+iw5LHny+ke
ZtuVlafIewbqi+M74m+QCKapn7/4+WZ/6a7dB6li+kHwQYD9uZulY99gk/SZNDt4vHuf3zb6xfA0
PIpke2FRL3Nw65L0wO0J2qNf6kUA9iNtysHf2N+KuJqXmcUJAsjAKe0MFpSJPRn/e2rCHs6J18MI
ahH6/nUdxDv1F7w2cU6cUP9+MsF7fVVZ0Rzz3gqinFurPh2qbbB38o/H0/+Q776q05854yBeJHdj
9YM2qMxwu2cTj0f4tjwuZEXGV3oYNIYecbskqgpzvSWAcc8N2qg3vTD4adZd+bQFDe152kzZ20Vx
N33Gexr5PJO7uF6xM6Zm2v/QhKJI/KwHswfSRYmritOJuy+uFfUI9EijwkrVCpT/hgqSRo5JuWxi
5YyWiCHMMKbf4VdZ1Cg+THlkoauvJh7Qv6mOvELEkSRK4m1duQlwkYCrVH+nU1XaC+CJ1VlgRoJO
SXcjXmDju95pv4YUWiJ1DuKjyma9TaboeKk/9XLlQZzrNo5s7fqjDQmHgEOi2l2GqTAu8v16Mgqc
W6INPLFsoXBhBHY39ztwzr0TGa828mu0liyyl1JEmtOB6ZL+P6v7pjVCw29JSchGq3J2y4SzxWgM
1iybbHOl+2QPKAf5azP2/iKadW3vpcnnj/7OHN1XoVZA4U/kKjFz7B9/04Zn42Mb7yi0lf38MvDJ
mcs+oVcvCHOxW8uSlgzHizzvUK7uy2gbMPlQ/NQ4xDv1aguydWO8f4bOE8vW3ulqmeFcI1aw57kP
kgNdJ7o1lLNQxR7OoZapjP3y+7BoCOpHe757kcd9u60Nsbr+2FBCha9dBxo5jpqyFG8xHWiMFtbK
uyji/twg/0UqJepr6IOQdiLuPRNyRHKX+oSjr03c55XgCQB4wA8m/+44uXhl9fCr8yXPB3vQrkyk
Km0yXXstMcghQR3tFuDJbFtmNbpl878JSvV3/kO17yT4+wJH/JKw1GoSME4VfYNlBWB03COZuYth
eAOLsZuaz/WovlVEgpbmLLtyEHvpd9ECc/oqheRt4FkHFUydfLUqz1ClvJ6lQsLtqxGjEghe8Ieg
9FnsZXAWWtzD5t+e+GV5k9HYqstFc1ZyLqgpGVeRY/NUUTxkw9tjFXcDnZhnFGwjhIwAcxMDzYaI
rom6uf0zVML1qX9u6At5t/8/QXSrX12nqOT9U5n7E8zvWNBLkSSsNPvFTXYQBPmY4a/QnjJUzXn/
wPWUN1+nLS3IZPHfcRuGRWvtCas5YEJLwHzu0PNLXHFneGRCDJ12xB2oqyII0cT6UgONVpDfuTx/
nOxaBa9jN4XXcyXqpCpBlFlz8o9UcI4KlYuZGY1jWy9vCqFJqIa2WSFSXRxcJhhKvzjdu+0Ksx2V
UpP2AAO3GoprC2tJuueSgqiJ5CfIgZLOck5d8SnQbYsT8rK8FuE0BJses0Bag/lbQW4q1u9gZlA2
kVEy8BmnvTRKGosaU4vLqKDxCu0UCLOhM9D0J8OHYZyKjn2Kn6C/P2HDr6ofpGVJtWi2afF6tbRj
xD7LKlS/7AGYGwOmUEiXQyaTGLl8qeLbxCVC8EKmseQ0qAt4qu2AUu3QDdA6WR2kO/uNIJbrCvwb
pLIyC3pvuqdR/SAsIcC0R23nKfoLi4c1GsosrRxACO9OREAiSFa/euaonZvOAlVDol3xVXvvuUdm
uk6G7ZoeGS9G1b9XAF+qSZFk1zYPlRkQncnA2Si3ggYN1CZRybSiSdS5DS3s7C4Dh2Mv23Bx/R6m
3eXTvobJNuOVSnD9ZrvMcYx0zmdlKBUldzKKFDaH3U3Ml8vU8HSHHvlO9GDlRVvEQJohEhxBe2qO
WHPd6p70YjPE8UeLZ38wcaOS6pYd5cF2jJPLFUqC1GGXATOVLmM7va1DEMx8FhRhIpfKkBrf0Q/d
27MqEsPK6HfQBTj0pDzzRAFarVBX0tNK0qG4ohJQNsYJtq/6oTnYIVgEeH9dlSwoBL5PoGSsJ95B
aPjKHu+S20G7zGjYEXJpdrIyOGkANErCMUy3+lfifNS1IvO4O1ydVhCCdlQN44QgXYi6eOQHB/rM
SGAp+BLgf4Wz5R0BZZTKv54/f+JuIEWU41CyK9sayDVEQPLspcWR+/NwJrTrQ4BiGhUt+Vg8Jsm0
HgJrGOWBMNGeR7O2GJM3rVO0RJ4JVkRig1BxjdA+RoWznRuM5xWoEn6MgnX4AWUfJgOy6MNjVhvM
f9maXonlfG8yurV0e6SxjSaBkJRz+nirA5gBQpYQQ2ssx8u2AwB5EZchm4rJcf+zeO6ll3AQAbXQ
Vi9LiBnPqi0YLm/eTQSVdXstaryj6ZuOHQBlhcQXoBU4JnDt4E4Z/JQnsN5klNP9+fWkeF2dx4HA
bQT04jNniUN+aczgRECavV6JNN2xEoixTIvWUiYJzZNE6rsgYkMAaEIWznnA2lXkaGJtx8I1xe8E
WzV/VlAxXsL0ka8a+TXp5+R7gVpdT7IfDbzGyv8z/11RQKglzIvm5rByPTGxRZMidDsfTDgdM5tl
n1mVLkABXj70xTGTcKMu7zY+oo8w/+uJWYKcT3nYpBsIwPuX/5z4h3WgKgLvPeGFm9BpS7feTpDg
Mor8c211QWF/nCSCQL8uwCo4iQyRW3B43eqA7h3BfPiiFwBkvY7mHxg2vVkaiLmAK9GLywX74H5d
II1eTgB5Wz1noPNcIR6MCMoSFUxZwg13pEtCvrBw0tQaydM5NyhTL4W6JRB+b1tFb4LMQHinDbVd
z6BpBRMm8NkbQpMT5Ac2t0wah+dg5dekgl13/mGM89Vlz86AdO5qNMAAF1cNIjfJQGQvwsUWKJ9d
fI7gBTDTGjDIUboSydUx/PodhzY8GgOTN9unSF3C3F5MN1TaZ794PPK2hgsTYpku9hX1mZINH6Fc
YaMHThzDkAAfbXUxETww+c/AL8DZbv7CCLfSmeRS9Hhu0A+MvB4RCpBeJm+6BVP0uha5iwJ2vJC+
usvQlf7VkqeISsznq3wVVEg9IhICcwL82eq2+lbexvWWpMxC0vO9UK1lERuvA5mnftPqKcwY+dZ/
ixbp7SP/9bxcBf1olyCflSEsG3Gv0b9AvIm/os9Rm4lCufTVhV5wad7dNiZnTxJ4Fb7cBsr6MIG1
lZ45ir1kgx8DnZO6WC8mmRKt5v68sE3M3diKnoFjeXAbObl0QcAUkxQ7A/pkwTAiUFX1zUBdrX3t
kVq3ooxTfkIluKt3IJtbm/w79a+rmPM4MNWj11szFxE4a+znJqMIAuCwAofvAQIuKzEK1J5I/D75
//W+w0mDW/t0elV256/Iwx3UIsq/9jLXdGQl6qQWD9FLMp2KFOKUV6U4Eno93tkBZMzDtIlM4Duv
twN+YQMIEvcisH1BhM1cyMiuLdQyswFBpINzZkro3rmrn0mAQsSJXD4rBjAKSU/bk3DOaPnHX06I
mLMnbWM76Y+/Tqgg8mKYYOtTnCRncriQyVNr7cVmq/aKAPiL8VN5gpU6z3lPYVMIsNHGAIUflWyU
W57fCG6GC6JYyNVhJ6WfBvTGiJTPOgY6atkIG6iwC1hxv2Py4NNWkwatWg1TGISaeJJX5SeD1o42
mE1OE25YgRumxQvXmzEaANtJ2PAs7wQeQqKtc1unIUmis4pQgrTUdmUdkM/22MPzvxnoVQsiY8yM
aNT0wf60RegpEhU7i+T50nPRibN/Ct14OY8AU1/e/IS5/9v+2kqCPv1KIdppsEnalqd41JTxPyWC
A69TbiQz5uk8RAg8g9P0kYXINFQ9I1frVMFjRO/6fdDCgZ6bVQXakYc53LDDCsczZfWu3K3vgfDL
BrVjedxqKV8b2puxS1ByC3e/fIL8/qIFI3mIUev9lKBorbLYpS/weEXcOIMrO5t7Vfw3CMU/YP/6
UBMRsjXOKpk6rnh5Afl5OnypEhmB1SPbtgjHM4g58VFz9SZrw1ip15yzpjk/SYk1ez13oNszMqCI
/cR901eFa5ooC6l8FbU3WBmcvom8yLlNzmBv5bJAwk51wje3I9Yd2kz8BN+x1Mb4gweDwXhsZEOp
NSVaISy8ZEQbYDojZLjC+dwlgwXKrh7SwV6EsFSUnVr8XmX3D7HGO8qz/MkeoPi/o9ByM1PFf1Sp
yjZP+ZqPB7EFb72JJOzx7qSsoELgaClsCNYmyWdiu+mTkvJPoxSovOQC9oTdLoNc7tyaFfHkiGds
8LrX+yT0ujlRcoJPiJOpi1UWruSBELGPyh6p93G9aB8Jl54OuYF7Bymgk3g5QJvQzCu+TZ1ROwsR
OMwPM5oIVqSIdqmdnqazfAbWtfq46VMNKZ4Pbzlq7n9vAA393hUsm1ruOzy8dL1hpQfPtFApCRp8
vclDRRmAjR5aqiIphZ0j/A7BtnLFN8G4/Hk1Hm4iD/b54QDM6u+kG08AA8e4KazbTVVvFBNmo9zt
yDgCjJSbCgbliqiqP2n7PCpKh9iW5ckZq28uXq1Nasbl5fOBr4sgBAdc5YwyLWOzaNN5GzoBB/ze
5cEBuRYc/KXsv0OuSipgGswv6xJIJT+ghpOoqGT0a9F/DEP5qTxcnvb3KDEI+6p1c7OhTFVOwtBv
Tv5jfQi9AqLAvWchu068vQ4Ts2rapA9gZjP608Wf/d3Kst4NBf3nXgw5tc9n+rw59L8r/8c8JNUz
vcPMXduenn4HHDW7ZhFvuaBLjbBLD7CbDrYUdzMWTZrW5BchXtYqqPYo7DU3Eto97xQn/xxVb72y
yQN87iaGtH78YYDgWn+fYAUPJ0yuF0zGM+B68gkmiCSO3Wc4swshvHblpWtRJaDVzATMniHGKROc
PPoova7vtvaA+7AIUHmZOw+uyeIKqkPCZgFXUu4Zpb26cZBSKtLbQzICOS3tAIgAinveD8qjzgQ9
/HUiZdX3RHXVIlNcQKQfygHG7EpOJ1y6wifznH3m2ZhBM2VXXWZofmfHvx+QDywWBgE/bHwbbOEG
QtCo5lYYODeiCVuSWvEnZX4jzT0vjx6IASLKH/CNdSkf8rcH6LaRqQBkaEd2GP1iWlgIt0XL7qjc
XBS9YDGsFTzMw8AhyebkBtjVeV5pqbQwsxHqvSKw5FRjnmNNxLCZfTFc/whrPaAul7zkpCQM87Za
GhoMo9EKBTjOcNwkH5DcH6SPL1+uTRBxm7zZnNz1cItj+yZpMEkbqYdos0eueYGt7CKRrraBe6eP
kKxS+uLgWlxHn+dDdyEo5NaZ5mCr2ZjJC/4zL+YXDVzAS8CWF4cDBNguIWobPxWsqk7vW0aSRslq
sLcnMTt++XH0+ewpNcxfut8iusbQsE2rKAzsdjZHqsuRlJ2kon0WGDOJI9GC90Be1/bZkcE5JcXf
tiSt7taYKeEoHGfDCj+2UyWV7QNc6FB5qu0t+dQ2dt1LIGZglMh2NAecyo7otHwjL9eh0Keonq/q
mrKkXFPfvXt6TYVYjXA0GB5OHK3lLrT15oplFdFzJffGtNpfYIMYLbfREgmFWQKfsWxKsmtjpQRU
pkgEHGF6hiGJxeff9KvUWyPBkSLMFJvv73m1wHAhHp6NpgYXXbz+ZHK8RvJKJ3Wp2YWbwEjluA3+
tUWqdAXOVL0ghE56l7zb3REC/dNoBkZlmjODBlwbba36m6G7PIkGJ+d/Odf+Osnj7tzOO4axaqee
kzQKWh+lGzkGhL8Bmoeqcg35WC/xY9ssQ4VLhmWc0cifCDU9T+0ilIFoOhLXg56v+oQe+jUlHGHB
ZOWJXgSl9oUhnh6GSOrr5/mCHh4jKKLu5n//lV+Z6Gtu7A/GCirTfACAfhYRU7uMLZ5ns7J2LhFJ
NzPZsc4fsSpRlw7pKf5IOvaJoNBPEj2r+Enltuu4rSbRVa3xW8A8oFwu9OSQBSvErmvu2RPwNZlt
t4EZTLp4+wDZ6l63VNKCswLN+j77jR3tDFtCP54njoIYaohRhnqWND6bYIMs7QbnOfaBEkh4xWzV
3/N01c2QPLBMN/tljc7xeBDrenkyWqkuVS9hIU3zaDeHhprQaHujBpjCkbCXf7xBPS7C9cr//aOR
/8mDQcl4brBXi9UhFHoGWwtUU/iOjr2iVUPIGowGy012bwK7kPWenB1buVo19xVHvYA7ReXwZbCQ
+L6Zqe5Q//2hwNfZMx4qSGW5GnWYoNsKK4y1eyUgV8NQMdE4wG/aKK+p0LESHWdek8NcEzqRkee3
ygSLFuTVTTU4xi1XkkoCQl1o9gZh4yNMf4vitnZE6TZF3gV8hmWri4FmzENeeBMpxAl3kIFfli++
h6U1ivWFluPZtGvGxkRZj6Yw3jS2Q0vuyS4qh9OuChZChi3PDX97T3Y7Ol81BRNwAqqJQ9YZTfZk
DkKZZm/pAugqgzl5f17n6FiC/r03O2PoC8ZUY1H3tiKaOuOpfMpHm6rPjZNb46FrSyQSSe0qZijI
yhCbl/e8WUpDac1avbsUhfK5X7eB0TgtGEvt/kscvpA2B5p9axglz3Z+jW91+sv+AE8l/oU6z3I+
igMJhsj1C7r0k8Z0vG/FmJGtr734yKjthGHjgMj8UILSGLTiIJrqQbfbpUVkQxIS9dz0YEn98c6e
bZvpCnuCVMQI4DmjVhw13jhKcSaATFoDGnRiZzzhgzlHK5DRrQg6obJIX5ykyHQOCjjNR8NEGu+c
WKyA3gqHio15t1SFF+GTFWsUUpvAZKoQM1R1EkyLmFrTArkFMD/BrM8Hj8DjHwnq6SDuh+PjAvXx
s/k1QPUwG5GVu5YRHVKnk/2BT+pP0SGNu/fvam6bN54xCcbEUvC3Ds0DRAre/xR5TXwsu9ZTqcpI
1czbsQRzCUoODN1q5r/LJ5p2UTdi5Wc94uT10qWSmPwV/MHE0PCdE9apjspby7o/HYF+buW7InoK
7ulTeU2WNPag7FO+lcCe29TQkt0NmBc5wyd6fT9x1VH6liRb/KHViKsdBi9CTUo7xTZBbi9GB/OM
g+BFCU98XrYFFOXKg4+uZuQHUXZPs6ZLqBb0/yAtZftMKtM5A1rT98bZxqtgs2OysVEu7zHTfjEW
TEECXcLf49az+oxs6J6Caj7pZdFMSCDLkpqFFC4aGxwN/vPraKhbJ3uuqedbvyxAoRpG1tuNqjyM
kteHXP8yr7rB2baNWOXQuizSSMWVqiTSEff8ZUgGCtiKqTRDtQEwZkYbYnho5JWXuedWA172Kiwd
DN7KSROmMfov6Dh6+REBZMv5EEEQvgj9rqeBCrTkvail2IkGG7hnsg6v3H+Y211DyTIrUlye/kKo
jbxM0gJMB0QN2z6Y5HKGFkzaMceGrD5wcOkfJnPbBODtvbmWDTIcLfyZHUpnva9ssYEysFFFVjnd
glOHgQsrYg0sDto5ojomtN0oKPtZNCe6ULz3nhrBOv/NFj+eSrxSxhi/KlGMs3/5/g1Yrb8fNAiy
Jt9ktC/Re7vrgNpa0zvVGuO03owrq+fahFJpiJ4t2R6C1wP4+4FbAthAlOXpwCQ+zTXWrihdKpAV
PAImWQLgbXvT6pRa2BC9vIfUjTbICQWOxeCpc1czCT3uLxAo4jO97KPqWwC/P+CPwyswPZrQJ8l/
wQ7bBvxif4IEo8ttEpNAKxRPqfSMRWserPLx22xyY+8y0pK/flg6KIXixyxQctn4NPIrC/dsIdJo
iTpG1R65f4W8AqUX2L1WOoI9d8RYzAJXcdfD4ciyts3EbVl3FzjvTHMLi/7kJVyRYmVyD6RCWohQ
d1RhoHxzIq7Tz1Ay+Tp8y1PBwqKIuu9hLwhONULzqWZENLHstq8gfbamQR8wGlEto5pVYyHOKsZy
ogLIsKkxS+S6J/j30dIZBn92Cs1XaxEtVWCLlEPlyUdaea+Ptp14L/4uYgJ8yNXydrKRM1zbI4AG
8uY5dFBNEkeFVWG5g011YAqz2mhnLAlMr524cH6cPT3P4yg2HEWD7+Xkd8nSrdi6FdkOXFXMJdic
90nqXA3qTXyFbaLM/OlTPHyCEBhWjUAJ1qaOH0hSeD6BaEJ5nhV5bsLiD1lYDfjEfkMT8tmtPJ3I
vqyJGNBXwOmAbMzAH2D93aRZyLbaQ8XVXch1Z7EkBaLtRgGNf2xT4atvy3gYAruoCVBTAsC1Nam2
8+UNNH3XBFuAZXLvsDii6QKNV7v6T5PI/l6a9CjAPw+ptsaM1YqfWTSQ+lSX74TUuxMwsjX6wRWn
/N/abja9b1b0XB3U+bnLZy083Z5za8WMLcBk2eXInJxaC6iLLFQsMExtsCnCu3igc0IPQrVNjXxN
NuxIhaB57gAInBihf3RV55IbvYY2K7JkRdtiexAENsD2pTGKQDI9i11O5NaLQharRJcJlyMfJqSV
VgP/O1u1ec0HWDyiP3VWyMZDxGOgr7C0nd3xd0q+uMqv2tsvlsmcyGdTsDUe149AduO0IxDk5HgO
U4esRpvDw9T6wDgrRMdAZXCzONezqi22H1GlIVduC3vlW8fGSciMye1/MmyKRfReybYch2zNre4x
97FEJ2Foo1d9X2avjl5K0TZ/vvZtbrB9IYj3PlH3EuFTruTyjW2M6BANL6h0MXsw+rEAik9uTy62
nSQwKk5iID5gfy421lifgQr3L+8jOOfSs0wovsXX4NwbFg835D+geuq0mTPI4GFyoJHLuTcc6IqX
F8uu8S9GLQheKM/CmwZ3M3/WXraene039YNLTf6LxLzxrKd9Jio58yJunwCy/8oc6WJbzWhALUqs
uVMpWXcOfITabP+ernAm77A98pDS7EuRenumQ+3H6sYBkUh9ZLxwH1as8QFWYwnhZAJ3cLmL4qhM
drFYS3PWvzIne05OyZ3WlbQgnimCgHmT/H4/mLlBPlPJb2ERTjsOJhnysfmMdG3k3oJAN98Fgexv
FOnU85S/0yEPHq5ru4QRxr4KvNHbCUdTTeVP6GZXyv3mKQY/GGMJAV8CkNP7wMfKQwEDagdWWCQr
zfgp+2iN0YDidDwtUVp91e4YQQfYhCqRoEywHxW/SDHvXfrCmzxatBZUZhenxqgdXkWWXWTjyKOh
9e8syQBNqt85iU1qGP2Lgg3NOZhMuHCeQvkA2MiFREfwaMLvb4mVi63CHO+hqKhHRZyEmw119rKY
JTy/3ewgNY4GKMyEt/reSSIOWcAO92jVxEd31YQuumMGgjGagUCR2le8YT1m3dQqkJ8FmwBAeSO+
ElhbSurpcNtt0rz8z9aovrCdu7e7Ly2hm1EXCdW8+zUPzzIXqDFA1bF5pVapPFHuGnYBuB4Fwrgu
McxGB4DhvvL3BPBsxfJrrKEO0giLGbV3fQxbPJrmVhmxSG7j2qARByI5gEyS1p0diQbC/gNcu315
MSayKGRNjgtiuF/xkawsiN9Tmux98fV2HkAo4HYDl+hyhuUaQgFrdt8IfWSbq3FddKGS+slvHWDQ
9ThnJOoRFdiejh9eyqlpilwF2kdpU6L879fSSim40aQ11dPFq5Gn9GOU9kLmINg55SGpyPoENRRQ
R10dxFfDqpBzaHTgrbJ6lEx8mC8FJtO40EtkOBpXSiZN/43TJ39nwUTmyCynoSRHCJrEdbluTYCr
0b+24k6ifAcf8uSMftzXn8jh3JqlXhE8Gp5DWDjja+2TCQdxPmWdTT0BpzFGTqo6LpsBdh2eczir
d3dInan+nBz/OgKLdDuj9gak3Eg01M7K29MvpsQwH+aqd/qw7x0uGsYvYCn0WYdRtAdXcrRDDwSU
qafV1/g2iDtZsgULAgGrZ6CJgWd+FYMIaiukuPm0O9dJPUG5D4VVg4mfBkQNEjiixDf9Cfdoc9Mv
djZbV9MVLjrfSoh3jjoy8PbCxh4sKx0aHVMIjx9BHmw73LqX+mlOg92r13Z/1LeeGuCxcRfRX95L
Oa6/+G7t8hVUM7Nv+I8jIb2tkxchL0f+bqNDzzHtnZkoI8r9J1P13HW5ocG1QfEIwxrcX1ucCuh3
0MqpsmeJdKJ6LNQtZToijPm+AcM9Fm3cZPfUYNmwriDfjA6BW3EnG7oeP/sjrTsFG1csX6g2Fw9A
JzxKg+naq5Criq4X2vmgnG4vIn3RlbZcSYXsHesAYtNYZfU8U7TvOkscltHlTCWOmTnVxowtmbsa
6/Be0rpnu+Qvx9yxNaVahsoPlc0iU06CBDsWh73nU2fejRAT3tiINpJ7GUlFTm7Up7RTa0g/xfm3
uYCkBbu/Y9svWg41EqhbJb2ImpMxHoFksr7MqcmQfnKl0TSRFdL3duakHvYfDAJM0ZgooYAHTpm/
FRQgzhYkDZU5MMwqYYI9ZzdyMg6/WbbvbN9vIlGz0S9asvjp4uedYxT2PtqzeN1qp8uB/MqAVSl2
lnHzssDBgv+23jrunzXSjSQYKQ6X1mKy4Vi4NBXcbYo0NQYTyttX/j1lHOj6NMd0vGM6Tn8NWI/K
RqLOd+VBrJMrqzqLYdoGkZ5CUH78OELyvLkSSwwgFh39dcrsg3quQccfyCiG6pZld9BXD/MAU509
Fi7FAyne4gOAC1cIgK2eGRcF8yrfiPwDuYQvyHyeoSGzMs2ZZy/t3/2bT/YgBLPpwiyVuBh19oxK
vUDiJvED+rUgxQVJqYPC315UJSgmohvlqVrTy4JbOy/xhV5aJVg9JklewA0XY0gwKLgH6cRerkRa
f6yBJnTLSDFqXaVxZwD1BAraKxTmhsstU5o56sloAmcQLqFyyCaQkaUuCL8Xz6bNL579UObqnpCX
f5uA6UQr25sZg26DS77HI0idzOu1FapflvHVIQg5zaYzgjbxxGwHgGQ4Bnm71bGm1MxCb9Es2ZGQ
j3awMnc4vHjVPCBLHhaGLXM7AYoRnpZZiKMovTCghTI/c4sWj5DemDFYlS00A2kKVpwF8fmbaZld
IuRVueINGHsOrqLFne1jCCABiwyvqALkUmbHsQbehTNFdB/is5iylsQExg3EgsOoh6qF/CbLVLBK
1MeVkZIQbbEc7JEzlXSsKVayTCyH4reVK4TpvfE/v5IouVdV017gKC7FcXKX/BhSIn8OFKi5tqZ/
0jIiB5gNiFV0a4cVjuStz0WzzZN9SobWL6kI8l/MCixBTCvdH2YLNO6sEF8HcCGF3Ce3079lreoW
1MCy+3uyvVvO1jCCX+3RF9DeNf4z86lxQmwgXFxdF8c6RtudaeQxFtKzMhLMqwJnLMvWnlzfvamZ
jvKY09f+A1RFLDxdzv4MsULwRXRy/0nQFC1vydXc4zIA5lGafAOhwHxvgqHY1SxSKI6IJ/XHmwaC
iDrwp9O4FOefpYFhTIdBgOHqdHUH3aDSEY9JuC0N3TpATamuqxnlpWciyBEDip7fQ6fX0IuMiaZv
qbQL8V4i4MgyJjuVOB9d1e5S195vA8D2yiqEgADHk3Ly231T0EaV/GCMXWBFyL3l03NLSfvObliF
vQ7ILXn4TJFwZ3CBSFI4uHVTpqoiHCu8ifDLZyrt1DiReL99WkP1PpG5Al7Tm0/Lb30vda/4joKC
qURFLg50eQVaxvDxcjNEJyUC0QGv6a21+P0wfdKj6Hp8H7UhyBjPLvLd1wDZexlQIh3Y2HF/012p
SYY48fmQ+c0XJrFJTeNH+mqOuxYBbdkwR9CpwnHPE5Cslm1NkzTiHGoqGLUhRdd5OspE1aPWHhAp
yVb1tlNMpCBymvf5zfsx6Kt7Oe+s8/wMAqevf7Zr24Li0Fp9KkO5A/69NLv64UTLs72SVMABEaLQ
SGCK8ELoYYL59GaR16TjLJ3JiWiWavw9FSpbb3osrav9VAZcjIhDIcsRZJg0GO2XBaglHeiudwTL
lMElVHVaJhiVDL9jP69g1GP0FK/OOwTr471WEMRJ4+Vb+45XbPteAQWMts/yvDf3GT7pyZ5iY6+Q
U/erYr+N21BhnwbxWbANAE0imkExZ6eeSrODB6Yzqli+dEmFNjOxx3V8R+Lt0awx5MvpEO5fBJNf
u9kJmKjsIRAmv1pdZK08gSGBBtfC69ox/X/BBQkWOt9LB7M7Rrgpv2guEs/5Lq/xzR4es99bR/Op
a7Yb/1SHXzMNEnxXKncsyc31q5+NOWVq2Da9yOXQjluIcI87v/8NPIkSHS+ZDbR5la6nB7wcObdS
I1dcAZYaWOMvohWArIWGTAKprNxiKhsma3rGPsdyB4klL8qJUZ1aB0yXO28XfsNbUlVN4RrHUxJD
hZTCbEr2anb3EZveMyPwCTWZ+xNpSuCoh2gYjeL3B7FC4OwJxvKLti+cwCCTvdacAm457KchienF
9nKHrsipU3Q6IzK4fNerOjst5F380LP9FRPxrs5F93anWA4D7cjOL7/uwqAeRPqOPOLH464kT+7u
yvlKO8VBSUCTzID++fNk9kZorYuCXAmk8Lrr6ZERqt4ACLfOztZpD1yBS/isLUOntT8RKSxkpX7q
EqD3ks2YB62lsm3ZyCAzmYV4zkopTJCJT8XoHAX8LK5IxStl84PcL0QR/nQbiQCcCISvxFWaETgi
mfgQ73DUj3dnIKYQdYfyycK+z0HXm7mQLYOqKa9E0D21mQD1GIe3KbfY7wKdlxBDJYx6ezv0Tfor
ohGwINDZzXYQCI26bTJQUmVV2DGOmO0ZKvmK1t82ZyECibxz/GKhxDQBbCPYMqSCwbB/bAPoYg0P
wLMgYcsYTu5wtWPDbk6m98XaCNxUhBmv84TrFtDh4DAcGvB+M3ZeQNm+UX1Dw3wBiCpmOsJyYF+V
mctZcte6UghpmJaWktKCFC0H8N7D19igfEuR/eCxXbH458lhVc6S3kUvSfC+gklYVP9km/Ou/aBI
u6xBcNk54kNLbjw+J1QakF1TrLKyisCKmEXnNoyUbctfWv+63lx91S0TeOrerk1DZoHqPYHG8c9q
ZFvWGEi7LQsgS1zHJwoGYPhru+cz6OBl+Tca8EPF21vLJK6i196+p6qaELK0U596dffMEDTyLxr+
MEpCZdvb2zjBRyrQ9yn+Q5tcWgl0v4SEbc61DAVfmHhZVR6c7uyPXDrcmH23pr26NtaLx2Pa+GUg
BSHj+Nel2w/aIDrDKzmflMLjcFkz4zsXONWhk0k56V9rAX6IHAYCrBO+1GoTJLK6MUeKBOdhkk/d
0+M74ktHjtyy8k1v4Ntx37FMXCeXNpTvm03UFaw6BlOO0bd+on8TwhhFN62Jo6nCxAesGYBn+BLk
iCTvXSYLiNdL0TsD+H27BuUH4ixJqWWcPMz2ZPHO9MMlS33kC2IbTdZw1psBtpkTdCWdK0/cr2PF
zh6iaz2NyzrHsZAdkT4gjwVAt5A47TP8ro2jgPga6J+fO1w10+O/yKWz1zUiTxEDn/RiSN4mgGus
nMZPz6lxcU5+yW9fz4A8Yrb8T6yDHzzrZC4tsGSOsxh2VakeOmQmUJlro/m2FB+YRp2p7Le6ZdG0
t4Njd8PvdvgkvCLiUDJKo9FUEQTg/tmraNkfI3BSWZgw+UbKv6AzvparHsXbNkJTbCAa+SYVNPdt
4NpC5M75/IAQk/IzX0Ixd4v73YRh0qEnMiTB3B24e6WhQmAbi02KTNYriXc05jD7we/GEhVI/5og
ibAZ8CupDSkqUeou1V/bqn23YcRvziWeHkJf2X1nWbyYu7nOFU2T1QYb719ahiQxD+nyzjRmrIf2
mMXNaQ/agATforoQwMXwps/6LukzVtx4g9aXIqu9EMQhxEgpmM2ch0o3ayRZW/PKM1kJFpByh8Ab
SAfm8sX5VG7IYxYg+8fOGL/PLC8QHTpr+M6EyKNhVUaNB4kcbDGBR5fIup1cOyIlYLIZyLWSzx2f
t4Bhn1UbkoQgmGwb25kIQIN+x1Y6RLq3zGa6fndsLBkKgv3xUtFsXZ6uKhyQkecckbuqGrQZaKGe
JMAhR8vRrXvifFml07LLuTeEUiibalGHvpUG+yYJuVSPTPoQYN8XG9HDsN5OH1YguBau6GWj1UIZ
1SKMS9u0Kejfc3eoD022G00lQvbxD5t4rIJPjarybmvBypvPfAqnqfrd16Zf5TiMFgoxOso5xAzU
FtCFGweY0aS5h+iRzzT6RuKC2eQHBiSQPGISa6h9X+j9d/GxgGTHkmFivLi9xy31gA1MUNFBVohO
RENNg3EFjEgI3b5FKalOi7KUVIOohxeq/W3msNW1KDdPHRFjy1MPIgUwueZ6M7956qN03hU36eJ6
hh3T3xUQQfmi2vKrxZxKpNlijBpDsWRS7dxUazLmSyEzFthfPg4zjfLda6ydO5T3jFXPbIyersI5
l/AQowsa99tpNETL9sUtgj5NiSrSQD2SCuaa2kbeiLeu6noRAbvsQDmlhxqWzgaxVCoadJH2h2v7
dXIFuVDJjsOdAkUyBBcdCxmu94SDfWO/bV+Wr6gMGIcXS9YcpU0KR/gi5cDxfxolDN9q85YEiExB
O2woIyUSsIs1WdmGU0UtXiJjjJxwzP9Tgurw68HgQzDhNLBO0CdAcGoZmE1BsQFIhcAEX3yPRf30
tdlPBs3CaE826eIRLKA1J32ONvo8sgEQVAKau2z5yTzGsewTe466q12semGaqHKE/imvzYcrUEUg
uulhGdU8dUr9Ij8kEmTFmgeP0tbr+5++tNmfi1luWhEwkLc0iGglEd6iLI701HbwybWtdzmYjeGR
LUSiiL23c3NGiAMkU4zEUHLk44KLt0uNuwcRErgFOZ8Q7LSLhtntzvFquSaNCDkkebmzYq4yN8GI
DobRO7W2wWfGZG4KX/TE9kXyqQCcassyxq0wbTAGH522PqsNSgF6Dt28hG4lMmGisu5pRFWTjFae
F4B0TA8NSkyPqLjD51qcpb6pZ59CjsAx8zqhFGUDD5uc0el5rw2LEAQE2WVE/a3cHN97aAAQ8XS/
sKIxPMjm/NjsaRCpStZYHqvEjwwlsDdJL4BYWXWeSRVFOFwa3/m//Y7JL8vTCsBbrN7PITB4frHZ
R3aNkB7ztN2ZGQAFUHHWLqzKoDAdSqt2495smgrMSrfewrKME5QL+ytf5T2YwjSTmkf7LW96EOpY
rMP+N8J6mnulbX9BFOeU2rVlKLAIPP1oXD4oanD63GPL11dJhlXoOMDlUkOjhn1Zkd4dCQiOSrtT
aWHs1awa8OpN89yL5fmX2rP+yzPOsk0eiFTkNKYnScUdPDR4GirKRXl8FqHrdAAHryEH71464vpp
tjPhNfwpu0e1vxML8NIlP3eBwtJU1RQWk3fxD85mP1nosm04NR1LQAVJnh08cLSjvu1WHBaVTIHB
eZC3wE/MHj3kpxNeTpRhTGotZ+1VJnZ9ogbxWYn54DkWzNCWcyM4qHGiWZnscurxAfLEe1ww2oZG
AhmzEXcqa1GPtwmCVcAJhmmRNVgYcpgeA0VdsD4xQwL8TRf/SnxAM4nGhrqOiocGmHUXlGhMT/IM
V36xxeZvWLlIBbF/H1nFJNA3rlkThDEg7uuOw/Jkpvv+mJnPRU5D2HWs/FhSAVJU0k63weNjMbi/
2C+WFFXWBOkAAQQeAS/2Vez3r+DI1qWqMbQWekyIGYv8CVg5PsnBiU3y/8YNK+4S6PvOIDTS0/vd
5d8i8/ueVF63dqjFj3vyBnXaZUvC3krqiPvr7pyvsahskSjQmRfirWz2+QS07YzAEm8Yug4h6mn0
FXUg98uQyBCPbKHxcFsRD3g6gdGUUW+i2RD9c7Ib4EgjXgyrrNKLeCFtmNCS8/ESG01S1b0Q4PVg
L2kI60mSialSNMwNx6aORn8AIwBeIaU3y4ZROutfB/B0UBrg0YWE86IpixaNr9iZA3axxvf2+tEC
Sar5nRBzM6NkdE69463+6SPItu9yAInkRduE0nGwMGrEWgSUvvQf7HyRWoIJTBBHcWRm2QoeXzU1
Vgc5E8qri9Q3tiUN2GOHmHNIaTzTizt52yrR0G1H77a7XfqZgBtQhqyebRWF2piP99LdRYXwRfrg
icjvnlmiJBNOcpM4sBpCu3sf630pXOrOJCuKZxPHwD6NA+4hM25ed7oOvH5kuOLkgoIPyzGcvpb6
WtY2ozdm0S/AVxAhJYYGurXteuYl44NHtuDK++df+UIAwHCx1RLlHI20YzN+QvH3FbPHmNkK0naM
CQgmaUEtcyNcaKg/YKAXOtNv8rXmAvqUwVSL+P27U4HyKAcEF33GVL1wOASIE9vXhFfNYKWZC4sQ
1k3JLI1lx1O3/sIT8vgYQonjEesjHuTXcEvF4eWKGIPud2ZV62mIDzO+QyKTse7rqZ5+DqApwgYB
PgIU0+3Cu3m1SsYxqcQdw5Gttfjy6Dn+pfXPCHRF+7D2K5bzk1PM0o7lPMDy3ykHvIwZFampfQZ3
rGBg6PXzv4qGchOLevRyvNgQhud0juNw/J1UY2je5eq6n1QJ73+njo6onjbHuxM7vYeft7yAVsEc
2toS1N9hrTpQ1WJv9sOsObUAQ00QIsyyyx5BVGKAzy6h+Q3tWP5DT8AGyHabfAH0jROGEudLX9xR
r35EbH98Rf5gW77aS9GYIEs6MYkkPWi3fwYHaYcSMQn/CwVXp8/0rmGcqt68d+3niVG0Szzy+T4k
1n/c1BFsSFpxi+FvhF/QFQ97ZXjD3q7GupxBKEufsgasLDsyZYqGwNCZdNdoBZkLlazfhwBDpAJ/
T4jlwBAu+8/Q+6RpzOAbpPkFDgOpnuK7Iz9vDllDsT8jc6WMs8q2kYC2xrgtxlbgo3ATU5iQ1UHu
N5CE5ECej6lKaPkroDv1mqL9YSkjOLmKvPlsa7B1g6VtvvoTB7lhsKcCNHNxuugQF/+GMvw+TALC
4HB4/qC6Bm+cAGtY0AQwMWIXdbuBPpwNhC+88oWkdpHgp9AIyVsRUmOCViRI3DKDgDQsiTnkwG/2
TGSlipYu98+d/iQCbFBSUHAI+LVxSDMRPoajqbUdaUnvxin66C6g4V0g+IFiWPGd+q/DtGlM0bCS
ezHzui7B36ahUKF4t+N6iVQmB4il0rIjzj7371av3D5lBJkbLAK5y4eadltF96x2/yMNrx02HcX3
rM/ckAehKGyqu0NyMYlPa50KVp7WX3r3QUK80n1yt+Iw4ih5eQMKBd1RYgMfgNkWF76HwFRcqeSC
p8FvQbqV+aJov1e4/0YrS07LMsixAHDZVqk5Xj/PIQSC9dDlmJNSFNy8SJKpi0QNmW/mtOSYFFzG
LeeZbtS80dDuIweeFe5uvGLtCyXiApIHKR0uV770aN6MbrNDi1IwhRjFDs8tzgRTlwIMkbfw5Z8H
UzOuNeceuF4ERNmu5DX0i7ceoHoqGslAzlF0yxYsf9tluze+VLfE4NHQt53T09XTQoCg/UfqxmjV
qTSiRjA1CNGLqH7w0I9weGkrtVbvs+XA5iaKfsdi3eEjYe43W1taZL+q504P1EDSYSHu2P6QlZeF
DCK3m7Pc0edoN0nDczUAloiSZc/G+syod+3+uNWiALeGGaqc3XeKU1yE5pQl/jTSKK7lzxKUHewT
7x/IX45BKc0naiEYjWBhMfQ1SYPx6il3r18iJhOHe2g46shgO1n+eiQHU+WME8Lw2JUXlsaFg3pP
zDs/PLuxZZ+tNh/Ra+7DOz1kPwRrbxdSS6M78DWgq5zMTym7ahjpwfqdtCLrXvC9F6zGeHvRGxrb
k90wMln4BaxNoJLlmNecsBam15Lz3LTKKqqkowTZvufSbn+hqTur3syVLXj/6x4Qj2DyxR++pdDT
Xb/+SBXuUe0VP31QB4LiBokoBMqeLzDF4barwWtBucc/QnIDB/yPq6idpDlAAR5YpFypZM0zWTxE
726cxFtLiUhmkGHqbGuVAe/BmBXLLViT2ptly0beDbkqk1nDs5w1AELCLIk6y5cPh0qSI5GvtyG5
YdS87KDYHac8XDTCe3K4Jm45RnxAytiYE5weU59UzbzEQx/8O+mhUo5/15KgvAgCWAz6oetY3W8U
1HeG9QAReazCkzpq+9CPmr+5matpSVMJlg9ZnwWA+0x0rewL4UqkdmFUjzJ4/k4GaYX8GkQs6PrG
3vLtMJwGHWLCNxmimjArqZkuFUGxEP8YTkTylPlLKPprv+qpaQbEuz5D90tVA+vRRZspWE05L7Kq
gUbT71O65wa7gpy4WRrL8Da/o5UnrhcP0IediMdsSjT6Fijo41FrgOPYiIh6qnNuxpKzlBZ67+oW
fan8t75lqLdOxZnn5rCaR6eC6DvLEAzPFPv5BBtw0F2BBH1n6+EzoQ7Wtpw5SZrK7s8YB8XxEt97
khReBeb6GaLcrmIbXrcR5LxXPWgsrfLAUgUF/3wRssI6sk+5pQ9xm0LZqA8jlDhZt4DqO+oyBn8M
loKn4U9sUXZSBN12EDyUorl8YkMThh14YLVaP9sDAvFhYh+7ES7IjrGmnmFXvulkxMN3uWoW72Pn
ms/O5BEpsHiQMdk/vlUFhGh5yQqp2YChPSUOlvV1rfHZE83PTLho35OmVJXHXS4Bbb/FP6CnxR1o
zCwwL1KM1r/P2DJwCbO82GlCk/V3wPbogADRDpKkQ5+M0U2GPZVcYR8rCX9ZfDXJEgHnyhIcZztq
YmCZXAkbphaQm3AdzByaDgRdQG7L9z4Ijw4wSg3U5pXHaqetDdAsgrXmV0LIYk4wjhxgFS6uvfR6
OpbcGyQjnBN3CwLmZNd0Z+cTWk4/44dANdQkbHMUfu1cD98UMMQz+r4R+4ssOSGVKfWKMEZiB6w9
w8WOGlMSs6ccDotsHpuaoC/Nog4NqO48C9iwm3z8rLgcOnv25FLalqVMpNyHKage+OH0hZ5kXt7Z
f2gwC0yNqwWQnAHmEj/oWyzGQCwKvqbiYTq1TlE4sakXJKlW1eNaBLpv9+m7ifj9kvOWZV80aqPZ
xoAUW6VTtw6RcCPBqR2aH8s25qZBEdSQ0CPdnS0HkmD/WyYawyYHaJLQ89p0o76xlDARHcX1YqcJ
nUIbzNcrctHHK/EsKn8SizJRAxpE6ev+eheTylDRqQTEykO9z813UWAfXUWjQgAmhoKLb5Wor01t
c1cowgDoEXbeLe3NhV6W9WZIhT+x+XyIxnLBVx0fikXnj5UMqueOTSBFjQSdsnOIUSVWOm99Mzv2
rlH0WNvR7F8VlKIglqyzMpqGUAgn7DOg8RzxUKhUINr+CYH+Zt/ggybCA7se+60J1NU/kBQZw2XX
CWKPVeHjNeqgsVv/5YCzUira61raBJQSR/5du+EHNpTYNY1ryr/eTshMU8FFfP/E60yq/stN+MvZ
MKXzaGoIIBKUliEO/hkc7bHAEBmXsMsE59wAUi+Ys6fnA3kljHk5HBRRo55jK2zbwZe3vdf49CAO
iqbFjhf008j1cSee1WsI5sLZFhLuDpf6X+r5VwCaxX1eJZ4/rksa1KJHEq9r2RA9V87mKR4yA5L9
1oYSwCFWxv9jIw1nj+BZsIBnA6Qmu560fUnDmxRsrdmwQjZLOkJg4K86NA52e413CDjARGYK+aIe
+MRlHkL1PbaS7DrtK0KmyXnfIrCP/qHmqpUEe/T7eXNqTTTTZcPinNVuLUY9l+2hG/8m8PUqKk2T
HNaodYMBaQdXJxNTbDNjPqC2HkOp51jirlOrww0hE57n+pRgRXuRSBQPyRc1AsXhjjr1/FQxdmDv
X292I3FDoRHmlCbrDjyIiO4X0eaKhsSVX0JSG4YW+ZQ2tKtTKVe+OTUVDPB0MtEDcLXqRXqzjpY1
haG9WKGbkgbDljy8/2xTJ4PseGv7A57e+bRyTNVdw8gXK6yXl7ZDbQEV4PEW2h9XTBzXzmuD4teY
RW0QvxdrIolMrz1/lCkisYJ/aZoHnwxZhyXi8NAPdhnusJmRJ3lWNtz//aBkvZ9zjz9VYfkhmaGU
oZZXe4nOZBYlhqEw3j2Kd6HpKSAf81vqghmQ40jI4eztHprrfgqohW7Wew3c04cRxifZadaNaWDI
iqsbhwDCDDIuo8GY3NpPy+MgN5QGHWUVUgt5bcyh9a8Ah66Fv0fUsQC5lGqew4phI/XSjDKVHFx3
klsEjB2fXoLwp6T7uCMZGyIy8tHZLZfnXoR88dw+Gg+6lLtdHvn3e3TAG9VZtbmkmjOIHVT3h+Qk
pGaLaslCDKR4EN9XNp/BVSI1UY9bCJkZIjrEzQijE7upICg7x8SEXh7vyt9MkR8CjOcVQgPoExdy
NAYVTQkErcYJSjF2R5qHMivIUafAUdS2xEQGga3W8ui4YneADMoB1KVVxoJ8J6bh0odDwwsMNDNU
jqK2zIQwgrwvtoVzk9ID7af4P3wUbDeQBNQq0yCgS5fONf8gDKxUcdvKK4/JULjUIoR+aAmahRpH
kMkP64g5pffBxlmpL5nm+Spbj1NnSI9X3Z8J7uxXoFtefBhSzmG4ny/jolynHf0/+mtJvekIqFjz
Fw0VW7Cyo9FsgVLl46MpebzIucWjkYp1j7NUtxDgLkSNYFV0K81yAQHittJxIpKGjhlFPuZkRtiB
30qf52FVip7JnmCUhHCt1fWoYfcWmTTFjjvF2P9VZMOgBp5W0qamGUdGKJjWrdRPBDf+Y8h6YXa5
aHWHsEn4XealBlcFAazNW5IcTdUdZEzLom10yiuw+z9kzrmU5QcTAFOfdEUiRk1o+3zi/X4TE2YU
vZfbgiHCkknnKTHuE6VoTnyFoguLnBoXkJxhY8BZYdGW/ORsNkb1qF8b4S2PHgt3dAV1S3P8RlBb
ncM+MeH859vMhmdIdneit8aeBwnVm679/nPTW7qsqvBjiCVBSaq34POHH1Rpssk6DtJoyVmBn1Mq
E2vcK6+2hO8KbTOaB4hh2vosY2N151SSpNt6AoVtD29lNVFmgPTVS9lhxfsLtFMjrH2KZingO6vF
lnI8163ynDKCSIFiq+XHMqq6vzQY5QhoG75rm9eGrXsUy2hf/QykGjY1nS3idZDg3YP81LK0Jv5H
4hsl57sipYPcXJo2QH6PmgzXnKX3t60dhedHLz9yuBAcfUPw/K+YiZCXskVA8PQTRRx9GiiDJbV5
pvN4rMnVAxQ4SOiH6GrapfyTRpdy25BISMH3c3HW00dCinGbHJ/fIEafKTg9+UFEPVByTcXUF08e
OoVUhNpIRyRynTSILF6UP91xEvHsJsLAf2g5aI2oVBdQUv1GFWPAUyvXuZ4XJ8Kt9S0Czak5aFKx
f/hKtHYC7VJFlQ1KWIKRsj2W9oq62dzMUidDbcBqnNdjWud3ftU0n+8qLtYfMppJfszeo1ocbGQQ
Nkudgp9ngIVjx6GCk7GEfQk99JmUVMh9Vf4NmPvhXOVkEkZIwVBC8RrQIWkpEwPAwNHR92msUApZ
dA5V6D/KE3z0E6Y3K3f+NaT+nq/+DehNeeYbXpoXaGVL4GA1jIOmX/Au+D+fmFM2q3JRbEt6nLdR
41OrC9ufqAC2rPw6T7koY2f6i6rSnDfY22iGAv5cBRWvpMzJ2ORtVaMygqgfwuQAohq8s5Q+OS5I
NA7A+265OJF2wb/be9Y1PtJJLo31XYOdLQUovVvlnkyXoyAOqABXzCATXNgHESO3b/b0ygk5XO3D
n3u+IQtKT/8ZNFIlmkzfOtdtEz9pgLlxjQYGSKqR3d0CH7U8yMSMzXl8r1/p+F0s4MM/7oqlPeWn
O4iRTeA6+bzTO0ULnqRGpcwFOC2va+Z42PlZaWf1oKrzgeCJMl752EfF82CN0dxOYNc4DOjZjbVB
ovP59HwFMfIF38lymQltUMLnjnfNNBPcq7DU0HQAQijxFq+g9ipPw/bt/ui04oRBrCxMr/NwDrv6
+F15WpsQYpFX2tneX8cRBFLeNF3xePOSgUVr5glWDN+2jPdJOPhd5vMP/Ogch8obHdovXPsWbv0o
JjREYoJgbNjYRxeQz9Bc9vI5Q4xBP5k3ULjA4SBZ+OOAZtilKoI3tNCZLhaVjWHfzhP/cuym72PS
FQlBsp7V9ZbPecI8YPfViurjBnDKvmOvK0ms8P8tHw3DQTF7MduqZS65kthLzNMXPMaJNS50NwAg
Kmxkzi43G/HDA6Nr20UO1N+MtoA4sY7VdSPQowd8DjjtyZ6GSV/3XWnDGgDBpEvsOsOI41NlEBCX
Mz4YtxJkgmIvR0sNptx101Zr5+uLJDD/pb97vs2S8YGd4WHoN3vdJuHo0S4VjT1boUSzJlMh4o71
JmUyN16yqgRRF3Eww4fBHPLr9ZszdNtZYOoeWvL8JY3rak6RDv8PV48fSq5w87EZ+uOlskXII+7S
UXW4HXC0tb6xFCUPr17y3sLQ3CvOYN15y5SqDa+9/lhlm851f+2Oqy/s74c+7uhu8v4tDyMXCZ8P
rxSRugb7ErzAHO3pV9bgu8sr495QpeSdye2tzVpVLK/y7rcjEslsHP22rE0q1QJpUVKUHz8V53FF
WwXcGdGCd3y8a3ZSnnlch7x3TFnMeOCI3DgVxrgo02Os39kB1J1X7BpZPS+Qjwd2dLoWeKvP5lhE
xtdIKqYi7WbrjeINlafvNKB/VbeJimU0WgxZ0nwn+94c/eIyTVBcr9tJFZmoJf/0i5Lxt9zdrNv1
rB3vQhthvnxsI0M/AU8z4b9KtvaEmBglQCkY2YFQrBK8qZqUiQJzptd8hDWW7SKEeiBFlFqLGZzv
V5wUuswOVAnnVTRBhATS8QJSSvDNhivTZEQ1RhVxkI6RnAX7sFV8GNKoDyttppCsKSu6FkH7lDpK
LlptSVzMMXy3mBQqcRdxRoJxlN6DPMNe3p3Y35tyregBd4ZQSoOYP6skebIJtM/dbp3CUAQ7zudV
4xx+krRmLWJiEpuRqfQ+g8f18PYLL1hE80P4C5I5GmvwRimSH/9dfWUYpEMSiKFpNtkvw55nRw/4
YP8xGJ1LMf2ie89vq6G0yHFf30KM7/v9DbZGO4BffLjktQHeGnimWJ/LWWKR3cuIhPOvsX764wc1
Huy4CLsgnuwVkooijXPGxZVq3sLscAAXxixFdc2B34VpPa3tYYGIVx+hx9C7WBtnUc9qqvgXay85
36KKS0Rk7E3JSxBQlr04dJmZUYSFmLsj4xC0ZLwLl7ddsQFYwfuphr6U9UyYBLBAOG5DsViKyNzI
0HMcFbg1DdM3/N8+l2QnqxoOrHL32+QU/docfgLBk2h3qGZ+im4ZBBq1BGMQVU35knWt9T6DHz0r
cNW16VokaEXxjbk6Jk2ikoxTIuHjxULg0H4lXpEfdxmPAZv7HTxk6Acn/KGzZLk1aPK39Jjbw1BB
KRE5DtvuPMBL6NR9h5tuJJK5p3NNOUL9z8lkFPaGZWatwi8Rqr6frKx5lmZMrCBwbhyB7jnt2D5m
WnXB5mVrHO1pXEXEo9txvNjoHXZqLxNWHFMiyQZyy/B4TzDRwb/fU1nvwQtSJRFy14fG5LeSP0W6
/Ms+7knA6WvY8N3jmYE2tex/I9Yi8CVTnwccQpxcaZ1DAynGSfoyn5a+NIsmMPhwrIFvl2uJu76Y
7p3DUCIrgsXQS967S6e7nyRwCkR+4CrOlVMJIRX/k5RDtPSYQ2OHWYxYiWaLwCOYVPlCb1hS7OIw
Yc9Qdl10KC5V73L55Pj2Nv8It4sWHrvkk6plQA/48ZOoRgRBWSwHc6miYu1gcjk/mLeRdVPP5z9u
TKQ1Gywj0vwGwKAbLWJZ2NeceFQ9nxVVVynIekIN+ryIwbQ6w/dxtNvcFmUefhj0KTHvZQCtsm3+
9RcmrkdK9BJiKEZLfN7qt9JV8KaP5JicTB1pYretd9VJ9YGY+TDSUQ99jSPI6qXNIIuWr5wNV0Hb
TvMc3DI7gbbEd8jtcBODbdk4Ted/AkKcO8mvs25avm4kyjOzKj10gsLwVQsf+086gTy3WbInWMrK
ds+t9eEcX5dVIqbwJnZrShvlJSDPyu5sPiu1dxpZHoBNHCycIKjZB0cCEcmYVCXwGOkgPF50MfEK
yY6fn/VeKQTN4YDi22w7iXRJL6muv1JaIt7s1cLGqL0+kfO1TIj5/kc2HYIlrT4eNKjSUrP7uF7J
b2FMbBahaf5tviZmfWwYnu6WK6/OFP/HMRdpU78gfen37FkzNSR8fqniTwdFmuUdw1Vbh4Yn16L6
LtdI4AjgTa7uJB86yD+0SSDuBJHeMc5aDDJ+Ld9N+rbrIbgIPuaoM3M/kjb9XILWGXEUZg4sLWH7
jJpWFQB3SBgeueRWumRpl4CzSFbXl4OFhy/Sc3Ect4qCF7t4SKe/AjfrSGJndgHU4ltAvuZEsuty
bfeuwT6cWjUgicHKuTk3QaGuIkgBcXTmPBic1QHCgy7bq71KE0aIj5yunhHIXEByPFfN2/S9OXnf
IBUNGUlZZWTTJAqkO3AHOs8Ievtuq/sh4vdBi+NgDp0s/sNPt9+j//k5ojVf23a7Yc/NFZPRaQ6+
mWk/JTsrr3KZAAv674YKR9nYWapgHYydGf1jXnzmC/PFsoQ2S2MBffMTJ4+L73+yPEfGRppmvdQx
QIeapJW6YdldJNeTVAAxA8VNFELlBkbocn+wPR7hSM0+JxN3UBmscC6DYUFm2tJTiYmPHd/hHe7R
EdV+xAif44zxfpRohA6tLyrZ8Xw70Td676C01978mh7JmwoIXq/EoiJW5gr7KiLR29BfjCThFy73
I1f+o/Zkey3+5GNY45x4UkYpOw/aZbFjr4LoTSQXnGxtM4FI7VzvHU19W2UXKbJf0h2hDWuL3Idj
bb2/b/nogdL3m4XGkpXIL8//g+XEAD4hZuH34iZDKludzVXkAEstet3KUWkBnh1ilZJ4BQ2Oihka
aQOv6hOligZMKRcuxrz6NXXz2XaVlTD4BzPwmaFKU4kJGwaaJ3F5KztLhgECqurXb0lty8aV3kEc
K/WrjW3b6qASZuDi9oHVq8U0g8/KEQm41Hvn9bLke7HsCzOK59unwrsh/Q6nT538QJ6vo9oDaVgc
GrPSKjhy1Pqh2/+GMRX2z9P+quQmhft3uSBv8IvczkMMmdUR6boikBrKJdJBN0QgmFsaQr/IL+8b
+Xu2UX6o29FWzNXYz64w52hy9l3HvE2LoHh5UxfDRvzzePKO6FNkxUB4ACGuosXQU+ww7Msrr+qy
FkPpmREVmftd1GbGDdAFNP2aA+d+qXJIbOT55BUwAcuC63STHkpcucpi7cBkyCex2uzOciS1BF/i
EmMBL7Fn4jS+XORg6PnQiLXq7Sx6ZfYV/8mgViZnC5EMj+cYOEriQT0u3JKTy+lM0DTgkw+qlUrV
LuD68pMsdZNd/M5zMo0Dhl4731UatQr5+crSqfNpVSsk6G+SB+sIhrZzn7NZ8MFg9HNdegyhtT0e
nebmZ1aa0dS0MZlyRUrXYz8P3tCH0Y3/+6gqFMfMA1n8uuZCc/CrFKwWbbZEXzr+zDSgZBLqw0Tn
kFFQA4Ol0xI1jJb+uDHWDAv9gvJXaORL/JXjTVsw3oLb9L6VGWOSxS5i3mprO6iwEPLGsrAZAws4
rbcWrM92CMWgJQe3KvlI33zqpXqrxN4gXDwszdfhrJnUsHjc9c0oKQQEa4SAJTqzrY0rQ8cK0FUn
zvXiJfLMCYiJVE8mVbkf4wM0Or56JyqusJkV9B73miZHbqrI2gyOLiHyyaZwYaOKJ5eW5rURKfiK
nW+SrC3WQhPp2VZJb9gMjZRF/JUmzATWsuQgX3HtRDgCW++1ff35lezNVgSAU7LQJTTJieXaCVgC
bo7ThU9RpgOJScx/DQutSUllRCSmpwJ0C+frx/6NUuR13pZdXiTWcTYaGRuUCHO7my05ndIGvIFA
8VkyeT/pVA9xTcGvVAm/in9YiHje61IgPslPPluEiwiyoTWygPRW80YzoeTHybxoTYttig9N6vRB
bfD94uU2ocseS3BOF+1oVwBIKM07zMLUA8EwBN6bcB8Tn6RdKc6TLyY52t4V/MgS8Eb0EuYPrjNn
b0/w3vmQa1a6Ko5WmcLt4YVZZEy/FEdHLvVygZ9LPVSS4VyMlr8qZ/B03zoyn3tKZLWcvtd4PMjx
iFHhkHDp7m0KeEedJ/8Y6WEkVw3Ckiu5/+ToS0GwrAIx1RIAuQuvGgxrE0JEA23lXjYcDySgpbaB
sE0nqaqVYGg5ipMaJTWf7Em+FyN9WVMHOUFehZktU/LCDhZTdWljIbWy3lrmy/sx59BWEGPPN/ab
KLziITzAQuR8q3rqp0hypVumggoiOIK2llhQZiYU30zFL5deU8SaHFx4VCykupLY4Mpqq5f5i3QA
oTs/PK3ZwxlhzcPzO3otG3KRH+PtJxoDzmqQcdcScD3lCooYY4S5Ob6j3AKKkfs4F8tjFNQ5hFMf
cgvcvGNGLAznF1VJO30FUqoObpsTAHwps+5JB6USw8pchaVCamkrkS2kDpsjKW0XMO7pqn5DhOAF
8KxCr2hS96qwlLV9hEFmF1CJtcnNiu35L3jGVKhuKDNERTV5ydKBf/wtUqCRIqeWlELMVx5qEJhJ
6+2A1Kpgy/JnIWrGZSfY3alm9v4CD5/HyRNaKqMlYaUHsOiWw0wVUwDXHYgtUXl0W5apaV802I7j
yQ49IC0h0OMV2xl0w2nvuMcJPGmvb/cAnZmUrV38ifHxMrmcXUzuhCrF8sgN688Wntvzvv7RthDl
sfSplkO2l/2ADfJ2u3tUFdbkLDbkA1IZWpdiA5DX9ezDwcpZnx2HOxbgH5nebVdZ+ws/A8JGEQMH
+57ACvf8MGUvssHJnzNQVhBJ3Jh0q2eMeldqYaVe9SZ/QfX6BXvf933ynrT/x/UE+CQO7vZpMBzJ
TKSJRVs5qnOczA/6WHrp1YIq8baMt8JM2O6ubXRrpBRlpGINZDGSIFqxoL8OxaTEgKp7ofV4qufb
Px0rd2xOGJl6wvNidoS2Qvpr0WsoSaqyJYpwf8Z8L1uA3aFJ9m8O7PGuFEDZRdSjtRKNxESunXEU
cZo/m8iQi/sTJTxqXpIurGzP9yW5ciTYVC6HAvmjmjJZIaR2Hjs+pHnKzT2H4IPoaF1lvp5/jkD4
sY0Csjo25Ka9iDosY5UdZYJUc37CSqsPtcZ7BK+RnnlbHFulsSADYqfPz0BZJHxDwKSSuryH8ygj
boR/rqeOIBJP2WBpHIu70k9vC5ZACgQCdChSE5QA/7n55qadQLH8JzSyErcJ3TcTcPxeHrViZqfw
PYxmGem8awcK3UAFUCKwRx8KawdsdHG02nUIFdfPorkzpVwz4tpOKBOm5aVOucnnxbq3Pzh82TDW
G2N6I3cmmIysmHL7oK3ESvLYCK+68NkZ6wMQv4skeb6dOV04XeYEkCQb9z6RaBoXb1gJDTJKWZkT
rCpejdMd+F+NjKH0BpBxEjtA/F2qVmN7pebifz0S0FnWYVDB8Dha8nBBdYkCaHcRkr92yte8dBCR
7LFoDtNjWu/kll31xwwDU++5YnrtfXirHbYeU98cZxEPbtnBdZtniZnr7sFP5WARZk09ywPz1Wdb
L+uTFvrOJYfQIpger5jOvcip3J1atao2yKkHUYcHAqrbGVrQc+a268HupGfIlkxE2qO8tteCgkf4
IvgbJZzEc0EqTIg8fheeEaXVld/lSHd1oU/B37vr/u6SNNv91iUEnLnXThANHiViEzaSkxYo3grf
Jw/BRIrCP+GQZGa0NdgWxGYHsSkJaeBmYav7lklPvjLZeEK8zlUPi060deys+xcttPpAs376BtqY
iP/3KE2vYt/vV7Ue6EesMH3zNkh7S2S4HBM9ZINkp6wKaIUYVM/zS27/RsvZLdzteMPJy2s3Uuaw
cy4i1icEsHF+ERQqgcwd9eBbforiPLfd3FBfzbtAEbwoMABi5TGxOW/xH/8jj1QK2K25MaLFKorB
kDbkOAbhSDwEECEdhkWABFnpC/rm+NSydEdSB+ZhUe19aqW+SDJvIpgUKiY4Tl+mQBTQSnCHvhYE
w0ut16xlUvEz58W8hBEZ6STLBM++c//NhBbrr1/T86jjwzvpTKbx+ZryW6cvarQX02luikBg7Scc
kwISe0DTSAlAiLJKyYDaNh+3zcnv1hFrchI2WNm1WKlEec3NhdcCpJYvgSd29OfnJEOAqq/xbZUd
0i/X5hO3hlDQ4mssRjyReR0nL66fF+cs1JTTRpbI/T0PnqNYuZkCYBAQdxqonoV+qA1DnueblvH6
hQCE9YWwI+fSQ8tYfILHdJKu0LOLY+4zlP5hVD61OPSQemkPYggDn5nvqZWUS/2BJvint3SXivFS
2w6PBDv3e7SIe8pgepiL/9ppHycw1c4KTtT2TmcMqH4nJm9KTp7fg60UWXRzVNwORI9Wj+qBZiEU
hx6Ww8G77sF3ftjjiSUCoACsGEbToXrZic+RvVkX7AGtws3zVPTOOa1qh/PsemCkBCnHC91XOeBY
avE38SiTRtecOPDTD132imy8BD5UymFDE/QXBI3C/9iix1zQlTEpGY/jg1l1aQb2GjUOWblueSxA
V9b9WMoj0cGn7W2RBmyujQPvLVm8GSPRjz6cY+xFaaf9qIMEQGGXCt0GbZ9d6dprqknNyGuzdk0I
t5csFKJPz+Ex7mrKvAvMAai6ME9PEQWsq+A49UklHeUo5WLXbDpOc2XWS0gfFSNFBGJdMGEkR/1/
bsu5QPHjz6aZstIwBldQ0C4pGneC7oWTnMwooeD9PXJy8GIJ3oYb9Qj0NRHqtPc36jEw2vlV5aH6
GZZl0mgE+myEkr1OtsMLimTRTjl2FAHbP4s4cpLOz0GhKtvWjXDjvARA5XHLkRHnUD1JnEjOzESu
one+9DD7aoN7HBHyIitv8HuHsuN2JGdafeVGYFfqLis62YawbcI/VEi41sTwwv4l86CAyI9oPg4Z
XYK1qa4LUyamNLpBMgElGmg7tE1RyfhFzNcAqQau2OvozRRQEpDd6mexO7DWvL6lmoLxaEuJdxTR
ziC+sJNdyiWGGb2tcNzFx6LFShLjT6x+kuumKoL8eBChJzZgFIXjMrRG4aaDlYpyYzKivP3yWLUY
D0rDdtJJYkDKpIQSSxSmGJDtkB9im1O/+XKwsMaIvMa91trOK953piNusILlM+zjdZkh+hy/DzQn
Nd0nc5K73YsvkGqPUoR4GslnrKOmKPVQSDqBiFauqFyJnUQIbe45C8DQeW3Wqm/YkE4eHINjRrAg
UI5POQq40WQHjpPyEzkPRjzVaTDJkMRCwe4Q06A9HNvIhKueSJfmid3SOvJO8nvUGHGBn2t1OV0M
nL3S0nhH193yICaiLRX7X+v0MgJy45zqi/fB/hEFGyyccHyA3P0qnAl4ioJqHo1HaR0r8R7I3hHJ
jOm3THOqSOM1G+8SrSjYLVSrw2BauMbGzPdA1u9TV10VBs1vi8FyefWnQWd19HDkUHnDuBjV4YnG
+Tf65IXv6JX4NjmzTOIQ3Rtdz0LO25lTEpkC7d+c4LFIJXgZfojCS5EuYqe23qRBsXPC4IoFdr3R
6A/droiOg+hVvlQjOsCEc6T2IQRutri2b6py+QHod5lCkuTqhmK28+3Dq1PS/f81CZgCjwUL3WVO
uuPxEa94EVQwBFuGIsNWxPplorxaO54wjkl5YJEB/3iv9VHx26qw5DGOrku26wVQzQUIfvbiSxJI
oyh13ANs0FKbxpP7tdxgnpsEjCmUFWZkCLewFhVfQ2VKOZppITh1LxuEHGBgW+0kmY9d1m1xSf5I
xBhL7LiMV00XoUdd7mDFyJi1mRBVQOwhy6Xqwex93w70iD9Rj14pM1D1crY/q8sNkiHsaj3D9lJt
yu6nX5NidLCZ6iR162FxVP7+ImW0BjbegzBMh0wqp3LtlYAMDCrpXQlzT2CRLZFlv8q2F0o4CzRC
FbfFc8EWFI7qOsga46uVr/w6cui4uCzgBrvqbv+brY4EmbJDkXmvXPcMaFn8ZRo2gFPHtur6o38t
lCZ03Y5o7cAO6y3FcmavsS5lZWI+OT3zRqIXfE/qxf62eSpnzEyaTmr6pEg6KbjFd5+onox/CeS+
mnyPksc8kKbSm6oUqNjFGd/Rmjr1+5+XgBqVCaeeuNrI//zyGv0RnqOGfjWoy6ZXZr/qY9CU9FwL
fdeZGhtxAZe0VNdHEjhN2FiLdDbIlLayr5Ky+XHZye+mrGwFn/x1YwOeqruH8GV44mKga8aeRpU8
uaWHbbt+kPfJo+35wFYho/qzTb+CZaZUi0WP2z1VPmD3Vnj2daLErOP/fkFCcZRvMiueK2XZ7NSq
G342PDZZyQj3laolKw6xP7A5YUZPbJjjabgrLoNL0cx6h87LZfd98z9OeGtejfPlRoOdkl0I3tKC
2jZyc6Ix7xuboQHLzEmrIlT22msUkAN3/R9hj4uy8dTu0XL7ANIrTqLqgBbMNB/yQplSvepDH9Ru
7/TviAFzBAM1rA/Vc4Kh3AGgsLrT8ywNKHxo5DOeQ5vi+l2kDm/65kzBwQQiQ4U+sYonIy9pEDFN
OdbCHJy+S3dTsk/5R7jAGMTtcUUmHo6dyb/h8XQExadYzJ0lGwclRo2Gh7WrXwYI0SyFpVNGOq6e
fqqJb+tm3R2Shi6xC69LD8QPYAUcNOFmUNHLK0J8Aimkd8rfqcLTVYz/dK33JUgpjQ+xGYn0yPE6
XMJMDdq+H5kCz1rKNJOX5bmYlpOwAz8itZPLneQEKDbWw1TYLd0kmFb0E2tcaUrqKiGBqt2foZZJ
CvkrJsm9q1EJSCatIJgPOZKgbhs+E0o46V990Yu3SOukYWRW0DTtdOFi0gppGgkYePUMWIpCwk4W
W0oIepPXaIMT+zfIjGIOvpMWDhdwm0jxlJo3+/QUI3Mt48X2R9z29gHsPt7Y+hLz1NX1/zirnowX
6w2iJ58Nus+saPISQJ4EMKchwThQYoxYMAvumLm6BlwoiglHkxtslS51iIVqwq0XPty+zzczXEox
q/fmUtJBiGvdneXFyaD0Y35Q0HT7BV+NYpduFD5CBYhm2mikIGxGnoUFqkwm0oWlG/J6+2REbvaV
q6c4ZbLMpolMNAbd1LvHGbU/igwHU7uDknEWI0wgJkQ+hFSv/ovbTxm24p8eJ4lTLqo/DQa/1B+I
r63jpsX3hNvVXAWTsB6FCzEISKZej1HbEWF0J/JpFtzAb+Eb9R4ST4zFKv6SB2SzG/dJgkSZsZQb
H9CAcehkQ/SsDvkPb0+zTdPfqmC4dcRaNJNPEscf+tNGzl8WhIFqUK9CWXY4QZpxhPamV+lXankC
47Q325AD/wWQYVGnnivsTWC6M9mTQJdzUOQD3ccIcGHzFSMD9EZimHcQGZ/3G6IoEaMSDB+E2Skc
8inngWNPe4Mv1Mg9icAze7RAFw7XUdHDbiNPmS2WlMa98Zqw1+cUzaZtnpja4PpoQNUH9/Os0uRJ
5l4Ba9Eqyuk61SCS7/nmMUJ0c4Q/7+PYQn185yEsz3YqhLg6wlECkGiACUxOh3jZ7FS/v9ND2xR5
E3gPZ6tTM07/lp/Kw3lL6bI0aG+kZ93VxyLsKf6mHv0E8NR0OKqjuZLzyUJ2TbwKtOM0GmF5JTvF
DlT79AwvE2OjV1knzGgNFJ8FrFv2lMBjkdYGjlnLxTLQMm0xbXL7uoSOZ4qXlZoGUYn1P/bW7cey
e844aFCgDX/gAXUrXt0QaNtKPNutMF+TAh2L7EZI9cX7HkV/zOT0DsvbWGkY57CrXAksIQSSL99v
o/5ENAeInyj0f/Bn7MihZPW8Z++a9LZ6FjSKyV8HgRG8/wJI1x3G74zx03WO8kBg97HqxNEhx2UF
M+v3ldALPOiNXpFtP64myVldiLemiPF99xugo+lm4otzITcWLBkKAkU5bh5S695cKMdmkkk1oE7N
wzofO3BaCD/jDpA2WeBkomCnOHhVIUgxO8K6m42GCTI0ylPMrd6A9iW2p6cNB7+nyeB+62Tjxzxq
nNGS+PeMJPwm6AdOHMBDb98j77ogaAxQMBc+nAS2hsj8rXBxjG96Q/tO16RzqHyh1lF3asNsxHQb
9zM76BGhr4iCes8PIxvuJIj+H2TVqJLAYXqOYBLmrSGpS7f1hawbw42+OePdiwATUMHsG+qrATbx
pDndhfZIl3maIuns2ymFWq3pqinlgQkW5dtCnDv2xgdqvO7tHsjy30qSE/DCLHqkP7WyBiiuX4GZ
nzT5F51OGFRX8dmJQbTzXYFLITtUlHUD8sOZzH+y9aM0WT2OGfO/R/ebV54DGzAAtcrVwHJfWBFh
I5AaqMnVcEueno94Fvv/QWExdLwZolOVXC4pb1eL/hY/Elyu66fZxtoEPVsIO3fEAtqRC/GqRJXZ
rFGogTCERkE//439KJIxBGPnfhlworUZdcDX+8zjwo8HbpeE/qvpt3mlXunD6cIRDSdOqRgdxlSD
zDhLFayaZ78rZkhs3xc9LMMpwr/I18h81OgQkIrEKJfsM/GZDguuiVOp8MEAySCv5qZRVmWb8p8/
krk0Y8LaTAhDI7rVyAcJRxy175EOu1SKknSitk4DXnlfXDkt/pvsPGMPQhVSFB0u80nzZQ+PJGLe
mYo5wUlUXBoCK+VjW33e3C5aZmiRCOqIUUif6iwHE/XA7jF5lWEiwB7nIsguEUlRCSdA3/V2aJMo
e1BR3CeNKhsX5N//GSkNkA8R7X/r/3KCmJC68DvvABxV4nW7m5q1DrVbIGJnnGmKRyTMtrNOF/KR
97sSN0+LyGOVMQbruSnRM1FIGdm7Jz1Lj5SopJLfklpxRMcQWwrcqqir3R03WVEdE+tkiSjulAFZ
LOLzTHw3eNJsX26AxiEnyP0exCX2wSHuZne18PeQeZo6pyTrkVtOCr7+zjwXJ6wzpcFtJeTo0blA
Mn/J9nbFYBUT22so5jkgna7UkIEAi6neUbQmDgGFxMZxRWAv+xjENHwsXSv0uU778t2fByYb4mey
b3l6cPJJu4le2rcRjj0GPmXjBEheZZoixc1g/9awiqMgAat9HG7K2ZAnWWMiNQvMYYDdqgJNS2ZH
W5uPGR6f/dkWctMK/pyichfVUbxjlUXVyhUoN5McSA34uF5N5PXe/a/yXBDKHIw8AE+3uYje8ZMt
2T8LcsSNbXL607zDxAn1bqfo9zX2nD1et9tH/JFcPZSz9g7ARN/Kw8In9SK4TlbU6ZHx6iCmdUdH
klAdSPWziLr9TBEbcP6OBElyQ6QVP4GNNvUEaYLnwOf0QYM9t6cCfmqK02zGZwV5DQJnK1lULvfF
w/xwzGz/6UoaRjI3VPjaZH8o8Enl3fLdN33dkLv5GdgYZrnxZJdXM1u7FsWJRHQxiUEZP9atAAqw
zLVvGvArCAlllVZsj/wpshtp0U3L6buWQ3nHUAkzJFTue4kGfY9zjQKZ5W7irc63MM47W7Zf2Mk3
wkOKv+vHpalY4u6rirm44CAxdTZB+fdK+BNYaNJQxxE1cXU0j6yfZ0UbQD+G7Z8l5P/3ie6ghvlm
aWPCTwFmlJHV5DbO0Mzu4u34cZZvstqvSQlwpC+f2NnBIAjqRltG1THxdSLQ9WnYfVrZ3FwvrcJM
wrHz8/rCt302pE+teuuGdJI0a1vEU62+H//y5jrJYkendZwj3bNOZdrE2XrCnmo5l7BukNk97snO
NBWWpis4+g2kXMhsdhz8IRas87k90Ffp/fR9lJXqAA0D5CqXrKdgnkAigl5fvCWi4QLyQRkgGgKp
W2VfDB+gz+BmhD5VvVcRaiHqUBDkW9Z0csgYNFMg4Dk+XYpXcOpPRuVNMpKFMo7GdFpqJy+5+fJY
s01hJO7MbuZZROe8oUztsCpl6MwYYi/Ix5NBwwgI8pZt6OEXPb3/rPsdtX1VN9TzKt1pShJcJNim
V84d3cmkBZq1Vedv1GA7FM/54zKnr8dhu235Ox2R2cjaUdbyL2BJ5ZtQ0NwKs7YL9XJwy8j+V8TL
vxB/8zDYumj9tQcO+NXk5upfMWr6JZBXJhVMXG+BhWlS5ZRGod26B60v2wNevFDRsUNR9FBDUJuz
PqYYySmbj/RUfwOih7SFK1mD4kTTkAfxxvgcTYCi7Q8BHcIPnwuIXME05M/CS8oq7hDrYmvysdKw
3HVo/7HWZQPa5cx8jll1RSBl9kUPETmiSxEDz3CipMREMvknI577vmEBtFMLlQZr6i0QG6S+2Fs4
jvnwQr5ZWYYv+SJPCyuFKwWXHrklsdF+GgS2sQlax/u5G9k+9Mn7cSLG6xqjVUvmKpAdM1wK4Piw
qgW8S6h1gQNgwa+z9U/8C5nusERTtQmfdjBIkgRYyiqFcLX8t0VVnMxXvFHR3u6+jyqfpbzdv3Xz
JsvIbFBuFKxlov6JDcR99w08P0Edr++W79fF6TTp6BOJ7TTx4BhF4CQSz1zK5xHTFnt7Ig43iOly
OYkqyDLLRAbo5wwAu74NFD+Q1ElXQHToWk00pJ6ZQq0Jl4ONxsSQYxCQ4zwSelBOHnZcGw1q7Q+f
dQt00TPUVJSKGCR4E01jlaqbZjBrwNvtY+p3HC+6zNLfxZLE5TmFs4y/8AbGmQ4EPeTvaf7XNVpF
RIHOAFItAnrpLoLt/aV4GMEQYDBwE1+sw8QcuIde6dgKyd5ZoEDlUH6Y238amhOmt4tqQPqAAcUA
xDXuyrYxSqvL27eG2FHMr6NZshMpGOl0wAoGR5SMtwJRE3gZRAS8Kixjriyx9A4fSDH1wK+xKbOp
IRojbWwb6l+cB+YNKzleIZul3NF0vNLTm/+xF83f4phgq76d/S7gT8O+T2fjYzns07o2lMi5Qz7y
0tbD46E6VzcpdlnL9htIxFt5281+u7truCQpnoCXv1KSwaRsozgdBJ5UxbivTyxQinhK3Z2HaarI
oeUEroJMCX0uiwScZUAAQAmtX/4hGaI/s1etxx3p2zl5ph4SQRzluaH9DMecV5yeHYtvLF6ASV21
ZTEwBcaf/Zyk28R8jpVXwxFk3QyDrjdxfIVfifgfpREbp5KxngYd52mdBvw0okX0zcUBfpNB2uko
5sgQookAHCOJREuORXcycvjgw8bO8FxRd6f01C4omFHVC/epArudRg6W3M9m/2N56AFfjDCGm1aQ
XLIylvJB/ZgBPwbZxur6z70rsdL6q77MoGAzs6P7IBbi/DYWfaisWIMZvMp/mEfS3niGWHI+B7E+
bc2lRu1Toh+qC+zzjsYhlP4yP9k25EEl4z0CuH/BPnc0KQ7QC7U1dJ65efxy6dr989UmY6PA+wE7
sdsbpxH81X9O/EutXDzfZyjhz/5CyAwkhb9/hDwZ8cPaWNo29trVbye2lyqoS0bd6UCLw8W+MaFa
7meIdFQjCgyNjDSCm+2HVQP3Be7lyiYHpb+seurIhScrLh8t7kTdC/yCd+2Xb8A+U/zw+B4y1y7m
+LnSzkLkUDggzpASvNATHeCqzGLu07dYDQyNsvodwFr0b1UGzs4dAifWZ7FvXbZdvPeV7HtdYfk8
3lAI4ooDKruhxox8cq1TX3NkQH3f3e1yf6QI7hvfdh2rZaejZjjsuyRBOYKAmZEVkTfVKE2jOKvY
xtryVEuhvbvhIU8gG9gWB05uleBurDdax9Y6rqnOJpHvgMLkp4tqtLtQgY1yPZLZ9dWHqp5VIzBT
cD2x7KO+xgue+XCbz9zELA08YTwRe/QDpoRR+smkqinEjrszihntirRNVe7tS7cOsX/G6rVjzWc5
l6ITYAu0BIDjRy9IB+7AdtAn5AwVtuPbWi6kn+7NnwTbG+RVf9+PXFWSFEzC/pRrtyq0KdWZ9AHX
7NY85ToW0YIFuwZu/CRsE9V1pLrIIunLLH1ruyD42nthe4M9E8jGfkc/UUVum44CR58NaAc0qEhu
RwQVF08KWHW3jQb3z8hlEaWBstpH7Osc6Yim7jS9hPOXvElyOMh4PL6OXj660jylCilKI2k5jGOl
c8bbrSenDDRYVbyCKPhZv2hgdYis4ZpURxiY3FJilkAC7tItoi1PdZQOizRN3gveUA5bf7GCcg3n
K3oOw/kYLnBnKtuXHZhjN0498tEt2SwXS3dQ3dZGsYMCGRI/um30Vkg0UYM9P3xURVa6i3ZBShyd
qA9mzeR/f68QmumudcvuCy1AVgrRlCn3Qwg0Wpq56tfZQkwxhgizgRxv1uehYh0kOxBZClAJqcsb
FaNDyxFjsNmKwL9+85fUy5LpHMsjWfWL7+iCPvfQwxPyVoF2eHBKC0xA4o897JGM7mDw/S1hY3wb
RsDyYdZ7QzBvv/kGPsm6uWLaGHy9nHU2W3iJN5WGyxWpCBWA6fAPFJor7cPkSwupYpU246m8kmtz
rgbOAvoM5V6a5+0n1w7dWHn1Dd6kOOOHzgkpZGyEg+eRimTyIfQQV5ElEq5SRXh2iKPUSX1rYy7w
3imcc3O62NStBlmPsVl/GVSOaiSqQ8ZRPR1YU1r57ZiSDyT4CNsCN0dijAEQFo6bu1UXsL8N8Y/Z
A5tIaDnxOtfwe7ntPFe58DFEnYmViu3RrL5Tzu8E3Z6e+F/Ye0Uw8mq6DZ2b2NrPamY/wIdXGyqa
ZzpL1IOwpmSz1NoiDdwCJpoo6dmvApoyTI/jITjKJRQruI7crirLfalfeTQIPqfRwnnpr7VtnraB
KjA1+4ZvruoeHI5BGR46xfPtWI+4+L3guGnMtE7idHKg4DLhQe6TUhkKG/fC0ZbxQLrFGbRUG8HD
citAgfWKPJACyuGWvwlSb1IPErhavj9KY43jB9dK0uE4rdOXN3cHI7X7ZGTNxhjD39St136731RO
TtATRCRrNL+Nubh5iBQhqwlpyABUXiYqh/IYE141/5xF0Snx2OBodcpSy5fY8Pu5NpC0xQ1VHgLa
RVn4NPaUQYMjWb2pnefPoU6PHhbe7suJMdx1iyanHnhni1U2eCGz3+f2GdEOeCV1DltzLL2W6i7k
gHrE5zKn5bEcRv2T2BKpYgC0hnZjbA45ctks8RZcE5PQnGyPi4TAbN2g4B30wZDk70UVx6JvQHAX
oMqe5UK9MYTbqVbK/HYnpC14IA1DiVxg5NQ5WU0LTEr79FHYwA4yEfMw35VXaCtyXsDFY3mbYpJZ
Vt1KUcoMmHizcmJQT7vCC/Fx/mqxjTWU4c9q/pY2osstYBX8kPU4/Ff1LNjCBVD2d715MhaqtznV
Xfp/e8WDNG54iVFJ5nq/qopJDX//fV9+3wfxpcrhchHB/0Yf5jsR+Uzr+Auby/EnU2/3sKh6fqHh
cC6LsL/Zl8Co3RwHL0BuB1Nwym3kEdhWfpM3vz/Dq7y+VcPEqPKWm53afeUuyks/4l7JkILX6Vhb
p8jCc0OTr7HW3Empnv4p2XYvW93xOuLQjyKol/WPV76mzIK59s0F7+wLiG2hz42DqrFkegRSKu3E
iDUpD0NWortGKvstSt2VoiU8lldvU+gZc6LFQAkCg7QsxGOOlD+CduZdzvKwU/qlJqdJbBMRKdNg
TCsyCO2HAH12Hh6dfbilWPajTh2BFvucClS1M8tkjaZbzoqHWq/eV16E/H9qR6VIJY+00rj0UFdK
PtrYZcBfPKcMt7MJGYqiHawtW0u5LVvft+B7L0DjvW7qfmDcHvJIRnpye2PXJk5drJq3JtNdT1MS
Qz9Mk1pe0qj3yP9faCcd8BSiBJhKqqSaSeN+ncKZjjorNKNhAr2UC2QmP8oXr4GFkTbtVgZ+wk3c
5on8yJ+neIXVxx48OkpEx29eHM+6F+49W3IFlkoj6NXwq01Tq8n6PmCt33m23OJhtLzAKO7Fs/8t
LzLg5F5ccDDAQg3OjcS5OH/ADXwJeNfdlb+Q+zxjQouR+JMzxBExMrlfJnTRTQfiD61peT4urSNp
BLzz6njsNtA01u35mBNZhSAveABJxgfgH/Xloh1RNQCa5Eg8CaehOQKd+ysHSgAVK4sB+YpZ5+q8
CaZo+0k2RthqTsZYB/5vjp9XK+iWrIiqhy1rsgNNgJ2LYL2sTc4pxkJ8Eo+1U8MuPcf6UkEqqC2c
t1cSc7+zy6t2aHV7QyYbt6R9UO84zUVPJEoBfTTNgcVW3t+pZ58R0oCWozmmQb0YEOqNGbO1Hvs1
mZaFvqRBeFMSJNkX90O0grOHR2AKqiaB/HjvlCO968lK5EZp2ciJf+RW+5e9C9DsZzKSzTylWw/7
WQ3sjacOW4H2JjWhC9ED5PSLkiq/Io34NGeo11tPqRSH0QRYkOxhkHes8HunFJn1SYQnunn+pocp
2o+GcyXoVHhY/LHEV5YL4rXUj55gSwYl3NAY1YN4Xea82/mzJNPEOVs7Tg0Ja88BnALnsyIO8in3
zYSnhYtv9xa1l/i2p9KkQSZaCJb0s3Y3jTg1Q8I2GbJgJZ+GFsEX/eyPsCWlM7/a3SNMJf3x/aYY
4bq2iyNXCTf3C7JuJXBDt5baT10psIB89ibhakut+aEVSx0fhFmL4q3N5AiQIul3ps2islOe0Vpr
dTVVhLCptwuMAiISnAG5aTOQscZrOYIzn6kAdz4NUjMM+6SQk/yd9rEHHgBqZdYfz1scU7+dyLzc
HAUdn5xAAQBI9l0TQxXPR2lj6JdyXpFxvuapvarkqvJUvaNcPLbu9KQ+imM85JcCbSOJASl7giII
oiGlpDyMVXh3gcLCPrdu2iNpgyoPtbfl3HloayLdbyj0/SzKaUYWFkDluhdnJkotlb1xs8ukFLmm
SiMeunvC3h1chK9fLce/dGZdy3RcMMGs4RquAyoUMZQ/g+n1YxqiCQX4aur+dtyhW5SAyoGjd6wM
TCN2uGGrlQzhKpEVSgZdCYQLnuWLZea7ZMix0V81Kj/mFaGrX2ZmJwuQN7vneiVyHi+zL3HAIgk6
l5Gq0IcQUC+r2PvVTvbR26SuywehQTEzhosFWlZTexXnZx5pdcksC1rahv4ZG8gry2heWB0Yixuv
0qfhgqcQr90mNpUtC6arx/NQb96iADMDc3t3b2njMxdcpFL934RzkogZDPjfDtUHgFdmoTYQrbek
QO8n6zF4Jyfl23mCPEiztBXwOPvdIUMUWmPqB0Xi4mO25ud8S9ysw1hfah40NXAjxBk9tXCfS7dD
08VfTNhbCKVeTZcFFdkYeGM164pZelN21NtanADvReYuSdoQltl/bYsirwnhtCxAYxdTjJFyRTOn
U34eMpWMft4PKWxggYsf2exzssAUAWkeI38ynZkVnhg4OZYJGiQta9L8n4IRTQgtpV+CLBVxbxHy
midMeFP8vVZcVDDoeLh/hmq8GpbheoG6Q1+/lpeX/q5noMdlJgqIAv8y3Iim228tBAoOSn7UEKpl
Vs7o5mydh02Hlzjn0TVVRVjPxLnL9HDaLO2aMyLDBt+oNTpwoAVej2C6CHv/lDA5GiNugDaBGd4N
8co9N28Mv4q7jCd7hv2q7wWKxlTwK5qH5Sy/AJ4s37l3SCw7Hfkh/VS2hbgshb0GS7k97lBG9PNb
aeykwPXbjfYtbON6m6Fe7Cmj1i9STK46kkJIhTKc+xjb0wTfdevBVrtzzBtKxVuKA++iSjt4DPkd
SeAM++LCzQ27bmdAN3RlO0FfLa0vnVokZcx5/R8EWrIKLQt1V9mcW06GGEev5L+cTkSbJyOlY7vx
Mi75Z4uyXS3x9p8q+xxLIfnn166eXmzJNaYtygm9L4l+VbVdSF7YPCn2H2/fW1JPx0nu5s8flAkF
ysmaTrjWRibI7SnuZAA844pFOla+6Z67v7UfXLJaNUJlghqFnPvL0Aq1MVdONTTmBBUWPX+uQood
DkJcuKuvXVoCm7WJqY+Fp2E90wgDr1Ox8i3sidxdhP5CLlS80MNc2YDzSjhHAi4MJ/qvtafBOfbT
UcZIg0Ds+BftK64CLZZHZny8aHpeDi1oCtLupQ90NtZQfEE/bZIrqUkT8vlg8vxfjYRRdhv7Yf8S
5g+pwBch0HsboFSmSDTrbaFLgwpR3vwIMOvfwdSbVAM3tb/ojM/9egZkhWnPBO3irjErqI6qQqHN
PXIARluzq51l10mj192FOB3KQfCMw+ffkJmppR1R+VmZsC/78yThLHxfNDyr1rLLn090YQfQ/Cm2
MaO4mifLVr2IHZSsaftIGg06gSNp9fvwgdjucUZRbzkwjD00b+N0Az5PEqcsxZhf9ETg39jddhHY
jYK/m0ctwbdInXKMw1E81OEUTRBVnvQkY7PGF2MDQnJRptTU1cq3GcFzy+H3e34JL97xwPyqSb5I
c/BDZ+2DoqpXAssHTMGjmrevG49In/tBIzfdOU1F/LPZpzpIUS1KaCzKo7hDfkKXZSC9pKKL1Qwu
pXxdj2ep8NdXcmCOjOG4NnfDyZMYR15KDxbUc3u5SubTz6RrzpeOnuyo69OwC7epDrR4hfL5MW34
5IN8rrZRdPtIGfB1jqHJ0dd0RXkjdDNYx+btNxRo9tW6fKkLNfYefgpWnG7LQ/ZL18gwEl0NWtAS
sajhA1w4f+XsfJyNEwPtBvIIOQzEVhyn+0+sWhX2KmtqDp56d2D69RZeIyrArquw49wsp+gyRy1o
F6LoHAX2bpdyr/RVBtwNQS7wLZS8l8j60UMrYMUI5pezD4pFAf7hJ4ClgAmBQJYeNAd4wEosh5Lf
eWU0Ca8ZQsB1FH5KWj5UtWsmtW70QfAe9KnoK1AklQQJTLh1eVprngEXi7OALqJK+35AaGwN+VAc
gQcp51KhdHz9fJz5MKnlxdF7JbRhxplis6WOyI8DtQaCb7QdfiDQQfKBieoGRvZMdWqF1Sfb8mIH
NQzVHgP111qRxlMe6F/TlG74FvVdcKjfrSQAwLU3+//azcXSaK3L4+gn9fzln9VK04V71NAzqzUa
uZzmhDJdTFiZmdOHK9eDEb/pF6msCcjEZu1ZKewvodl6c+RUii3rMr1UdGGKZKf8iySLIcSezaiw
+IWPFoPFw4RcQfh2G0FcHc/th8k8l6b8kYmzwMHCxhYTXVPqbT04yIxZTAG4Mz/d30qt2UE6yJQR
2Q23040lds13/zCvfbTeOqi2FMliqcRJ5JTZazSGfQ3bTRCEngJmltBBpI2UkjDedS3DZ06Ww7l3
QhLkGuI8RQDUm7KJPsGHCOoSVJMhH2Adn12HvLh0+Pipda4uIaNaUZLZ/XT//mqJ7/nnHtIdnJ4u
Djp2FDY/6VCklc/0p6KJKzRIUjutxhA9EBwk6RlUHHeZqyX9hDDbXZ1kAzZUteeSwhJdFcE/yME1
yiIJPmCd7o1BJrw9LEH1aS/jUHYo9eHH3EjCsEBaO0sliW0grP09AfriHFGbgIbyr2EWkbNhoRjK
9tzwkJMcaNmf0MCCeSeEoDXVEo/MU86euflA8VuwrQbG3stHXOqe9Gk2mOXwxaYi8xrMOUKN9iml
xrccFD4QiZljhBTDn77GKC+qjPxKI7M241Ph5H+mTzekYxifcG1wSzAZogNWmXrsxEhBp1m8+6vS
geDvC5PnWg8gt2VnbaJRYfc1XArcoRYzNH0XJDm3OHSwd423v+8BtMJm9kuQCaz1SU8sdayVJUgs
sotfAQJGCNN8+GNltTYq6vBtBDcQ8/HuJX8qkveus2G8e36zKYf5vJ5Vss7XhzrzWlZLm723ErEC
HGhP48A60o8QgcgFHN+gK1zfCuazI8XiMpHU3JEs2+Mm26M6As41bKhTyF0CDCbHfwnwdniBea/I
E2wL/B3CQYOcZQzDO8Ca/9eYdMrGEktWg8S0AVDYg2oKAZ67DHU8EvcHGUra2dURzJynlGo42vO5
iV1x32PUx6/9CT7WKQyIEHJHnipCer03AyxOYhAnrwmxrSvA+004KPXDya/vaxiIaifUuvO38IdE
IHkJpzjMhOoOkqUACSdtqYbK6pu4bBXQrD15yMEJYzvAtBgFmLrwcIpmpOln/wsfOFypbDMc9EXa
UHdEmnS6SRVWItRYICBoG+pRSLbMygGMrxsgsDAzZ+HoE0Zq7ZI/mdNxQyU97M5LkYq5sZmZQehR
dhWLb7CeJ0qtor82oPLtiSnRcfTIbh45RgxwjKNGBbwWANQJ/OOWjBKkriRkZcPmHrBqiXFCf8AL
vAWU7q2tdOrfDKJLRbXbJgX8i4dxP8JMQ+HIjcQnnnLHBQgt3hQUN8ChQMqeqFwUl+Tg3FkHoSs3
cdcfP9r9eTP0WLLlZ26nW7RwFyDJWtGU0STxtjU7KRt5PZSoTumvoMXRwKGmAqVDYLAU4D1VH9MW
r05iDuz0qJR4lFOb99XCLmQi3g10rDaLo/UjfZ+fXLp0y/KChRn1V8Dc6CQB94KYirVQ5WpstTb2
GGUROUZ5qgYDmwd8/r15barr+U4NXpagGr6C0XkgroVfWd7vT6Zcx4j6NPXy5Nt0WXMiSLOaP2eo
XV86gEMrPZs2bFOP4GDOTfgrjYV9e9urm6UO+rpnj/oY+1KnEeHapSRQUjyeXPE/VnMXX/u03oxW
rv4ZDQr3fk2BuiF9i6DI0LbLKSejaK7SnHaeMg50r1U/X28PP0Bu9UEsnkwXf55XiqoDwRmb1WGD
IhZj2ZHEKjLLZ1Duw6VKWrb3XvCuVe1o4DyGzOTnedhDJGAuWDtsbGSmOJDaJ7k9h3NM1H60+pVq
er8HGV3zhglyDqmrwfY7huVnBA+8kDup61mGMC4EA4EltEjLh1d3KiwPYG/8iJrvexixSfTrliX7
uEivFlUfxHnltiIA6PPhwKGUtAIjeFOsyrEGaVliKYbiARdCDzoNHybK2/cHRWDntY1vxP1Hcbdj
vzba00tSfSucvXMZvMylrNSKI6XCdJvB/U94B41klUmJ324jtQmwkLTqusFS3FL8TBaPiXpZEf1i
f7GAXVCWM/8u62UNtEAJHwfxSSTMzcHedyKDUEAQMvdc69URDTD6FiWXDpBLhdLd8+N7IvYZ1Bl9
Ff+cPqVQ+XOWchZv63mtHaORnopwT2XOntTW10RFYaBYv8TAA2lys76AJ/2QOA30KtQdUBvc9r5m
A7K3LIWtf7ZwIMN3YAxF9/RiqJWaEM492oMZK+VQE7KlYqNLyxvw9My2aBZjtLFbd9DW964aoqn3
SZxmYRROlBgj/Nsbx3/UmIFDuiVLfZhSJr2B+uF4VzaJhiErKe/16yAxOQqmomVcKxPgkGHeSJbo
tAKheElcVRsh/0+cXQRsu/FYmrcV66HIWgynF+aDv1vdF8PCdnrMxcBEXYIGkybrFo95eBeS4CdX
R9pV24gjKNwC35WRNMP0GI/MJaKNdZzVqcf46TnLgm0Qoy2XEyk6xOpvifPel1El5N65n/7tUm9V
HJiX9JMezlFU2rY3oXqr9xCKUtNYzQBaUmYqU5SyW1w2sqBCUNSwRzT1WTiP8PTD9724JNfGMlS/
JZcHRIoCyZZkvs6urAVuAeCCfsCEtWymSmJo9ImgbZWXsRBIsQG46sWmkvKyRap8i/QbZCSOaa1F
8G3XdxXPx9n4JbUNt7bBILKInLnAjjVdLlv/3ALG/8GiuWoWVd7tJ1vPxY5jSBX3arHll77bP8kc
F4B7TiJSE1TrxkcTyid3l24FoTIIytZikC88P1KdAJ7G2nDu7xVbIMExGV+A/YMH53wYsdFvk9Ax
Z6TcCZ+hm0jtHukNowo6ny9vnYiqRutJyBzhTeeQ5rjfG3q29CEI14rL+aGeoQGTsuO50g45d7x0
w9Sg1/YS24dScJ3RXIALAWbMR30ajvk0WQx0FqRo6vsP2IS545fDpg98KKEZNTE4SAG4uwvowj0P
RiYb4FINmlNmDhQt8ivbO+NGxPj4RmNyvqBNidq/6chR58ccD1ymvVKz1iS1OYNeVt4yi4TUVzr2
HHTVlDbMr5iMdLnfPNG9q52iMEohh00AjPCzAK9O3fUeWLY490sfY1AGlkAGalCXcQxfzikKF9lC
ipQVmw35LuiKJ6Yce0L39BQYJ14v0j/Mtr0uRio5+UfvZihLU2GsLS+xYh1MBSBM+nsBb5q2AXg3
s/stx/PIJqGYG/HruWgpqJ/+RrUKutZlhAIX5TBwiHaFC7cVHQ7/Of9BSm8wL56CXMzLla8JSljJ
zaA3thmVrzKtYUmKa3ekIbDLpjmu7bVnh6QJmrFgqvK4uWS/3oO3rEF4aBWoCA7ysUFUMK0IBpl3
O41sGHQ7YGFciOukTJ16cJ7NvSaZvJdz+3Cq6WESkQ+I7L52IQx90C4BurUKF2XXFw5MBd0eaIgM
FGAai76jUDtCMWO93yvlayoC3qw8xRLWQIZUeYt0XjuS7NyZsEfvrh2jB0YnBmPCZFtg4BHkm33j
o4LhIgO3Gf7JgQ2kbGCVjbJAGIg4ZULmILYlhoQbCIOGxM6KiZbXTiVQfQO+fIqnah7yl109lWF5
SL841sqJ801G0WwcJaM8Xi5nAN6QBP2LTcR147Xbp4yLiYl+3hodufjHun8/q4mxuU3IH8ocBCoh
RH4HVkqmAle6UrQcJzELThtc3vRHpcnILeiPKMC2GkVvmSeBS2EvhqIs9FOnhXM56OUsu0XuWXkk
anI6oJM9UPGqRCnUAlb/f6aPg9PyGG3KeEhEIOP8JISmooGH1gl5UDNL2vWLhgMBponVIZMJO2Ya
UF/kq1aGZZE9K1EIiaVG9XTn8aFM+QxI+nxR5Bw6OkvquYrNJXqweiUui7XK4YkZaiJbVjD5lxTz
XLUK87bRdNO4Svdx+xKiaWRVeVjWeMqb5TbzJwD+h0EZVscvn3HYyaFT35vTDXi34sN/c3ABY1Nx
K/+RGPlB3hhDd96aLRMXJ1sJaumKmJAKs52vxrdZV3DF1xuY+IrJqf3jl2m6Dxtv3Ft4f8ZUmTWr
FKtocMIB683Xecz6fymHGE9p9UvymL2v0chqk+HrsMCanql1umAkPSQG9QiBzyEuohk9Te5+eip/
MarEkWO6AmZ31WndZJ6Xij+oMcN/KTntjSiJ6S70Z/OmnhgCz+CNaSmb/yLpc1lI9Leomf7LDjE3
jJZ3qZqrmYP8JZDSQHyLBl3mfjLenRN39tMJOHguU9iGlHSsM0QMZGxOeE9IR/gfTjcYjN8BP+cZ
YSh0BAiVD0xXLPVuTb+tnghP8Wikw90gI7RpdCjH6LYsN4bpA/vVBnfqQOfSDvyaz5A6OiXKabLg
nVenD6m5u40mbAvLC/SIMsNkmedR8zOgGX5JZAB9cbQrMVt78LI9JCBjmPOVxTohe6ZLjU4BWzHy
PmJa5xC0U0jXSuQ6UU3bDF3CUllGDOdoPdc9p2gVY/3NG+wudaJYvOORMX0fIReFTGn5GFTlGQ8Q
fTGVVEEjK/twVrBvKdM8s/yb7dQJGLIlFYitsFlanA3nE+gMrYIcjvMDRVmQJMwkZ8+fUzES3viZ
RcW5zHlHDHDQq8Z+OI5rkCwyS9Hf7iT6+baT7gFnz0Y5pdAc23hC1CU/R/aX7d7ZvdzlgnBfGNIG
gzis/eojA0ylVfER/FnCxKgvUd4FeVytQXRIM9P1q1E6VRWkOna2Su7lLRgDGvJWCEcfiAS9wJnU
AUD1nH9HMTD4CvqY5WH4i3oujc3hU/kO2NzGwm90rJJeeFiZxVFw666MYt48Dr+2jzSPzpg8kbBl
u4VKEZI9pSOJiBkXBI320Cw7dh0Qu5pLJ+Fsesh6mUsV7SZxcOvefKD58rTkhGB/bqZMOx1Hd62E
8mtjS4wp5OJC49TYGMYy+xlX1gz63TdIzn76n5klAMqwHSuRQ3fTSC7eJcYw1kVERoOZ5oZOKAaf
dQqUTXKVhN9ApVY3Omt60YRYgNCoqNtHHnqFk6RuHbuW8HAEsycxHvtJKq5pWB9iS5/OEdp+YzkV
j1QDblc8WfBbtRaIkri5YGTCtcMKx7Fso6cf1D+fDgA7op31Av+lLtH8JvdaBrgJ57/GD0MACDyQ
VKRmNJqZ1vv9ckEmBAT8e1K0NDDi4rIzzNHQUz/oHXnZoPP/6WCcXaZ3u5CS1/vu6TK/iljdw3fH
FIVuLKgHtLZZ3/FYS9zwKdIAvWFsi7VX6AHGNs4eqHyuGhvjsQSFC8JGzdlHGq+zIjJFKbtAxgYJ
6k/JIeuAk17qrNsmG4rOVEfJmmRlIvr/agKbloWWH73Mphusgc6gGuE6xR1ko/Jo2fuO0p2fLWDn
VP93cB3zmlOQd6fMaIq02aTLJQ/dz4upKN21MFZreyQT8Lcjjj7ox+IctpwytdghR084OmIBH5yH
86s4UBm+4UGo9iT5/qOAQFA+AllExfx/XeNj/lerNx+mKzl5gDjim2rbwlJUvuOrcU29DAGbqSi1
RMNusi44vJqKbsijyhh68nXZT+2Jkt+pnb5HqibFfgsE5J7+TqoQBxlgRUecONH8jzaBRYdhonNa
Z6nncY86r56k3NX5/uwFM4fe3Rwa9xBpu+7jNoc2arPUmAsIh6/FjZe03V+1hsRiFZeNxVUarITC
9ubCh2RvK/71bZNJxiCoklFvkoxmrjJwzntW3CizLlT+vKfILp3aHpPMilfpKNXKFMT8/narTGSa
6TwVMRYY6GF0CJ2YEfze5sWc5QNNCqWn40RdS+yTamCmkVowcQCmkp2/YWk8A3q0mlK5ZHaHSX3c
5NauYIaXawEJI5omCeztax3unIJCS50ZoSA2eRm54/UUodEiIdbq7TeJHUOwM0zcxRBsSRCP8DNL
ODfKBATmMbFYbUHSg2fYj/yXg8IPTQPl/wPU8dCrk8iULP5EVgvNd9mqjUgm8LRhGzLNaRMDB7p0
Ax5hneIPb27yBWkCxMRD47VhN+49oiEp2EV3d2/u6/bDb9/N4s6upnQU/sL7UK2Mm1v7jVEmlspO
8TPlM6juLAPkIuegN1Df05HL4MoI08G1rrWJ6p+8PsBmq8bPL2wpBaqE0T3bBCurIw8MvE2ofE+1
Se1VQU70agSupfJQFn4zV30tJdPV2EdaAkHryrs9JZ+rVBUGMTxrWMEzVyffDPKubQuAzoLDcg19
/h8hpJ/aZlpHz8KfvJd3Zpilw24aKCO3Aj31AY+CsDTelKIV42+EKQHqSyibTQsG3wzgiM4iYipq
/80utfezCdJGC5OMtr1ju/c33jBQgA7I6r3Ws4yobolWKGJms3KpTFoOgr5xlxwI/eA4P2o84Z7H
5My+x08cXp+I7Zm8KPZBL67b31wJoPPWcfgyT9WvlzzaVGJoKenKCOv+KgD1+Hp909BuDvY0yzIF
j1hMLsdCAcOBfFP21jZveqMyIT4DqCVQZyECxmzcxEtP5PORSgbh5WY8FpPVj2AwhE9ao3yGhNKs
CQyMeb+/DVRj3DT1/xW10Ofh+DC88XNLV+r1/KCKnt128zwBquYLUif2wHGDkS+1BQtXSQIW9+5+
dAENwzmCM8lq8wwkI6YMR7fQCxo70ibsObuWkAXg6m+Zg/GwcrnyDNbiHJCZveQTjezueo/ZGFuH
vlxMS4dARtTXGcuwndWm3+2d8f1V+X/zAa22o6rKC/0QWJNhNgOplNDfLGrOdPmGUI9wsgHAPOJr
G9r/E+3wJGp1RcOYzxgfIgHs6TLBWaiWzp0IQzsQ1BCBnENgAsSZI+N1/Jo0Y/9i8/j1Bx5+6LBP
o3YSsH0riD7wJlBjBNJJJmQoUxCXbQV+70rHJQYWFYp1wnhD1niC8gupGng3FKB3uMX0RnAS5w9Z
oIJL6WrMZjHKNPeRPTm8F54fQJ7FfcCFAEIIhtciPJf/qKVxTJQvpyP5iTqCBYUqEDdjjheDBu9x
UIFLyFphf60Yys5Hzg3eJo47ztU1sfcHFhSmxY8xVzDcRumMgSr1GbKsorivTMMeVVnrMssLwjJO
jeru4POraMVuymvbV67y4BPb4YiQ+S3kVfK5Ordju2NcCHAL67Vsk6SN/zceugzSgDYxxoizxSRA
hX/aCN5aVhv2xhvHrfOdSema5r1h/QhLTPf34+78uX9szNYfBF/4l+T8nmY/H9//S9jrNwjXFPfK
t9Fd808+gz/9GvswGXgxwgkafT+n2Zai6rO6avPKsv0lxxZIqbMX8IGkT+qyIAGlIJA0kASzH6gi
cLNXW6uhmTjyQz+3UH8jeKwKWSYtkKisr8iFgwSleg82pw7adfkz2GnbWgiMvH0Z+mJqOEYRHi14
PbIhSLqSxvMIn/hd7VGA4c+QK4ayWptXTJ5tb9umrsy17OapsnjVuQ/lfBMToXO/yMcfy9jTJHqb
0we8HIVoTvb3aOzEKZ1Uw6/mArHOg/wj/hL0TRw4fkSehi7dIDBo1N688SjxVQLzGcrHuXhErELS
LFk1yl9o9lMPuW3awC8vMN4HBINQVlLvlJk697YM0So2GCdkjM+hm45/SJTBq6uyTXVqm6J0I2Wb
vph/puoxGgPk6AVz12wAmsLrVuRUkh6+qyBDevgUsyGG0BGaN5EaaZj5QWYXxJmlhWwbfENd2OFs
uZ5wGB4Zosx0YFmP3g3oz5FqTS1cwwxGzRk4gmT1YXFEBsJK5FykaO63LCWvh1jjdzitFcuqLqe9
l2lgSEaLAeVZbF4sd53om7+Ftj+FxgHLVJpMk7rnSXwNXKKGXp6M6/eXZtcTV7B0II1aQZMCPvXm
/vArNDa2KFNH4thfoA9DNNttmkJyclK8o/Pa/xcB7dn3HlcMtleJPqrEYddnk2VeQCrNl9GzehH5
BcIH3Fxo4IOBFgGzJqZsD4I4ffk/6/6W8/deQFXJ6NqvI24XWswn31LwA+XvIR1A8ZNfrfSwwF4v
UZc15bBnZSlpchLuW3gMGzkrkDjhipv3qvNCM9L09ivg3xjrS2aXGR1kLkxJSVQshGP6HxGHnauR
1ADvavkyPbK+3CbDLLXsm0BuWaPtf+mE3YCOsQjzbgBOqCHFy6lyJW4gmuYB6VfERSXd4Nu5X19D
l75/GONfV7+uA579yZurQoaIts+Q9/krHWBMudngUIDOz/O8QmR2ifYY0nGt0Q+zFhfdLuoIEmFn
j/mgxhW5mNqIRg8vHkP2D47CJgsZn6OHCTIYYIjF80Vw/nubpj1n80eYhL+RtkHGV0/TUUycnYto
ZwdO3RUu9bLPB8BuJs8LugY8TzV+lTcv+PsJL9KEgQkfzcGRpTkbKSNuPi6+0jMnW+2QKCn+4303
mbWfgowbFKRqQsdoxGk7tC88eP6l7Ln/eJpAnBI4ZKAsd6jVD+QHthxv4QRUp/ZYl99HySS/ac+M
YVDvFCVknBuPiPeM1X897FV+gKlzpHhRAPoIUpPwsVswbC7Qq+4x8/twBAoPR+UnzjIMI9wjcCZK
QtIZSg96M8dqYAM7xCN7gmWE8hi4+Alm42hw0D6ujhJvnsU+ADpsRb37umpSv32+N7H6fbcYFUZr
J3fsHouAa5nS9+Q8xtCe0iMV8x0ZiJR4Vj3ldyAQRj77ImC1nYss6eI3MRDbBy0Y1tWx1QlZj7mc
7m3zwPsLDc3uv7L6FFngfz02k9puXyVOORAj63fqlVJ5xRM+rSWF4SD2cclqChpZq4WG80ULtzgS
DxUJVh/aAWip/rm05L3GuLaLBAm95xPH6fnN/5dRI08a6JQcd2NFy8GQAFL5c03wB9dUDBdFifg3
i91aHzrVcfFM9jQnLWTb9sw8hJ5Xp+9+Bgc2/kWFjp4JuvXOpClhfZViAaOVy/pFbSzeacgQL3Pz
YoXUCZrdSrDyPDG/aAtmAO10bQYqkazCivnSXbyk/49/qe1cJ+Aea9EewKTopRRo6LFrPO+Hv7qA
qVZYau2kxVFZcFNEPXFAoaWH5iR5X6+1HOKbq5DtDuyhV+ENiCK+MZ0zoh+9YIaH540A0pW9YK39
G09E0ABhcZfortjIBqYY/22KKDfYv4jEUVzNKYR0J5h2TrlogvpfCFLjR5wurxK/+2txOWqFn997
cggKShM7E4RupCiF595UIEQxKZe/qYI78Rc8ui2kCZHQ1Pf+c6YyY0cWlExJwzRNrU63IVgPV85T
LmS85GiVBhzgUwKsFw55tuMnkXJZJLtzSTWc5dc2bE8ac4T43c+iy14NmZrdwrwIRVm9P82YIGCJ
Sd8ACKgEYT8QJo9AIikbvBZKX2PvOi/H9JEzfNtfJlfzDoDYLjXmZL0YMeN469kNshhGrXcNwj/k
qDZl3vN7swfTO5E4jDuIk1EXKtVKZ05csvU1IqYFOnz4lsO+PHAqn30KP5Gmnfds3t5UW0T21Cas
HpxdWN/23utewvDJc5W41C3tT3kOhTuntQXkeLvQ5/Vu73P5IPPycLK9MerCYwQezPPL+JElwKsO
o5vjlcRzv14Q6NMjEJFf+riymNEgZMqfu1hMUlgcI6wdIQ59sW56EE9l4u13Km4m85HkZkWRwgez
CFjngUluqOmN5UEZPa5ii6psXA4y+xVdKb+DC0S4iixs3mxXXf88ofa7/4Gj8E0efLdbZMIryArk
1n0eQb3RUb0G3fPzvyZD4eBt/I3w5/XGBccPLtoRnTxpEKba6nUPXzFxeGwVjmh5rlIu9gCeX06U
QpN7GM3ISBJfuZ6Ju3CnuAT5b2Fk5tRrn60cU7r+ULOJsCFZgrES2qWMjyf9dmb3EPICx7EYxw8z
syUtEn2GoZWCWdds7LF0JRoXAWlIlb/IGlXSiLqy/IFIZLJp6eOEJT7WL2mJfCoJIntuwJKRwK/c
kKW3l6NelmpsOubkNFTBLczWLqKuYqLGZyYxqIN6Hg3cw9WtR/8qkOF7bGw6SJwAXVdA/eiI3oGn
ynLie54h5iGu4jPVsAxXvAROAHe1AZmsCJpZ3jmF9hfGdvueT4HgXmd2LbkwGeBrvd8XGY07qzF9
xuyApkM7TgnvJTaoj1Lw1YzWP8zcXgZ0nM5MadR/jNpCm090xNQwO/fsuVyt+Q6zJqDZyvFyfHnQ
A4dIO6RjVHU0+yBS4iziJtnEAwhKQPZFiEulpj0zqIWZUdJVvushjsjQSB7eBdSM2DBp8I31RrSG
23fLtvbWNPr9EAqEe1HL1fDOGw9Z1hIK31nzWqRNaYWAM14jnbbNO3wRDwicFDPmo+Ki9FkXHlWv
/otKJqSb0+Y/Jar7P2SGZy5pDf6oUA2wiU+Omqh2Pl2kv8rTtC9Vech5trSCXnn5rfZ3+G1WiJtD
kt8TnOC4p9GnUXej6TWYZAreJnFpvHOAdpRPPA3fM/Es8zYWQwV20DIv3STXKV9nxM/MShS7cK7I
fL3QB1ALrpAa8nsz0ML1zccjGpT2flZq0VsdrApZxcMsyzyaUB/vvkTf1c9AxzsX8SmZOrcfCJAc
/E9XusJaJE8JTIgKB5CxvxOAKp25IaUdH/FXylaJXCN8HUksl5rcNEBiBovvzMWakeCIFMqbOUSs
OLAlKQ7dak05KGXcEdzxeMqSvzf+QINbHx3HUKsxmb8iq3jk7WsmL9ek5fidbj1oQhGHLuYXhCty
7B7cIABqB87erb8/g6pY5zOxM5GaAAmck97FXbo/F1EDyd3zheqSYR52jJtNcODqEN/USj86LgQi
SyV0FgmaCmBM1ZxtiQpzNjFDY6h4r7vDGKuzB6YQ/Y3C8P+NVHBAHMdqRQ1S8jF/Wmvda3o4Vzrq
ihOK95EWnGq0DjxxGw9VH0mfwPaQaaGniyJZ2WyCZDDsu9Ie3eG1S11UTPX7q4CoKWsncFfWqyLz
ywQdEXEtOSVFiOAyZyY+tLVj3HZSGlRbBu3gYFU8HviJzbc8F2ndZV7K/i8a/KbX3gnVjWjsIigz
NqSjv5jBdwVoaEvn6i4GZa7khexdu66fQmStd3LENGKnQ/IWMu1LZHmEybYGpNXTYpbKGym/RPIw
R9jUdfHCDp2MIX7oijgtxy6uWXRQzBMspbG4xuWQTAkYAgVqZcFXBlfQH2ch47CCEY5hVcxQWysH
SmTYawAUGF1GqwezOWStX8Z5Gwj2OKw6+yV0+89g1UDS6339iNkJP8Bb9aP+6LCptaDeACBx2w8/
s8w19SBFWucYffSXmUVLQdyqyF+qe/U+1jGI9Ql25m7IvYkG1M/nRZeYI27GugCFUjg/iQRaayfq
FJNNY1Nlw7QJK8pqqlAYu8CJA5Gf88U4psntR2Zxrvc/bXIS1Skk0F6btQnsz+SjtRo7kdx3iEzL
gZmXgKcNkRB+osHE6/T0mgLaQwdwLzQrS/E7H85qiF7o3vC5Vw+KDKt4Q1Ard8mlPnim4le9Gu+N
81QLpEYkKI21ToqaWMeTuS5Me674OSPJQlwwpF4b5wgzas+gboRQ/BZr18RioCMsGmEbwb7oDhPT
VG2s+O+IUwZsqEQOHKq/W1DQsPu3ppLSRrVwuNNOIrLHb9V2Zu3vHxdOeSlATIfkufX6SbUJCPwj
2eXEEQPMFC+mXhm/FQ/hsF2Fd7fer7sqZLcWNeiqyoUNkOO0Q1bALuF8yFeYBofrjxexpnhvYlGi
aVQkMNKTWObdgZfTmq58eCvKmSrXxYQVTqMAC3EApg6sI68xGRbVzBNxD8rtX/TG/iGPPmC6bnVz
cEdEwdZtPg4CN/mYIn3Z1Rbtn9Nfge8lKQ2k3XMr0Kk8JPAlJNNsSph0WwrSizCKynoAyPSP8Tcp
tmrQAmeGRPkPBqSt0to5w3O6/o2eNCTnSTkiHdgYmiJ4BJu+YZn5RUpa/ssu7uRVVKSeR1vP+XT0
T/KzVCxqVHqWxbHoYV4Cj/PhiiT4+QPogw1KV32tPUrE6h8lS8Y0kzrk1A04Xth7p0Zyqqbp5dNo
QUgkAVMheXMDpbHwbSCGzGlm598LzPS+ErWATpNuDhsy5AQf83mJPQVytb1kD6nxdtJZ5N1J2C/i
5gCwTw66ktkhB9vamTjl4KBsP/8hCk+W/XLb+RU33p5WiAcKehAzdYg39DWXm8v56HJoHpQCiAZ/
GdOydxyXAeSIpeJS//Mca7UBp3Ud8bqzzViH0TDessaWoKJOX3ybAJrBBme/hcU6ASHMTF4Bs7kT
lHfPuJ0J4HBlxga8N8npHcev2K0SK/atI90xMg63R6ClfKnPxlklYk8QAvxCf8UnFASTCZ1UAz2C
Ma3comrX/qFhuFZrlH7ilKE3oy0vr3XUStkC1aag4spOdm0KaVuORuNhT8DzIVuts12c3yE3HB7b
TLdeaotRUpovAcKcL4813lpc0K3x+lrDkIgjJvZcp/1UygtmSgeYu20ZRATaXlbXsE7SVxZw6IGq
8fozeSdA+5TPgadhR/6NQFHY7cZOwRNKyZifAgL7jm/hzYSc7mjMxr3Og6QFTY7grmUnuFydBbM9
oFYee44SXLSYv4obqZxyAHfUOxW/1F4TKTbFo/E67G+OT2tqmLhhuAxjKT9Pc5RM2YdCLz/iB/mk
zJ5mwTMpKr6IxgkAXp36MvvHEraRGGjk26P2cJXZVBZG9C37W9VfM3hO0wOl5KV77QFTlDnABz81
ramaCjjQAjUxtXJyoorjYtL/gM6bxhSXQg2c/Ss0OlBstrAoy8ble7Pef9iCDUoHbTql1XRDou2h
ZqIgyDKGf9pcJUVwpkXg/NfjVreNRrp5EYE2H9/roJJkA81e3MNvZDtCAzAV5Qt3xKPJLzTmpJON
U18/IKfRMA5IDgua3eqXO08LFW5Agec/Xj3W1okYvUf+jK8tM5Y6u+1gc1EBlab2Q0epTmuXuNcU
dAGzRbF8aHnczvZ4Vvtk9q9E/mPSi1/eZdiNordGcmQ0dZRTVtPvJi/PSX4ac26sKOTBpFlE2k3h
CVGhXCLa/pO2FSNGuYkOSYJbPhkPaAhUVpjnqZz8YeNpb+wqPadd5TcL7Mn0f+xMD3E57Zyo3EHR
fToEm0mqLJbWcFI4HDEiP43HyE2uw1S0Z2P7ACarCdS6nU/y5y3Aqog0S3nm5zRoIxcaW+jwhWZO
ufmw5MgMea7dEOXjwupiNpv7HynGsdFuncHl/+UtajlP37n0lVrFm9dfUeKG5qgnqOJjulH72NBF
YMJdR0Tq9T+ZCjCymN/lJ8Uh1BJvSrV3s6zy9g+wdA7yrlty1TWzKJMBDmOEsHy1TFH0tM7TMsVJ
waYjaM8P+dmWnCnL9v1qwfWKv3cp5Gbyyrmnt12PtEnHyWdy/HezFx2UOgCExUwLzaqnEEiyGezE
STQzAJUhAUCOJKF1BPXOMzPI52vmlOZIQlrzOX2887GTrGO3IhCPB9CYFX3mq0VjHJ4Co/bF+u1b
EcQD1H/ePbwgCkJGKA9im7woLb3bA6QQ1wgSnM+PXzxFwbJSUwW0NxioI/rBMJr884YUAw/M8FfL
3nkcXLK1Ka7M3QfY1w2XAPdiv9L3bOHjnJtkXW8PFfYZ0xon7uwOBWFMejXy0CTIqBn7ThnX5ylc
pdtriFgANTYbi4EYNnKdE9QhA7aVK4ma+iXaMNJX1PMRnzvkZhhcpViLzUEb2GvabwPozcKV5glf
WK9reOg7vTcbBYIAJVHZ/lxqo5lYDOPxEgC9k8E2eFSWl6BbEQRoBMG7QwFDbiCcoSU80qxnmKxm
79H2fHswDfojRJLSokGGgiJXKttySP9CKovOE0xR6bVDktJ5DEuwdvrzNdScrlTccjvwfq1FfDnZ
szGRYQgBT+MRZX05WtRMAdYSxhbiREEeXZRBopl2PbrWa/ZndIF075uCCMTeRJINqPqdoJWa+p6W
EqQqHCAPxItSI2ywdrixIvlpH2udXEhR0/oehlEvNESLbnZFFyX8rb0Uu9eVKLi+FJkNmT8SIGHJ
LwAMczbLtiTUIoBZnWqfQlokc1B9VeqRzY7Uha8ZaKoEP24KgzTkyTx2VzEsDyzfdha2EBbF7hOR
uPzxyzES8pt5P7tkCWyLaLpA3EtlHswh49z7QJTXfO+FcrWvlGanDG9XcW/MF+ZDiAL+5fAPIE+p
+LedGYj/Z6XDsZn9jw2mvdBYRY9P40rFVmZLn+pFN9cGhUwiN5DnQVX5qlST0RRF7xXo/0AEkfMZ
nVmI/gVWTusyPYvzuEG/JMKvQbPhzsdYA0txKmx0pn+kMusEdQ/PYsk9OhYWvsk5okOrrTGvbOeZ
9leBvcz+3BoseOP01rga6fDc3IBezBp3drruvVF5i4K2hy9gnD/MVqr+ni8HKNAt9GEA4knUI6eE
QIsvftu9QeXq5/85M7Bgco30+pRsdoh9onV4BD8O+/Nq7N96cNloGGYrBXR4bXTS083UUgf8YYLs
2m27DicU0Pj8bWq9GaqIKLn0JMefhnKiQpBge6QpDJ+iPc5wbhaMKDpq5IAHHQ76v5XVJclE5SCZ
EkhoWH0KRdS6WaAy0Y6sClvX+pVBu3RnWRBpGORY63RgdHt0JjBXt1BbdeQAeUzUvHtVgUtZnRfD
XEk3aSKutT0SSQPaJ+dJHkXNxdBomeoY/aWgn898wKgIuZVuHFBcxkeGw2St87JKNH83vETxtGET
L+PNntU9MLh77uFkyGWsICq/hGUOzD132FIVR9TxEcvLQd+abdetITpqropnu4RxgLhSOaL60q7k
pds5KdaGvEEgSJnGqkYGpcz2a+jxK2V8csgaj2UfKlQC1ShQx2UjY7wRozjZpf7+BibjlZiPQOtI
TnbKBm8r2oFeQHTLPbfXGCHQFTvP6wmtp5ApL8PAIEc1PSv3LP2LmVY0bH5kKoYKLFwW/LjyL/dw
n0oolPSBHtdq5Ket5QHaKCihRTbTrDtqHTvIBxiRnXePaWLVetYf4b5OGBLgk1Jk77c42j1Wjpl0
yeXzyTp2Fpt8NAiaiDtnSg43+UCeSJPzfPR+wWNnumIYLD7pXXBV+aSnDKnFWeChC2z7v8kcX9Sj
RUcC5x6WZJDTCHOCGglbDTtzvYtKLfFr0xov42beQRoeeLU2HT7Uv4R+7ZUYC0WBaQ38mkL0Qaiq
8D6ehK6DlXU2JfvBg9UkmfL0wzrqdeDdRNO+bmkzLmZDZ+wJlLRvjisThGoEaUkN7pCoYn0vYA6n
EE/ITCsB7HWLinPNebkR1Zki1AxARMnOl+BG6bxz6z4GkfiI3EIReyqyaLO6V7pdIwc3SMpmpO1l
chqF2RFtkX4UPcWSuzGbclTP877u0KR+fC3uifA2f9dk5bTU8wST96OrDmbmPYYX+K1hNAsO6dH2
aDnpoz9iOFETktDY58wU0xx/0ZBUMpslQDgCfPtJgXjnMB+USc75EcUdCZ8WICjBLN8Sc7eLpxdd
fNpM/zkjx+r0qLaHneyIMv7L1HkOui7P6uYb7deV86c1/jboJQAEWwhs8u9Xq3zfNU1Pcl1IW5Hy
IWe9Y+0DjArF6h80H/DDIDfZvMaC5CSjLA9fJRxQIq5pHNE+CpI0Z0dk1fhn3y5N5xQ3nn0Usgy0
bpvnwX10tgsF/BV2ZFapnGnmZYaiQUHMalkTtHVTXBs5NNhnrODWAX1n+y8KUnU2Fw7bnd3dQ5BD
kg0oiCiPfXilsMirj1DeG3fvlHYJEbFFg9KzV4I6VXdlF13rarBC0bUV4lYBfolD2OGmACeJ2Teq
pAeRMrqgQF0CiPJ23Avg3nffVKGWcSxIjs7uJkcQhpIxl5EFsOk3y4QrElV6fsqMKbA6JyoTW1l+
9BDBod+bwhgsDDZscRfRZJbZUxXYzmksvZt5+BYUQt5gjmvKFZEzdW3FSIAGdVbWDwQAS/3NsDJB
keBQJLZWocbiKlSjzlGg9ZM9wD26JeDPNJQ3pM7Bo7tD3/0agtbZpWQFBHw3i2rUI47YmIK+9PC0
bQr/wuApEJa9KjyYJzXjUMrgGPmD9OUb2nVtpIF5SUru3NgU2VIuDGgLKG2b3cefMNuFQHVMTTRj
ML7Cn1V5xY0ts7yfCdj3q/TUca6CCYlsihRZy2bDzsaUsq7tGghfoAsDCwUfPLhSEbYs816lA2Pk
f8F4+KFr7b9rXmqp96N1UOdV73AqkcQ2yQ52i2o6UnozKVxI0Pt/MyHKY2nLP6SBq332toLjigb0
vWCzbvymFEDBwk1uHcCeB4XgLwsb+BTlw0e8eUfbDaL5CVLVn8taRbGLkmjoheneSU1U4tPkRQqw
n+V8K+6kK4YW7tV8PvuJux5lNtJ9xCFekXhSaO2lo1+5hqDaikQ3J2yBqrFPto7X1/OsCoXw5poK
3ww7Fv0J9QTHpCw7Jllxoqpb0VgX+4tGdPchDRmUvLMFrrXZp7DhORwtlZsv5ZAjzV8s06wHvjWE
VKvh4ydHehXLUPaVEgRKToyKpuyXdV4+1DuIuvJVHxeFquz/bnCMLv56PcH03LEWUlVY7Wao18yQ
Xy4GSIEsu+eVAFZUZZu2pSrY6t/ab+vstwJBU9OIVMZZ2IQ6Gwx4bY30GItPsnKv+XcYs1OmtxBa
E6OEwQqf2mf8uUDzAHv20MNKNIY3QGvzWLHP8APJCvr2YEVAGBMxd1GajjbZrKUYDIyDF6KXVUCY
KoHCquw9Z1fuy486XczP/EagJNSYo51PmrBOnjYW/uHILT8+5uqvxtVM9Dfg+mXeV4re8GbIbn/K
hG6/6cYhaoNzKNx+54Z1Z6Vl3CQABuEzYvu+UFpC1fl7UX2BpTD8E6R43//+knUuXtb/XSzkfIrz
Xmygt9/vZSjilrfloLNCnFFYp2SP1T5IdCfY+e/53xnz4byG4UKLRUtYefTwASR+dYMECRtfxEul
VxRWPkPY5sJ7YaWX2znpWk14/jCzGpD5/laTtFqh3gzdvXuLfEUSbv4XKqPReqOOlcRW+li+zXSw
9+DjtYel+SrPpHn8CHPMcfpcE6/XWBBjVQ45eoFBoupQO5PCrEvvZ2JSm4wxDCknNlo7I0XLBsuO
pxyCxUAQliTtno1VevXopZccz4s+CHOXT791na5L/I08BS2uXAjOGBJWhp2yd0azkC6K2a9I0iJ/
dv0J2Ye1KtUsITHZHkf0bNScZJUIFy1ipvBNdNp53Pu6XkTBAQCbVAjUxgYTYJXISZUPQ0fmR4mT
Fwq/rooSxnXR0vqwKl3M/VWfrf8X7nMIaHIZqo/v8NV7/JPchaWe9/6uVpVdd4jzFqMzs7ym3e2L
n3RK/f07iZpdaqIaqCilRxQiOyIr855/FP6KSx2s6g13ryxxqg2afQnt5BVdk8Il7AV0L0kqdnll
pRQZ7yzzkt8earUmPJnLexDtB0ihdkwb6V4QQh/a04P7y/KT5KBZTvJd5ltNqKliCXybROlr3Dbt
G5tChUgs82/pvqfjrsuwd4wwstIXK1BXvfH4kDXf7Mu2d1QcsnRFncwFv0/mKnWsKmalO4fgtcjG
4RquQ+8Z/iYrA8MVKrcmy8qLqopvzDn7Kw4sOn6Pph4UqB5VEnqrLOdZrK0Ml6rPrCDPxKnJO+3R
e14pEGNb+vQWG5iLdGqPAnvyB7GMol1qyRPCC80M75KV9FbV7Jol9KVX3Px42eDjDBPHT+qxd58S
AR0iAwVPbx8bIoRbh+40qDsugrdxjlUorms5JFCV6FEMUHVBJZLNW28nO/Vd50g8+h/USnkPEdUL
RovcOIa2X2yUOtpYkOr1Im/6BjWaV5Bq3elqVRV37Wi7ahQBVySfv3ituljtWc8lQ/TOKpssHQTh
ho3Sa+9oDJ4OwrXkNm2xNlMZXbPwk1prJv3CvzELqksqDz4/DDIgUskpDjrgkWkFH6Ui/8kWFvnq
RQFvELxNUTedaF6fhwSNX0Mt7ySDbkBOBdYbL2lIN8HJiRsdi7nq/cwb0O+4lg7K8p2e1tQW4tEP
KLKTOcfv4xbb/yqoJxIrX/kcf2d3jF+WFI+v73CffZ6uajhUY/6mlQZ4MLHBnmVnkIjx3tDbo6VA
+idZT/v7OpToA9lr7Zc8ZpwM6kvHv03jtYUzYdGCz06HmF62L0MHb9pC6xDzZ2OZgSRNpBPY+Ajp
bOdFN4uXwiYJ/lLx8HB9aYA0qRG4tIjmafO0Cn91xw8INNsxZSfJndctKgYo4MHxewXezPdSHCFh
Yymti1q2+Ui0MnlR9aqfSCBauQEh85CtfyPWgMYBbFFRCyADuxtjoUwg7LbraaGZH+PNB3oa/0Ak
VMgGZmA3pnvHcJVvlHo6XkP9OBwtfbew3y8SoxJW5akhAldX5HvnjtGW3+henr5YLJbBDXCqwfDq
MrnmQ5SD/eLALTz1TAVxZSvNuPEh9XxzQHokYpadxGalDE5Y4N+NWFl36LYHZIaeUXbO9QwABAvB
TTVJRtEtgYDVEGfHBKPkZ0+8ozOB5wFn/ZILv55GbcFb42L9ntCA9Yp4r3jbRGrZvERGJsHS4wOG
BsNfbQdOEPUbb6sZB8rTKc1AGLMExlXjbko9YTzSHQ2gDV7pqsY+CUop/ZD0+oEVKks27wFLyfWW
WeLoJzjlTAzIQPs4Wl+PaOrDkNVJwsvd0GPW4KIdAMd9xJxjnAVP1fFsGf+EfhlfKbsOpzLEcohD
KhhZZA1bfW04gVQZbfPvwA7Hq827JUZiRwQDo0Mcb2yxlZOPs8xlPxwCNMK2v35cGAxLuxo0gBDk
5lApooa8cVFkq4tw4zRP+9GGe3NfV6jWF0ERMvAeX9zBQCk1AM3eLcCXbrpPRH7bOPG2LZD1eSOf
tHUrmK7HHiM0PqvuqfYOE0IYhbHGZqAJyaCj4o7edALumNNT1STEvbHGo9tEW+v3OtCYyY2E/Sz6
XNYP5POXTo/3bL7rTMc20TL1Q9OoxODVKvhcybzebb18jHD9yDW32545RmcLXWaK55zgwtGxyvKv
5WwHqOZaT+ZZfb00zhPZeBiZZjGeHpzJpAaVWXCgqzvalB7upIJUj/sj9udJ210QuMVc7+acWjmY
4X61/V8qLjMGCS5Yl1jA7O2uKCmykcqRewcb7sLwDf9qPKJSEXx0BkT3Yg34RoPE5baI1gelQpFz
V20zYS26ET8ZLUFhq06jzcMnFlO8zvywEjzPPCGI/hvebvv5jqJ7IZPPN8e35GxLZE+I9N/3POyv
WNdn0M1hVnOvx4Qa98j9ETXUHsl8v4lByGHkZX+uABIpd1in7acQj67u2O/Y2FUgQn8ij5raE2+0
aQRqZJSvjag40PHCiPkbtH6/Y66DOsRnQ0movpeIJW/5481R4Ae/HnIlHFsUNrsbUZdQnb9RjjrS
xJdVv07bXwJxNYjrS7chqXNocmkt9hvgXCYdNdWhzw0IZB/LH5jozjRUogI89HTOR4U31iyzNbcj
5IqvHCSzfoEpTtxJ3+qXGznionZE/Vav4boOMgIhFDkfFZt9QZ3HrNOuVOrsIbYL4pKOpnb+mhSP
F1wx5ZmhCO0MMFeYrmlocJcgj870Xjz3Ssv6IoZLg8O+360s9Ez+I2CWpPQSUWz/IVeGdfdl16oY
Y2r9royy/6Z2eBPaKgPT6rdnwl0G//tJ8LtHqTroLZJhUupwME4vpVQwTSXlkOGpiPsfFPCckN/g
MFE65Fviyk/dv6tAKPZlA/PZ6Nf3Bq7FRWd1UWyWWlV88gBp0PtnadZ2vCo4TAvCoSzx69ECXTU1
GTdAGGyniTFz5KZEEnQvaDqgfqqxHUGZG3ZQUdKefhuZHJ0jGQpd62b34aMAiQbldqGbSsuAyuvs
OB8MzpU9WXlLkE0wrmERxhbkhLmx5X43ygFJenmZ2ue1UcBc94+mFHv7vh3PjFLQeROKHrnf5/Bm
jzmIaBn33STpC2lhFvhbHFHlko65zKaPtm72toOAvib593PkKOMFmclqdxehA+Q01KmPWc1SR4rt
pAyiOOLk60Nz4Y0z//nuIJn43I59ddsMYdLKjUVnH6LUVjDRKjUi4CZQ1n3CY44R8Ba+L1/Y8DBY
HwxKAuK86l3y7noz3Lf56jKUblsrcD84ZIqDKMBBOudLY29WLLCN5O/aHNm6rac1KAKiTXhCbEnV
+diYqmR6NmiJ2fyLZvBX7I/kQpumrf0rza+O9wlgUvS6AaxPkNPgNL8HvaI0U/L3PVboU6U//pEA
snnGEuiDKJm5u8h1lKEobOPfq/sizTHCAKzsGu7VGr6Pyo0YozJkym3kzz7yeiGnpnvfgTiIxyU2
65Zz0JBM0g84+qUY6vYsZUcZSxeXfbu5JIIe3rFVFqwd+i0d7heLAX5gLdlBpIMeoSkiLVr+3Kla
2ygSBmjyy70azCLuXKaR4O32+9vp4GERiGzyzptzD8WNoWVxYKOQcd42secvPW0dBXvuvU3KYT6Z
TLOQG90eaxozhE7rF50Vatv+dXULlOlqSTb4294ZUDy2PLWYvyP0Fh1ZPu2Zlg2uInzIWJwbN38u
LE3T5DNWt1Ms+CS1dV3sNAYuqc+8VmNu6rhWH0XRj6vlqgsDrlTth5c/iQmnWf2IfzIMq+W/F6UF
3swPwEDlWdFbqInm4tubtzOEzv78+4Wsxx5YKbNypJGuXtZApeKtA8ZANuVyw1GdT1OcNwBWewpR
lk7Ajo1Ybt/T7nvdavJR/dt73RAKE/W/VpghJn0QFv0gTRrxyx6WNFaN2kYbPnLNRHirdafxgnYz
Ph2XVpZ1swjYmWJoUr2EZyNXSx2GJBeWMnyy+GGwVtrdL37hMuderOmGZId5YQ/sXbeSsi/28RA0
FN+ASbCgDAItjc7VDqG+a5T1vOyPYw3iRyh9QUEeugTk9WEzYh7gj0qfz82HCYfau3w5igRjief6
m8DZ8YT0s1N5aKnl20XVIzfH67vHBNVdDH3JSmll32dJPqreM8RmAxzrRZ1NeWlAMow/6Fv6JjX8
dyiXTnMf7EPy14bh3AZDvPKdO0KnO+mxXYHBeipEl1MuGnNJD2Ajldq9TOPOgk1tarutPBadnHtr
n5ZftdkyGhTjJPW6ZsHPPxdNWyez49pLYbOtrXzjfRg42g4hlP5Hdd/MkjPT6AUQ2Rn5u5qg31Sd
v7FRH4QNhqHTZYlYaqZUzyrJYIUCwDUzo1j7DP/GcpG8jxJ2RgUi8+NHgc1IREmPgY0wNOoTNmso
DNTIEtVUtx6Q5d94OFDzComau+xKb9dA6XreKv49xwnZJTMJTEXRh14FlNGQNv03h6Sgx639zAah
bDEE0IWx87GZNTermYsVbGywzG/LkZfrAU82BQASAOq6yM3IieIOW59vMs3kGCtqG81S1DycHgVf
Gf2UkTqEBt5QXoIfajGn8J1gaekClh+Ea9n4Kuh1T64w5Th55qDgbxc8rK6n5e7pRxBUNIEUSHCO
Lrr0niNUwMuL3+Ef1nABYczb5X0OR7h8lPzGEYQvA+wMo0/JhFaTcMiq+x7ucxnTfNo73LuJmJ23
LprA0QWSDcONCFHCHaT9+qDe4jkm9MYorOwse6GZBMtNZp64pahJH4d5rpYUkSLJuMY2yUdd6d9X
/lRRga4bphJLXxSnd3QMGD5YvNriU0JDwVi5c2P3fr1jjjwsNhMZIob6H26c0Y0w/6Av1ETFFiEd
8Pk005YeacO/T4szIj+26VIFlEfv+Q8MkTE9TrK4OWU4B6vwOP/QjISS8o43/e1S0gL+Qf369S+i
OzGLHltn1OVhDVjiKYGxegcdy9neLvNgI0k2FIa0H5oc+tfupZT7LE4w3VQRIXMmyTRn38bB9XT3
mqgBfyD1fgTSrSnzZfpbmwUYXVFUHZmLFf3YhcMIWeyFe1gUZqK++sgUqqAWZZYJV5mC8RvX480J
Ei8aUYQGZqlJuPh+UzjGmLueSNCdLG/pMqflOalS2iRsywCWrhrPwOWsGKnNDLueKBlLMhoojB1J
cudQFTNhXrFyCdEoKL1Z/MI68+0OZ79wBgt6ghJGz3aiDPptZrJZvhpKJopNhUWlWE9Qu+OXleq8
oBfi8tmz4GhWSjXZBUPz0QD+Xmx8PECjuBX8zv+JAwLAwLax07zGg89Nb0Xx+22jIhjYTkRomjQD
eI+8Ns9ZP+KhmFEv7XMSPtxIjAyVP9ofz80ZpH/GYQWaXKNySFnc8xPYVPQY6pC1IutH9E8yTcbb
twTbKWybVAfl3URpJdZ3lVlaQ3x6TiknvBbwZ/wgmNV+g/UMQByED12lPWFWzQJLwflhdNyvXRKW
2LQbfOuRafP8TFY6vcqA9Esk8rbQvtr8zMA4Yd6SIGRIOYtxJFrhpQaqmVOHJfOmS1Ek9qedP/qG
CTiKTQoWXfVtwqHxkZ1EWWdWBZuP9RUWy+aSqFjs+NgFr8qfzR/zZPDG3V7EPkbRV3AjwhL/J4uB
Zras3vsIqi/ZImKJhqxN/8LXegnDSUMIp4I8lDTo+sRZOHQLebgpiltYCFJ8uX5pjwpNoGgz9yif
D//FB55bRr75iNMIKeNidjdOyOnMI44bHWT0hKLRBnzsxOZBztKOgejz1iLP7qlJQAAvg5LdM5B4
X0URwtwmE9TwHAFgELfuN3qqwIrezEd96NRr106ldLoZ5uI1WVrZQYgj2UultauRaFBrzG8w8lJc
EEOUCbCg2HHNcpcOutweCJDCuNfYT0+qtyPKi1xqtp2sXL8A6VMomPRBqyqP7L3qRr7HIwAVPEgJ
ehbn/9wQKPdzIO9Dq/sNrKuzw1ZSwTgy3d6CM8MafbcVnhQPVd3gIWHdjjFpKTsKQUZVYfKO6U4S
CnoRZg4BncZvUQP3/+FbA3gJhuquhlynXquFfx7pIBBdxDrVOYlebi2OH6Eh3kGyDlre3mF4M/4i
JKNqW8CrY+C5eSbgchqbaRgHtY8yiKLswEfxwsWSP21QVQnppq6kEH88YuIqwmvwn1bTWf6boYCB
B/rRn++hkR7KcVZvJeY+5gPkM9J9WfiDfD7b2f3O+D0jdmWjcXIVG3S/D7NNZN1gvup/W946PABJ
POrfQUnYnZYgPhu3UF1JuJ5RFo3aEYBdYpyLloyqGGxAAPYuafWDNBLQwzee+nFJ9AozdlHZ2CAC
AshVPz6sTigY9OX7NvrqAczifGiEPJv0cZul3xVG4nTCVEHKBZIWuXJ6pq7tP5b+spODaW0HfKkm
F4TQYGGiO1nGZCBsYs49BJ563JVEFL40ILKmwuqXs08nkDk1BqLXu+q4E5PTGHb09uugSDk8L0il
74cLDgDDXdhHvTbzwqM1TnmwG9tjKyJXfEmeJuDgQYhWFlaGoA1Llicnawc/74hO99RmOWMf8e/d
Do7MOVY8B0Obwte06rcRwLNvqkwGtLeEPC9XnLZc/TUde1jzt0821X+571Lf6/oawc1vwkM0Yqw6
XRvVf7eQpOOKLliP4tgnzAUuRm3Aa1MsU/309vEO25BBb+oRZNz7vLm/tywP3+FoINMtsrkRSroz
vhOdP7jOIpZaaVV5pfumoJxl+rvlvdYZhqmP4xT2PA5mBOE7+mw1D/xSdag8lzk8Q2lNFKudaGx7
U0ZpAGdrVK2mRWnGzjV39m7x3l0AqCl0Ayt3mc/lGYGb7mHhBdqPIQOtzxnqyrVio1PwsgRYK1Sz
jpo1p/vYlT9j8+7VuS5EFAt6T9XiPgnJc1chJgLooaAsf6XArGmOkAeUnriUpVLmhgZUjHcYGdfe
taAy7rS8RkcGjeglvZThI+WJZ0/SmumvilCwqvTOX08qJLTcQrDxvto/XjTCvoG8mZnLsYNDxDJD
QOTmVw9ihoBSvCxVs1zhZ87CMV99teCDw/Kp8DAXtRuqGmX2mWCPM9qtHSRzXFRFATDEoFEHdxY5
wkQDwn2zzPoyL5hBb0kGiQv36OqsLbUlCvvMcU9dZGJIOChIwujp+zbnU+fCNoyQT52qSfVFI5S1
CXihFsbnOZifu0H5sf/EXAbgZvQYdPh7FfdG0CwbVPR/0fDLctdDDPPYA0FZOxg70J+BA7aVIsVK
0uwoUf3d9PXdIlJmVPM1ZME1ObHNPR/JkcI0L78mVbwXwvPkxAIHPdyFst77MbjKkGx7vkWC0fEA
rTxN9QNFQJAidbowwaymG4hl6rdwU8NRmbjWahWtlhiIjMTCn3vN8dp5o2zKZKcocqtD5frize6K
Fkijyt8HN3a+l5pIaAnKxF9uIuikfgKKCxOYC5bTg6eC+P9URteH/Z2XmJJ8WEwZR++xMNw5rdQb
Wmo0HpXQ/jNJdcVyCZYxUf38NAP2AKe9FYX1O9a7j4UrvTTmj0uoWW0vT0c723L09aI0QNKrZpt+
pTHGGcKjaK7EZ1yPJyrMSB/OdfCuPFRbrP1zX7Mj0HQv2xU0NV3/q5RL8j4WuztjFWq/iOnUtSI4
bS5Y2/uOdMZOa0DnBqpmyatW/JPsO7ysIXzi78Am8guVPLIPrJa6JqcYjayzgrQYDnvaPn4r4hHg
RSUaO+ugZkIzxl+ZiordCo+i+lKUSQhmsisj0HcdaCS5ThQw/V2/TsiKLEZbNvZAcNh6bdx+BMDR
/FWMMR8NOI7i5Q/k2iW3SpWZwbTf64+zo5OHoqvi5cVg6/0zKdxAsEZrOffCsFpJHnCVtXdu1cW7
KyTHIDSASgOk14OAlsPU2QvC053ik+h01ARs2U64VVtL1H7jwZnTdN4NSJoi+IwU7fj8wkBc/H+O
wGA+ENlpCYZHEG/WuRa/9+LAN1lBFacevaqKBrhaU193RKsEu2HdBn0dH8Jcy6yQL5xRqJe3gVA8
eDq0HsXDkUyloJAPpFKrNOSic9hYJPxwVWYB+m6nYMekfj4nZmCBG70HEIj6yAjwhWDCnbTRsJz0
rY7qoD8ft3f3uNi+zs88haE3Ua1SUPiiA7r42xgM+DLot0dUbb9Ck0R1Rpm1TnWrYdzEG2CgMDAM
JStCCNNiDapokW0AS6w5HZkw8FTahCCyteZavkD7C/bkcmBGaJnE+Ivs2QGT2kiaLQtmhxuPdHch
TMVFbccQTDqu8fnJnuutioyAJBeUKZPd/9+ynrFB3jxd0H09CUS2+BXzPhRdmBPDn6LGGtycO8NO
GmfC3YKS8iX5WkziPFRauLgoy00ZlG3MFSKUzGUXl9X1KJ9qqZDrUbgSuatfq7daZnFQZyasnxe4
wD/sY9bCY/aBBITKh9A9dJE4X3FEapAu9oOEu+/sI/8D+km6vXmzhxSYBc1s8dOB8ZnzRMvkAkV7
WuXOd1HoWssQDo75M/jXbH00CaA9iz4KgDi2EFemB1GICJxvdpQ5e0dNaFFI8oK2EJig13Ow2/lr
TmoBVMvZe0pcDMhSV7WaAheUw65tlCIkUKks1ovyChYrP3Xqa/V6UU3J2ZPTUfctOgjO3jIBoIJY
y938qVn6DBoMVkQZd4FzF9aEI6qXyon30rflFQyWSMZOTTzCEwHpTLImMSWJBBVGDUE2YTh3eVNK
iaHz7vsmmcLnU24YOVTGtL/y18zJj6Nzlcj7ZcWaI9otx4XSKQQAuzWby5DkVTC28d3CmeTw2j34
m7eXhGshHzi2gIY7jeMRWnNYSW6Yht9kn6KUc5wLauuX/hUc0KV80pTtjnrk0/Ismj7Cl4n9Vngf
zTmqVjkU8gDCi/bQAgKJWrLJJyAOEfJqpaEvoCnUlQBx6OuTsiHDx44p+QwZzrH6BFA8tql2xFUD
mGZwhXROyx0Ic3ha2Vyfh9AH26CFDOyiyaKx8OJnF+xcxH6Zxm4Lk7anJjpzhRKUFooUw2H5vJHi
GDBT2qszHknowrCRNxC1GhE3LFLwiCl+iDDye04FQXw5szuNQmK+hkIWKakPWk5HAZYNBTBWkBfT
0PLpYw1Y2cYNKFEzTXrqRONFcO6piAEupLV4ewZb9JPx2rB7K1U/0Cf77vU+1f/6Xhm/aPzqVnRh
xe4xFJuwG+0nMkeb6q/pBuqlK+nofO/mU9ZA6hunbXid8Pk92tcNquFw5Ke8NZ+EKxZU5ozj4RnZ
9DylhVU3UoPHFo6DmhCtWXXXEPFmR2pSIvrzB9UdvE/PXJ4/Pj/3z9vl+dsgvuAzQ//+jRcsgus5
pm8r4iLvIs4LMkI59gx+QoK9Im1Om+yE3zALKcj/FGX8rNQJO46vWzh6CmqI/xw6DzWQfGzHoWKk
9m8mmPdHY8XIi0qLU3AUv2atnrozqjzmKvlDMACKbVl5UqSGk5pZf5faE5CODmdlOwMjqM8DQFQT
g45nHKyKsMWOaSKNcOMBShk50QtAI7Nn5Kx5gokqbItZpmKPvMoNHB7leE7zzlunu1d/5OlQvxsl
6EUMQZgrFZDGap0AhlZWQSn87fDvcYMzxk3hhLI6A7Oyc9JQdnVwAAceSPtLToPu2xLPowfpSeZP
+01JiqpYfGdb70uX2+HXKrZTWfReUCLsQqu52Gyme6PDI/4Reb+9AUdYAzkYt//8Wm9QzpI930m/
FQbBB4oBVl2UYKMktAiWX64qbIDVrY4QWvOUg38HUXq7ioNrYZkyNZPZSw7ysIJs72Sjifav3eaH
M3bzP+Hd2QodpDK//NM+LyRbuvC0siTc30XGYM5atTTOVAVrHPcRp+T2qYn5pYYTS05cblsj/e3/
JYI+PQcGCNMJeFEFASH/x/c4UXjJfij+5g+X/2Dyc5BGki5caHQmHR5mPBlICeGKWoL2tpCHBvJn
BBOHml7fwSkKJ3qwALD5Xzi6cGeSWqdZZUP4+zEGfu7Pes5xSScCA328wvYhw3hi+OaFuJms5Yxr
wH9Iy+1Jv3pVX18ufO1cOB6rD6j/487CW23GA7ovo0p5p8OY070SsYC5O1zzsp9NfG2zLmHb76QP
+kmhvaUd4IDKYPpZBY+OrY0Na/dl3t5sBoiGI5IhOg4zYpzpByDpkdzU0uplaXx/hF753TJSXwK6
BqUj7/a1yXcNVofYAwcyvIiQFsmE5CkVbEf4+RKXpw2Hl6srIMQPV+qoRnJ+ErrMqOf9gzyBQyv5
0Qr4uz9qQoMCQqGXkSAR+6nlAG0Jjtk3lygDW9vHCHVnFP7zJ8UVs7kLOgToH85Sh51kACojT+U/
mjjubVW7jukcKsE/3gWV1Qg7FWaugAB/uAhaseMOBj8xsUuHqACqOm3zPnyvCENLqEZrvseLKXjL
dLPGqf4dQ6iMxjW3Mg38B5oLEiJalMLGG/VgQFcYoAMNwY2yS1N2dQyJ8nSGAWbWDyPW3KgFyw4a
J7suPy0lHD8IOt3mBcKqyx2Zt/G5J3hI94uaGyGlqwzyA3ryIn4eDIMc9TmNMXdaLspXfhfjt3IY
SVYc29v+T4kuD7NW4/RsO5n4uhyQssB0xUgjcGgcIPXLv65j397EjjXu5xJmiFZLpGapTw2c1dg5
fyruA2PcMJT7h5e+0Gb9Zhzc+wlIH0qhJleaIGQ9KgatsKqU7Y2OTNXkRMMkBPnPBI0oEq31Qp0U
RL5MdlzIiyGpJlMyD47EdRtD0XKaUXd9HqTF3u2efUNFYpJKtkC7vCtFfCKNcs0GOnTxQLn1tSkR
xgqtigCmwtdensh5sn2JExMrcCmBkhRR50ZFqvQgfBpYd4uXA85LCHyMCp/lmyMZ27aJv1u2Wi75
t9HibX4ceToyQZGbU4BdBWWYf2VfO4o4jgjqqn+A1qUFD+zxrckJkiokeXjl+HDKPhkY5LSrYVMC
dUAbGlUu6DhveyHWG5Rx6bxFMO7gX3JFhQbr8O+n+V11CITNsJMU2bSL4Zuc26OqOZvwpDhqrT3g
Aq3F1uSieb7aYP8QZptO7/DP1MKrMn4pnoFwd+Mjvg8zxzlr56WIPCJNHCwf8RsIR4jmJ8iZCS/Y
c2aN4xqgud+Yv3/bwyODx674BmFvfF1VffVLEUvVVe6DLyewvDcyC9pYVMPAwF54PLi+/vrCRafN
e/C/mIsGmi/NtNJSslMxtR0ti8VWCrDpoHQAn5HfacATBl/AovCj40ttkRRl0lDvf45yqYOhmduR
nu0jeunaxzYJ4KCIHibVyOzNtVbHccoXLU98GP6CiKYrdRf4lJfvI5FD53duk9lvo21rxTI8anku
XwkVEouDz5bIAZgDq89h5G1LyggP7pTdq0GRcOnLDaXHCYPbA9Wq4y4KYx1Ti9IxWlrHoCuoYpcx
LHzCWUZAaX8cpu+oDuj+Ta9civom6bweVu1xff4lAb0YaVrZgRWl/bWIAGVzKOHUO6CET12HskZx
eretVAUqzbbM5ZQwR7RwxHArfegm7BseM1orh3CIiBa0jZcC1V7mjUKFzjnuSWN1PN5cZZ+W3kcs
3I+VKS0nt5g3DilWZvfGfZv4vzvnsnmDsDVicMhPUSpL7fODcUN0o2G2WSnMzuTuPeNQcjZo4HwI
7QFB7h8RrCUn2G9tmPySul/sS5jpEBkJD8TVMZYyZhULg0zbOB73vFpordgA/MUWm897P7zpUOk8
N12lmbpAOBV2zaKohKycCvB3/iphYMrK6bRyKOsFTgDSLM6jvPzi+yr7KQxHInjz/IfB5oaQeMrX
rUR7mCLQbuUoDxS5s4gn6F3XorV0R0ru3NRPmp1D12Md7LBOnhIH5jJbN6Ao4UFrlrtE+a3xfQXp
RCZjHDn+bhi8IEukAtqrIXa5YPrtdKGtmiwlD4yzDKIZmuwIYb8Byx9ZM2vcB7DLIvqLQP6W5hYp
iQvuwQukSX8m0qp0vhFlkwLOiraN3kmNGLugacqkNjm7tVlY1/uTpXMLFGdPu0SBivDl7rBCrxXc
jr57da+KnpRsVWWJgm2l3FxuKmCkikoAiJ/rvHqjFz0UuWC//gfOpzPbEgDialWq4E/LyNGG0vYz
/esYVTIrxC/JZl+WNhxSuRmHOO9lsHm2G55MUkMFQEy2poQ07jGH6qmXEPXAEkJ2C/lnoeVLEaid
lv5X2pflsiJDIOZtFsNdwwYPXJeI8IdrAjVcpkXM0IBofslTyLWwhVbs5OWjkW8Ys7OIwNgg8DQ2
+O9bcePtNYkqNIy8Q/+/OO1lx5lTa0nFuUp1IJXuYaQfuIyJ/JVE/f0VtvVFxxXj+kAoOyw3eLTc
Z0ELQBmO5ylSHNHR57t69KgoxiEL1TNu4XQdFKMfvsaPmK+5XmzVhU8c9qzLnZsX8evoYYuNFmxe
9WgHotpPkYfPPdtxgPGgMmov4LFmLFGv/L/o1WxLN1Y1DrvMtaM3qsVJjYXbbTcowxFQgrQCDlXv
+1Qe2x2TTSBuo/+MrNJOAS7FMvwXvycu3ZKAYygo703sA/dyA5X0J5NjZ4qPm/6MESk7ZxJPAijt
bOlRtbA81sGBJQaoAtnnD+AwCB2iqymnHyrCfdQaVB/MRbuHbwwpkESObVjBymOtL53XvzXFSCMy
uE3VKzyNFIBeda9bajDY7L8XiDTxttcAc3aTvIAvJVIxBoP6rw57SJK17j9JDpGtrJjtLlomXgZX
GLyDgPLoahZhf0OR4Ve4KbPG7411KUEp6+bJMxdcQLCtqX7qV5C2wr5zaVijK1SUbXJFgzFKaYN8
RJucOf2o+RxK3+LTqc/oKwVxOAz7HnuIO8izpDKGOeIBnRlfAF5rWG9mKOOgnI4+NFQ8KtP7P9mN
GoxqUQa1OuaTlKDGU1mBa/fzJONQ9FvNbN6FQsrchOJA8mWAavj8C5WfymaxsGvQUeo48GrILRuG
ow1T2SvhjtN5l6eOyvt+6fvvQCUxj4zlVfkqmMrc6jMNjWwmEZfBheBV0Lp8kg9t4i5lBCXdB/OY
5vePgfPFbrY2Ke/DZFwSyUsTUBOSm9+9WX9S17ejajPjANDYAElH0QyWHJSbKFbjXDTE9cQTQx0T
FapJLiwMfNq2FuSWwvU6X8QZlVOF1d1upbm664xEseDjyrrHmq6KxOHJJ4Yn0zG+CJ80jwgg+8hB
AGMWMRZr369QUdxyuutVZdYGICTcwHgqBD0GxVNYHKzN/vSwFt1CveOJZA1sa7UYoWvshyq+LTlO
Usf6jqFOEsWEcIYcqH5RrIAEiSy8et7PxqVNxIJvnIx9DYQ1G6Hx/w5cXHtZtDdZwzCCYias/Hh5
o/yOQSbhjAFd+uWINXKeHFksGBPSSawXBzh+hnCnnMhICMoWmxzUNVgVPWFMVISvgQ/ww0jYHhzJ
0l+2Q9Wrk5VH5f21NY/vvn+2csguJVrZVlImCx8x5RsfCLQ1q982PCBn8A6hGp3UNX96FADs5tiV
xTHD7SVKiJeHmeuLt5P7kn31E40T8jK0//hOQiysC5CzUmAKfdgPiLrmNwd+jDF+7usSJwBJFrKp
DN9LgvhCrxHvksXg4qVhxoNJqbeNXkloVc2VgkERrlQpjwRMywf57aeHniIymS5Tt+V96osFQvu5
MfmVzPSNwjGqpvd62Shr8Bj/Z8RwhTfySyVQMt1tYHcJNYL2ZGszum1sxK8jRptkYW19BxpT0U/1
phSbDC1wOb4S4p494P+eN195O2+Px713cBnpphRczlLq8SQgn7+Msv5cDtUzFSIokBsuJhQEuV3r
rQx7zWiZEEFC7FJmtnfPnxFADfyMSnTsqD/ovl/Fn/7EDDbdm/WOC+6CTeu03MY9C9QpgIoo/dYF
TjdmqVWPl6KbWDaui8J/lRUrluLsBqUvB51fwC0rjAzdGK8xz22qdHxRpcuOF6q3W1XfQlbLr75O
aU9ir5YLAH+kv+v9bgijajk9Z1rFQYpOoD6HGE0STI9qM/wTfZj/SuCm12LpPG9L4lG2JNLJomaR
1i5rOZ371JQ1rrwxY20KdYq/Jy+KfTy64s72DUtaDnJ4vkEGDFG3lZqi/4AWiqWNxxXr7YIIMAC4
cKd7Klj5LAhcToJ+ZRE7mbarLlgvqb6O4T41gV58CoeZ5P2/9MkKJVIN/Pg6CC62OCc0/n2Lr7yf
31gfUHXLx/zOd+WGrZJXrQm/f1zT6HwX0WlRJnzHhGCcYyDIKnb3Be2HEhKcn4NR5l4rRFmOkyLP
L5C+9P1kYkYa4bihlU5DB8TxmicWiD57YuaWgdiYXfxJEpDoz1MtOVOIdUAgg55rNYpI7A94/miT
Ol3+bQv5N/EcIRUCJqO5Mgm7kR8RBNTH8hALk2ajYHL6wFJ1Ymv4ogwx5FCOyTqHQQ6gyad4Anh2
G1INQp64E9FAw4VQ0o3Bv4McpZEhQDpcAEdNsSqcj56HlgHwGoc5u3OtxX8R3yXXvHRbsLcY312D
fZ65pBhSQ3eZai3VyDF1/67uSZnxZ3fkYwKtQA7B2ehZtOvwZoaMTandyZ5evgmcDM+kKd34+7ql
br9Mp1Vrgxb90YXL/i6shU46nQxaxU6RlYhBQn8n5UQlA574fhnFjs0lYJZv6R59RHNkVZlajvle
O+8UR8W+umiKkyWlbjIRK+4AdXdZyI8Nj0diw6dQZdqjNPrTOI2GN0TrBFEv0PGbxOQ9DECDtJ01
MrAFC7Dd2Muh5D02cvFg0c+2fD0ogD9eiB21UAcz1yTC84FjxUSjARtgJ7irQ8ameVZN9Dzx7d8g
DvEXKVbu69Nd4cgE9HeTSuI2DuFRhRI44BHnlefE0mNcIkHLM2U+/YGMTMWHyRCRBBGjxSUbn0qC
wpGSV6wGTUu58+ZwAemHVKkfPdhRA1QZ7d0z0xgaEj+Hz1TZBooPW3isLmMLZvvXgzFdmSeivcrN
PcdlGoV8AaTln6GbmJN6hSV2tQxzwEll6WxOin7C3CuwpmDTSQMpqEftWQOMnURxj8BiqB9ALqpl
aweGuFlO/IDODJ8WescdzNtj86C6nQDpqV/305TCUtgIqrMLaOzCBB5EhUB/RZyShrIjEr3kdxoO
OUirDv6tEkOTFacpQViPv6UZLd0ltCCVNJ5+VUJYs0xIJvjkD4f/LScHeT/fw5AYNDbVmVPpF9qo
CkUXDzmAkby83BX4UewyWXk11e+w1ARBZzxTNoLsvCZPqldaRq1dXUAfPK/Tued9sjQrkYSuamph
KXvWF68xiCiomHo6k6pSimhvodjfm5Y+JNEDAAl1ha7AJlE3BW3BCEf/+6jqYWqHne50bnzlQWXD
4O2eUpcFKD3li76BzvQ9kD428CUHQmPJxy/gKkwJfCT6q9hxgwfZIFAuHCAeRK/g8ojAO7e0V0G/
dHEcH+dR57Z3SpjvJ5DKzbSZ6/FCpHOsKc9mtxS9QuuRreHjx2p6F6vfAPcx+6QU7MMCrorRjbD4
JNs3KCyfMEn15JGfMu7zlrZEUEpOlwuPkLVQ+JuxEj3aK4l0UgINVktQEwD4qNjUL89fxsZHuz+A
EUCt+f2Kca6W+SlAl0eGvTy70OS3R0K2aJh6BdFvaqF/fUkMTsYuk1mYdP5uGEi41cunBa6oqdyZ
kicx0577fjmzCEpndrcompLp/jolWg7qwaJftMnYIct0rfFWkb6mMOqFYTka4iSd+lKFdL2rdQ2i
MuskKGYiUj8gc5CAA8pMP+uMdFrPxQLM82iVBs3dbiuVHklPA7b8h6dPQU4E/GudaGyhzv4xpqlj
qMGdm7EuasA9bLVeSFKROtLxnYYAYX2/DY5bW3mwJNuSvG/X+Ro4ZIrvpNc8TYUzxdtysFxZYFxa
jzLp5YAkQ5363im1tu7cSuvOjgbX7jmFqdYOxfKSxjrbDpJvEsPy19UZxbhqAJd2QGejNpoHlKbY
wVdcg+U77enHK19VPC/PpQL6R3TisHd4t970HRNYTiWZPqVL+xB82gMFSafDNeo+KhaKUFnPQzjr
qqM/BydcJyvRInJbCuYtpCOTfF7ZVQkDbksU4xUbhBROcT2Q3KhF3Baa+oqlgyBUd0RDhorFsFbO
BE2dm7PQ4cXLzcdFPhxAqD76fIj3BxArf9wDHA8OsurxWfzLhPEkMzo1IlP/ZmWdASrsrGy3r0Xp
0lrKVrM958Jz9rR12lftkyjdUGHCgze6kRW68puPoDqYBOHNsKNQs2FMpG0VTijzZEBwaa8ilFqM
yWzEjWz71lHfqEYP1I41i5RmQxWhnzHZ2/av8gJPii0se2bgcAresFgRIZ8yFRICJmQ8HgYAp8M3
Clsj9RmKeGMNXWm2vHKuL2HNOV53kI+Xlw+3DP7doyvsf3VaQVheYJaf0Ou1o4tjuXDXOL1QY/pn
d4OyILXvHBqEaq74BjVc8QklqOJ4d5lfNpMe6kYmBdCZvcnTkvRn12Br8SJCDwAL5LoclLGCLdwR
24kgPraRdzQNtKyqlmnag3KcudxVbEGXLsWdGD0SCaJi4VLdzKNLNr6k5+yHUVFZY5ThYEkfxNZg
+d/TaB6zFEWGI4RkPcHdVutVx3p16OxH7WS1dhn94mA5E7k9czGAjW6u2x3yWXuOYL98h6ge0GjD
K27i15IagXnugjpyHYIHYUKZGyFzJvuRi5nnI1CZdl/pyHBBy1khTx0BB6/Qrc0paXTB1P4uSL6c
3TI7UBrHbXEAaOHfhnzrX7cD1MfqIUFCNAmYPPaNSkyYAj7nfszJ1441JeigG7zhMyFv1NnWMDrH
XSdUdB++ZTSQQq42y8EHtCM4FaIUNJqRA0GWrOs0lY0VZlAdDfwNNr2DWAD92jEslWSawLIlrhLq
qizwqoKhtXs9XgVgPwf2EdkzYX8w59JhIsfUpWsFyMulsVR8g3k1Uq5TuHm6SNZ3CeHs864rhxY7
VN2ZBb4tSHVLZ1r3oHKDUDjcs2qtt08LzlVvaUKxvOe+M6ZQPuK33z0KWHX1xM7VH1QZ9Q6RXCAv
4se8Xj95Bf2OtWbOqAH40MERacXDJXPOS9erLmxg5yP+/ULVtiGiKkYAFnVLzjRFq4TPqwBmCXJ3
sNgGr4p6cWAxVTWxaBd1bPdZ2CZLJji3lzQOok77SwiSB1FLbJ4nBopRoet7e72/Su2wfE9bVjzu
Uc/yBheymtr6R1JrOwBsAhmEwd+GhG2nu/+dXRNA5JklWcK79e+thRS3FtimC6c+H5IIKYO8Ei3w
s5Nv9FDFiLAPcIMapt9aC3HocgGrtCOn/GYisX3pb97rOLMMs4utNv1p1MknCQa5i2S76Pf/x70Z
IoX9gxqENr+Ax7lHezOXSYZIFWwe6KzBAKGE8c/GBmrj8LMe70ZVOm4bxtFHp1YvNl1t6qCy/roW
0HD3z71V6AB76JO9l/OysnP8EzytbUrPbiNdWUV985U2XREr5W9XjPSLfnh2SNGyeeMZFYegIZN7
9obEvaMKa+voLODdRjBOzfLx9oEJtcbTH2tS96AzkuLC5cTUqX1jQB9eynpsNDrvWknQtX7Rvtne
My16tm7q0AekYmsC+AgZWM0+aHJcB5/YxdnSX/Dew8agWuj3NgDBU2ZFSYVSjmV/m9+mw5BZL41c
qo4BM1tg9q+RU/XYQbPq98ICcRNokEZvk1D1jNMym83Can4btYmxaJ+96vbdaiejFTgB14BL861m
YkqMT/kwsxjEH4eF1/zPnH2dXyb7uZgXmQ9VT/UU6Q7ey2f2sfp0DOPsm2W3EezeqFAHZARhMQD0
OWNzHOJlHglX5awJncXqgVIFDSQjm1++86jxqqgmYbwRvzKG3CSO1FJXM4tExs08tp2i5ML1jKdd
rU2m4q4Kmcakk/p0qML8KI1EJyuXrMHrEC2bloNdOgOAzn451gFSd9imxIN3wb0+hgkGrfXplkoc
+7YK0ahz/FpIQtiypFn/gz7LNvtXcsX2I0mUeXRGkGLLL3fbOGROkPuyG5Wva7et2gpdRzPY+qkj
+31dobFrOOVqzMcwWD2G8To9mOPhwVXxBr9Hb9QxMRS0Y34vAguOr3ScjdyFhB9F35nUUP0Q1ef1
us+d93EAfgZWg3a1iBtFbL46QAVq65eu0ILG9foUMMLvFrn/k8+qiaxzQ5PkW/1qDapvT54rtcV/
//F+70r5SisYM5Xqt8NTAGrjiLgeBnSEK9btlqjV5/VkDDZ2DUIfTHMhozGBt6zqpp/lBOmP+SAd
ZqYdkFu7UiuhmN1vjTR+2o4QHL0SCWn1th0/UZfP78C6Ot0v8O36jhSRO9jr9sAr2ME/SDWP4oaT
ZlYNwzn7zu3EEwC54RRMCqX1ol6fxvwVR70Oexg+ijJLJNckofE83y3RbZ8LB9GJqW5t4tg25T/6
nmHriTUnIrPPrpyMY2zrAXpV2Fj1d8x6UpfhZtygF6ikVDAy8chvy9koogTpdDwT5Du5kMvtb1II
gZXxt9MZBNXKWIb21AadH+M/pSnxy6NhGuFNBtzrV+/3q8pfVkCOqgBijcsmvzcEEMxc8kBoEbZj
3/7QPkuY09YMzEudMINEaRXnIJk+cqnYU9/boRwHTFP8Px4AOQuYMacrF1+dqp9awZgp1GeVkftf
FVuIhN/2UFFFdGtmCGeV8WsIQC87dNhfVjCKb0/XgGvERTWWxDlVggNz7cCOETbPAlkNCFy37bBU
qfsOa+8+ReuhTDyoWxhfb3cJx34zvTTgHFYeEII9cOQgVUBE1HOSiLMiW0NHVOUBgmz+hjIp+urY
qzaBj3VyFgzBhcoU64bjuL8OfDJlwsiWMGS11KCRj2rJfDcNdMO6ILLBpeIa7dsD2z33KMbrwLeh
aShfKh8ntPOR2HzbVykWimWyVrSU3NnUoW8xYjmiIFyFPFUAxZqY3i6MqaF1VVGxh3ibQthv09d8
KxBTr2JeKwltij4VyNA1OHzOUClZI1FEfGH5wHMddYFM4md7+HgOMZgiKuzGOW4gBL6CkLxrwS/M
3isHX9MsccmYs++CX70hwjKnfhvoI2hlaVN9q41VUdfcBy15WlCrG/5hS1MkUmg0r/rENgMd2vJG
pRke6Xj7QVrRY1w9MTb2CP5TSOK6Eelm4HcUxHNbzDipF3jqQfBcsh8xJD1V0Xk8m5duB6gSMBAp
24sGbwfyy4BTd7Uww1AohTJUNy8WXHS5YWce+D4n9HpHMrkgWgXonl4APQQ4gmZjGyeVaW0kJG0Q
eIgwYPm6XCrOVrAzZ6+rEhNH+EWmtBevtLtIMtxCul2HcgO2HNa/So+oADAyJI/3TxxBTqrNzl/U
ZmXp+spDFXRvqM2VmINvKnG9Mg2NtdtkbU2tILs2YKXwGawct0ABChEO0B8GABFObkcwUsFWQBDo
KwQzhPFMVH8poZqY2j0heS1UB+5nCL2vrAfBupnZiC3UJnWr5QsZS3kqeGyDri/+c6n1zyEXJ6BS
Ag4x8nW6Qe7iCpgkLSXW5e27eP5CC4jSgbMc4ZsR7Pg4Ez4BG3zNNqRBI20GxGLgoF/Xn1jD6uvj
JCiEHJgjhmVIX2nrLy0b/c0OAwKs/j2CcqY6wtiiNUyXUsSsus2vNV9NzAz5Oi4fKB4R5CTRuEs9
feA9DzrZu7g8Kfona3PBxNLH4qHj6ziQQ4+uEQvOoSVgEkP85QNxYr0djzbPIomv/YKjmAZA6U18
l3TuhRZQlWAivHEWI5N+CQ/i7ZgRozyNFcz8nlprLNW9xx+sUN4vxnph0EA8y9yCMQNaEg4VISVh
6TuNqN9AEmfIY8btJDoV7FZMTL4Nw5IgH26EWbAFCkKOXDJyHuA9/fuYulI2UzgeGyWdMsUxMnT9
JDo6Z6JVlnLKSeeHAHs2KG11mx3GbYs6GzGfW/0ez8pLoxtF4wLrefswja27SGlrqWbYHqdNLSqi
EEb8swCgcXdXtILoiBBMrkPawSZmuFNHctNbqBtUwwJG8/aOx1tZKHbQPfkz5qHGh6sMJNn0PlQR
A9VfTAqCYCTNq3DITswhXSpoKwnjShhTllpgsctTumIh2hAi4NudF8qFKCwNqDsHOHF2yGwh+wNe
Nkx4Fv2K9HVkaJC8tEf4JozrLcpMVO2tJX6/W/Kr5Uebav1qFio3wc8mqb7WP8m+WuAYWwW88qxg
mcg3ELWl5iPL7ThWPvb9SBdW5+NmX4IMw1DsvzzmNQGGc3vHQxwTtvR0/dQC5g+frWnMjRA1feFq
Dwv+ZdzSnOx836la/n1itP82YIjBMuX8GsiYhDxL+Ds7VRvzwGpfq437o9Sm/es7Tvo4O5DMPk4K
TOor/4gzIDxfyFy/OXRRTSBgbYPXU8wH3lMY4kzyGnfsVJ99ir72DcT7XikvD49uhieujrVhCyRa
ouLr+9VtYAS+jmUjARWQU/32b5pgN/vZAqWjCbpvhbUYKcfI2DLPJHkIGdlSgbi6og3GZJiR6UrA
m+n//dlDDlljEwC1bCXI97Ex8q0IChx7ZeXYfu1NPrfqpnMuNFFSd1pBxjNs9Ww8bCHSRrIJJKic
HGU4KbYP7vo697MQ1gOAjTtVnRT/Cv6qebGt/089tlzMNXvQu1e90mfYaGPu2Sh2xd1Ythnk589P
5ag5ndUU1mhpmHN06q2r41HybiFcLMh62NhPIzLLBjJf7AeGAv7Kr1V4X5m8X2HnOpaCEUXQAkRu
WY2LYm3eDt4B1lDrzaLmCl2Ppz7s2PxvdF3MOcZOQuCsmCnDgHlJM65HzETl7Pz/YFSGm4z11KBv
iPoMAJRnB+wVKgQaGo3/zcG/TJgrHsLOHaMirxDgQQiuH+WHSQfPdHkaxftX4SFqGSjP0IZMbhqc
yYQ5l4JJBh2FKImjhoSa3B6BNnCFLV8F/Wx73FOITTGhSCw/cwmTtw7iYjupQ/tOSbPRQa3dkLs3
IhNFvhq/j/B5G53jnkLRGOxDDBR5N2k5XwrGJcAkjjrpE6D4C8165b2B3CL7FvHr5RiTzbRxsT3F
4tB1qKlbnlwu43cEk9BtNcb+hvJFWqm1yYFvnhCDBh8jj5zLcsh7EU991AZ25Cbnk92uwCu2Ljzk
BzZkYck5g7OtNGCgjwi9bJm75F7RVILBiTuztvrZoitp8CCFRejGv6rvjE89bindhgrwinOwosME
qcBk71/RRb8szVOi04BL3XrLLnSNaiWQ455zfuXuInUiCs2fE63gWM9JbvHDFPm4WrN1aVm/K8ld
PocubOF+RMva62ppuIZ9/kRVoVFmnXNByIeFWW2Nx6jE5hheqKSg5RDZEIUOPLDqMIXtFtNj3Lsw
FJAulB+ALB+VShZ5T2k7A5uOHsFnPno2SmFk1yS8F11RvwZSIuGD/5Vvd/zUULo2uP4UlPunddAG
AmF6GdNzzkT11uVIrY/2EkuECA5yBKNGUANKZTe+9Sh41DiFeVZuymvaHnbE5+LVyAJlwXMjOOS2
M3iaOOK2au6Q6g/KCHhvXR2KUk5zkIhcWIJYyU+wpAYJpzFcTZAADreJODtIS+kNxFwdRgW0E4WG
NR140IvesTHeyAJdvqYfOEgEmgJerBT1evEyri5BjykdhWAT+sDjx+tBajzIePT1Q/ZRh+XgkJ4T
RDfx2E2IlI6x1G6AP8PnYsm0hFXlz6TJL3RWZ+0rkKkJ3TgXWR1CRZ1o5IY3lumjSXjwW5OBWuvi
6yQVwI/QrEKokgF9PcmG9dU9WPSPUspsLbmbKAmI23Vxc+duJpnB0scYftZYRSW5td4ODTPXgJP9
JvtD8hiU/WcuQc2sjn9O8liEzRF9tGUGKPn2/2bUCGBTAtb/uEi8iVZuV2psku38M5j/Vi1CH/Hj
0XiKIIHVbB6cO+uvRt3zHKjjyjAC+htx1NoHnpyR4iYjjnNyKrab0UyEZYXQ6qalj5sdEFhmpQGe
BPoEQhoORg53ii1a/zN1hy1VC0FXsjry6biGZHTIMqcwENtjV5MWhnwgKuq0BuHB5BcL1RPnz9vE
8El9Smmfz5iFj9UjUXW+/PaPC3neFqx73NJDZkoBHLd/+6xvfjTi/zUtGgtlXIEDs1Q/TuL2uoPp
pmFoZwtY0al6mBhj/eW7+ep3uIzUDR4goz62qB8liXEYegOevaoQelsHhQvRImWK36xiBEZz7i65
16pA9/rTR8Jqkwc5HkHQSyS41NGE5ALUwATGh6RZJ8o41Fm1/mLGv0LZ4w/+sN6S9B5vvjEqC5hP
E3KcQIXrX8HsIv2M3Pa7xAqiHpAG+1xUp2wgucJ9lLFt/lRjQbmsFM+ThQsqYjJenqvMr/WUghAc
CA3j8Y+ePTpsZBpnaEvThlbVEUgmX4FIfLWaF7Nn2hLCLncP38PgrSbMEN4hm+JMQcNn20KM7w3s
4r6XotTbLo/tIkSp+m5nhGJ2rea/8AwQC4A7kZOm/CnvpBZm5fb3TgbP8HDhCx4rprDk76OTWTtl
azdSjfYTnogxSUFS0DCP84gnjp6zsNOpswGue7zskJWWg1NelOpsYubaEBKoKMPhPRR8cRIK2ab3
nai1Th8xZ0sLMbyBamPOB4NCQ92zq+LweCx7bomd80FTx/uoKPmbZBMWkv0LJUAkX/TVFyjcNQAR
uVV7bIo8Ly7HB6dgSNvQiuLup0Myph8RXPHI2bfCFPi3bjpmHvoEf2JvMpqL9iKEfNlXLaQzyHzQ
XfIu4GdJBGbqZ+Vnx+/ghg69Ooz5DlIPVwBSPZatt7Afr9Ql1Otrug97CyW+1x+f19HFcb1kwXpJ
Os4WE4dNx03ubvOVtUolz8mGjxQoBWxqRobrr6W2+RoYSLeF6Q1HlTdyhewqOizndFJadsTeHj/b
5tiuB6iyO5ku5KsozNLXKBnmUljSI1BY37NzRPoP+TfF1mgJk02xYdpP1slBI2PNmJQYFSkg8s7X
3ROR/yyzPbAFTNZU1b+xIMpG51bhc1gh2D5GPew34mnadAoLWwHfOdFivxvHpUu7k+RcGQJ/ConS
lVCEx3/SpYO6Z3pJqRIjadmeVPXnCHBiQ0bTDuH1As/C8mBQxQYqUqfUixf2LAOBY3VBi/nLjKNX
VSDgGiURnRlQe7Nvoy9g7C2JdhFvK6vtNylalhn3u4WUe3aGyKaiqsRIXF0rQyiqSCl7qyFDRwiI
VGNPAeFzVUXWy7lUvJ7TFZXzT+x+Z/n8LoiU8BraDnGDlAo1IiUk+/d/3RFvaDYAmuXRtanU8Tf7
K2NIu2MTefKfz/f2HAKXZolo/WsaYOTAVvG+c4aK26US7f4b9rJ4XY/Q6unxvNWDorMplcyfFVU/
Qp81A920xr9pNQeDfXaneFFACu+vMIU8GW/eQJLd3sfUKouBOO64XawXho5YNuhVjNlpgPe9SAwC
4kfCR59gNSXAwX7b4yD+AQRylXwiNOP4XW31upyGO6A8T2gLpzAGPocJfOTIHsW1M+yWqU6vuX0L
+N6/2gnIgDCi1iPnYtfgDGBOv0Ty1UogjL4o4WoKBVdeAE0poq3P01PniM+OdvCoOiuluT/Y+eEU
x7/7seBaOwSrEumGje+geHnCCpsTxcqRxz0YKK2kMYaNVpDGF7ICXubQ0vE02sdO0z3LD/tCEFNw
4onzEBWVH4mnTZbIIwUFHBbtAxegeM4ju1GTJ/2E8ydcCmQDFFcNsq8yLUxVtjdRN86p+ZiZfw6d
qEKyAR3Dyds2sMpPJlxACMa3H1XuZVh5IG4ChDCFAMzikicPujlGUcEo47JhKowhe22hR7Oyd/Fp
c2R+akW2VfFlYb3AuvFaj/7YWI397d16IXWLEOeWnSLKWXPsCFfCS75PsxRyA54shHxyrGuLbNuQ
MMnvxlxbnhgYCchK4IBwCOkEV1OqL1+sSNDwx7WjZg7HYdd2feZ6c4YzTYN9z4ZAqfmcUC10ZxNZ
xSETODR3cv/bGyVVSn3AoQriRxROe2u3ash29w7mEbV22ekd73gx8gyAdMKsrJjgRGbkZ37qtEFi
IQb+DGYts3sff72NziyFeSil0odGaRNpBbbl7XDh/S3laNN15SURXPtDLS6IqzG8dz5l/LnxE6OR
S190Mt/lD89PFflIQAcpu2Uqdf7lSa2O4SdoWQzouje/p4XpMyL0Osh9WOZZ3o26+EHTFHoYbSfU
o9wJ3Fe5ygwohv0TI87HXbTwiieAS7hBeWycfkKBxC3tW5300yLkCXWRopRS+D/JjeU8lg5mzxus
+KLtDPXydhND7bGUkGz4QeXHEifGLa/a/MzGx6mA8N3UViIOrrUVOjG6rpLy/iGs2B1s7Wv4Kv/F
q7gCwh323098/mBcq6m7aknfPjscwiN/28vaZJVZW++kWiClQZlDZ7/LVm1jrHlxtW/raYR7qrwg
7uUzlJv/qxNQH3PbHlXU1qKr2dQZlvrDqvFVNFMslJ01X2hUUGQPLW7b8/t/BGLj3RPzd/Qww66J
5MoqlM1sY7GOpljOe90gSKdYmcwHfKgVBDl6tXf9DUI1uyJNKo3OfldkwxGMxn8Zco+msV2rfZte
AptZj4x9mVU92tXqDNUrSBa1ApqRhiShdhug99HJ6ooL+3gOIXxLc0o/LZB/TIa8HvtupEk/tKyS
eRIiNhUnYnOOeDjOA/B+7KJrSDI/ueLS9nL68se7qWlNtw4y+TKUPORt5eJplOyXJYoOihPAMoCi
LQ8jaBwmgokmytx04cjVlP/k7apd6H8IT49Ni1e9MSyAd0qBsNmePiMHg4aRWcd2VAHchdrHtOr/
Eo80PLTaRxMp7UPuK0MbkcZoanYrdTRxJZ/wVi/2bYhUAMFNPMsfoP0O5ux/DmSSK3CFZ0Xiglat
p0ZP6PzfuBC8btpBrkSzZ6q5yHShgOZJX149YobsjfCNNnifR+s+QSVlwJgMPnAwNhqa1YeUS+9R
pzyDaUggp3BnpKGYVh9Ur8e11teUYqaqbH4HeydX5e9fBPizHEbpY6JPDKcyx1tbkkx0xuxc16gt
1AYylXETu4JSzMQv26pUlz1VJL7oBitzd3lvueVm7NyH+UCfd6lwXTF1W9U6iUiToBIaCEpfftfG
KyVeDNiOZeLm2hfszbkVz/O39pN+FS5uD4DVJ3lJ3E8m1byUWbgq7yYaHcnNebI457Gxh/ChB/bK
2slo9Jf9wx1IJhqJCIghZ6jLiKOH8zuAp4SMTAWYdzh7cQEkgHw3ftRyTuVx8NsBMOr94Oov469t
AQpBV0r9uK/evmyp+HZR3wVyykyBf1XmwcUI6Pmg1R35PfUv/sz3z27W2Tp/hVLsaeFrxOdu5w5+
1K0TwOC0gJ9suYrWQCT8w7pMVkKOwxtY/V2nSpORyNjEThzgZ/IEwqexrTX5stgF+DqwMvHBreIw
JHL1J/M33gmnFV0hfUNxfM9Yr3kVnoCEXtM9BNPrGgkgE/rx1bEK74LHmo9pCImmUJvExHzhQxOb
SiddmWrCUNBf/8eydufWQjLIgY+BrA3iN79gjv0qSYzpUpZCr69rJzVg/KWfIVVLz7GR7kWdPKga
eUdlpTbyDhq0Ctkqv3uRQJWgcBP6zEwuBcc/8PoqC44FJf/xc5wQFXPLoyHjNMJdJuPceZASytuG
TvKIsMPlgcelKi6iyTBain08Tc/N+Y4E1J1sFrkgGusbhyN6k5ZHaA6nUIO9NcxmVwkykViXe0ux
cSpnFcYJvDYVMNpGZnK4bZHJWtSwAhUc+p1UKjAR/SAzfjAoXtwZl/wDfvNs3g+zwOKFF2jw526m
tim7UWcFxRVRfxNnN3pfhsK/rYvr5Sv8nTj2EiDdy5hhIO2V02eSCbyCYwD19Fkt1Nv59S5/Jh9i
1R/faEu7+sUsmlRSnmFqYMXd9EWT88ABmlyLGzdNBW8pm/1RF6dAVrNkjhZIkXws5uK78l+/SHnV
4LUA1QDmJc7vrJPjS0GwrA3u2FAK2myd+dJTk8zQzEGv31DSVsIrGY9mJVweyxYJrV5NG2cAbV2e
AzCvlwp9AOY2WUgPMj2ZPzuH3gIWfwTW9omdE9JK/32PKbS5Ue1V4eV/j4l/kSmGQOnowS6ney8p
fnigJUGlU68/w5zYBQupVBV4Ur14M7hBpGhbU7uQrQoPxBy2mfGzju7vbpJm6bcHAW4/9J5RbCqF
ch4TJWQq7Y7ENYHyX2kW658arzvq+BCXVe5C8KrQrel3fgoLVhqInuAywMwhJXKBnhU7GKs3dOgs
BEATteSlinhgQlaNeuhXHzhUYFativMUu3YWNGVGUWDZerQjc2It+ogYB1BcttLxadV+DF8x402f
tvYrkRF29/r/LVpquk4JIixYN1ksStO7pUIa9vAXYbdoyvyWR7Nrx6Ia1PtH8tQs+tgp2HIS9fmD
JhAwNBRT4gmYZI33xQ4/dsA4UuJGa2gMtbWpKteLhjY0HECoWJBbW0X/vNNJU7zXOatBJ2EuEFbk
w+QLbVrG5hVncb1BdH/WBTTxoOMnRBT2mZo8sGjPU3sQRwVV2pg4OQUZzQbX/JzfOP8rluEkEY6b
Bb+MiH2ikh7U4WBsJ9WylcNqPNHYMOdH/6FEk9Bi47yHYb9cyKRnZp7DpHjrXh7i3w92At2wpJiW
22TjMNyqBl4q6noJR7ntL7ICqesh66R+T1clPHNxT1ON0NnMMTNkkelFeLweVDIfbXH7aIaoXpoS
a+qxwJ+al1x9lOb6cuZy/MtD24EWzgrtSUEE5zcgqW5lmWayFvfdhZxR+o2sZXzVZQWCJnJutOBC
nyEWqUE9BCQQ5mJJ8tyD07al5c+nX39jW4BPGvVEhSHa+4jlE+y9yyKvNpiGkSSQNV5dBAvM/+u2
O7jIvrD0LLjiTvMjakgqhajEjO8Rq/yn4aACjD7rEEQqHwPDRIEtH06hnUcCUkMQu6BbFST0MB9n
QcHVp2YBF7t2Ip3Q+Trs2B4NVlmLFrivID3re2jABXXn9ntpg3tXOkXn3Uhh6B+C+g7nP82np3Nh
h8yZ4rmmoJlbmcIRVoDCqRV6vwNGfSLBxrLqCEMQ4sLitHT/5nkIf1Fu3MwtWr430g5pM2mm/1FO
4jjdhf20T8lftbp7yvlfOAt3VC9ym2aHWru/KMElIdAV6Xw4OWySvpTiDY9lYknrv+1g/jOPdh3U
xWxtkHkg5mwrNmGhA+7sPM9BEDP0vYh3pTeoB9G4iFQG4dlnsPV+M50gpa4HpjqsYqLZE3fQfzwH
WxmHdz/TLtnRybbIOiY36x6vEorNcW/IORRGP2fe81EdvKR9N9mXYgyfynUf7sLQSJ00h1w3tz4N
/X7fGVTi+7EPc1k7Lx+L+GbC1LLow1nX+PS7jI/ZHchRXo3h0eG+NCPZEIsl0WpELDqrK/HfOeVo
lc2lXQTE0fOlz7HLAvsxhXjMy2lkZubzVxPiGrd5tyqwU1EzdaNrfLfKdCvr1WdEzXxKlU1B+gpE
as7UbFtro6oZpBLvitKyTVO4yr/tNJk1+T/5bCAEOEeq1jd25rHbJ6m7DvZqGrQPpppJYFBjPhHX
XkTisvFUk3tB6KCsdh1ZfdObvy4XwcKYi0rFN+yZU4UgMwUQgomwHROoAy34qhmRYRtzDwj3+UJr
n0C4A6XzjfOm+35HXjNczJutOyjnRJ7kkuRfPrq/tPb8VL8pt08DO6q0x+Jd2n+0hbxfs/6Hfw9m
1pzuy5IQATc+tgjkYgELGLbkNGU3yDCi0S7WnatwZtBpQT+v7ZFz+3sf20N0UzATrOIiT5m7pvHq
DfrQ1PG2luOci8OLwb7Q9jmNucMUPV9NvbnPgfeF7vy6vO5L77LmdgY2nvsm40eJbflyTbmUzbGM
N0WqqyIiWDhySKeZvdCSpifraSlRsWN35LzntCH98VzjPflRuquH+HVqmhE63dENzWYrv7EPLEEB
njobb4gXirGIfvKWJtp9INeuGmqbfM8bKp/H7U8JYjgJJawFEci9AxEEpW59PoSqF5VnHHl8cd8k
qPycMvsS/3qsjvcBED3X4aojMqZoFosv14vNiZsV5c66Mr4IfESmxGu0msPhAERsl01x4O6mWKfa
VP01NETi9bCazWfrLRoTX4QqpG3LPTPZeejnxj7IeLofYiODip3Htdfun4sSfqUse6ndDG3HsUy+
g0JDVL+OFvDqK0aB2MAoQ9UUkR9N5MLBLMAuaKnAsqY/H7nsAhfhQgMd+lEZ10VGaSZJPOg2T0vH
goeJSz91lH2G0/OJTofkz9vLe+XLU/mtgxDzlZrBiKyVpqW5UG5Co+L4zg3mDS5LYmjUiUxsujkH
dBJp8SqJ3eJ03NB0Uk0zafC9Znuvs1kXJlPJoS6VuLUnkx4vWRhKCM5WiLOk/eCJSf3Xc3ErwNSA
WLf8sKYAThG9CILUdPxRjXP8PhLRYblWL/3xmU/E3t1l5VNz8n8KdEZxPXbwlEJs2i2c8R6ZJMfk
YcNCFNTkY/qLOQbiQVW/uN5trO1vJt4f1ONFPBtozZfIR7VDNH3eMSlWiKTt6+Gt1s7T96BIMYL5
2m9U2d+e1+Q8fucGn6uTPZ/5DXuj9n0STp+DpUsyAN8bzLwJyoscVrf12wRB+Te/Zt2hQ5THCUkt
UXqJuCAdi3pzkXO863GXwU3ZTMAZf/gxn4P/q7BnCf2k3oNX/Y4pDDZ2g5YINfFDNniv6QywSfQM
/ksTWaxFo2K5bZR7vHRvDu2C+bMdHWDZEPWNsUYWOEgoYKSa9FBHsKB4UWyA4m3+NzoNXkaAXerf
kUzj9RVjTx1wTc7Yz4QsYBr9eJZOajD/WjSKLKn1bvsu5CBfVi7YkeWG0cFO7OHbPFuYYAMQ5AMO
DpayGP4KjdzuBSN2GZX+GgY5EC5cXruWCQNkpFFZJNoOBVrYX1WUYlCas1HtCi9UmVWqRQCBTQr8
3mXDJcGgDq7egXw09eYwpqHdHtmk2pkYJQFLYpAnJzwJS5lbXLYXrrAOMAi//1Ko3pxDgoF8W4Fw
M3l4J3GyuERMmefqXi3dw6nKChmWkowCh/Sl052TcC9k5p7Q8fpacif1Oh4zQ+1Hx53Zq9kPXkXT
zLe6M9FocOwirOxs5XsBK1Nm28v8cH2hWwdQbJ2RLT6OGgXKPZDadBJGlsbchXfb7od1M2Tns21l
qOFbd6vxkZUUwFQCjSEA3BrXSyaRgv9Wj4u5Yh66LtVpYZUCedHcjfuznp4NbEaP0FnucMqZi0wo
0YFOJlHFqjk8JTk8MIpiZtahs3o3hj+6NmYzTQxhUSkcPX0TSlQdU27ahFz74G4L8fZ8cZY4mZv6
zXvvRYh9zhXpVnihIzDTs7JQk7Pmr5qhbr9XZN1OVXaC9Rqed46a8924EMC2orLoO9i3HGJLDIVs
MeC0dYl2ODx1uC6xJoYOenhuGT7iWzzVBuH3Vo2YcN6jgJdBV88FmyLo58caLiQsSVaeLjpNs11E
rRhtR3EfHIb4HBCual06PxhaHUlTPLhH/N8lSVs6MRQ49Ip49RMQ4pTKUPSml7EqfZw8D18RfMQD
cDjBQEbvOEKNSM8tigz3YBhI+DBVJJ7SjQUK0nMhTC/3hWZyULSXA+wjqZJsQlTPqfJvTYMFdUtW
REZQDq2PkXYPVIYYBoicxhqVV/3g18X6818uB010ch+zmmIayzjlX0oOxyWdfHR5KGFF/zQs11Kt
YyhHOr2t3pM6P7Kocsh2/SfHCLu6A8yD6lDwsI1fhagCtPdIVwgnfpKjcnhm7R/+pBSY/k5NCuUG
pkZ1pGhsEA1hrz6gkoMVGM/xWvYlnvajpXTEKD0EKiEKMILNsooGf2sTCPzfQFhFxTpune5iDIhx
mtUyRksbi+8hJVgfKvhwWehYBmSv6cVJZqZSOp1PthDQctKh+GL1eI+FL+Q8pnweI5hffrUW/veP
7A6ygZxmh4C5rfCyqYXZsysrZkr2uV3reIWgwbQ451BtH6e5sQsna/bYCuD1+DGvjEpD0uRZbFpM
CyB0kfj+SBN0dnpavfV6BWH/aNk4TviT6qDrzOc+ErAB90dDlQDP3f03kLn0rYYTL8mHCez1O7gB
NRbGkwl/s/u5SzjPuHYuraun8VYmC6mKX8EMcI2vyAW/5ZC84j8/MTyxfqYGTJdri4AqKqrj2lzF
wYNES8//Kco3HccfCNbiNKGeZsTNWPPLyzzBwHDGhmuFYdwlEVglSIbVxtYZ4apk+2Fqev1hjmda
fhyuZJehYrRiHJyP+lrsMtkqJZUHhCz/JtBI1+RQHnhwXtzaPwISpEdwylPvrfTJxtXbwy0iN6bu
Xds2sNYf2K7BD5PiJxra1CoddyEaTNZTZwI0qVo2itnB2gIjHEpzYE+k27cBZ1rQZCt+KZ78K0hK
fkB1sJ7wG3azYjhVCdK7OhpPKHE54ZBUDqOjHmmQ27UJMry+p90OB5P2W9JDoiPodezGXe+GfaOQ
lkcREU9hXDfG0N+Cc/Q6QC0qomFG8P5GfZYpqZmok+IZzHTYuBoL2TPvFXW7WNz5JRthsWf7tSpI
9RJ/C4VMpZUWltOOUzfCi1iJr8S147QdRwSHNRhXdl62PSsjPy6K9GYV2FT4oJV/Nc8fCXJihyo4
u1ZigCnBe2nbKMvO7Bgmq0rcKY+8zJq2weh1I+FUPZ2JU/i2WkP5UGJgUAAqJwwRn6dQLGXPpx37
pYsD0LO7nVwjq2ORh7VDVbVTRlDE86PbtyVWNP4URHwt47ocyOxMfy/ngPu6nSZvx/kIqM+uUx0j
qhY9tsegEU+GmLgChHsv0HLvZs49eCBFp73K0YHW8zSZR7TUpid8+dS8qKNW8t0w3TrXdexVblmO
eBMCsg5PspXQDI59o97K5eglf2h516ybBRSQ+01ez0fUzPQ+zz+Vdww2HNofj9wjMowPUvymHHH0
ROorw+e3HIrYixxp9TRnw5+87DhKAT393a/NqXijqwgVY7mn9t4Ip+Os1kyvty/nFjOFfzbagElM
SFWcsft7H825e4H/F8qA3yBv2Y+dUZVvjfaUAUHTv2afyR8by7YVNqQI6TnpgNWUQGSV8w4xn1rL
Y3z9T5ygXDsBc/jXlijWqqe3tKA3JKaQMEI67gi4SO8QOV9Z86RMICopqQxdE8GnEdTPq6xj0dwK
zLcz9lBP+vQNrBNcKBqhevtw2rMtI1djdp2OwkSMGV0gJG0HgrUvMwKvQJRa3Qk7IyftIqG2WtyQ
KGrKG6yFwDsgucMc6RqJ5MJ7SiLePaT1qZ8bOGM8/ZIbDXiYKzUudc8ywm8GE/PwGwKfxAp/q6EE
jSK8LlPsqU+7Nm/8GaHUqn4XHfz5s2X2c8mfA9rK2nAZrAvFifxepHzbSC9OI5pPCmqyvn59tj33
1du94BYu98d1W5IdMM8kJaUm6Y+VPATqx0/LGJkeR/EOXiQy45ezWeeCYSnnYIJZ9T9al7elCjzr
ThCURTxYfEkdAZWbiAkyRw5byrbRxfSHrsJqZOLTuQ1RCy2DHssRzaaHakFwhIT9qqY8rmOK9mjB
T3uIQWYpOEVqhQrjqvp1TOxJ19oMDASFeyCxURJPhyf0klccQczclcO337P2s1Xs65F9uajC8RWM
tVdPvTbrp3yvzaXUcdIWFdeCIckGUKQuAt44YR0tEh3PK/Lz53dI55AiwCYmXcGcSikkmAOAmdhP
jiHzxRjU1eJgm3RYQ/A8eVUd8S6Cy/jMo3VtmjrjzIgWam5MGXBBiehN4DwNUAEHjQhcwCD1UuLC
01BBCknNAdDyi2fvekUcUb+KubKZxFS1NvhKIXlxkXt7ak/LlmeqOufnQ3EykSBRBycvjckedUna
ogX+TAZp+r75RM/ss8oHoGRvJrFV/IaWxVTzgHHz23xbWWiTADudEfnGmytpXEfhic/sOUHdeoFI
WfK/LUDd8CoSw7W8xyMsDVNqYFe+af8+lI20SvoTXNpMHbQP1eV3yJj6fyVeFyzy+/BHGlFygp3B
qZznxl18e/m0VgNb5/aO+rpd1wulQvdt4x7MoAaDNdUb2xrzc+yM430uqe+1yeMw8s3c+apX0548
vireLGcImRo3aGwOkLZFkg8Yn4sOlLiUfb79MNFw4ZMRZMNDT6djnvR+Ract7/5JtV4zWglSzEKx
TVhCUXm/vVfxMtQRsyhq82PjopJcwrUDotQkPAZksmRMgwnSpr8S4EtS02r2WF3zlW6pt0LG+Pr8
XnrJjt4TlwQjS7YMmK0oGkC0dzHIlq1eorgPKWzC+wUb+g3IJI8owdk+8uf0ovXoLFXuHmsZ1+IO
L9ghszP1jaoUxPVMqiLyNnUxhzyfSr3Tps1NB8neaw5q7zv42NTbRi+lAJZ+vIOnftgm1F8EwcUV
ac4cFQOmFbIFgkUmZrghxTvucV3tUnlAx3Rw1jfycko2PyKw/I2AYD1PqOBVH9gMpqbstaBYeaFd
du84Elbha++B1aaFULxtvQGBuw/ynebjeRzv5igPz6UeJisO85u/XBoXoi76lxb5m/lxwaCOwQIi
Jd0JRoSE9kPy9f7KFF7GXkyXFVaz8KxAOfFdPRKMy9GbRGMbp7W1Ix+obG+yTf2b7v1+xc0WtfAp
C4pptK1HGeTHmWhE0NS8XncsF4MfMQ9/ZRTmth31InKL50owBhHPUFwb9eOXQVnF02YpskgoBL+S
p82Ebjq8s/6sqQRRDzrkcqdRMH+CaEum02SMyc1tFPndg6mGjr/6kvebLjTbpyKBgEubdHqIvtpz
buDaxZwMjxFijEgFCIv0p0rp14sRUNYplwqHCocP8FPHfCgJurUxcrw/B+g8Dx6B2DQTKabrr8Ml
98etIgDn3BB0+LX7zLsgJTTtV5sy9WGIFr7E5jg49sN3iXhOVJW0aj5SYcKdeE0I6kIx34Q2K05a
rLfVMMajbmRnQpCYhHe9gsokRB/EdMN6Qy063dL3J/6KBzApmbnvkDW5cQwh3mPKWNg1dlkgiQK6
06mhSuw8LkKnq3bUPdx+mttP5iEEQnpQSftxhg/hvMrICDZv7xbntrGYn2VgQji9ZoMtogVS9NZD
bK66jtVBZ6utpD6xsWwL+ddKttzUoon4x3+23x3AoI1H2RDa6wqp3UsYWxAMxLJ10jAmnVYD6rDd
BO+QTnPztcl+Aqiab0gXSMrZhP3oqJVaYrQwjQksGgTGehGGf7JRuBlfsIuWMeSEU9fCbl8WyVle
HsLFnTFkEIjnSJ/bohueu8QzEb/Vt42oxhRqOV/4V9zYSIB24wZuuRWKFWwDWvbYdz3tHgd+7Fo4
Nt1IR6KXX473nixmogE05CiHceZsBSQUUU5Yoe7ZDDQjn0shIjBtX8T8QOeAME1zooQx5ujS1Tb2
jKdiuYPZbeVJGWmYvf5hmZ0jOrMOxVkEjEFAV8QjqhTixBGbe5g9M+c6nr9H0RHVnddAJODJA03W
8IQ5jjzI1cJ18fIA3a7dRGA060DckKeC2x0m2XFFNs8NZatvFbI3DjK9VB/5s9K4NHmkdG06Ly/T
xB0P9a77VOBl096cQ8JCBwza1MaNR/Y3mS426eBWSdDqTNwNzXELfv7GXv/tBvJLRSb9jztgX6T1
QXrMwYrghc1NoVEbbIXYire83UqNCj7jA6kVm09/H1ix6k/TO0jbeO0uQDcT/WYAgb4B5WGHMnaY
/v3vJkH5U85hWTy59ax31UhZt3bvONrxcEySDOcslISPzph5DydNrnptFnDt/gsNt7Qgzfn32gr0
ZTxVHHV01b03KP6pmwG+zCwviYDJ2yqt0QB6lHT9hqTvmyBAchEnaQheQWI+KTO1z63gSXcK0Ld4
j+DWVHlCKe8CPOzJ3GHSyJfh0EFzKjc2YlyBNWd9kEA2rfVMtzyVj/J4lct+5pLl+Vl77wTGP0z4
LVSfoSnWMCEZLSU7yKawitkKeUs1KVg6ZAMsXXSTSxDwqTLhrFbk5pMXs/ZCrdBS8gXz20EDlGje
SVB+9gUAXiLmTKOY8rLXcTfV4kv/0poqn3aYlM3Vy2UNC6N5M4fXLrfRG+Ptte5X2CpqOYL+1Eu9
V8zImR81kgXZACZtdMnfwqB3o/zHk/0BBGH8rk79CBUylsnDKrkbOTekQNw+Zik+QAZJVbHDJ506
TmzIE/5nOCMH2arpY71AxoRGIsPsNNvNax0FepAQpl4fBXlyBFmo7viZgJR2XIBMOascU3IxUJdA
h8EctqPvrgLtAlo5wM8rsX9Ex0ksi/2ZF3bwOIRv4xLKcn5HOjfiizaDag6Bl8TnxXWkXfijhzcz
kBIWmUg4PADNdZLdwAy9V4RP1wlrC397XNWyCZs5M0WxK/yewWlImDO/HAaOByL+zMtFzY0O/fvB
MNdkTnZQqMayJamvdyDkmd5MOhlohBEiW89g+OtqAPHPrB55j43HcZ5CkqPr58Dcz4NbwaXBI2Ox
/5kpHKw2cQNn9inemSX7GfiEud6+eoSO9Syv4AN3urwX/m2FV4T6Hex5sE6qEwaDg6aBilWMfSJe
VwqPe6Q1zdv6vI5yPhHpkJXyFzXdRBwuc/FlvDli3JXUnK7vC2vewm800eKrJSm13whpYPSAbVqK
s+gRt29fNeUJV36NaT8OqDi5VELr+gl4U+M5+lqI/af/I9uYAZHZ6K17pTZ+Ob7TvMCQWznpISiQ
auV8Rv6HmnUxgRMyG7K/8N2XKToK87Gl6DMgCIs6JgX8xkP6AJtTeYXeNKuGDuExMcn+np4lox/l
rt+tRkENnlS1Q2SS3OZZ8ZNudDJ9/51TlY7HB029YRs//Qz3WF6y4ZgTx0sKe1SodigfU+Bogdag
TZOgpXSW4GxVauC/qM9KaKugnGYRLc6VYuWSu6sOgaYZYa4wnZU/COYtA4mujhTm1Ib5F/EcMspi
2GJ1BAUPNmwl9oTwTWWkyfhUMk7w1+T8E9lFhlNj30UysTDONLNbTg5x8fFrwki3zWCW2OnFg397
7sZwtEdgpMMaFSFLQj/HHnpSiS5jBDy15Tao1myudJTg7SbSU1sXjcNZsGz3w/3T3vk4K63d7xlv
49PLa2cvhzeQ+borXFBZIO1PQkBVZR71SP7Of8zxfDzbFUHnDKpT7zbgq9eAoAX2UOdY8I3xH7Oo
R3FBDEq7sw7umB2hTIqlzzyuoDBt5EPR2zVA3DOUM3kWemrsp9YThj20mulYLDwrJRtBLOaZB6dD
mSa7dinqsHje14uXuvH2WepAEpwQQkl0684VoDf7sakq6lXpm+VXG3MyEwwLjyhaAsCYC3mbsjpE
mLOqZ4h0En+75nbLPWMUjVhtc2VaUhM3Gcq7BNZXPm/u3UKLfFYuAIgL9iFNdLlbcXjoDRgMQU4+
rIrx9t9y4hk6XU4DDBiuuNmNWMaTfXYLvQo4RYk7YA1I4OZAh1EHfmm4GKLfcPvq1+Gkg1BdIaXU
noiNCuQWcOZ8mTQHSlLVR5huBU8nD45rZMu/TbS21qHjlxMFhYg5dGiMxXOi6Jqaj6ITz9/64BIB
9prlybeeL3qwZUTdHKsx6GK+WEJeK0cCFIEwCJduD8fj2O2fpIRN6LVzNLVxHyUvAQDf0jC3Zx78
/JFJ9Jb+psiHFl/T41BCu77pI1EWHJKK+zIV9q3dg8XRfn042f+sbJK1rDTysv/JYx2vm4vEt6NS
RXGgPXdvhIVCP8ewEAtgDz0USr41WjGdOEMjAERgN8aPVW+oy/tB8Uksh4o52aLXnbzcHKiVd9Rp
bd/RHSuaFrmnEXS9eecjj0xgX9b0ZnE9yuBPvwFek0rs/oi4F63HsxsaFGvNc3WcqwKHbfBbacJM
JrvEFf2tdI7Ru+K+7KjNx06djdMzO7znlVK+13mawLtMQifUTspPIsSN0roqK6bfgCiiTL4d5mNO
PjR6RWhbqP1iwtkSc2RDnX/kTDBsA6l+xK60gCMSH7ogqItKonYbhJTFBqNpdNtRog2G7jc7YLuc
VsQTmsmjkqIuveHe9rrg9udkefuvTFWa77jsWrCPQMLGgfiswiyY9RDhUr5dV5mRtg6lSWAW55hD
3eMdGin3G4kDJhuS1kkKRu0bT68coR7Bk2cecygLv1U4A/PYPN+2pDMHqJZRKH6W7QCwTYRgyVDJ
1Q7vV7zHBkVKWeiSJxKEMaYpqmZk29FNzlfsJpLX5aObcH36xKuxKtYQivClUKUsECjN3eam7knS
RWxRTrjRvejtak8Qe3yZ2ylbK+NvWNNSHHAqv0FM0EG69e/i7ZXPA6MvjQHoqBy+GkqlWo7M6u/r
K3IRW2Z/v+bZuQ0m+jYuFOgVnlYS2dySIEUx5bRIcdV29yZGOUGIy/HOqdbRIN8/FZEt5bLDGhjD
/SfSyOiZxaa5JB+CrHc7FWjAAkq6WfkWYiF8FNdztZwug30GMyP5nr0c/MaeO9G8lbMHsnIAcnlO
EmfZJSo8HxwQhidzOtGmoXM3OZduIqSy0+S6cnCkLfteB/QoniwaQb/jhJl7EIv88JG1crCdG81m
g33h7Uk+6mT0cr00OyHbz8Go/UtlXo3KlJlOZ2tx7rMnd8yD4FSfZ3VIbrwFfjc5brjxPb+8RULF
cOsygxBWDR0Z44vN1KIX3PpCf9onggzsUtrbLFe3z+kx4LYT/NMUpvFsqH+4s5rMdA0O/ivcNuBO
8PjQZscJ8eSYj636L2Nul7D6VbTYrjV5aVhMQQU+ufI7s94DemabWczyQYt1XxeEJMyhnGfc7RvK
3aQPMjz88N9A48XMwFs7KrulNJT7W+8DfT1LR+A9ETZNK/vpj08rsOvQIASZwcl8NgPIB5ZC6rso
zu1BtKFzpjr7VVpXB5CjzJTaVIwuPUy+/jpJ434FRWvybpcLxkEgZgK0tG6SQKVnoXJ08pgLGFjZ
8JcVHsYWivizocha13KMdFjoscdpE3viCY4JzW7J/Z7a8F9z4PHftJikvhl/FSj0vZl+/Ewb3RK0
d/X/2Vp4ucihhKl8D8iO86ecvVJxVD7qgCu6HVzXQicVork+PckHtdyjAKX+4TFkDpLMmy8ORaeB
wzlIuJNOS+OF95scOT4X3EpYfXU/ER25pfiuKIJKKhCtQiwBBF/QA/vMNWPi/iaBB7G2P7EMd+mv
piQ/JzAxrKUn57XN9X+BaYkiseB3JoDZyXMdvALRxb4e0/yuCXgKeYyipmCSpPQ523euZLCYtn5e
PD2LB4m563wI706KxLRFyWeRbt5260b7oMhhpHdMtrMKqNRyJpZtBBYOP7BmdO1G8BVqXObtera+
NAITObW9S0v8IBmwtq0E1DPJTB/ziD3SP2MWKmXwpxzh2vwkQOoUbn3cFE9VGE4jOuZnS05evr/m
KbYKhbGXnsrx8b6JZjqylkFVAfFP29EYYZjIMwhdrFKpMwOpedEnjnv7hRxjtlqp2hWroSIdtfrq
Znpvg9HkMBKYdDsD8BsK9jxIz7Cbs9256a0cLplBkh4TD6rTUEJ1P+iHgm+3jnvmUb1kavNQ27ce
hNti2HPd5QWMUkpTFWWkzRRFtQY33XpiWQeggd4pWQEogj48YJN2XVN8CTKcNIlNfkwQrqi7Btp7
0RirOp2LKdyWkA97oaoAutM/hovKMVZuY+L5XlJbejgcRLyGwxGv3vuMFT2TFD5eePksCx5+VQt9
olJoS6ZTfwNN1yzYKjqX8b7eypc/MSb+3VhAbUgzDZ/Rhc71PThPfOLXfscBGOR8AVl7d1SNMxK2
N4lfvgZqMmmA1j8Cx7zfUpHn/G4eYJH8mMuqHP2eKzUZLNPNEt1qevmzMhoQZlJoljZ+j6Aen7O3
Aj9hbHbCjUrPWo6kQrn32n26btNNwQNZXjyTB2RDmKW/0beEQIppYXl7q8AK4HzdMBZg5n0PV/nc
ajIu2brzDuxwDmelIpsKbStgb5JjoS/nqH3V1mt+Pz6BagRF0k4Dra+QbRISqpC8nqidItsv6wxF
7zjkqEZ6UIYfl5ZY09fXPuonVbR17kgN9W7oN5hfvXQimcyOiBGMRpRHoxlXC1BJvFMt8uVY3vr2
9jiYJzv6iqbX+KGrqEkkip82ARFeT069bOduTVz7QWKCUZrGm4cetYJyEZp6URW5UNdEG1ls2F8B
61sXZQn8/UsFSTAPnhPtTA5/lIjwdBE5HHKVC19OpejdnaKTNGaygMZHuN9Q/FCqEZDA7XbLtxSv
MdGv0Vb96l9EfB4zvXcGVe2q6yhQOHH0ztkLefYGgXLnhxuT35ds6FYTrxwOd48lWZGo6EbhWrJ9
twYqdsIBAeuaZc39CH+o8xhuFBn/85YklOEXQ4a15/s2mNFxfaaIUy35cuv1vsfpB7Y56W1lLvb8
zij4qftDrTbycgNN3td0QgCJYU14lET5njClyufLNS3J2I9u1DNL3YOrRtpMDvAqlP7lzI6NsSOp
kcu0FxgTQyQXdyTOXQd4HKoBAasUq84w9WqdBNoyqGC8eYrLPeZhQDrGdtee5Rj29HSbywgIQXw/
A3ES6/IiZ3poDcY4NFpbxLcnfjAI8PKEYRnbDPlz6Z8+4UHj+FUoy5OgWn3qqar0hY5gvU8ulVMD
W4x2SX0YfyrjdJf8pRghO4Eq8QKQSxzaA8UQL+iXcVfbSbMBY3L+wZEG02AThGeBnjFxChFlot95
3OHry+F1oXz0BZzMvBrZqfHJZja3paHEs5thNKo2VOfnVa0rcsf8eU7lr5ovt00+d8BIB6o+jGvO
z+A0UCTaC2XOKOuh63Ryql9cc6P1uVvsiwS1u8OiZ64TQakJuYETtGOoBolf4vAA6FnWxSarJCyy
DX0PzM6uPgNA7BZ2Y4ycf6jrQMBa0ku6rGl5Xp4l7+r5JNGglBELutLFBSKUPvSEqtSR+BV2D024
Kj78X0GI42AgjA8tA9sooFiO7RM/PYFoPwbrVR/v6ZgCAf5OfIZU5tqsjPwryo+3bn0ZZ/xRuAKr
KtEK0KWqkZlbloFSoxDmjYcieuhYxCbC5KCEYsX9NWWcn7i/1oYgezk0QjMMBPi0+0APHq356VMY
ANxr6o7ZyoDplxMxDQQmLfACZjTMaAyckMYQFW+g5ZCEDal2w2bSBUpgCfjjcosnz2S3R+S5U3Ve
LmvYdAAwTpE0GiZgC3Vq+KIs8UyvJUXE2AeDdbMW3m0iqtqfYwbvUQZMDrplSVWx2CMqsdP2gukz
xv6pThQd/DGQSRgChUc5O5JixMYe46xYtQJZGU2Q7RsVxZ7rFguTtLxag7fi/GxXf3DGWJU1MN+C
JCB0vMo1NL/jjijxAYf25TB0GUyBvqHOCwkS7qLH0TFDav88AD7SAkXe5XZlzs+3PCJQZ1XKwkvU
vRgHIy0/dm+SovKetBnTuUB6aiDq1xqPQnELiglM8jkiH9bvi7MrmIosMZCHu4aut5DpiOhIQGVz
VXugPUJXg+bdOdCsLOMS2sZUTwOW0lya91RvGI4mJGYxy7pTh1tECXbGuZwfsIUYJJ0CeclLNYvt
XqxFcBqAp3woOGgQWzcPCXLaRUvmNk5nVpdAI2O15ON6q17pMFTlLOHIWW2nssegSfW9HP2cUpfx
b56eoItTaC1V4dLSvijKBstYzMPWpWqW+ad8Jfc+Dh1ah4MmeITLvi0hcXoxwl9Z/2GIQwRBHhaJ
I/J5n9KuS0nIyYj9KnWWlTt5sOc245bJzTyqNzu6N/rRLN82ArWU7Hmno1XFkkA/lwQYCDoizcPy
zxC7EWYs5s8/MU6RQIFlIPI8QW7sKKptwq8SnyAfVVSA8Q9Lr7mClBfCY1JvPkARbEqJLnSzIg3b
zRHloRmubOIHNkvEKcvhoi3Tn0GbBqsEIpLxWRMTNNf8mmnHVc9ki2TnbuCAPf3R2qtjA9AIJ47z
OxOyBlridsl0qJ7VsSd+cjCHt/SFUIIz38ZzXyp51KOw8vqDNTAXhurQB0ebehN2jrQmpp/LSEZd
7kyLhx5frd/HzPUmoKA3r1ee0bHGk/g4a5Uh3KYAo5ZxiQ0ACbZRF4sh9Q3VYJMAAZUW2qHaygwS
zCRvBJd2bZlwIBp489s/NvYeOV+4yprfs64AwwelaXoKhX34srMCaCxaoEBf2o+cjzeqe2Jp2R8n
7le44S2+J1BjFNBIDHCyQI/DtA0vPJT1NTlvRWsUkwsDu+yvVXOI7YcOE5iCedXCaYxAnVuRxeDY
MiYYrCEjkKtdJ5S8LFlufJJP/erJL6p2dFfJEj8wIAgQxYN6ftQcxK9bHtpUtJd8L/D3jUBav/1H
+/v0MUW+zsorS/WrJR71y9/+xJOG50qplbzboinTJsxgJ+zfTI1alOA8reDpdyx9EiNY4alxGxGr
+hev3GPgfuFACjEgCBTskaaJlvl8sLzsZ/VEMt1L8SnVpOsLhjvia/r5yx1CXhO9zFtzOinC8GoA
DC8FliYUHipUJelAbhnidkJ9gQ0GE2SSBJJkKNhVYrniyEBV1GY4vCuT43OBMPGie4QeYSd1W2Dq
J/1cLVmro11n3FIDDUD+UIp8tF4HcNF+0CJo1CP0fuaTCnNYgZfZSsNlW0o2n2knZwF6qQCvnuha
TfilJ6QVKI86hYn81s+DnKghYugTPn/TTjVZjY7N3r7AdNICDmbG1X8an86w5LOFSR5MKUgAs/KA
iyjFpKQ7dOqVWvolHm5Xt4Rt3QSYQrYBYS4NEaYgDEiwXRWrwCM0+tzsGFbZtXH3uG0ZbaTBlkVa
ZT4SvcWE7o19sNwmrgZncsIb14RxN7v16TvvgoV+MJfV1TGb/S43Iy5gIueYdhzxajVD6+Fu6mlF
/9QwhZQW5kOBbbAe0NKMbzBIGyIwKG5Nr4DeEDe96GYYVbsEi9ZpcncCFF9B5oP0p01Zud6DNQ48
6lq0nCxvNjXzevW6u/DyJGUejAuEPcDDhvfgS0VZEDr80z0JvTwwC7C1pzqZcDT3ktoiCfMIG4iV
eMfkfudAQeOHmXeSlk7B+dPZAFqlpBF/3D2McZufj5e7Da8DoxDosHM8mS1lkvffA9JBh0zGpefm
Ftwo8Cv/+BscUSBKYojckeXHISOD+BcvDyTCFs7eaYs3hKOcQUcDJWc9TZSDzgPgLQY6QVOmMYQW
DeZQokfyoV/3ruZqO9u6/Oy4oCNQTiPDmvgf6/krmd7Rq78PVFYryeWEdAgCBgz1CsZQeZLGDdPB
x0fGnKoeDWC25OKrXJLy9gGVEzwQDdtjs7Y1hpETdFun7AR9AjJLXTPKbl8pEnRSKPMK/Y6PamFM
d0AAFwnHMr4SfkoPUF+wDU45pIxTUAl1k0Q1QeRtt2dYg6KApiMa7glIkXoEd9iaFELkVM+tgNPQ
SoJiG0bPeKAlgYU5zC0s/R/ZzuNDR+X276Zak+RGbpmPWq3k3dIRYm0HccZ0gu4vXtCHDEKTkr90
gOG0DWXIqcUO9775LRoeVH5rWvcjBmFQ/XBMHXfb3eITwwq26HLyBGtH9dmE54oe040a9veekwhW
B3IucfToKQmuoZwXYKOcujKd7Xl3TXste6DZ5OMri6aRZLftsvwnbT86OJm413WGzSQM/3/bwOg6
VTA5m68Oh6KSosFYyzFrAYPUaBSszVTqltxhaCkyhSvtcD68MGbWo54n2N07vMSCOCj55XtlWRtm
eYrPH+TP4fifAPT9BiWtAmmMMH0vFpzyDJpEz3EDTJAPhP5vtwowXSrR2dYIFLCopaPpLTJNHAhO
s8NKwBDZ6l53J+2OKqL6+U1vf6vbzmkPC4rFJF9z5ml30y39WfDcu7rVPx81v0d/qOJXo5r0f0ER
uej9hzQxYLPAjrnSP+qdahjmK+5fzSpz4kr8hA4kH/nq+iV9j/dD20v5ujpieNhWjre4DuN+k/Fb
dioD5BN/+jOHqB4HAum3kdfy13UZArxyfrjSkG57w7DXiEyqIyjq1E8UzZtFvirkPNIlIqmOdH+C
2Di1aTnAjtsEcDY2kZcmbQSkqhd3RNlHQb8G14SrW8qjXdMhzMBtG+BdbKXbgklVWfcIR+6Sd7Q5
GkEbYvGzFzGcx48FYeKafalQlPjbrkTM1gel2StqRt2Hl2oGvrDOKcIicMp787R6sKaTwS3ERfjs
LEXsFGWIGALNFaH28cX5rky8yqK96+dvSLau9Q7LvLFQ/xC8C8ry5OCrXKysSU0p7E3O9KK0dO/5
mTOZ1YeF7L5NKV0l9r2LoEnDdeLKcCzIGVsQbBsn+VRa7h+xCA5r8O6ulEMGf0fff48uQfZn+QSq
++Ixlohqwh6iZmbIxBJA7E5h5wVlQa6suagywdBM9IUrbQo5I45xyUuCkJgpf0mnuVH6jk38YYqq
E2Q4go9FIMlZqr6EP1UEQ/I4xjX/KQ5Drxnx+i2xCFXuddWW+oh02sbcQ4lmMcjrt7UDrYlXc8qP
zJww82vCFkSkzvxFe15EeZO76LNOYPalx5NqSewpkNkIZojOvIfwi1J1VnJe6/xMVpS5rBu6KRvV
KBPyX/Pb+eaU7kzli2FpS+lRgTGNXkW/Zzy0FSBkENcTTiu5nbaNWa4nZCM7CCiE3WdhqrtzHi9D
pG3Tzok+bNczkVVU+C0/19Q7kUM33VfYOka9+01p0YD5TTNfhTeK7U51iku6yCzpK4JZyD+ubWVs
4SjTGccvVpsOJTDy4Qz9DQ0aIU1UfLZwuJF4r5zFPtUq0e+wG1tiOlTdoRRApsNmdaE6TxgmbwTt
wURWcxegsaJMPlt+U+a0fZy98BaxzH8Jbb/f7EmmLNkScz6kYJHJ2cdxnEF7uejUtPEVVRrLFq0E
t3QZDov18z5K2RSevoxue1y92Yfka/exs1ZNC6bjAKVGNZR685AWL1h7nK22Te4qXbt8KHQR+Vyv
y3yKKZjgKUxncHo3g3AofrXHXNArqqHYGAqmrPk9ijymd68dUYTHRR2PpxuveB0Wn03WryY/Os3J
1FFp+uF/IP76Kmv2dWgn8sPDjtWiYAi5ZktPxoFbsWvZA6qri2kR2B1JpFMZI7Qwvh86KelPQHQ7
liM4sKYTJw4OCjPWCV6RgX3Yte4BqlTA5342IDy/dL3LxnYtBKVtHkSV3781mz7Pcn5SqX/FuS5c
IuhqFuz7mPiGuoMdYHg6XbFUA4bxOSOouClTpW7yRT8IEoDJINy8IigejkuKUszPJDN4MPkA+q+A
CjT6p3naXgbspea/VDBlG75JkhiX4vVfUwPolc9HYclu7Da4+GMxvsATD+xmMSWA1V2PPkEC04/0
6/O4CRTVx7oUD/XCA+f2FN8+KHnJ2Tct0KScZRCk5TLkUfezybV6adwZ6AKC/poP0mwaNEFuXnTg
q/Z8fOjgcNTT97rx4gfZTDj8+v1kolvfVTVhW6CGSaxJai5nbcBaQjTIiJzoFfmh4jeE+Wshn4++
ALFOoigvkTVZmTauHSpVJdwpu+rlzrsJr03s792C/6xmdarjUo60R3IFTLLwByr/GNtHZM5hV8ma
h64+/4A9DqxXFpZa+3EkJO4VIZgHkdqEQqgCLvZ0VhAjkgSbaQ79edVLEh2zYNEXzmq4UdR4DdFA
AKlNqwlaFLHH8CtoO1MqGmmatxv9v2mxsxeds2KsTZUeT7qWeHPufcVOKaqGyJxO/1efzU5rSFwZ
YBLwFfQXWYIO3Mo6xCGy/65H/fQBMyTxLNFwqsOYvl/1TK5k76liXOVHHsY7HsJ1bKi3nI480eBw
rgzDeo6A/REMNUi9iT+13pudjthhYe3kwN7V1egGYT8h5isvHt3Eefp76Xm6XcEkbINzMAKfbqwT
qgfMW+HccG/6qis36WgUN+briHdD6hz3zKoD2VKegvRQjROzQmVhUAX7Rnn0tJgssQrTYxICoVuP
Re7zduTHYpqihosAwefDZ3ONYQ9Dw70oL5oa9s0SrLIlOowaZd6+ck6TaWDbH6GFP3Zyc5d1FoCp
BlinN4YzEZJr9+qXZooMCBAvp9j4uFKxruyACmBSWWeTf7y81UOExD0waFWEVPzvHWXLBu/mFueK
YWsDNZgNJXbt8BN4/3+Ss8dF4+LNmVL5gE6VxKL+G473f9rGDPRizFs4noPJuO6N9nOTXbXeoA0i
pQA5qO2tz4kJH7qvTkLPSurSOiLrNOiHhV/rciXZUwrsfMAEMLEYtW+1y/+RuJsujmwRL70V86wn
DyPrD502v5wcG9RrVNrRbko/8KBoWRBq+JSH46XSRJ8VE/nTN9mTtC55nNdC02hY4Hg0ZYuZmKK5
3qMcxA1kQm4A6LMJo35a9xKgCXI7x1ADcE7onIvnP0U2AkuBopTjktS3NC13bVJqWCgmpBrM6Tjx
75n5KCSxTK47WBhhKFKYr2mBMyEnESEpKEz1iYYiWVpEfR16QZW/Vww8ZE//IblHp4F5BKGG5FcE
vTsrDuLWMFgjxIQlI7r1+EhRCGL/XoQaVIIOsISNELmYWe16QRcUOeqZlBdevA0bZjAPewzWh9Bx
w6qdNWu3OMuf5E/LMg6OKiUmP8mgdgewJ5eUke/4ZwLPxCSBsYHtWrziyAYvdKqECYseEqwGf90T
Fy6NG5ZCqBSPDEBRsb1KzutB+3Dm46hsK5m8edt/f+r4oqp/9+zQ01vPCud8rC/MTmJz9PMzCIeS
p3id+J0raK+PDP7RgREjbmIMfsSYsqGqOx92icV6hhEB70EnrzguPjZa7mTAVvJj+ntw7VozVqe0
MXV5pAGDCr/EKngM2hShICFNB8r/hSO2BdK4VVC/ye91qdELHFD3ipWbF7DhJckwUt5EBZpNJlfP
MZehvH4iX7JclPHhMDlM9PG2482g7SsM9ZqzSLiL7ndqNDoA1NNNDCc58Ijgd1wbKFt8CRPrJ/QL
JpX055XlLiLVmRjuMpaL/vsZxYZwpGVnTGBxhyndt/n4YV2GmrzFwc/VQr+VgQhvCvDVxyTjSyqX
NxZ46QfcEtYa/M1+UMxQcUyiKnBLUGzih/iVV/QRhKytVlCgwPdbGQC3eRgehB4R0INi84OP5PkX
FzL2AgLg3OpeRA+LJDZpyza5B2+O+GSzDMnaN6l/QqOZsK9eSH3moc84AgJaYm78TAKzRnuTkgSI
Vsgbxw17u46vuGhBptiJ3KPg2EQI72/G9SPtznoc7byLkT0L+Tn94HD0rnKxsAiN9Y4ZBSWWRq/d
v8C4V+LPSR9OP77KMj4O+y7CnVYg87V79f5PV8gkCfBaVfjDp76i/VMfumTuJv0jv3HLbkVGZC7V
yh3D/u0mSbxbCtzFCHxSSaKYCx9BOovlJ9vFNPptjzOcO0l5EkvTjtHW9PYn8BgHRdC8jfSjUYxo
fe2atsj7iHI+feqWipkt4bIZYp4VynVU8UwZDHoEiQM0vtwpaYAbCNj75lJQrkYJ7v3OIO840kfj
HLCAxpFI8TY5tNrSqtUZrHduYwJ/j7jRVVvMydDXpP74gMnXPsj6HT4L/NvjVW26Mx3wUODqb6s8
ICWTjyKduvSXoqREKx+PuioOtQ4n1/SzT4k7y+Gs6WxobtUrX5X7W3OSChcrCOiv7j6pN3mF+w/T
PwD+W2U5WR56DffXjpqXOs7qE+Bn/kpxnoNI6IIXMNret/K47YNuaPujUO02DLgTZehwKs40T4Hc
VG6Cyj9aW2hWrC2ICNHG943XPQZNuwG2caWZHNfMnW2fTgbdpEgx8bj+10cdk/CIO1AAX2McBVIz
3SAhcBb0hJ+NtCS7zMiseyR9SxTuBRsjJvqQnuctssJNBdR4/k2NhEm3ux80CgeU8F9TXveO5bV/
P6wQ15qGmwMBdkUi55JacX1c5a9SzXCJEtE9XC1EFyMPiWnPdzmIat25/mIhfmQwOldVNzI1CbkD
sN0a5zzsncKb30yhYeScy82Ma5oH/bzV2YPoczxDQVZH8gaTXEz/FvZAUc/rY2u247Vf1ezNvhwg
4qwdGMO6MoCTfCqs9C5ETrcmayQ/uOZDSLFc041L75F1RBiDKvVXSG8soVdfRmbL7dYluYfN/RVI
F4g677ux2fw7OEq/PAbBgCWDfZhVanrj4UKaDTmukVsM3/I29aQGxXVLQu4AB4c52u/vS1jQY0Rt
DtWLivaSyHvjVqUAGWuUKjeCPXdJEjsyPDElq3rm2LiNmykF9vtls9aVZdKsqsH5HE3a93vicKQO
BYWLv86a0PEN45x+9eKdzPXSPaX5r2itvdtQo3JoFBdtrr3c+QbcewOsCYFCbXyr7i1OLsjMLYQ7
3L/8DJEgohT8C1hRAkpQxIJ6blZOllq9JRioDUYdjv1vqksGA3vhbxOb4xTSaVShXYGtzSegqUSn
z1jOBDn6vHWX32aiLQlmbvnrAUF2URPfkLJGOFDai1ZSgbNn9V/CKSh8YanuAeW39CY/hBOqecOI
QUlztwk/ljJjd2VtZBstBhZXpV2WM2DhctJbS9nMZ0YCz5aRIQHE4cF+3Q8x8HNnOpteY9zvzFqO
8sT2b392qq+VoUxmP1TSkgGKAsqa4YJFNsgfTG57KT/+UnV/hprQzIByyT2HzIn7q100uh5f1ksG
/ctl38GL3G/B7YT+6lsm7ijX0C2CC7QNRdKx51vpaYf5CkgwMKh9f2hyGOdnYBAieCeuN4/HtDw+
cLQzNN4XlwXZh2rrvAueaXTkjiLbvQOaOWuxdWtcnGL92mFSl/fkXBGeS2ExjUBwevczsvufuMk1
QF+3ovU5eVXNL+o6C/V42fMJeGi4qF+ojoIJjdjV323Q/aLyXqGx9yNADrAq3cPp3m9KEXYbfl5s
tk7fBlInhLGl3Z0RKGIaAzPsTdi6sW6z2AlGUplCMj19JMT4Ll8Nc7wrquDTyCRQUCVNyKI1qJAn
TaeRjQr7KI4kzw3Nk5p4TCVPfsmgAOEQwL88II9ZM0FNOI5I1IDM4iOnq4rPIKpZ31q5HI1XcWlm
eeAW691zB8eYK2vcQdu3orL/OwCDHP/T3EefGETF51kiZAibApzfDL3p9LB87copdD2AxEFJqjWP
n7bZw6eW8Dhc2l7I8zyXgiJylOANt8ms7+iXXwgHd8uc9QuEmGd6EBnV/4YxL0J8WSsGhiBfdUc7
31oDkCvk001M5Sq/y2g3hKJkVdc6dKEse4nYn9zyJ1QEEc7DNnX5sZsjJXjO8IfnWEOsXGf/g84e
JJPpcL1jEaKcB0acAtiMK45hQu0oBvmLIj6FORAse6X7H/UZhxjo2KVCIdoNUeZh63dIT9OcmpdJ
DYIbFAkTwHKY/l2rh97Dwf67TQ2IcZMv/5x6mHHKBk1HdGOJfl2xGIIv+iyECRkZucHhSyIkSTYk
tvZfF8A56B5DibOiWZ3JzkODBkOFVobJNjB+hc5piS/tQxBu5zuB5fL7m7Omz/8WSJEfNO6yvGOo
3cLhH0zmwPh79qQmWeW+Ds6+o5xjHeDkdvYbytdfqlXDm0g0eOiwkOIbmBcTbnOD1WhbDbmuMTpd
qJry+zHWm9ptXKLDphVQcBJDFwsZ3II7Bl5FP5UGJGdKydKuV1ePRAWnB3ZkpLzj4XvwbiPYClLa
vjs4rA6NTP6YEPwc/RZKHl3lQQL2CO4Ikl4ANy8R7qrPCiyXxHB2jOH3+pmiMSgJRY7l/PjG85yQ
hCplkgnWIK87d0hXdHJ5udxTI2wfpyi4KtMwbGjd8IlB6W4XSB0lULhxgCqNVD+Vq+KehGM8t1Xa
84ZucRTxbDmdVeTGM2d1ng3rbeiJ2bG8y1qCtgfDeieZKE/RiXV96/Sq1TUYj8yQ8S3hVn3822yc
oVE1iAOzO5Ql60lOkU7PWa5Fq6UKgeAym06bE8HUnWU6y9IA1voOyGWPMSELetphgYMJMa6SnSwF
bTbEEdLl1xYZ6EFwDnAkK5axvRyiFxghQjAKheGqdcn4EZ1+ZHDXIHqPIMXiqSZJHW0Y76WOnnum
DqT0Br74MAWsEcQjHf1hlRdQMgGOwX925Broc4BU5A9gqT4y700Cm7vq8kV4usCiJYullFFWDNDl
sGR9JDfllpFjj7NLyUFuAnNQrKS0t2uuOQLgHSExVHfzASMVw7tfzU0dswW/TYry6ZKj8pcE2ojG
SGOlbWINDu2e/xCkjOwksbbY9oR1t500+GEYHywfF8CBR4InxlR8ngowVvaxCLf3X5L4PjNBeIyZ
p2gIHKKXi9RL/5QwJLzy9i32M2BXnarM+IRy6KgXcUSHUv09q4kasF2jBtVR7MOTRVGuDYvUOGAx
WEstJXID196KKg5sT7aiJ4lU8nj33mI5YQ+yme0Iz1o/Of1nabPAxLKzWhKgUXzs+B2Y0qzxsvGM
Gx7qs2CbSdd6+9ELb8awGYHhAJdoXecjR8mqvFXfeuHkXwMlMiHoyRIU6hcYO59L//1UdYowIcAC
DR1vnaawTqKRSBJRgmKhGihukYLfPBjcxuido5oLvHtwD4E3Lp93uwIvs22bjHkLCY33ggRIi92P
GAflMvDA12oPBO4HG6B8R9GL9x+iKvAFjTFQxR6mRtVhYiacHk2pin6Wp9gSNQkShQOZUfqjFAFY
pjhVmoLmMui0KdK9VIhvOXo0UOYVwn1xa91opVVNXcruHyOwCfHNOqPKeVU+HmDZK/eaW10IwGt9
nRCRNmk+Ig9dS9SOZbSGIXDeXCp3Xvd6YfFo/ESQxHTU/TG6EH2vEOaUgTxR3oCUV5xR1ewhsIQX
oK6eaT2lvlA/u2hJp0mLZbv8AVvzhL9h9CIDK0soKtueGRfHGl1Cl+3SVZpWJPMEx7dJCoLPCvqi
Avep+MtSM/b4dWeWZsl3NWzQ0zWqwliGpYx/YwbRFsQq+jm+I1rkjvfb1s3P1aVOGeUEObZ34W+0
h6WvYB2/IhdL9Gf1G3/3N1tB5DJmQmqXSPv8cHqk/g+3zlhRt5eSlakGO/PQ6zwKtsHwkdTJtn83
EtS1NffJ5I3/b86zYbW8XCDA6sledsEYqJcTokBItLqLdD5G7afzieBqhy7igbSID6NhfEaoDjUN
NrTTNqTUopzxbtEDUSzSuJnECnbH/c+jOVJIouR7qg0T4Clj/NlEm3IskSVhW5skNEwINJYNxKj6
IN7cRdtWvdynQHhqCpIpUDnZEX6puWLtYMiRKan+94ivP0ybzr5dkp1rIeO8GaDxEUkwkleb4azr
GxduxtUH0oADyBB4Bb1fNTsuEIpecysLw64mVwWMp2M2MeWwoDuUFb2ojCYPkC5tHsH6l4oPO8hL
0wfhK00BWUrYe42WAci+tpQJaVKpERxvP3WSnyY7ALYNugyIlsz4WgCBhbac8nJ2TZrU8cplKmgN
0sJLI8Bt0PZ5XnN2Ph69ZoLf7Df6PlB4izxqxB5I0OXrPhfMbCuizj9UyszEyunkO2yrIeLbt4kn
XoYGYrV5b8g4HKWX2kjo7BFsPM8a8/tG3ABDSCXVYk84iLzf13076bHjgCaOMetyMeFeeLOgMxfY
OIr+OAqD/2FwLR5gLbAgBI1MpBZinlqgg0UNo+QT25vm8n+mQpWUlr2AzPw6oUUmnx0GxreKEOys
77+W9gTv1stasw4tBN3veS2TumjYxEWqckf4hma/dL3eZLtqoB1U5sKf0l9jCFvl0UR5AiWpcH96
IBMso4c/VQz/b/xH4+0L+T+cUc2b4o4wXM7OMEaizWzLvLLSyvsgETTeg7g441RIk2bbQ7LrBKN9
meKDBE6DU2G5JHDO0glpM1saNDuuaf6Q+2obq6SkPGRt+MwERrovXtvxt3Oo+JHDRyqPKJm1Tl6U
ltopxEMKv1wdUNy0cuEQOvhe7f+T8I5gGTwFmtfdGdDsDW6aBawIwsnvtnNnk7IiQ/DOyOlwwQGb
OuKtMmEhOFslZXA9sSnytpVCzLSs7ttQyyXNJ+pf2sribgToNcG6RRM4RXboBbrRDUazTwwq3eEJ
IR/LxT+84r2YLh3BtQmEPjNg6sjajWWyVGoYmq95KEybHsLfcOj+e+MolbmCGOgVQqzEYWhyzwz0
w5BY1EPhVAcIYW4gFQ7GhSfd/U1hAtc5tt/kPGhdL5dfJpHozbkhVairwIP/3VznhfWjLFY4s06p
lNgUIN2zupCDZ4lrB/yIu89cxDIS6q9zaslU/8RMRLtPRZjeXDTy+o70xo/wd730/fFbnumbaFK1
I2/Q/oE3RXjRU1ppzKYP3/9G0wCaBVF1I9cni0cz1cZUVZOn1WRUuZwQsUjg03ieN6W7E0fUPIoA
P4nHqROSnJQa+FNlHkK9mGqB3+ZjWC7uUM+OmQtk42h6rCzw0gl4CoeybEn4ZLBBTcTITR/6ESRT
KRYH2nCMQDawM8onQpi6oQPER4L0dOb4YSIJEcsx7/gYoyP5m1l65qZ71MvkkDRh0TA7DhkfLyph
wQD3je7YISkKu8F869aq7vQsYFIYYEBWA6SdctEzvoMNaCWnfZ+3hJxX/wdj2QmHQyLgJIZEclPw
mhrt10GpbhHrdVbRleM/plF8C9kghwYdH/yLNBhOLU3nRMq4SLPcROu/hDNXpD7McFC3PLpWVarv
up5SHwnErnWiq3Nfo6GFQQu8gmSAnaaUOR0BQZ6hHJuW1ngivY4/9B7ldwlTlHv9MPkFNCbKpj/i
Atv0dbbtd49GSUYB8YS4iZ/6PmRhyj/ddNzNsMCf6646wDznRZ5peUY2usbvN71g4K4oT6NlKSM0
CiSDA4ZV19pwo08tvOpInGv70Ds51SzsMWQ2I8q6pTS899ePfRQsWiEIbc/5vKngkjt4b/cQZryP
8wOxfevlRv7Y6qHjFYoJL7JVvPoaFERb2S2iII1rpJmX320zgo4q7L57/bdU3GzLOOCnUTvS9M9P
wRFq1rICI6LYKxEn1kWRyCOGhb6i48w7r+GndYPoUQh8LaD7Tbb/LG5SNBrpcTqNl8pcEOn/mc2I
6b5k8Q/td+MtSgqARX8asvumcgNM/GLZE/O7tARGiNKypKMi+qzOGLzgUYocT3em6UvYTXu5nHSJ
bLeGkkneWjpmUG7ml+SkECXjMudJ2wZbktPelLScFx2sQ3aROoDsa4s4NNL630fP+PjsAMlTKsko
Wk+bM84iS1yleabju+F4wy0WCKYibIHcYP/WQtR8t3nk1itOgai74E4j3jHbWq80OBiYIYz/Hud+
ny49DxT0gjsZ5MGwvEnJ3KzjoGYVBDZi44RmlMSzcuVFyGiCc5Jgt3pDNulL7PRB32qBFTQRurO5
rMOXRpm8O/rnSv5exa6eBThd64bN2SkzWmiwuayS/RV9o5XjeNdQhP05tbRYBkJj8pb/AZQSOC+c
E31wX4R37GR/YcqjnAXUl4/zAPTuuRVXwuBZuZOR63t7aqBbgvnjDv/urjzUNLEHLA5imNuUM1OP
okeDg1Jo5OblvOPbvgfoSNEfs1QsM2idaiRjMwDq6E452X5rNQLcHf/EeExWYsb9/kDiPUAHA+eG
ynHQ3pgbKZicJB/EDtyYddOBRVuPhS0vXA1mr2UZyeSynDvR6sjfX3fI6bdWqsH9Ne1xGyJtyXAd
AqEjZ5tQ9p9atQNsagKFUZ+NBN/0XU7pA93sYNxjRh+ytq9WTxCWL518FVZpDIdySOGOocQeFsxu
fCGW2YW5aJf046ZhrmICHyQ4Ups6gatjpT+y+sM4DqXHAaSaX330MTY1gelNxd9RVnzYsbgydwyi
sziPOxSZv7polcTfXIvLKbSEOXNDDuZdUowSQpKQ0G7rLb2Kq3lNSWq7ivuKcAdljidKs3y/JrbT
l4XUEtWVFXwZQ+fMyQRYFns0sTYtrjiTwsvB4rqDKdw36oVHntD6jUTdATan0fgIVgHu0KcBX5lW
hS7TJAUC7T7t4qdfePpiWecqV2bXMNZyPo7F0yk0psEglmC1AzLxIOT7BNCLRR9eJwY6T8uQwDO8
sXFjLQNHqRpWH5Rk9DVx/o3OmLCoa7pprgGrC5m4syA2AOgFKCfLB3//KJXXKA33RSoFd3d8IZxE
DJ5BK6w3LZkrAg99ZSc6IEZGpj1Bu88GXCfxSUow8KJIvODdQjCdMAlepkGBXFk61JFkrmI5po8j
DOwYXsk425VLSrQ5p4QWC61suMq8EuNzro0gm2kxHaJSpA7L8W1hCnqLyWnKO1W5wV4lF/CcTdy6
zVB8G+/J756alDgGwOeMr5tUbIaAZwj5LjCheRjdEEwSfaxSVXQ49EapObnrybIXt1yaMqe5R5yb
EVYLjy3zGi29HJUln476bgXHxdB+vGNY1JDH54S2CZ168oG7/XgUK19iuyVypaxf4pGeTH3GPMZx
vmua/jq41+ZnuvvOrn6Y683X0OfURTf8rsnvuSJsOdPSgtR6Im5f/+9Nfik7+zVsxd4PAj0Uz0tp
UVWJs7/kWyIy5aBjeXASHgDrtF0kLQsIR9u/UbasT9C5qsA+ulFbI+0JjBSaAmNuHjTBMqXQF9Iw
qKmZ4kD+BA/z5k833b197hITFULiisKONfILag4gCHtfXVk2adQ6EBU2icPWrPLu2K32OnKhfKm0
5e1FVDUx1fmnQK0NDg6HBhiIjVx9GMV8lfFmefPqyz24ju8bwQWR6yzE/vY5MmO6srUztmjoJJEQ
P5Yxq8MImikaZbtfk4aZ/duy7VGL8AOXMaO/cf0+V61LaeBwKP/qvNVTkXxgoyJCZZ50ID7qDjJa
79O4+cT5vOLqMDZBOXwLXDsiWQLHdpWvI+JGKL07ATUY465jKVH+fsulOFiD5jE8qPmJPgE9tJUp
j7hSIAHH6eL4RuFAssEapQnGHQUbST/w7AzfFNrf0i+aHCU+Zs2bH+R4mwlfrB1u+hgWLzarzUkJ
GGltyRTZ2BgXPONXYK1gbimPDowJMdped6zQjnHcDQZUdbfrR1n8hE6vYrSc6R2h/ns09Rqpmmhw
yvQJX7Ws0aKMH2aMHcNIm8szPT+QslCJqZkWQTOMapgTFAJLyteX5Vk65phlfql8tOZ3CbdkEBzd
ZSsDsVobQMz1/ExExnVdj14dG6FsdruFdHSgp9wT8cruhKOFaqjyZXu7yhdSggxdwfhSFn0Or2J/
iKcUgWnnHcLdBWnAh7bbcPcALB6NV91OSMzJll0e46DdAwWT5F+00+ZCnIfvcdHBxhJcEZLnB1p7
fLkZdBz5bFTw7HUOPUYAU7rJvib9Jl5aSe+HzuFxrhkzSKEJg12mx0QwU+04/T2zM8GvIcpwk6Bo
HZBo78tMyULuxUef+EaE20a/9RsgzUKQOjMvcvrT0iIcHonTthMNELJ64DxGSybMPpaVLNcNNA27
dglWCxHMEsJcYnF734ykDvwarfI4QEjsGV6TCvezfCDB7v7H3eAq9nbUgY1VZPvYPo7VTjBb+34/
QwpOMm3FmCkKbBRqJJf8mqF8RHxn9++8cBUlorOQK09UJr6i3aZ/Yx9zMQ0bpTYAuzmz9Uhd7O+O
dCeCj6IF/gykabyVku7cKy56XlCZLE9Dhfql3rXq4jXaEfViIf2LwBhrPNFeJ1BXAm5xHAR6X+6P
YZUEPF9rPHrCVjU/dufAJx9AWJj+HwIoVTlEcmu5kcDr6k7mrcKRXEeLWPYpdIQvWgibw+PSy9H9
J/aRKvSyPXlA5ztFCwBI7HwWukDSCLKByIDs7hBWISRotboLZpg7JpKSOR/oh7LYNPBxKr2l8w7b
hTE7p9+KbiG+hVWNvPrz/NcyvyVUVPeqHgccAh9gQsR9bD9tAWfxZ5uq72SNWoayeVcUWRfDDAWP
gJeyBlzzl3cuuxhxsJNpTuwN593M+lgql9WQXuCtBhBjya40CbvOa5X9E3drzPD7Sq7mJs0p2xW5
KwUnVumR7zdWJXHh8i0uSSyeItcwqSSkeI/49ZVaE72jJ/b+a/Wkkg8Y7+XKVjShk305x44Dt21n
NtClbMvzC2rUjMZaV6X7IRSTSe1G4r2vFUls5ZMOd3WoC2EVsijWgFqZBqU8/hGJ2bKGKd5bTUaR
QChZCgIxP+D0LeSVdiR3feQJS8XOEYTx/Lib8AfD0hydUBzXtxfz8y1znV2NItjScfc47xj2dlaZ
WwNVGGK9FQtJbOeu8QBbov6N4tF2piwqcBnR22xBxcH8fLdhtjbltN7k3P5yM1nCrSLDZhIfRIlD
qaTBFuJhHhDz6gpGJmwmVB5ShiL/hcwydD7p1jzZgO3AhWcrd7CsHT+kRGC4rn1xirPA8Be9mm3Y
ijgpfNyeg1xcCRxJiHX9wlWgssH/6fUMMiMLaD/fRPqqK5sPAzHcruCZ7eeFhAn1GKi3MLDhhoTW
leNU2X/KB6XITjQJowO7HCiA+TwjybLCzVSK8bLj6UZ2uRoo0Dff8VOwJ/HF2Jc5e6m1LOVYAlCC
nuQOQqCLjgo9APXFAZvedlriRxbl6cM1pYmDLz2SaJRyO6s2S+jgTLo30T8fpUeYdv7twfWR4Xen
G8O4nlpIVq8SXGZWF2tZu40RhhFI3I5vALGz+LBfNjy5rPMVkE/R4c6XAeh+930Je6LsS41odvq3
rIKMmOnRD3A/CESeKJY04DKoi0FMOoMeyzvdjh4na2Aw4j1LZ9MUMDUbbdmtFVrZdkUI3CPeqUH5
rENl5l9NLXBr+A9TREt1ukaeLpVVEM2lENuD/Y7os2zPmGBT67YzR5RZhGOWq18ollb52ZpucSqZ
ouG3Mz14RRn03bNkUm25zhL9IVRoRox2//1gqm4+DBK/O12ghfdazseP+1vxrjlDvhVGBAGX/03G
N+YTqxA8Uh2awqgReCLnCP6zQyYWBhSbloB5C7m2NvYRKsPBGmivh4rbuTlUFr2iUU7JfmX2wfIH
xC3CSJvs2los8Xo5vg0qnVCJz6pGbiUvyKLxJtmsrFBxO+XRJpWDaoGYdGo5SShKlIlHz+RdBrYF
i0J9R9q+vLp4bNgCoTFqU5JnuZUTlM/aXRa6+Z1s4rxcff/gwe5KrCsxPaXBTsPwNCPbiLBS0v9I
QLZRwG6OJLhDtKN9VORlpyQHhI2CTH1pLww+yK6YGwN4lqSip4AhFrvpcOBAgPu/cAMbV2SVm/2c
kxq/WIAtm/CVtBWofIFIR2rX0pxl6YsTZsMH3EXfgRXPsDVRr6v6RJXda8p9BokdzIeYDxbn2n/o
fQITPUl5+qSbEUnQBIbmWn0O4uah0b87Bzdjh+qRKgYhc3LO3pAZMiVsrnIhpqz7Az83H8xsZ/H3
XVCiCEUqYCe84bwCDMBg8rrX/7dLxibkKLXV6e483lFQZJlTFQKnk48EKY4K9vwhWfoCwDGaxYbR
ahDt6/ssDkMxm97IrJuq+q+29KUh5Q3ZROf89n58dsR0RByILMlLcGNn+sTj45XkJS0sKfrxEtTk
nfzb+MW8I88dEOK5A9fJn22FRLyQQzW95FHmKxfoWzdvedsxtjg2X4SubCD7oOHI1yGfIWI/aMCe
+UkoG1lZwbiQQ+geOjrww8r3V51Sa3GaNYFVwjnhmQZbyJi8A+rGGXxYls5ja2aaloYRVoUX0rBM
g11hVz2ornhsMomf8WUTrirYctv5zbNPakkZjBmYWduTbgfHa7UeShfHEgZj0kB8Yd3rUKvJ0Kdg
osFlRjlVxN19xstZdDrtJx9ZCP02usBurJrxpJVrp7n0VhJVFRv4GP7OpSJIdwPiIDHVczMMRxFI
A5DAvIU4QzxAm9hKDSpnM2/Oh+KDlu+JKoCSeufs5af+72hDAOmJQq24sxgLOxs3CSlrSiBRwLwG
petnJhMNt0FeSBOVyAZb8FkEZeW9RNU6p9R+8NBVlnRvDILGtYSJWyvonnLYwVMvKAeiplrDQylU
RlTBSwePSDkaCZi17JE4/Tz3Q1CO/fmmVc/X8lT0JFAatnKGPlSKA1/CS8ExNwbiZE1WUXO1TUmV
5PXrTQfs/7Hw5jeQcXS2/F9kDRJ6tCf/Brv5IPfft/4AJxOGtnoO4WeGSSBJR0ou+JnwOpV6dxEE
Iy+oQDyV/GcyE/nVdRM+EAlwwx/uNY3BG+eISHWjhqRp473+uTbYwJVkL575KkahBMBQcFamlPtj
B0OXh2ylvma1adfNZ5km96pJGoFgvYsrIZUjs/nwKptiZ6uIr0NbK8zRQwNKJnCPwf1qXVhBdsZC
NnbvsSk2claYHgOTh3qJ0qVrudyvbmA/60AmNbWk1cgbnPd8HTraew7eYFPzfcoGlMM7XGd7lagD
2U4CAJGkpoNGyimHfJyoso+1Z4edvTGHjgFxyiFJDj/VEkU05Pn9BC5gKBPGepQlIC2GSW1H7R4g
SmBWNbICluSSUSkOZUqcLSKEmcJhSYemyHET9gTouW4WeMaq1ORh3X+TuTzZLqHdJVh3fT+DTkTW
agZ/B1aiCD+z5morzu26pY6t6aiN1lknsoAQGUDDtuhZwSBs2/wcASZC3KUo34hepSdkkHEr+Yq1
A/mCDO4oPb6vyvAhARm7TUdJ2YeFFEAwfZl3WzZ88ijrRdcKmDqojbaBeNUy0QjNeJcKRQxxd3QZ
mv5iVYxDdOBXPIkn9O+95arK7cW2lO3xZrd15iY7wV4BaddqkB5y5bHUDtd6kpjF0jiABbmRupG1
jrDHSZ869Yq1AADHwstom9qyfrG/+AxENA5FCkrnRhyG7/WdQNlbsFTpuBPeQQRTq31cqbVQN65R
vPdN0g//F7CP/E7BmxkH/1hmEYRIj1z/w6dXxgWiYvY10R+RBWq4sjtS9XHY7WSszDyvE6fODE3c
9sFpBR/btrx8m5fjTlxQvIlm+HDLVEr5zLnXMaO+KogbOyWcwtQfukeeuDjPQy3f6F9B2buuEAAq
KIrDLCBW3a/oCJNanJTVgBYTH73I0B/QFe45z+yxLw55to8Y191B8Qe2Rjr/8u+9Dmfpv2suke1p
pOTHIR8PzKTdnWRMjke9y4p/L/KkkYbYG/EOme4RMh9PcI2qDJmvONOlyKt0funFCJg58ED3NNux
kvoQIuNFL8IqKbazV2VgZMcIvHKWISTamNAbIVbStEyb5KwhSOyJhITkisSksZa+MlRHCxtiILZS
+wMb6ooEH0kgwdKkpG/Sq0Md4AI3jontqNBWrUFxo5Okb41iyQeYFIcjVfqc+Dg6hKBhe/+2gebE
EvAUWMsr0gNAl9VTiyW8U7CyI2bQnOv4Gw588mxeOAN2PJYKUzudKB6r7ZD8k3v8WruS5+/Fcynj
IFo3DbAQXydXcCW4WvtopTu4j8p6F5JSxwNPHAXoyE2l8rR4qr/K+rA1j+WPB7JjGvQcYrVPb3ls
nkFETfoBr5dXsb0SNwBHtIytioBksku5ej90tH/6DQW0XnbbpUwwZpdr6H5E9QsV/V51ba/NRfCj
SU/J3K468RP1uT9TLKOwANYHKb8eCdwFkGpuhP/Sv4TfgKxREAvCZyLh21apdKqkjj1A8NFIvDBd
C8S7fX99G9mJVeqfTOyDpduIHrRs8CPHczZ+SkA/vMYbZ69z39yKouGjJFAvS4xZjWCBwf9ESSvG
b5svFSW6ukRHh64ySYWtUOHx38f5s/y3czHGSdKbQdnw1BMaluMB+CxW15z4GIUiVZwdXBIcTd3E
SQsNTaWx0am7v2oL3QUnRAptJdDqG47Rhk5obtpdxWfLpjbk3zKrWyugq4QFa0k+eftxWyt/Q/qa
jXMYyv93fH+ud9PmR1fPRk/nsviLSqPfX2KkTguptyKozOg/tt+oUKMYUqi4456bUWOoBYtjx/BT
pLhOvokVciiAWenEUTPiJy4amN64Zdorn96TbZ+1B1xM+H9r1X3igE+e8aj+e5UQaRr4ByTafLkx
YqdZLtJKkMgX8Bh7MlrbKfmcwMFoCf5psXgZZNen+TBnd2l67KlIef2SOi96uAlXmQITRzsiODmn
af/7BXhjvC/RTCK0iD9he1W0/2t+N1tDIITmT8csV1/140fl2L9LM4lZHIPch5kre27WYfy22eOZ
bEAg/CEwiwTK8s7UcK7aG2Je/7ZMJfAeEAtn2hXDaOQHm7hxJbFjhQL47pJTrloSm5FGyFHdVrsN
fOLrpe4urmx32Q4GO0IsCPVQR5iOR66odZ7UaoLjfRiXDUiPPySVdjLA3v+MaRKmaD7L3yPsEbkW
P4XQpvJIV343pxJJG4qX68FBKdRrV44w+6deEW3w2JGySqyESj0JNkIfGw2vDEKzyIp0CO6bMCdb
QIEeF1y2Vm4+N7mfDkh0dtIQOyKA2m1cyKASGMoH5uryx4lwCwFWnG38Db7MjiJPwfkGqq+1g9F/
mLltQ3ZjIgP/DESzqRo4TDSojA6lQ/Z/BZ4ghMvQn1xhrebNNUOSPnCxDvT9+Xb232aJlGggHgkw
mF/V2meA+yl2kA1TlwJXVnWKdpUKcTCZovmDWwVl0vrnF/ZIRyyG9sUBhLb9lo8wMnz0fFgjSUJl
bDWOlOU4RJ1g0oV5tZlCqFCWmqpEGKXOv9/CqaA6VMJXSOVXkXu9dn+BhyW+JYE9gLxNYHJcTHLT
2ndq215fSPr7zmDB7EEm8zHL+86V4YM6uMTDQErAuZ0TByLHEaJvZtvSH7BUw4oJA1Xliiqfb8CB
j3Zw8Q79smLcLPj6xNMX4Ps/9gcMT6UjJ46XqNwfoZqy4ilOlJlhb4h/sDrp6M7Hd3TgdhMLnQyx
5yOUBTko+LHAqtKVVP00Uor2gbH8c0DQxf851L1F1DgKlNNEmNrUEiOJ724oqk14D42fqNywL/Pc
IcRUYvaRn9MRkjXQIZqTeE1Ry9LoA1roXtbexcnbbeHBc6tplrMjDHfbP7RDtSWz5scIyFIjSk5a
/q7f7rTC+hHmRYaZZEoH0/5yD4WlnTapl99wl4y/GoWcqnr5VCncWKlWygkauA1Tu1l/EFAyFJLV
VoE8i8Lq0sh/iACaDW7ap/0icnGG3r83d1LC25QXIF1KnI6NhVZHC10Db1rhBd8njjztulyZxnb+
VbiZcYqLzMXicddpQGDWsdwnxSqZq2Q6Bs+3wAnm/jFbcDUrZKcR+rx3Vj8jgdfvsWrD2B2z9CQj
0JkBL1uYBnl8bqFsnxhjYZnzcWMmREhG6vAZvUr5lcnIiXX24Fw/wUYLJcrAqc3f9QO69hS5OJt8
QflDqIJWHabZX8UZ6ZH0QYZUH/phCguj5rfokBqTtmP7L6OHhNgq/u+3KnQ3liXX7f/dhzopv3xc
GFzEOcyltmf6AqP2ULjj5dRxsZKQPlM7No54XtxKCBCTFs558lS3GE9FzAnzYTx3So1mUM0hqFAM
9Npo6bx535t5Hkyk4Ng0EDWUL2LAiebbPVCxdhLQ6DKHuY1K++rCsZ/px46jAqfZ/PTSGWMMG70H
IdRXYkYHsgP/vI2FkVmvLwwr2EPsMfjsoiYfJqgDCIQiqphkLvPAI8NSBrkCYP47lBpcLVHzx3EQ
ysQ9Ad8sCojtbHNoXgphXFf9wIZorHKPmRHpeGnW2icZPepV27Vp+EYY86scQVmuU3vH9Vis8oyU
xVbeoLuWhuNBN+wplLBKwkgI220nsM70tsoC02d3m+ah+VtrMNcFQF1uVMeRS3UpT3220QDFYSPj
ds7hw8lcV5z63tsyBdVgigB53E7AR7t/TY4myGG1lR4o/a/jF1QJMwuP4HOFxLbJZyEd5cV/rV2Z
Qcww0l9TZ1hMw3i3SvX/V+nHXKcjX78RHWZ/cdu3yCS1dxHHtC5EPkqq0tyZHXldSrLx4mO4bAo8
fPHLCSRS8YpLv0cAKLNQJABpDTV0S0ug2y8sx5TOfxWOD7Hh0qeF7MqnVae6nQeoc5Qa72B40UMZ
kg2/HWCbUacEucS9X3Says3v66P+KIBe96IPDV6Rk9DsCh23oGYASLCvy7lOsDSkkEPIMj3DfHuH
xy2Yseajm3xUj3Oh24M6tEtGfPRYGjnu11qhrw+72+liyDYmgipzXsltNPsErERG1CecGMJ6Cm1U
4vquokP6s7lZa9GptPGXRluxpz6SUWtDEuzTrek3rRNkdqWkHiHrkZ12oUFXayjJTCqtA3qwEjv9
N1PF6WQkg1C8WuPSdhN8kIXxHFGEGPENqbDC4gUyqnzGqHbkmuD+Lz2sOiMOyxn1y19Rr5sRBQ3G
5gqXyA2dVfCellmAYwhIqNPh0VbuzO0+uL+enC4/l42MGV34tOAqhXHG/H4haQRx1mqui+g+EQz6
omc5+jnTBwj5ZGHgcvwE6XOkBas8sgs73OVi21vcvTM4rq6fNmicc6S7tGRZMCNWGTnWF4bOoVHQ
MYdBchdJKvxi7Qcl1rLzjMZ2E0I6bhOWMIHQwc0W2Uccjom33dzcy19ymy4QVVeTOLL0DA/PPWhp
oZeNBaf/GtPoHfpez02nRYd+IRHA/gJok+bqVw+2Pv68ld1WNGAvwHdrHDSCHwyDRYFKvMC9F0Rv
SeXwcs18sHIHnvR5J6X26VFxQKCBm16OoU15qrD/9hpdMJvEWQjn7WdSI/yybmOjTMHkr8fRoZvR
SyVd0B3iKhfoA4gVIEKdsggTKu+YZfoPh221Lnhu7Cw4KrBCf9gfYEn1p1lNiOjIs9BJhqEPfSs2
KYMCIEVnj7WNLAELe3Sz5Qo2JuTK3n4wJog68+s/COExl8CV5EDUIihiljU7FXhWzLAqLoHl0sMN
i3nEcqRuI9Sk6HWsp4pSRbWhxWmuKPeSuzhZSBlq+BnEKTxbIUlkuOClrR612Lmn1Vo6nxlfOvPC
9qy5G1hm6/AbKEL6LfA2sFmGYuLoAapYeaGdMJDMhNh7rYRKkShV7yxV6g/BlOvoc8pGkdJqIu6n
hRVyB1VEGnxqd0eslnEbyEWV8XbPJfu68TxuMaUGeQg/PT4qnUSntTVM+ZP/Bjr53iDxmBAPvtyw
uIeH7E7ErQcxzJ8v3FHM5n5fTn9E6fulX8zuQ+eHDczkTnSvRIAlcRRUbbePbCwWlt4v45UwK7GS
yG240qCsdEJgZUGKJ1w0i9V17aEkHkpVPY4GyholG9uo2tvFfAjSNEtkI/7X86Ru0Zs2pKCPOxgu
AtAQag7BWDTEW4vtVAycZesuIPePB+Pa9TH+GajrvUfN9+FJBR9hUg/vRTh475B8TAcxzQUcUtBr
ngj7D8gKlcioFIVoPemVqSCu/l5Zyslh8XDlVjEhaHVHUek5I6NxbdSUZARD4gaSHiU42yOd62Cx
JsTcwWCS942pU5TQiJnWqkPL59P8Odav68uz/zAafn1QzSlNivWi3q8Vhpe0P72KzHnqVhPAFoNx
Mb7NMSQO+jqLKYGdw2mbdEgBUe2leODfPRG05QQ/FAL0paXYASSAZajq2zXw8gVWyc94EwRH0SzK
GCy7cFkXYmHzBOHTM8KUZm38CQRNv0bpQ3vdRZmADVi1ADnQ0zh/LkY0W60EfHeSCyHEjOqNGXAW
hjSPCZFOdJ5hf2udNvyA8TbbH7Zu2lcrOU8UN7yb1bIYMByRr8c5zncyu1HRFARn6v1SMulfxdf/
cs9ThFb6NqSccH6XFuB4o5xcmwqPtvrKU7fwlwldEefAIJ45tirstS0mA3xst7/TxBdJvg2kWhwW
TvYRih4w80vOVvgBNtzRoDO1gOSW0ZNF+u+3ZOTrM/XQ7W7N3z5KdH1bF2p0LwWQ53/YG6AH30zq
tJrU00upNC0CHeGsWy6GvWHBChvxV/Xtrk/dRP6iodRyomw8B9A6bxqkRr44dP93/7lqtILi5/tl
r7l8rXKXgfob6kMbfFFObS8rdriSwSqLlisOo9etk2+kNqVgGxWvMeP+q0syRGL/odoRX+Te0wQw
d/cCvRGhBkon+1V0xyhQvi9npgmfZX2tcPfeMKhxZP/vdblUKgj/Ww2EJpSQcoTSHmQRq6qs00C8
7+1t3HttTK7/RN4DhvUZFUuFVyagloBQELU3B3WyyumrYcOKWvaHUXU5ipRhlKOCsLMrijIJqUns
spZzX2jRTS4pV2PKe8mKMmu6HCJtsSI+Gn0+p48KCUxNcXm1wDW4sibIKLbg/PH9xDbvcQ/Nu+NG
6I4l9qnEXHHMoRcT5T0qX8pklyqwTVi/ClRlyQ/hrU6fyof9lsiCv0kL0eMT7/e/w4YDGZSSKs4L
BMEDzDJMlNjKGMzXHXRWTyaPHhKkRjW8vr6chRNG9E/OgCkM0hqFBa0hj36B8gR3vWSQhxjLSr6O
SDlhpGKReQKfbO/T0e6af5EzliTTRXnlJOLjqQS+N2q3FZipiP9dAQl5rr+wOorKsv7KAmX1dt1k
fU0WGWuti9q5MX2N5Skb9AwCXGmqWCe1P/cuT+i4SjtKbJYD+mC0v4XtFT6B4dKbXkgi1xYObHro
qSLl9h+qtKWPAihs33CrVk9JloGEX0Vyg6UjIyutmDwSMzTbHqc593QbmID5T65puIHIkcRbMIn9
CK/ay7CSA1hxMe2rJsewMAAunq6XzEei9/Nge9rLkUevmLZtANBy64DctcZpp1Bi+TvN6RHm32tQ
eYAxKN787G/gOeiylDnjvU+WMy7h2PCFxH7+8/uTPZgwPIEzSIfpUnj3/zliFNPDY+/Fc1sBd1h4
GfgTui8UnpkNpbrMk+ALv0tB5jnSgfq8xWRB8YsY2UCtVnVNbX0s0UhNyw8aMK2pz/5bQdNsiAvV
bYoc3Cyh5XKete4JF1USMKP0ra9yLO6K3PqGC9f3PSmh8OgB4NjKsqv7o8lNg/Uxo22gY8r6F2Fb
HAVaU30FLzXp8qVqc7pgM1MeL1e7ChoTDztC2YK5b2Nyqos5eN4jj95+xswN7BsgXTJP4+5mGeCC
V3Iq5K+yMQiVEbQGBqRU6GZFYfpEzQXAEHgqe/M2tBn/OJtHfFyHYUMO5t0pjshrQAyTC7dH7yNj
U8vI2sGbVhY+pSLgGT1P/N8GOf6/H84lv93n+rPug2PtliuFH9XqLDHbQKqtaSjZoQh8Bkqp2ppp
mMC0SS40KZM+/a7+n9SqBIlAa2JuBXgz9efrOp5zFgXuj6l2pvS/yG4DrSgJDuQPNBJIkYPanK7W
+CE9saipcVjcswsGzzILdl2yKG4u+kLvomKa/zPaGPR0O5LFbdhUdW2jOXB1RZMX/O6U+u5YkCBb
01IOyi6LH5yftn3fjqt0vXOj/lPZw6yr16yi1uoqRUdW5KnDAlsuHBMFoGN3xB6f7bgR871Ceyww
kCFPcvrk+GH5o/KmEowi9eln4KJWhrhsX0aUPypkC6IIC2BB4VYSr30xzWBIk1OJuszsNSUM6DkD
8Yz64xpSfqL7QZsOUlYn0102qWmi/p0HnlcwNkFgxGqf5nikYXeijPIrD2rZIF7FqAXB+wH0KMKw
e3R9AZutIr0Jz2fm88ebJkNSofiIjM4hZJJUfbo96GyGrzSnr0q0Z8VnKwqapo5Buh1q9cZfajhy
ZYaBmqIKK3DbT4RoIguCGjo6to7g1bpTy9mdmpMMbnQptTeiKlvbz4NExnhNVbwHfpEVK3Z8jgHY
AwTaTGsZRaAyv3BxE0ZSXazIjNLqE9gz5nMXVuhGoHiCiFUNfOb8ONwceFMOVC5vBYBDcMfIxEZy
FkKbpKyHwKP4KclMaWx46waKigLHi2yeLOFlTlC6AcWMFLTttMm6Se2eGDO8Lt8F2Mq3C+cY7fcj
V3FnFMz+4VXN2LqLbOaxX6h/JP7bVN0sKasxDCJ8EN20sEdt7gQtIPiTpFjMI164VpPqFDZAEK70
NnYHZxqlHTlz8NiAahkPPjO8qL4tkRPKtRs7nsHzpD/ocuyGVFXeNSGF81U3p2R9Q/Tppyxufzy6
4lL14QsVR8IMlsIRsX68AyNT6YZQ+0Oq+aTaZO2jFHDv43MzXpCe05RHN08jXx+XNvuP/vUgv51s
xOL2dfN9m5nz9J0VcsecjZisYKfY/LEx9mReZeCiix0M4xHIrmFsSZl9/Q9PISVXIq6N/KZVNyTJ
CkBTphIKdMKelNCF2Xtl92ALFRJ5vxaIRi1/pcV+4CUsB0sMy7nkXJWbL2BZjqkiDNHMrOBV3WLG
YOkkwlSz1YvYlDKXOBUdvWeXhTDVAyCnvOIxwAO6Kq05QS84kbqC0YYyukwkvbJgqdVw/GiQEboT
OuBbK9NQ+TRFaoNh+BwD8C+hY6hq9F8CsGNGaaLoc+aDr/3NdQIJB1BjBfRlkKQKlTR+Qk2kDjmE
lVm7T7JgmguNUsjmFBvL04pYn2j8T+cXB1fYSp3KWZawq4FflzgbeHJ7qV2W1yXtq2t8fJtE4jKl
eXD1z/+vzNvHaP25pT96QS0PmNpwOSFKOjO/1E0SwZMPaQy+N2cbE9dOviV0w2BLA+aoUNbjkh1k
ZDrXD0uREypnKrjP8xy1Ymh0OPZ4mYoQzRmw5U95qJBAf4PVTwzPxEa/X4okjNk+mK17/VmwXStl
4291eBbQgWyj+3SYQ8kjYn8V6PFL+/ocgmF4Fz1tVcMGz94W0NTZNjL9KasHRg5elJe9LUgm108O
bze0noeLDLHZv766bBAVaQWpfjUPEH+WpnUmeXNXrfanN0j1HIsg/2YkphWE4EllPVG39LzujzlC
Q9w1GmM4BE8nO/N3vxed28taZfQ87WNgr5vgcqEI6XIfgcakTxRsSasAVRPOoIGR7pyJ9XBwVjot
quPIdayqDmDiIM+rlntIOArnZ2ooY6bQ5cFXseZjm5D9nPRrUamdSOGAxqMUlTL5cLTZzjMn8zFB
fN07c6UuGrHnOEcJSzqhvfpKH3y9pgX2S3z7nydW1B6830ZaFVEFVs6DGvLufc/VcDuifp4elROr
3qjo9aslpZWi2QtELB/5B87xQr+SM0bAr5G+pFaONHIPNXaJJksBM1ETlIFkR2Q5zmt+56L0gvHe
fLkOB6LL8vW8dI7/JNU/UdWeK88ybhBrXS8vP63vktu0d4n2o1ZGCi7XCLHrMRHvaS1RIBFCAqTN
jxWsZxD5KC+8KHoOzbtqWPX1nolgfAIkRkgvu57Fj4b+/b4tGhdq2eQPua8LHWZHLBbE6g3M4+Dn
keMBkrfMD/pw40boZTDZQyhx9ITh/gGj+ii9KB75aDC5iYGKRhLcDuhrFa71nhIzqVujTw4+IdYN
6e5iLCmTR2rHp9A4eT4taUaI4aGGoZvEevecWmC1GTZ4p+zHFeXBSYnBBFHhEgJOkpPeNANI9kZC
O8J780WU3PcCXVzVDvINPY2kBprJ6l6RKjf0hKGfsc6flJQSqkvP9NFqDaqL4HGhHdn0CtZfd4Z/
Is6HWo7ImX3GI1vVkCxyhKerXJaf44MpcIswjJ0EIS+GDcySjwKQ0PT6/QXYReFrjxJiF6NaUacU
Q0hjW/+GW2sMZND9NvK81Nu27Svd5EslGvz3FvBV3oPHUv2C+NaL5DJsgrKbp/Zk5UZl2W6tII+Q
9JzoRypefE4gaZr2+rJcAiivZcyPLpSM166ND2Wp2SXbvyJ6ZeqKEV32gPRZ+xWO4MA6NUErUo6V
t0Ob5kvMpmeEqpAAJYVreOk231lES3xVjTn4j4n4D/AhlEUoQ3KndmmdYmxxhvCSr92AGanPy3Uh
yjNqhCeAODxkdc+FPqDe99FpWmrsVTBghuT6YBRNsWrEhsJJiJIUZANK8w8Dh2hM3Zvj8INbWZy8
vwkBGwPZ+Flfoqx7hIt9n29MWlCp5wxu9uisHxMqWqJiyKEhmychUdL05tc2uqn/rhjtiXLYaUg+
NyJwAmi32rgGJLcRrO4+7ADu7xfsT8KHf9UGj6JpEGyBMjgu4mhnKDZXJTYrnWAxs4XcNK2ALpVn
awzOJD9+BZw11xpGWr2SdCaNIBdvtHclT13kL6zAq+++yjnVZy7dGigJzAWP7++CDqarlH/6o/Qf
aaxMt6iftxtAnBm2UQEWLWPwVB+OYAIkFluSMOlUwWWRNjbdWFSVQdRGc2zJdtlPb4TjHk2M5vT8
K7+XqiRke4pL1CsKxSgm/MRkVLgbOPq+kfooQkcKSM/B2jEaSbfphb3wETDSolrEU1MKrsVPCBON
aNtxCHQ7BL9exAboCZ4XZmQSwFC2m1m7C9zo3A5VRHHByIqgjbzbsh2aNTQTYLKDy/hzn3jxl0da
Ol5G3a8i5UcYCgpfqoHF8cjkB2LHi+Dcicu0Y1fFfc0JTrWYCiVsFCh7kMGkHqNwLpfnRYeFjf0j
xicxHatTlkNF74tlxYAwyISkattOLLq6sj6JJaVkYx5TSNYqfeSKPsPrIUzv7NxAosINSNvGMi7j
6ZB2sUDDeFlNLDeoPm80eEsVwdKPcFwO4n557SepvB4xLAjny6xgf+9wEZPv2zI6uvCvIKA4Ev1V
faS3cBi1vqWaI/nXmQ3CtK6r91vFtoiufvoVqYFb21GcVi4FoPZGiYqmsdUWGRUtEdvKzARINyoM
ntO6VAVqz9voGVJoyjiC+cy3JN82Z/QcjNZ6H4fm13BcnHN4UIimn/JFfVmHtPva3mxPeazjodNq
zEqGr+UijyCQFmNFS7Lv9LjGMj12NWLrTPf7dVG3rFadhbyLtAAia+7ZcLzpOlMoj/MYiNyEO0Hy
pYa95gNZZsRIsFeAGAYjaRHuUKSr55BMI62Vpvjdk/ZxvuC0oP/5IECwWfoQ3W901iqGcTMDKIdL
jTIeTHH7ycFO2YbJUXgC3Arl0QvMpU03Y65kH2CJIVZKnfRJjba+eolt1w13cd5BdDqyj6GHZmuf
fnzhEZvBg6QEfaF3nGq3ZFdaGfBzqfq2mWtS2PSl62kmoBVOX4QFdUFzSDtWpo/EC8eXQBpUNAfD
x1QPqmgoaI5r6h3lz8PpI26kwD9fVlSCzHveJi7BBrPbYuFPShICxZfQSk+kKkA68reIe590bbio
vxsX34wMYbdfxuzaQZNlK4FyzLttfAEO6E0MtDlyWLCgfcXW/K2Wx+c+T85RQ/08UytDnwXq0Yca
34U4G/bjIY+KHg75x8CIiskejjnol2VivzdOmfp8slV6GQFGh+/JfiPwj0gozHfP1F9H+1Xa9UOx
kYXcNvtUzbZ+vQlMeFeMU0G1F+4Cj3SsJQscMv3uD1ZQ7qQCYe6b4VV44b8ni9MxH2SSYPiIEvZ8
wOXSN+vSzt5d41AWrPY4EPHSu92x7acuyIjTIXQHs73WJO+IcUzgiRuP9vpJQWEYf77dBhip90IP
g3Bc5FttZ+HqUgD+9wjeNnR3q17/3x0eG9u+TeszA1fQzVv+z4DIWXehtYAbYLhbwKABMXHFXCm2
DDIPYhiAz7rkochqu1rTIL+5D9FuDZnaY4cVIuvzcSnvm0VdLnHaMAcNNEsaL+9o6C0POlzA/A4V
w5BVyc/MFYkKmwnORa85EdWQWEaGrfHxP6XVnHvGIFd6oTzI5KSbQ1AWKDGIRUZMjWytc+qWDxBD
pc8uN+xfYF7U5j4CBAs7kzfSAEVysy8hv6OhYUNRGGgZyVI7RJRdl9HMfaICzfzwuNbiV4QAjF8V
QN/li90HmT3nazNYm3tDvG+NTVldDZxaFQZK3y9W2ukb/TQAAXp0dbb9n9w3LUj1UU2GnuHisbdQ
PyZmJBsG4mUtz8M7TDq77Gyf1T66ArvQ4J8IltzSeGTBfaezIRkVNGucoW5kgAxLqVahJkPF8fB2
23FqE4iOt0PrgfbP5+37lPeH1ctJqZK2QxciQpa6aTfEyQxNBhY2E98SkyNLObLkw6TA9saAIx58
pytF/lX8WKotilA+f6BCG0b4e9qEY3tqgvOh9WNO7975QAsGWj2drDcRdv0PO9vAfLyKZXI4DLVr
+dUJRbkDiYEglbJIk9U5TRbKqag4VlqxkuCIok1tqq8BgJ/cYZXXyzfc4PtF0pqy1NsyiDi9lcJE
XQqPB9sIPL1EWEqX0eyKl2hntrdEWQEZpXUXn3VLRltco7AoGE6KrkIW0psN7Q72kUKVoM7G7XRD
LaXLyibkh6ZQiLFLyd3dt6Uh2tPR50tbd8BXsu2YHPUKkdL9WFY9g0K+i/hi7Q0ODxlcnjNJmkCD
D7AxlIet6K+ktao01NlPrDvKEHxrkKg8L5SX6Mqb9KyTAK92xFKDaZ3n0eczoU+gIcQSDuN69YXh
sj9RzcsQAWgJ/Jf1KpzJN/UPFqvVAQ1Ssu1m9ppo9PyXXZMP/oTsDtRr/6x6vN5wwuOOoBrn4FDM
F08Fm71/swizdu3rRv2P3td/2BgnR/29Fe78eCLNA8g3THoQM5xGPZLOvTJap70kP2DCtLoV2z8m
F82XOmrXcks69GY1v3r6cemVOJHiBGDs/nPhExs+o1JAuL8zdHsNDz7cy3VMj+mrTrCLm3XYu+gJ
1oaQkF5frgOI+L5zap+ZCqKno01qYUAs07YJtz8v0KaBB7hrT8YK2zEDkHfcenRMcJlBbB7G0UGZ
IHKV/dZ4xz6ebzm6GV2VmwHYsOhfpuoRsNE1V4Kx64bJxYqz6fUodpdAW7RAlH+L2S3iH+KPJVGs
uoCum8McD9G1QI4BdpEUNqyC+6gUMwqtb/9VVGWs928QvSpMVH2H5Uf0Iy9h8qh0m3vGpVeyE9RD
N1P6osNg1eUZD4dwqa1jfmf3UdoGQiWmPcbpofYT5Sm3dghK/O0WUEi7P0fnYYvgQktzYh2TNmzA
6/sR2AMRZCgvF2zfFSSupuK4wKLa9EvZPC9/Za2PmgG0DHIsqi+rKqM33RAtobnCnD6pgBNPC7Vo
kGLl/vemE/0Wy+WbYhvcdiuPp0vwjqRTtkYtzajleJm+2g4xYGznBTXQXpzTat5+XsrWA2PsWvZr
wK2oWznu+76nO8eCUXLV17jlu5MK2SWnZeNSXYEw6axOiNfOuzelmDFm7rCzSXC5IUXb6Wkm2PkQ
zvixG7vrUhxXnblxLGLYw85rJ7Cn0ZdfHmfJgkTFtgD0wXfPE6bZkk0kktcB2JyRPB2Qoe1B+Hh9
Jjy1iqenDFjE0sYw7wKpPrBowmcjAxGvGGv7aarRhHynfmDvrwxSj4OMZtA0woH2egnoj+FN3dUE
RSuF32A37lUeeGBgVmWnQC3hSyXHSBJZaZW0CkrdxyCJ5+juT3NUVdQhRd7yW/XkYVgSbbmp9bAs
ob6rmyJdKclYsbjbwEIs6ngjsKSM3xk7nkuXSjxXVHDvXyzaZkMvArMz8Tw45/Won1umfmvHSnSe
I2Hv6ZROrYdXGmitI3FjMMlYqrR6gWGHuSOgwhsQN1uypcYrUgEiXJ8TsHMhMvSztbjxW3pgXUXV
38liSP5G0z5Z9KbEfvXT9C3Vl1xndh8vxFkVYJ6DaQseqOrz9M0757xdhENZWnWfmLbBADudSEne
iQOo3pLZaXze0HooC806/gBBupRxb1gBRtqVCHWuaWOlEtgzLQHGBTtPVh1MXN+A1Bhm3jFKUCDE
w/XE09Rm255482oA8I7BLflhSjmYnN0Mj/tV2hBQkj1hjnRhiGa0/49kMnQtcsqge84VAJSMc0pu
H3Gr8d/1acInWxkSF9A8m4e2KU3sJ+u1E5ujA/4qq0GbBMUU4Mzqknj+6n5nNs/xsDrNdcfw80FP
CqztHjRQupOumR82ENlpVWHdTgXTJbGuvgUJdF48BrL8Jmmm9cYO+9h+1MGsp5eqMzdo5jIAwFlS
Su+YmGj4SYzwssQc7JwKVZPY5VkJk1sCVxrBDO3tSCAkPBN4VPHj8ltaNJGzbEewoXu2k94iK7wt
YhDedkMj6W/vhHjn54z7Suais3rqBYnOa9/HgEuX2VmtfFIa2uZ/TzTatIhpDkgByW1LTIBArG+z
+fi0YxkKiOFSS3ApdK3GMqTQzh3Ri55HujMO6c/ghSMkJezlN4f23vOzlQH3cB9BSVAVBJxlcy8+
cX719TuZp3X5Rtp2egiTtSv1Qfco5PqdE6NErBV2pG52mCYf0DOA5kaw3/EraOwC5nNSsFnFNj/X
7dUzc/W8XZtJ7UgzUUTAKVvKjwjjdEG07Qa7vnM1ITUhiN4G5+wsRvIeOV8gghfU4LYbIUHs6NL0
3FrrhSfjBeOD+xzLzYDLFlWlzzW6kvWEH9In1e9j1SPHui9IopgveT9QcpXMBWYeb/4wXX4u99AX
AHCyiQPgk3wd30nxycPGgHMw8tgAA5casohON9YreLbOxkBrr+AeKorJOwlmqWO3ppe9ZvgcPKun
c/0LpvQEgHGVMHi1+FsrTprAKUxc6yyfSDnY6HBfbTq78A0vMjTK70gnwgTdWCEbR5gU3CW/gNOF
0Sg7fDsrTNM5/X+UeyO5UimdZgJnlIwtVRM/f3Nuf7mBnf5QoioxgaTBS0PTBjJ8nn13ItCyQU36
rdQ5UIc6U5R+O67Xzu+6UYDoQGYoqXz1AU4cTHFtzFz/B0nsMeFW8J2fdCTAuAXSzZx5Zs/SM+Ot
JvzvvC/2wq0Jf1ir/h5SG9GKTUn2BXOXn+t93fL0d6KeLahQt2t7qjJbUgibUJlzqdUsAVQZGZmS
jNeTqsc7Zv+hSpBAtWnvveXxIkg/r4fvQiC+vGPjIS5d721pwafxItw9G9xJIJMEyRYgvsi7T69w
QiUTnEp1fCBux9hQu2d3yjKapxuVRaLEeqTsX9uerjS43fIP++ZU83ZPoaJdwzbqpoBPKwZ0QF6W
zkpBkhaOkTcrHi+w9E8PvwG5G45Ke+pnmQ/8GvAFZr9SKu1paOs6YbhDukOjI142iqFmg21u9+Hz
plKS/HynbaiYJyiRPsjPsbst619ZEeOWEfK4TQ+H6JgwQ7VpTL9pWAF0Xa4BLL9k/9haJJ2Pna8Z
8zTCSAYIdYxgN1N2VBpUzmOsMz6xiikA7poULcqP/II6S80yqqNxga2idVR8oL1mE2RicibW68ga
I/Q+0iaHNCBY0Y3LnCiev6ty6iLdGEOTac2GI56dIKZrfNSeU19UMeJ018Tk4Wn3chin/6PTpxw2
3qXBDC+zT/XWJNlIOFRhFZFyygAfk388gXyge0/pZ01BqwU4IvZ3dg2RQjthuoYuEtWThl2jEhCu
m9GRDOLjlRLCJPT70Femak48UaHq3ReeWvp8oX/ePEEF+ozUugiWZFW7JdLIo4fv7jAfrxU4kOSu
1JqwfITX1ezvxxg5Y+nfd60y5LEEN3caxoU47QRU80Mp728a46Dyegq+/ZbnDCifBzNtwjdzLeW7
W0URXT8TXmulSRWESzBmD2PB5rjU/SHFX1rPP0ZtdFFr8RD8EM7JpYHrGmM+LsreFlqUxYx++lpI
kjIyr+GpWAoBOBJNLBXCUZgLH3ZqTwRlNXSvfmO5bRavK4U05zHeJB16YFhUuPqBtemsxbZDSivw
9TfqIN+Bobde2BRGbmNT7YX0z1slso9n9YA/Sz+EupCJE4wrR9coiAVoJ0WEHBYPHLR7UA6VUCjr
iyryJAAnO8HAhHLvOpwauF86wII50sIu6Sj1+hg6O98TPC4yYJUxv8yByXjGqrqu7mAWTC7oo6rr
Gn4oGm6Vb6y6WQf987TjXJ3DJqVl3hAQFJOCq3rw4yhay2SnJjP/x5lxkL4kMSQumUggWZkAdhHz
TBisnR/MVFlYESIukrQHrSSJ0/x7khVMBQrpjbWg7E960PMZ5Wc64muqAsfYTnCEZnJwAWPn33o2
baeb8ee7Ff502W5WHLg16UJ5QZ6REcZuQ2WWIuCrv87NYPZep6JTgjWEmpij8NZYz44lE1joBxi4
Sff5bfXspELj0GilYAPiNZN8Pdcr6McB41MV8tfrp+zOWaJSMuurzVcmNf9B7sGzJq8u2N6E05w2
TCcL9EiEaXAExA2pHwN+XJwOm+L7MAHD6PfmUcVCPsabilgPwZJ+KowkPyZ8IdlpNutObdc34ye7
pgnt/432Ya1wQsuwW+maJq/7dOIfrpsQzMxJ8N12ZraURqqLOQIemgXYJalgxDxah7/jH1U4reLa
wJvipOse4Ff1s4BA1GR/aZKvbp1lrqEF7+p2AAk+nzZK9cNhWPL7Rqk5MQTtAQzx8Wv8tvincrMy
v6DLcg7LFrXh3piXQJWG+L2NgK4yMg/nGL1jQQeTfCi8Zyt7QKFD7ukPEYRvzxVbKf1CVPMu7eXp
rhb2TrCqip1vBod84nmEPuMQt9f2qoZviVYID02sTp+tBoXbmhx2fyJnjXhK8aJ2bu0vYyuIGwud
2BGGTbnoaSox+q3E9Nbnsab2Pz82gQ5LOxbexWhpq6MfG2814oXrrTZ0tDTisGs2YwasnuDbKziB
9dlxFWDeesRUecyIpuupeaFqKKT2MLKaghdHowykEYoYn0v+Zldh8T7nSnY56xEU4ST8J2QPRYeU
9hX+CmHBWpwZ8xXONPp1CyBTB3WejFfjnj+I9QBN85X+GSMRjzU2Z9jLEsGQddMmrLKDOqWyOR2L
aukHUOekUUkenl0lUE7voPXvL9TX9wWXbT3L1je5E9egm9HwDCK3/qMJ6Wez7XmdAim6btcjfkUf
v7W2nFXfxDFw0Cg+2gxBeAgwxt6xIMohVQQM8uATob/JVVm0Pth5ZWCAt8yNT8TKOAYE1bpCg0TD
xKRyU8Awy7cy9BWPwRGsAZqpSJlNk8/AtPeiMsgtv31D2Pvbrn1nWZmBbTEWyOVK91fOHTBjrX5d
eOTxdT1LdjP6RZjbZG8niEz2cwvyM+h/QpXGmeaykjfJTTwHyDvNyaojm+W8DDLFk8Flu0TXgtQE
x/3V1uyBL7TqL8VA6eaopxIs3JUWDmBSaX/GuYnNc7n4CEWr34DfX95MPZDJkyoBl7Sq/G1ILUn8
8uipHJrGH/jv4EQ/3WtFg/gatfgkO+IpC6bjP0feFM41JXnazkFe3V2a31HRnODyJe12j8RCzEAU
yHp2FnqA9L2kwmJrTJe3hQH00dmJnHQjjDhanU4Ru2mhIn2l6b8hyuaGsan4g2z44qMg8QOiHGOX
YNwJ+wp1W+TX/9ptqfQ6oj55Ywv/ZchTtUInjulYLckv7Drk5GeniEMC/J84Y8MEssE8EEr213n3
hcHNtOzO5WuS8boYX2WpvHOJjKk+Mdz0mHHPXRVIDCFFf4rn9+TMVGl1UowtT+XntcOC9ZqapH4v
5GzjFC8+k+Y1eGGbisbqYWJ8IVAjOwyWYw6diXURqDjeSSlU7fUgdO9bo6aLipjnGGE6Om2VtgWx
u7la9hqxwWn04yPi05haVkloBp8nH4gKTr/YJQB5NG3ewYv6y54P382VOWSRNjA3zSP/yY3Bfoym
Dx2dKyEmoaL+qpj67ZlUEFQNIccbpxRU+9nfwALZuA7vK/BgGIV9Pc5r2hJ+rW4cYZh0PkS7BXWW
bB0ZtDufsErm+nhEJ4lWBRxo43bDzRaXQwg95EZzoDLgM4gZLWRwIIOaE3x7LDzl//+NYZxBx80Z
ogdKl0/QNoOFVrn/KeNIMhfIicf8Goqqw728quLetNIweKFTdJn6LTI7DbCEFd5d+v6/VoNWeQjK
OpJWPcoIXA6Cl5zwFwUqsr/tZWNJqSdB4+2V0TO/dcAthLsgbhOobAuGqWjS6G8mEoP1u6eDoaGj
d77YtwLKrJd6g21oH+aZIeGMDlAY7Y23oaUQoN1olQF6qoh1G2OUZ/c1zvB95NEbLLKSWePMUxYa
jshDo5AbVDKB7CKt2AiySUzUHKKWwO++fv/mkfz8NmDWLhtja65jVnvKUJPgTSD5oy9thHkwUoTi
5lEgXx4nmKBzsFpdsOhQIwHbVwrC6L9frWWUFXgS3BI79C0nDOtDXrwyABsgV4/6VyGnN7pg88/d
e908/+OXHUk9elzs7fnNbNj0p42GEs59DmyUGlt92Ne1SywS3NAuaW5UllWR8AgZmqvdPJjAURxd
LzzI9XlnowlUALuqsHhpV7s/pokhHIO1JKeB8RjX7pPKDGKR0EwBdMTzjbzZVrwlHcDr4E+UFLHn
ryfZR+ip7CXcOHIgDFsWfSlCuze0UlDgBLL+p4WeLFk8bmdfwh/w9FLWLgUYfAbfMgW+N00DeCqE
ST+54lTmc4cBxVMgPK1h3QTpMSS6yIzQRPp/QbK/ndWhAz7cnYm7ofeAVBLJMjb6g9s2IdOlOYCf
osArYv2BCmK5FG7uPfQazlG73KifxYet91N58Mv4+VZGN326BxIiv/Vni58LriEP/BG9YolPF07X
lovR61eTyEw0d0AGC1fSm55dd49Q6v/8SGUq49BjaL9nfb3uPWPOP46eyPTv8F+tMm060kEdpJ4E
FlXV80tfisDRB9HnNU/hTSKsQXZhYhegvCWcsirnHPaEFNgx7Wv4RdLufUylGCVb7gbN990J7sLq
e5po1NqzKMBBoYZuPcjeZOHeJHHupvCb2QSpUjtJKxbnutR5w0ETCSycVdfbOywxpBV0eCPoGiR6
k2vAEaWzcsP8+KfehGyp27A4XyTAHRiJOaU+h5+CQkO4ofpCKcQP9O3xG5G6KDM5a0eRMfOWenoo
UEZ7selBG4o+QDm6Nf8MEE2aIt6su7gNxek/tYLhdc9abu9HvcSdUckBvoKiPRABt2RvgW+fb8GW
11Ph+xd5oZMTt99k/++/Wet/HluSJI0q/NDbkaT834xZ3NaATB7xHWH3fO2ym0GaaFwEkwp+T10k
UCq1L+qEMlH4HkH2mz2wvepygQB/yXWhEP750gFZbllm9J48zjIGogZod19bpstlr68Ypvsr64VG
EVL0/IEPdoDuGfiOZvC2vE1BgwJxuAtmrPZcfsIqMPRk9oJY16tkmlyBShnUVVIytXFAsGQ5pAR2
YPmkLJHUbfQp/gfP0PksqiSSZGFvnp+gtMiC25ZdL3WzXB1TxR+tmOAym9f/ij36AdjP4wQC28qf
uvX/BHTFydiFZRjiWIdr8Z8t4Hp70Nvc4fEa/WllmguKmEBq9NljlcYMar6InWJgsKPvtBMAEbZ+
5gjvQqR2NxzOm4D6uvUmiWXjqxK0B1coG14k5AgZEqjaEAlLrPFRI6JvGiWizj0UdZSFgxIxw07h
M4RJhaimcsvnCyw5ekFNmBcKxMgqTr/d8VpFGyMQ/hYhZUMV8X0iyqtVCvfvxhbvMxFd+9YqMQ2l
N0PQmJBIPyHyXqmcwhNeESHtvScFZWDLoqTLPnsWt5lRn1x+lKe837tvYGA37vA1Vl9G7fxeUNU6
bJTtil5MIud3M+0MuhJmiApfRBvr1ZKMrOjCIyNaeyrYBTx/KinztWe5JBl3R9pdEnh3VDl0kpBY
Pk2KMoNpyhyVN01V/IllOv61J9IlQQBro5RYxGo2AmH2+ytdEsHv545haISqX5jJg732qSPwZshj
MBFq0PuM1tg54msYru/cM/kCwfo9+uV2B3sdHSPmxLBQyTnAGVptmKddy+8186JpMffoClF2ae4s
ZiZz7TXbC/1/iHqDk7bRrgUquXv4khjvrNn1odYS6VEZhBWKvEJAECfiOd9SvpLXRMIQHD3K03KA
pnv/RdTXZHEgqcD3lUwuzU1smkHeV+U+aW0uRB0w6SPVT00bAJh5t5CPaCtd3xVJTX23uCJHfzZ6
//TglYYHAIfnVXL03CNJpQSvLRwuwgqPtupVDFMG6yi9rvDvJExmQMFsSDi/84eDrwbTXxj8IjFd
N7hl0v2jXgKdb9x5M1qsJlwLdlT/sQ66itFMm1vFckX6FV4WABzBsYFX2XXfQChOHBJZYjEZrvGK
9mv+z1FevGf/dObwoe44GzRmOdcY6gdzXBpdhe6bu3OOY1LFwCVzuBOJTLTfufyZjRCNaJIftYZe
Z5m4wQLW+ePlzL4p4LGJQlLb5+2NShqQWm97/3hiRYangZR+8AGp96HPAdse7/4/85eMJPe0Dlhr
8hBKyUw3l6kncMbUxrwL5ISsuZ2GxreOlTvOK6YLHN5Rd9iesXjsHFPGn223Q/HHu3wo2juJ6SoZ
hyockEbegYdPOp5UxRHCUaam+LC2HpJTzlQUG86xzSr02XY2OVjIIVcN4DIhVuNv+VF6sU1SnULf
pX2PMSWbQ3/XSeGiLimx4m7WHm5xQH+H9v0LKYGWdatUXflMsK+x+S4cXmcYN4YOmg1/+cCPOPB/
Wxy598LNrwyIMqU7KEMakHL4GgsAf927oudMdDFYwQAwNlHEsB5U6HUlbd0f3JwG8+DWnKgpGato
a/+foNze/1yxuNkPKkUHo8luZ10LD2jUBbsep8+tLq+DjkaRGf3eXrEEd+BdGmIJZSSIPlahsVXX
8+xFLHTCw9nVXPfP0nkNiqmyN/nqN1ztqSNEEuLHcpStU2SV2D9pX5bS8e0kRzP7g0kyavyLGHBK
UAZL59h0Nx0x6zqdh+S00tepX88/AzxUiD6/Swp+q2bnl1FI2cx0rQjtNPMUQ1FHI6U8IEtfzeJi
R5YvgrMyLd9MSfEUFb2HwEWT3zLR4SZu+I6SfqTm+oIZ14ArHINHIMFVHrOTBnoS+zdPO8ZE9MGe
3oyEFXSO1uE3GWdAqQjad74N5KvXIDpuLn3IqhSNFBkd9i2b9UsoOtAQVDGPwUL6Zz1cPn3skz74
8/XYJXb2DiJMCOwlC6H951UrG4zOZf45PU4RQ7bS097vZb/4l86uO8M3Sh7MsJgGNQTvpl2NfQnU
+jDs+iKK8DcPIUmi43GL6aIBZt2nhgDh+B4TWkzs/Mv/BiB8J5MyccL0/nuwHMZBVd0dI/YCuKOx
KqYRBZm0uE2zM6kBem+hgxvEdxdYdN1G9TVKw0bIHAfjZF0i94AXQC+mfE7ODD6C0BAr4/ZrgEMl
bkyLVzSsOcdYd4SDc2xlTiEWynbImHeBYAGeshQqiQeAII+9h8iueLSb9/W9YWi98PklYNeiG773
7AyZ3/oN0/OirGgmq9xdd6wv8DGB2qFCjgXcryX7G6bsWv5omeDJW1jbOci7L6yziho5v6IrdG/T
5pLXLh7pFiUbH1RZn0KwNC1Qw4EwnD3bF3XSiRq8AUSa2/vIcGcnuxIr8iV09XBideEl8NouDb9P
kxZFujh4fz2UHH3BmQzvgSVG2tja1piz48lqtn4xrHhJI2icpKEqQPX9YkwbwGDTqOCdxrMe/kW2
syul2DZnjz1AItKr+Wpl1WLLzKlJxhaCwz08oQAjG1MsSX2UYySWMnj0sjDEHUI9yLJ71kipGxdG
BXppd7MdLiSUuY3Nv7Y+aQh0FkmNcoq0o3mXlpAkASnSCGUZWphvALhICiO3AHZ1rIhxRRbtLK7J
K/zXO39+DqtIk2sTQQKpKa2Oy2lDMd4LGZ8Vyx8JpLdBgShJ5grRbAQDrrOQT3cxSk7WAf+Z0AkN
7u+q+L3TM/2vNOCwOlltoAGIEDI6oUUZJu2zeDcKvbVsyNmrSk0QIsHn57b8tdT1GFpXUyUyH/J1
WFNj9M8uxd02LNqko5tVdJG0V1yyTrGoJ4WqaYhFpLMBF3qyY/rpbRAATKTidSfwN1vfUGyNuHXm
9DZ+a+g88ULqdam09+HsY1dNsCs1H6LZsnRpLFyklOG2nLyceXm01V0q15vOpTjKQ+2eKNbewD9Q
Xtcp1Yp02SdQMNsiivgm0Kdp+j0T+DwM6+bTmOLSaABJU0ooW4grCWBt4egDDrWK/gy/6h6tDDe4
LZYpGRpl8kwB1UYZGuYSsJ0p6wUOmDEhjpWkxa/6tNYOCNUd5RJcmolxfiDVAcJyWFQOkb0mSD6V
ri56ZmQgxjQei6iIIw/pO2CSC5+qu2obHV+YxF0loHRz2M3kKES5+UdUqi5/E4Q5jlZ9eS9FrAv/
c1tc7bbhsCc+M8aATwpXpHSsoVlcV9GIFWG9x2WtUArFAMkngnX8taIssQmc9lDMTdgyUHu5dld+
47GS/xi5XU21voI54LUgHCkYvj1qJBbu5lc81tADjLTDHPDby+9NGTiIGN5Lnnf73Wusis7Sjmh8
quGUQOi7jj61NhSTfOpwBKCxPI3VkqfE+ziMFcAVz8mDvMZOg1iudwigvF2YNNlzXSP624tNOOZ7
vB0zpGBn+2rUKKCuJpX/NzGMnzPzddd12brFMqmXGlY/IkkVOq2fgQatTGMjOLehpWzJVfvjhT14
eQiYzPg9BBO/HCcxnfwgIawaaQiq3AEUQgvpPkMKAG0sTqEstFJasxpSSo1j9BAkMglqREoEJjOI
6YIt9xYCxfF/fo7SXQhttwAKJmiPSX+4Y3oaPTLtzttbkO3PGzNITE78x22/E9Hwi1EAx2tqvxJv
pLJnVTBc8oZCVHIQUdO5QfWx+B2qam/FSw22G7CODCejtRdigvYmJHk9cm71rCTJDzPGuOHH19CA
UnNLg7A1A38YRM28cseIRODa4QoDfwaNzD7AUgjaAQbNWmYsueyO+HbKjwEpf/eBh3NRg85BSHQr
mqr+AaZi1Stxl4Vk03k8W64jX6mRbZx3rFJqOho+wMDfALD2MNESbmGCFaXGR+DVdMjZL9aSawRa
SsCKHi2CE/QNISdAPka1PzSFK98NVw9uIjT5VEZGtSph0XIYEySVqRb2ut5AAiwyBEDuLyiYDZ2k
iA8BoTa2HWdo2kJ8PBfGb5r3sg5AQUPhT5rD50ZqpLOFwCa/Iz+IzfZCOsjBnfU2IkmAfBSGY2TC
sRTIYnv+ajfBZlOI1c+A8iPv+lD4px46oYZru2TcYT0jueIUyStPQMWScEkcNDw0+0e8pv7uIG4Q
FhZXO7Vvuo9avcklXl6SyihXB4/ktcOXutGfGKqK+3xU1KRnvyiiZjPmXHHNMx6dmzOz7mP9IAzM
CsVc45Pjd9N6QOFu59UBqCWtaqvyZPWOzUzYHZcxDmrX0WhFMuvTvlKJ9nt1bV2LTsPcyOx7tmne
e6QbcDuXUNDf2PtockM+RX+sWMMPDjcB66ECssUgDGKjATxUddO4mXErbkvuOR/ZJ6PA6FAqOuQ1
qfvAX0exaLpcpHqHFs+3zjzmFShIoWTQvMcHNriVD2+w4vscmz1rmQ8ezMuGKKflJ6qRwQAwrdgx
cFPIm2w11y1fx8LNfjY1LCJ4s4RDtuADPrF1BDaG3+/umAvB+70g7jclR+WPUJpPdrwytcOqKfyH
ywX+pBTRyJgJDxa3FYrzhgzYIHB/eLjUOmmzNtgCOkzlajQ7owrekTeCI4zhRf2uC7zwXcnkiXSZ
qrdAcvv4uu9uN0QHyneaEhEVSWbg5650Xo56ZgnphF0CiBK/9Dgbyc5BNFADzE6/4vIkxa4WRcQ2
mPcFTMND72liMJIjISl3GBaKwlUrjZPIy4meWrvJYwTK/YQ1c/m3V8rEow7gwz0naZwgFH0DR9TP
fAnAyyvc6kL8Qczd+hTBmFAo97l4X6fcHqj4MgqE+64nTu3IV78ITtb7aE49yp6USRCwoUB7NSMU
IHopCbaAJEh3aQPRRDeVattsNDKfyxMT9Y2N2A2Ump5EhmHIONUkBcEkY38X4woX+3uyKDCG3zqn
n+DxVP8uTZ+8kcgwVEzmG9LGMCCjpSgiLE9kWqdUXwUKX3kkM4RicIfxa84BQs6S4X5UqtEcjwaN
zUmP8MQlgJ03mhsPlUeybw9ZaEQQy97v4HuJ8FUBLwPJsJOtOGz0L2zoTGJu1JUl6mm9aNjjF0Qu
gAYvPyemCUbeWNs27SC26ONt2uAZcRcj0ZgZs4LwMgDo2DYmZJbB8lJ4+grv+i7kfhx24H7eqN+d
6tffocSrIGIRVgE/22Wh/54c97gSoRjKSU3pYG94QYXT8JHS3GAFDAdGLLqGfEljvCSq4W/I0lUk
5bn0TgnEv+SSiHcWpI2IAXszQ77Odro0upSNRrCpOCxXokccPIP4aUmo5Fqhxnoxsp89ypNQ4MC7
YeftbCnKCgPPxRef8tqebw28Ab8N+cjeY8pLYYL/2fh2yFDmTVbvk2wvt4S7DPvVhwUFhmPTKDr3
9KqoTUz6gP3k/wavebmPX3dR3mBOQpA5A6a1O/mbv4YUs/gRlNWw6yqPPOZ9ePnEkc4l0I7ov1JY
amJAJ26kQLLmHGy6lSCbb4CwHRBYz50tUzJx8dCuvfvm17hNqwPWhi9zEoyOl4pkmU7nF4TiNf3r
vXjB40EAbXOoXHjODfsNbKnZAyemYqxPNSCBALOmyBL1QbajCNj2AubhnnZ5KYiAWxI+ohjO5ARb
FykrgwQL2IsxKZfof7zxDpEPtLnIqor9CcwlmRxj5iuIPCfKaS2igHO9fHtOgVSLpwaITw2KMnnA
QjesfqG7NAt8SnF/OCmz7RyGghCb7EIfwSwcEJt6iZV38H2h1g8WFUTTmuQgpcTX6ny1eFWJ2gY6
TAwC8sP47ILnJKt68VQ6TZIfH3K+HHamIjfJ5sX/WjVXSnXAHukuEJwgQlb9Q5BU9+y1oDatDnmG
imfSlqaWIG523TfJiI0CaX1rW07DUArt70HEtW9RO5di3fgtp506JdjCu+52X/ErgkidHDZRNaTu
BMQSKCvO3+fJpsiNahKvdFIp0cu7OXnzwo4YFFwpgYtQ5YLqKeUSyTlLJjuQknEFzz2NCGpvO7sG
gZ+E5VRXUeezdZ89nlw438stba6q3IJVCEsApcM3eRud93y/4OSEHpZuu4+YwoAvVIrm8JAqTuwL
vwW0efruPikLHuxdUafhKsCO7gBHwjSm0jMK6r8IQs5XFgC1ljHaTzr5tUGRSmG8iFgdd92RhNUk
Mn5fsF/vRhfPp/PHKfuT6c+kOkKQykP+IGbltOlqClNRRoQlOcsEr3hjmWQQGfyAIJNDKokiIC9L
NWNKh1uGb7gvbFU8bMWBAAZ/J91dNbOPatVmIlWGnF+b5bPx1O3UacbfXUqtL0VBS3hr3Ogl2lya
dZSdmBfitKyyHYlcMMWxo0Y6HC08eax2lompnoJ9lTJaOc1N7aDqQHQ5wscmQ4HkAfc59PhQZnJW
CeMkvTsVQJj3Ciy7FAHBsaIVNljH611PCXTX97ZH1tSZOeG/+cWXQumL3SoIdMoLVcLG2R1G8iD+
6wC6LaYFTM/A2V4f+W+h0CHWbBVWpZD0UNZd8wuD2AbmX7ahX1FWrHUAtRGitTyAXZWV07VsurT6
UT1izjMJr6rTXNS08u0T2a2m+IsZQ+by4Y0736lhM72M5ABjfOSk2jAcUc+dI5R/rq4/ZPXjr3JM
0B/NUKAoWdlVMa14TmSTcWh0D5oNVzXTAXISPMCL3Gth91dolPp3WQa4pBNQAC5Lwv5Di1WTRu6a
TFOE5R/QelrpHmdQsKexocXx9v+JzvIDwbhwd31UHHsgqxx8jb1S/0ZN0TTjDsBUfglTipOHWjep
qwQL+N+U+9GHK2G89z/gHH09Q6Q38OImKg0+vgCkn8DXe9QgYyHceKOVyjU07YBMVcRiUdBLuLoX
WJfvPYnqL3tNtC17yUIHMTKOpX51mvXkTqO1I2Hi3jpgh8qnQ5+uLOhsu/SUqqGlGZk5JdRwVgW2
NmZZPn3BGyW/J1ilLTJNDf4fCTPVEdePCxug73/wTZmnq1UmXihHb2eh3RLEsOkF27yohkkvgx7o
GYyUCuoR+R/NWvgva6nbk+DdJyCuDVu1Yelybthsz4rOvB8Vnkq2uVo2t55ucyvyfnQc0lKlZmf8
iid9q47gbO4B+KgF9MHjnxP/pYr3JxcUwC+L7TIlcWITy2klCRxw+DE0pSFEcIYZuVW5PzuXmpyx
QrJ3Ppe4R79UTHhHAdCuPzq1kZks3sAIxDKOM8j+JJneykWSYuYLN4pgQLJboACZpESfNloR7JAx
rwsQ5kb+u59ICVZfMjfS/Skdj4rMBEpM0muXqOog+vllRXXzHOa94kuFRf0xQy6IldPTWKEX7vxg
fLNLdO4l9+zN9QlVkg/BuBBy8dTuaWxHGR2NIvf4rOO8etKT3Z20ztOLv5qm9ZztQ+roo75U+FoO
XKv/Y3i5RcWXzkibadiwxSl7lZHlGsQHrOIIANHjwbX4P3YEZ3XEfN8aFOTofqR+AJwm7yHb7zU7
sAtIou4Mteb45KU+Svl6O6nLFRNmRbmxWTArRql3gAdcKMSz6PipMUqjZlW38Y0QbxxRKUZb2bDX
Vg4u2x7W3lao0+dHmrPa3QYg8uybnRAesWtrErbzHd1P2rVYeMIgig7scWGc0LcXbHrlWc/uILWL
U/uw0T4oNUyeAMrqiRs8WGTi7nIQ8b9wdJ9SjTUemlSkk8RuwwfRm2Rc/deqEDFMXRdWE39Q+47P
swU4OECH3QRG3ORoyHXYrveV40JSCarY8VQQZ9//nZvtfzBtqIgRhFc3/tUJcp4QeRsPag1+hR7F
TIrJI0aDPrnKLwlj54bxo7MLfLxfpCjKQcBRp+xP9KTBGf4J4cbRCwFKm0jx8MKgClZqhnr5Djzz
ZTWfhQBa/Bb8zQzplKPMlDpRMOxF+Ly9ORMQc7U0888a2VaOn3QnNZtpyPeqCKrAvjn7oYpJkQyO
smhXoNI7qcisEMeHenLyE8L9KPksvF+UB9kqnUJoj7CHCswFunhC1ACkJOOFEOZx6SIsY8jEF1D2
cBZAbjBpPbogYgMmfpcMxm6v19Kk4R3mUCsIuvrZOMNZAoCozUqRtQnGYJ+me3dI/y0GyCjIdF1d
JHEzIUUa/TulokJrL31qB+xpNbqnjeXP063Y/bZ1Almk0q3rgV3YLXWWKLgTOnSfE2C+3cswu+/F
UIeEcn9POiiT9XAnN7WQIIgfXu/BQbmWOf14xrturOznzEmZ1c1ConxrsPYFRp02FfoOgh8/RQk7
48yO4+32q0VF/Fb53hon5xF/O5bd8Xb3ZzM76NhVxGP17ff1sYoIxc3lNJH67AmnSNMb7u34JCVN
KOqt4uj5T+mJY74CwfdTWw8TTW05T5vG81z6Zp31tzyGVISNSYFR1Sn4c059k2D/qlkIbp/BQHyz
qlkGdTqcjtPFcdH79He3pnzPmqUavODvfInWHttlajCa4bqBfDcYBFv+LSsQaCXCJ84tcXlTiWgE
JCmWbtDBmBK7QWqEfD6vyoV3uWWKIitFV7c9O9WQrASkOvGr3cQBuZv1IDudVqFgqRFWxP9gAVNf
wlpFC+NjMPNI5deMseryuFeCJibeHZrtS5tIQSGK28fjeKqloINp5BY2IQybEDcYT196AQtjyHDb
skik4Iu6EjTd23gkgM8NajFT+S7UX1OM0WFbRZvnPkpPdFdy0vZozzxC1OLFD0GZB8TnsrZgHOPz
e8JQC8SsJDEbPX5etXhv4Y6Zly0zr4nKBMk7lI92moiZT126kg51K1fr08RcoEXVGUtA9w5+5PS+
YPFVmzMWrokrzbwTqVIqTlIMmmjckkMdR8OjZ0ladeO4wakKGKh6SLH51R2CCvVLWLyB3XCyIZSX
BSXcqdKyeiDTQVQgtc78c8Krd/k2iclV6osbNnZGNapb4iT98MAWE1i01p1u3gmEcvCWYxi7ifNO
RwEJY33I55M4JKhjGmDun17oPhuzlSWP9KxHnLKGksw2sTt4IiEFSVMFZjqbJM+KDtPAHfWhZynq
+taEwr/n/yVSFswR8VtFpdKcJqj1vkG1IlYt9R1IB3lXtrOHnKNqx7/RzSiUcPKdXG+wi2dx0tOB
2/c5rEaSQ04cqUatOWucbLaOiFqI0kfkdEWdEbNi/XmyUtpHuAMaQ5so8XC1vKOcu5AFjOdcZrh1
UsR5XFPc5xh4wuFD+2hOxD/bIi6h4oDnvfbBqCv3Pyr1yQKXBVj/hcT8aER1U5/5ofeqOFDXNkov
P8yGNjbiWy/dFz2gtSbGEYNk6bUHMiaRuxl6r4PKGTVl0EDaG2sTnzWK8iDkSndBSTBvmB6m1+ZL
lFOV14WQIuyJ/LPsffxrLW68t8NhEDYWas7wcDDxmHUDX3hQKTwtpersBPg2QLVCTq96M40K08Zl
jcaowXsx6MfFnsY8FdBSyM8CBiqgqzGKik9B2fh22wJLvIWOmrEj9YsHlsVTCyRr5fKZbFVVCC58
LCRmSItnvcOWwTJGhZkEftqMDsuDNqFjIyy0a0OBdbn2+pjD7jhDd7TQhHUghHnrn0OwV51RrKE3
gYAey4K9RWbfJGbu1pbw4yAbbRRX5BvThtNs+Ww366TPXKfbCRx0ZWdzOtBP90Z0op28kwve0FXS
6QG8dw4LKjz277RDx2RtKbMShZx+IngUZoNkx0JfKxzKhPh9gxloS49a0EPDMMsjl4odWQ1E0v5b
DInQF5V83TbwsmcxyEeV+4psc73VGf6zncgoBC/cFELC7kZkpfhYvK5RnldVBcB/CqVK3vbK18G1
ZeOcHiJwlXvf25FUTFiIIMaW3ICBSm1yge2Mp/8J7CX8DCs7jzCNWDiP8dz0SJpAnYqEByzjw8NJ
A1NkBDMd7q+FEuJhV/GvRG9q6TAGORvAevf29F2V3JtobLu8ltXmF27ks5erZOp93uU/sZQaJ5uu
Uk8ox57ymkNm+29P5zaBnxQ/8ukGZmi5tB00bS/fPSOU8WT4sZFnrJZvfAfofEYSZvQfKDtvtlg7
tqLdq8d35gizYwmj32PCawfNOa0CP8SmZN/qDzsdS3bA1rDuO3At/rYQ8PP7SEMTijkVL5BHxTgp
3un7uIZW+1B2rFhyJjBkTY3M0lXMhOE3U7adWk1mUKiAu8ZkY5qAAhANP1/IteqMm8qAAzXFvpdm
KuTfw+aVpRDK1pI3Xq+IOJ4MikEWZw1SLtfy3ZzzQP0Qlx5XytPdRsQ6j3ZbIOBo4iI+OOvS+MIX
TV4crMrpY3lCbElexyG24Hv3CRW9d2lTlsSSXmTafY9R/Oj3NuNg2UNr0U5XEtIbsQoC3P5rz4ac
cwMF3ty2dpxLa6FbS+1KCprfDB9G+B5V3anxSdBI+RlVKSXG7uGHD8I/FGkxmdnu8hxHtFfnZxBJ
BSiRNmJQjFPw/vL/Vfqxa5FmeBryZhzlQXPnHjr6irDlcYCFBeNxRC9CAllX3m8TPvsxSyoPxbtH
HWwqLg5buF8V8qrp5fdXWV7vOmrCqsM60awwZNfuUzO6GcRksCc+wjEndJtCn6abRshxyQnDQhM7
wGyZXcbbmeOzHLfGdSawPVwJdBXIHFPFuik19r5etfGRhJ0ia104+MwpfOX9WRZ+MXY8+V2tuF59
tWYbbxXtQfpPwXW2bw8VpdUaDTtnKJXj6Uh0dOd1KgCyCHR67WYqjt0E41/F2rNn21Ss8FGawTW7
+Gvj/K9br9qrVYsn91krzGe9xjvp9l7Pya4wSPb7R8ty+kkF0UAyAEiKrC3ByM/nwIiwGwf8ak00
TSmSu8TaCGqA4N6zRMmHM9ymBGWZouooG6ge4EO3BWNnxFJbx/Wdc28pnkaGsGFJRZXgNStxt7qa
UtHOkuqOSRG//J97gbwJzr5eFCqN3m3muwbSKZXQsAZisOR6EcjcTPixD9NDFv4t4tq7ElDxzWhN
sGiOZJRnRb8jwthXGwma0Zt6qCbJ5aws6MZtMRbBwPwjnWQkxWklGv7z/bv/J3DueHiH+GERql2A
X1wUB3By8jbCsgpwb4e1wdYtzvW3O3WgJLPssGzeTtjVzYlPaVZ5JjE8gKrG3xlub0zVzK3ZBu4E
vzMHAzSxrH8JMyfHs24IbW3b2rta6ClHxwKpOqEpl7FnDeRg4PwXFqkQp7+wK0OEhZ0gKe5GK35y
iol6H/Xiiw9QYVXnX5OO36b0zAeOqk4MfW2FLEx4537F1E+PzZii/u4FZHa3ELreY9u8vH5EhIX8
xNc7Xjg9ohAoalTK4Nx3golkkZwWZpetEqtPWs+c8DCh7Dh62PoSuZgsUor3cxWsXGEGOd95voLk
4WeSf95QVSWtJLiWRuT9DNrrYel1SonqCSpavZC+moI1QLthK5HS0dP1zlCsr/I5shMdTF9zUL8T
6Q5+k9jUKH+adM2zM/v5VxNIDtI1QYzlSTa8Xk67H7LqQEqu2uuDvfKegvInLTbsT4rsYxFTijev
7WdK9BuLEPjbAKhtcZqR+EZvC3QBwO1uaOIN/ofjgZ3Dwyohtl9i5tM4yrt68iJiZVhtWDh/pnvI
xUU36uWR949ti9JvXI+yO6eFAcrULM9zL42aCQ4Lk8CfsvvKFhDeNbnsN3X+l+KG92ip4PJ48IwJ
cCYY0uyzAca7TkpG3WugcLcFhSRIbGRBLB4jyxdiZxLvRFaWsMvYDCCcVii9NKcOQefUD6835m5C
+m8RwxlrMNg7IH6PbEB0ZevHMTxZoPTwo8NrrbxncMLBwmVSfYWTTYJ6uzL795rG/IayMD9jqKzw
mk0PyKh93uDaqDW6Wb3ojp2p8HbrEKRn7voPvfXa3T6Maj1vlnY1BCJfeMTyO6K8ufdgjKKLO6la
H3Xm2f0BM0zJo1pbe5AZiH2SIj1eTxF1GHmZ7loj1KRW98R/6FPnbLwQlepQ/gXtRiXcb8fL0i+h
tR3+TSibHyRwfyF9jtOrb2FE4JYU+Kx+V9LLKxoPKviuL60xpkUdO+HTz6tU7qMtDb9WXPqm7Tcj
Aj+XC2N5AU/Mlmlt73M53DVWthKlXW6HJcrhlT7K/Q94UlMahzn4lHL9R1wX9vKCk98WICj1RHY4
1t2IWJxfjLbnNToY7ehwB5uuZcNHrnCHNTh60hWhry44pw3swV+zXl91+QnzptNWPVqbov94Aju1
cNeCc+AmlyFWHwpmRRnbwQJO7U1ZWoMS3AXwGiQJegMmpMXVfWtbH2wtcMa+U36HTy/Ee30hofuB
wUjPOlFNh7kq69CYo8XPRkKeBF0RzJy3Yrov3j7jIperaHD4fleKr4Ryzq3qjOPXCWKHYiAf/sJW
+bWq3GRiesLYoqXESZeQ6+YQOJZtAqBnffq+QONe59E4x1iRrdAhCqRd66q4Soo441eSt2ide/8K
oZWkRGBB0B7UhyQEznE/bYqCbvlvv1sDPk5nMHTA+IAMzKW4O29ACtJi2bqK3WCUoUK0L4JEfByO
VeuUbSPCnQ9a/RNpZc/BkRe+ciPyweT/8SSl/XjO0p9m3abSPkKTiewfNP7yKyPyPN50brzAQ7Sk
sUZWS2FgwBtYG0viqvcDWOFuvgbX085Xb0rmv5D1ecvKUwB5ABjPdHfQ1Nrfgh3yNZi5dOhXzjdk
ahrJCbpoUy1it0MOYRP5ELoYg4GRfocE39RaZ6q7D/0s7Dy3mcP9WHSOyeHkWQiHK+bxLAn7TI8B
oCeoYFRzFjdhcGhEm8XrYC4FUcmgOs/xRmxMoxWQQkQ4VopAlk2eT7VIyTKQwVCs6ZZ0RhP/qQOX
PK2gi7N1TTHyLMQpQNdV5n8+nM55ujYHut3aW1gzSnShVt98CkKjcvPRkNnaunMIdGCrb0mxJbYl
J9SUKjTHLd311M8wdFUejAXPSC5BVZpFA5EiIpKwoMcHLsa0faTr6s9v+dE1UisyvhuioKMpZPPX
TWsiuKkajEz4i7yIXvOztouczrZTkOzOycdllb4+yvz70yE5/9LX+kc0NLV3TE+1xyu10XFbWUbw
9tDzMOySJXEtI5CRb9MWarpjrmq6CzcuYu32as6isQw9H0UIHlWCUQJuX0F2BwmsiNoC3xBqdC7A
Vbm8fwWWRJQI82JHmXsUDPmq745eqfcnC1fgI48qKajFM/Kwu6luXj26ykxOBGEvII5+tWv4X+Ew
c0X4oAh5Cmk70tMNZpO+jcZN5WYdgQaxAETBmb306kSzuzuFNp39FYc+jG+sHiI30ZPL2LDbn+dN
bn/pVSgkdYtw7wHZgvy1QXa0MiO9F9oqIe6Dg/E+eCT8ZlNkNCUAPkcDa9bD5+NUddmg4gI+o0Qv
zrPGC6PPW1kN9y+rO6WOO9w94XWQI/ZPFKVfVl6f9AEbXvxwjjBQYoQJj4UWnAWs30YAWata9wH+
ofbwsTqvCn9aq9iHMhVZ/6vvbHMlOkRVGiJtCO2HCPRMaUFBZkL+gYXn2NkAcN5Mw2xmE9rqoqr9
fuTIZWjVaLrQkopSjHtgOJ1Vnx+6GBqRMxBuu15wLga3z0GmR6b2y2mO+OzPAWJyY7BSWoGlJF+f
3f2+wMeS9mFIbRh2mA2WWlhsLwyudc6JH1Ey9+r+Fxe9AlDcajkZ9ujv7CsysbnTIXlDi13bRqWr
PHqm8071oeLu4XgznMsmiPLLPP4Z1s4bebB3aJrbemjsf+iiXNGL2F0U3kcpUgljzYOcdGqgp76F
202X3gP5Yy7dvf0N5lYvISHiNsvcjx+XgRVBzA82hcrBqYce2I4s49WdhfJQF5CWxJmgCymxTt20
fRkRjManxli86avnE931SJKzsVr45/9Vk6pPT47GRjuxMqiSeTl4m6mm54NLecsLJSNPUjKw9DID
7CtiGE64OxEWSsZIOmr8zGl60+RnUYYiWjAnfkJONoJWTeoBwFSs42D/6c4jBnqCfddehWJabnep
btfC4pl9/sVxEGAPmE4aaMzJ5iPNN3QQKXPzmXzq/o2FpjSiVOjBnmPKbQA25jIcs7td6R/x07vF
yk8HdOjMWBlrGKFqLX2Bq3VEmp0Vmb0hu/EJ2iQVsekD2ejVUINe6EnHR9jyNiqLVku1x2CG+pNg
UBX8XzaflP7NxWmgkAoYCPxDjPYmraj7NdEjHHDw2HavmWem+1dAiMn0sJ8/yy0IIGhGJ/bLp+x5
N7HeLWdBTaB/DvKiE5wcAqdnFU1Q7mgzMTQ3hgc3C7wDLFq6nO9FZ40+G7mFovGlm1Lv0fInDlSA
af13i7a8htY0wcEQUB9LqmY5GOsDwX9G3a8CbPyJ/nF0jMpYdV5g6jKqKWoEAQroOfxRLXbpI4dk
g3HZPDoMP6m3WG3ubYFn7L/dRfx7JjajW5MTvDB56YaZfZUW7vp2HL+YC9pjuoDLZtWCYUxlwHWK
cv9pRjjz+VQC4Jr/e7v7WzZavGVa6ICq/kb6OCqWLafPN0N1wxzelH87z14swWGGNYnkU/9R4PUV
LB3W1hcUxLPrOeRF0AoEwKZ3gCZ7V6aikTarcWhOuxZN9mqC2aIZK4OXFYpsviBcnk+SEKh1jx8o
Snx8lzphxtV5alACaaHngewKRXMVQiKpxcuO4rRyX6OQxF7IBuiG5AQA44vhfGDuf7djxTAfWuEA
e+cXtetASHAWQxKdwPrDt6CiwgoRVqBFVQTQmd/mIWmDR06eobocQg66aIVxptMr988WhQHtywDF
sF0xl5A06mGbz19Okv4XDQrWzsReTYXA09NNiUnvAQL5EaodOnu1+6A+nUU+qWgnzg5CU6YGyxj9
yjpcmrvoUPHQeeRR4VID2CCM8hHbj/473ZJl2GDHI0tulFYidagNNck5mLrlBYjL1mq46w6/7lEh
QAtg/3HQb3ma9X8iV/Wn8cP1y0xUwu5V3YKz1CpmvDxvflp8vT+Tmg7dNHm/knOSyOc5k5j7r5M2
9nHKtsnh04sguOquJ9hVJad4MPaSFmWmUGsgdnOYp9Pzrvm+8LT70oS8OLnZ9TCE0Q1WenbU9BoW
JhPro5IWFlGU5hP+p1ioeM9ZRe3vWR3YcJiDtcb3/TY42CZYZsyKxeKxLpNPR/wzYWHgaNfQUBpY
APC+8VyDcccmprROEoO9jorPkzS0LDCTsrPsE2tZuqXmW62R+EtpkXZyKhwenGKDtbjDfQ29dvhu
vF8MRKD6Zn5ynQUDt7guxrG60LLrTNB88RclTwy/vEJ8UDbNlwfwD4v43mi83VWp4QsgHEUlj3KX
PNYJwrtbzkkQVcrr/XfCukyh3BbxZXiaSQwiBsN5zoWz8uFj9sLlCzkqmOnbMe8CkvfxJhuuEua1
YyVmGuMfxmRW5S4kn2m4PvFsdlkhpeCjUgV1VWsSs1jnuFbz8HNAUBeLJfRzLymoHiI4DjWzc5J1
q4YvytjXBN3BGbkfwKWghyaGxbqR+AYSw/fYBalfmMbMvKzqzdjXRDSK7Yw8w1WJA6xRS8/wqMA8
9Cm7yXN5o77qcWHiC6P0IiS/ty2aBCE4bsCdb4UlJ/AEQO3FWJp0lIoBhC0Qe1Q6pj+pxs7cnX9W
zBZHDiqknmVUsf6oQXR3YppASe0182B0Vid1LMxEzLZcxeEV/0bvZoZwQoC0R8T3fFDckAQNLO4O
t9lgIEkuq4DOz1s8w6djx5NXGJOPMnC3y0LQkIrf8rgwkRoTVNwq8N/wUJrR/Uds4iKQGWOwGRce
JKBTLdbHs4Qa5fm7dZLMyusJar4sMlOq8fC2jFmbMPPkKM/fLhtPRObICviRUvdZtHSdycb2XRDw
TKr5rqqIVEiUPlSxRROVZaAvT7uEQfRkoiCvdSKykhCt7htYnI0qZ8SMmYBnCdOqaC+YRnqLCvdl
OPog39W8C2epZLIM/GEvwBz7b3fCZsd7sOzBNbl5vcvBf/Fjf+b4CHQqxdQRt6CVLOStgv8lhVsF
OAWbkvDRIKMcQEIYjhfU5tozk+zGdSmEpXglNr6Wvzke0ezfKoVOictoChsA1XalLf5XusnDSr6+
XppiVg4hAQs4ajkpynIbWybk2Dg/QoTGDuOSlpgOfyvQxdBPsNps90gU+dbtd7hRa8OiWmQNU9AZ
z3D/4abG8F87GFtZ6l3spQIYPB2sukPi2W8kl0UY6GH/PftHSlHBmBobgdZv5FHYcIAffc6auh2p
OscCza7BVx1AUEtWuwY8ZKZ5fVPqjh7GXcZ+Ae2msOI6wzQcXUxd3mYAdqfj38tbGRWj6JOB/2Kc
f1F/WiY1duY8XqS6BVIgF+Ia2M9A70SzeDzixNR910OqqDxsQ5BZIuqbwIswf9QKnMxPe7rEBKU0
CQpgXBmcGN72tw74jq3LLN5RSMcPSXxh3EvpPUcPRfGZJypSwVwTAO8mIYFaZQGy9+r7RhCiHN3A
ZQlZ3csKIAkJP0ipILkj/YoeV3tDRZlTSi0iDEQxpeWHWF+T+FuxQSIgJfC0ROhBZC3bGq3q7Exq
X6DSskVFV94WQIXnocsrgQbAeIzDYcgbWdFBx2XmtmfTcLTeSrNMCKZQPCtiDCISu9KcXrkqhr8O
Tx0N+z+zzn+45bBJewei8UZgStd4ENOB2btjYE7BI63HMFC1vwNiiF0fKToPs61Ge43CUJjGEl/W
RzC1ZVT8Ex5Le6hI6kzQ0qAouT4UaMdJbWNCdIt9h7DqsGEQvoBCRJGauGc4hMdWte7gm2NhQ+qM
Cz1kxnWp0RExXNxP95hCB5UU5gPKC601OKdUXu9cfekwsA5LdzAwWtJa/XkKrjNo5IVv8axWJ0II
z5O7t7x0paM8I22eE0rlEhklzzx17hr/0Z7Fx5WsALRKVtkKuRMkv0jzGLHjLQBorpCbrcI2zipL
dc8C++XLcwtJfPyIh0AW1Y9nyC50YlJpoVtxD/8UG0W3rrfNFcUygSwPlBFk6ykthUcltmBR/mzr
2KkdavCISON2npuzzO3cO59K7PsYFVRoszxupaBQOOOH1++ivxGxJuJLN8nAk3+p9k/6sApdQTbG
LJq8ERoQ/EeUnAS/Mqz+Gr828ReyIcLCnKV6RXA1HfYQ4djyCH4o5eJI99fyuvHf7MmYddI2SMAm
HBuACc2kKiE3cnvnw03ea8QRDYkz6MobP/w0/iYhTQddIbzV00DcYBVBN4lOtVIOvtM1v+SKZ8NT
mdq8zEc+5EjFg0J/M2n9xGDX7At9fTKhMznLYXLhKLTY83rgoa5DqgkW0tQOwMyYgKPCSxHwGWko
5r6MDbUhLe0nGqVy4z32W8EsssIAZv3bgiR/ko3T3Nag+YD2fm3Rqz5+/iCCMsgeDwE5VUzvrsXj
JZlYkmNtDGzbiGtjl5NKntJXbDuXo8ziIQBUw6NEX+P5MLhqHOdUcY25LVf7LLHrDa7bG7Y1uV0X
7vhd7cPGAZUXgI9A2qZks0XgPVLAOLa/Lccd7hF1EHk/kJ3iIdybaq17jf+JSxm40a8B5wifSVkl
aPJVZ9p55pt5bZUs7GdVY9+xLj32uVDz3WgZvntq71UAyDx/2wqDxsOOTim+lvD68bHoNEh6YiQ+
GxJJyUsazdmezJvvwuwHKAaJdmCti0VRRL3MMTO7/VzrvYvo3+E8Q/J71ftMS11bN4JZ198VCi1z
qsD+o5b3SSoK1qHpWfS3iQt/v4mM5+NiG5ahoaYg1W0EtxBRM44gqkmrBg7nh1RGEqcuSy+AJG7q
PkxDEmQXzSGQdtLtk97cFncEiQfYtdfGAuTkWyVRWrusqKhZkVRCfiH0OQJ2WbAWldcbkM1kG1+L
K/I84IE33LIssNjWWd0TTievtAebR7vOuQNnsB8ATIe8r2YZaE8LB0fxeYaFwyZusXE5kCNmgr/V
GD7K8QxcTZyL7z8qBHsHadGtlRZOUdJ/AypC/vcAgFgPXmSI2xbHI95v28cUhk7aW3pR9VBQCCin
TyxLb+2tf8vuAidLNuRTTHq/+P9vYlhSWKxo4dQvE9Fpb4A/kujvmo5Umq6lvZDlu48aMFFkW+M3
ieHqJW/S9ZLR/qcLEsczfyYMniio8Q8qSbt9hwXi3+Zg/D1qBiQ7RWSyZEb0ztXuyLOUOSspz/My
NP57lVxl55/OqZrofXXkalZkFiBgi1Pnzz10uLzTpGFxLWDIRd2uaGe6+h8+IzbBB8NzEP8MaA23
dGBN1YEjP9NHF23AKxy2xGnCDJBJ1Rk03G3s7+uj+w9kdK/H1ekY55B8kwzvWz8adbRGMBStjNxF
SdZG2GSeSjODeZVGw3BvSugL0AWI8acwyIC9x9PqFairi2Z2eMKkLqcXX2RusPAYX7ylU7Y6MvLq
HIUaXqtLqo+Kv5YBThxj5ewjs7tPDDgn6EeEbJGZ9FKcllyE6xQWxh/ZRje+3ipGN5meGmsneI/V
dRiySZtKwMiG9SMTvdOsGASDf03OdYu6+qqIXqzpQTuUcolcz978ujQFVnZy1wXrg3d4guZgCMQN
SI68YwEUWhWal1XjD7iClRuWAMrfsVm+AmV90tA355iHUDlt2HFHrJap836hHiqWjQYbskhz1Tn1
jFDbBMuP41jBROEfCEcwIwDMLILocqieI7MWhhbQFm16GTmG/6wfGEQYzvnLbk6hCHkOE5/3qLwz
F5A2fOh4iAIPLwdqZ5PF6UHp30YIB660jj3xzxg9CFuMrlo02GRrbZ+UG32TwfNqFZearFBQYXPh
6XkwV6eEgx34yJvefo+AJLnHMY/SO1E2bmtWrcMXm8D9/p8XZt4QHlym14FwqCvggle50QC11dcx
xHgia6WUnq5VyOt1/gQd74YzfF20Kbc1H5bJCOySRVyQ3Vj4upfs5lC9L29Ro5azbXCvg9oodSRf
wHB8JnuqJDgljglkmsmwDFNsqyC0ePqw2QgyWz4PrFg+hq/o8OkudMXZ+f8miUXcVbFmHwoQ/wko
UEX/8ABLjdLXXiB1NnW6iCqWs0jy1MZnHFZ0UhWYdxtNayqAdJE5EY2hY9T6i3xPixrGm4B3Z8eE
Qq7hAVhi5+sp2ihBpRro6WVfv3oPr9KM/WSllDJiJxn11gfSFV22hcE9Wf5Utvxq31ZLypFGLMzK
zh3Ret7BcdBXfXDmitmETyxh4ELM0kxLG0YPZmxb9dZCBA8bNWQ2XmXWEZKkuBkQ6yrwk5+pFEZV
S5shjG5ix1kW/k1GzMsWqA7lglT/0wPOv5qLuZmJe78gRzEHvfttYeOQ5gRFYKqH4QJbGmkn2Vwq
BBWpQSECFnc4XjS4IM2jjUpwQXY94gyFjlnvtzfLqo5437+WlRqJKo++kGxi9U5RJOPJm6nRi4bv
xobsmHjHX19Hq31uDAhg9g9KprrZn8+aG1s+f/WHbhQWPIAcmW0gQvRw1mpwNP6s4J3neXytwFCm
Kz4izUP8m3fQYXsH4bKCyhdVQdNncStHDmUC6QNtoCyQKWc6J0p2kf8vHokVuVjXy/0yi1y21q7P
SWnsYpUiFE3i9zwGrEHnYjAR/Z7IxNkbAHskX++mHp3lJX4Hmw0Oy/cS+UA7WYCfxor2sYpTWB7y
ttQdI3tPmvQ1OeZbvsLoS9fz2CLmTfYKxuVz/02CecO3HSp3ovVYiryA/BrG7SkeDBsb+2LikTNb
bAlAGSs8Qk1KeH+9lbFf3+UzIAK+sa8H00Q5puyACfYVXZ9j0RaTO4GRbr2cxt4NIBFrulOobxdY
ffR5ZXPejHIaRyTl3RqRM0MJvb27hc8PkAT8N9lzBesHQtCJLTfDg+CZosTJkm2DVsRp87H3Jh+e
So/UpSlcEgZDpDREYz/ukyIATAwqDkBOL/XOVAdAJ/YWtr+ZtOd7bFdP7bXS9vXlr7IXRIj+UYRs
wyySzql+d0npUA85n3EyYJOBMPr1OPsokIh3JhwQ4VrGtu6qrqIkyyRsoNrm0mOhh+NIa2Dyls+D
71GbffZJTckOa0Yv3CdHJBdb4bZcaFMs6zgj4q4Y46rvFJmjM+uTwxNpvqD6x2jTNrVn+h9AqDoU
lz5oqHgOUlAdndBXix+BH/dj/DEizsSfsnowF4YyNNrdao/QxcKLb6PKNIzKHgWxkqNP1aksM4w0
2XEnHDcP25vvby35s2V9y4lIquFWYYOJ2yYVrnKFEIzslx7UW8W/pJlSyolc+3b4+6R3f+CMcYDI
W//RV1dyjSANpa/5aSqt/b0+ZxNT/iJ2KDw4kWsZ+3TrsFq6Bpg65nY28X1/dT/NE7Owi1XzA6z6
87GLbqRrll3AIE6LYLe2ygectVGnCrO3JGZB3mENZPR6j2qvihA9cZujKzF/4Yls5ToL3FY5M6mh
1NXqbCqydHKVFWm/QQ/KZqYNiI6Q2fNVE0Vqb3K9Q8OLnpHjrv7i+GKlEoYntgS+Fcv1lWnGmjo6
Z6Y/oIlaQYfFpxMzv+HihHfq0udPLdASslIxHOnqVED/blMI3eYCtYCBvSUNWmzhQp7+vCVGoXGJ
n72xTm2e9+b/JjBoGc+Nq5JYDU5ltkmEhVmlzMxSHvDTVDZVbFs3wnKE8prFkAC3k63OC2VGtuD1
bXcBPoMUw6IJjq/RhYwJXAaai3a2ChDRqmd/7NYwPhp66eVI+E5oeTw79MfLM8KEVCvXbhSQmm5/
9NOfitjtasolRJ+7fuxv/pmsHW/cBpqOmsPEJEAkri1phikiIMZ6ejLhM9cZ+pA1K6bnkJsi7mvP
0Ao7KotQ+KPNHF4jIX/0sx1GpEH3P98d6aGZVktk9IKvhUktDyE1fjsRD+zzAosNrgQ91CsDQfN6
qKdtalUrif/y7FmsWQKw4IwTIhdL25pnG++j7wTQTn3k89Gug/jBehTFvAOM3lkB96gNtnBN/fVv
/8dQ5w4oU/8ShUTVq+CCus4Lpxf6oTaBN2plVpFjQ3CkjnKkdTBMHYkIKAMPwrw/V8JdVq7iDUn1
6l9tXLqk7n2vRY2XPXtuXQPKkrDobPnzTHNscvWw7dyHdlTZPhS5SijpFmyGLfQGcGXjQtKrY2sf
36fufDApKp5tAq4f9C2pQeorRb8VnO1yOQGksMPxN8eWKLo4w//Iuboj2rlPzsGvOhY02XcKpHwL
9EIzT93HXT/2/DA2dPe3krcIW3hT1ZBoBVbRSX3CJs0NlnI0by2920HLPxYkScaw7o/GUcriPnd+
OetUFe26bmJo1GGBCQ7TDCdCM/inx27KGDKciIekP2f9yVldADSGVcsyef3n00nSEABbrRWpu54q
HRNYaBc5aO73VXZ0+pEJDcTsOknzXHqOsl5ybOtMqu4a2WiUJLygQtOdqdmd5cLftMuAS/kXuu8b
OAn5Kqka6os5DQ5kRf5ZRFWOW2mbdvCwij4u9DQY0Khm9G0SUJKJOC7SGjMi5LNDLx3sxvvrxg/3
XdtUFFtNXuPQOHew1o6yMK4OJiRZ9urE1Rmrp4BZ9oF+5pZqUqrDXTlQ1UFLOPbarBmWmU4EplbG
V3jwwisWAfvjQDMqqk+gJOnEe2Q1N7UspG0FaQO6JQQ1z6ODFqr+pgoVn30rtxZxVMMBQ2tpqD2R
nWPQXc92/Bl5MCn95zpTQUOcLiIRoDWR2Cmb9y5eoOzuFBcgJTaQYwpBZkdVtLYtjEZogGEczeqT
X7vkr9tI88oE+yRJUBLn+DdQrT9lguXlCu+jC8QbDSLYz/cmaVCDZRXCAJJzPXlqOMcgnSdUxtZS
S6k9QotfIhu5R4C0PjVfwdAc7+Hl30GMR/de2h1XpYE5YI7YtLQoUhXzpNwwyV8BvRiLpJMkMadp
2H0OYNspOo0Sx0IE+xVNufcHrzzOS/pVYUpjT5uLocuT2vEHy+RDIwmqxMhR4LkM9u77DysZAzd/
OUx1fQVIrgw3UItG8BnN0EpAcT50eOaklQZH4Dch+AuceBq6VT0YBYldFqjr3IJovvuT/zxHylLk
srdp66TTE6shJPGpWdS3RmufZW6DGlsnsgppxwitJkwVSNZrrsY7OfbMTN8OlTLN9NtqZ7PPt/a2
esr8rI4HXkTrbenFVQn6QwZKyJMo6R5VA/wm+JG8C2AoCeTtkpbLZ4IU8jusBn2e0AH7Aa+qUT8j
lu0+CVSoRVp5IY8a06HcF+Cm1uB9tol2mfGqrXNlmRR9tVNdZqOQVdOiWQ67jOukEolbUiU/Oz2F
jlf3Z5V3SAG9fklmNjvMNnrK95UcZqaCG5uNUoIMegBq1+/wRXegy4i3i913tyfarRwJkSoMGjiO
3aniSPBz+hfKN8ogBTtSHXKspk+R2bUm4pVzhR2eLhTGd87fDJK1npuf3idW5L1J77YflBRB6TzX
ZOz+wV8cRDlmTJbPg1Tvh+jSxKrZQRQ0OC850iYD2BtG9QPkTIzOwUvf+6M0Sd8FoHIu8Lf3gzAX
4Jbt5EF/bMox04buSNwn5PXxx1dZQcGGenoUyBWRENnVoPdTnAWjWiU0ia78oL1tTfkaZqqp3fOr
EFGwDWsHcx+MusSf1lDS7R88P6pC1T0vNgWc7fwT/AU0aEKdtNtlR6xD+mA4BCJlff8oLeMr9Ieq
M0kpcSP76oCYEnBKAn1SktRfa3XUWM5w8gR0kEz0pfGMs1XzJ4LVUlax8zS0jrxu2RdMi7J+O84C
s5jQg4OfmDqT3BZciTRZwOBVIvEE+kmtQFDSgEXpaP97GqzaYUPcLdoRd458K8VzdTKq2grx1gC5
WbO9m1na0ZiliZfvf/1uvCuj0qQzn0u1DQiF4+PZgYwhgycaHJZPFAddEKNLVAluGQXhtHR9jhN4
9H5SKNcVUfdVoEDkiLSGCU0vienSdzBI7gKQY464eGOiQcbiW2haY8eM1Gd+DICAloJ0QxQYWt40
t5VWhmEI74Aqqm2PD28k5IgHBTF5ET8P3+WWs9W1g8x50yG5M2vJp2k3zoiJZ7uv1Fql/e8jSlfW
qD0L3/6MfYnPiraufo/WhNjrRO4UtVHjBTT/MwMRPKPJ6H93PDhJ05AEAjhrT6YGGZS4kPTEVyOw
K0+l4IQarLqTFwXqUlZO9ayKZdBkystnNmyGSpjuySOEKDJSAqL6FHIE7uthhR/HWjR3O07R67d5
m+8J974PRPi7SUOiHJzMegZw16+/FN9PBd/55En4nWwunLfB0Gm706MclRE7EOssLlqxF7jdcIwn
dXj+kHuAJPlwuamIj980S1ihtLvvjjxGmlxuh4Voc4l9DsQzD3Ty0VoNozFRvrmfzHOKcB59YxNG
OEiI+/khLEBWmN+ViXAemE0hSn5vYM68p7meXNf5oXugBhC0aDESkHIPF/ocjExeFbcT1G3SFJUs
62N5wYEt2SgpQiMtReNqCpCq7qhMNXjwRIQamWC2oBFb5adxzOiSdPLMg8JhRbnzyxHHtmeozdg7
kZGG3ubHp4i9viGJY5E86LsjkVmcXgARDfQRTkMvG1LU8nUw5pj+l6IE/PzfTA5Srzxwb/kjAVIm
TmbCEcig9ZS0FukyXE5dsiDUPeJNE7mSLsu8i1xHlvq7w3Z9xGwKO046X7atnCwbbpTpnprb3xUG
L7XSu1FKEwOKhlprBh6QtMGQxoY+txD0j6VOw6uTxY0Zod+BzZXLvLTWgh6J6AquIzfwMdriTvH0
v6uVqwkKE+y1mHAVvr/roXmgMRttF/GdtnAZjmuESQTIZpy4uyCV0rbCMKVqRtocow2eMYMJg7Oa
QYjaBHXzGDqHSFntMSlpqlytxLTvVnrVgDLOiZY3T8jupOcqHfO/+OC+sZ0QeTu5u1LlzhntCbXj
sE9BzD9DT+Mnnq0qxnqjCw41K4DHVa1IweFmeZihnm5T/b8ZRttl7bnDQTFajzSmVGzzsKVNPMWD
SJeifpPn7HQQJX9vxebDgaaEkGvg3ejBtWrNw4zzAjxnsXbsP3iPuS442D5lTUnMC40VO9iNfGXy
QWs2FQ4ImmO9tQuf9d/Ijtsn8s3wAcws/4thh9bF2BRyY9DYrMaYKolUFFGbKrKZooPYCD71wG0o
y7Cjx0eDzv9H5PplRutaAvOiTdGUBcsxspNuvWf4ZbQIdsQHnNjnLBugkeru/dQ2NcFWYGCbOT1b
b+DfGMjp1nwJKdUTFAYzEIWl5Tg9wM3Jn01sS0PQdnM5+H1AOevFRB2xtPqNUGDXPTc8Wz8ffI4K
vX83Mxh1qWt9+TRRSy9uwRO+UkFg/QuM9xxph5lUNUJ9VWN1Q7lqlrpl76QuZwhdlGZveIcmXROL
w8smuYY9zk2eZY5Mh2Uq/mdJhV6Wt/01+NQwL6YuSmn+xJB8zL1P0oXgnUqQHkiUnZ3+lT2ZlBzZ
1SimXpeh/N4Lt1nj91qRINUhjtbPEWGPMkwZobx4hu+2gEjwrHYTOS86Xsa8Zs5ZZNXuhfXrPXFi
oE2pGgliqt47hb/D4BqVNGYUmeFqZUGD8VZG8FAFfaU5gmrhwc5UDN8ipP/bDSjkhw//BkXJB60r
fdSzCrBLpS5Fb591yWCU+5Kh7pGbS5bvRqpFyJx3kU1rQaZ/F3xQndNiw7HjAAje3s8sWjBDbM21
hJEvFMD67tYMb3FcKK0xAtWoScGF9tD2fnCZeQJDnhyJhq6XdeiLfcH/36ZlJ/qP4GhV6jku4Urr
HVmtL3hrxnQO6fterI3WGAmP4R/iape+RCXG63cuIjUhtPqO56bz8Nhut4ELjXmGqgjKrERfWiMU
/JwGY5iBiVqbRAR5Y/JhtiTGku1qA0iN1PAPSB1HH/XjUCICrJgAPvy9Bw5nVJ4xT8dzgJVeYzn0
2WFvc4qkSE8o3pXRoSQ21QMY872F1gmi1bsy6KhuTWF7s7TQNGZaS6T0ebu9nONwwl2vDeBscXP/
l5b/1masllWS8V+5ipfc90ahtoVorh6eICSNAwyluNJezf5mJRdZyZD0tKOko8lXQ5w+u7Wsv0oq
gcMecCguLoG1hZ4yGyvVtnOla8upE+DOuYCLfNghANBffz3Rf7pwkvn8ap90jnERzm8of6S84HQw
L520zN2i6ben24jeiQD91GtsdPRd2wc85UwaHgwHUZNhepvf59wZ4K/P2V2aSfH8kbTIsGgisNCj
7ydxyy7r1C0qo948K3nkzqEJSdB+I0r5h2VWzeLUgYo/TLegry/VOEivfTMbFgATUcVLjWNnfSQN
aGuace29+y6jHxXhMD+K039EUj91fUT2LonAPSc8pHB7ryNf+rKa8Q1sc5DBRHJI+3uSYRVeaptR
53tS1DqO3WmLt5HykXYylJI2tMLcCK3hBA+jonjFaEjUAFSdK5BoQdXcZaX1HyYULC9mEHLI0jir
Px9bNwTgp8fGHDotHO7Q0s+I3h6LMAxiS5GPRAQUQEpXkfbKvt3jyFY/Qmsi/O1bZhCiNSWxV7aV
FvFolEd2kHFGwkq40uoEr99IKITa8732ZxKi+1fqXCqOJYQ0j/TeIjF6ItMZyFR8/GJYwF+8d+fA
FffzYbsEDH8eka3esZXz4C39QcS9YdYFNmT4V4+0cJTQa2SwojGFlVfjfRzmrNxTTHT9sub3DGl0
SeI4Vc0yeKLoBRi/SoUPtv0uxqeID0VFSdgmo6dFx84RPgWM5v29RO4V4iz46uUCdSZYFKx3szXj
j7kdSVOtTCCQAvA+wlO1V1hg+tqpTDdJH+ieKWi36RkHWzkxwwON5xFkUq5f9503KAeHyRkv04Z9
ENZTM7qGdwRzq5Aj68vhLN5jzxodXCqDCzrTTbduk4yPXrL8NPECwqyghjJyFkv1TjzsyNzJqVF4
mBWBcrDbhQIbWcJwZwO1vN0LVBCO6tbo38HgchajXZjphlzsmJ52q5D5giQG9Cm73+yeZfhUubHD
3qiHtpijrnDQ72aknQDiBLZeaF+lHIKKpisY4Eg24gOZPKWCP37K0EyYGYvT/d29DMSck3hXnF4f
Xmjr7VaOjalcaZrwN4sHr6+h6n8OTLu+lukMD1AP4xhvppQnVgv+y2JOlrQ0YOOVtvasCPyuu2zc
VEJwH6Iff3fg0ueCmZqd0/HM0VL/CsR32ie9FvDzoKz4abLvh93zGXfv6OFbg8b7Z1oqPjSMzfXJ
AuJY86OV0wzGyPAR32lyDUCYD3u8ZsAswi2iok7GwEafOdSz7MdID4QRJQYwrdw5LwYva6Mcly2X
roqDyKiKiiKKE3TrZpJ2VU/23CVqe8rgXudPdnGXPiiioLKMnZQK5BxBPmMdR+Ah7n53U/n/bQw+
9CCuqXfu2nOQ8IxUaCYeS/gtBWNOvXPOKDlXndVn6EYg9vzQMc7d4Myuxw1kteGw+iBdPu7krQJd
YrfAeDRvTcZXlckoqlAyWpAJascGWwYqu2v9E5PUSByfw3HIGq6+4zPbGtSI+FkIqxcgkEJWiUDz
FwO8JYmYDlyYupG6CGoaxmFKM+FwnUghu2+6mhY0TOEGRD+TPYdfSXWylIP4Rx47HlE/O+0mdaTP
zZqQt6GPnhOQaLwxgojUjK0VU62V9RVmWJc0A4XXe0mThmP4Mo8bMDUcoLVJjmcB65YmyJXjh3qW
PTczub0xmQPgAimqMZ/e48i3vRzIsJzUXDmiosBebxF8QaS6vP7ZuRjsDpQeBrc1YKWGi+VoLh8T
u2sQzPqfITHMk4M5gpF1q0yk78DGQjERL/ogh8MO/jQ6KRblfwFd0y6BKfZggXq+8+03yaDaqsP9
2gCKHf7ErOXfTyoxXqfTfj/mwJuf4F8eLuLoKdXk9N105n82+bmCIlYVtekfPprEJ4e233D6MdeA
ED2f8P6F5xqQ59Df0bLyjHpSr91LFqTdTFpVcYD2ASK7XRE4A6MwDB6lKIwhs/I1SDFXz8W2NXKh
pbTdPBFJGOE/fDM/nLLSe8jwGUg6ADH5Nq2E3qgipOrXZvtllSNL02j3z2iR9sxKhn6/hIBlITag
i8yitdmEWwmLHE/17vga0uQIgkWdlIwKm/KEEziVCp5oyd2HDf8/obpTcGEiimrYIwBBbQ7d/2at
uu5DwlfK8ZVafqmPO5JBpfjVHP20aYjH+kWaikFVKcaq7ZN8L+uoZ+N3JqdOmp8ZvnzUCJYmBiJ6
YeGQtX038rkwqvXczoUZji+1sFH0awUvTkMxdo1LQzmO75umhZxtaThCeEo6IG8n+G6Qr2oVvz4/
tuiV18Ye/NO1ZuyQ5Vj4RUL+ju6bLswHoBze3IqtNVSkyUbAF/FNxGibXbXqYC8kxcGo9f4tf6sb
RYYeDtTe21DWF82Ezav5jsCscvRKcONwNep4CKdnaMyWmomjzBrokbCeAt5+UntshSRTBGTVcBuR
TYb+3Zf+IWT6Dg882xUh1t6vsxocI1oxRdeFMsTbWL5CGDUvfQ8pJdpeX9OgrPEJyiY9EPW1yYYW
2GbgKkqrPdVRe4m/lHg80sE2PYsabmsPebazScXcIIYfwLtwzOAZWjL1bGGTdaH6L3zoTIzqKwYc
02h9BgYrY6K35SpvGVO371g87rbF6mF+uhzq0T/QS6mSGJjgrMxktJzzZrAvqr7nhuCrJ66M0nUH
Q822xgWen9ALHs5s59915BmhZJ4M6BU1jGQQPA1qu6XmaUOeSBjkJAadWRl8K9un6Jw634qHiIJL
tkwnSZ1HzaRvcwAXu3jln9E0ZlDRKs2XZyV98JOlv5OywM9lt/4nO/sKr3hW1sW+jkwlyWrJVIZ+
BVBaLUTNKTZTbsO7sKh7suCJlKlQmkN16aqvk9jNOUr9PJIgsdH1+M7Oh4azrgH6SlTopzWaecfg
K+sZzGO6MlG1IMxiWuvjGh8RA4Au7gZGv/YGPE+wMaeHIWcXJbIm7V503hs6wiPGsjuoTC0Ur46E
TxZdA7A2ktMeL1PzEZKuv764hLU/2pC0XSVURWGUpopywgAOGFM4IjQfzSE0fOqN5R+B3MwKVOKI
J5F0h91VAycXpAehx6PYs/Rx/fjarLI4dT6Dwi8on1qs2/AkQAnuEJrYSy4rNifWOlP/E0kun/MZ
VBlWwJmpA26ehx81iUc8bqtCJJUBCbFIQF0xftaketSjxpwAxg1pPeEbtL5+5QTPtCYkMkb39Mb2
TihoJOcVdUADxN2q1O1n3RGa/zvNx7JGM1yQR4i0/HGr/awqjkmsOXEw8vR7prVsrD+rsz2rEjl6
uSqw6Yvw9iYJKqa1WpC/5Z6OfSvkO0LpyiqE9iEBdatYp9s+R4/tZQFSyoD4qWPFpDZ5FaOneMg5
VJBB6LwlFiipy0JBam+U3UtpmiYAC0RNcbn2iGy1fX8QtL6tZDcZM0F8fwmBhZmnXgr9U1ntvyFX
QVGy1KZCkKixKyHFksNy+1GIHDlGTQgCAZAwLKhqSfMOSv+/e+lAwFkLgvmr0WmcW7PeKYMUwu26
E+F2fL9mpFTFIPCNYlnKXkt7PZX25Il9FBiK6qQ9JrPBD0k48Iv7V5PIOYm4yzDW4WUEUuI6c37b
rye1z4YDBRL8DqY0YNq4404rbsCYKuOhKWpV05I9oTkMhvBlmt0+68iNCjtsQIldP1TO7k5YwBma
Xfr7XFo6xJh4UKmp0kHHrS732tI138by228xwAMt6zMzhg+mbQxt2EBPVrnJU4EzqYp72M5VoMj4
DYSH/+sJ7bs7Kk2zMCt8wFIn71Z4phLzYh3uc4pxGLNIFYOxFAi25kOrtB/ZOCVvgkxAW3nUuQoM
nFZeIBVFO3lq3KxuEhLOM5JpsRHNAt+8yGyn0eK4QN2xtTb8NA6PXATEj1Xzyy2PTJ2+K/m0iAqX
7gpL5CfuB+3tK0ep6MZMjcmu5D7JeY5lI7/kxDag3/u7wOkeZ1599AfRzCaonHCWvB9VEJP96JfD
VL0d65WmeGcKZA9alpOVtVxFcD5SGOHCtJg48jn25U4qu7zxrIJaAfXjsvDaUBp0UbMY2I/bd4YH
zmxgynYta/zKva00b/CWKde7VxQ7/aYSwrpQ7d1/rIKyu/NuNbfp2G08uUoi4mljvfjJDgWQa4Y/
eqnZxumYLqaUeq/gbcBwO23FaCQmOyOXZDrVWkqQUOQ/SDM5+axtbjBqXtHarP96td8HQrEg37Q6
5pBrjz8U0cJe6GdWT3b7nJj3nC5uKJWNsJwHWTRLOoy0ygTiIEz7VhrDy21BH0+mz7fUIEAT6RS8
8VQog8WPF4C9zh3z6yIUtlgdHLWXQRlE3q1qe0SHD3NGCTPf5J+MZYS/5uuSu3R4izD1iErtFtx6
Dgl/NvMqVQeP9zaNDE8FkFExHmgdl7u+KwchfM8H0JHFYuOuWgJqNkYybf4bUp4p1vauss4XDrxT
fT3AHai6BIGZN9cJaf6BMTABTNJU6Lj5IAfhXSqngrrO8Bafmq9IC5mt1mCdkRkhY7PttArYH1BI
qATQv7U+VF+2u5A2nKKuAk+obZSbwwQszrUOj+M6GKLeAEZA5KwkJ5iEksQ+C4TEunB9yxkYt+Hg
tYnSUGLKeVpBTUNb0dhb35Llnwu/UYqSBlvRGD86cRr0JHQN9rgR5GlShwNTczwU0Bq/9HIht8Ym
5g1y3a2pCIfOEXhRlTGYRcAaSFSInZY8MILD9rt0zOWwDWlKxGN4sZKx4R9IKKx4yStRtLbAIXHS
5g9QZY+j4lZ0kgcW5Pg2IMBVMSixquHCMzYYfURsTKX0ob5TUTMVnUh9apZypBb0zd1a9BEMzqJk
Nse4s6jRhqsTC4oSP9+OdZcOFYhDlizrImZjTQkZUt/EfSjaFpUOV1JcWHDmpkKpG9LRpLg8CISE
IEdXf4Fjp5YxUe2bcMEramjB3I3237UDCcEY32I5risrQUlxmUpF0ktri0EDiruZzQHJxGLBPP6M
jLWFqLqYaY84NBvzch7LM1elK8UTwfiwPcFG0Ok3nHAj+IZg1Mo30RzLblFDTWJJdmRw5itBiasT
SnMMRhAsHnYNaxRqJ0wXIxYttYhpM0C6sQqk6fikcOj99OCD1ALoa8Q/OtEKVXJISzuNSOre8/ww
fE3VzBWhk8mIXrmX40hbzKUC/5wzI0rKVe8rgTwRo7Ji0fJZ7kPQ98qw3mSCen+dCQNhMxZMNJFb
t8t0HMJmm+Bnkg4Z63LQ8s51NccoZmwtWOOU/F3bkqHfKeOS+AIFf/JrLx65338Ni1Y9PRwiszf0
uHnc3Iic4w9EyLriJtHM+kfc3DP0j4Nz7WCKegD548MbxsiMXQaC4xmblUVQ+2JI2VABWRMYw9o3
Xu+WUDySw5droZrhIXFGHSy+e20aZO/jSFQTlkcWGPmxUN8yWiDGkmpbIbOlLmRbwAzn/GesaMEx
y2JgT0FQDTEXRhfDXM4rnj3q/ck323yDaSkhcROHk4KzMuZ6MHMkWsBTNMf7Jc0RkOfNbWW+siG3
rZ9fSlSs/yJxzE7jItaWBFVT1dvGgyyOy/HrTLQ1vBBAxJA4XTo4y6Wi8y01mWzxrxqxYnV84Zok
pDIMVDSNCTq570dGl2jt6LgBrvgJhemx4xEQldd5JYETVgIeTQmD7ekF1UpOjGP61gx3oXvmvpk1
6QS4U/TsWXZsu7wj4s2Y5+kzeu3R52XcI1uEy8qONhrv2SRlaDsroy/gmMgAkjrBC27kglJg5hQa
nELp2d0Uw51n8e2mOEAY/NWBPMQXUa8rZBdZC6/ust+GNRZgRTnwtpmwLwGC9uckqhJSfz69tI9R
zsS7nRsiO9loTgHAW0/SY2FtfaaczLDiSBMGZa9QX4SadkNJzGVbYts345T/FhtVk+U14oAgxKXr
bCpro5/UNeJFdykBMEjwy+spLFU+0oKNyfFfwgWCkQq8n9fakGwXiwFN/dxKlmCXOrsKBZI8FSp1
gXPhmzq3kKCh/gznIx5w9t7siEMVC6z7Ej89qVdxCJwcHaqLfsnMIXHoifAX9SsIVyGqCs8f5US3
SiY9acxD/DUzB7Qxnn535cDLAsX9nwKWpTjLujMd87+Fv2QYMwKP0volJG1hN3+T7LrGAiHnICPh
pSZ4N/wo4pVM2zVTSmDjTEyXWRgoN/T0k9zocKaOB8A2/weA6mj/TkEAHibWfHVgAlsH0BTJaSK4
tlsrxa6rbVt7PuXfBaw6eYsV/XmGYRz1o8zHYPIGdpWWAk0RIgsHOtqLBOr3tu5HiFVKRtodPPE0
fcB4VUjMm2Q1Cjdx/vY+sY9ADXs9DRlsb4RXCUdPL7kFxjUcbySeVGG1bSmHa7LDj/nw70nmtQlx
kX3j2ui2Zu+NH9KHliIUWOEO5ai1Qm/QrK7gT+X4QoenjIHFIqugodAtnGU4kdhKcue3MswNWv8a
85sRB/LSiTIO/UcHyXAsmluOjCTfK6vOFrpGOFAyhJavq3FL/QkOIk0QWLvkoj7NW/JEhb2+dYtF
BmePR1XYog+7y3muMsO7tjQkXSStNrWPJi1RSbNWhOQokOFfGMDCLQGLl85WIGPRjUcr05QqjevW
Yvj61zfNY3GgZL7HwF46nIDu+zznhABCrh/yKwGaR6mfFEUFnRZPEb5DTcHWvmXsTMIVRtf99+RY
bwWZexjAp/i5aMqJfqJ5Me27oqnmJ2zj78iTq/1fhCegKFUPpepJ8JvWzgXMo95MAtbLFj1ifAVS
17zhvhH/GYHFdU1QjbojIlRmP1BaKEHq2Py01dOVX195SM/kpQCmeiVolNzXAtDkia7OT4Yfxv+b
hsC9l3ed5QuZ7ORY3dMU7UKsc/AhGR74+8CxC8/Wj7CBskEFF04+Z0ASbbXX0kDt2+/SiBBMTv7n
kwtZQukb6E0j4WpdBqFwuX0+w9Z/W/NYhnH7mNfDGDXHmXiJvDjp5pphFIeodLyBUwMT6fiZ7xkS
Hcw9cuKdfLs6RHifzyOiDkHuzMGtzibOvObmeAMHnHclDjh/DKD6pyNHY8PGlDY+yD4qAoJZTlLJ
LgSFDeJffVeZppQkzKrBUIn6S2pNngnvx139oeASQt6CKWDFwrMtw5LHkYbWgeIX6hlyg8Uzugv3
JKtWM0v4lxUn0qs069lZE/arWoyqxyRFC1DTfBqbTvaXsfPuym9cnqfrvQr8nPNajq1At9YFZ7yv
NHLSZSGiwbvHTXD73QHN0AY9v24KqVRmatal66nUgx3XmgJWElhpnilOwNM7H02JkxU9LK4Tw8hw
2B7pf1wmyZn6B7yH+vBrpE2vQv6nH5zbW2QmaUJobTm83RP5ciB4fEbl0g/DEbg74034z04ipizX
8S8dl52S9Q+j7DGIrX4tdTvvTSQ2zZNdXp2Vo4lxgvF/GFNdPGwcBWVwIHihNY0+jJ9JataDJ8qD
c6YOgBfGlpthKKkN/i6WUgf3YSvc21chGTYMPTIjmKM7RkX3pZpqOSQm3qlN4rCXFaWyYYwwUEIZ
vCidYhm+thhbnUy4r6tHp9bvjDW2fduLoy9v8mbFbiHmSzZVzWcHX58IEbXIohzstDSfV2aU0Bxe
lwGrdhMDtJ1LbPM3VKlshfqWODrxI9vuwytW3ITpgGm2M9pPo4RGRaHQLNSbZWYowFXeVH6VsD5h
gjrPK2Wwz8XZMHqrVc3R3zloTLmCWlWD2p0K+9fpoGzYPmp3YBp1RKWMKDVLmmSccfH6ZAlMB6ON
4v4V/wQ4JWJQswtZ7zNBQzcZXri4S7YYxh9973nWPs4NA7EmEa0YLN6A1v9dqcBJvuk0MZVcXNSp
Co3u35o6rRCKv17JGzz7RoSw6WUnAloXzg39EjfQrmZev3fsIut1/nWaRRjoA8rd9tzLEftENHeu
SZ6dndsPMNusO0e93aHzqMeMZ5nehSFWvlh5tgW9kj/dVEW4hhfsCr72/s7GSb8f3auZuYszw9Eb
L6jQIu7R+P6XNPAeY+c2Pc+NsIRmiw9iaj3/9XDMycWutlDS8T/m4OUZcYc/KU5xEZpa+iK+sw/C
0sRklOqMJawfXJaofeiG0SJbuNM+AMWyURPYwfCtSOmIPG96hhYdMwHxVHhsj6sjGdKzNwcJYgBK
AyZZz0MOSH8BH23+AIA321OawmH/z+qpoPhmSAe0fkkjtSyYYsyOIhZyTS1mrouOGcjChBClA92x
89WVPO8n35hZtAB3eKgfUC9AnIZHyjjhYVwIJu/mI9UsH1Dse5TbOtrJJi6yP071pVb78AFfUZHA
40zkqokOMMid7jYGiqPqhezPsObfs1UE9rN9hZD4vCOfd8tYGlHycB6ELD4qgNOtTFORZ9VLrQPo
uxpBdBc0LSl8JWUwV0Z+osL6k5MF2ch7qBv9aNyAjIF2e1EGTz8viYCPXjhF8Kp8VN/YR7AQjK35
pf9MSi7TcvPY7TINeCLwtWONFG2KkQ4athdkcE+zphRh6lfWRpZe9bscBd5QYMpKklHUgFLKdNis
FFYpQnOZeRyjCLpfbt8EZPw/6j+8RjMTpxQe6MfB07yu7OO6vE8PsR2TY8jHk4CELVo5aFHBq4eY
X5Bq4UiOWKKJL3QRIIRTS3gc33gAVjZnKrBAqCJTXyrtjk5EqIv96rtH9/YIfH/6Wb72L6nYZXYS
86XRlBMyuDFarTcWcM7sQtSunYz8SxRcpfi8mIRE+n9YGoUqnFayUUowT7a2n5+Pop6MIONAYAdr
zcMtLV9WaYYu34EYiTU9uBMzfHsmMH8kP8FEvEDOH+OI7LYYwJenELBfHvQRrIhTLj0yCAYm+Pu5
EXuaSaT9Qmz1eS2jXgdrsrHFp/0QBsLmjGoISqaVLL9NObk2ip/5IXzNwue2R3wpS4yeO2ncSWNy
9XjRIyizUQPdYUOhjUZv5WhGswu4mXyv4ckkAu9uSrSqkggmKmJY5P1piGoh8yV/5UYx0TEDdCDQ
JDGemdqkEi+x2I2EOPIrRiq/m3d1+QUoWMmU/K4CEL8JT+MnOrSeejCTZWzbi+OmGRHU9/MfiZXQ
FJvkV1tTllCyXbyF32+pEvUFoQ4/vupnnsm91/kLJMqlqg9KWqlf8f+atmyMSOnXcT/MXyOLyK4C
eHHww7R1Q0fprYhHjC7J1Knztvm0nJBv6FXhwGsFFk2wpDeSCQ+CXEadun8iWJy+2t1urZNWkZJa
vRXOAn6S9GF+rJlQVOrRoB7HQkKeDYm71tkE4DdlrHNTfh7vwmT7EMuV6gCGFGDP7SSacbidV82Z
K6xnMA50qjesQ5ku9k73ltcOFlisBqdDstmGWX+WfhfCM/UwTK7VRdLwt/rFbIT6ltQUWQuWWTsi
s7TJrqYig2gM7olkUfFVHUAqTSUJerECxkOBKNXxQL8MAbEauLchJ3uEwqrJBEFwvZvVxN+N/Ygv
71Ct+7w/NkdM9jeCI8uj7rFWt1L5cSn0Yt92+9ug8y/vty+MRM+cw87Vz2Py0fvcvsucYQM4HRAh
C2EBz3y5xikbisq+rczd1OmB8qPpHKO92nIhZSErsyBXhicCzg826GqjVs4zwV3zukZXkEdeNLfs
/nwki9XePb4AmblBKZSkGltjKNFOMteB0U/xerT1+I+HJChRDPR9JLExx5U3uAmI16vCkVXSTXgM
gndTqxFChcfWpcxKyOC/Oqz8nLchL+2/ePAPdJguz6xIH9I7uOmt4LU58OQLpERt0oHG8a02XFuc
2XmYWGZIVQGCfBbJh0ycOUpdAtfKkgxBFIao8QWnUtJ/2tSZSTi6mVjGof+z3JlVk994GOCUZ9oz
J6ay/OS+DwVP2Ez273vE6Ol6dpg51ICa7pLW6yAIWFC52Osw7uyzJYaDi7jtPXCeNl23Gbewn7P0
p/hXAq50DeyIibezhDNJGF94zeuqv1csuJFSJI5WXSXWF5EFgniQbSKAIxI4iqOPOjw0zec04l+P
513WBvxr3kzytkUmEWfe9ZxkLMY3bFp4qcdWNrGhbDdcCzYwly8BwImqj7QTzUKnJ4Z6jT4Wt+V5
yV9PSKG5+cvpbr5m5nMsLEPjaBKaBw+mXkYvmgBEcNoks6r3ZtCTfLNVVIOmnMIkJnURAJQLYx/B
9UWYbUFqcsKuQmEARx30XqFyPfLSN/Oqph0ORsHlpTiAXOaZuiLs3hoIQQBjGmJTz/4cVKHUVgZ3
y2N0KPa6FO917OrB7vBiFZxYTGz2WjX3Mlj+d+93/dGYWrlpJ4T/eQE6ajB9KSSXrB81xfKPtRM+
KAD5d8JPjY6J5zrPl9kg1P6V2WZNSzWzNr2Foof3UZHkSt9hrKQjDYdLOLRv7fE30iwKMCuw8bT+
3tcFirfvd3SSIEIDvDrKQ8Z72z0W/DQH9QRLcLYUTFgSjFHe68VF9RuHe6A2SAvun+oLV89goWFd
EfRqhlaij32Dk1ral0eqhZ3o1f611eb9ut0Ba1V4AJwJLkqRFWvTDR9vKv5TkSDMAIuP/ubwhXHU
SSY9zLzELfDGK8fDRmD9zam/vhvyXJjrkof9//GT/30YtmGJDt5n1TJgqIrZ+pZInv0kPZMvIK7e
og0HOlQDTp5TH11Qrr0+zq7dunHDJtj+s/Cwh5K5mTUHpc41rIxGbpZC11/4+iskXWbImcdT07Z2
EAO6MeLnieGS6RTB8VMlxY/iDfgoZ5tfJNlFBv8XEzGqhYar9CAyr4Pl5+E8LBowzjYYqSCRJhjQ
1dOjA5DxFnjQWdVo3/bCo23v53jnYO+wq/jN4wqI+ro1SaGYnYv4IE1c+t0fKzokkKaoS9Oa3bS6
dkqoOhvv9VGt6Z2YNLKA1VBLfOccT5AALdIzTMJ0MUYXAVsjr8NgxuuPy/noSZSxIq6GcMCp74oY
XqikPQ/jVMfZdohN/aA/UHf2x4yCH3VJjpPbypjIS8zKc8YATAbT+SY0BAi7W8Qpnw0ThN0JEbB8
SdaRjMgbqEoivDXBsb79XO/ZYl6LJ8O0N4ECoYFKh91lR5lx+vkJJdJmSVIDJBUmG4kNXNlAcxkE
SFLJ5ehZOya4zpQmD3HgKa4XJrgUVut6WGBUiVEQXsV2yykS8Apt6Ji92XktDkPQfevO9/xqkah3
tmc60qHXkWJIXL5NjZNa7b9C+UtYiWev+UdP+6IEA9GP/ORPV/GELNapeUT4Cwaz4TOk28LJ235b
1QSSsMTGCTvNF8TENAMYBZBgtX4/zIot7Yd8GHoK9OWyLteYS6DnO4zmRIw0cuCPohbX2swgCc/P
GVctVsyMcaTnnr6roH95UgaOxdnla+mekQDoGYpDuuWfxXs2VrHcY8BEYkWMorUcfpFY+g3ZN0P/
nvNfLDXOGp8ePhfXURAzPsd8MxvE+sXeoZnXHul7RA/6n32tyAgY9hhCN2r25wMWIHu5BRyd5dg6
JK4Xa5fL/9LIdUGGWfyQRFGo9oqdk0Bt6ohLj6aJHgT4CtvPCyNzJ2gPZkzyy7nZkbZ0A1YOOnqF
3lcynuhPjJGaoalXuJMi5XLypvJ8FdmWN1C04deMSn9K2XA8gRG+VhJz5Ah398tn2fPeomSqcAVZ
7G/QnwfHPmavZ576t5pBO6fchbRaGurv0PhIvtzHLFBfsXr1N1oi3M6k0IswGBO+HAodapR0VtnI
RicNN9TDhnkqvSMID+PaOzwu/iDlagMnF6s3WuE8lyCbk4bLMNpbnRncvpnW5hW6FJHnQkVYF/e/
kyrXl4JWUMAg6DHaZ8Oa2hUctlW7T/0zqmH86+nu6eYBQLEmwgpw2hco7O1FlZoBLzhJONb6Z9gv
9o1t0c8bHheWDHPnVmR+hDXJAwnua6npdUofEXybpJy8vd4SA2SyyO+xST/vrioJmjPlmpzbiax4
upa6VhC9D0I0znjJpx0ki8vNWjP7R6eUOLm6ACFn/FQwouJ7TwmhMTyqsT6s5zJEIpYFJn0iHOEC
7WRoTU6t58mNpcQl3Y6Lx6KS3ZFDTMYtDzVRXfOUnYK2vsmLBSCWv8f1POhBglig0vq+M8xOSvbx
QCg3DfqHlKJwpYqbzS6VV7HxIaLwJqB5wz8orw7RPFMq09+ljD0CPVz7U+LOXZ3XpsmTczLT2TRl
klnYei2Wsqtm02C47dlWcXl6NHeJouyP8wIOUpsvST+76FjTYVS5vri/4RrgJBw6vCBrS59oZVTU
hy5ldxgF5gD+Er7gJQSmnSjGHjHRnoq2UhPlgFIiphLNlLPrme6YLPx+LJEn/QdAcEtdmorn6ydb
0mQBKQZLhGWzQp+yYTdpavBb+wpKkN1n26j+dakDJZ8E7sCcVf6+WIfKi7UB0TqNNbeOlkEqoJuZ
h6Z265CN9TdZW42chsKZtlWk0bl1Pt46/er8KoiS8u4rIkmPR+I9/1bfiKpcp9mn0zGJLCQx8Xoi
UOzDnFtp0tQkKBFnZPL96H89yd93qoOkZGQpxvHog6oddC/HZVGBIz1XENdmCORnqEnhYCUpW3fU
F/vU1r0o4R2fSs9rR5itZHPENLQSfhY9hJh6or5XV4Xnc5IyB6h61I6ClxVjsCcbXxuG6piZYk8E
zjvd/tRaruHjRuYkymSLEeRgs62rYnHAaVUiFKKvogb+QbyRJqG2tz74B+N3uALjEL5/gUQf4hy4
7E3sAVtAbgX2QNUubiQht4lX5f+rYWEaeTcWWi3HCdAOfj5ttsbKTDFDH0qTE6QmHo9uI2IKPHhz
K+Ez8Vsl7ifJt2cxQKcXrpYh+zwZQxOrTzCxb/CdaAHUHhu1zPwJh7r+mdOyqiueVVIH4pA72SEk
yc0TEkMT8SvfFzGpdMhkDfLgErTjLI0+Ev2aVJrSEww4vjuUQdkctrC85jUobZtwJME6kb6CzANS
ZdxwL2NAEk1zwhUN/uJLWDfuekkqJqn03WR8082mAKh1uedkPx7ycMrkZGk8fPZkFUikfGevda0J
BF5tN2tE33gSSy7QBEcP1xXZcYixejJwGE+4g3fyUfUOwf+B5S+So9jyEqojUA4q4MyRCDMbZVot
8T32QWtbzaHfjKdJ7Uao6jRSW2doLtnuj23kN+h5srPLxxLbeW6GNF9bIQH3KbvRgTXd8mp7YOWB
w5dZpsUtSXqQTZ95AwfQZl+Z8j/KGInRIk+mwbZyzRHjnpXwN6R8Vfr/yaHNRIZBiyHSQcSY8DmH
RQrTFVhj/DDMiRLHX6ZjNlyGURUpuT6iBs/nVXOsTZ2MeRV9P+50q5QQlhJczMX0GFg7VkmfXPm9
DNpMiv1gL/ho9ByQqdP2d2YHGux1T5XSuuEK6KI0pL8icgwYt93uU/C56UuoVCDBNc9zFGQTt0le
0kOkszfrn4q1fXP9oAA5cITQU8qHuwmqrpVAZHSX/7b4otZJhiFjm/2l60WLj1dvihaqdYzMrXxx
v+0FSrkVtRm+0lGBPkp0baelkkxfWQpp3Zhfi4Szd6WRQASFzOZSmkl44r4pvfrlrzKmcjP9ljk6
m+6asARefBsOWZO5BSft/yPnf+1iV6CvvTqAnCgScdw7+i3RRTseEjtGyvVoreahlMtXJjQ7USGw
kv1Jl7oCUB65lo9ounluAFcfnmo/ilp3JmJiIDwxiNsmYfQ3QbdNpx0BHsDuy4ORlr51IrV9tEek
OaGlY95q46hfqSTOh4pTmKGLyc9+QhDqDyS+kOvA9ZIMyEnNZ87weC0LcQ0JPxz0y89bcJ8b9f+o
vk338ZLJIewCjVkKJbZGMYHc4ANvSirrYZB/+J5buf81f02na4VkhX/EW37iVJ9xMusHvPPzazvD
JVH78kR2wh9ezbIpCU15y/j3hQO6mqt0wyf+ktLCmuSREN0FKffph4VfHrNIfS4tB/WaYSHD863V
DRTWk9oPtAi+ql1OyLQU68CrkfkKjg0EwDHl72XOatRZ+gIFsFd+gAWkgy8RhRgZN6zRtY7Zdn0R
1i5k5uAxynQtl0aSHTGsdEbkFtCXTOzMRtTtn6h0Wg9HO7ze7Pbz6Vmzg6+NQLWCR/6ezMa0BM0Q
k8Yb+2tqVqV4ZxLegQiCfjT3MCG7tZ1Zaa0AJauD+0WiWmQy3XPF9jikF/TIv2y81VsDIdl6UPH3
a1CWS825jl1xJlAxRHywXicwTCidczCOesuZ/oP0S2EXILS+W8fUqcRvBfU2JRrq967SFH9sjXxR
Um+a6pRQ4UL63isTcbDiB9IyizakN15/tX0Frbd68RwAhsDARgNMm/ns6zlvsxnX+3ebyMKP/HK6
vEcfVtTk/6btaRtX6TQjEBnA3JGKxnmOS1XKZuF7OdiHNJe8xXvECavyR4rpxmMnc8EV/Ggt+eV9
LyzCd7JbnOzza2B3dTvH43ET0OoEgPBffvxYf4Vm3SAO+C71jLgATmCwDjN2hC3swiDPybESjT4J
bDieCzYnfHYNyYk94GmVXJMgyQYitbufsxPnalWVaMFDusU/CpLWmbljh63oq1eIrx/g8LAXCDiE
v2lM35bKXOqFKcvHRU/s5doO2Av/pcMiQdvwUKebCUEjjuA/vjhCaBfX2/WGOaKR0MrH8TUeuR24
1TGnO6L5ATxm3J7c8ekS+SVdwFCSwSRr4AT6kM/OBAnuUb/zXHR4RECkvve1dnjzBh2T6rXqMLb8
juYrkT2KU2CZQ53jLMjGB25dv4hKkbi65ZbXASAKJpSP9Q9MEU5gE4mYP/0tlR+RJUbKq+02uXZa
VwyaK+455GWzz/nF8cZI2bMBf3yQdI+/7mCdJSlkvHIptPkIxYVr9MzixI5RSfUVJUui/F2O//F5
b127KzvlUB6+HNZVnjmzngozfqJOfaNSMQurrAovr+PyvRUD9bZt0lAPvZEzyVH3pL4F/zumeSTI
zLeP+pii+EkBulqcx8NPyOyOHOPgaZhDsR0xi7MZ3MwcjePrvfEQ8/qnrwPRhpdkcl4zEtH6HQBF
20wdJiutJyYzASDAeZdlTm2UJxCKGVQvsE9RwzujKI4pX5OqgIQKUqvBgGRc412AtCKrwH7W3uw2
qvEcMyo7/J0yvYr9jTko08IIdkyaITbj9hO2CHXIbtrEv+HAJzDzcTZRiHaspT2TQ1dP6O7Rb789
p613gjqXDPnZgaFjiS371wFqC3esw6B52+50q5VnrzpoetPfo/eCRa9sVTNPPiwzmpORH4WRnv28
MYAfr3MdFWcs3aTEDXQ+xAI8yxmcc664FpSBll6dG8NQ5LS/fbL5+dbo2QgJXkKlw/+1V9TPIIcj
3Q89V79NdZv5TC+j5UoTKzGjZz+zk5ssQ21FnRUhtYzBEn7nW95967WzW4gWa2TqFAIL0afeAmNh
FixiKzOKUUVr5y1oYQVdi3A788O4QHyCXGSiRzhBQrhyJTrGivCRHhhhIvkkoOEEjnE9mrrO1Ln4
t5DuDRD3wuNgkA6KfqYf6A2eOav4dNdLK5EdAdHDLfilEslsqnCRTSDzmwBazcu7D6XAyUG3oV2Y
LPICINRVpXLBa1sUfcYQa74KdOWoayQTfXmJBFPNFeWrGiZGvnIR237CVH7cz68Wb0zMLgnYJsMx
AxL0jrk8CjUJfD/m33CjeCzpjKIzb5Ogw0jc8wDM0xx5KGjGSS80p4w4aoZ7Ea1QDRw60RlSWk4v
///zbEDmv0y0DK8J4yX52VC2cOvBXYXP8cRVRkvg+YX1L9044U9b4eEN8YQpKohbEedmMjIcsauc
n5VqwT0Y/6ItGHLzpXe/VTQVIgGOnPbuaDGisEHJh0dScMA3i3aihjxMDVzMAwuE8iSgfm6f1GcD
wkh4AjKygCr55sK1m306DcCLzjTV+2eFz2KOO7WVKwUsmrw2iHTyiqx+9/wElgp6XG8kPsiR2t1R
P0fM/5RKJ+tbBdWaqpRxt+KnxwY8+0PXsD6SzXSu3wvJdUGLC+GEmPuFgBuZL4iGfxbqv1Hticn7
6fTzPyQWjmOW8XD6OXTP6YYbWeYyfPzimcjWHDttdaAlANULTxlmDvCiV1D2/7ANr2vbXAKJW47M
P9jj7wiVqgQwW7Us/0wi7RKY0go7BxRGihG2siuD5nRR29BnhAtil/Q9ekBjjuLpnA4wZwvwQMlI
+aAvNEpKXnbt07f+sPYDJkS1NjjBynftZk1C9jfHfHmvONv3pAjfx2pmQ7CiVRZHp0CvYnWTvPwM
RVTN+TknyhgVHD3ks5I1MmgoBRfqn+MxkLn3hzyHCbjsWto5qhlipV5+SibQHKPwiKDIP+oOUXj1
N97qkVcTcz9t6Ubg/OuapsndqnFELpnEWTlOnjS9klzZxnuQLqQtOybYdVleQlHAPvu6TPoqT2ML
Vr0pHv8T8NlqaNmvE3Ex91NDZN0aiXJ5bF+UDXDFCBSmVNkLQouYnglLFKpGM7GbqU68QRn/ktFX
YpplR2/giFsbn+xi60caz/Kdt4ijo+lkHtSCY2RHy9mf1++7IjEMQXqvLtQ1LYmwKiHq+QKjwMb6
ozdYzx1N5lxcQyGCJXxsD+GcoRA+OHtJH9XPc93XEHQ8DwZWPLhd2wy180lxOVIFt6OuWK8XLdhO
PCUcmWL3VIrqMZfs+Eicp/wG4gvqBNcoOxnEqPKvCbVgoiK53YJHc9jgkIc5cuXiNC9Bm/0na6CR
qgHfWKpHq+g3PeaXGSDeHxIWUHyQirIAelgUPlynqG732eeNyWV06919uEdpZwThzLFipKdnZodG
CLS5GHlkDRs5WhPTQR/wX0cVpTs/heRaIrjzmHKAZ8uOk+sO/vxCMPNaq8ZLw8vSFkNDsn25IEkb
mWA3CMV/5d/+A0gPjPVqHhd3QkONz6QTU6XerTeXJ1cGXZcr3clDnQ2bdobt3Dn7X+p9Wx8TJv/W
n5Yc1gLKWPNzFwVC/NunvrUClgZai2vuQJwALbWrGKHEn9SeDoNf71dGj+RFNikQuxtRhz+CZ6A4
XN2WbY5qwiqik9qwW0+NdzSszVAsRLaxiw1jyq8jqQtiHHBkKXExI4Gnep/Vry4tLcr2RYKL4NTp
+min/ehFMeTWQ+f+gUbujMFyrid/Mpcj9gROaT/9IP2pUBVN7GKeeCd26d842KuR2KH/iS25wu7r
ShqkzdMpnOOvqC9vzwkEEM7qu6wiFYzuzJbSA75k0HH5KxRU/6hnm78MF+XXCR/5mVcouN/JqZMR
5zgpfwtjZiZvhHFShleae/MBWK08OdQyb3BxKmHngV19L/Nbk4wRx0iMXmq4y4TuHEyGR+uIEl88
qO3mP1uGRYcJXxeVY6D8VcHNdgS0tNLpDSM6aZvFBO75MGqsoiOKgd6MZO58rj1c/fP2PZNh2Ntr
PeKG2FIDfQpKAB39p832o3f0wvWeIBV04sJewWMjxwXx5X3x/FPrdB1e14QVnrxOeterHeDGM+xD
rgRmEB3jiLbpq4L7VH0CJ4FEchiDtvSXcMTl2iDC7WLnCRXskN0KTeyOjmbfS12BSbFz6eBisfoc
JZ9BrOnHuDvzJfGEY8wTw2qufk1R2J34rGNJJy8LcksPworfNLiDXa/2bl3FxKML+wIYtULC8dRc
IbbP5boBBzPR0ms8S8z3CfqyOvH0e00VfrsT4utvt4aPFWkJqZC4flLAWkJG3VqaOk7t8429GQZI
FF6i4O5FmXFTEuZk3I+//cY8juP11Ck2v9xlOvXyGvMFWg3dCWhRHxGdWpgOdv8HTEO+dF+4hoS0
4f2g96iNn7HXo8TnUJ4lQhqpdjRWPdEkvXBeTFlBmLmcsOhqkj7EtetZNNDLMie41pjvpOpJEsLo
F8bT/06sj1vmzTOerCzSp6tvZBtiJXUTv1rMkLCYzEut5L8qKJoG4TJYzBCLwdHdc4/h5ySus62v
OjvK7yzZHaDHhTJefkYAorKDZeH3Subs2MPMugLvVxdN/1tnnbHhTnQufIP2NRo4NmhLapJ5hF/7
UQ9O5c2KcFZht9bAllPQ4rwwAorsmIEE24ClKyCGRL8+B0W0mdz6bHBDV9/YlH0ALKa3W1L2rGh0
yfoW2dvxIGnmxjf8/TuwcRbIpspJxrUusiX6BEzsgKTq/xdxsXsUDN37OpFb9DkF6+VjzIMfED2Q
VFH7bhPlOA2e+PfSYSPUHxaxZRL0pFFT5coMsVYO/p96RxoOfHYPjTDBRaI+eYT3Q6Z6sRrWYfFX
pF4g8YE2MQ0yRYuBcFWmgQ3oTmgdtsX+4DIdodKo7BYvYyQDEPRuNOE2YmT2OkYsUoud6aZrlxxO
p6R8AwiHl3Y7nMeCIPB23rwo90Hr8mGl14pzNa0UTUeaEfblTcTxOZtR0meYyCdIbM2Q8OiDWksJ
CvDneUCsJ3KqdE2D8mgQ3Q5mkj3ALAqy8yTH7ApGa6lseGlGGhfjLhWmqLY/sDrIIeh4tmoLfCK7
ZGSPAnFiKdXPL3CAkSaRyLXbuPnVMB7LRfm/awe3RD2bx/gSV5ZZfjnrpg5g8E8SmDy2ilRLzu+c
op6jhm6d4D8hL2FxIcQRMsFhbK9ODGmAGQ0EQ5IfaJxClyfHWrQWEYxAxili61HSbp8ttNHR1szq
P+Lfr8PHtO2xPIkYQcNjm/cZCHBBOvhDMQoJN3MYJcSfUTWNZop3rhr4mbP11nWRkpnpykiCYXK1
So1Ngs9yNQwCNOHqjxcSoR+nYjAnmRpyKkQXN8DW61lJVLNDAbZ4IzrSIzVmqjmYq5pBXPqpo7iw
Z3VEKukK7RxhJjjt8SLhQeJvzdh9ZFsX3+zjPUeRy2SIZVuyKNqDUTXoWNm+uft4bsig5Jpd3Of2
kG0N2FEDX6mjtynpism74nId+F+i6SVEsX8pyD4R5JdhjhxDqgDGMcecp5z/ZbQRmvSRm1kZWDhn
RTCzsqIUzbGPDDQoX8g3zmoV44ip2sxH6oLlXLqEmNO4LsJ2J+1Ec07frUXLzNpychBm/0TJjXb4
NgJ4zbO+q+9+w5TJb56963seqtx/+3gYy+UtRf+InaeLQQJrFMmiHd2B8I2JWD5poHz0qpuFCns9
h8hkdoTMa1CCSHAfQYtJ1jP9z+lWgVEiGMJ4edjen138pL35i4ocHwd9eYYFlqmc8zBxYEBnFG18
iU2RaFFAT4C37zEhKHa3Im0/LpfxhwfD4k8rS4fKsyxy04P63Fe5+lNfcWv7VN7U7SU0BFILDZgS
vdz32bZbzsk1Fr1NoPtiCKvd0Osa+fAqu3l+JoUOXhgc8laDn++g/5Y/vrDIaJZoxnukHvVFXKnD
/LEQt5webJ2/RdCl/ugbei+fZWhM66qf1mXLK/3tJjHrRpyIXWXWhT/uZGsG7R6/FuZ31BriFLm1
1zxPRoqM4fkce2iMx4W6MLfITcjaHZ365n7zzxwV98+UdZ+VCLEt/k/xDxWg5hY/3hpy0TrKaJsH
dc/iR4XeIMi5LsOcvFrKImfSinSanFLJ2i01RqRElz1VldpWgrxOgq4cnfzE6T0f4aainlkVFHL+
J7XD8uOk/uGoney2v7K9eiksKEuELHhXnNXFygQXJgroAGI/Nxp4A0/x1XRCImu3jXHyaXznHLYP
qZTxNVNSrQkVJnkUP3CY8LqT44Z/bwNT1FKwK5Jt/pLD5sUFo1zNZJKlS4UmOWtLfvPw5BFgmcqB
JMdpOHKUEj4h7GM5vVFhhyxz3T+4YmEt40n58AXaJ6rlCqTzU21BS0fnbB6q3ykm5pGv2b9ZakA9
sGBQTyenPT8HXEbzSwbxFZUloPfTo71atfkZolPX5AFnWspUYeWTaBaGu/wFMFdJGGnFcg/2iqdZ
bU9MHENFFWB+8rIb26Acp3pbUEVX2K0DB0ad+ITtoHbobjBS9nR4PZVI4lW2kyKFJSINwg/Yj3Gx
9Rd18igrbSbMHHKCOwfoPj/zRYNmv3mSZVOpA1z2qLjKo3c0vSWo8IfxKmccoqiraThtNzBhlLRe
Yn81pScv7jBTOF9DTnad8HzxClUZl2R8xk6ACQ1qN0InWFukFPd5epC3feUoN5PS5sSqpioxaav3
McObBrgsR4DBuhhmuO99Cb+ymDm49CeMR+K1JvqOAMOT+YeLGKu7kXZtDmpaBtO6FcWAfz/vBa3N
fGWMnIWPN79UCNmQ4pY2uX52Zahnk9e5ignC6p8aDJgCu8euyuocRXu3VavpRGQxT9brb0ECqIm+
/bcxMnCdew9uEmTLBxeuYGAXa+RHl9OhEHF9ZjGyAcau038rtK1iAUP25WOJ/o0OZGnvVhB2q8AN
qmMrbhBTfkUTRmB6FmnqeIAgePYjG9TCVBHfwwhXrksmPtoPZntcMIoXBsXZtee3lpbM5q+1zGZ2
SVfM728PpYGkKKS7+RSU4pzOkxnWnG/3nDwJfie32dNndZvs0jEtUeSjWRniNbCZLlJGNOpni5SI
8R8LTFQo1mcFM3r2UB/RuickpoPxYdVbx77mv441tKOc41G/hRD6dx95wTyIerfLjUyN3tvwxSGW
ijQVCcBc71w6wdx13HcAj4RTe9AaSo7TLftEgtqp6xLsRmCNG56qW6IOcHPXNQ9XeiY0O0mPvu5S
68qsZ87Q+9bqVaKyabOh0z2Xf+iqP2azYzbPSFExVbG5poif0JxmyHWeL75uTG2NNs32dWs62tel
Hq1/xIZ09448a5a6EOQm9NV+RS0EfoMsZPiidZYQRgyas+Wt7JPvN8Dte/VRXY+yT3oS9c9vCrr8
JiHRT+qTZ1seAnhsU8Y+sDqyBw1Eu4IRjOzHyeDmTyC0gXLq7DB85OGKchT/UcgaqvcIjCdW6JsA
qk1wtEOwptua8A8fkPG/2CEx/l5xBk49bTefdP3H5jlcRmy/Io1N6ab4bwDltCJaX32NMhZUrrna
QIVriOykioAndt8a/YpQo75Pr3NVNuGE3iM6tLGIlj952W944h44bY82dLWkaRF5H5Unmur+Ehnh
wQEW0aT//s7LNRJiICsutKmSaJ/QQKN1cSTmfj3274Q2cMLEN8rIZP3fUzR7dyFbDpm5cLvhwB28
DTEX9DXRHXjFS36xSJluVR4D6EwVkIx/h0VT7P3q1aVZ/csw0i1IHvkC3zQvqMkXK8U97mD1SD8p
OHup80gBVP68u0/ox8+9AAygsdYgc6YhZIs1Cs9pIPNiGnhXayJlrDf5r3G3VcEg0ajR7lDzuMWS
4f6J5swEcTD1GDw56diWlLQLyENGKFx/aM/wFSub8M7W7quizCEXXYGnaenHZf/lYknQMOmzSZY4
iDn3Cxx3wOw/jYMvgfp4W7Hd/BkK5/o4udB32i+s2BGBnFgg+el43ap1Us7QUMeQBP/ATXQnwsXI
QIFZ9uv4KrTYmy7jVcVYGDLFUHM5DOkxzQ3+OMWFQEO70ZgrZlFnxjtJVyqDW1Tckph1jz6PiRfK
B3GjZLG9G/yTeXi/2QcTGHOuV0VgpV7sR9cM1jCx6NqzMIxITJU4f4uEERKAnzWnu3qAbM/EXdd2
AYy+lggeg547cZXAST26srFpUcFb+pub5HpX8d5ZdtFJ4I1L0snKbUo1SbQi/rVmfpc5kDy0jhuW
UjlwX7l51En2sxNWIrXndDDXA81xLsqcKHTWJZJvW7EXYJCYFMwg3qOYSCLwusjXmAZH5hCcnujN
prQRIiJFq0L1XobJ0ZBQ7b/GTUCOL34Go8ncCGhOw3cxMVRsySvcji57ywD3yeAl8fBYD652Re/C
RWAd8Nyao6BMETj356Xz/vlzxWp6gdT8m+MmSRfehplp01U/FQxaW/e/Yfu/DAyFKsbQuDD0+/8d
ljeDlGigw9js9zxl0gie85/ro6wAiJR+tTMIKYUcNDN+rP8dFJhgH9qFCNSVQgM10/L8q7FJQHy5
BqBrNQEko2M1870YPzF1pRmCTJhBSnnujeLrej1X2DvMy0HHlaI8a0dlm8lpralIukzRlfl3CRs7
r+kn9c+pM87pJtCKAtDX3ONn/spIiTUdpJIBeXpUFaAhd0ho84FhnUq0nI00Qg81KNWljUEW8Rc+
HA+f1BTAn7AC+ZxzGJCTVFx8QujpQq+UxF81KGoY3ZL7ddKQugH5YYFqL46E/bOThuFp9yHZEqqj
rv+lrO0NNlzL3w3lXW3tm/7kad2DxAALMlufjc9sSBG4cQuWSnlT2SMhQWLJ7Rs6nzjqrKGwYQnL
+FoxKbzgZASbZ6oRS9/PO5epnyfLGydZfahd77h1JKMP7a0b0UDHMDXPCcl1iq1WD1fHe65P2mk+
GJp1qJQc8iFRF0Nq1+63bG3yH347b8u0UjW8w27Tvrm3H1HDbFTtDI1demUMJpEpMFIvJsZObucG
/UQYb5RbcMD7zUxQGdt+wCVgYn/NoG4v+tdDdmm0KBmdl1gEViWktYCwZhOMbUfDSYdpufRskMhp
win6bcVB+mqzy/gyYMP2CtyDm/XqH5cLeCQYN4yo3gMr3K2w9XIqnk2pIRWcIIbaxpY/rd5gR8xn
Ak7qzTq3y/a7YbDiQGUHhMJ0dF9ZPJk60FWYX2EwmizmbYGaFPsSc1vTl3uvQENQklJLIMRzRg04
43WZgRsRhiXf5YPLBeVpWTuEuybS+eclgTtcDQa461Qs+x9wzmx2l7UIMn05GpWWT7r2OPY0IGAl
fhlSS1idPjH/Ux8YhYsjgKPJj4EU0VubbiCCetTjweqqqy4pIH6WZ5Nt0iWJq/qUSG6F58MjPf7l
krLjzHY/YlYgGGrbS0LUeRiVfj6hvFP2K2g8zTQ18oNlgL5yephrYbySDQ7anlxqgWHaFlZFUMbN
cc8Qod25sjwsNqluIU88kXOpuRdroYyKNomyGMBHt998kwz4qdUCW9CrUBeZANngGuizDWKadRVj
0KqtK0q+XKo+LuiBuK8ry6MHUj20h6NKoBDLo2V1pYkwDQFltuf3iFnzaloRHxjkrD6coJt5OuhR
czC+pSPUAiIycQd7AN3CKSkc9QKlVhTUw9DkfM3czI8V9SYDvAduzeZBEfi3P4yJ10sRs3vt+peH
+2CdF8FSUJVTaHtC87ZQU00aa/3jmC5JfjBLvrTDU4JCimSdTPD8jZpOlXvpdK0Ff9/1A0/IOSut
3pPXdHbWFrd/ejxGX67UFsLHH28wu8badAD3zepH7YxB4aOn+pGwv/FgcZhKnkYpteGOqnxkeTjv
rOOgPutUPNgSYBETFkwd6zdPAyA87qEaGbl1y/qR4s1gpEGzEUob5NdJdn+ZghXfdpKvoCTtvdD/
6EAqVpmRdkp+ZGqzctsBbCOrYmJkrDkyRaTEKhddZL23LHQl4TlQl6C7uciai84tS41OpK9RqRbA
rzcB3IkL4dd066AA6cuV2yZdtZRMJJXVgvHe9sunaA04jI+ZRKdYECo+ucv5fbmyfpm9AQ6NQCzI
eWPGRHjOubq5OQKmclJg+294e2PqSlTh33NMboxF8F3NHHejzrvfuhp9bJyD+UcCjbY1JqXhMSTs
qTOG/ischbx0Ne4Lr+bBiGZ4qU00Xh0eDp6R+7HzvPwj2lkzvV5VOzZ444v8THojd+0yH4stgS+N
S+152MY95TPkJ4MjQU7Su3ytXl8Ix5PpaTDjoSHmTGzAmBfA+yvj6fStFp7GHJrbLjMCxXLVMpHZ
nNN9Zj68eyJuRD7E6eplAsYQP7KfFUYPPBPSin+zaUuIeykLT3VEdN/xh6+YtGEpXhJ/i8+raXcM
4ZCvBRLEoTmRbM/H+s5anW8f8ivB3FwjA3OQE6h45VQtVgkVIzJNatz21VNiDwCjQZ+admai2vdb
FjgSvidf/IcznIsDdbF4LLQSMRjMYtXxKdwr9Q9PiZMuJu5VGgZGbQ+w+z9vQN8buuRA2D7t17LU
5wj3bIVt/YT/682t9bV5W646HQvAQXYeqQl6gSQk9hoMOD4gPGKHVqy2INUdgnhWo0dorVr9Mmxo
4vJCqw0gmiSLPcdrB5HQh3DwVLwmRar6ObQQ0wJh85wNo3H42nJHjKTnrZLh9TNPHa4E8CQBJDAR
+yMjXPHlbHaxk6YxOkCxFp3hEDMTZvHTWJyMjo07D1dWH3YX7X1raMlUx4EbI83GIhqeICzlOVCO
vLY7dMP3HTNfRwufExcVFMkilJQUk7peCEh3lwQ1aoc+2bqkdia9vINJMtHXXerM7hKfHFMcAyfB
pUlnK/ciEUNh855dWRHZuJPO5P6oGSgaFQuleQn2rwgzZKYakw3cQNkJm1D/M+NCUaudq2V07wBm
hWZFPwcWFQWFh+/gaXDI3tyVIWvmYQ1q9QwjSRJnLHfWSPeit1Cg5de8BGGCXvXu+ufnVJuuxGny
Q2XVoBWoPMfmUGMsXzBI4RDZHGhPStv4/lpf9DroOYgdR50OlaHABEHtNRaJ20RyJ6jqdlz+KGGj
vPTC4feZESe4fvXwFDg0wysk5cJwrNNUrtWCtt2RXYPMx997j4w80fi3VWp8MrSp3JAD/kGK9CSd
uvVKBkB7HVjoXvZjwMt2IZvM9UcHTitdHUOsicaRmSs/8uSuL3LtIdCZBXESc6W/0mqYU0TjVDQh
e3Y8ZjIjOGw5hm+oKW44FNMaiHUOjfgYkcRFUEuCuY22CcGA9ew8nwHDTDX1iXbTEbZqBdnK0twV
Z5IEL7jEyOBEJFVTpJl9eWB+gp2aXxKNwySFC06/ZopsoGrbnrfsLOwlK08pE8GJ65Oo2BXaGkaZ
RSMy9bfP6fAXCtL6tL3i8bSS50aK8/WU3qKlkzibANbbxz8bEz2dYxd254u1N4qjPy3GJFy/mo9R
9etWnx27DH4C0SLLpuCz6JhrJkODW/U9hqEJeT+u87qkM1PS5ZTjufbfnwQ5iMjaqT/wzDDZk/lx
pVT7k4m2dhsBQb2rS9eTlSRMtecGTVQqMv0pX1TbKy8JR2RncEFTH72QVOSr5vIT5CugUOsSpUF6
XWqUVp28SLdPhTLVIG3JrVzMEcTi+3d7NhdH5dOfbmmOQU3vMq7+ll9qGyt+BW4V1dsTTn8J5c+F
o73Hhzba54yG54ZcW6pcvgC+yFWh7QbbbYESNsxjnrQIPZ58gYHWCBRnBagFlFZw/dBIWyDd4gyd
pjnTkUc6IKkRMTQNOr/Jf2MLhZg4mj/IBoTWf/ACZJb/xVNE4Z5S4oInibdAo14kPRFwYBTAcoYT
fNb7EO8xZgzKjgKEuUVWY4G00kzJT/aah48K7VSuCD+p4sWEhEl3ZmasY7doEW/q997aA2CDGAuf
aWlv3aHyFHtYBFtsjrvixb68vLNsFgmFFRMKhy2x/r/giYf6NFHprGHDOlZU8OnyKsZLCtVflUJE
ukNdWsYaOg6cBYF1MY6xSxNCCOXeM5270+YP/ZVoC+nkcIEKzPrnPxY2Q/NZgB/zd8Isn5S4jjVI
AGs9DCB3kYbqGynhALXkL+WJyagjj7chwQW0T2tXy/J41097m5eLXzDhpYltKPDCjE6r1oV1iNRz
bgyLaVrKbliljSEz0xcDmTZXSFED1kCnZusxwb4xb1MFtJJbrYKBgKdCxkcm0ymrZOTUO9eqbnIN
5NjI9iNDoI4dEolS2By++j/gfj2b27fyNV+VNd3WEUUaoOz1MExe2Q51wXdQTwx3ErBEmv7hovR0
DDzn++ahtlakJjCDe8FEFE8200S9acSGxNEKCawstjm2JzOkd49lM+6k3tubYYT7lZB4iPmgqAmB
X/u9DEBKeMndXKKjVEMb6L1wCsNQXfrHGTDOgZkDno+uC2z18a3q5rK2VSeJ8EVvOSRP2kYZBZSu
lveGr/0OQu/I/0I5VLzGBALk31V7aTvG3Iwpe1qSR0QNFQ6qkfEfL9GZtqbYgL/qLtT6ERxH3LMJ
B/JsYhzgRuXMGcuEQm381sTg3MeJK4HppK8BI2iZz98oOnzm3dnCmD4dNR6BXxn9dS1YuLwGrWCd
xHUSQOL7MN22RiM5hRUCovtWQZ2k7K/6M+LJytLUKnQeYTYwzsSA/QN112WbbtLQT+fMixsKAzhh
xuOHD3tFmxC7XAfl+oyQEOe+hni4qLHxUWPeqxxjEEWtDPKqJUFQ9V8ncKff44pmZf4OlnBKQy/n
MDvmNJF19OXjYKaThdk7JwqeVrD28kL015KuffFU+isy7OzqNnvINw+zpKvaI80gg4UIq5MeWly0
tojfwrwAGgahphi1o8gUAtppX7Gf2V17Y2lOKFRGnrTnf3DjZ1gbHfD49TBW6FRvtW2bSlSWVBGm
HL7nvRKD7R7DQgTuJnB9Q/64VBApIki1AQpRch2YIAT9EgSUZWN9xeCFmlsruh3HiyjLi6YXue7h
JeihBBApvtMJaxvofBbeaml0/jhA0swLbZTY8evfX+NHRzX2ipV0ZbrSqeUPgUXz3A1NA2bzDoL1
L3klYgvp6W0CFy5VHuxzxuZkrkOMFNkLd2MSJKL4PRITRAtdJuCVVhIvZgrHFlRkepDKeDVUd0Cu
Yn7VWMXBlswnIh5/JGKW7yDhdeG5CqD86m+4BEJA/OQPtPHPSav2I5K6CPFL9zh/GZPBhEwiYjTM
lKczx2qV1gsPrUrsx4lskS7lPeit4aaqwS0m6hek76BHWdn4I1alc0P7w7nY40xq4abnDoMw0ODS
6xA704H/NhqqkjvfQCt6InEjsJh9/WqHJ12oT8ouXdwohHOfsUfLdg8OkfxTV3cyAa4HZDjw6FO5
h/Nt/s4gbz5kbAYZ1CI8eQ7p8htB6xcpZuR84YXqcZ+iDyKV9cs17q4jpLSvZxpqWpiyzFY55Yp4
e5P1V09Ie0ufuObdeKPDx+phQz57vFiS1Yp0NtJEymik1ti5kdj9ye1Ho9wnaehX8jjQrLiAs8Wy
JkX0NmAAG9afpggoZ8Xw1Z1cuNS8DfDYXYwT20KDqk9/tRsxZogqRhCrD6LHll2wGbAIo7FWvbBi
uLvi+Mt8pUZhWwJmpW/Nc7i8IKxhWy1TLcMhU5D4//0pW0q2JqQH/XGSs488pQXCTRinQi5UpIeL
X0DMVxuFlkv5767PqlgZ99Vxw7KmHevTAmwk8c9v6N7ge05N0wRsatyyWvHiMPemz6EFooy9SE3d
lXbI5RUItmTusPG2lSS2HaBf7yYn0gLNkwj4MjilY9oJKiCSxcRjMCPFYetdGjXy+UpAaT89NVXB
uE3RUKQfQvmDOS4G5eVnwc3WrnNrmb0FAi0XIdvYGnUGaMizmqS8+jEY7jChMoy3jFb8TiT4Lqv6
fzwxyKNl8ccUXPmdlfDP5kPTty0l5qFiI/YD8KdDEbS2C9SJvohg/WT0nLg4ur80aGlUutFboCek
/k9VVDJ94nNa4N/betUmcQoYx4K6sab2fKd+LYIQN/OkdCtaf5G+xQUs+RPVpyXz6G16UdTUBnCD
8oK/+phG5TUsKesY8Ai9Se1rhjHQpgUY8VnXJFc0pxj6ZrKoLs3fdiL1dbnJ70b5kWq3OATL+8Yv
WtmW35O60SH6PPav6FoAomYgdlTBitKlOjbQWdseXzb3cG8/FSnil155E4Ux5T8uXQdjeKaBk5Rs
cn4u1qMr3+UpF3w05eXHCLiQDCKR9anoaT4vgIbEmmJuwG2ks9CvMbn09AWX/yR3nh9CNi7Hys2P
Apk6t4IkWOcFQN+KIE81/Fu5P18C4Ez6GQqoWvmQ7WDzxlkb0lJ6T52UogOiC0TtbSkjyg7dfJlp
Ol8YuMd7e5uO9I7h17Ym/12ukF8nc+Hjw/mWxxOLNHKixkudtmSUDFCHzM9nknwS49dcXI9Qd6qO
f6lFOhUrGixmfYDjyRiB5RlwUYQFFIRTdRRveashdGFKKlKDj7JdZOi6lN9eQY9qLMYyxpFlYXZF
OziOvbtP/J6tOFgDqts/djBucs5xJx18FBQkCKTCGG9nB2spz3xyg7So407KNd1kjQyQvP/s4yEQ
b4qp56kT0YDsR1ypluhtOXXfSFrIZjweskcNF4xwo+ULxHOqqjrdiOuvZX1lfgakN0CuXbV4x6kB
/zGqT9LlfCha8DjgprofXFmVRu8K3wlzbTen8dJH3LWIxp2MYeZSELi2c0pBB6SRQfU+8DVqOAJ3
E1mbSEidxXMafe57uRN+bQhCG/vfv4qPOHD9+Isor+VKzByVWAS6Nvxy04ub5fuS4qu6HdfLE+zs
e1SUGKDFxVgokfMkx2srlWnCc4rixZoqoVFK9sxtrhF204oGnEEgk0OZM+mVOgBpC32YDq68zF8V
pR6rmdz+qhShf+DA9CZRyKdtcCgld7HvhlgxhaohxR1nDjjwD0CoeODhPUMGbP2YrUGIKBoJYIBi
OKdEtJ5P/n2xnBaiPlromXZIubg6BAn6v+HRGG0y0VaMhgmTCILRQBoidO5hl0dMCZqCkSdFkeZT
jeB07YJ7MLOonzkohNxYJxN29DNsC6Ob3d1AmnbDTW9mLamILX97tKEP4/uzgGC6+5zdUpCqKlU/
uB/QyUwy3z1onOLqTYys4BDvL4YWQqB2suCxpTQKynMrVTp0v3Q2usblXwUOM5xUEK3S6Y51h3Ss
aRak14RXkUSI1F6Bxl5EsoF5TBXcLKcwMOabL+EICtZ+yDgnki+hXEe6xVS6lQUh/EqzpIMkbkfs
0G8eXoanxJpx94x7MZr9+gPELmUyPX/FSHASEELeuBruW/9P+uUm0rcLCbg4E/S6X3aQ6PBy9eAo
zQLq0HfVN0KoTiUowvzUE8dkCbHi6sP+HQXZMrd8P9rKULTXlRl3U5yuRvDJzdaZI+n7ZQXWebNL
W68iUzukfIyafzIJZVw3H0BErs5SoDnmDkdFrdzD+59yqxKVNeACygCOvF9eHFDej4ZqupLt5uYU
Tyn9BuvwY+8G5JY0VCd5MUiOwMjQrfbhoPMbZghPPg4u+Kr6Eshi7Egn6RKu8n3xLyx6Hb/AmbH7
a8ECfYV9mTFh/E5MxyfjiUfyxkWfThW55MxNXNCpSJ0PmKJywEOrPG6sv+AVUFY56DkgU7e73RL7
Cnyps6MzVPoE37PeYFxdF9hWSKhF0pemrmzlRO/k6Tb152Co8fBmo/7TWvCzqvLpwvGwe6YIKUAI
RzNdutjuTqyL3uw1PGLdlZDUtb0MwlP8Nv/wXnC+wrI2D6+0/cJJ5aVPDrab9yp1x7phUwEv0qyD
HzateB6RMb66EPT/hW2p+h6pXUbaeTORjllO42jhOoKQeQN9tN/Sc3PQrwyI/trBw4P+dwxwcWMJ
CPB5JBv9LlN0owNIRfsq6wLxB9YLEdy0T6aE2SuGaCTzdkPGmqQaR9dOdIifEWUrJVxMGnvqtKzG
L4ThlMwMryeHe7F2wQHwV1EKovZXzu86gOjPL4oYsMH5gaSXjCInBDSakhuRO4wuRYPTyRw155ni
XK8YiZvVmfebn6FO303u5EAmgj5RHdKckTklPT0JRaGFW0kEE5m1isSWYAsfxao+UalbaqjBlgww
TQrOo5XQSPLG/fZi+tVhsyqMrIsggQckN+xg+qGTVNPiQfFcb+Q5IPW2cO84e1uhF8V+iif6uDj3
A0IeMjZWzmX+jhcMiAfqI65cFgaIKbB7yA9KAKDYIm670kp6PXy+IHbQTtVqeOq03OAVB6SsNL6+
IDuEfI8gVZYKEgydUVLQwHTXxbPGdhZssFLBOHUXUbqrfyqaHzLDO6dpqqKMJSzStxzNxwiBT+b/
XnCvfsm8oBTWqsMC1kFHWZBcgfLebG4VXShxxLcWHpTqHBzH5qMRCQe2T6M9w99kiA3+LCiCnxs8
8Oy1NqIzKK17wpFy9ok4+/071aLRVhK06lMVUo9b0LaLtWL1we0IsObNUtkjLXRIxludozFAZd57
RztnhDGUlgO+NyZ80uoZ2vPhSRD7fFb0AJyTbBo5ImtVTQTZf1vUr57LcactZSIDlQDM6R3ajFKd
X4g/JSvqt7RXQxDCh5l/NHp1VlBLlgRJxMJFhenRXyJsPua4npFay1Hdo9KDUepTmTdYPSPXKacW
L2cb0rNZTz79mI+ET6VgNd6T3J+C9CCIzk3um1k6j6O+53GSgao32e966v99OmUOM/9lHhPG9cZw
m6oM/VL8k/n2KajUp1WkWsdXJTCrNzmsnCKW76LUkCY2eD11hKLlo5+OfShsqZak969+7TlGiTWw
cqpv3TZIj/qgX1msOx8m4ISZ4AYWSm8AZtAxdLDtCDTGH5Jiq0Ie7frQNcjzPXowg5rFlFkM/qHg
Z/s3gbD4PCqbqG5vpGHICZiknu82TQelO2l4k6H731LA0WTHUEnaQRKD13j3e8P/I72E+JA2JCxN
xQI6br1K2I6uGPcOq+N/U6X9x8el8PRCUTO14KcjEt/gBMiSzpg/1l81zoywG55/vWmQnro/nvUs
VZ5MilnpSE54rzqTDteIy6RWDC42jh32ELz6lZ03w2O/n8bO6ynSGvEtdzOuEq8B8AOJlHeoS8kY
S1czfIdxiPDXFmB9i8xVRTWgppCzHEKVISnLDZbBm7bwOY6ohCoRVRbzgGNbCbhyMt7ZsPZkER4t
2ziDP2xRLdCpqasoyEkezJDSFoUNMb91tWdjkS2EpqFf7DMl/0M98egRxMfJ2U8DxDJzJp9k4RqQ
PigrkldNGCS7cVn0QOjYzxe7s/bCQQL71dVCLiDRhPUvFYIUi/A9Fu595F8AwPNk3IoO3xumsUDF
odJykc3LnyzZpRqLaDSE7Y8Vwc2yRVgSOGYFbVF0F53fCUbb7V/VtJC7sLCgFyFT3NLxSAicPF0O
hEipZNQnNswY/iywbq5/Xle9kJo1sYTIdmzLp+/jH0hH9qU+4+ISOh7bprtIDi5if7sfXhv41ixA
knb04zazG8sc1dbZdXg4G8E9poxqrzAYFRXHSdHSzbgX50nxDoJNLQlvNyH4rsNWzvVUe7V7eHPw
RNketP0RU8ae7f/NuV9RNel8HZPbRrTwxSRXm1J9t+TYq+YDtNubE9gHMpZSKa8i+Pzo+abybxjf
e8YuJ17YOOMwfOwEQeN+mTCcBhBsUippKIKyikc++IJW3lxD9UZSxIT+5XOUv3QCzzyuovrayhBj
2CNcXhdJXTsM4T1DF0ZMrLUncTGpJd/nlroJhVmaon0ugqy1pB016HDi6UaVjy9AfhCjf01ZZsRe
owaRV7IPePAX0kPdv3E8S4cOIwp+7csy9q1/KN1qMd1n7ABEJX5ljbzRRLYiYQb42nklbaAE1eHU
6dMiNfHm2Wvm854Guik5fOt4hzdEXMJOGIY9cu2Uenn3rAvtF94I0YYML+ExcyXrkdo3c7OiMSKE
4J3qf1r2x2Vb+TUV380hw1lgf4uiTcjOfqw+rFTXqh7VYfL3x+9UcHj32AhKy/fWdwI5wLI3VrYm
wafoWB1UBBcLiIt8u9c6mC2VifKHPyy7BFZTRj4OoNUkkvhesatKNdsQr/EzyWcHCihsgtiGwFY7
9cIbXbI6WIJywkUdakyy3aZg2YK8+m8h33zu0e4HYVkXB4vwOw/JRUifg0IAXZmU5g1amfZj5lun
fyDNETS5e63GKLujSmf3e4abfR4cC8FXuzcxhmiOvFW2n9NrJt3pmD2FkxbWryCQHIVCqZzeYSW8
Bxecu6kZiCfRFhiPFKLiwuyYH2QVOx8OJcLOM74tG9oMFmRJXyqJHPOmK5Bd1/gA+31n72GTsgXY
u7ZxInC+DvdvLGZaWJzLo0RscKITW1zlXs9nMNw5EbXEANdu7PlSj+3QEyp6xsCMbNIxweqvRe1s
ao/xsFSPTpy0Cj3eS/syXheHLwtB0d5ncj08Q7Px0xA2Uo1oWPRF6YNliSJ0kWrqNLUJsmEX92HC
E1fn4oKJnPSxe9DrH374IhQsyrhNSRnucLr8Wx9OmRc8ua78VLXK/lN3Lx1kUbLtsdqWW7Wrggf+
YQcq0nk6vBEuTxKftPeg/hXx/PZqgQ8Au7IUjjPYFXInJ1qfkFlpHiIodQSys9GFfRMPcaYdT81b
zkzWGeWQwsSyA8TBYTfscE/34ouy/71rZ9I2HgP3PAE/65aP8rn3/RWvDeFASKrryedi2HcRZ3tp
db0FvWai0BEk3KQq5O+AxGDf9TefYIqD3QmnAMTrk2sxECrxFarw2uBmZ3HznupHAuHahLuXBILV
x/K9lBYHMY0u1nuTWUkgRlFJWxLJjMlAXlHpv3aluNPuo0rL6r2V27Y9JFZZHqbVhfQ+VFOcjDVZ
uC/TZac8PPqqK6l4W43DiMFEI4iT7l+SJJOs6WdqKXa2nrBZKuJUmRRumnpbET491Xk+ImzJunuP
5Ckouxi9Ykr1NUmn5vhR45hMOOzAcB4AIFqp4rYcbjUCYoAfqSLRHR1ISBY24xXJw0OiSSTHnvyL
D37zVd5Yqv7uYaOUkLQBIvDS8pomOxqqYQeNI0KjzKGYTyt2YD1mkcEenW/20mPOj+33vwNPhkIY
1/nV+M2Ou1iGb0eYV+skQgD0y7ipF8qR46rOV0KZMIIdbkT8e9IY/UHWfvjE5N9YT9T9/dPx08nU
ImB3wTdTUNtYRf4e0Eog5FuX3qMpp0IOvyjnNhRkFeHnx5ob9cCIp+qNFP9mxpqt90Ju8sZvA1eg
wEMstwQ6wMNj4Y/zJ6r9OFiabXoQw9eG7vg6uNaIurnTGh1wtrdBA12KDS5Gw5Iqt5YUIQuZM7xD
EUfYhwSikRl+xwUP9a6FG2vFO4ar0hzSYGF5kqXa8cFP17+ILupMfxrpJyowUq+vMvx+f+TOW8SF
21b4yzVKjpFHIH8/HGmUmts+IsGAnhKuyzbeuXtE5Y1gzifWY/nGAjAypGSFFHZVUHVCxwRGDK6x
2Z2S9hgYO3iIHfrouLXhJJBQv62/rExnHikKOyaoXheIlpwvCVKY+j8f1ThtNVCbvxaCF8OkM4TT
VFxv5AjRR4cNHnESjVNjWrLXNCUE1a2CgqJJZrBhOYhZl6442fV5nwaKeBl7f2Lf+mtZrqZTYL1C
yqHvhaNKEnjcD+8R0YvQ9wEa+HzWJq/3aflhgmdAamplPo+XTh7vqwgE9PSGgn9nUNeCazqI2qHl
9ylyIBT3YcYIfcjRE7ZihFbvGiwo6Q5wcN5WOLBUdbm0pvwlmuKuAGPKi+RgFwFO2i7TkLPR5Wo4
EYFyBxaV6OgGCGm+JHBX+/RGMNcGBrvPFwMKoKBxpuaMC7TLnNV/t+ZsPdpyeRUDouuC1PP2fFhl
Jn/uOuMrvinCLUXhC06Djic9822kjWc8Cl/3OCirmXDr7MAJWgP9BOoKNdY6dq3cVSHo3JT77t39
uTBoeRmDK0MduJVwKW+O/TKhPacHSFlFBCcl/V9Wfnat+kMu2MbLoiVxMNlrP5p/sRUXt1dqv8/H
cKjE+AbrzhQmMpTc3IERKUq75cai6435Sk76rwuNcIzsyh6dw3yozlRy/JHD7tvniAxGQAgq0X9t
kc0ZP2sCidswOtkihOD0EdkNAM2RppR6aZ9hyKZgv+ei/FILlbW+wqZPVsps+LpZOPpGO2i24pOx
qJbUhjGO2CPg96iW1DkMlpU9Da9Sg3yvvYp1NccQ/3rGjGhpptFni5jy3AkZZEaEstFS/fBXP5uI
gNrwtr4R2TVwscZh7d8AAZjIo1YRGTLZyd0f4RQXvWAch608wnm6p6KbkzP3N0bX3/503bm5FUNC
h44vZn/L5NDQEUTImESWuxM0uQBkRGo6SvsdpMpXDwpD7Z4jwmphDViy2Acgxy0vrz7CM3rLWfQr
c5Dqa3SIbJyUN2qnMU8+hnCm9lShhcqFf0fUhCUuC0Y2+vFGzjV1kSHGvpcg8PTUh73rcG0sK1CW
7Q54iqrGECDbVa2G/PxmCvk8MQ9BctWCjJU4XmqmdjkT0zUR2WbAN/Ldp+8Z8KpvOEWXCQvVcpqk
X5rAzpQKG2W828NV2vaAvvX34OaMadeb715mUFuCvv6LW14XhicJhJWJ8xJXelR2+AvYjLymkEfu
aAStF5iKDkej2VFB72uEhe9ruCnFVRpbFqbmRxM6BTyAOejxRZIxWLf2IhdUf+z8g1nIujX6Tf8W
7qRHbn9+Dr4bvEy8AgPkKAy678MVJWelPT0gF8+0BE8EyieBRQ4HdhGv+WRPk0zI6fvtPRsyGckC
lZJtiW636fsUjoE4TT7556i7e2wE17jsbvnmwA7fTRRxrU+2gYzRmfvxRhntUhCsD+2oAiJYD1RO
Pp08T5TVfWBS629chbbUuSoGRe0bug+1BOwjU+LEBgy9rj9X796uAV5hD6oD6mgppME8i7tsLQCp
/9Ciu6+XF5DTbAYHZaAXPmT5DjNt63sFqJ2iLFF/DZWBycM3dUcH1/V5MX5a3gIVpR3ayKIKLUwl
mw9hEKLU1VvkQB8bQu1WNxpWbWExiVRHXPGSZfLHepgiU6TYv7gpi5Aly/w3qlikZ9m5F+4vZCAQ
Hf6HzUG2HjZvEkpLMtzyoFYZig4oZDR+OvOQGk7z5+G8BvyffpjBtuEfkeM8LSLJ703TxRfjVaDl
R/FKW6I7ywuSowxnBRlGwuqEmt3pQ7wgb+TJjLQi1WEKmMS+tIVpf/dRb1gK6mx0n1IcdQVeN/KX
vuOmRxij1Q+Vx43L4ruypqq9fGPETRmukTNp8glZEgp/d9cpIf6aNGPUXxIHNp8yckVcZsB2uZwj
nhPeMvIdhceC5/peM99PvKrZcRVihTl+2dlYlRCswk3gWeXhezrgtfUm9nsss6wkEneHNvS5m7QC
YiDZTh0rnbd+KTjp+IUjj8rpGBPC8hk+MNIov0L0p/mrJFUrblzFAXA3UQaWbMB2v6FmTJyjMP3z
lkKmKEYopNBosl5g+bSCPDimuUZECF6aEtFI/M+PL2JM03EK/m7JrIOwB08AQcCcCt1igSUed1Y0
RS4BJBOgM1yChZpN7aVhPFvoR5Me0XHA9vsA9e5mdbwIKF6RjWgcPi6z5jWPEELGDWJ/6P7VLFOT
V4Y2J233LqqR9w+8RYb/TkDBGtY/8Vw4+hHLA2n+hS67D4Xdq95CuOKbiZQSJNd5sA/1i6/nGaRJ
auwXUw4zXkrF4T3+DK4uVWyAVLH+IyLzkwMilzMPajNY+odrCi6qSvkriPt56Qpxu6Oh+V4zQ5Oh
4n1Qy6ZAlrTJo4SaK3ij7/lFq8voPZY3je29YL8+S8qofoM4mxQHA4bY6TNCQIy/phJaPlZKLoeV
avp8aVxs8AUgo4Do6btmDCFofheKtBRBR4/mNsnqyVdJOIePv0VzOQ3NJauT3ryXtoADdhH55Dou
Uq2djhyJE81B+Kt4NujTFRWMENK+CYyi7PNDXCsDEoRsQu4gpKvqigPTpLbf/85XtxR+lyhR3pyx
c1WQyijvNPnSLt+zxZazC1vpvQwHY32XyikAgGLaanhzD052MxgvmvGrPqjeHTa0lnj7pZrY9mbA
aPXW1w5W1JpthAzNDyHRjQY+n+v5DPR/YJ3bjNHxYS2cOh+QRYf6GuwknfB0LvpT5gyx4jYtNMeX
Zed+PCOPALVQMp1wqRLcZgxKURooQKUWv6HjxuTscyTNt6cqIwIRWibxz3qCJoXHHHFTLH+ILmI3
O7/B5NmOQUHW+vffYgqmBvSjGbdotHQHNFhPW0zwh1IjtVcmmF1mCdufQdu3Z9tqe5egKtZhYY7y
gypfQv0E3wLNadHJXV0zsGTS1WFxP3lw0VFouP2HmSkXpzLJRqPT98pT2zIEVtHYyYQKzlbyiD5M
P1kVmEB4uapr151aLYn5oPzhS2p7Jqv9T0qfz2WJEQmdQdAdY6QmEzmkr1biXCTY764EF4Lhvby4
i8zoAtW0vzmF2vmp0Dlk91hyH2URUEY6BPKRWemZfldJojB+BEPsz8/x4Cb5r3Agkv5XeOiI07lj
3LYw+OfEXuxhmHiuogUVKhpPTQl1zhgi9BSckLNvAtdTH6XCD2bQHUrOfZEZipWPmMrfC8DBLHRI
WwexfisPDPwUMJfHnbyqnVxWpRCBYefyHyw4Zdq+K5P+oZ9s2Z0b+eIbIRoh3j7tf4+bNgY0WfAQ
wb8euVPWYnpwNbrI6FT1LR35ui40G4qgKZU0/nXMoL0Xzemeu9+8doUyGds2FrS5w2W/zZi+VacF
9C69LG4bpcphR3/tkB8OSitfYVFNRzFX6Kajjk6Sm0o5f+IFhdaE5vg/5tOx5q33q2ZLQ7DxOMkD
IM+1cOz+F1pWEcPNLofpW0YI5+Dyr18jzjC6wx3OHCJHXPRtvJ7yyWy2ec6x/9wOS0e0O9+OPtW2
CdeWSr7oS/CP138obKfcJj05ilr3ps4bJdsaGFIAxyhM4XOonhi5Duen8lEJHEAeklOJo4QD35gh
IIS8nwQ62xchKzDJTMIph9ecsooL/nx4x4hwwS8IK6O89EjB4YbDzp6sH2Pp2iwwk9uC8SihiI6D
pRUwCjxZNc7egWoZzENY/4bY7050p/S0+8FhrxGB7CPyHcHL396InKMn4I4IL/4B5FNhZAbvL4k2
H1+ABAFwl/4HmKMQ81NO7GrGUY6MTDp+/1ocSNxyNUnY9L3s3/ZCgJugips4wbMDcUMJbfY6AOX4
YxWdRzdMvhXaa7REYrpqK/n0DEl/W/Y5qZE2subV9MsZ8D5kW6LHf79oaMuBYMLuWoRdOgN5tu0T
IBg2g1Uw+5yrnBXa1HhNwPqfq+0ufgxdxwL7m2ojuWa62cCw2kzw5/dklul1ZX8N3TCH8OZoMo4b
cbFKh6Ie5ajks31OHLJ3b9pVRi2N1G8uPQoC3ZYhxIklxKgehjpf3DPDD7+rIVtUvyOrntzjttlM
SxUee2xzItRlstEoHiTHeeK5qHTxaKRnxNy/NxSoj7TOXQuThJ191oztVvw9+XssnVmHaiqt/ebJ
Le3U7Izeb9LjToBr3mqpGvhtH20QdZ4ROmxfIYwZ7OyvBoE/iueXnmWqlIVUl23cR+c9LofHVgCM
GBKR7izWftubwaOLviSObCq5cMUAvUD+z1jHv6wauer3dXpIgB/uZr1QbPLac2HL8mkU+HrmNlRn
0IV5gv3eblB0XmOfXchOWNgcCk8iLue4VF4ha/umPqlvsSw/Kxl2PlIc6P+/XSW2Y21SYl7RBcCc
+ZJ6TmUacoGXMOc7QTMIKiOjwnr9ZmtIQXn+HxWRL69XWsYjKM2wSzUt5uJ5r7df9AXqEWoLxhFl
MxfQ8UFCctpowqeq/a+riFqvljCQEjiKBsoeEW68CIXSfolYPNjtM40Dh1YRdIfPkJYXkfzRSd+a
zfqLxS9zYuciFDoDxfqCIzAM739ccOMTqt+21AWjn2KV90lC6UrA/07RhIEmMRrwEOXOzaRWOaXj
6LtHAV2TGX4697/TXO6sluVnRuVSgivjT6+38iIUKa5gk+KnoyUOjPvTQPKx8Ku8hAaER52PgwQF
4PN2gaPtxIal2/872EAyJvl3Nzp27JlQ2tawLFLI93so/kN6Zh3x87Z55GJ7ar/+3qPzfnkDOeKc
3R6p3tListPs7eLKqqmTdJkRBZPLcB5uGVc7nBOQnJVpaxLs3oE6aJppdCosY9gQ3j/XjUf1N4OO
eQn0dGYkT3+MeRh7j9IqZGu93oQw53gqW54v9GX9pTsnyHGlF/k/sWntsHNm68IqAJl/doYl4vIA
WFANiHR3RJq3h1UHFy4h+cRoMsHd9rQqywnvXvgt1jNDtvyFMHmswSJAlXXpd03HGxGYEpuBjRyG
6GN5Oy3psMFWfknAD19vKH532cANuNPEUm7+WRgJX3UoecpnNvuxRjJLhH6Sstrj7yWZgvm7y3nf
a5lAOTZJ3+ROuDNW3WFOuO6Z4Ww3X6dB/dZlzuebVW5Deppefzacmug1e+XtcmQHqYNlh0vPXTn0
e+A3L2DW3lHRZr6inSg5PSFrGU5GLjj1JwTk+a/9JAv9lpBrKw9aG6qRbvFpAKFMhOiEqR+PjJwZ
vpJNb7s911ee5HpM5xyZ8QiCKAbZyv//TKGULg9drdMKRQep5cFqQtcYMtXYwsboDA0liEiikp1+
kVc6hPOZLywHdn5BNTTsLqr1GQiwRwh7YcAJKZWRFCbGbpsJOEIWjeMCRy7uQ3x1lbjtAfY2EzeT
df39Js6oLzoOS3eWDV9CuumoQEqHfLuTk0VeN+0YaJzZ0KzYhGFTMGqiMpaibegjVXykpKY10ljE
4naXzFVsyuctYGhpinBTf/2NR5gFQTWPr72VDJaYd8NKOWujq7WbbognE7dg3D2n/nhdWo8p479W
Mo3nYlFz1QF2diPjHOF+v0LhrAiAJCVMmM3eDrvipZ26Di/eiu7Fgrs+a+CDFBNRbHrpBCKOmRaB
MbDaUwfl010G01ixR8vCl7g29F9S97EUP/+z7PUINg90vXqvwYCyiLDNcek53awDceO7eLEjZCs0
z+45OPQnhD61OcZYkeCu/OGQw/rEgCK8MCrzC+zf+AdcTGG+Sw7CTnRux2w6t1zJS0MhN0cs+xkJ
7+jF/R/HSd1m3TgLhJQnr0jQxx/fX3VJDemKAEZBV8/5CtuxdH9chSw3r5+Ta/0Xzx+XX3EwVOyK
fBpB5vylqXWyFq1Knn6pnzwWM91FIcnI2c4QGyq49Osch8vKn5+AhWWChLJFEMRltcqA3d9HhCUs
2nHixi8U4ZAsaq/RspUq7rHiWHY7y9FYP2zZ0pEmMCb5ypDO3hL+xSb8TW6dXdD6IpL+HaI7zUQM
YfXu58Uz8AV5AgTL4Vw4SJaPz1vFzpN6hZA0PXX6VSmUGi+61EFzIxjk/0dw3uR4iy0gNiCVIZlU
aVTE+vkvtyyrUaJvvd1qJiM3Xk3fj81/ThXcBRVDXQZvER3l+ULO/9ARnAPnSQ1WK4GEqa7qmPIn
wn2attITRhKvUhrqdrpiMgaTVu8N6m3h/+YAyT5wX+nvZrdVg7eWpT3V73+Pk+Q9i2D10W0a9AM4
xs01JQph4ud8hXg2r4RvUH6a3BezVlhuHOK9hthtJKcX4GFxDEE6+pGxAsHVOF6IwOBnIMVyc5FH
4LmbbPbxY+nugGVTrgVPDBZLDPf8ItDdZO6t6MP2rRwxD8L/9GsGazu0MoepknrW20xYiD4FNRcM
bVa1f+F/rpBlbYnanzVWZKoQhUsexuiyVLz5GPXMEFN9j/FoLbbgdGdboDl18Qsj8mdQJmf5r/3x
7n9U1ustAk5dpQB1+7UH7x7lJNbBXtN6yag5xyGiMi4/rPal+PJvt386PrVWGeFklOpiC/94+tnw
BPWyGytO8tuyHVIrGLL03ExA53cX0BAMvY8TEGDcHpsyv1LQCoIa8iCDdAhZWnGjh6WDS7Jrk6vi
cXkZGkYD9oDBicH7mtOCf1gdCkbTlJveGwUjVp/K9ZEGGxXuf4ul8sTCel+SU7532TDbgR5L/SKa
lUnqcfsjJhaP4Pvy7QmetfoPJZkyB13lFirYIabAW96HTreI9O2Qjc4kvse099GYn8Mmn07RNW+J
u5FmQ9AVyAWdQREfVB9nY/B+hkPx83n3mI1IBtRqoSjPIaLIHDQKEOyE3dYCmbG+ICOdZevqkLRA
+iVY1b+bwX67a4ch8abkRGajxzUefNfxfIBOUBKOA/2lrSXUX6nZEJ/GNguuoDTII1TyjnyidoI5
FjzT4ZFxTcinpdEx4VaUwmIL+pcRgLRgS8CHiH9tJfSgiWi1TS3J9qhLclH8QTw+ojAVReOUEQ3D
B1Pgo1b9081ThtU6U77exzG7Ap7C3nfQP/Byf2orqeli/B+2DolkQbRskzXIdZQUBDJ/SH4v6XeW
ac4my9TaZF0cpC3wM3xIR6NIxKxdt++yGjTHpo5qGKQebV4/6ktwLuAz8PdPZpXTFdAUbwl75LB2
g8dZ+GX67mbIQGOyMx8h4usy28MAWX70nmwBjy03gp5OGQckpCFftgx7Jll2MYTouUACr6XvHifg
3l4p8afAPV0qY6gwQHmd2IHsLwnytZko5zYRytzXrcBQYqTB/q6Rjso2X8y4ViTorNRdWvuGUznr
4qcu8owQtBpsmawO9HfikPfSZwA4zr8Lee7l071dDgDHy6qpqs5KRDGeV3bFy5JxFbfma85g9fHh
3s0jNece9OHKHXQlIcaNZlA7y22kw2W7P2u9+sk1rD7iNCKeHSTndGT5xrDB3h3F6p5VpxjItfiB
w84pD/f+yEMxy0WaTJpr8JD8CcLIIRmuRG/hdmw72lUU3cbLCvaBMw4vfSW02Lf0RR575o11AeCk
+Dyh9EeI4eUPcHhK9GyeVZum77nKBCB9wLRsvkiWl39xq62tSXg4eoN4AANDOhOcPt3kPSyLQ8PS
cptBaj9m1G+XXHlnqKsxsFmwXb34IT4qho8y0/AYFc4V20JsatZqGV9ApgAH3/F/0mhTTFBQ7jXH
PO7OZ65hdmJVP/zcBHCgqvF5bQgfcFWW+vkX4u3FVwXpFdTXJanHgB62C5K/D5LXkMcPjYCidBNE
ONGSiIaA0DekOhh2GlxgE6fU68e9on4u1JJZUoJK5S/U5m2oDNxneq/whXIIFO6rZ05ZF6V8U2tC
j6pdn+bIJkN1x3qwusyRV4E8K12tPztYUYQpZcpskLW03xV+cBs3h4WOVxaklJ41GzLwlbFNM8HE
k2mbUCG1/k4VNEDrNFF+WyYmmg4Itj1AwhCLcSISqdh9s/hOhDJA1UEZJN9LHejimp9rLu7usSsd
hISvn7Lpux+Q/ktzDQ8y72T1IYe7ZJ2XSGCZSMPYONkRLqaP89n+MknNZSX2ZpG/S5AsKHqhw49y
kWfE3tlwiJnfScg/WCgVoVvlS7AoaNbDcLKjFF745d5i8NHAd6U01l9g1C/jsuTjiX+E6hvyXMTV
uyUDJiqjGhwGCgWADWEPcxeCl2BbU28rs7ExDJxbpAZKydXMWnjp2x/JlPX7BeodTa1GgSbippaI
ZeyO/bMqwyqyM79vNQsuI7U5spPEkcZNkg4UMw5PsPtLpviAAjf7adMHGp5G687tGch0D1f26BQD
TXdhPaRQKI1L3uS/86aNCggoeC6YZlptm8MW2hap+hhcFlOKVlH3nYYASsckyKh7IJXns3nQLcSn
QbIa4s4Cg8GCMsMMgyFykGJAgFgKnYR1o52w3VaMvbFaHf1Ee2s0yVYSBqT/X0iEW53tHwxWwcC9
h/dfq4noXy9duwDq86rk9WL+UeW9Zhfa8Oo6R3GqXgTMxmHNCT3cDs4qcVUcdptoZxYd1GLNd8hn
7CgWvYVzTtnf9irpiNNj/rBFAdHa6maH6eJbC89QA6HAbckN/Ol0sp+fl4+OgrpaAfeI8gfmMZmv
if2GHYFptHmsytg/fpizV0Ol3rmHGLHdOLrlfb6YOu1aMyUO8y44YU0/0GfFhyFtWoDuRcrIReNE
UbkVDzrXVfuuYEj9w8AHuUixMq+G1nt11LzW+VKt1bH7eujRQG5yerCdYX656zrhDL2m252Iz0dw
oqT6h9uYbWuv/heCvDHqUUUZvzrmwnfdlB3N0IxJQUJnAKgy/xNr9gnqvbFrtWlMT8xDMq4z/90/
UqT9Da4mcMb7DmtZw9lq49+ERPYZ3hVC1bGoDm9+qtcGA54A5NudKqnUBYyHRN2p3LGA29dJyr/4
EsaSHBJGh5HLZiM9wX7h7qRtBMWGprukI3/od0EkwsqQNK7sq7bH91rEaiLuEAN2lQ/pS0Onli51
AIt/oOiD8oA2X2AdVNlLby4y5ZLqCcWErmV8FpX2TibWiW4JbCIUTlpsRuIxH0PygVU8tH5JnN+C
TGs0K2p9lbPZ6kHHrwUdhiquh5oNU2J1IgnH8RosfsbJcTeEHkJ0XQPasWF8SjioHC+sQdfU5tpZ
up3/ZbP8Kx6efhhUNNHkbqamaHC2t0gFGDgCP/GdgSzdOB8VP55hbJjakQRoWzp+plGTVTOdszAH
M0vzgQrZ+i2jDJHxpXYW02krtP8qTT4vgZA+u0d1EFsx9Xn5luJSr9FM2rHohYhyoFrJYVHMf+El
5++O5iFNYseMV+z+K6v//eTG9r2QdQgQAqzZtCt821SRPEktjfqdLbDGJAaLrDXrdWw1dwKkKdb3
hE2MiCQxj+WSjYawQPwnyxJgGVDqg5Aci+0nlnbt77befhwtoaL9QF0ApD5Yx5bNOdlhi1jbviVM
MTcqXk34SPFRXaJ7li4sV7mCYtHGWtRjahtUBRE7j6WRIPOrm7C3k0BzVGl8UJqBcGZXGk/ExKPg
cWAsy8gcQ0PP3OHD6+B/vQG+FsR3mNA7DSQlCQ5VlW6WUt+WdGwuB//tZIr7OF3iQc/3/MXu4IrX
RZUO2LXlJiFAw5MVlRfEumsesRwKSfbzTMxEnaSP0RY8k+wmMdaStriUWIWTkmCMIvAr4dkWdkpA
flXAX2K6lOcpEGfk/JCjIuketQjBBWrUJJwGh30u6yeVDOWKToFx2lALbVq8lMV7Tt9V1uKovTJU
gEHMGOuBI/ghYOQxZFQY0JV/cctZiipFhRvre5ckd4OTPLBinxaCxeFQJaPQ7BqK6kVSIgB72xao
pNSIjrhxGkNExLK41tSZCAZm1chTyRQhIaf7wZPOmfP4R7PuBcJfSh04RG+OdViPVHslsIc2mbuF
Cjy45FOoBqee15Hhx4ExBGDkGs3Je018GouqZQmG99Tr9E3gukao1NIBnorLPLYzXw95NIUauMo5
AWhX3kt65T3D2aLiCsdorJSkIT6swy84hWV+IvcbAkCAEshv81sTBC+PuaCW0SAwkPEE2Ylt86oA
3DUb4cIerf8s6OVCN8I4r3rlu4gpAUJ31MCtbMzbyTDFBaUxIV2eVJ/D0lllQHUK0D6bSjBfN1Yi
eYaLg2RvtCp4MeeFb/YOUfG6OXPS9jtdyG/IJA5hmsLixGanRa/S+LJOZjypLHUcZ5k9a7F7mCB6
u7qV5oBk/rjioQNR05PdJ3KzEg+yY8BwLRPXoKKAEX18U+/dlVjZDMsYDc94oZcSYbNV8/u6NRQI
/fbcNewM4Db1It6ui3jzlBPXe/YPNmPwyEVQiQfsz9cOtXlQHRdxB+MP3+9QayC9+Wx4OLAC7Ryd
lEAPgcBSx1/fpDp8JEU4FAJSMMRY/SVtsWfmO2KVzTcNLduub6Q0zKt90vRhWm8TeFfzLJmdafvT
0ul8yc2X7hoPb/VTED1l6oF8QwUZ/QuryfHgxz0P4ZOu5bHlWF1f7ZtrCX69PARuGcXDTosdTpUQ
49zLjnLm1s/OoFmGuTWlz5zEaI1o7M0n2InwPe9ys0+s04R0xART8eJv+ERnWwmmD3jP0VCVrLYg
0L+pMsp8cHobKwSCfqP8n8CK+aGbP/G8cZOYTANar46uNUIowJr8fPCPuvRDRE55H2XxXrPLbu5r
ScFDapPp4VD7Z283huTZzyKt3U7ohkFQPQAZKzOnvyCmN4Ch1TuTn69IkE/mQ0EsYgYVIDi+bQJU
VbYg+K5r0MMeFRMnOGhgQbIUjWfdT/R18nXRXhcuWstaMJIMBl2RdCjIzWlmRe98p+k6JgQyDn7C
Zz5P6McFX/dQP/ZmycTF80jgooCkQuMtFC8K2cUPF0fbfXK6VCwOFpuGqvKY46q9owQ5JevXZq5e
jPcinO4S+ZHTaFtvoKvIHZQIc3Ppev9EbNJ6IYT3GsJss+YDDz/Jj5yz3lTEqNBSI9t4P0N2Qjvf
iidkDp1CZpU84GJ0jyeJ4s7BDMZS1+y8SLZ+0RhFhZpri6/4++UWBz/EBu0zi+++LJY7D92nWJd8
+oJdgtWh9xj5OYf306+aNsn/jCQ4ivvj8CHJVpp+39scNPBHvSp7Etq1+PrCesDbxseHPqR5RMtG
bWmlJAFZ0YQYTNF4i8FDtgzTdsuPFwOHOL0oB08Lp8hR6cNia9NnVv150poRbWxa4T34quAOCz+4
Z6F1Lxl3cUf9m45luRCgLUNwV784QLCew8vxWVUVamxjy+CiivZdsStQ0mhMr6gKKFIhGqLyWSLV
a/xkxV3pD20p/BoX4ZnTOECVeYV0VMQb08H/qL9pVii38FEnA23TSpd55D+/ize0HsFxMsBHTaht
d3d80jmLpVNcwybM00518JBFtbGXT9jBfCLQbq6vbkGVu8ZZrNKrZ6azfpZXqxUebd8rBNe19LGY
7xvnoejJgr7q15i/oRdIEu5F355uUNBkMzhmbJhSHBXJ34TpTG14rfii3JFquJUd54w8IahYsJRH
LXjrJg6JB5VFBjpeaoBiUyU9pj2UkcHjjQqQ3UnFYl52a/TW3EnhUJ3O6XAOHLF65BdpiirpHVcE
IiaY5lFjw817L6MzbDBomBpbgdFwxU8k2hZy7ELta3hrQhHAx+j3TWJ8vFcigBigoU6cZB/vChBT
0o5HMuj0Qk2qnmG+6v3vp8Hv4VhOdE10edYii4Wzo3CucYrhMoWipZmQgYyfuAUEK813N42tzolJ
IZYU5HS4VSRO7zNDVJWHzr/BKej/5CIYRpTU6ELo+Pd5RjE3ab31Qga2hnmBmYQBh3uoMAQmo4Ml
9oDUlcvSCgyngQTd1p0vNjEPtnycJVZltv/qSKtPG+2StgVD2wOLUuPW9Dj7WDyCOWIE8cKdODDz
ui0OreAYwc86TqYyFqcFc/6g6Yl6wsVrIpEWv5/lKhJS+zCFqqxZ3rPKM/MY3fV98x3/LenMr4b/
X3HhKg7vphSDqOyUyJbZ2hiWa6us1vPIglgWvgPVbDvXdau1Fa5yKlkTpvLDhLyn4F53bLfrTT/P
px5ZjlWlLLuImpUsmHsZfysa0Qygo9GuCLmSz9SBhEVuAHZWSO8I9VWVhWVDYEETELaa54RbSJZy
QiCYwvTYSkam+XsN+CmA3tEV4B/RP0lib71E7+KBlZBlNXwB2NBP621N2EQIPhmMMjlUH1vNSwpO
gKURL/px6fhJhgHtTsZOcmSn0nR1GBP/ZS4Z56JGoz+mHyw1ayQAD3BMFtFdJLNpHreMs5KiH/+5
RAVhZE4Y/o+U1xW2Jkzgc3TPcfyyop51wSgjxdM5muRby8V+0iRGRe/REfRaoSFZhyUSvfA62UpY
+qbz85ibWpNihKJUJOGujdcj4lI/4cwtIEV07ZTxdTRNjbrKdu5D2aLyZ/RbybxNyXz1jypSrN4b
RBXPwocT18ua5LXgV6LXMKkgNesbiq11190pn29UCFyKuUB4Bwew5tHHyCQWK8ANOgkymQ8XhNUY
YJKqEfDV9W014Be6xAO+QuXJiI+he95lDws2sjGCY8giy/DkAugS5+PgV3yGc82OaSyEsD6YLwac
TVvvWdNFoah3cy8aQCvvw/vfKV2XHn/kQQktZyv3vHf7VrYqYTDktYeVYflV6ulzVJDb9X+1mMc+
hazECWY2pPDorpIhX0pDj61FGx+lAkjfWLou/jQ7b0ceJeQYpNXGqWQDzHy43GEhPOzCDujc4cQ+
Dr90YiXlhDnCamctw23ghzfnsKpxSEbe+UUOEps4koEaiWTsuehR7W2gwlaU3aL+8ORkNWXtIV3J
C216iBasSiLr5K7NqQ0cg/2ZX/PWe4o9+1goznvBtBB44QVa8Jc60hdQbExLgf0ba8YfUQWWFcwi
L7MPqApMCUoyfgtFZcyqQ4U9ytGjcmD3C9Je+JV1UDDkP22Q0n3ST3nHHuu+MlVt1g3Wg1vpPs8e
aGfmph3PeupIHo7FDuEcnrzgN7MwshfyyOjbbdCgzkcF0sOdeKSjbrqOV5r33feZTA3MKrPEgjki
M0mG8rK0BktFOrvRKAMuZiDbmZUr9RY9OE+bS2raUa/xFbBo5bpSu5ndWirIptJ/E+5ESYHl9jFt
WYCqSz/x6q4O3EreFkghMO3mw2wW2n+HINVrBsf4zP/qtJTDvc+vhb5IoeQAgPhY45M4g3xaEjD9
LP9uLAjEE6klbScW9cuKPfnAZyJXIQUmKduWgQe42G6LxEi6BEEeqIXiUBOPTb7K3QVQt3hE3PUU
Ml4f0KDSi92bJlqUPazHynFhYoA9vH1RT8XK8Gk5BDFTRBD8ihkJTUiJkzEG+Gyb1n2+j2fCYgum
lLUcoITfLQLDDtWbN8fNRLkg5ii5fCDmY5SxZMHCP4UHg8TQFPjSs5XJ/PAsrZclByzmqWC+jByp
qX1AOWtEb9YiSChHOn5vQV+zuubiX1yuSWl0H6ZwXsbL/kdkjPRMeWuwFGZaOOuyZ+LFPjW58Va/
vi2KRYjj0umlIBb0oO3aatZ1RF/Njd9q/14Sj35w3hK0oh95sMfIOtfdKKUGiRNooF50YiNIapUG
0Hvso2n0E2pNTP49GfgTXusv2t9/9F6acbbSelfbbjAWIqcCaaO67kQuSnRxK3FQilqO+bKWnlpJ
ZnyUnMf2zVxRGeZuZxOtzErlkcpS/JpHQtOhq9DEpCL4pyzfgPTVOSHBaP/XhkAri9Wyt+gQOFHH
OAlXKMu3XEyOTMojebH9Y9lsp2gRbUl1ymOlZrAk3Mw+lNmtq2dN8ZW9zCw9dy4VCVXMhoYSsWu9
IUPDO/gRUU/7BOEuCkpyyMXlwTxKNfe8LLXOqmc+/X/8OXvW1jUVsgfSXY8LrvR9F88nLgFJO0KX
wwnxkEZ0VBwsr5fdFDKTM23m5VHktzOPs28a5Kq/dDbTqCDIqjNeQ6MEbnOMEuxWRvJfk7S9h+ZU
5mXIdLS/6FNlxCvUdtnYnuM3gNL9FH20N+1J4OrS2cAvMDLuW5Zn/qRj/7mC3C9yMhi8XhpHJIuC
WnJZi1fq4g6MEdWJe+VpTSn3EBTL8oebZ/at/WHxoEytuyqqk87IWEPlWrRqMrk2OwZr63mkRkuh
+k1noKa52m/E8FUSogV1hFa004tuOVFphz+NBfkq8i97aYCQ2eaqXhOkgEh61yWvWAMFb8Qtt4QC
a26ws/JbMema9p0YcZC05sgDk4vQrMIosELEnmlBc41CtyGKxRhCnFd6yfycTKeu2MEu73l0GnPZ
7QLz12918SPh6groN03GnVFHE1q5dSDwqAju3yKBvHTK0C8jU2UbjWcneuBteO6lSBdqp0zP9Nug
wjoGrXmHTgfOEiE26SkHFICjeRuu2EeyJeXgsODBzzfO92vMyx+ompuZJHFVD/srYKs+fDdVZok9
DeA6ADvBbKfnxoK/3dE4gg09lTYP4kq+FujsaQ0roTiJg6j+LuHGhuh9mjCxlIKS5CPnTPyG4uLc
RsZuvaQ635AvkBLvz8KlaIfH0ZFLfW1S4S34RMfZmY9lkXCSj24rbOv+EOzfKnPwll+zSTBci27k
ntTF12j4UHYjerVBVlPiyerGpPtCI++AG4mufZFx6c71qrF7gnfn2vV9Wl9Pruhv5NJdEKFeStvL
BHxKcTpZDTXX6nqFeL4JsdESSH0KREhhm6VSqmNEOm7PtxV1Nw/H2BJLCfehfG3s92/9s2PtsFn0
Q2EuxCPysjLaJBdaXdGLGiw0YZgtLMFaFys7YJQ3jd25I40HDTsAgyZslA2A/ZHRbi0axL4RcoSa
9O/cQx60km6kCyPmqSYkZcZqPqo0M4/Up4S4CBVbsB920Zo5ChShjisp1sGaHWhkkmrZWeMJHeS5
rKAq0eIh9WVZEOuK+2odRPkWrLWTqyQ1Kh5jS2WmFDSTuIUmxuxeV1pS6ewMXt8EMmQcKAG0YK8z
nDBeUiIlFsjD/+DKxYp/l8GUh9qkof+3Kh2Cwze6Npw9pyxhWgEkuoeJVr/I9t25e8YAsMujm8Ul
rYOp6n7J9mO/Xml0zSlSNVgKMR9OVDdCXuQHygkS8XFif9sAa8nntlGAW17zkL3p9gW/wnyHIMmP
/UPZzneiZZQ9jWk/wFeMONZyHObZmmRsvb/l5pZNSk/1OMM5GARc6oTnFZPV6Oy5MfvxmF0nH6gx
NZWWN8eHRpXddOknR7voqQnxsQidqOfcEEOSugIFYo9g7gKeXX0154AIIDXkkAjyIoRBdD4Ir5Q5
WwtwPfataX02ebCK8DnyutOdGtPywgQlcLj1+j501CnFFzQh7KCCzxpYHhuNwVi0OuLSOd7R9uuq
n7ICcXjAh8klqNtO/1nRU2QIsZ5/PZ8QZNJFuPqUfvdPrgQOARfCQz4dD5Xb1xkVmXD2beAkYhyo
ElDAEM/WH5AAsdFKoAr9hOU36Cmkb+ETwMBivFtpy4VmdE7NMFnd+LKqI6pZ6X30uXVaNBibGZOb
+DXqrYeVoIwwzs6RnX0vVsXRcwHH5TIG5Ipv+n4OJGq/D3rb47l0QRIV5zOwk3YgsJnbloN+ibzO
pDEHO21/jJyTpoF2qZj4BsI0Jt6ba5x7YeFEbOCnu784YWXAxH4tuau2hbJdv8abQW9NERu1XL/c
M3oeyzeHEeISJqa/d5Npzwe030ypvjG5bIwlKmeblXwQW6f6A+XHm+lbV9cEuO/l+qHr9pz45jVf
SzOtPobHNHI99eWYhrvwvax41XF3DkrO4asb/IkvBF4qlHsU5MgjWnDPx2LCYyr+ps8Qr5CDvB0A
C0mLcDuU2WeyEem+m/Mkjg+bCDF1jtr4MptWXfS04cpCqt1lTNFw0bbQSbt+CRZygQiiqcS73Tdc
qG3dJ2LPy9dj08kzRnzczNwPVPMz0CGKgZhrRM4KuxbwxEBpa3vtbRIwxVwtAoPsJEIdV0chIUs9
a0wqliU0/Oxof/bOUXzahvPHUuxCXTiWSCay0EZtvSHhvWevw4yGOyotbw4btyhh0TtcCxNQoKzO
i1jEHiCXKoktuXKkFLxBK8dySBdQMRhqLvMbCO+4U30y47IyYHhReUvLXAJsSOxJOkLTiYIiQtgX
8+FRQhA0VSg0Te8Gj0oZ3fMNKf3kpbHbI/J2/dnS66t4ll7biemSfafPTOdap2RrDcpm92bX1D+z
WbYbN/HoMx1oxd28r0Krm3KcFicxgBZKqqsA8Xx6tlC6/ocjaOXvJ2nAce1yhTbCxB7sXSZfB5lR
WARr1lLALUVQT4NeYp576IKs2undzoaC4KULi0nSvPdCIVdpIQZ8fPiSsRg6jMW8y7JQ88wxQryc
UvMbhR35BOxZggi3Vi8GFKbK18cD3RwAvO05YvOc5ci5oi2C1k5OpRmtPHVaVleeZHmOh0cMJj6Z
5KknnoUKY+112kJWI285A4qWgEEAQMCuxk8yGh729enWzqALDXBstis0MBAjFxaiDqCmNSLeO12m
jqidxiIRleuT9yXkQgmkZDrfAUCGVr00xCPptditIRrP1GJN3Cb1ES3RM6RH3GW8X45Eu8hLsIoE
8jGD/IScWe8V9/2eOJxmkP1hr1Px3n2dBcNtJqYKZsJwdK+LVG3RWtBlzWBKVcktoaXmrmhclczW
5++APRNcyCdoS6r+pgCeuAuP6qUMSukZVJUtHCu4wfro46dDnueO5/+IXyIOzlKybpfRkrnzRzfB
9gKq6HreaH16kWHcBDHT7G9wR5Xxxy87/CguIRhPr/kiXLICWuJZQuvHxrVwJFhSPTGgTjEuSw5s
NJXp+lk1++BwUAoUu6LgpNQ9Tsi5aFmRwFPucS702WAGSgCgcIzo1M72DEKCAWGcN77NoYt6zt3Q
QTvQRkwjqnJo542M50H/7B7RHX7sMqx1sSbWlYjRDv99CYNfucQvhIOsmHhGl+M1TL0/qnhpQJF9
IL9dTExJqX3ibngP1eh1PLs1jxli6os66132weMdwtALN2O7ierpAQs8924LDKEQyu/sjz78QGUW
K5nTCNTHTTZ1yZonLRbppy9pjX33t+7KDkXZZ05czCXLnDgkcmeRsPToUXXtzT2nrXLq+gzECQt3
mqnwW4f5R1NIKAZNqcmXNTQiliusGtUtgslDVFKcQLOIAv8T7VZeNnYvnmRURsXd5AkwmjXGdhAL
jvzZuln7Vu/XpOeFzsvgAjfKTjsef60RZs+moPeVOjCPYFIGGpaTaosRXUndqaRPVlpR+zYp3T5F
iZyMXKgygZjc+pr7ia0mdGMtxw2R9N0VnLPzB/XQ1SxQ5fxk/9m6I+sX5Z+yzDSc9jEfnNMd+80y
zWG3Izvx9jpFrSVKUO/dmF0fVRqSWTCE4OBWJ+K8IsisYFHjfKfb2lqxqG5YBALSRFI/wDQlkh6s
8BFBHJxnTLVyKYq6zFSVnD+YaQd3hxwGHVUODW94HKpgg+eY3Da3B7XCxlNJXZ5UG38+JmNAB063
oF26XPXKT4kIF5NVx3tzF2QNhJhimr/oQMOV7GvYRFR3FTvdKUU0KIrpDxJcpKJPw/tBIP/h0inK
cDgyHzeQJBDKKo9x70dtcxbcA7Z+ARnD5Y+SyTTTHgZtJSfmal+Q8Xijm+ABNEWA8Gl2sldZoSHW
6Neq7GFZJ1NV4zaoxH3UwdY4mDpyQwK/VyjnzpKrtbagao0q/iPwQ8GIn9qpRpFXGqnn51sGtwyR
dczxMlcrlmkHNFX6AgbK3DkVJRcO6fC9dEYugDD7WAUQJLXWmxzWraMOOQ9ETfMvjBQK/umRpLZf
Il0VPdPD9jx8zmLXq66qonzgzjV9Y0SQskhx0+4DVVVWytMOW1QRHpyN0aFvkbWuSBB19ZW0Z9o6
ZZmnIrpG44BOtG9ACPpUtm6SvxCQtIf+8EpEvfow3DwOlhIlq4XlzCsca/a9qiXML5rzIQh6W7FX
Hf67MMRsfYZhAIrIv7rZbOwh7d9/tzHXOtbeo4IpmAySa6r7kCbH1yRS58a1BcGd3bSfIB/lc3FV
2TYZ6INrSfVMSLfyQ4mLNO1FPS4c1QwX9SM093r+WFIJ4iSo8Iclkl6dm/hW1gQIe2cqeP4F8vej
b+AUGduduwwTku7jB7tPtF8Z9ewJo1EfFKzL9KaM2xyYYQlePIGwpN+Xx4w3IRt5fRzFXdqElpXX
V952Qcds1FyT+lrTbw2pfAr0Qc9CJEm4hvkN9WaE50BtxDCRQnd6cBys5sEN8cSa1+AMtbQMHtZR
yMGK0uJoBicyCRsfPJBRnKPLc0b+bubLCPAqfKAhm6EyfOm1TtbIviw/Foq/slxZm5t32b/SA+Dk
ULEZRqreR+JPb05KykOIlTf9YozByxGV7aNsDaFBXfAj6n86nwhoadN+pKdYuBdvGS5mTH2hDDey
gWxgtXaPemRUh6jRjoq1/JrSEWDHXYzv2D0/JPjK+l6FJxjQddkEIV7tbvHD5hfmBjRU5dp1SpzN
+jgMEJXUUEINSzJNWSGxX2LG1EGKsj9q+zzczlGRf20fScjylARkwGwa5HSNePxW3ILaBZnQipk1
BeNAvMZRDJCHuFyIlDjIdfgqPRRSpcQrbzpB/POgCWHJxfjQdxxSu4K13i2ON8liAkIC6bBhITDg
1C8uZUjz9atqV4YgAvlbat53ISk3s+AFvU/KnEMKv15UBiXjF26aUMuVAAfOVf43Pqj4Hh562Zth
wZ5Z9qMWskfdNg3HoB3kNPBQr1XKfnkbQOC7iSj/5PvIJhNspW3zsncYROKDfwkPBVUjngXqyyf5
/1Ot61Upf0MHSENqCZHNecdwX3ETYiA028r1++bwm7NTo3merLPWZku0w5H16+/gtIisjG9ONSq+
/2yPUyEBwsUtMQggMhA7oWlVQTcK49ZCBwZPBegoMVx95gHsh/Oyi+J3z7p3fp0LTLcL6aPMI+Aa
74Du1uIPRdepUGPEqHswvV16qHt4T77T52KWhHx+i3RxaRZuEkG+FffK4g4Em3Jc6TZyiKQ1D8ro
jFK9iROBAkZxvrvm5VjWfQPPihmBezvqYw/G3JWPWF9yB9pTsdmSsyYfRzeyxEkGcTlg5uBuCzOu
x7k/sbw4hAhRPaEzEC7BCKzMu925kdM8MQ6xK4GG32xLtn2BBMPOyRiBqPFt38+oagfxHYHkLg4O
KFr7cELHHBih2tdk3lCg6Z96lSpdjNTbzZyQa5e2rjrdPUw/PW/ycomR1FgcFbiP00rs24geZSBY
7znuRelZ3UYjOZ5sLBnvhfkLAfgoiuUgFO7XleLzdQmo+UIYwGEuctDw84C9ggwLcHXOh7ErLjrJ
5U1eBbpdD6/l61IQ5IX5w596fLgwqAXBawSnuklFIsbV11HIW/ETI9kIFgvNM7ZgA3pnEWJALncE
OjvSunzVMWsOBn+/G8cH/bXzwOJ4b+/pOYIDLgazoYtpYe6Qkl1qB51QDMxFATF+Ar0SSxC4tqT8
gfwXaBw2LoN+JQlx+t0p/0MlTSdet+BeZj5/vcqFrTkhZyNJqD51efvCewVdJV+KPHyx73pzQiqs
fIrxh1ZDHgauikVqyxH9eeBFyRV8YJQzQxZCrqgGsC0CkkqLPdKBI8Bkv1VAdXLQ458MQd927tuE
YBmgFBw/THt4WPS28Q/0zb/fsCL34lUtu2NFxXUOdt3Tuz6xmnbSqVtOfgq9VFploArYUrQTQlm1
Bk3Tgf6PfUi9KYF0HGq3KPFRCLNizYCohsG7lX72n3cGwwxaEfLZ0+FjzCX31XJRLB+rZTnzBB83
QmN2274DXW4nv2jDsbumjvTEqaBoRfa92t57BHxyA7Q+JBXJzaHqNoyLwR5SrpxQfRHrRUXmtyzo
oU1EILHtFvPwRiPwQ2Pdw4LSGhT6Bf59oNjFUGBRSw4MlCFMr4gGGiVKVWCDl26Rwc4zR4bdEVJh
kbLPNGXhxvRo1gDdiEH7KoT4scDhY4PtAf0ODJRvtJ2RuOn4l+HxgfCZfYCI1NcuPzZVfCp5AJ+V
DSWntg16K1OObX4BrJ5dqYdZo7E1u4i5NByCbZuaPsaElzePQiGZPjcuj6dQ8qQZCP/1J19Wjl5+
aWN1Pu0ZxL1LqkUf4H9zPnqxWSa4DfvklvipEBwAazBXKgJ0e8UIcNOE2KbQWyMu6zia+tNFr/bF
L6/K1LN8NK11kO0ghTffm1IZgnQ79qaVumuo/GYswcJ4p0HoU3QXbfIdZTz6DK0rrRv7ngDaveR+
51rmDPmuCG+q/jxIzmkrS7QpAE5wbRn4yYxLS/wyUt0lY6SedAezUOKHyIm5kzcXmTemYRj/V5kr
BcYtVCVpV2px9R5qWUFD0Zx2hKnQAQnHU9AV/Gwc0LwBubcZmwoKOWKCCHgJdTQ9kuw4S6LAvAiM
UdPz5TUb4JHfVOU7wbJUhUJK2yeLDZWWfZtL42x+oYKbtHn10bgs9JH0iki1AXe5ou4YJMmzEv0C
M5N3nJnnCgM1GseENk7KrYvz0Y8ZD0tSwgfngngPrZqRkAbY/4gW41LX920mqpkIkRGcBPu9Hfaf
7/XCedJj+kBaroELYjP1EO+hnIOKVu3FoSupVFjS+3P7Xyjs/FWCziKAIFayM77dDrQWRCAIOMWf
x0BajVVztXGYmlTAMCLHrq1BT6NIj/Qtkk746kRge7TXQPWqoNxSlyUxioZWq+pCNfWwKJeG76tx
VI1Ch4rQVSQWwVVtrG+0pNAoddZvoPFFXTwBWubK6WE5lOBJ8yByzhVtzq3YOZjnLruhO+A2PZ19
s2pcsENdSyYSvb0vOucCUBk/aA2mtt8qAT/4Ods1k9fYRwQ2oflOFke4wtvDhP63uBJNtmeBmGXX
hyXbhRZ8K8ltOvpU1ardpN3ih0KvZvg5nvkaUtk8tWruSp9Uc2cbSztWN8b5FzamqJlSFlwGIJa0
QwEAj6f1pylEunnewy+L1rqIYS6c7X7oNDRONJFrQoAEw6KbLyeldFih+BHTA297+VTV7Loyiybj
TplYVR6SM/FFHVtEZlP1kYNr8UR0di5iKOyHgYdWehTyEqAQFJn7ltr35GGkZ9iZQWS9xWFB5aNd
0nQJdfSGa5uzfqgIZf6esOYaR2bfP1kyKxgVU1bjVKiXym0dMf0ltPdxrMgFf5Dz1hGw/Bskv/pA
If7gle8ZwlWndqWuvJ2mR+FLrWpJ/opajUjqsNbdxnJ4NqVwtWfnwXoU3Z7Mh9+b+bklhgdL1CVb
OTq2jQ/nN3VtcgLMru0cCmvJbW53oVUbj7y3KlUr3N0GVWtEv2Fu1yhSZJHex1J62Em8TgZ3a4o0
2DGuytgYOtCqPBbt5aQGbF45y8WUa8ZU06gx4FOk/UZC17rZgb5d9puKZ8LP9zQU/cehT9ehlZZI
0+hGou8SslDrzWJ7uJSgqPhE5IcMqs/3Cw44SpAvc7570WVQXWLmwasUPNq+2+RUetJG+jboaIJF
TBdv+wD6/LI4/fitv8kGExB3v2kljEp7qXwO2596UZpy8IxuNBh8xbxsD0BDRE15vpogK1SBlFw3
2rZc1axgoaWGAwJmUtEkDtmZvJuG9OApnmpIoHRils8axM+HxRo0InGugvDO4Qh6Db1Qz0Anypoq
25Do9/lIpEwy6NEd6UtWJ+v1kKyMO+2++aViA8LMZnKBF7FkhQXkt1401kpiaragta0eYlP9P4t0
7Pz6d7ItLOOiBmmTpMOjgX9kBRiYuU/Yq0+wa2kWsxbN3nlaGLV5qr/WbKXHmy3ZN80mbb1hHIcb
4jsWuLGQOlFkZgcPp3BogImMuW4gz5y2UfpMECwloS4MpMve1qfg1OWSaEy1qrLSr/bWk/OT/mKb
I6ETfrJb7Dsbb1PqjF6tcOJo49DtJMShvMBlO8XHyOePHsm5qosGp/l1s7pKUHl1f1Sace1VVko8
XJG2vCiO30fnRYKyI3BQk5Yan0kHxTbWDhx2r+uL2OWbuO0+7/XLCQUsZ5ce6lP2ahhwkoV+rGJ3
3bfvTywWsaz7JI3dNccz1MlNTnlUB7XnBi9yLg5Ym3V9JhJgzyk1yHaNPPeIBh36SISDETqf9JEc
9B5O+cgj3SAjhdFGndIPF88YW7Q/z5N3U5Cs26yHXKKiXDXUrIu8yp4NKc4YmJO+croGDchEyhOx
B2KDU0jrkVPIqMSzezxgYDTE59XkKgPSsgOQLjjwQHI5NIvqBZl/DoIZH7Q1Q79IN8fMndE37Ltv
EGYCWxNLHc5D4aJBdHjm9cziEGCzxCd2RWgTRL+hv/B2O5BvzI6kJBDqYQmPMPk9aNUqJcCcOj0k
CQeVMLek19NpIApM9yrYKWSCURGb9rCefuZBJXWFkGWDgD3rLJA90KIIB54bsDi9kAhzsph/eHEo
PAQ/BgcaSsL6cnUs0OBkf64z+sGOw9/L1xznuhL13Tt08nJl48AJ9/8tTmDnagec1cwuRWSjBxqr
VbHFi+2iR5/yiZUJHgLuoGyfCfBZXVi9/XC5FQ4JfMcqlNsb/+kSBM9gcazQ4wvBclBQNak7psep
HENKh8OTo6mznc3gE4hOIauJrVb7ZnU1CZqCn6tSlYr2aWoIv7CovMKdVBo+X9viNbeIke0UJMSF
QGK9JctjVMSaRu/0sZKcaFrEH8d7XTXsWlxac4VetULfNMkzrMJhnsK8C+YUEKisvxrpEuIVQuna
4bHtUOQGSbk0QemEcon2sx9IguzMOwlTMGusvdWj41kkATy7iWytXjFWEh71T0Uzgh2w0T6TqT9F
sJdcMSmELtKPkCIFOmUCvWClnSWJlxRWJ/ov/RFc/UlvCUANZIUPc5d+DtKYMKx+GbeJwqcZQKk3
I2FmhTr+7Zs2ioXgG+vV14o0t+kdJK7kbi4JHRP06utraaOoHStTX+80nyxWoQlHgxT6GN60QoUq
9txxOOi9rgeLQ0RxwaY7B6QTN+eJVr3GCgOzwNOlc7l9Zs7vS9WPYEXUVa11zmyLdLOyXzSY1eDT
E6A1jKqxtZpdhRCEF3QC6oHUIGXb+P9X9c0b5PDeZxsxJqTNFxVLxejbp3toMVl89YX35ZJH2sii
X6vIVkvBqsicjR1FemgRERr/2+jd95Yh6+8tk6wmE3dHfdrFFHsIY+zseVxqQkyBvHIFti+D2EjG
aQaTiX0oQMHAlcOqBC1QcG8jeyXQmuD+HBBwL9MEsV/fc7PWBXrmeeuQiiWcP8IYWfG2x2FBJZ8/
80dfyw3JqFYHhxaXHUWZxf7egJmD1pwnFxY/j1QC3LAYrBNPANc7m1X+A1CpjNxEbQ0cci5BAKrr
MlNtMojP9VwGbrwAO2aGXoKk35aDD+dPg8fYiZeVJ1JFOQFQYiCGVP7ZtJR1xjzXeNI5iYZdFUwy
qnsSockV8Yu3DHcmJ3zfJ1BWVXLGmmOc9uuf6euXlmCZMX7n6+TeVdTLJ6Q/woAcjYlfr8zREgPZ
Nx/OcFIjRCUkaf1k6tbHJrK+XjU9T3aqOtH1M3IhfRYE9RiM8N+xHy53K1JKkAxG9KNhdRgumuZr
Pv/6YQsf30tz0qgsIpYXltnKku7X3brhbegH9mqmbt2D2w1yPWTPEHrYoy5XWoHfSWL6lJbkzm38
R6Q+m13TOrKAjLc0i/JQtzdF3POoZLg7fZ2k4YpSQGBWzvL2bJ9RXc5QrHTBqDRgQw6lAsw+O6/d
FIYyfiNtEEBKASEPtOLR2NZQ+sc7p1yOiAlJiJYGSKF7G0+cxCo79H0MZZCHqRFON5Vklaa/7FWI
k6X/4s7EA8GsFt5yZt9XjZScsrGazyVfpFFBjNGfYuOQeFRAOcpQGZM/xIwZjw69oHglTVg8luST
lvUT5S21RhQODeYNCRL+VT+HS+8fNRFDFqwM599fWAaNhf2sUWDbiIsNVovmh7ALF7Bdi0lWP4Q2
auCNnjXLYEKdrvuY6PT0qAiaKVaJ6MON2ImTFDZo+Wg44fqryaMV39gx33vqXifOUG62aEaDnVW0
Nz9FiFKMZKlmY7W5k6XyXt0b1yjtVrIxVpwTp/1iiEjmZFmYxLfZETWoA0YONkrUjV/ETYu0wrrh
gUID+yxfoQEUWW66QsfzlEPQ/NyKw+giJC4LdhmOwGVNc6cKV9+q+1ZyIzQ4DQWyVUotkLA29Lf+
n6zRHIz5an8/IzXP4cZuD/nkfOjnvuhMyAPwibwPTMMQN61j66rfU51JB6blaejpKQdJLZbd+IsK
e7g5dwRv+QyN8KAeCVbqeEXQmIQvJghler4JPpxmst/llGpicNvyViryivNGBNC765lTNDoURkk9
zQl1WDpxs/eM/+xq1mOPCLaeFBYYktko2YDZZhIpalwVCuwWsKR8PR3dUxicv2yKxath3irioCcw
jc8M5JXi8LIMuu69V9iRzrfu95kGUCHvI+3Axwf7oQ7k/Sf7CNVkQFxqZ1auqMxjNswYhoIumb1B
xgWuWbwUohULNSRBdswmpINIIKftxNIZkewHh3uqHMGC9ahl3llRSJWJYgSnbLPvQhD/vtSIdoWD
3+l23AcqYtYTlXa+qWr8eKtwsvz0MlkzVMtfDdCW/lUgfTtKfqdG6mzssrnVuylF0/+Uc4uZZAFP
pTKX7VTLMyzcTWP4MXLzRKshNsr3FGyRGrU/J0SKBlYPWaGQM3xuqwX9MF0g2/pblMG4C+ZZJNUp
2KkuFtqRd1BUIQTXEpjFzm+EEnuHBZ1rtYoyOFrSuMEqZPR8F9zPR8NKgKR006JpTHDRkm+mhHyM
SaJzGOutnwY2UckUK5zq8Gnl58Dv08XfbbuvBCqfxE3IOhgEkaXCyT41g/MqG8qyJKpVLwUd2cqd
AoH3gp0Zfm2UK/4ScVnG3tMgiiK5dHdJ5zsZq2CR07H8+3oHDNpLVjw3ACBgCWWnUtOUOW8GnmTH
ZAMZ46fPH8nPZUjpbdtBFw86yATYnGlALwFQt+kPx/KQl/meymj2svMZ16joKjqz0CP0uGNN597Y
05ohDTWKC2zqgZNZq5Yf7FD37XpFwrhmqiSkkzrwX6zUMdJqPeghI9VkXMTZpim1zIDnUYnN1pyk
yEQDSWndYljvJLm9BpKVSqQIH0bNBzVy84AhiqAwODRHmtVQt7055uvP52OOxo5wQSfEAVqu7Otw
qTA2XBInop/L7xlnGNFxKjEvss3xPQA2NThIDP4Ivlna/E1cSoY8j1wQVP48bNqgkQDeXJWOOI65
3U7pfNUaaARuC7PSBjYwckvIroCTOGPvmY3XB9fNo00tEmWE8kRgQ/7+5usDuK+uuuWz4wT9DZPr
lJn+QWlRGE8pmf27D+tqaMBKZRxJBqo8SD0oen76r6xvnScmYzu7mxV9HD4EDhI51Bs4CFZZFTOq
lpHO1FYNnP1ADx0xxg6SwmVKhXjYb7f8iWp62W/4fFCPNM+5cf+GMHuzMP9KGC9E+Hist9OzIcRt
RFPaXsF6zhrypK6ZZLKGjygCd9TFeVPK8MZtKhwf3ZH2GiX5zKEmeqcjOx87md+pfAeqBYsiz1Lt
h+a2YfpJjiOIRUR74ZIPZdqR15ZMrG8rr5vO1o7r6rvzKRZbpBCFVvvxXHjEoefVTG5i23ZGKuWp
EF66fhp6huMGKO3MNmtWc3Zm/exaVGodTIDJ1N2kXYVnX0JChLNRogoMsMVTJEgAgEkHcTYmK56D
OmroyCrDhhfrlb4Dilu++XxevGiGLM+avo1GJOrOK2J41VfsfO9grw8KjFIQIxsXHXE1QeejVDUo
fIlUYSSZRYsJnmECeaXPILse5zrWJmiFt48IcTPKsOal99HjhEXCD2KDUdVQDPEZcKsVlEIJDaab
u/H0hxuRcTR6QyddRXa+7Mgnu5EqrL772hg8dzC4oO8duNfE59c5HTEP+DoTEkWu4b/V86e38beY
K2nZE7mGRfR+uqGpFVLb7aM2+vxN7B9ZtyCneNbUEPalMw2BaEVwI32oIUe3El+yatTj9+4u4sKb
+fBb4TfULtT5E2v3WC8f/c3VRWGhe5C0Xa8tnGd3dwOfbzqWaAqBXK5yADldvTHgaEgxdwygNrSA
JpdTJx9Or2RVqyEQolXWEUGjLjgSPk8Pv7SNc6EmSHfLB9gEb12WQG1NE4ORysy8aGQqWxt6dgnI
vJihakaiT8V1O6fIVXI07vuK5I3HQe7tgdtWfQlWtDR35NUSSKsIokcT4oiW4BLZHDb9hVaFDZg5
rcom9m/Jn3gEHfE0EVRPzbFmWkgDv0MzJEdlZeTSR5Cd05qHcn+c4BC0c5C3ewQQakezgVqYE616
jMrc52WBs269l+e4cEOMpy0ut6ojZaVitKpUq7ljpKyWIMmFyNG9pDgBEG+2ovmxIlN8UPcOA0mC
kLOab4T3FweUwiT/+Ser2ZB85fQ5vmUgL0U4dQVpBV4mV0HoHgEhQzVOyS0zxmjSbU10jhlvaxH7
mH4EtmgWwjsB15/18bxnck83OeOKOaJ9XXKLX66+5IDECu//+4hp+/HCM5ZXhvEBCYCMn8kUgmc/
G4TBmhDPlkxTYKEkeLjz/IPE2imG4CYnv3SBfsS2aAUFQah+cxkQo0l//Ublj5XvzHkt6SboZ564
T3VxhOaSLB5meticd2OlRIhm2PG0640e8wUaNP/cZn6xF+Nqm4eRrL0cCyoCNrUP+DxkukPhzpBJ
Mvjm2Sbakdh3bPl2lN25/GfK2CFuBQJB6a7ivmlm3xWv1LcH86s2qLxyTRyWAcH71wgDJun695Xw
6dyfh1J3GfMjwRjKT8uZqIONbRdRJ6yO0waQYDpMkneO/EN4w/o0Any6bjMFiBJPozBYmiywHNht
lM/M8lAXmTldPJ3XzfAsmv0ak5s5CNT0VF8PxEsOqjGnjqohQzHNJeueJYwqrhrLKVlTVHOaOdpo
KHGQAwCXun2AYU3Gr0C/fO70gZjmXwmPr5ULf5jdN1SMoHU59e1iri6UVkSTvmGfn2cFIi+3uZiu
Iahn2LI/Lt+u/eYrkAedR1HrTXzFklT4SM9XqUVh+BQRVE3PACZqh9/xupIvqME+NFga/f+6Neaz
Y3vxH61t6HHtGiy5Qtm6ytyAUOqHgCqocHL5LxshFiCCKSBJm/rOpBGE4FM6z1BMlcwmZGQXaPrR
BYqpax1RsRZidIjzhF8T7eWm/5yW6I/wef0g3zd41kMYmiAMX2Rom1M+C4cQEpjpDNcFQcE4XPTt
WR0tnKV6mzVPgCjIwxnt60fkQlBah525NHoYEmRMXB0EcE+Lf9/c1JKXQU5HdRk5bsSQ7F0cBfZ1
WBB1C+9cdOYfdOAzgbajt2F6mltmnk7I4hHwD9EW31eMe7KNuLL80Pog629J7siw3JFLaEqydvCj
llCJ/yXEbsfpKK3IGuuuZgJNJ5AN1dniS+17XBlnU61F5HceKIIejs7D1wgJkOgD+hpaJdp/ef91
WU6/y+zEPt1FhSxranYcLgEFli19Na60b+2vp04wVk4UW5duKkRwqNLWg79kkYmuiRSfh2SGSJeM
cL1Np4rodltgnq7OKPn2OdgDBHNXt5QTB7PLE1wky9R7iA6nVqUMox6sDAYykjD2ehfQOMIHfbLw
JFpzrGMlwpyNwfYp4jhH5scvDF1CCMQGZPe56MVvXLPH2V4zAPLVXGVXApXhoTRhU64BNqYvXepB
qhc8y+VqD0pWvbpqovDh13LQGwAuRxUYXW6k4dZLY71fhuokz1tdKRSSrnNAuaJWvxloWPot0LNF
VpBPRiWwhxEVcf7nNitsDOts7gbnObk8j/dEkdqzJKlmObc9TOl7XrngqxPBrA0Pnt0B+c3yKUWM
r71IJfHFuxf/HtlZorksdfxaECK19knGTdpiuwf/CnLmlEyO74iUqZba3Gsq1XulWxV7xP1iPt9K
Kwahk4nywZNF0IsbDss48V3e0PYyOEKN97jM2vns03L+jhJe2KKw6Bwa9BI4NLEnbjRuanmtcYR+
5XISLP1UFuy0GUVm/wnvuwsMJaI6kF7bwHFByjAl2R9nCaoEs2/MTY/YEdbwVp46w+/KTg/ya7d9
W9PTmqgxv1Ojogsp/79EaFEE6eFzvp3Vn/Tvm+YJKeNQSzP0uqIhk9LnN1tazYhTMjDXTalwXR2b
2sJKH9Shy0Rq9aDS0hwr0G9jKRsrTjcxjq7XI3e/r1Ob6s7Wcr1HsXih3cyi5x2DxBN1wxeNoSoV
C4wTRNLzU0rEq3+qhY/WIaxwrEFQlMdz60Gbv2h+2wbNBaLtkDUbR+2VV/Eh4Cs+ySfmFtaRNiPw
lQKqjqkNg4/cNX6AEDiOtdOWf5NDOgFCWi55F9KOM90s5QIX8uAKVyZTs8iMtUU+D5dAgY6bErKj
DLPwSS7uAvDZ+O4Te9ONKnwxUBoHoSviM8slLqyL7X+JinQmdwzHcbUt9ZyZ4wh6PwO4Qg9K7pHH
GVmqmurUE9W+hDE9lNYoiDuAmhf2NNhpVB15rkd/LiulcWERQbQL/7uVUy5hvsBEwZY2KTbTitMI
Q0mWtVOTRNSLWtyKjqy3MkqF3PhEygzpwKaU2upDX+jeNrKSxFpkVNgQ1dZXHm26lklw/gSfaNPS
j/eS8sJXTkRJjJmYoD+pGSgcvQAqhSNgPISuMNRB/kdpibMyO9pI8XxydzQwwqkxptNrkt1246JI
cJIb8PUYpOZlk+AvM/gX4rCMDWg40aGXhjUoGjRc3HvQQ+dLXI3wB0BWuhUcocD4QuW0OWWiU097
qYtfDrVXv0nI+cZfTcfgjxNFbfh25orgoMwORgT771v0ibRpRMg4VSp6jc5agv6mY9qbbQs2zV+u
iEE1wq3m8nRDR2b9mvc8Pj3mJ8zq3yIAHe/9SEVDZM9wFLzVj5PU0lDm7vHYpF7uJfdTnOUEoQJF
LlWIjPqxDFxBuk9w5QjOxE7BvmGwJ5l43zvo9mGVa7NNiwGkLXhZaqIXFRf9Xe5Swy6t1mvrq/rp
H/JC4ufu32Su6DSi40p3KpkqMS7iQUAQ7SnGwgihLG0ZxFGylaMoxIDdsqfiVkJH1tgKFNlC/JL+
s9sP8nbJWKeWHFEPPh3+B2tlLBJ3daYnYsNfir2gI7HOYINp+lPQ7mQEkWHmzOi8819XZKQaDZIA
zK86mmMM3Bl6tdj5I7cKdOVj8khaI1Fml4eDy6+V6GuVyhYhkAPDm+st+kjw9OAj3zhcVsHYZozS
JSYn718jsedxx5CudcA3k3p24bEu7eUJb0AqobIicUDT42hXZCTEaPNfJGhXPP5cfNTsWUrzebUq
8Dr0lZJZHgPoSY29hXzFGju/PnbTyi+xOcZZSejF64hDlS4KDkTScfG/TxoXn7etnz/Ixd0knwrO
2npUAodlLfVBew+/LmbNJ9bF2FhtAF+g9z1HwVuFG9qXGS2OfAgs6SVik5m3omkEoXjHUhnxe01V
7ATs9DyYXV6ivmp6n3RwcPAT6Gb9A6pLgh/EdOC7YEQYvEXMmfwReW+CuBQdMXIiNHTh4nIR+VoM
bklLfDfXooJvcOW0u0Tq02x58e6fKLSTPlc0b0wrS/AHbdf1FfrJOjSafiw4MW3Bhz56MdboOU2L
QQBnRvzR4K3CNBzG/kydiFZoveBIVC3YfjZ1/7BCVdlfRWMDiiCBqHgk2LH2qTe5wq0xa9pJvNRr
+o4v+dJILiXBRtqNTCW0cQShIH5OqPO60w4QPUuEe3S+UIZdRB9Yh4MIIVjLyJnPmANXJYEmgruA
fgxHmyZqNWHdNJktz1akdR1XGAWX8+RzWhIp1LKD3I4QU7RSZ72gSzET7kOiqxs72TKzWiFG0tKc
DB+wx3N35ZDHULpmIb3lSqoxB8oSiixMsEAHEJ7XlCm+82UFBgglEGUIXe9Eq1qa14ZRo0ac5A4V
v/TxrCLzREhkCYN35KipZo8Ep2bQeCBLcr5nI3Mdd6R6njBG0j1EAn76Nsgrasv0q0mgebgq+9uF
ZVs+WoU3jNgj0dIcvjB4DFf/p1iZvclAqG6oAjWhtWiJe3fkpmKFh/Ilda3QGfC9C3EeNcj6IgvQ
z2CkcDkjzbsroGfeJo7rbDT741zoPzqG9OAZeIQ/bCMZDEJXecUbSRDRnIroXwFF9ylvCp3uniYP
ov/xKvC5UkEm1BLnMIE8OH49Nq1pJoe/uCUQoL7SVx/QbfQiJp6eef6UnrI4ec+M6KyUY9AuUKAb
ogwDiy6pEjrzo0bwk/1q4obx70XFxmI/diewtP/qQdQ7NIPglDLIIs6Mv83SYH62gpK9PLdeptp9
0QQ3WBRflX4RKm7n19/XuZx8+NAzov8hCHvC24iFgIVFgvwFQNGpd93zUu7OSE7L0nWzT7yC6ujr
7uPrr3ZW9gQsqYFTM9OCIKLqQipSF2XLi0Dq3pFRz3ImPUgp0oLUC8SSnuLFrWDDVCvNALjsX6Pt
iZLFbLXJw8sl5v/A2VI23vImLENERRsAJ0WkIFJtgFMrRgA0Epp8KQjPgQolzTJUoH22ATy1xBri
KnDFon2jWf6KpawxNDG/s3S00s+NDE1Isy9nvzhdti1Ns4Zfo7ut/ETMYRcMMAM511E5WcV1nJGk
WH5yQH3gfw6BrVbgrQJUXY268ahCOu6jyCW4F8iwa6SxyPWq+pvOp9skwhZp1+FpOpS2KxqWCgCC
qgHdLBcADwpWjglVwCPRHJlZSVjWhggOZaAMOuW5nXnyMV3oYf/e88dxgSuIxiJA2KGBrjGceZaa
Z5cRuevIVMKIOy+8IrK4xihUGYf+VDAlNiiRdeCQ0L9pG7xdhYyRdmVQH3DHGNfEEjpziea7rieG
OvPLWZYcv+8fFHXtEPMUNqVx/RWrXvFfv4kMm32M2ENKIwMhptfgEtJZSnawwUT9nIRAIcK6Ex2S
XZC20F10YbO1G2T2zkf7thjFKKe21AcoG43Ae3JVnl89WKW16NO63JMYr6LUrn0sUKpJQvlEl1Hy
ob/oYUrJRSmRqabO7lV5tihk+GnDSvT4ySAJ4/VCBjxa5O7/6erTYL4QT4pLpK17L9Avrrm7Y9e9
25IObSXSMLeJHZluFDeksC+No1j1t6GfFm1f1GOYFM2dAGo+ph6IWBYCTtr3H6S2/zfn0ICiz98k
ncEauRr6YVmXSymVqJn/HtWzdM9/aFnCeGIjEtPgF3whxKaTa1aFwqKsq/AZ0NfVabz/cYUTsKiP
hIbxIg5VBorp7DDDgedRLXzVWd7lfZMNHWRd4VkVek9Hm0R7mFXdtbTyJXjFnCvsXhe9CPeV6lQN
USSvnFyB6vKydW+gx9RT2JKFCfn6XpDWWgFCfU/YWc8A/aiG8ewOKinEwzssoXmUJoI3yMJlwMU5
Yk7AgY+IleWNC6xcrMxmhiss4PEibTUOU+VgMrzu/hMoSq6AhFZ5MKWdtdueCFhPeIXEvF/77Xtk
2BUhHtySWVfgOAbwTVJ7H8FU3AZ8bwrmx5o5/6711KUtOUzMwB38pKmoGnKryFB8F9BX+ZfZTkEY
EUP19VCx9uLeJg4SCJSa3O1uOr20gO7MmFEuEmjw2uClTCHOWCuhgYDv9dV2MnWGg/D3tbVVucEy
12jmc4OzBI7jFEj4zURjGtlt2DN4dufebnEbRqc9RzK3WHvkdpme4nJWsJDdRiw7nFkYgOediEKX
RqCmTLRdYq/s7jximkYBEXHYpbBRq8OQV7Kt0vIUCaS/JTengPexQxcX9M9EdfNsXVj4eDze8j50
3xrjZKdqca198CeQ3MdEpgGEJz6M/A7abkNA3Pgq7EpO4DvvR4Gz/uWjCmH6mTqCNJMR+PSy56fE
I59CBnmZOimVT+oXYulasyE2IaRQCio69EeJteFY2dmJ9f1TZQyaTY+q+mA8xB8VVXlTVlzJM6ID
gGfJgaKqhtVuyH/NLTVvEGFWlK7tyUxfJ7mLw3yHk1Lwt8255BbXZ9XeQ9lVArUAIFkxBQZpPgzj
LRkzkXgFbVf+Laa+f6zeTc62mRlfTwppy8CMB+Sydm2x9iuU/dZ27H0SJn5HwOY7tdEWJirP3Nbb
ouQikOmStVacKyVumog9FMWEkTZs4B1PpqZRKUJbZFEYQC2bEmM4HoPc+MGU7Y+zLBqwZXBc4QHe
4xaRj8hRsDVJWu2y7ofa89EzGLi7vTdKIrwOStGdLE0VfLy3mUhjtMxP/5uRY1HQR2yzji48oqBM
ZLRzZ29khM5551uJ/3uqedZ0tBH48CQr/2sit+T3HnjHlOItKaJHCxWuntBWucOM6MA1w/Cv7u1M
e94VnjKCavOT1Eb7eD3Ar3IvB1oEUM4xKMYRBAt4LVMPUr8kmvxSUrpwL60aLdgZOo1mxOdFSoUc
7rORUiA8wE9a6EatuVJ/xjh0KjU42sKeUvl9t6HfwKFiRvWd2iAVvIPO+mFsae3QMo5UBvnAObiI
4F9BX2yrV2n/Du+5GRUmkxzsF/nrhU3RHybX94RMJgAv9Ui96dvavyjQqF0LNEGEO9AdzCO/JGBr
dVWdmqp7Id9c4PkPx7U4U2YuEa4wN6yrTd/pFayMdlMsIjivkxK5mFMOT74Nm1/6FtojJCXlPPis
2XDnkf+m5aGrHgW0P2i0SMnFN9jSHap5K/rL2QS2bupv7EiSiB1vVRcQMXDFQ7uw7ByGyDZZrLBI
Uhx52rwDzHX0i7RuF2hZDLW4c5XyDs+7UdU6JaM0vXEdsPOv5ao9e+pN9yvVO8yxR2YIogLraLPU
liuc8qtlkp5pOTj53aknvJoajLUd8/BDiMk9ftxEwrrpINljjfZaiMc/lsLIKSlevNU7ye3Lfxnx
SNNPfdzBTmZNDacuy2yOoWWDukAuTAAIyoKVD4IN2wGUjUJqefqRnoTo6NhLZliiXgtFSYMT2yTX
lLjILi4GpiYStNaV3LJKe+uqyNPwSy3ZR3WIOYk7RloGkH5lmGU/UC4Kmk15UF2K9umROwAyjDLl
ghobt43mm2SiVZm7t1H/+a2+e4aVVKZZhtNBsQHRKZ2qZEiYxG61O37AMl80Kfh+5Y+ehv9LJF53
ufoMHQRQCfqWHBfRZD82QDjFROcHPSL3StlGyDT3VDE3MkEvHnFNRaF31FVCgheFYQKxZEpLVyHM
tVzElYrV3Vl6yLQYW5Lvypw9aJm/6VWjj0lKVpxKyKF3OZnjkXoFmzlDeL2rhLL/35iTHPpoHfWF
Qt8rbUhF6XIxU7aKW3K1jpVvyR7TWd6GRRBLRRCe6Eh8rxhjEALt72vG5delyBShvGKHEGUe8rHk
77OPnOoHvGdoaf9rE2UqD2Bylk2hjVACDhkN+Kai2amujg3tip6gv2WIMnmLGh3LwMSZ5+uZxx2r
dFdUdoxBigvVP55743TNccNJxainjCxcqElJI6R9GIFu8MazdFmhxOkfYdxyA3XWLOiBr/pT2yR0
tdI5O6IzrsKbgaRR901RAdAjfE4vg5AqomU5dMgUrDi5O4Sc+nEQ/b9cqMIVywVteBoTCu9kDRhP
lD8pi7RnBgJS7/zRiUwUwNbHX3SsT1W7+bZ5oae5selCJzRAohZw6zJCm2u8HY3zMVl1vcr+Mk/7
e0wWS419jWWutfppyDdrYBovJx80vzl6IUmQDinbe4thpuD/5HC5D7z/Wct2fZttYuVE1cbgYZZF
jW2K6fQj4pZcybOx6vna2hpQdHuANz52zXelfcn/9ghWY0cd0dOMManaag/oNAjGf8SUiYv/xCNu
cVPTQRBOIqrnO4Lp2H/aTUsagrfFKDZ1ap8qV2WJnJj+4zRxNZX7Gp/ycvJMFhZ7hIlUnSwGcKEC
CwuwndsOBEUQtceFkb4FSh7gKotrxN+YmqQPEHzNEjZtfaQb2hAGz2G/BFncsmTGA+9XhnuQGy4c
bvVJsbkKuad0ZuBBqzES1pkMs1e3alD4yMrtHTl8sNWfFYMt/itnDM+6zkrAFS5SL1NlXhWeS6Bx
6Z5HH5tptAsmfjBHY+5/csmTVH0SYOmtf6Gew8qZSbzgSwxiDq2z8Zi0S2/3cm67hK9qLd/2HYuf
uji/Q5OfLcWCng/jqS/s/OZqLKjc22+L07lk/Lw1y0+3mPZ7rro6RTVIaBgDrCAAS3s5g+CdBuT2
yuPx5Mt21zA7fcnK/41J9MK4fWbWxPK7kkj3vQh41wCvUCyRxkMAO9O5sIBY6PG97SKGloceAcON
J5/QfWGnyOl7r6MwCTrOMhvY4X1oXraMbtz7ELtbnIGGDHKAVfAJCT932dOkaYTnehO0arLe4635
G1hENptKJ4ygJraLfe7aXG8+ldCHQQmjscpD8CMpwLJy+qfS0nwJd2dcUU07rB6MbEhjayoDvtW6
YXdc004PxNl8roMxdVtYV3DhDvPjpkpSqcXN2PokvtZ3GFvsZhw7CxFtwFqKfI3XgJPgmTyYZH/p
n5lRf9m7/z20JJVx94Zs4pu2181gnhxLb4/jf9gWGFSQkTZMSpAvyNcjoEdS9WfieXOhgjuUlUWg
ti2HCMj6XLa3e5vn11LrVujbpAXvGBrMhkS2f4X73ZPmJOuoyAQkCNZhXIIfT/qb70qaQTT1HsYd
dmjUVGCtQXT2sDbbO7xGnwUv4RHR54/NBpElyUK3qUK57jSmgcwlgVlcyxOCvhQOs/OYTRG+Rph4
bzwBg+PMX4OZldhCDy42/RcOperUqn0BIqWInXqK7e2XMTX2vSrUMmoTstI2xxABvEayVAAuxusi
vW0NabhVgppUA9zdZccIlKdRxGmmiO/HTJAdDzZQOPBGSkYcKuy8yjL6AqnUuOuATEVSfQ4+hS0o
HDp1HkRooHIoiGSauA0Q3AWVQGsYX4Wxx0HcaQiXdwG6HBkMb5Wu8pIu6WknlbOTwrOU16+PF4mw
yuvXdrgfKi7gQrUeYSMNhS94KWPl0daLo+bRVybEeY4sxJl1e5q7CpKoc74lJUSmj/cNsr0hMdYk
VvSPIwp0WoyQ6orIlU30mzN4i1ARIqwRbDRK0r68RqLX0aB9Y53HAA9+LhOyIEK+rv+5cf+cWIzx
9FKHHEBn4onqO/JtFHyYf08ND6MOoQq85Uiwkn4tSDlnV5h0xEW1XiNJTTpdFwI9LmuOE/6MRKCb
XdzOHuUA1bzXsL5kpOipQpcNpZHQQ7jt270OIIhEZEcjb621kfA/yK4pxP4+55O2G5qvD5zQLH+V
Q4KvDpJbifrANZRxFJg9uimlC176u9281yyTLCtp6MKjnxQ/6r1XjQN66DpEUcLRPmMgFL0NYsXG
MvON9ZPLgFgc00+U7jmx1APIcG2dI6ojRzra8LJ5vq9DWrTasQhkKIlgodg8lWUjAq2sDKHBrH6b
RXJdRvUtNlf9O4yOcoOyKbShdOY5p4IjmbzYR966Rm+l2WapQ2q0J7gDS3IVMCm+D+rgMZDAgGYT
zoWhgoS4gw8xlJrL0+4zlKcwoEgjg8o5fEXrQJvCtEWc6VHhwQSAxXbH9r1M59YPjOKJjJSHQKuW
dfVj/7bR0tp6mvM3fUNgAH6CyJqfYBf/OLtSBNPgsR6L5RzuSMTpf+Rfc7C1i3+boBquTuptVATI
aDuKmofvFlTUfQsuvTTtuV3rsZGOhzLqzz0Lb7wuuut/Pj5/Ul8pC4SbTgwZh6ZnoJDo56239hEE
1DpziSdpvNdFtZqaWnrvc3ED0gIjZcmJUEwmEpFZPLIrRT5wxau8pZ3Pdr6FruhBLQrJXUeK4M67
M4DDR/fOW1tYYsVa+rBUNl03Mh0ngDEdA7Jz3xfxMApvGwdq3sHaYRUzbgmR91YB5UEnA3ySU66y
m9oe5nU1BvIqSm3FnfvlGJ/6NyIs98J8PP2mKiYXvu8dRcBSmAi0BFqmCZf4QF0ZTs11xxsTgTcW
DCVegFxne2ptIrXyfpmzvq1/dWiLlWAwlFLDSdN3fFV6aVQFZ6zpxB4iA2ynF6LFKp2bPPrFkdSt
0qjY4xt1J5VXShg93IutfLICuU1PeRDALmgoyNcKupp35wdqjRptxZW14QDT47rj8ofN5i+/0wnD
c9N6Efp2VpcRZR4d15Np+NffEJKWuH4lP8DAusUgeoxuLMD5Ey3rQOrrD6eG5ksNou29gGoa3zeg
u6qnybiOLnHG3DZWGo5LPdR8Nw054FEWCm6t3z3iBvmnSN6u/SGeMElj3S/1NGwD7E4CThUOrTbI
nnbbFaArE08E6yQGoOj+KApEtKoczTNZcC6uD1ME/4wXFY9jzkt03qq3zFQDGIualNvnWTcGvdze
9BUyxgLT1YgkavM+se8Gc6g027p1DM1DBBHSBFkRjxk/ZkpLoxQBfvnjxBHLBOHRFbbA11Kq1tDG
8TFkXTiScDimHFIRxEriipU1iNX38zP8zeqgN5s8Y+N5git+es+RjivkyXkxO5R5lbj0v2z/I+VW
+gdh0Zq50KxFU1vQcxR8Wuc2YzPrO618bF8mC45oV7pzxTze1sPsUURmXfWZ6zSwOXMRGgFM2x/1
rS9o8xRAS8/ddqbLtZAjKLBRaVE/iNgxZA5eYXW0TJrIifIxdgTMCEgFyOJBMcrTmJMxz3FMoGPu
upjPbTE36RKg2/l3P11BXMskp1hWpxd60fzw3Uz+PRM0mhfkI1fVi4AIoIgarZkfvFLJtobeLuTC
pxOArrQOgOpG705TOGPsdTKIxvZ4Z9j0VZaotF9Vrgg4Z6DAQ6ZUgN09PQ1i2bSpfP6Y7fmmft6F
ttpSGdoDVpijf8UzCEH+WTW+vIwGc8t+iqCoQyRNbn32WwWV1puHXr9nY7juFpHWOFCDWLLq1Y0m
me8zgC8H7VrXZ8GqESNrRWNGdGoQcc1ySBbUKlsbjkoUuhWfTnkPXkzekKQnVhH/NXip+huH35F1
s10eKIRIXK/C58huqTEAwvR+grsYbM28offty5hQGO93iu9b5Poqj5u8yXgriMmsW1vk9VF7Emgm
m2O/RjOFUxDwaH1MFSzuG6Z/hjlEGr3t0xgBPgzxxdJRAtLQW9JQ7nJdKIKkfy3s8VOCC1Qz5xuk
ptBpr1lH4HTESC7KeSsllsYX9Orxev62ZIhg0E4wd7liansU9hg6ABmbqpfDr0eDRVS97beoW0ak
RSl/1D1NpjutDS3QgVO4V+9oR+/FHkCsSsjKpPFUhNgzvDS7jzpii8V5LWhjnxWcFzWPbsYizHO/
A6a+2JOO6qihnMpEUGz3/jdy3J1XKr7QihN1FvU0PEViihCHPP68N4u/+OmO/RzgUfO3vjJONq1t
JsmvC2pOYu53AQKM/3FaKCxBEdqxPnjsil7s0WvPmlV0v5L5AuiKSiTomLRYEfuDSIspviuMLYET
SgHZh91EpyKigYKIKuu/AftIe7Qiazw3M+H9hhuhLqZySJGs4yhosLyyywU8DR6R2qXvK+TdPlRc
dDJLsDcD6i2NsM6vqbolAh5MUU7AivzXYA2SQxEXZTJm/bcHzHGrEvnVabSDIjtyRB3BTXeDM7Ur
VnSR8Haq60gKqx/+ssbdgmJ34U/Wz+xbqLYgG9dSGxJIA4xtYYJdC1xgpqgiknyXmo/QDTg8MVNp
Vo2gsTkPPRBhCFQd6qSt0BHIR2XVIrxd4yrdjlW/T84w+t3F8e0VueGwk9CddplhvHIaARlFoSv4
aKFTeHA8k8XkOO3cJkEA6zR0fBnGk2FB0tInXt+H/BfQGNx+2tPiVeYp/i9RVOSWJeeD8Fu0HpmB
BW7koMBx/6i2/upqfOoh4Dbsu5rAGtzGWyMxRO7fDj+0jiH0XQX51x0GMWUJ3SqZe5+nOsOF0sYk
itvRMvLZtT8luTCA8X2TfCTpU4B5WqS1vKlDIoXyN3U4iMsEVr5d8udFwrxO2GUyaWsE1Zdxacww
27IyRVRB/4ezoq/NunT6XptDivEX3N3mXLthT8rRE3Z+pPVn1E29CKeOqPwjas/0z9JBCI2XKiYA
yRQkymon0SQD2BMgTADdBB/Re47M3243vB35ZXECodsocPCS85NTAhDLrNEkAFUj/o6Wa7PrfMix
kF7zjr04o69yU1c3pK29w120AsmbsgGD2x07fbdj0w5n1hxa2XlOwOPJv6zguYMN/xx39JbZX4bS
A7CO5+SnpgLt6CAXeO149vFyxwYQ84GJphbr0Yj9dWFsZ8SwxUUxfC93+uGsHFp//rW/9rIOlNHN
PEyrOB3x93GnuHsOPGnWn4HYvdaryZs4QWGxHaToaw3aFy4KOyu6K+8Nmb10zHcDBPYkT7BcaY48
qYLsfdtXDa8l4XfVHC1ozXmXCL5R/mvvO8YNuU+xGoZSedxe8Dn3yE16UnaorZI4HdSIODXsgD7b
c/OJYkanYueBKUNBgqHw6XWh+rABoiHWpyDSabUmvebQ1TprIW13Hwwn5JKX+hDVnekverp8g67U
RqDJWui41MVcrIy8wb+kh49/goYrn24Z+vkqxRUb4U0GC/TvcK5+lhb0ZxwGHg6HTLkgS+Kp17+b
fE7MMLvZ6qiEY0UpiJfYdMdXTgy33FXH9eF7ijZnlOhsEZWHyV5lxVgJLWZHiu2PPvjOYjFZll0s
4ht6gdVCv+PGJBc8WeMKBDVreI7png4pBcu0rTEAmSRcxNDcouOq65pmZeAc6YgSaohFrHnXRDHY
Ds5P2+D4cyXkap5dlfbhqR+2PdQA+7qNTxXiY7h5vxvD4IVxg8oD3/G2uWdRYRYphlitM63coZE8
buLCqwr0RGKrqiY3IRFZQCTGkEuim0eY4BuTX6GEdzoWGFmmHY2laHlnrgOWcoTfz+nh36ir2QMe
G1dX7dsqe7sqt4NYtXalSofjqFT4LBpDjelh5H2yBZV3HsbvoMApy4U2pDt8woi86HBtbUXS9r5J
4cXxAQZzpCJYOjTl24m5Pqh64iUOqPEtr4sasHzyGCBCBpB6HyAQ/cAPhWgcZhmgncq0fCIMy5w/
weU4ActDmOQEi55E7qi3grWqjHKkx1MsW4QruZNg1wvTOJOTElLIAaU7YmPSlIhKx/AnIA8z5FhY
IoTF3n+f1EAFkUTbrEDGtCSljfJLAmvwbphqPjFeSzd5UxvnB5bYbQhY9ROH08dbSIhiDQoHuV+U
XmKsNTOYdlW+3LFPtZrsMklNlODPx8icR/00U+ynzG+XJP4q8YqtZzRN+hbfPK3zYDTWb9kUywVo
odLgC8vyNfrEfZC4IcGOyZx7NNWwvQlulAQNZaKMCXaD4VtA2Y4YKDha1caGfQfAfCu37e3dX/bq
wQOuSM08tnoaPhZ6VMnHyBeLr8P7V/jXdK7D2XZW/XfGaBHrAe3/V+kCbmYEAuafpDZZtTJeRwQp
yZFHisC7a37gQaDauv5KIddYd1cdeGUtrMiAng/9Pu0Ml6Exl4yrqKTVzQmEVNFinVS0o1qZ3UID
Y84oGt8OHNarsRDEI4E9VTnpuJOP5unYb9cTR6IlKDPmFBNGAK+3hrXv+zw+5x1i/gbVMeFncUPV
FT3xD7zuC/zmX0eno/Wg1px8S1UPBhbU/LbBQuZR26yg5KW1aWABKU8iObXFkXPoIyRRA221+l5C
AVnhYmL2OHdWlx6yAwIz9wvFZ2t3oeQir8GL6xqHlhQB9rLjlQMq3eiUya8Bcyn1oLMY/4xvpIih
5VUAWBNpATgMW8pKTugDidhe27Lpm5ZWU/bClhyz1NYsu7lvZsoR9qn8GZPYHswj94IhPAcaSOak
NcJa/fLJXT0PJuekfSe9Tosc3W5k6CnLucGev/glQV085UCg9uIXUTbdGBZXNm3WLyvQTFvoKzzH
ZvvH/Zl1GINitkTcffRnB9AuWg59ps84xsR+552+/zxWQItLt+NVsiI1Ea/PETCtD8ucRcgQrJGU
gDhqB1AicIgxAreCsrmSIbF78/OsUhTZLkWjdtONTc3PVxrHIr/YAKtFQybQi2VkxBoTFK4jYh1Z
pbz0U4/d67yIUN7OPTOq+SvvclNmdCwa+R0tb9B0ClkzKY1eP6Y7W2z3eVTBlW56JXXabg9Fhs2s
2UgX388GsNcjsC4krcc0+O8W+SGoKCkvJnCOmsfl5CwmPVxgyGgsnZkoWOtVD08+iMC/XVlqY3mQ
ORTIPkSyxkb8X16AWHhCy3HHE5Mp6BZV2oEM2TS+ODGUMVxUibZA0kU/BGk7c9PNGM+afXsdjhi6
ZwR8Qp9jTDB7cDh9ewK7iIUzcKXuNRbXo33+oy8NX8d6MQbUYyl0SO5fsm7gnYB9e/Gw2NyHZuNE
0CZ/jElnwoE35Rpn5Li4CCAbAV5Q/H8/BeCJhhsZNlwWO3A0vYEtLUO7Hc3/LEUbC7vPvCZC6ux8
DyWKRSTdA2CSyIvPGkPQv4gG7+lqwPDf3AEJqRp7RggfcrXpy/5OEio2WR18czgM1yLOGX4y5nU9
kU0bN7HiyUPIt+0Bl4+U8TGEUsu8FNXoHxVlUrVwbZnQLfnvs2Fw0swdXRZrgoicDsEJM4bhWwZt
3XQARmtYuACdOQLkeWYs5ZjhKuHdqWBoCmjRSOg3p7g/BU/Pu3yYp6sGOztpHJZIxDg2gC2lIzbH
Syw5uueoypQ2t7ae2O1F0Of0Y0Rni72W6r79cnXBEI44Jq4p33E/7DpRUFVhPzguw4ijMP77YMZk
g1FrzJNyKWWFfz9ozBM1ndgBGbTzDSJE84CBBU2H5Z2z0Iw+Dt0QojTY2fvWB6yc4MtlwexOjXlJ
DXsWhuPLx9Cq0I1Vh8KEb28rczxi5IV3NvBmQ923MrEUWNMCmq/Gl6d/37ZDd4T2hvPAIiO0tRdb
HHiuEBTKiLpJGuaHZkY0dEWdO2wc0KrF5oPH99jv0J4LHzmkD/Mc+vxjwSW0WioB+XOK2SRFsZFj
g/eC01xGMWY7pwkqvxfNhnRkMvmH7ibmbiHEXKJC7qjU8tjVz9U/mLDu0B8TRxOOxhS/3tmIRosQ
vtIA+/YsHBP9qFxfdnVRb8WzxgDvEqB1qYU2kwmHhT8C4PMdDETUErqGXd5ECwF1E2Iy77lpH7xn
yTqiNSzNoALb4Kg5SZWI30TEqEFYbVPSmeq18OzZrY2DhsvFvAiCvy+FECM4bXITCJd8VR6drg7W
N7IjotQHg5W321QhJcv+UOsaHM6WHEX83Tqt1QEBjajfBz05929qFlgjhxf/eh8VCoBSy/cwDRC+
CVR1SZsyX78fxIpEvhAdUBrh0iOHattGMPa3/i25wh1CW9QfvNlRWF/emzNV18kbRlimyn3APKy4
JYDaukhUAYRVWrCf3AsSmPta62aJ0SQ1Oj16GED6hrhFtb5pNqRyY32/ySyaYnFEhf3jCB3HnNCW
hQNUZUDT1uemTY7AekVTHmObS0/OnbQHxlsBxAYbGXdOZAWCvICkYzWO4CfSdziG3RdaRi2J4/nL
Lq/Fv4pT/O6OW4DdYlka1a1FYcmI6MbVKlGh7M1NV6Kobm5fOGlAHfVyd+O73UBB0ZYR1/Tw3Ffn
tLyL2R5v8uQgdzUG33PIUxMmtE07/1p27Cmdx+Ay9wHp8uIhfbOPI9nIp4JaU7VTNShzvDaMjj3J
1rrQht2v55FFtaQp/VG9FIfxaEETK6N5KKr8+3m2rgPmGMpVdlf8Ma0Pu029Xyo+xpQEDNuYi5+2
PjqZimA1gXyZtRXKzVvuBk/yszMZM0djcUNdd+IPFHY+yG496yqVafkaQCKBrgyyrLHiPl3SA/Rn
XyDjNXu939/S0tsFeGwj5Brg3NOFXf+Ebw2V4ZzzD0cP+j1LLY1Q20ON+evcbl/L+sn14uLBFBWe
meTj31wUqf6q7plJhDWj0Op+IlOgbSg5iTEQPR56bkC1AYf5nUrBWRdyt4ewgDjBJoWyAjC32rLx
gk+WyDJoGvlcNgeOkk/ezyPCAv+Xl63aqQIQL4kjpNAYgI2rhFrm3mFoW6r7JUcmPLesTBz2JQXP
9KF8b0AJs0pz73EZZNLSh5wD91VPA1EcTjMMURWaAcZAb2/dq2XYKtV06US9I6iya3rdUxT9I3rb
uLEg1+MylmDtZzaNvUh6MLyJesV8aRPO4duPGajJG60JTsYxd78UwAXxcOe8vAhmsxcYIEZHp4aR
PZXlcYSUWc+sHFTr0ckJou5XzyFyMaM1U/tIlaEo//wOs7TZw3ROBZk59dl+pw8R25GZBXxxHqFV
Qwg+Wvq/DFHJfCYVMryLwAEYwdB3DfK3p5cJpu9Lzh/z9+iY3+Ki8fbERYYRTtYVw5c1gwqRNrhf
L81LJC/HxJC0J9svUSNOiYlqbRJOS0b/b3Gbbc6ovUxRpUy7r+7LQ/LGQI3jJ1A4s8ywitnI+IU5
0k882dgVTNBQOd4GXZh+AdVt+vHfOYs5rgsv1HBQihjb1QmXEs1Li/USt3Es0dE6kKasB6njv7/m
cKmVj0s+iQX9CpbOVIAeOop2RLUMECuaJNaoMD6nIM5+b9eXfCscG7WgLoN0eocFtsXSTTMJAdL+
5Bn+eTeY3Iqj/FN3/zWDS3gZTbBPM1GU9aCw2w5avxWRDr8pP8YgmwCK1/xuT95PljiADPWeqxc0
WYZBFa6TDeUNzOHtpfO4KpsyjPMIG8BQts1L4TlquvCptjPGGFZneoFFbLgxsbvyUm6uXA9CU+Uc
2uGhz03okS3PFo8NAYCHh/OjrkjoOJSvu3SA2hBcYfL4zviX2zkaBRqKBjLxK/omaBPRDwNJzmwl
K3gX+bWqAM1roUUHABoRWEo4LbDrUBSGyqzTf0WqXzK+uEHErxzMYpf3xPVC0BptOr/AnkNX9oci
J6Lx21xMnV0dTgxhO7+bHobzGvbLIRmFHzRADV0FmkmgBofZvqzivmnDcD0exP1EMyABt7hWkF1T
6a5Fb+Zg6RNKAlFw4EyqdxU5ndoJWxVBQF1zObr9HljjhASDrR3e/RUGmNB+R/LeTDSEC3xWfp+H
40XJvriWAPvEV6bsOEr/lRCDJQSEu+SHwYZYnsRo2PGIGoSoExJkFuQLwo5Hk+/JnbUHPB5zGWNd
gv2dLoCk9PSnp8k98pbjgGhVjtID8e99IAUBEdFjucERIMizJF9YYNCtUTRWbX7/60JOXngPxG8X
AG75GBNcn6VSl5B5+ORZUl2uteS9Y/7H2XdJ4c15WPpsLHTRcsDUyvgm5Cx0ULApzopVxS2f2j3T
oee8z0aDBDevDkW0KExCJ7bOSDfiWV8x+PP1rO3VQF0tAHzrfbQDRZk5RrZtB59Tb9eHz98z7ocj
svfsNTqYzIwaPj91wIxz3050MGHIAe63vfY2CO1+rimYzMnarwkamhC2tt5BWOHs/Ipc1W09VDTE
xAv/LflwEC+7ltTbJt5/Hlb+yS9/Ao9VQg6pDNbKLvyNUtFnSiTzD/oroJZnGqM0uP4hwWbO4abF
zjMsUxJmOBMOYYuW8mFi1lCCDr9YpbNQ+wWngdpL1kzt6wBcuoRBMrninzU+u7EVTB++JtdtE9t6
Rl+1IZ/XdHEjcK8vCGPL3iJipAn2t6E98WnlWiLs/JggYmvaxrB4+kMIjwAXsFYPDW2j84Ktlvib
FOzAHFRNHzO/x+3EM+UFwX3AwCNsvA3rTDdHQxb/+Kfu6WbpYsqZFrrwVHj0FnTOw6ZjEmkDjdJ6
cMOupNXI0hGbeXD65TXu64EnfEtUT9eiXPatEnOu1ZfewUneoVGjDVAQQZDkk0yvIeNna0DtxqaA
CYmbuFi3UNxGixBCG7oXOCy4m6U83TlC77cHnjYVSFGWMqzXwOW3YH11OTk8DmknJkkEV2yP7X3Z
RYvAcxwl81/sVdqPGipN8hJ8W/R5YmGXxnOJQfSLPaHRQoDkCuA5C77HCZWDJtNPvw+dBWx9ewNe
xWytGz/HOGJLenyfAJ6PXFwHVIDmnxn/R+nPYijVqd+VWZaCefaJkawx3w/gfYvpK7Vw2fVnSuxC
EFaUGjLYcbETy9ILd5Qzrk8MdrJM3BQN7uJNVrMCCPMemytXZImGVSfNVnfR+yqiA5HB7WIYoPCi
HWgoxZNUGFVKj0TtDg6ssiFyhB9JNLvMXBM48qGP5hArQd9Am4LCCwb4evpditqYyXBsFzTmEBXs
Mgj31RzVau/MjHzRDm12GuTGfjsyy5gzyCP7UKpNLfybR1nZYHUZvl0sDqBmA4zZRVgPhrjQAgkm
IWIqm/i5Qz5WOIV+SWmHA1+yGZL7hbXBnx5bNAp/BTfWrO43cMTJG1Rj5cMqN4lklU1ykTQQ+flc
TJIegPhNz8Y+eLJoS07a1/x8jd6j6nVmxKhzW0hpRlhlKUF1naFU2EmNFtT/0bnSYdrnzb6PDtaF
f4zgKqGeqxfFRtnynmgdRsbQWSumaFh78bGAan8YYbp3jIcGkDFdG5N9ToNl1PjwiNyEm7cA8AJ0
jvU8Le3R77ZKgLFtpF+aJ/cxxrlED96bi/vbwCQ6Y4wu2Pt87uGFKzBM5sBJYN+8uk/K2Jcnb2Xd
18HXGemsNkKUR22axkvXD6tZLwtuYEsA7AhL3fDAXkOdB0XK4/zkAtNJz/TNc24F5DBqYFF605DJ
P2zLJJMXGRbzsFhAcBjC3kSnGgZYt+UG/SAfva4SC76Pus7Ce81+y7yjCCg0dOe0bc3z4VTiZ4X5
H5CXopfVxNbCeOlXR5USeGQydC/IJoi1nSmfhuunXUI6ewM8cR311Cz8+mjibW5XVLIIMYK6XFIm
NXvxdyKuCRItrgO6lJXfZXZgWuNqXfRKCZPvyXXtwjhS7ShSSFcFB4OTzVGjXV3mkLiLnue0CwN2
gaZAFbb+kPsyAow6MSC03Oq9vyZnJ2qVddKt+YmJXWNudUZPMt4TtlRmAZQ8Tv5mrryVwIRwnwvr
VobrqeGd/IjQAdeHoIKBXqoUJvgFU9TPx+qae0MeZNBX1imSQmq0qsAeLdKYJH9S8UX8u5988/8b
HAnGZGb2q5g9gv8hRpybvFxKbK1UofHGDGzgYlqwlDwnyM0k/FiAhc1/K4h2V3xBZvfTDjGPlW5M
raaaYT3e2yVANhF7pCuDpuVlspMqwtyrG70UIQ6i3Pnx+WMq20RHnaLGgWE84GfEmVc8fAl/uhZA
31V5Gdubd7Bu6mk21//5OSsZwtcgOB8V1pqElH6pATtI3BeR39CBVvH2SMCc8YaX5c5cMK5SBvRG
EQu8WNgvYHmRvwoHzpsMFSQF6Qy+Mqv1XjWOiPLiKmF/J2K2XjzDE0XJaxpolkpcVjzw+R/RU6rq
1mZ//a8YtYQ42kWWDvowvmwXnOUphBmMNYDjqtiTyjdlom/OeqEHH9wbD4XKLTtAs+XoDZde7nx1
GvsmYGEHOCsqgfzpiw2IfkqzzCWymzRpijrTYdS3XJcCXZnZ4r6XSw1i+z9Sl9gcMrYSXwmhLQ+U
wL9IysKUztj+bs5EKZRp6mBs1aPp3D8vjlnbNcdMN1mFoj2FJztdKLDRdh/LmkIaGQ+xKbYBcHKa
O1E5B3KUUJvxMEnKB1XXyVa3Kvr/wJpjQ9uGASkRyaeHEJdU4TOHzZeur1fPcYMU4oEVU8GVtf1K
oaG/29KqclhRgL46bOFX3ZvjSv/UWNmrdiNNcziX3OqiCkOhgnXJvlZvbigX6ljExRbJMDbFIDIG
qoTPGKvZcrhE+g4YUhasazBBsVFVPAX3Gk9iAmPgChROQ374Myl//BN0A9UWrvcs6LsGyGdlgKzy
V4cyUuIPC/GeaPQhgZ5Gf67vmAxFkwhQ6Izyhy4Lc2dlPoilABzegXgSvSl/BG0hNM7aWKuzNAgB
y4qD7YBI8QjTuteaApqW/sqLXC6Wz07koT1gz2C8Pu3WfthpL0qyF1aVOeEz/GHppey8+qReDDxL
L9UDv+fexEnjslOR6/hxEpJJS+kqDd/FyDNrhyj7Dr+5ox16j/x8ZHFyG48MvEuCt+YibNHQQyuZ
tQUYVFfzR1KF9d86qTOWbJsgFnwM2iup4TPm34yaVwVpdLmCi7KpRC7CQ8278reEoyhpUA3P8ia3
8iQMOSQCxABIqcDdOlf3xzG+cMlDE4gA+dGt0Z2w/C49gcMagK8+hwhglHMYUUkHF3YZz48HGySh
uD6nv5tNKvHvZFScx05s97oGivuEmLqJ7RMqQdJABQJT+IqH4m/dopTctfTNxjbJLWRBxLqkSWMH
DNXMOtaY7C0c2twZwZq2AVHfK2+xW2s6X668rAOgHi/I5onNJP5rWgd1XmkMsImZ6oTxTkO4mrRu
OW6QwR5DgVJpgZu1HZMbPvPFyS/WykkURX33ksLbv1kfOVbdT+gHmF8snZ6uEeEnJgmlyDFf+XDM
WiwUdfsDB4Mys+V1Ck2r4IFBF5lHBh8NjeX04VpZ7y+Fr9l8XzoHLgj5e9zaGJqZ7CxOJz4I2a8j
gthijbnCxy2HxsM2FLcuXqP4MEjClR6gGQdCbg5VsnLz46kRq0owAEO3DXSVJon0ksOBBx5iAvL3
4Cbu6W8JG8EIgTQiWU0jGfOsiMBgMDtwhrlE1YrpQpIIYs7Hzk9KkCkw43akigGxz2WUEmnzzddk
/4UcfyzOVdGaGIzneGGwp7VS9ziSoUE6erbwEH3nlG90Lj7KCWbqmUVHvEetP6rrG9s8pTIfeTiJ
dQcyMMKHJqa6IqTOsBX5VB5uBRsg7/cXkGxU/k+CfQDPVzUINGngpv3D1dFlhriq9EvuJ6dKPfy3
kC9PSbM+XMzGg/9ueIb0MyHgeN9ya4cLK+EGUL7c+XKOJpHneVPB7AqZrS/s19rDUtUEFzz/ZTVm
06MGAHrt/3SNgp5Sm1p0TlmCzBCe7DksHHPwU1UvTDhQrwPuuITBLj9+0rcJCGuZfLW98imOvOFa
TRfFyZ+EW+AW9UR3Skh8y84JmAp21e6IS9dDuJn0ixm3x8W71EkW3rzzOOQltc3y0mEniDTXj+oZ
VjjuWbxD15hq9WTxV39bYiehbuiwlz/upvy8FQE6A8uiZD11YTy9HnYd/jYVtXUPbVaudMSVHoH7
FHZnHLa/NRJcMpxPmAVKjwb5/TimhrgToVnXNJuyu59WQYbMVzrt0CdWiy6zvQ7eFOzoo563oyVP
Jcwb4WcYfoCywkkrjUTv5rSHO8Q+f4alewteYSt+NZd33O/wBCwXAuRf2FGb+nl0tHkbtxTNBvnf
lZUTlSDV0e0XoM+eY580Yup3zYRXBwNPtraK7jTIikPT7G0b02hfNZs3CDlS0AYpqO+4I4n2KfJK
z/QIHAyQmtboVI2iI0YIHaLFG3SVN3Nub7Rk5cF95YtfMrbDpv9or4j7BOdqN/5KsoLHqgOH5gZl
XBCDsYq3mxZMTeteR499K6zhx2Ir1km2LgcbMaEghR4Yc2Es7eq8jr7a/UhFcs+2mDyyRrzqZQE+
DJEdRGbXpymrsn2uK5QWj8iBNrGGcHNuL97nfeIve8XXQW0F9JlXqa3j19YhC/9Bkf55omaRmtFI
3NUSyN3usN29u/XX+QbXFNzGKSZu3DY/pLhlngPpUVRdVURFTsZEHPnFTp0+tlTXt8tzevZtc3a0
v8FGpdRPs/wNQXEYOqDy/t2wNZU8ZM7Hrz8WYCjz+sUAcaPTZZEtsxKoE8uGNXK0fMyOL8Az7hzN
iJZAlHHY8Mlz24jsLBm8qwYiX9cHqkgBsgFs/6ZwLJ9Lub6Y+liAg+s6F2e3pnDsQnDg8ZDYlhQ0
ZqubIO7lQXDuMgQmL73IkJJyQxFpqSaE9pgoEt9yu6oZ8YMPuC+fGr0LE5HDzid/SbKleDOQPd4B
B9i3w9ijWjUoJUcFEkdXM9pV2vdQ20mU9p5kORKO3TseFWwomGKoZdofS6vH0DWIGYZbYSFsCq5Z
JGw/aEdZZ+oKp3lYTti6gzHX3Eyc+jI4t/jdt2vb0QWCZloYFw1yqJmt3mPI2URkkYLdW5VXZJrW
cT5gdgsNqq/LinDxhxW+VaTcRjKJC8oirXq26carfn9sUj4070V2o82o83TghD3f2HLwQlut1PFw
OHhw88kWS2EY+Y6B5QvuHQVQqIsKyj8R1MZBQxswY2JjfZKUXmP5RgeTsxi/j7X8oJ/TVpVi8HaK
+JirHWjnDZwJ0VpKitBWTnV6MgyCdF99hDian171cKAkcG5i6tTxtOfTRf/3VcwUoswYWNbzP/Ok
J+d5EYYdLYo7Ibq43LiBTvA0ikbrZus0SmRw2zc+NPEn8JX59PZNRizfoZgiGIXMm3gT58DRcXg7
D4QQLFhSRWPD7gZwRrkqaOrMtpF6lU0t0g+Db7ZVUzsVQRoHhWVMczARhPEyuNmBMygFBhaGfpQI
aLPErq5mkUi0eiR740puI1phCL3Nrw5f1aO5vepNOYSq4Sl65HSyPJ303bbkoVErnbP7PW4er3Ox
2OO6QQG1H2om3H5twsSZlEZ+v6sXcqtbqK0cD66/L3atdA/mvXG/4eU5Mkh8bzMsq797IP8p3EK5
MBaJvIwMaedGPbe25Lo4utHE5sZJukp9lZGwMbWLiz7IaUdRvY6Dp8Ur7agewV8/Xfx/E0fYj/4s
Zc1d19RX/KZa9iXj+3f3V0qirbuJzNwC/qcMTZvOyg8cOMW6cF6Crc+fSPOx5EPphGXx1x5L1gNq
s0ObGpX8UrS/2AKGlJMhWRqaxO7mPa5CZjlim9OiVNADMayDAvE9v4Ab1eC8MOnu3D/Bt4Ur2byM
fBtmMb09++i9AtZMdEPKt78Dou1yat53IJHedvvUPgS0KJdhfAekZpr4IxDN1bnNFgFHYWx2KLV7
a579HYGhOwGBMBaW4Z4TlP0tli2Hesz1MRt7R13lQxQb+j+hZaArQCHakwQ4yuWMV/ySzdSwgvpq
jqfCFk4bR5W+Yahjqlo3GA+ETfS+11wab/Xx5eX+qqz5ITt8md3Az5Jf4h1puypplXKUpPaGC7N4
xM7By6XuDJX2u/UzgKtQUVkcmL4JKo6IDJaX2I1bD+eY8e6e0TmcqDufTOjXGuIEARreaggptMoA
Iuh+S5MGKXuXFac5OdRV2zFEZIZQAoOsKFWefBdOyX3smXCg6KyYdFqZe0cShAVdsXlyxLBtAx3e
8bikyQHvB5Q6TnS5XY/d7/pG+cS4zhzqPvI+kq2dhTHetYfCTBvb1KrKvcwgfwDqzr6C5EwRijSh
krubi5pU3T9TeewYB9SaF0YnN7nzSpkUDNDK8LTS9/HH1OYPdprvOro2vUiqQiuBCWUeqtRBKBYz
0hvDcficgX1xLgsL7cXh0RVeGFntaf7DGx3pa1vow6DMO5bf/0jFV4mIprAfUKBROcmiPWtB3THT
quEkFpRZpeAyruYtppSFuvHHEpFpRjLTV6Jzy0xl7gvWaAkN+9jg5zbrtoI5rxoQ+ifmoL8DaFRR
HM594QwkPzvfbh4G92x4/fhknW0ZNpbO+xdvSBtgTLoOM/ee92J7IrBKScx89oF1IHKUwwoCyZKw
fI1Nj2Ihk3Upx6U5d4KVaNTnsKMEqhxfOQ2BQH17JaO2QUnSjYhqYaGPDS6AnYO1Diyi8VF1LO7f
cg6IXrWbcVtXllejTyTh/shPlLYBl73oIhahtv7nimavuhN0BvoFkPm6OK7jUV5SIUuCGw883sfw
JHquni0SZ6o4zLyk0t5E7ffEJj9gh2iQmNPFss1/pwBcke8meF0J/l1l2amRd7p+iy7tSJyS4gbz
aGZKLUOOw4R+qBaQWMBrhYLz4zAMAVlRDrNrNJgkXhG6H5nOJEywVKtf+czRaUfKgWnWDyYB22L+
7G2r1WkV4q6pmtXV1Fp1USH7eolb8zmQqeMj/tsanlVeTaNc/zlF/7GRDF80HDuR+iv/5cil8e1f
H/IikYPZ6GZq/kFxXez2qwWEaEE4NuE2mRq5MFCUUu47c7Mh73O8OUZu+pQobKTCKnyDvQhnayHW
BOe2fFh4s6xeSrMectklv35foQVWZlr5KJxtT26i2PcvQE1UcKYq6ucHlhi6M1k+Wp638CAsgakx
VVnOy1kGDqCl7cMtG48jJe1Rfxlyu+m1Kpw4XB4MwmtzrLu7Y7zZTOuHFMIWjxsIaq6w9MqFhrJD
B/edCBOREEZIu81hZQJMxJmzjqHm4g0Ty284KkVpJrOZATSkocVJh4PmRxPvGSjQNgAvr2pinf8I
Ct2SoJTQAw+6BxX2eUYSuaTzkbCyhluJQHPqiJvi6vh62fC2CqvIlyhxVDQTwTsxTAdveQ7kgWRL
jwnPRpXumk/xBiiZe0otNOH2zsc88oGeR4CoQNthT7Dt+PK3Owh5q/qEQ2qhrD5Y6ATPpJkgoXpc
aCKq0HXJmbHvKub5O7ZdlZQyF7OXMTFgeFUFBkWeDnafz/2JPRoOBJfwJbyJ9hp5uTRpwfH9fzRT
JCs3U0sc5IlvzGh0O5jNW7VhfDWQCLNi1EgGpQDyeTswVId/XbP5sqr/Cy86D7F5wQt3yyi8P10W
DtbJjRFz/OPDie3NE9ZGKqDlCOXQYNgxZv5tLyzLR8fiDIbz64v1Ub7QnqUAvBbFBEBtr2nZqEbE
ShB6Na/hwp7iJRwRzOLafrW0HSxXkcH9Rzx9e92k2ggE08lsfg/WeD6BMqDJFn0ebz1qP+1Lkjev
sXuO1mSkCPWw86sy52NLakKnNCFuZFu5+N8qP5s4xmB4lJiz/jRew+T1EndnCgjP6kxttYIvlDE0
qXSGtWAP4I79R3UUrnNxIp49XgQ8NshaL9h7aZjNFwLrKvQLzD1r/zTxcPi034Gnjw+dL3kj+kh7
ISat+lHe18pdrrTilfqfWARTTTWkuKUL/ZSFoLTgPf9YVpP6n/smoE9MlJmGu9tpcxjO7bHqyEo0
fC1+Xez7tOkKLSeNPswJHmWIpphlwPffd0KiPgKHRy92D/5tlCoAR8De8WfnvXsWICnHaBlCDKvo
46mwBHjcwGgZHsHhaiUnyRzlwRyPD+vl3yWnq2FSHApaMyAuGFBaWc6cEOXuwhLDZ1PtIOANHGC9
/2aglO+CeFDsT9jmS+l+HLun7ii6pY0YYhgOfJG1OHyuyaLZgIFoDzEO1DUnv86s6cXFaHD/KbSY
m8sXsIXhrHJtkyrHr0bJaSET87fHndIbEUODTXVC/hq5U0Oe/KrlefeIywnlJcYEJCa1LjRfax4P
EiYuUyVhYWgm9zr5fPBuXYL3EfGJPB6qO4Y4rm8TEbSZ+UUszrufdfaCtL/zt3fx/WCHGxKG57MD
pcG2yO6D6lMJZIZ71DdOOsH5K8vNZZD0PJzshWBOuGknntftGSHaUABFEpeLAsNr+1FBoZ1bzslD
A/5hECyuAAj+EJjqPVkeyUf0Ydb+ZPbCSOv520WplIXT+CIYX14zCKB0W4/3XGQzyJzMp/ApFeUC
fS0MUUKbc6++4s8n4DXHc8LFLfI4K7glfrqmOqcOaBE/gIZBy6jdnijWT0/nb/Ac8H8Or5itGiqh
jU/gKGmS+/XQqsSW/uKS4+fhcC5LCJp+QWx+6KthZ6D93IGmmciRwN725mM6sLl7XYil+aokRdoG
ZUpNPjuVPTPN6A9JjlEUjYM7ajPy/1zXjcLxpLSe/EtGBvQslvt7GmpqsdiPcMFkmechvLgc5g/d
cvBm20juw5eQRrXXFbDKTE/p9iLRnKkrLqgLinikt+hayBD1Isq5MpWmEmqY3HauwdKMvu+NCArj
DR5vYym06zAs4dsVQ++lRiZTsQm4VBMmwr6uOYXxu1HMqSUAGq8ePkZ4J/SLVyvd9+3zKGHoK5O/
TD/PNYwBo7CnG1RUl6koCFs6HpQaQduqjK18+JV6/X6QR1uILv00HmD7ns82oXLp22fou/hRRW9U
4wDLEJ0a6LZPnggJBd2cCtsL7PlAUkm/sV4EbLAeZPRLB90HfliP8X5pBHyYI7BoRvG1tYrcSbPf
4mV1hCEp7i7R8ZaBpGVz5s3gWSou5qYftbTjnP+m3ocaXqQkbGknZp/AxiTLiGmTAB6W/8vBlvML
joFNqMCkZHeXHjCtyuKzQ5i29tIGXcOQ+EApD4hoZox5gClKkOI8QRBoBeMKlSFfgPS7AiGS4/0i
KG30HZEcma5KN1kzX/xe2tdOFiTd1LEaColaN8vNbnizKnKKDzepO6GudDQwFvDvRQ00m+mzVpu3
FtCBqb9oZa7PAz+YBEb4yPTqHo4SuxCjVYPz2PbzGaDBiaU/ux9i3Zc7nCbtOus+xNGu01fLCZTk
2+NBfegdyLqLk58XAMxb5oeeAbP6xiokpukQgVjMGk2Neaq1aF1rK68oDlsTp9a9ACTWAgFlZC34
yViI4ZVSZG61Wecrb8OlgqZ7zqpa67zGIQudgKoTPRg9jDsp1ElY24m1wWc6Mx9yMiNbBxwiJ+2I
l8l2J8QYSh5hDHuouf1mhzDL4ciOkivaf1SrZ2QkQlcQhAoMw0arDr5ovElOawnwIzOrIjWH0GAx
AGBjkya3/8KRDiblrwzomvja4VuAJNcxBpLyZk7Nxr4x7VgeVZ0ufhKeOFzaljxA6Fr9wOBCd2q7
tuX0IOl8SnIOrXdScNcVplRKsuEjta1T4546i+1lHzOjpVYl1p4o61QuG7wz+l5Zb1N2DsbGNHZq
fEOVKmxiSFIyp2YBAXHdsOZKTzi1vzJiiOYPkdKSKxu6nyhx/PWpTcfn+06xF5GyGww3YHaW9Zzh
yS4RTEygShN+r9jn0QhCWEt2o8vXIbRxuwa4JJNRXoCwaNrCQPeK+OJZu88KUIX+NZh+9Yo3lqFP
eDzYq5RvzHIxfTGhK/NEG7BFeIiaiMkvtku75LXorXuPRJg2i3Oe9VOQZFbW7f2RiOrc9G6kgvA8
sFiMC2pAeghANL+ofD0Oo4lAQfkmdvIYY8gE9Q0HZuldN/NDov3Jp0sYSZX76r8PchvA10glupEA
hDGd4f9JkMrNNRkN3J7dhXkihA4mfdyZTK0QIqY6yylJefk3UJ7b1v4V8Jclvx4scRhgdVfSiFoK
qMOb3qm8REFfi0sLgiwwXXu2LISY1kEgWJrO0R+e04u3523tJcQyTWmjMTFizKeKc4mKuVx19JQQ
LAiwBdR4v6PKfPmg3JED3C0P908H+0MlsuFXjrWeTgujfVzfecHyyo/b9yRnqdcQV/69eyt7OIwL
gwzbt4SzAnEJOieUg/RWf1lmsrCKzg/dKr7dHan/Ei6fVBnn4LsHOo5tCf4m72w2wlcyZf4SzF+n
ja409fc0Ddv27PGoO53CL72orB9yP5WotkxSwvsa7uNxpZW0JqQcUzlPtZaYAvbb4isJhsy1ssTr
SbSv4cXcwXO+DnznYJv0hM3T/Z8+M1ZXRzTnD8rAa4+6vjKsNcI9EDPf0uY9UckCtdB8CgU8S1bT
Jnq8s0DmkJGj/4pt1DdiYxb3ioRp2v2ppMNu3H56vIUYKKdH/69zc3psU/zC3gOLCV8CELFBdI9x
rM/0VBGJlpEAnwPOLOwl7XNEjd7Zn2n4NwRnw7jxwakDQ237Z7BHCl6BS5wDETy0BM6yN/OIddAN
Q14xDvD1om1JWpFJaQro1DIdYfZm4obOy6PO3tf7dp1VsP32ggVsaK2YOATY41JIRdETd9E7lLIZ
oR/XGSwe11Il4wtmj6iSTtwUAUXrS/OgiledTE9yrDkApvEopH9Z/UzYXPUScHGSsQm6EGwtuiN5
PNi6EqMPPNqJYSBXhzhLoszKYMp2fqncS/RslXBGCVn277/aF2cxarCcRereYyR9xwyGQHlzWpnD
F9vJGloR9e4+E6ViIktHYw/uqadz6evi0llY6l8E+imcxxf0ngMCTLN55HYPEb+eHu5RZcQPBPfh
nHgwMNnCqVmNyiQrcmimy8tBvqX3lqHwbFhyrZepZ/gnxauVkEkew6rAxeqPHBhNJPRW1TNO1ngk
AWts1tkr6qytQ5mLg8J0ehEpHUm1jeAqKRvBOuSDUel6+7yLGNpUYpdpTPq/RXhACfHxTaP2euNo
MNg3gZOBorQ1SU1mhy655WA+ocYceyuS8biWNiQvFJeFS6Rsw5HT9y+BSueZISwvhqJYw87odq17
+pog4Ezyd7s3ZkW2u4zzjI0Afca8oPPTFT6pBpQ7QRsTBZ2ON1uhMKpMsjux1bNG9F0xP0DrYb+7
KnH+Or2+nUlHPS8Fnc8RsjHeTbH3+Au93rt86Xqc4vWcbmGEh/FL9JkxCfjDVuN6rtkHnawveVGE
7bW8eXGloBlP/JBCJ31UW2ZQlJNSl5unVSwNQ62vUYGrTQH4+pgreUTs3Xm8k2tEGfjcqM8zsbE3
BAhn58xhYBFgWN/dTogS2+VY49x/ofJDta1Qvq2sYkgfA0aSiwTpUF/Jem8MKC4uFG+dRggFTKCb
iDhgr5FxcTGb1eMcOjZhfHUKkh2F4hKACjTlRnI8An22Yp6K6SKItCzYAHZcYloimag/RkSmUCez
xDxv4nx1UgaNiEkjRVSfkXrezuis/Lo3xNhGIh3JrRA6uyyXm+0oqCooEXadWHCg1iUXiVoxmC+v
CXjyhtHsxjg1R2++P4bA7SdzEMJmdYlITRRBWjPJo5/4gz6vEQccC4ViP4VtPKu99krasHJOx07p
AtyPyg6jbX2T0rEaYiwt2/npwa9MuUv9BmIjUYq1NuyoG5WvN8USleXZHcMigsrTH0qoP4uq29gy
6R7yHsGWIcYw3QShAijyoiCUIw/Id4l11aBsScU67hsw/DrhloY67qLYi6tgpJAi5keOpkxEvwV+
RWYQY3CRY5jMB5FSKTrDfoBgVDM+b/nGwMeiDxnS2BwN08LfLQgN0oWjezej4nMkzUoJ3vxzsXlx
xvHsO9pmWT38cJdpBg4rqn6IvJUbPsNBK80y+d3w7eBgnpXMZjQrdjHZpI7EVoJWnE+jor4xREL/
Ny0/R65DOeeb3+rSY7nC5jddlcLLvvcKWZfcHEUiPp/+SB4+ZUTu3LWzMcyVsvumwql1taJQs2a4
X59MvuwG7r5KtL0RG7bViLsESoR8uyjbPhv8cwhOxmGHx4AIdg1Bq/GKhHnyR3rSJ++dMsxZVFFD
InzcZqRDTBBVYNf4klDss6q9BlyZD4fyGpyGjeL9UKKgo2X2zhUhW/MPq2+74O4cCfr/61e3Xlrs
diV0bLKBnCMxKSuxdlC01YlHSZ3AbquWR0Iw2lm9Rd3K4lsiR7/IRR/2n0QbLFTNulkxioUGagWO
e7Uf7/6tLceDsRwYHsTlda7nsuyZrRzEEw713gO4GgGRWPDfA54O7CO/z+WXtMHWDXTArg4hIx8T
KL071QpxOQ+XQZtUruHMJz4ZtLU4xSKxh9r1h1o6dGNX3p6JcjQwWnAlD+dsDDQ0ikfkAsoEERhY
udY2KrkSrglknykahebmTrzASrvzAM4XrU01sBSiLxrKroF4+ox3A5kvpBoAt4xsIXLg9ZpK5pP0
yfWATsgQ/6SN2D5jEEAq2CiBVey0gxdTokU/9M1I2BKixP9bP2UJBv6vfAarVWjBtcZgBxmj/WW2
izk/AbU3I4XvSSvm6UZrdvmlNSB5xmrQsA5d2myZFdeslUurNdR6OMgRExSe0TIK1pDnjgtk2hqJ
GQTcKsmTc24pjCbuJu8DEfrXkqnZx/BSS6H+OAZBhPzzLwiAuZ9exroHozNNCcC+wjBWdSGugxOw
NpdBGO3txdF/5WZ8rY6+1buENPej6sZHFepAM5aScsq5n+VdYXxsXxdE7Z4m4x2EJOiufIVPUxvv
yszCHlPvIIYbZjfIsKAAtwYh/58pbNZUbGCcHMPNA02hqvkPwAfgNhfQl711SuPJN9wseYI2wq39
qRejCUGlhEuUM81j0dVpGDIeU3Q2sXt+ldNYvpTe8GbJdhRbnVoQrXolW2qtgTsZqtW5XAerp5Ck
bZ+p8sLR3VhmWHaTeRNPxH/gjQKuTS/JcMwoXb74tg6JoXRvjRQ+v+XO9ylfDjQov3jYkj0x8BHR
Es95AI0PzC9KhMcEaxhf9vSarr9bLKhKqmSTYKWJmHXltiNHZSeDrrRsHD8+oe3Gg8QKZzptA9yR
OM/TZ4ZDosK2evyz4uX6HLo0259f6uE0x+YBZKkS1xkBDsE60Tn9N/ClEiIweJ6eTNAq1BmuPBCY
TanZBpirs7gC9FWrqvfI/NB9+f66T827ZgWh07GhFOHn14qNitLHSbnaW5og+D6YaUveblIfLLU+
LZDZhNehgsOijVTNzNrIu1jvr3ZuN9XPD6mNHKrUQqizD1JVkqNNPfLje8Nvzi4D8DqhygmTvJ/q
GGzCapV+gNi4Ag6J4FXyscre1PvwG4ghoQqdFC9OvNa/pX5PjpxQcVSYx2LuGvgfi5CaolmrcvWI
LoVRWI3MlpZ1bZapdbiQPwWMDiVLHlF6YOXgp3C5P60dCX8CtV+eZk3ggJj5F6zTCDaXgd2UH8rT
W8sQMCUHzzHAgYPrsb2tvjtMjc5LEeGRX838EbPUa4u3hqros+z32jqKmueNFqZ71gmZhz3V3b9O
pjXFpA848saZxVqiKSQIs5aFSP1gxiPjLnjC0/N4+9DSm4CWyVJgjvZ33wjYDLltgw2mOv3/vfj4
S6QmVjQXKkzN4zMG75F339FzI74guf/CW8lJ6vw4A3LgEC1SsxqgoVyKCZvT4knfJguyPSCP0nXs
Ynp/B+wMKc4m2HVIA+WghE2ebenA2GFsv492Xs5Ywx6IYSoN/NcslP3+c6y497oDiwF4jnSbQv+X
5lYc4Smq3WF1/etVDQZV1wuuFOjJTFdX3leljnQ7flqUSqd+LYkFTOuxfe0I/f22ySXxZ5MhJII2
t1fe+YCXFZUxo1KnMIxUq2bM7GDWWGgmtZnn6nGE4HZ/gD2V7yqD3cnPN2L1dNdScGwC9yy0XE3T
omm8gOZe8OR/EJnfrE2sjwX6s9jnLNgyts9q5SLBm2/A4t16D5YN1m5xQRClTaElkv3wuQHB8FeH
L959vLvF86zLckFzWblU+ihlPbkMwFs/cfwTl3d+W8XXtOn0gmJXwLyCEHUUnSW2fRc7VRQAZ0OI
82rGKHRuX9Zda32BwmQaqXNzjS5doBV0AFWeiSCMop1TgCvO5CMAngKrlyGT05XKOoXoV8pDY1JO
8Qf7JHZchdLa+k/U2ASZALnpckvfirx0/OVCkHit2MEkxQvOe6KhngJL9mCd16H4+Itxy0GRNaY2
8mMZowHMD/wITmSDZeQXSVH/mKvoIuuiXw1veDPv1PS9MYjltWQKHcBpZaLWCg11W9HacLiYzOtw
70e3ESXg6vJWuwRYValpKrD4GopgsIX+dzeABvDkvmFHAVVSPm9SJJlbMBsdJx6A4rOy3l34oRvX
d/zDd4U8gD9j/UVMklzmBqYVxi+ENoMYNDDFPDXaY7ppqZUcSDr60mdNEbkVlKBYvtn5FIGNwXUb
X+Ita3qZqQttUrqoXIcrCdTk5D7DbZ0EIB3WvHGOAxKwwLX2ph2gtdcJVdC/L91dMaOYCxxhyxPY
6GSc/Toaqi7gu5qpwwussIZey3Fge+iEWo+H1msZgqAYn+IjY0n9LuNq0Uo57E+Lvtrdaahg5DNl
jUhLxmy7DKh/TZovTxA+WgfyVPK3L5LZcb5xpXHrf/WKRWaf9fmVBXSbG8zpIxYS/qkGXqXPs4p1
kS+0ekPo33pGk9mvZHAchwqh/lTm/luR5TPFlKJT0tNY/fByyG6Ep000PZ2ZycLhiO1QcU7OoOGl
HXP6DYxmx0L9NoZKuIlAtQbfTQYajbCjTVl91YbmBMGnOhOiCJOvyXPAuR3BSVnqULUk4V7rofxF
fKLat8VJFsu6G6vi/A9D9Od/9mzHdTrIZVr1hENPBn4tqoY7LRWu30VcbXCiCcX1h8uq6Si2Gu8X
A0dTqfBmRjRWIdewMQgZL0SopP2t55VOj4So5UgFLN5D3IKzPOMnmcmfkx/zB7Ys0A+j2d4S61mQ
+CyXZt/pCudF3b7NSCjiLdNoubkAUJQmGDNuFep4ydVdUAU4SDhieN2q6s0Lm98mp/gC6NQ20Bl/
rznSZxHv9P9br1fUDLq27Q9pnL23UgTzFoAn1z6PaJOrBEpU5Vru0L3gNancF8w0jEVscbe62gF9
lFAPS9Z5CQanfPrqbzw3rjCa8T0DgpvCpk4iw1gmg4G/3w9C1fWLQfETwlLcjhejpwZ0BWpfGhQm
7bPyZ5qqvOiuKaj7A0dpeCaNwz9EPa2ClZSrySo8pBbr8oxp67dKgkzkM5vpBi+dDcoIumhAQEXs
SuBvlnb+sKvHqHm240BgnYz8oFulVGcR2oX4jNPbRx5kwPlphJ24S+vjtt3ZTU8QQfcGx9WeML3Q
KltXTaSSmx4l6Qxn/K9vU3oKxkD5iEjB0nALwrA5a7zLnbtKYI4jM5U9BPlhApmDGOUlj54p+3zv
eAR5gbvBd2xTfz+VwXhqBvLOseOK/wSBKyl6QBxi7TCZYbOSUf/UtDDeUS6xXVHKaT6nYRKfVuZ0
rXUpAbS2+9QhLtWueO+I1toK5XmSOjZW+BRHbKW6yV4HX+yYWdrd7bAFSoFxok2zJA3zM5lnz30+
XROBJuVo7uh4vVT+eoJRYfUnG6BrT6nval/3/xfNjsHDhQcV/wJuHMYsyiyx6Lgn6LYlyMpmbCBs
q3S2Y+cw5Zw862kapuIW+j2qG8IJYdDvwugrj4qQtB0ByrFxPV+y5EBL8k7YLE2VGyVyrL8/eVwc
dh8exzmX+m6Ev2W28bRx5FTOOf16PNDSXJNvACSaEJHH32TdmcYb2SBO2GZ0Q/8rTP0Oo1zwgABS
z1WFfBQOAQT1jgPMUfIR48CpSA5GpA7Dip+cZ40rhyf8MoIqDEH+mlLVUWlToiQcmSdeTWg/b08i
1BtqUmusH6sH6Rogx81Q421laGjALOHCuUYW70pjGzE/terRweB4UAdfQhOtwMfGbiBPeDw9gpmk
WUIoWG07xmciUtbs/mzKNJ4TMQr1NNRLBfAFo/UZTrW6nxOBk1q2RnH05J3A7WoREAEzC+clqpjT
pFYi7gTqhHZhJ9pAaVMhtyrZ7v1hz2pa/XrIpJYB9Vn0D82EhNJEO4bZxBMbqBu9f/qnjg+zPThj
KqGltmUldUkkKuN2+ojhnD391Tp9tTaa+twxiesfKRy7xR3KpSA26s/fFhjbD5Ns6r6bCwXDP5v/
xLjaR0VQrvtidYvXEj3Ocqe2Vm9hHNoU87S/Ut95nlutB6WntTTqrra5+Z+2MRdgwwBDgdkjggNc
rIwwKXC4eEtiTa54GLMrBgQoW9qtdNX23I0vXyJyI2oI+dm6M9C3hnq4rXDE4Yz6X+noJX4ODTHu
gXMdXzolju9HYM2qV2cDyu0gIGLvtveMVSnUwo4tfVsOeBpewByL7GxU96dsxBf+tpyKU0WUhrU0
P3Tmj/Rj9wFai6edVkKLgPIgYemK0d7EKpVI003+fDxu+kC+tL6g0uyj5cQNfb/j3d4TG69iq0n5
wVLd1uQ1G8Y4CW+dExSEXverDBQ/Dzl6PwpQk/eBAzFBoXyrjcDej772luvmkboJmG/3YUKsx4nf
rZNt9Be4g/0cOyIXlCF+DD5EMWIf6JOG/g+dcbmoyH3sRxMiHpY9TB/AVJ1RELzUvwC+vyL+sdVK
ga4ZRb2GBIdCzw51JV7VAI50buqxiUJu/HDuvK1MYbM0RliJnRv6Xvj2bQO+vaIWW9XDQtYEl70N
9eg5NKQANM0Zy1/B83Qu7W58UesXxi6aig5A/l0jdz1oLHx851Gwqd3cfaG06JNiBwWebKqWokjL
FD57/cQmZukCz92YqAF1fNPxJAQSkVaB4G3xVbn+K8Yfd/oSx9kCNh952k0YCF9dRHdbkF83O3bn
jR1Tffw9PekXASx9bcwRSMZtDOjArtW7Mp6OvZUhgTk9McDiGd+w4aUhb8Z3KLc+Sb9JmzF/99lt
PZ7WwmasIqAjdbn2yX8yYnCc2hYnZY3ErZA/ZaI9WjnPDamkmteT+EO7wnAKda/KSkQw/lnSH2L8
6MW0gLsU5K/MkhZpG+1lkeXlITWsUdfObWaaCTnKppc4dNrM+47I7zM9mgaj5p7mx1AU/FzjrNDY
jN4bKsKF3yGZQBoG1nFQanrgqAPso33MXZvC6T5O/noM5kFBAHXDyVtNEcpo8h9Q/PKTsjmNrzR7
xQDHHxqyYcrm1wWNvBTY2IPZnD8150cLrGctQJWY16cAf3oVESvc15DWxE5hl7JcfHJef+DVQC0q
MssGG4SwOgXWPQlzjStJ53IeixJwco3R/+vUqXfVg+AOj+fJ9iwk+qVPOs8nu/WkOulM+jXDvmjV
UTU58xUGKoctM6y5/85rFft9TgzE4s4Yn0PZrmi1eUxlUxutWICl63lkqKuCwzbxsRIZHQkD1flh
pQiyWHeMaaDZoo6E9FM9a1hF/fJxaPMs+s13OnJNxGlcSTj4f7Bfx82vBHq8bM+t5qPXJQUTtu59
yVg487CanvOHpRjIzwQ2IxdoQBg713j6Mopl+2aYGKq3XozBdIkC8uR/aoyJezEEvP4etIa0kETf
85kIDKwp2oDG5z3Gw6+hJ+f8YcPPm0PnC9ZJmAWHLDE1dk8YoAwy9vcZ4eOqp/gHqD2h77qejGU4
xT4XkgXwY1jPjFt59kGUBvFNvMYXY3a4O8hWNHgjk5hW7TVN13g4yEt7ocnCtXvggMBlSH+EicM9
R5tlsPW7Yvs+/LstMalxXOmVzaSEILoqUiaUcfcW9s9XZdNRJW9DCBVAaO3vZe0LwI+6PSIqI0fj
4ebe8F5cJ2Lq9yaMFok97k4RNTaetbLq5T+H4Ak4eJiijUfz46ZViWk+XbjGkIg5e+qIqwbJklXz
1l/ss0RLtSAMbOlvr6pmrGpakUYfZ842nvA7PWQdFIJLfqY6VqDswh9AwCYjtKcXe7GjiJ+8IVmS
oCmgisG9rqQOwTnlV0q/XoDkSfbscAZwJaxQ4kydBBwGlnhh0fvdj5bZk+sScr05hwUexBrGyP7d
VNnVbfRHM0wFvrUdflyJX83Wh9vvsNqKRhysjcZBvahgARgl3riaEVzfHBGkQIB3e8WdBuZHUYv0
ribh31vgVLbBRa66xvmTPXXiqVAV46YEdF1UxTpCZmc0/nkTFfoS7tLnjYHebOYvBVXV+mLvtAgU
/CWmLAJrXhonAI0ERncxodTEVY+wNTBFTvFd+50SgdHb1o7nP2optiJxFDwV2tzuvyIra1hChFkk
XLaw/pvwzxzDEJPDeQd9C5QRnw2hvRIEN75/0NesKwwBSEC9/c/l/Vb6/yrVfv6zd+QcuwZNyMQB
v2rOLcaSiLcx/JEJjdvSbhlgA1Tnrm6exF+6Uc2R6q2pFGctpUi2USg+TYYq7/dcsQTuJS4EI9JL
as5VURsZI9YOJKW36eFRX8GIbQvYJykgQku2Zeffc5eYj9zxLXaR76j71ZSkAlf9kW6rs0+sAQlv
6eTuE/pt3uhTJVBMKUvP0VQisV9LB1hWNQfNntf8T6siHwP679lD0cwp4Il+TXjy6433VqLZPrGP
/+7LXnABiJ+bThEBm8eAlOEBsPOQLKaQ9MzuakDXIpM3DrTd6ZsS8czeAw+pwy9fTd8dmG7fYLpf
X7myOwwfR/HAfdYHBofQ6rOM242VEQyzV5iPWt/9OJbf8PfgfD/sUiedbelavS+QnDgKntzOr81d
8YF2g0f+xyH5WgouNXkvD2TzYCxcQWu1xSb4oJmo0EQnQbE6mfp8jryGsDZKs7x+dpjo1ezKPl7e
9SUNPGvO1SuHrMx1vj9dsXZPZJx+TmXg+o8Iyy5RfbMLFXX5kxKLaSQnQ6QXlYWq2aYXDQedQG3x
L/cL/oKsxw55y8Wcl+va4n109X4mdE72mvHzPizBT+bbFzQpXyDu2ujEqPFc3YsxHfHJVgMJ4M98
Ei5q7oVuUTFL0HUKFFKiNTbQDM14fLGD2Xi1UPtHud3rZlG6UrYepUj54y+5EOMZ7sJCQ+OddEtZ
tsVNHkpJRzQQrZSJQjwMfGfaSg2KoZWHfSRvptOO4AGglO43QEHSJKFlUPfjv4ngaifrWXA8nHLM
3F+RSotvcjqtXTqnGrPN3gM8cHSBu1/fybW3f6Hgf+IGhJWGtkKRvcPsGPqX08WcQDF4dKVj29eB
2XeB3MET4C+6MSI586VA6ueqLiC/dwCZA2ybNpNPILgRMRLOctfbd28ImZzObjp6iGO/fB3H64mu
w5wZCyHv5sQomQebdSmXJFFzAcYRt9mi8ZbEAfvPlO4MXOXJ2XOgOjR0OrWuAtPw6q+liC5KhS1R
LXZ51BeiYTno5bh7hE4/JqMPVSvBtXW9DV1pcqAqV9fMJIHH7+w437rWG0sLtejgEtiYj/Jvz8+P
J+PXJi2XOofUBPP1Td4rzrbH8cxoYD5/zCq3bqge2Et9iFnhMR6wP/icE9ukO8YN3phNvf6+tIh2
ksdENgLbDq9k54MoDznMvar2aRiA9CfylTmqdA5NUl07lz31a0Q/dK0uqDxGCW7xm+sJGCrhSFdX
lvRdNSCixTaTzI435PWfGgtue3o3/Dzbnr0nXodiLWIvLJsLueR+SMxv7XlTyHyByii0MQQ38oWv
fmFGmkR0w5NFPosCVRpKggpsoBOYhiWSnU79amEW+S9Xuog0LtIaaGJA+72l5K85g4Aafloa1IVn
0yeFH7BCU7q+JYWLWg/2UjWJckFbH7kVvff6l8hoOovWc/5HKh/4EDsjqE57yuxTs65D11xFwZTX
+NMVGP/3Irwc7YdNpWKVikog0ixH3/GfwqxnJCD3/ydt2vf2Pgg1SwJFGoygxLBODwR1vy7xGHrD
qGCO9UVB/8+TZ/2ejoChj13aKwQ9nf10m36j2tRpVPtKh8Yeq4KggCw39n8NPhgFf2qGktXizDMf
LAvxDHgUF8KCRF9N8I5hjUO3sTL45UE33Iwd+iEqmb/Tt5DEZs59uCwCf+3/hyg+KJ2Hi/thJgCh
1+3GA5EhXdFUQyBcGDcm6/ADth6AXeU/k2okIPf1oF66yzob//dIWl9xV6IsLnrB/+M0BCJ6Vj46
Aj9jACl+biBFsttRhc9vob3kQUNdmokrLZ1slHQOPMG72K3qNUWi0X4Jgs6iqCy5J6RnHbFz338g
AUTGNeIwjjClrtIKtsiFM/jQCBDD2rk8WvyJ+/yBXH3T62Jrp/gFFzc5XRhQH8fmx5RVb0PNjbl2
kILvPGdzQtRrQzhwtsaKoIUZ114kIbXYoqzNb9oXxU90Ht1x3KIEOVUI8DakXzpsQ2jOP6Q+i1Fo
5lh0cCjXes3eEIbfGd0eOclSUrCG7QjkOqpQ2tdzliuUJ/AnXX/pJNSyp6XAxMNAnqCS4g/FC3+q
JCZls2tvma5gKZeRaIT3HM1+dJ2xQDxGSWR1yNoYSiKYDjhZ/n9KGHSsOhQRxfZczqES09mB8Yxw
amlKkYfV4l+CDIB0HTGstsfqnQ8uD/70CEzq/e+WA4ePAx9Ek4xpUKO2WjS7RxOPQ+MrlV7t24EF
Bg4ppkNctQi2FcHpqKz4pO762wlmpLrnBeehppNE/tWWKT43ha7FpUcVAAk2+h3N2XNfq/xlNyP1
oNNQ3k7w0beRCfJJGZ+1E6qGbWPUhZcLTHPdLeMaU7wQDUWLuqsQW5AFQ0wI2C0gvFi5GhyQyKYY
GVcFaAF9fofkVYNAdhkVxGo0fLK4wP1gfZ3Gkryu6/5Ro5EZeJcVxZj64R0N4EtKUa/XEarrtYMK
YbR9aK0aMm2KNQrHetyPVBBTUrJXp/qVtzSiVDfsMwb+eC1oNaSsEEpAo3z3CMa6R4wcfwYirPlG
BAtLndzbpf0+xdlGU6eRhRWMcSr++qoDj/7ipML+fa3CJGuqqfVfKqMieYCwIOoyCvX4hZLwpDiX
EA8DvfiYU1aC8mPoTBksqtpo7uIlbP0NdB/6t8dvJzhHY2wTEiC3wwYRAx/eqKQaSEihoT40hgZy
jcnA1A5O2A2XYi/rWFpH1dzrF/qPqj/N2sLYgJvfEvSrhMJlm3xI4QvpkQhO2HOT574jfGj4WVpU
5FFkucqsP3TMWFWVqM5bYj9/SwQQqarw6oacXhvoENxwjWZSxrTu1DghTg2Y2HFuCow52bJhASCF
1shRqQ+rqTX0uakYP8+XXx2u9Z7y1D85K0Mw6zW4kGg401Hg+5rJhKFp1NkHf1LdZ4wbQkFtlkZd
977XBF98yruU+MVVOcdeWAfy5eWA4pQ319NioXCdNbEGHEI2QdtxisgNV6r9QLXzF302Wj/TR97q
9QcuAlJFpCni7RYrwsEcFDaycJbE4bYhu4WH1sX664nNMUYYGLBYQ8cN3b9VPKOJO13OOUAYLfyy
Wo3Hb7aYdOetrdTG9fB8VNgjkZ4b+cMrgOwExODORS4qddCvny2mrpNWGm97qE7lzsDKMCx65jaB
ADTnXSVeyPg4TqkR4rlpqBnBKXLPCwANUkWQ5iaERQNvIAAulIY+Lu5ivFNNcuLsWD2P2GdYUM7g
7QSs42VFGNHnIlZKyrFrFwZevRzWEseAGsf8jizPY6oVW9WZwk8HGWKQfA4OW9x+w+hgJsjKd4wK
Z5dG6Yftlq/nRoZdx8VpgfmhAu75A4C62/02o0fnGkuHw8gD+OX3VSQWNWkxuKPaqTwLiGWYquc1
rJ4hiBvRgkYlcnwLLRIX6T6d5VYlxoFhe73bxRnAcE0QfOF3es9IE7CRj8dhtGkdYN3odMuX6C65
Ga3s1FxpsYkhaTxDMVBFnwU+yF/xUiQjQPBVvc5nAlfcXXTCBG6G0O1GJuG2/SooxgXbOiTe/jZ2
+5MtMbLdqmbwm0o4uWF4PQDfxpNJ6vMw/DXGU1lT9Y0tdQEwouFYPhy8ULvgoqBU4kiaUhuWkeMA
Vb2LIRi3fL/TE6lf/qst8VZB61IofLw87qSk7PMpLYfigCmEWvN6RS5MfDfZoAIlUbOc40mRRtsH
zHImbG3DHh7s8FgTTgIDjCsNI8pzntjD/vWaClHh+om7TV3J7v22KpKjVTovI1Zx/BYV9EjlP1F0
mFgJlnyu2kIkcwqBAFzIlfeQi+8CE0ksvHq310ehROM2rtnh/ifTCItMN4JmvCO8DtF49YRW5YTf
/EElhn/vdGwIsfTfi61TziFOAO4b/aQEI5clQSnL/YUdL0TQW52qmJ5PUeFdwas2nKjMKLHI/ioJ
7buLoaSvlCx3W24fh5jBYUR46CpwlfDeR0EghOFu/DSDszBORQd3g+rZxMR2OQNQcadabj8ADMFN
vPdm3TTCYGm5VMf2vuxuWXBII3qDckqs0uNTe+ahknejTxlqfNTUOCK+qM6XXYYhZkP1uImyraIv
lih97D8iwJNJ8n7ar4T+5jGCDNL5XqMo+QtHKxjbCPcwi95DS/nF4vQHEh8uLu0RjuNFug9ZyIeK
0Ct1bOHyU3s7KoWQra/V8apq9iYOZl2jDEyaGwTUpVCuKPyxUwjEfv1b3yyEzr9guihDbO4ZHgvb
1JcltA826YqLrtrCdEhEriAWKzf4Mz5eF5XLFnbtnB3k8QlDnI+4CIs8LXMB6xZJYeCUiwepOmp/
4opq9NK/P5GFCNs5qPno/MCCOYYyGWyYansWH+q9kv+gD0VMvQHar8UTmDpveEuPjkUC5at5MAjt
1mZ23BQ3dIchBW4u6msf6JVM0EM5pcKUlx+cEykjNxamoas3TdM9+GC37UyI2/sLc/NzUUgwWygl
WxPyR/MYhLh0zs7VYObRccG0CbIuN3KOEn0oATFElQd9ouk2cIe48f4Sb6QnS9oUbM88gknjiTB5
JkI5ZDKcrJS2dssAkgUZKKiyqYvOnlbstYSaxSIAfkj5e1j/Y9MH2PJyxuh36EISsOYbMbXBnrjW
I4X/kWfgqg/mMwqcFxFEcypWyc05kEMIFVXOswiJxPtKXWSso4sLxhd4o9dy3y6avPmcIsqQ/Gkw
2UYxq8a8/DVzQzyuda15z55hlDwvYcS9ZgZMBY7gbrjVdbAr/JQVtwlOZvVTekOVmuAmlICUs1Pi
HellGJGKfUX+2Pq6jvKH0pvnXTp0eF567s3IN0KpEMPNSSJd6zpQ6c+pkO688aHxEp/ortUsodcW
nffsvgXuBGtza+HcsWypnYuANmZxKwBV5cYFvS0c2fOT6sJhizkHFL/xTX6qpR+jTWe6J/6AIKaD
Qhhl4BWksxjNJFsLNHN9bBsSWjFt/c2Rr8g+pI+0fMRMnfJubGXGpuPoEGTMnhaJqXCAET5QR7JI
3hSJrz1wc6b/tjNRbO9eG9SwCHrPcrK6imQ1SaUAg+zQlipsScc2Nk6e++rxeSHCbO7U2g2/7gno
Ca+GMce6Ys/m7YP2WpLul25u5fTDCuAmgV/gME2c9yTvj+iGzPvvW8xEIT5pzcjwXShBYXSI1EmL
AI/E9zqeZZYIMG6gH+3xUn3hb9OFMHoWitAqQy7gcV4HsDZQDcVDvOfIJgVazDaHS9Ce/KWNA0wt
dAcb/olFv9+1rVU2ST0A3RL+4XzI6+5bC2mj7/jXmSUKWgN4w0onzxs8pRQV4/eiS07hrGodb6LM
WU+ihGWpRlBWgV3siU4AhbusfNCw1ZHiR1mZ5+Q6gvzw+mUdaxN1qGPm9CZBygBQr0P9P2jmHsIJ
aXmXPCajEKx5tqgtaN3TkMYCXjaLsmH0nQZfb4f5vjH5URjmyc3yzPqGYY7MBhIg6wXLRPmDrdxo
OsUIVPQ6z0mOZgPIvVRxyH2yE8DntDtBQeCBxQYpBwEsmzPpgjZYWTXxxWntgiIND15O/eqERvBw
NazDHq2RHq4dD0O9lJrQQKPRKu+cdTUiQuB/8iPCp1c6wz5dwcQ/kanVgIEB2nRN6S8EZP9ar1p/
WD5SJwN2U6ihvv8EATBinaqW9kp46ZD+Ar/9dsGy+K9PZ7/nLz14XQ3AQ4gYaHCKz26/thpY9VcM
zRyWH0vbqMM9uQOxf1o/uVD6ZxQSR4rbtuBIG/TG2FNcABHKDGR1u/FRQ5bKsYd8fLH7eHTBXjLc
XIwwsWytFx5POKFRWVYQO7Wq9tcWi2XP+Vl5bodFuv5LBFHnvY6VqOmlqi4dZGzg7Zntudu5qGqo
XmZn7cgxWnLHzrdluLSUkWbbxOU1Ww4mmPBS28CuPpUak39STfCeGsV5x6VgIinPl08TJwHpvWI3
nLnBO1sVxSN8MovrH6oUzzKAGZqVOxlUd7OTe5Ju4Dd9CWgJin2sDRx/UQ34EUvi4jaTKYnNy7fr
YcunX1t//YeBnJtbgHburOVTXCwbKFfqFGO4/x/KeGs7K72NM3ws8djAyrsYIVrsSsEfuacMW873
/C0jjGipCEVT3uaJgBAgweMlC74UuSMT8uMAufn6xRlcP0flPeTp8+aP5whZ0jRE4FmDnO5P01ys
i/6AePtv1FY0+YyEpZmI835ujzFarXWG3WsrKhFp2L4LqCBT4VZNQeymt/klnhxyUbYTO0CtMxOd
Fd88/7JOIKG1I7QtUGKX/GXOe/XoyFYSGrKB0JY2R1oDKnh7yAWSmPmqte/ywPUae/4JccueMa/W
ZJdRJEJA418GwK2raGyhy739D01G3vI3RoclRVJIE9V/eK/miDwsgiJQrRTNQyXxCA66mKSqrvrt
IVyf9phBCzE+9qfq6NV4g7BKhlGH8twTDUsI4AIGcnBaKjFrGMknZ7fsI/Cy2+4fyMaQncQSpP/R
7ffpuvctBhURYBNpydBWzJn19+xmq36ymtBy0Ln1JoSxDBNC6iUUiKIei6SEDKgOGSELyz9FVUsa
iVsl9mR+vhsbvrBdpPq7TuKqLGw0S51OaTrbNG8/2wPT9+rqYdnL96cN3z8GxulfAZBW7Zn6mimJ
qxVQOxfzSgT2+Dx2txM8zrnThIcVEhEZX1iYL6cUadRLq4pNEJRiJjT1N0pPoMG8KYfTQwqZSEW+
9WgfvZlJfvJhxnV5dbfuSlvZimohrallWqdR6iClO5KyeLWGtKaHxRdf837rN5UkO0Vnw5UwHvIQ
eR4uUtmAVM+Ua4S4yi483YygfXYM4piuFDmq0Nt5ZiDcw3PzrqkYc8J5Eo+VISktAKTaVMsJQmDX
h5ytaq+HQWUAhjz2p1gNNfGUpICA4/3tRhUruTmLK7LKqrlU+S9yygW4DyXeTi1FWBjl0INYjQio
iOMS4ywiOAqnwJYkefDgZ03aNAEW7AgCyc0b10Ay1mzyNfJ3IXKp8RAKAZIX9RBS7GJTdUhU4kCF
uV3zZHhOR2fQRPamCLPFm6cldjEzsKEiTAlALWbfWQTMmiaE85bZ7FQjcKbC+zWXw22Hwjedb3MT
RjiNlEU1lnX6gKBwly6RyzPxZd7358oTzkHr40498Kt+yMf7tQBvB7xKVxMI/JIMbu7qOKXdTpQQ
Qpx3D5g8aNBMh74E+0NJ3QRzqg0HNRiYmUe+0yejLJtzSMiaMcliP/27HeJC7tjMRGPBJiFHEDNe
5Tgn2oRlj4s12xCEWUTo7j6n9PlQHTuY+sqlupV3n9MvXjXIxiVYNIvwUul5NIG6MUbhMgoGxotg
I0H59SKAvZdOqWlN0oq9rGhbLRasWK/htXP89lAbn04PvyhRDk2y2z8EUU+Qh/+RPatyASWpEHWR
Of58UhNTptFC69bI/qqQ4omXLrCw9B/NgZq8f6JqDDoqok/EHUfi+/GG2BlPixTnZeteTxMhw7EE
oxpwBqHaMXsyhES/tzo/uLVkGNXY3r2+EHIrxp6YahFRp8OHBtFZGaRk5ERHphRfMnogBpobcZwe
uoFYMeBBunmQ/o/0lGXWdhteTya0yjhcdltWh6GVXBi9c3bWebT0Rb5yqkX1UqwToADU/Fe3lmU9
iNp6kU4ZW6gTJ6QEnmQFZWIbYFvWdQACi1/Bg1gsIALRkkfZEc5jHuahwH4HhVsxPZd8zak/Rl3Y
TlOZ93FPaXrQa1yM8PJUTza1FSC1w24bqYj/+WSyi2VRlUZYkHxsCWvqSn2qL2kd3o/H1H7JCk9P
SzAToJ7V0fIa6g1O3mx0q3cZP89TkRAWOu8moSa2k3irX6bOWaToXUTaitqCY/4w+QjuPMez8j1m
K1qrIrJIOaFy2ZBW/IjFeKPyfNYADrOBdCGy7qP8XRJSH1nRtQE1o07cTsYBZCMHQORftI65FqEp
YEPQ5/YZLBSTXgEW0pYXKkS6gHMZ7zI3/OnqXz949VF2OL6TFLR5UJQvAqTP+Jg5Gn478idZEE26
AjVa51qJf5V1OTsOk5ka+/2ZJ8Um+L1Lj+dgYVIdsxectgSSn3OothYoPXmJC5dYZPDZMHzXOwSj
+U0YGrG0TGeiuAlsVpirq3bpXfXlLg9ou4eXIE0kGBbPyGIWOm7Cl5zrjM3ri8xyi1jlRrWqapte
Ro8DUjiVfy+ixJwq5QidOm207ozHklBXcJP4h9KFPezPu0iWpqVpvfMm29RMuONe1sSYSb85Ywh1
g3+RWVdwe0VuyKIDaZ6T2hfXyAyzNvbOfKXMwwhh3oxaq5I9vwJipn3h/o/GK4wjzC2Ut7bTygC4
YuFPGoUQVkj4WiBduru0aZBC0VqBv5Uz7dI2hIMPIUypXbfuSGcesQ7zc92uOq4yCr/8u3ZAE7E5
pHxylQ3yFFlvsnVOhnccGo7jo2MIyAwAiUVPuGbyHv++LPNd97kajlkNcayVkbfQ9c+5nsQixkS1
/21Xfu4CTB23AJ6lxteVKgPtIc2oPfL6dEobV6IlNuyxXeZ2BVryyJzla1XfPgBvdRrOzqsOTAUR
/I1A+6YaumQC9HtaEGSrOXXkvvPgukze8zPsFYTYnoS5wxENzpbBuHq+kZCaELwU+Kdq5B6m2u22
S8jtozxix5m5XWptq5cpPNUms6MF3kIOUijSMktaKxZRo/h9utV94SdyOFM5Yiy/rpxqnkyxaXAt
2S6rVRw2i3wU02lLBYu6R5jgEe3p8s3H/MshGorklD2PdagIo+I3M1ODHH1xh3AfhCPRmvTqdcpg
5uB1bgGVPfqrtmwXNN+lu5tLVMdHOmHWMRuHmwqebEEzn7ERTAIV9Ppy5qGJHQ2dwwKE/cZV9oNh
00+I86ddD3VZOp0EvZqmoyvS7aDyUSo8vkRY3KJDx3sRy0KwAF7tORFzLqJW0gT5ali67y5t2CsV
GBikZymqYtH0tcRzf6War4aHXj3q+SbxyjwLgWcCkBfqPbz4gEfrY5jqv5hcUH6N19f8LLd6eDeC
5sd9HO0L1HfKRRDbMnpa4CtXjDrajfL5mHHEXjU156yfbe8PF5nf7nMgjsEk4mROWe8B3jF/4F42
BD0CaBswY1yJTqqR9kWZp9M/ZRN55Tz1r9lyJdjBQJsmcnVjFc/NHjIMmnZ9LEzZBnA1g+lnLxFK
okTJ5G9OmzYAEM7i8dop5q9uM0trC25IcHtQiO4tUhDjtRuaYg1sZWT3xIOKxLGBxlD/89f05bCp
jmhdYrwqgX52plmO/ajkQ3vDNAiEJWJ39LHu0hR0yD2LpoXf+9QPAKvtyOqWp+Asv0B1Wh5TwJOO
mWJ1HoTkzN9HRGz7UFwIno7zpNAFc8h+7dx9H9vz73db0TWrVlakQX4hlq5gUKPvH+EyiDnn3aVw
XapVbLnvQmHIu6TELxXQkv3c9Oy8X9lzJkD2yryc3i3VgpwZ8s/2usVgssW0gHrlPpXyU6sNITf7
4p2R4FwC6XJzV4Z9clg/t06TS1n7BEshKwDdo+k43WZ9adesx6RCspgUj50P+WAUDRxM8VyNq2I6
2lFDoqNGM/hYeWb/31K+OvpjRoYJr33lcd1lOt58e1HiiEgWQgzqmUvVyWc9XOZDjzGO+keE/WqB
atH43FdclMDAGHhhA53AZ0CRM53q0OOCe+TPqv4dynYrOSvgqovWFG93E+DgdsJFzc7jOt/AJXWI
fJU6V4Qsm0lAO692fK5RWPOthnx8knI3Sxp4foEDdE7/eNXZ44Y5My9VbYL8B0qvFJcSSVboLhvn
EJlvSbEgnPPg7VYxB1hmQP1542VADZ/w+Sbftr8a+vbdkO/nBFylzPpEQMjaNcpgAMfNTtg5WIF+
Kfm3QjP9ktrevlBTUv55wKtGjROOnIPyGe270/UU4umNRhcG1cy09djFJO74nLQGENdFjIf/lYyK
laF7sNOxRM6VmvIC+p9w6nLoKtw9q4Vc0o9/CzNb9UEaH/ofkc3KXR5PRQSPlurK2HAjwKSq5+xV
2Y1EKZozxvV0dU5rmrIWkjKdWjvpD4zN3TuOLPLJFGdg2i8w0goUf0sqBm2awNSzOkfDE3yjRetv
Y9e7ugT9AEb5rfpCVYgsn6XcZT3MqqFs2NQ3CVwYEWl/o0WIkt2ndfCVJxFubfWSuRFeIYjeLxNe
griiQlxdUaiWtLUSKZkvSWmD/9dnGhcniloB4W2NvnJRkDe4PhF/ZniL5heL1wcIBzYCxZjKNMXr
wEk2rpli2nDAqlfnFp1/6dCYuVVzCyfhDVzdNywgPKJcHxEpKDc2e+OO/eaCTaBwY/o1aQP6rYrV
tRh7dO2u6mK+pSoZXICeyMeiW5K/OKinP77BDDFMbYPJ3yW3We/ZYPfVzOoMBLGb+JjqzYi64sK7
Bpwch2EhAaYhE576gRpPK+iZgLbpvZ4Zwpe6GLr/mJBJyVy3tmEtrny33kozmQjZJ7WROUjBN5Oc
h7l5GQK+PPM8edaWn4Si666LlXte4oHOAyCeZI2iFdkr04UedhI8gAm5DPtS0rF/43S/Jj1xgrdb
tHmd97gp82bMnRCqIqKZ3CTrTMOgSL8E/7mT4xGjtOs/6x5x5FVEEK8sf1WTcTkbzssc4wmsdyEM
Y4dVH5BY9VFM7VrGYUGmNoTbVRAsXoPxUzHGbWJRvljbEAyokax9sK5qmIWLdwoj3lSrlcJgJd2a
wbN5YivgHY0QmXd+yEIBiIxFr7Yw6jZEduFC6J9PbgWiKsNbd5GcfF5K1X/VDHQaulOLXfsVFRc2
NE3HyFuJRX/GFXPWkZ7Tefaj2dv3Fh1mxb4SFKxnw9kO1utjmrEyPYcchFiVBVpWaPGyGv10UfUk
YHXnn84VchlsyLu9CX3ek5wP2QR7xVZXeo2v0T5EhKayPTvBbECx3/T5TFdq+4pbQQVrv/Vec1in
oI+k0YdXp8juXn7JWQ91U+47IsNghKXXhN4eQCbYFScyD8KknRgHhToV5KFbyyUvm8C8M3103xte
Oghyc67+9vf3/H1cQL/kwBRVsvvR6I6vSBdO/kcfVZ89RoYls5ho99H4H/fsfl5l1etLegwAbqnN
GzljlPrFLbLXhlmF8bD7R8sbLXOvZTgelNlFFdZePClXA4Xna0OWdnspvEuhQ2IPKMZWRZcxNeYF
Bz7HVpiO1hdWrxGzLooDFoWu7CiRisMdwBn4hwJhx0HsKt3Uuvcrqaf0c5GLbU4vhirT366jc14f
FsUWn+FtWv1RuSFHlxkjwCznqErh1zxAlMGpds67GOj/dTKp9HK7FYT2oM2mPwZOH7ngaixNzPSJ
u5pEo0BcE1WdzxjTfKPwkHw11bRkVU73OxhaABf+TIp5gDDHP8ek3DdUg60eegnW1JF0caxBlfPj
6zBh8JZtqa0g7TDjkXouXI1GBG9AvMdtCQ+gEibLVrgJb5vsM9wgOSaKAA8UEOwI1VLmKJs7UeWp
/Ds8Me8hPgOP16axkysO89F5KQkkBhThScY/8LEosUqOkS4RemMmR4Loi9OWpmCOp+duKUsKJ7Ry
OAD8W5i7RLQjsxL06U3l73tUiJ0ppTdB2M3giDY1ZK1+bQiu4U7l0m63kCKF3dXX4MDkzWvIrSOr
YCf8x6Kx+uQuythBXTgK7IYrxC7hgiuszkhRKO1oR6XeuO1iely+p5EOMoZSQgc+Xe9zTdyTjiLi
23GnDQSUl+XNLhUYv97WFh0aTAflrMEoGizGC8Jq2MlZshuA+srH5JMOhkvdhYdth7vUpWH7x/Mn
S4sze3Emn5qcMOGco3XazC2LZvRCLtRWByFfoNtFWS600p0nQ7IUBUHKpJ0+7y6yqMqbMyZRMolL
aWrYUtOPczLv0Uq2bhHrSQmMgcbdvjawc1KQBlVVInjTouLo0CIVdaoKYgd/ZlagfSL1eOo+vYXR
v6kPvVuwp1XU5ALHP6LDbcHHQeVzasB4ztGM1MfZ8ym7zqW2W7EAwAVuiEKQAwowMv0CfsjQ8VMV
wL08htSHxhVhOYFelQMQjPeEKTCEKVhOnoBd80rGoX6DDlpXY16SaaV4Fbm+0dIPKRr6S1JvcBZy
Y9CWbglxgP2k7GMXUD7ZeydgC1nU0fOOGnyNL45ocyVt8la8hREnsHLQ59McLyttswHBJRYE/ZEw
DoVnZQuS8Yjxe6rVGNPykUcMo9yKQpjgYYdrqxzf81NV7whVeUIyzR5zJthd5OTryjj+WWrS9idG
PIH7XGq25zOXe9xI/jsLnQjG3B3vgnCnFdrPng+9T/7t3uc9gIBOKpGGdxcz9O270Aec6BAC9Nu2
bSrnxcMeKELZ7B5pTCgpHDBsfCRXK8T084XQlsUMQPSj25Ms2/SEikdcloQGfhrhoWw/NEZ9EhvW
9XmYtAss2sZ/GbEIWzjM8dGXCzcSp/vVB0Ecuecponseze96ZiV+eGOqhbtMMBKRDVolOHFPErBC
4OP7SlEQKAY6lhavi7FIOycpMhI2UR+x1IatRChVv/i+8Z0e3tfbExHsRSBfXPc8417UbQBi00hi
5v9AStjd1gJW0phBIXgvGfdsQbOV4jzxWN8TCmR1mywi4w7f9CpJf24qsx9zuboar5XM/7aBbHXq
u2/BVyx4axOg1w4obQHVLbFfPedkDg+YCbI0fNAIXyZMR7rLsRtISB7dRO5161HnhzkcwPbhRIh8
vOYpwURe4vIKyjDT35I4iCiasAMyJV8mx1QxsAdwOxfDbUTy58Rrs073xBKntdtrsYx0bxnVP7hK
ikP2IjpNGDJuZh4T7ZUxq5TUlJv5HlvmZ40Sb4OH9KLyn9uQ157KqWJdYD37/kUztdCsEdqNbEyL
/5DFgxhfnBg5Yc2b4UKmBC2HOiXihrrz0R8fTFcdXY7DquyKLxr6uC7i02WbIOORcA+f9JRw2Kd8
iMNWfAfZne2+22Jm/U3JJTY8Ni36njYz5psIALq/loxnI5Ph8GYGFNUQyZoUCDGVkIsioMg/MSbD
YqzH6f9rjn4SU2cmkpdTWK31pMjXMhWZuF3l4Eq+N0kIbhrlZIruEVZvCcT97HKFQjPrfH1nbCZK
cmReN25UcRSH97OSEcwilTif+u9Sjx1HLHOL1H75GP/y5EvhhIJxqq6ZQUEV6VgJPGVXeNdb3vAd
/3MyLpUuTfZSQ2wed8LksW8MsmnLS/VmvTNowII763SvmOMX29A4Xb0y2wsHvv03L0XxL0qpDEGy
MYH+7aSsdtRv3IWvJqLDgxIOFCBeNivrWBFkoSBORfvYe2FKj5PrbFQoWNPP/vkxjHcn+ResAyxw
GvN4VKibbnkC3pd7TVlqkpcdsY1+dfIdumWy7JkLvhqzfeRbqOdAfA7ilaHcle4tkKojpE7EGas0
hl1bLGbJ9qo3sKsGRcToTPkog8WPxh2+IJXDBPopbAe5+NPe5xijAMU4yPwRUjnkEsOCsIqgWNqf
Qb7PSnIouM61N1CZhxEvSLa/GKQgWpqVh89cnQpbBxf+fRDZ7CPPBg6AOyXkwOYl3tfwvVHvWSG9
lYxofptBgS3NGpUfycPg5eLegoTHp95CxUaf0LiXc8H0vAryyWbQmj2CcN9Vrxr8VuZIfTWbdmxi
Mx9EtH+dAU5KJVUDba9b12PPiCxELYeCF/5UwOpA8gD42RpbAjwYyxNeKLua9KHXrVpM67TbW8yQ
RXp5yCGoN/i6ytj/cv0LShovfzLvv+oQChQUmb8VRfrPxKA+uAA8tdNu9MDlvpOBkyXY5mjDRtwb
+/oLll42IxQEu1R2wX5gujj9ZKEoD2tYhVF9ju6MX6QHsiJ+44yXH+sruxGFNyMVUexaM0vrKBix
nxZf1CfxXlO1MxSPMVlF5DyzmRdZ7SgSsk/Dc0hwBn5u17jF033EsqgBEXlGh/oSoHbZPo8Bh4ob
4DrWeyDezRBgzCV/6GOyPzLXcGmyYUIUM4yNy4NahOQp/9e5juak1F+rSrf3n0kmIX3sxSUowuAi
weovnAUvYqhc+hRbe0l3ouR0H6FD60dqOev3PANyaQR+ZoniDIhx6FjiXT/MO4iPpajuD7NQp4Fa
w1drmQFawKNHRfZqXuiH0gx7ahk0Ud2HEU9UGZBH25+c3H6UxyqgZzlifCYdQ82Tv+c0vTPkDvWR
XqZWY/Spz3VJYq9SvjE1+yzvAt1H0kM2KTmpTbYP+KP2CSHKzm8BjNt+p1SKPNUN9uOx4+G1hzbC
5ou598kctlJx9eG6drHlO8/gYPLZKkHF1A/zVMGRkre2/MaLxP/Obc+/tP3SI8HJ8GXI96Uez2Tu
SmA3UhEp+dduiEce0fuAw9VdPtQVtthrBIginsQaVWhqjRvOkzkaVA+mUq59QD4MzrTowqsB7Z0A
GFhrl3fnbc36WXvxgLuCPd1ZYVEJcpUXZNhJFOjJa50gejkcXPbKiavDxueHrY1SczTzYLPUw8z8
mvBAqtMC6jMr7/7V56vM+dwMC0vXiYTsOnigd3N703zKe+EjBthMWgpDWPCifXCTCqpeDKrHcKwG
bUr/J81MVQL2Ae6nAuoRKiRJPikNaNTv86Y4JjQSbw9/Ujegm3qirWixIQFStwiazvOCbp/de3gu
L4iFcQDKrJdU1wgmpsS+m7mOHr7UBZQavOUlAUQPlu7q3h/SkTxI13kH/ZABLJQ+V2o1pDr85kBU
rrTAimLLU9Kt+ISCv/5J0zTMJ1kmOqxkCJG8PzVpGa0N1TgReoVYbPwWNwjW7zT25PKzrG6oeF3r
/X9+Sh953wTRYZSPdLlOy+f7AxId2rGiKxmK4/i2l09ZCPay9mvGy+wO6zKfbWkhFVd4xO8KtSUT
qAcElB6rGd5JYaALc6YnS67F4v+9XYnm1TIL69CLbn3ZV4SVZVcG8kwzTNPaBVX+xwP8ZpejVAaK
ClpumwXPNvxx7edriBoRndYcbeitY+W4WBhpPlrJ9wNzRidUPCqQSq9kAXeegrjkSwOOhgMLYayT
dC2nyfuLQ3IaoPbK0k3yua28gc0ceVps0jcLpsA+AlmuxrXgM8dRSGWDIvopl4lBkTviAIH174G7
QoXYXPhWJ+0yqjtSfb2rHJEnbPV3uze9x2ARgrdMta0cBNjrUrK9HBVp1IUJboW46nGBi1GL6oPT
+RKXB/zUGrgl1RC74Pt7EXPPdIB9TgwHzdR/URuhcLfRqAtYWyyr9p8OfXvFsutaayckxv0oLoui
WmurVqiWSyANx8gdVWNO2drS6u/o5gfNZ4MBgM+jhO7dd2DvOoGqrzQGziN26ThiWBpn2K4cWxPp
kpn1xm3w+6bwGk1JOr1op9acQZ+3WVOVdpr2yatYotzbndvcbTqga1/QxQCzbqIzTPRyrGxRuBzQ
9xGySLjBHPrfOkkkx3PSenrdpNZR/vVnyvzTRoGTQ2PaRMJw/iKrth4cSNH0KdR8nIjJp3fIUD9a
jS1C7phqRByoOkIjTGovICDXp0k5K/7yx+4IkqPhHo9BpBa+SQbfl2cvPyMK7x0o6TYm589AfrCs
8YgJBp3VR2iUuUz+g77fN9lQXZDdaATEMDSC3/CzZWxSeaiu7bX/I87QF4iMgVJDEu2/Wz9MXIPV
RmzKlEsww/81GtEJBPQiYQYEwNTh5v3ZK7/leMEsMPTBnhDhgREiy7goSPIH9CRKaKQez+sh3jzW
ZV1qw15Hq8ovoRJDvvh/Y2G/9CrJ8JYem6/JkbknWNRp2SHSf3sbgulMjfBLXFdpuWKb9yIOChI0
6YqfahMu02gsuDRhqm+goAtvjNlbq5Of4a1CjmR6fm6K21IU36dJazo9HYKWAaT44v2FTcV8CiHj
tIsCWr4oGmx4W6MppbWxsxptNhIAFPvDR+1O0DSqfAebDWa4P+ABa5bLplJi0EKMoM9J1tNvyOh+
qJUTG5Q8ITCR0wIcqFiLTxsg/rPEd7jOHzSOp7yQ9TM8Pi5XMKfUGTN4Wrq+b9C4mTEWew6AyF9X
Mi1OFTsP3ydflLpgjd5Ky4yNDXv42D0AkwGNYEL7fA8S22FiT9iJ87ZXUTrhJA/PnSQF6p2+CmSB
1CtRbyO8pfGLfaoA4GdtW/OSM4T5e0nqSmyEOROp30snxC4PSaTGMWEIZntybnIvOb4iRbyHxKYF
gC8JU1+Zq49AbbhzJ5RgyIpE22ncfg+xPa1HXC1NC4sNoKlmU/rh2kmAAqD6Z4ri1dIUWPejBZDI
3B9qYk2/PPxfzWOdAk3DiPdq1sCD+Kyiq+pZyIaZFWoIsk+v68/xjgfo2bUE83FBcKGfzHdVojfn
x9mLYIMIcPbwNI3aRRJ5TOs7jsUqJ/ypPig0GEyuKKKx5q4+CWQ7Q4TDuF65/CBsEH9aAzVw9nHr
cl61jtaiTQTFQ3YIROFivlfjjAB0+DJq74zJqSOBzvp+JTsVt1ilpeAjUbT88CkwkH2nQj7nfNZi
SSQzweL6BA9HpAyzBsovURGESlCLNB9FzOdOjNS7jgwT//Yd9W52l4EHAgvfzlKhmEQBQrol9DnA
Q/xPPqJ4+0CjRWf7+2q+wKC2638Yo7IyVFf+scZ7NUHRhsdr54fbLVGI2piRz+FCnqCnTpdtprwP
HwPMMIWXrL2dmlBjhNmmE+NwrVc+EOFKSyTaz2hhV6Az0yXl+pRwKaFub9D5lGQF/2oPBqOC3lz0
uuP6wn/5WOgGcuCvfl6bSyaGpetR8fia189DsqeEqUQ96q8IIW6nJGnoauZfxbqoAnryeSl0fpiV
OuGb6dxxtlRr3qtzJyY5VtDp562FTJPnEqQKVwe2XodudrfQoklYlB0qLJn0V+l3BxwuOplDdlki
F4+8yK7T5uQ0SiFpoFvTpPZLClQoK2ur8wWYmHM36uRcX8Cp8scZ9Ho54AcMy1hVixhyJxF2Qimn
UcWrcN0bnFXC/BbjmiGckb927zAYtnrNjDHo2qcZyrFidgqxPpC7xJsMmVconeB/V+MDyukOuHEO
pa4FYcUjdlaQvI+bhcbdxRC1nLlx+qjfGWxOGtR2vuOwLEaRb4Uiqdjrbx637BwdHlCQjDMqe2zk
3iYFmydGB7EhrpfIMRVk45F3RW485y6yiGslb2JV9uMoPXsa6acewzVjvZ4BbVhdXMDz5Dwu2Ehs
BRmQjoUYHc71MqPZsAm3BJedP9+UrpWRoTQ8tfUs0Y0fdoN+47BAesy6j3UeiSK6CMvpOyusEECn
O3rTlw23kgNCltCiOE7woF3kRKqDxfee4uX79L/8zB7E7YDAmu1oWKy5yerJYxFR+3v9nCpWL6RH
O02wyglbQws79XFvILfhimDe2PvyHsi/MAacvDSdm8yyjyjY8YxseVgIV/Apf+WD46v2+UuXs6gX
pv99/byoOl/PH/wwgkYIGk2JcfR4LrknrJG1SQxGhJI5ktWylfkgafoFfIIm2rTms/jbwh5NJSWA
Md7O1UVtYoCVTdyW1ibgp0e93qUxxDF6/IFwmAO6WvAcGboMaUC6VNf6NW6ZpAD+kkfk38lKYl4Z
ViRD0ngEIP+KM50O37yYSNz+iwQ+5VVw6a5WwHT1tVvrlA3k7u0kewTkuulIbp45hf+3zKGmJIDl
iQkLyLW9iTvuwFottPeMuxwa9eRuF/l0zCRus1nqLWMeu7jk7o8B3HLh9bSQwHAdpgNfsrm7hN1O
jArmKmO+rl6js5VGTzb6HQ3ThH3GuycOkF+qJyQo0B7zXu1f4s5fkSjMJCzmoVV9hNmkZ2aGj6u5
yyor/rQSjOZM550kMefX59NsS93yi3lwV0zAaxdRqdwGoYPCjbR3FYNMOCQuu8OFINy4ipYDqxmF
GmZg7vZJDHQBEhU/Cy0WZAdmrRtj8T4+Civm58koJpdJ9JWTrYIYLMy5KFrJRxZo+5C56TKKkpcp
8KJBtLLNd9x7rbpSpAYwjw+JApqjy+AJx4oVtIhjHe9wgjhcGNcTu6cpB58gw1hs0cekVOr3CZEb
XvVhpDT/7ksUlXyGWOJvTY7gLTaqbkYueN/lWHU6GO3EsmcbB0QVMVTEU7b7F9Z1S7AYyii5VzPK
f4r2P31q33BF85yuI6fO2e8oqxKIhiLOmTR0MOJGJ92JsSjAM7ObQ/93qIWDChtQlhI6sVNu2dgy
XMZ+gYKzAecY9ZQfAH7j9vHJj66p8mGzCDTrEuw++iYnP8OnXEgRH2OsRrLI+Z+J+1ro6z5Q69zN
okde6F96ulOk7wDMQlkaLpokKjlmftjHsa5J0TYpQAmvg4idadLNEa8EwzAGiWlGNs3ZLRwCVFMU
ceM+9pUVgKLVt18qowDWIGGWeMRqT4DrVIGTgu0RlkLQT4H1AoM7r+ij8v99YQB/ae9V5nAmy1PE
BXxS8eueqUkU25cnVDkcwQpiiGqtHBc1+JDIXIPGQjEwfX+eB0P4XdWsPxjwLf3NHZsaMttIlEJm
b078RlVcsuTGEKwKNUzEBtX416E8NUo5YIXUVdJSr5apLIcS9ZCMy6V5G8nwLfUjqgkWKZ8wiIVc
2JEh+C3+uF33oQHsfxMVFVt6e/1CbmGJoNIIhSOMpiARZma7YPyFfmmHRrY6jJD8KCQqNB6ObDO+
yL+aouLg6kG15i4ycK6VNGBHoR704/YzBKQTnsChlBiRvKjVEre6P54689K4rE2lDZ9g9Si6xW59
oS/Stwge5i8/JrMW1UmlfNXQeAE5gtR6Vz0bP1VoFoP62OT9BqQc+k/ItnOOCYpHlZ6tHP5/yDVS
5NjZAnrH/6r3r1vfkRAT953jVQUBHQG085X9Xpcg0KoI0aYqihJvEwioftbulJ0LP4/0DjEG8aoJ
ObN7q9NRPUZbb/B/kNzFLt6BxHzAAFlco2KlBPI9empo2CvlQJ/Gmo1EURganiCG9Cw6FgnH3DfY
r/3GzNcx5cfeLIMhgO59iiUrjwXaZfIByo6aofmcWo6mdHj0ng+tG/DeuOoH4aKZVEfgKI9ON56M
XaSqkNYmxMH0IkCWOXyJOvxB6+du1bpu/3ptQiLMQ5JKxKalwQhLO4U4gz3aetMU4MrQyocDlGnp
7f01XR7wiMrf9T1UBVOBRA6EoWCYUOVvNXjq4KMBi60JmtjLwvMArXvd/YttcNbOe/MWiRRlOdIf
fYGRXusTF7GaNwgnuiz7dB18LJqquFWeh6lS4oAh64AoDeYneX99jPNRIX8bVHbxmzJKiaINcJef
FR1Rbhu/HXQ8zi2LO1NprkpsqeSIGZ3vid4E8m+ydnIM64NJrq3CjWVNA4tN3oOdBmfDcnAwQ8TK
qDmYNdofUYIb88iVxNVmIJLny/J8ilRe5n1YjGAfeWvZqaG1Va0+b6dauw8/ayUQ2LeCSQnzMsOq
Ry9jUOldH2zVvI4VTqwHV5DB/0FeT/+sXjUkgqbSErzab/jgdSaW6YzIxx0lXHWUtzieb6VTK9HI
54HHOzLV/El0Ra+MyW9Xy+1pd//PsCWMwWP2i2oZblMNVmYPd6HvrM+WHteJf7SyGfBF1irDZEXy
JiLW/KMTTIbohX5SOm1QyeX6LjiY2+yWbYcZVBQPKi7nBc7+2Kg2DE4HI59hMyZ/MIcP80bwI0vv
0KqLfgflpWnW/sCyKG+ZIo9vcV0ltBnzH3GY1me7mR+sBgWx+5g98thU2zP9F0GBKMWtOB+JeZ0w
OqEjC1cgs/n5An3+wrTPSJ601XCGi/NwX984+iOb/0/fJ1Bv2AbJ/sn8+/1sbLW3wpU4WVUb06pe
rctElIVxuYSetnV4lchF68RKSCSpBeiFJ2t01Fosy4+7czYOSA19sjIoL72BOMCSF582b34ixsiA
2/oUHHQuVniPqjB5Ko9HEhJNYpByvs5nVeGqyGFZJpTBwK2PsFV6JpEaWcSJNqlXWEPxiBi6kcvN
fr0IoIasClTFU9cAvF2shadq6mFXvp/fj/A8IfOtmO11UU4pjN4dzjKVSDvM1RFmHdZB9cp/hXmf
ISD/YucAX/nTVlqxWDgWJFpscuRbKVxjXJSTg4ILBPcRKKtH+Hp0ZylN54qvGy0w3lOzbwAVxSGP
uWQmT8IlEbL2LI6sMXUQFy9eqski6xyfO4qR0SNNMwXkIjMmk4Ht1sewGLyezATHELIMC0W5Rdgi
XfVl0qT/baLSUeiyl6gem0SNvBWE+G5Np3thio6m6jxl3X/YilV20C42VqRJgmRyJc4GFH1DUvko
md1dyXmpboNfnDWWAWElWkq9xAYt1frvdhOX3n5m6wUujjoUsyJBD5sg3KEeczTGYxx0MA9xB7FH
E727HdfWe178ZRyZ5ViVTJ0YAyCFZpIS1Hl3wpJTRdHZ2Gt/6Fg9WmiRCkZlXCsjMc7wvyCc6r0i
d2gxJiDZ4qUoUvWOUPfsYQSDjNncbmn9n/yCWXdr+d0OYE6H8n6dlIrn2I0oeWg/sBt/XMvMBQR4
z+jTzNWnHS1EHpEFNftvaXpzltsBv8mMrPQjWOU6poiFdMH1NVRGJpcuzWhCfZQMdS0dJ9myatiH
V9wxRLxwZGTzHzPgd2B24YJJba4VmEhDuRdIsu+WLYz8t4e4XjCrSyb9DKZjF1V4VRGYPACPJBGT
0+PYV4abeOAQpwy5JxFuPXpLK3D/7Ba4Ysy7+eAmenl43G92ViA24ajAjS+OlCe/7ns3M+JBv4cP
u8JaorbQtP3u8pqY8jjEN24329jIEezy34yXBVD3UHpz0KfsjaqFcbDNj5R23hb5/K0uk5iActVg
5Wv4/zG9RCLsotOaWMWw6C0+O960zz/hRgQNzgmAX8IjqPnQ/eyTS7xK4mu/Nx626oVytG+iIRtx
TYXsopV78ySQI4sMNtV87lc7ywZw9+b3fyWq9j6t43/v8AnfKYuk7eMAYR9DHJH3DptH59xRPm2m
Yz2tW4xuusdQqt75KtfThaF96eUGhJnTdVVEdkBPUd8C6iMj5iAxV9/l4zT8NEDX+//WKSoUcUkD
HYgJjN6DoRIHezXxZE69Y6ySFBLJbKRDur2Q9cdQaigxSWFYrQgfnsomvLnKd4E/FSDBr+ZfTqtq
bqMgYoloUGRJ1SCcPnZi0GNi3eCuCHtbxWSrkdi4Zh+eZV6FkvfpZH+qvRIP2Sj4dfS/idSviE3U
xtV3GLI6muVeEZIggqo4srknuOjYpLTdN/wSeyK/Ef0nVhs89jHOHQbCbgXWS+In2eG+bfHhmnqq
JS4iY7Q3A+b2ojvWpZnfv2TZpzqdXtckRM6nACDbKv7LL/uC8LaZkPtlShJ8vUyPEqrHNqiVYt9l
csbhNrJfLL3QG1rN+mduJd6Qn+jjjiiSX1R6wUKk6T57qcF2sXufvV9OP5sXIZ8JlpEtQdydQ4ki
JFZYf+pkIWdWVI6jktd0NkIrbVoiTt5TzRnYGnDz5xQiqFgf4pk5qZJhVQI1CxWUKd9Da/at56KS
Mfp/8Z9Vr7T78ffG7gotVQ3c4TpxjjKXMxqHrn8xQeBmbeoL+RjEohPsYjqRATmegZyX06mMDmTm
EZ44yep08PSa9Oj0KXa1Z2e0ajcmR90bs/YCbczCziyMy2EQmy5Jc4yqNeU0GjV05uVcG6EFJH44
mX88rYBFLlNOkeK0fvhju+UuZ6Prkpr2/aX0f8XPmi+OazG/pISU6LsALW45lUZgpeptN5e1JsU2
KuiOa+GneBF9bIfrnlgNhpFcFPZVocGRvVgXAPcjoVnBc8bL8z2keHBb+nWExvHsq43Ikznm/JXR
f3RUdpH9nLe2W3kmovuzbER8POLw6yknH2tyQAACXq4wNw8OnpUNi+jZj9exqdOS69khpkcy53AK
3itHb6qVqBNi5dqrDgunoma0MRMrvtbOtx+Wvn8+nlaXEvtFA3d6WStWGeQ4a9B0tQICz+PfbmxR
BKw6CWDIc7XC2rG6N1jWSCwDATUEdfnLikEvGnJkadcLFQndgNBVcyQtnvC8nwkkNSy+vDaUciqd
S4FH1HsLIStn+9BcDCDc87LjbWiT5+X8mgnfumH0AnJlgMRwmU5yu5Eq5kK+o4COMMIsLzSWrXr6
4oEYJe8gwOe5Y84TtWcLu991n6lPNOeTMhwjS8mhNEczmJdzwanWIyg0nw4fs9tH27evyFsEVxWN
+M2vZp+eRV1q428VMy1v359go0QEsT1Bds5kXxGDokZ3q9oFjemDWj8gfL7KzNgreYnEnkbIGMus
JA+KXLz9a1X9gl6Il7NI5zPJSB4h9KBG0HCjLg0SJo+s6UtbLzZ5PQ0i2upkq6zlqyE9S0g9NFop
dEJrrLaTPDDIOMrLaFY0lsnSOCp8AXGcRQf9oRyuoKFQ1zKfVRaEP41nPeCcU4w2jevs+ML3KYuB
rj8OCP0essMFO8d1veFPbnM83d9Ad7VpEesHti2rmfGV9KVnyH877j65E6xRNOsT3nWGHs4Tusac
t9U8oeAeFB3ss4SdmE821BQLnx2DziJ8pZfsps6yCrIB39mKoeCKXqJL7wmklugPokerX5DMv/wL
Y7DYTaG1AiBldbaKwFnk3+3kqWeFqYcltu552Cq8EVhJf//WUV0C01k96mQVCo2fuAvvWFQwtN1q
aBZ7fjD6JiHfyo/paAy5m5MihKzgI005agfO564x19piJSs8zJpYk+6VAETTwkAdI12QWiO/5iqo
SA803uVPJawdaD7Lm2KG2sjYwmSGRQqAFTOiSEul51h645kf2IND2DMwuVEkj5EWGkCDppFNW/02
UEePbgHVtwRj35WdoaFNQBCPDsUvGUMRcNt1j/2u2Wnh7SbmSGaYL8YYbwiUFq48Qj3i+Q90SRTQ
6HJAe2U2kS5oDgXFeBiE4Fz8aXZX3FYa/nwn4WmiGmBs1Hf2eG9wPviiNKketc48UyUBvFsx2fua
Rx/QivtIGKmZnQ9LChLocasMbZBbUPUQRCX1gZbxBtbWVWxVAehy34fxpHqYYOJEZNrJ5hiVWnb+
VQmvcxGDjn0ffUlYAQp9PeeahfnK9kCLNkAYokaYSX7PrSNu0WEFZczNXC8Pyy9Cx4cA977ufdeJ
1uDsFQiQENJAuvTlDJUbbSeUjspUbKuUIR9ILWFsmh7PErPnuStiBykke8MeyBonKya2v3f3veGf
YIw1dHbjkGaHZyA1CGHEMbTAfwszOBgP7wLK0jU+jcNKBNwPYrE0Lk8cXYxtDKd4cBBfxPNZsnxu
hqYZVYNWvgDqObu7CEzRsSnrkN2RJxB3k+Owd31ufbGPKzN7eC46mwvmJcMicILDqZJB4x54D04y
gv9es98vEPvPCvxb8tsEc3xwInQEeLkEMAXUU7WxPCnK0FZQSDY7hPTJeqXOBAxRDnff1DyXC4y6
huN8sXZGzReAEZ1Dh47te6drPMWrQg1/zgXulj/Vt+GLVC5zKA0PYkcs5rbKsnqdnhTq2F3xmGOx
vFh2xdNy/0FxuqblO7yEORkxkERXcB2lv5hHokkzT45uLksjN7NwunIjA0O5oNEvhHtzCQ+pMWUz
uoNVoXIKdCyIFKq7k7JRl1w6hGcSlwVTluH/otaBt6Dh/D7kiBr3O50x4nvFpviXkwfLbq5yuK36
XjgKkdU7Ewmtzjbw+1yEOAVy8NMrv3kWdgPAeOVsohc0wCuWIMlazPjURAKk+VWofwb1gAGywEIQ
0azQzyIC7eRJDPy9P/VI3GdfSFp+MqLfOL+E6RvSz7jIGUNlAiS8JImjFiVlMgaeCY6hBE99Zmda
DKlNkFUbXcQbtEOyq7YUQu84pKW5P7qBWaZkSmZPxLtWZDbHpIy5u/jItsSDsrpbdBNZ9XlU30A2
8njIJHGGar49KIJ5Nedj2xc2b7CelHs/MlOcNFtEEtv1HzYVTzqUBqORighREt97KgYOkdWA3bbx
AUnuUkzum113w+8fAgMss9427bMIu/UA1yFMZX2K6qY63X/Z/Rk9g14s8+ekDcANg5aC4SAmBMvH
ZjAtPGg36sQYq9LZydKCCHVSr0c83KkYsEJmGoWpzC3H7K8ezBwcvXwcaUPvC44D9JE+4iUSHveB
zp1U0KYmWOPBpklRrtXlbXNuNiSTGGlY+dGUdq+t/5a5oaoVM0+ODE658CGWcFIBL+WHpn8b5b1x
4opdaI5HdNdxqAOITq0U/UD+QlIsqqacudWAd/arRo7rZIQFt/LzQELUcsp2699hkhHOp/D8JXpL
yFzoDQFgUTNUPwrwSGK5OPf+oNNrOZJFJzbopmXHn+/aGZWvVEchpoBSFLYvwBSLZhIdgH0/wr+/
0771+zOQmocYmpuBftMCAJB0HnG6EKNDHoCJevK/ayv1yVEC8CCvBIyz2BG8n3Ccy45Io1mYNywr
UIr8/kTNfMHjqmuwA5D4pvo1q12t9hc8wGZRbc07tVpCCd30XUhcb8n8F6rwHYeVnWDSs+Etji5o
X/Q8x8wonWkXog2z73uRSrHOE0N10cmn1jie6OAOFoMVP4oDQkJUSl4oMNx+bALbV0tVPEcHt4Zz
W/UeEMLbVQEM8NX5cwzooE/sgS/XN3i6vCACxE09gXCLQUnAveXbBapLgOSgKMKtEx1FygIF6dO/
6LPYy6YNjJ6gRMU3NmiwgA6flpKjs60/8lwHl2Ly4QGPGCLybY8CwtgHBhmo1SflQLKDC3Pa016d
zd7XRFN5LsbBdSnxTN1ieAg57XAzq6kWDpYWVajvZQReTNVn0qVnrUmmvL1jJrX5K1Ofluv62FLN
zFR0Xk3NG8iidQ7tLst0D/5mNdAi12hx8QiYd0sUr6C5knUK/hbR43/M8hzv2atgBRRJrIWa+Ixo
pookDmq7XlQ0tCHXAaXKCFHG2oSa6iq2bMJg/oDbXf+w5z057w3mSUTYhS3ojJR8Fnw9Zd3+botF
gS3NkhAaz47kjdmUXcGVCoEt+0sYTh9DAJsPbaNjTXux3aUp8yDn1B5PgY/j0mA2OQo7kP5x01iU
irl7g2zGyf42Mlh3H8lyId3llTLmPMfnWc4tADnvinBI6NKagnNRZBsV9ZyxeIe6fu81UaviGCmc
jePY+cAKU2GQwN+fRqdcY1SN9Pw+EXvn9EyXUHUJmLAA9drhglHtCyxXXEAJGl+4Okkio7ayvKPL
a32uW8PXYokHbekSCzWQk3cVOT9js4izCPBn9V6XC3ZIwGlrA67gjbaB6h8vtvYmxJG0uWznnpJK
Kg1GCJJGnjajTFxxgZNpI2ggiUDlqg39I4usCEMD2IRjcCWH9YyhnxhKLbxxgMOdPnpOrDvKLaMn
xqt5eytDGKKkOLcqSFbwhhngjvxs7oYHUH4Zn5fGHfIgHd/gWF8vqs7LCWSPuU5A1HEBu4qD+s4e
7Qe0byLJu5Sds6J/lOmRusOl0l+VftOwjmY/FWJYN41RDVx/MU4jd15Kd7akgvAM/ff9MX7o628O
G6jbzjpkdhNRPsb/y/1knwxusmpWGttiFdZrXnXrtI0NrH0xtl0EP/Q+CjPkfW0X7zgvMRl3Am3a
50qOnHJ+3NwZlhcRKlFY1EqDGlTc0lu0mVDKmQ1M+chqyMB3KAwAEytnFKeDlQxc+G8bSmMjqie/
xCqzpit6V4GoARv2oHmZVpSDXD8hj/Vn5lYGAfc5FbgM+juhw2rTRmcqgHjpnc+VbrGsJs5wJQdl
DlE2DzUd7n5i44fZiJb9iqaPHN94IRKvGc7OzbWoFbWL46cClChXZE5i6rBfdK3Ft+cuYRiGxoWU
9J5FB3IGRrmuZXUcC+W14Xd+CYNvzgAMuyrLgq5pMjLXoTgDJhuFYEKywYQ22uceFyBUrJyueXkR
gXYthlmBDOCQ2X6K6QoF8ZKJGcIcD3QIQ8VY21ITLvaEMr8e/6cK0XMLKURihDXYK09b8hGjZykM
xoVN6PWCbqaIo+4ZTI1Ac06yimsnuN4Li2t46eCU2NFZM8BY2KnQMjC61g7BxUANGhE5G3ZXfqEN
EYC5LuG+FkT3oZJ0u8A2PAsjHgkeHdhFkBHoM2eouE0Z6/svaimGnnYEYz2vVa/PVPLW/I1q0p50
6a8sFS9gIGwm65vT0OGjAoDwEsg/GmC1rq0gGx2CzEHD7bEybC+2P2cqbAtYg5ijEw/W2m3j8daN
2NdQ7SDjAM2RkLJJfXZetp1wlnAnd4wP3bszNGbcz2enPpvwbz/Ev77WEzSQX0O17+lpDMFM9GBU
D0Vrq7FcqDgbVtNMVfRbUGt0Re90zUYRIYiDhzT4aDFeichZSkNvCd/TyIHaHmO1IsuqGXzX26Xt
S5pTKMTU5fPLmA+DBAINbHJTkcjF56fDFOiIPo1Mwx++1Xd2RVqYXdAOXGjhOmwMpsVIOChnsPNc
MveOS55bpCrMqEnzW0ECWt+/yhimHDBthL6pOvuSq6Y+i5WRyDhW48G9SXPI+ZzfsMtH1xWM3Tze
P2McyJwA06DtT1hhppaWuI0UEp7SrYjN22oZwzQfFTHuKrjFLWrHIbS7K6vDd0am8xhCWHtphlSu
jAzVeg/SE9ZxhH5CLch2go3phHRNnySdIKK7KV2o9tKt4MRFxY6G73ZNx6wg0PpTQd+0O213HWnI
eCWWjfFCT7lzVonytP6ngl/9C4m0Osadycm2CvgNwRBz58NBEVyC4f23UqVV25kxyl8A2qEIm4Fj
JgCJiDyZsI2x3OIilBh2sjFmYJEnnm4ogVzYZoyfcjUvWN8YhGhJgpxg+s4gASPQIsC+sBfYXwS+
LI4BSAXcdTe8U69e4P3mScb0lz7OQibiMRZjNaP59X/tuc1Oo19EvGxRd7BdLuday0x970GZnA8+
MTOJvlbyjh83GbM6Klnp3tEi8IBqK/4HnR0+3c0QqreJs0ePVU21zOKZlVFNu4C2vuQmhCHcMQic
mQ+kZFhzWrI4U1o4OYFToLVJGJLleLBomiudEdx+GAjcB48eiZ2teLh0yyCnZw/gHtrJl0ngadRl
dR1/8tOgmJtl9j/YU3xdGh3LUJpfLcgRYghhS8nz5gNWeCFG/cciKODFgdngqa2r74whq9heqV1y
CTnTiMTRe9PpmzJ/GA5foshqmeQ0nFyJaXhs+hOrxfL5J7RysVQlDt33oVpCCtYgba/ZbgmEnpB2
X4amhAVe+QIGVIHlmEEPAuXDjZsrr1LhhMD10wt/jmsRrJDNjjnFnGn+uEtQ7POxretzCw7eKOox
CMJt7Zj2RZPb93Ed5D9FE2CsmfVLDLxNCDkjPqrOQvFNSPTtxiGEHdgDgw4mnIrUmDOGix873Fz1
j/RjsKnW3R2fgZ3ntJfuX7AInP/J7bTILEIMB6GzM2ciyLBXP5rdAD+OQapLZmmFYEwUheqqDtGD
FVp4CQE2eV1KBsVfT3OszE59pLhudfm34Q6QFtgnt5xpU3p74sd3XNKzCRtAZ0u9QUopwEyYSFlJ
YCCmPN72GTwHQAG53K48RAOTB9mwkvRXb1MOuiMrKhYb+5jIB0P1TSKP77ArMGrwEueaAiiJ4BGa
2QVs8MIqBQzdraivS9RW8jaMHGemAAMpDO5rsb9AofMK/wbMEDp/hSsQaGKd5zxHQMyf9CDVm/29
J6wUn7G6LlkmMO/uj4WJ6oGbe7SwKkseP8oFxMHUEG2TiYPe6STpsojtrwfHmQ1URacp5YC62ZfK
opi76NMdLZQT/FbUouizyAGgjW8BAuE7eR2a1hLyCi9bc6CSdAUyVmu3ULhgAn0qdnEiJFnMf5p1
QDfeqDH1sGRmg6Ee1gQ9fqBCRMF6nBOHvRcolZVHHtP6A4kAordV/EI9pJP1Bri0MOy8EfIFhUXM
yNOdmjXqxvAbNs4yjri8boUuKP4c8MRcfMLS3jTpDRDCj7GQT6P5km18N89D+eymXqGKTbFT96tL
krVI3NXGXMfgb/pSQqfpxHnGLDWlIU7lcZMTGckVJa9Z7+qjBbG34v3UO2Gql4oIU9RRyC01f80U
a//o0vwYrLED6dZowpXBlPgVHrtBoueSuRcVb81+kveh4sVkP2FAwaDtfVZS2bb2qAmHfHd1xYgy
+gpfd14lby2Z3KO387R5UPDUtJiLcXJP6wf7sdVYPKHx4HhO/m4Rd+MnwnlK9wX7PYnT/Y6iz+Eu
MV4V3gNEwID4OTGCfbeO0ipIFIhBS3leVdyDIlU+mBpSSNVhbdVgVxFAyZDYwjeUatRuvS4k3sIf
c6IIWfeoBMWGNcm0FQiP5T+mVZl1N9MdQwX83HFVk5/gC6AGzw3vNuBKgDnBGkyMSQw7shGMAlVz
BxuWb8LjOyhxtHDcN+wjpRDSecncn4hbWhqY9a2/7roLQ4c8OEcXKyIgB4chc+0xQhKt10KL5wJ2
m7YG/qTk91+mmE/OgbbCgGoNCUFFKupVlS8SJ7zSzfPph+GEO+r7wqbGdxYyLuTLNNGBUAXM9Cmn
mWPFL/MOZNciGC6F2jEYMLSV8+79uLwLc0Q0xs0lcGAxsdDQf3d/H74B31lYrWU2UlGHxdUZctRr
GdT6lTMnDo1rHfZkADPv/lO3mtbuW+DEYCKkbRV0w4T0VN/bzI8bn5oraRNqcYycDcIJfcyPH+hj
IE5kcoSHOzDV3Voe8raKl4RBPxfJNNrljALVKWrQZqoFjkcy52JL/2sr/W9FnppSHN/fsBbcbymJ
QfhvUqONLRToGzztbw3JWbfmEwCKCrnE1JpMMs02llv5OwocX4brCnK163OM6qCtDfbLCudsEPE5
TxxEto+xiu28w0I8VlefUlYxnU6GySbwMr0spHc0IgrpQLgPq/wJeVo1qOkD/7pvnUkcvnkih1tw
uc0uF5cnqIKLSaQsa7miO8Gv9iao2VF75oxepCkcfKFmXewjY8xfNfDJcH4X/6tc/Gq1oG8fkEnJ
4cWs/oQZDjOiWk4c1bniLq6qmaA0XHvQcmIJkBb3tUQPL59SRDm1gzGhN62e7OfkSQK5MsWbzT9Z
J4hZ+v4oAcvuumD0r0bPeGsaPeSBiMRATaqvpLnxeryC8SEhHf7f5mHXmDqnKClEMCiD65mPcAno
9eJ3XUq6oOk77vqxqHFWCnu/6GVRaCaP3Xwoxj/dwxg86n4afmEPKUXEhIICcOP7IFm1liz6Ecvj
2QORkcehiHOhKySYamVGKjiJ/jwJJdyYIQ+sAi/0XOlh+CPEo4HIZQOvJFZddqJe8yBVwyPFCCgi
I4vgrAz7HM1wVHum7VCpL35boyGgVBjsfBxRl8ns+vfxvGhDvApaeqe9nwdy06ugN11p7xKgU/dj
PaNa/+b5XuN1/QjGUYELl3U72oVi0VTkFVbYDLnrgbfOIEri2LJPCayWtdNjIFyebtnzH508mr3C
OFnqJl5rYdMLObE6kGxjdJg8ifV5ItFz4vrFkyBY1e153Kl0ivruKDUR0au6GjGCE84O5ua7ls/Y
VfVuctcnKhHDImDPkNhEAfnlJ3ZTTuQ0QkXU92UbKBN5Xm2AKR9bNM/R4aLH60WsuhWckqvUS/Ql
q5cAoBh0Aan7i8A4GXzowWq642Q1cAWSKxHdX6AzlGtV5m6iJjlB1WNkwBPq56kwEagKNm4ze3y/
Z3gvY5rC2ckcHZK1XMlDAF53fhOMAy0AFIGAGzXUOW7Kr8sYwhs4LNd2vv/YZojf2QhcYYMMwx08
SSAUyd+1/9e+conyff2A9n5Vb3dmkTDldobmUoMJTdaUPJpbVKsQ+suSuas+T5hgRP9msRkayLBl
eP6elAbiZjKSfTzBoP6fQdQfPjzqQ1W3T0oBxS//HDPtu4Bmwz7H0j2Bf+R05AGxEap4q5cwSAZW
A1qRO/kGy6nCxp8sCI8VCBFxI/Hn4tPixjqNImH2+uF9YajwYzbNEQ7Z78TJZh6LqokUkeDttuph
MVCSVDeXSp82ZCYp2ZJesMtJIyHDKdWWjOAypuIlbQaK8lJ4T8X+J8oBE65gCv/RllOZqAJlzWk8
J30Zmkfs+firHAkdngC5qgHp3dZa9bhoVPT3DvETbkL3WDN8Q/gq3hRONDB6gk4PSLVpvft68AFE
jtLk0DRweTAz2vZxOARbrvAvJf5c3Lns+BmqT2wKJbeM4RgZ9fHbD+4JvDnaeDntyz+FaoQmYoB8
K+DBaX9PuO+lSgayIB981Jqegt7pT6TbESz4ZPG3ncHJLKKx0HtonVqzUOMaS5jaARaiEGz16+En
afmB0cJbx0WbT2pClRafGFxZHxZvhAG6xbpqEOG22JxIDVZqkhv7pEdsQsjwjmfcm8pgELcLmHFh
ecfBng9LEcoZFC5W9EloJcxNuomm5uLF5nHpbTi7c8S3+Z3XwaGW1wC5/K9Dh64icqBwgaluy4zG
PXyiaYlsXtCrzI2U8VVXCzw8J9O7wsydVjCgvU1Q2Dw6LATc9iVFEwwd0i/iyEimM/975CEenWKg
dfI4MS/PIjFEEsnArnxGfT8fRuZvcSyvGPtGTwlPG524gQ5siArnUYSiEz8ZLGIz5ggh8sWLfi0t
XDGhvSxly6nA3BjMstpsMxGZ/MuLyJUTbamqHXImTM2kDD7rJ2+7Sq2rkhXJEUHV6aONmqVl/Sv4
NbyLlzOjnAXV5OItIYhNYVZqNFixPTX7C769GTdohAi9auU8ZrtAzdZRGsqGo59G1mEcuBzzu22E
wCjtTUqZnJebxSU7+B+V12f+mgdcAHNTZY0RXIMWenWB1I6y8MZ8/1C+IuLsyL1zGFgd6kZvXZCz
8hv7FLNR4WC5JfpduOJHC0Z2eFwxVu/iyBZRhc22xl1RIqspVk3rX3o1Iu6lWpHK8SQkUM7pAOV3
j6qCAHIlSLp6H3z2OTbZSsDzh99Bn/XtV9Ou1xR5sz1gCDkc0pEq7BjYTajNBR4avaRTternnsy1
Aq8FpDtR/RPY3g041ARXgYTlKcTGqXhdQiaZi/EvM/pOfrmqGnW7Ae6UJR0PoB2Er70HoXLo6bmA
5vVT3fbJRSpRy/4AjUcO2RPfclJ5ZWOnJFE7cFSIg9uXWAfxXUaSeczoWff/QGSuQ2dmkUKO+tny
NPwrjDlsB0mcUP+kdhwVaWNSezvoJ24qfZlzqh7U2LqHETjS7wpTaK1pK/Y5kcZu9brqgO6DmpGN
9nmnvd2S8C3UOBiXYQQAmIgydGN4AdFNzUq1ea4SqZiX8qj7ndndiOYWwO3YspJ2+8PkR9W19qPi
dwprqxsF3p0OLDIlvxSXlRaoq6X13o1CjzFDNLDwNtbmNG+j0f8fYzwP0VUFphayxp80i7nZq/gp
QYO9oZj6QM19Dv6A/wbHFOKH0A98vtqVIlgQQuQbDecHE9dUtJ9yqfmHkoT4V5SI0IeCotpoxJeW
RX81O3CzvXhVgmAQ12pEx5FmpwUgg+Ak9dGyuOls1xToTzKuwHa84TPii7oWpHonza40Yy1N6EE4
gn9dg2Bv99bHyLwc8h48wNhiHIz83kTeTDZOMK+IW3kNCR/Rw6Jj0Q5ecSd3ubsW41ssOSxNhMIp
LBLqtpIHk0SyXY/x1YZhfjQGjPb/ICI1B6EWOp26w1O8+YBAxgpedbUfZ60YUMmTaJVq0jujPpp6
UR3YULgYuQ+IXgH49R1JxNGnfcXr/vyjjOX8z51ILCuAc8VB8+QVYvEcZGZ5bq/fhDnosi4X4Bsj
jEo742ju6gxztTRL2z1qep9q35+grMxYzOFqsfP+Whf+kb1LZJKm5EYlP+K7jvSwqfn/erktXje3
SeZMZwRhwB9ovsf3LQHtjk1/8nFmc9Qv2G2Elgo40e9h6YToCl5zfv64eZ3e8U0UF/FzqnHLKiKi
MULexTzAutyQNzYuNEEuiFH3moHqyTO9fTQns1sJtjVVKwVF6MBkWGTkyrj9cdp1/umvQ2MMn8ET
Y5fzQHXcuuXsP+ZZ7ZIr1sYH8Re2L86UZV4tjDGyKbpPpej6Tytl4D94l210iTWMTkHrvnrU8mh0
kqxZ55O6G86LLmFTtmV8qWnrO1XaCINQPzVAKvkg63h8SNQpJEfWG3Z4QVLQe7DBEIZuZymn6Mbu
glkO0gUULkXZLcyNhXfnxppP2euxuISlnyanpouVygINWxv6F5TzSAw4Pe1Z+TerwF6VlmNKfie1
W6+CAWcHD1quwirWYN/w61XGLHSXzfU43f+3ymcavF6QM7NUqWbTz2eyURcQQBZMODUbbt2iBwbp
4NGQ04uu+MzT0tG44I8ui5oF2En/sM3e06FAOCuHw2K1DnhKiystaJd++0OGO0i2vpDi/Ylxsuwy
fthmjfrvb8wgWCuKzh9E7SG6GGiBroYrCHRHH6TFuEf61labZawaTK8wMDy9X+ehOsOFwT7Cu9XQ
uBB+ymmdJyWzK61hT0nyApppe9f/zQsPYaX8N4n+l4UGKQ4qTdVJcqJQrrDPlQXvva15tzhX0gr0
Bub0kk+hbjax36+U68YdKE0l4i7GTg62ByjVzeerlj5qA39IweylVNvy8/NDMAr9jndKtl2gQrSC
2ZSuV7HCHqkAx6xVmyKYKKJgCl+bKJsL5eKqKaSiaJMVlHG2jWd+uVaTckFfxStWHQuAguQCytjR
xmTfjFmnCyY6tEVg+iSSO/4ZcD0fZ7nknfQQSybrRSNpwc8wAnOZ22qg9sEBuv3L4iHivl6VeaNY
cAQah/Yn82PX+jR4Z1OG9OEwlNyrMTsUtKfgrol8bxGQxKKjJ2hC/yn0OEDbaYTlUox7Wh+j2GB+
zUjvoIX5+vWzm2GQ8DVO/fT+7zdwcmclFAOSjdW6sAiNOTn3ZtBe3GAFb7YbI7y3FLeZ5s/X6qF4
vcMTv03d05kc8kPgL+ydSI31Ai+MRu9MjE1Q0ZnEQjyhctGlRDAXyj2RsTa+XpPkYYC9YXwEm0nv
fzdeeGaeJ+KJIjFchF8uCal/yxVUukiBdybvm7RVCPfp87x9ps/i1aOkWIWyaR/MNo6R5CVDsIOm
k+dc8sMh1JOgXryBX/GNV8YyNC5wJ9uxc41h4j7Dvg/U5UkCOPLNLYddC/vZeXbRjN629PDIH/Wv
0dGLTW21IfT3WtUibu/4QqVH26fnZQ+cPVafSgSzuey1/IVEnXbXjCKzajxebtvjwnSyPhIFZUyl
PWl7/uG/ce/OUl5c2PaZTro9yWlKTLR/1DvJlKSGNfRmgNk1YnhK558SI/DMYw0N6UR0XwWi82TD
bONbJkWNm3AGcjYcba/wSCI5awWqopxQ/UHGezBwIHKpSWNP3Amqw75346FvadZB4PTm1D5BdyNk
W5Fw7fjj52XNSPSBwJvzNFxpS29cKd38SCH43b1FwmSKhnClIgjV1Q024ZNXH03Vb3X7H6nTEhfU
CSPMII6Pe1MVIVTQyGChG6ISDquocQbMMh9fdnN5AbaXFIki3lFdxTVVIlNeo9blr6VZ4n/WMDUq
6dRUSl911YcwLDbaDniPOSt/9a9a0qSvW7PqUUyvanEwdJh5/A11wfAUT3qaXFF4vtd8uaIb/Ex+
WkrNZiJ8TRcWmpEdMd5D9n9Hxc6RPiu7yYnNy7+mmOUQWghs0M6ccFg5D8MR62NXtSOp16sCXrW/
YCvCZRoeJ0Slvfusmw93mXnJPTWQtNtczfS7f/1cqBWL7ghse3BzxL6nxYNjo7M2W5Tz6HFtp7/6
Q90or1UoWvFYdDbXRib9x61eG9IDsU56GfWQwQ1Jxk6JuYfZpY0YV21Aor8XaH3XYJKq626uq6Zz
GT2puMVaMagVgLr/8y4U32NMXtGAx9lOUPwONqZys8DiA9K3YVU/0qJseISrn1CsVz6iSLhXMf++
WyX9EYN3lk2NaQBSkUCNCzUgVR9MSVQ+NX/yFpyGokFpMXPDleZZVyKQui7lmvs2PhTB9T+EIVeU
2pKb1yVoa3v1336gPgj1qbkfASZ+H8qv3zlalLcthb45XTInMlCac99Ss2bdf5RfvwV6sJA1dpST
ZOKTJ88Zwe7+Gqayxfy5NC8L1urVEaLdzBddbD/Zr/FRxLSNYHxG1fC6Dd1FjHxROlFNiKfVYLgk
NnE65easgQmoq2F01pGdsKR7ZntqCCIDaxUXRhPk3xtNJr924lvkx2iyVj1Sy4oPvbQaz1xrgLOC
0uPyrJ/Bypa7DqtwAk+ybfAeK0k2GPrjdZRLeTCevf7kAsogXA6/HGVzRsREGstyqO1FgOxJR5ll
RXVnGgSt5NarjwSq6qMYpaVGTv/hYPUnGGRf6uGrVziEf53ZoFUFt6R9xuOmhs6h9T/2qhofGoHA
rX765o1R0/ChQUGpizfEQpvFbFDoE9cuN1F9hIZLKESydJ8TIHTTDRhboI7pkj0jS//awPApV6gl
EznMkK5Cji9TE1MRW18OJMNtmA4ZDiEkCDOlJWpTYo0hShJzI+M6pLng3Grixf98mmx5xzaf9P70
wJ5gnk+MHYEMA6Jzw0Kw4LlZ9fMzvLcyhY0rVR8Vliz0kIhbqUbD5Itg3U51oOuu+nCExo7TXfyD
HoLeqhncNsDIAhqZm1NDY+nBkNjlcEHCIanxOsSM5e1LNS2fL01O0u1pIR05zySjlL8GYJqShHy/
AE5FiivpNFZJcd5C+Boy2PeAB4NrJTwbNUuQ3wzCz8K9Xq4fDeMue9+oYnUBTyagZdbI3SBp2bua
R7uUanBBGgQ9FYZzHpf8lNoSSnEcv1gGcPSSffAAhLGO2BFVlwzJZ5YX6EeHfN7i3L76KO8NvzZ4
BXrmZeEha4wy8ypUiPggMowVVS2a5XvmuNP0/oGBkMZ2IJNUk5gtf8CMb3ByaOsLOT9HznhOZyO3
kSGcKY2I+X5UmEi7dLu6C65ooIKsBHlg8S8vOqP3EnFCZduF89g/Yt6pHzOnPi5N5gEeNikdYnOi
93ylaXOODc05fR0c68qAoR+xFnU3IVoICAy+qwxFfETPHTdbTX79eHCnfP5OD/YXMTjmw1Ka2lTd
q1uq8WQWX0iTu2aRKtoNox9dZiRaah6HTePLeSJegaSzHaQ6FVVUVjbBq+RrBvDZkYpGZCfv/Iqm
eKEkifTFwrtIQvKEK3WpmR1mbooIaJzzF2tottvosCZ9Cx0retOqmyai81z9aJJ8Adgn07/C7XC+
Wf2znZ25YGeg4bpz29LTCscE1LjafvzIBnHl04cgL2MnbzBsY1hiK0XZ/mNnVPaTq1b9iIfsZFDT
zoT+4X5KYSucgJE29Qm/WchwzMZzmCbVRvQQv3L+8/4/7lsiVJ9AjgspsHZx7yPUiQhBXTyM/KmN
k+Hte5p8AIbVdIt50IB6ci9rkv5/nJ/hK7lh3wJRm9nMYzTpebZAxmrpOb1IzcQppykCCz90T5sV
AtHDh2q4xdtJmGp3hqwpk7vXdkGam7qfBbg+gRRsZUJWN4zBR5Ay2In4UVdnXc/boQIYoLmXLv7W
Eb5JGiigfgFdITj3EQ1eRc/t+ctHUwuf7Xt9aCDHBEI6mqxZrhXtXZInJDV8hGD+iVDqZVt9v9WG
eFYp2VZRc92IsZ3xrlmMejMVnlcp8bjmgLTAWt/mNHDOGA16VqmOwmTKDDsiQaaYYcOES0VTnufa
vabzkUmSnf+bvxRJefrVb6Bn6yZHRlEgwpqMDcxh3DQBNjF0HWgfMEW9m2rN6r4rn5IkdE2rWIGD
a5zdxL5NShOpxB6SbNLqdD+9qzut2uKjARPr754Jj5GUmVsOgW9WOwCJC9zG4rivN1UP3GMeWpz0
6ZuyUJIythpf4UDKJmZFMPGUAB5W+g3tTVnsarvwps27QDqdoc6IKtr9XpQysG4oXdhp9lrgcFWa
he/txiW7OAPPMlsVd/bFEeQ2YglFqtOHSwRcleaJiuOrNBdVClcB09bZVyJRRqts0z3g/A2yN15j
Jl3kcpGmxaod8IfHrmtY5JrGYVR16DqXJS5UItDEZMnenMCyIuFjEdQYzFdh6oXoPrbZMjFYNZDt
SxYnAeWPCMRMDwTOTOmRad/Jlp1Bj0LU+i6/bec9+oo2cBl3vwfLOCdUHCBP1tHyGrjCL3DdIoOT
dy379IUtREMEZYLOcoaeVPHUTl9By3qpnpH7+b7gHS/r0Or27IMy1XFb/3AiPsWUJbtmIX0M4enT
ENTNivXuFI/G1LYx2kUYjRh02xjaZx2uJHZPClYlb0WZxyJ0ecGJK5BQZ9bxR/WcHFdnEurqEu87
Msm8LKIHDgbGvvZEqF5vSnHy2FEpi52jX5J6LVnlh9ke8r1GA8HZ3uTV5dBj1332JqbkUDetnsib
n1WOYOG59DbKtQsByMBu4/nu2Yik058ht2REYqHGN98l7KlOeU8CG+J5fX5mIaoe+er6p93LcIYf
X8aWFd8g2Kwt24KkNlOI55AJwfkMsUqqoiPUT8IyBevko9u+MPYoskeOQenSFCqBd3+c0QznQTnK
sm7d4CPv8EQ5hN01VScLl9Xyzj2tluYl8AVKF7ju5XmleQmXwb7adlp6MkwVCVheSlUloULEqsV+
/fyVcmUV/sshXNVo45Jeo33GE+pFIM0JBlb6PKAbflh1ioYJjcco9AJz0NJYRevYvpCBY5o0N0Ih
6XXl7Otocfwws5wCbyqFAYUCToZ8FinBoHypwTUXhmUngIBJ8eHkhOsBdOAS9V9+Jd5z2Sr6UkvT
zK0vw6gBeiEgtXJsbPyGsrR3albuAzeUq8+ZwCHqgV1wW2RepR4Eu4Z9wXZmMwp5gWh3/x12TT0V
bwxBAebyHqrH48r1QRoAqtGlwl4GtGDhEKjJQ/I9ZhlOtU8yMQ+ocC6ONW+qukNy8pCjYLTdgCaF
Lt9v3NCVd1BmaBnEDfvZ/69zVsofAcvhpmZmcmq/gRLHijUcqqnZGRkbg1yYv2VfgOmBakEZJuyu
4r+hLbgqLip7h9Qa0q4YMbVfnbfY5LH7OFot8eGaxYQWf91M5znTUug+vY69rS3dfulbDIQ1g+19
ffAHW3x1BCw7MiGS340072lUPW7KqW+dm2AIYWjq/vt4uAxmNeZdgYRHidHpK2Lpu7GAKAY2WF4p
dlgBujKqKhhEolKVEFjNSwyhVBn80yngkpOJmk5lJoylO7nLiSuaI6WT1ZPioIMOt7H6RSGGs5ni
gADoUBHzliOIsE6fOz2GQmVj9+x+w8S2o43R/243tMtGGAY7Rxd7vVFZHMlPWeMggV/qzfIdatCw
bY6a86nzR4WLsA+qwaLNgFPSa7rR8V3PpkYQ4JDTxbrScHROihPk3Gpvor8DdBvZEONSUqCpOju5
hnQDXgDzUNINzk5x1UtBciQlsihMOxSLNMp2RbUl8IzoZz9Bf+oe2wUl2yM+APzO8hvSVcIbN2bx
lAtGDSQp/EcripqhF0zJ9aiP4fo0Ckda6XEO4PgSz6ioJpAGQ+d1Za2kCTtIiDIxtxZwq2ml8Tav
jgBclGnFsAx++4Cf8SW++ctuFqFH1ze0YQGPINclr25Gg69MfWUaMIbx7iiops7MYskmwygRqHK5
EMIJPdtjSOcGWYDD3OLVzU5eq+j0JNWdPnpXcgMXwLTTsdgvEWLo1zexVBbJUH0PBlGqbp12Cs1J
cCMiVw/GnCm/LvwjC7iQpREAmZ6GMeZO2P93n0R2MBxgD/roJRIgSaVZsjEqF44txBxs8c1Hw+OO
BzgKKHhHdzauydh3AOOiFR1r6l4JYxHy5I0Ve8+zQV1HiPPqQJ3wU2srPfKuvgXPz4hnTK8OA42a
Pd6sdKdBhMHNmP1IwTvk9+qMkGZdh+sM5IdIF7gq+VRYm5OyA5sxqlkIYn9HC8k/m1hkePtIEDmM
1OqDptXXp9ICNw0nKB8E8OWrinocDNC849YoF8aBNUGcWGOitsAs/yLVP1ZmDMhNgkCGUwQY0v3t
T1PLd3xceVQy2+M3iuEt0YX/njOOUYK8MmALK9MbqSWIZFdJyLLbCQcTp9lmx6ACj9t0WojsoVrv
TVCiKlhJqX8Yfl9Sx5xDVliSvDQkvpo8Y3pw2LWH6kmdymgOworkjn+iXH1W4rRJK00BQyJpWBwV
Q9Q3YHaKh2L2iHDGFEzsPQiZ3nzFt/5NQawJEDH/NkmsIeq9BwtwH3cVTGq9DdWtW5dXjGtqMpRx
lMTGguqM/AltUbkiAxQU0uuBYu2FTMEs6Fkm5ZbNGe7m3CCb93PW55WE4QsfjDxB71zfBd/MGLd3
2xDH1qs4hpv0Mj+sA/KI5cHMdwBrxW1fFlxw+SqdwqbHNcVpJjwJ2JKSE1LB4SqqsFhI2eVZQBQp
5WUIQpO/b+yQec/wvzusZ4jFxRnVIFfpq2Q5WDwFJiP76m8AlzD//PUNNJ/ZdMyR9Uwq4i/DTf4R
qaGIJBOXguacEFWxEzSa0lxivsrAEEMSn0b/wVCcfKEU/SxOHgMhBzc4PtVE6vvTTyTS702gJNaD
hx8iZwwlgmcbl+EhgJsKRoKf46V+VLHU5dIYSY71MxiJ+9AjNmKEjVXOfjOSE+BTFAhypFU69mvi
lWMMO4+o3fm3MJwOkpzLkBSuXhLwbUYb6H4eLWrQAoGPyunYewixuX1KyUy+5tGc4wZ3DWSSXIya
y4UJhIPZYAIv1OVsB9GkZ2ZbmomzBFZmcISSDLgHP6tenVRhEzdJUcgh0yxExu0SuXkV3TDdk9ad
lv3w/dEipAGKXsiZDelbsHYRDCvsHxjk1swbEOzCImYvbUi2V9BaSPmUM3429GVDkF4YiCC1mrR8
dp1XcdCkjtwFv9H8J2L86wSXPUTB3NaIpRM3fkFP+cqQNqRwtDOF3Z2MpI9glCr0Kcp4YlWk4FAu
34qhVN6VZjZvDKif0i01yNpKqZb16/00x1CFBLf5JfKy13IYxLm7ysizoBJ+m5KKZA5z/hFYfpVS
iEMbcFhDmnjex0206gucaZGS0x0R/ZTtJYbqfuCkv3/mwgP5IvrL3k1Smlqzd/tSRCI2zZOxKEPF
HDezoFmmeevjF8X8YppJAx5LCrx0wxPxOO93z6/fRPn5jaGnZ63lXlNELuMYD8OOiq/GDFk1zPgH
YbmGNFj3GcHLMGFAfnVuXo6oi6IwYHQ8QMrs55JG1en++e0QW3lwOx4Bb881rUvzdkf1oJ7q8oCg
ohOlL7Ihq+Qe3UluAJCXiToonnDfthvkJoFBBrN1VkHQ5406TzSAr9LXfzO49GMYrvBc0G9e/WD/
YEj/OqCM2AKvUYNMUt15vRs/Q8pI7HDatN2wTZFC7+M6qoTH6VHbkaqIJhjqKYIoZymgKwV2GQZb
sD1jZliCvwdIjuoWhDvb8xzpLxkJNCtAVJfr3ocFMz2XXZK2PDWD5Tx9zKsKYzYhxvSbW7ry1LKx
GevEgM5PXxQCP81SfyY7VXEBbwCZrbHmVQMppOcGrJbLJRFIssUy/FfJjDWabxx/QTTCQY0zp2fS
Jz7WW35MI+NdJWa2oB7McqSP768T37yoqe5GeU9xxbMQGdQYqCv1z2s238xqlLAeyq54MjcigYKP
oJXJV2lTyowY4BVIbLUTdY6i6F7kv2hgL94KuylvnsUkYwbP48deuG6zjxMwLYmkfs91O2SjbiSy
koeYD7TX2mb6QzsneL2EBAM8TpDgcZdUC+tg7M9/NwaThUlIlyqkw5t66av5rQftJ+Dbjswb3orN
gisDuFHMlkPkgzNHhvxBCRPG1IbV6OI1vf2BoAD57ipA//KLAxdv7eYvOVI1lm+Pz+GY5Vbf3Iwl
j0Fc92Fss2vO9IEvRJbiHi2JtsFCLpylwiHn6KUitT8BLwphXX6wJH6ZOGz+iGJS7mvB+j1cJDQu
51AGXCXsk5PmR+gWGr+v+6YiDhwJXGlFlvScXdlY2q0aXn2oklD1Zry/tlHNkXCAzjQEuubG6UwC
9kLVG/AtUp5/EtFGD8BNuihqxH73VzOm38yeC1wawVExTxTR9Rj/y/TrWUbkh8I3xLqX/O5P/sew
jLS+PZUyqmCeZw96+q3fVmIjfNV1n7foBmvJm+HMDkdLMge9yNEqgf9Z9YHbupOkraOOGGyJLLed
wd0y4tG8X9wExXTZ0kbLoCyQ8jsCnccEmby+V/Pv8savDN+6YEI07pNPaDoGD5/2eei18YqgD/z6
oB94M07kATYki92oAHHm9gtMgECwcZ7bediHdQqiK4LksHO0pKYM4qjd6r0BZzKlKBbB9FG3+sYr
Y4ySo8tiDImCeNjoMbP27bg3SaQkSHsUTgQwA7RhsLtUo2Bkn+Ip0zpkng0KBkgIhNs6mC/RBqO5
GS86tN/652SZ2s24mN3otUphtlKrwclkqEyZMax9ZIMtcS2x8meKURJoTRtvczRUo804WWjwCSB0
Tj+ws3y+zt1W7E//yTtyF72hxo9gT1Gp0PE5hm33DVp3jbHDorK8Ro6FR//7TXy3m6ew1ekZABWv
ee84RtP9di6tyR8HfXS2rMe3wpUCOB+uhmMeQ6+pXlMumsS6ocGvY1qkMyGCFauW7cpuai6BNC3/
iaaQ4Wh0lMpsU47zJi9g0ZAIzfiMKYAzRvxGclieXki9ZlXndmSIx5XMcMbSv2amZADFs1pii9VT
+mglYW7o5I4607H/sqpb6vR6rQoYQOjq38i5r8QzW2qt7OEPFMMWxoE68WLvEm/l1aZnKjTcO0/u
Nv72quQnqoc3qj241/oLr9hUKJqacSEjHBFmflgr/lnF+QeJEFnYKR1FnGpmKiCFNCRwVfVd03F2
2ek1pNJRHQpxdhQegphyTG5Y56BhPhCVlyJSlfDFaqzIV/cZ3xb2djsb+150p2D+QtBeVaahmx/p
UJ3m1AfeI7tVi3b8tJSu3urvylP1tS+ZW0KA0vVNmUlcWn0qKtnYMji9+qiLLGpGr6YKM+YFEo9+
HFpL5Ae3m9fbU1o8++ui6wphOwZpzknMRDS8w+SRuyBDgt+/3MYsW8Pil7zyWQTh2O49k6pP8Ehl
Ze3Cq2G/PwS5yl8aG8C5zg93fWa14nqpAYwl9zWxgcYpwHHxviXGrjdiFcRtV4MLZFLaavy0Oi7N
dZYynzunuDMJsdJq7FL14fooZkEJrwffZRu0sz66CVj0jo8EehwFOSE2znG/3JyXu7x4fkZiCFRa
hIYK7EvgLYX4hWpBtHqNgENOxVD/7l+DU4blBD3triMidnLEM7ISt38+VILmhwrXM3577Oodjnf/
le7jspAg5mnJF3rPtMMYUohPqYJWl9g5t2029G68/uGzTImHNnHFB5HwIHwJ3l99lxXJUg3pyWmk
fJakzhewiVbjkTd4mqI/nqOLazA2cD/rC0Pgw6xWUkdsscpfLv5HFM4U6Z8U4ZXngO5hV/WihXB+
7OrTfHr30XLNl6vt1+CUpnGwWRb28/y46K+Ir6qtSVg08jxNaTq63+1kWJ6o/IUcalfQlzeNnveF
ez0As/Io2tIcppkfsv8/EyH+IKNTEaySI0a0El6dScZAvKb0Wfye8nQ3OLvaGCFOtCuGnzgaVqNJ
BhQOIGAGXioB2RvhdHTYH/oAcC86nwGHpYkY7CiN93bGUQ4s9XorciKWCtPouy2SWEGwR5yAs87N
NnTk1P1n9TrZzsTg1olFv/i7lWoU2NHZugyvplNA2jRA3gQa25Z3V16r6XOj4r8iuPic9bGQ5hh6
EW7b2pdjgn9iXUzIzCOBnzui7A0E6CFGMzvs324DEysHIeuaNi1xpeA0lZjMt7+ifDiSaqidyFJg
I2VLeCBThnG7ZIjPbBC7QH4v8Uvdwy5OT1vxkTlBwrucXdNex3QvwffdRKVGxuSwio3caYVqkhoD
a76JVAHl9g9YoIuzeMr7qQvGb/NiUzl+XIc2yNdgLGtMfZypYEGWcHdmOjcYCu2Y1f0gxEeVgLPg
FGVGexBZ2BT2y7cAlizDG9MCdee2x0hS4IUFeCo8JswFJdbFWO62R03TjQrOqxt7TgAUdZzMbX6B
VoZil8/CbIm80d5ZnD9O+RSuSiemBwv/vnKPy74djESK6VNoc0Ds1qPLP4rComXw+bGti4gwzWmp
J/DfrpqGIiDyNDK4CxtzzWyk4O26wsXV0Rj//8CCB3JF1yDVKMuguTNU+WwCsZJi3Ara7RIxBoT8
YwahVQ7NZqq4BaIWyOyJ+rKkA4jwdVxjs8RfOahYppqjcwmXPq+2AAicN1I2ICwiUTFiUF8Dafk5
Kn8rNa1H9B3Ibpobc1n/79xe25oJC5G0gVO193EzcIAQ9HuiFTIAgSo2nV/oLB7ddAYggKYkZ556
uhx1YOd5E+2kaDaTZBrJEoWEQTDGfBiE5LnfuupU8TEQTaaQBbnuypRnoWmAaXJtBDhYBx/0UWYj
XREu2RD/Ye8S5uukmDy9H09K+qH6bRX/ygi6iB6UidJ5MBgDnZ7UR7FJn7puUPYSAXgRzG/jHr75
XBBTf7Fd3rudenY6D3jtnl+Fe0O0XQRn3vqaQ+pKdnLGoa94vsI1N/rOWv+DPH5BLKI6qSGcRCHJ
YmuiKhs28u1t6A4gF6K9H0ZqfDcWl0IeXb74jYzVsurPwUYLilnihSd4YSpSrfFRBahOZ6R7xiUY
omQ17ZGDRwolbCcXWVcJJkNHVpSKTgcTmM03Rv1soS7P9Shyqp4tY7IZOwcLqw6dOQ0uqap0dnUv
2di55k9GGv1UJqlwsSfusk6xhlyETk3fuW0MEzsyDC/7sTlXV4N0OJ3kfdhNlIFaA4td4lzJ7EH1
X+zmbssQitGPfIgwyFsEvMIn8zoUr9joCWMtNPN61zlIGT8dxVDudWjrtlMlY3oODa67kONIl6Z+
ZBXTa19+XjKaIFih0bHqkqSotERiug3pU0NSIVahSc/KsWoLD0LlxxvykLPKMYcSspC4OP4HUnaz
JLzUCWiE3wdFlFo/LkojS6YOUQ7XjEaxArp9j+PlLlEUDmEMRvwP41XZZcjv3pdXQxiEp2GbS0wB
Mv5Qz8RhBuiRMiCxHNOWvEqQ3/Q1580vgCTW6uNv6lw+lQTH8THKstsi2y7vKuW39ej8Yo1xruSL
riIZ2BGmCnqLce3+dGqurF7Ro2X7YyEPT1Jf7PYb10duYbj0TSUQXEtqkwxat+7hsBGm+bRTtvDH
SpL3An9xmiJwMtuPn2nGq0P35CfKV9tVl7Wgc4yVKL+zn7VLTsCRg9nfo0STGH7zjoKuw/zBR6PZ
9RZ61IRC4xe49ns/7xatchZrovBrlm3uykHC9JGlfuuFj/xRLUJaFmBV7h+Qm47FGSi4iRHwUNIv
k4kxF0/Z1ts4TOL9loSWGtqIRCuDcm85S3UhRDGMF6dhVWQudWwb9dGNDiYB1zTHKjZVrzEM8T87
FyU4DR2Qi6WJtvHcEx24dBdDPvDoFFj21UeksV1P1q1a+rPrQtwd4gghuvZUds6iHX7zQZeq87CR
CKU/tKkKmFoiQEi7K4opLJl2k2XJQbYruggKasfqhcPZ7jrDpodA08M0hCkIho3I5I2JFXW0/gk1
zt6/g+bqJZ5p0zlPMb2oOYkdRN7hrolza+lup8SK79l29mahWa0KUThm/IFcoGpaTWJwEJ9P42NL
74unQOLISVfTqeaq5a0jPfzo72zYvboPhzTu89eNkUq0gra141X34NpDfT8hM5rc3X60bvvBdFwv
btxPQnzB1GhEq9SJ8aG0GYr6A83D0L0ulpUWcDQA2P9GD5FWNWcheUaMjjwXTVTee1IeCryJ2f7v
3vKXoKEAyTKRQUEKc00kDrlcXK0h7axZLKqBZtYYnpfxSiHR4zm3Nhm8pu1+LT95NWLZVl8KDtyD
E2YLz6wLgZyUp9gpXZ/Okm5ydR2NkGX8CN19NcJ9MCi3EnzZkp3k4qE8S0jy7M+Hzk3vWhIOsXs0
49Bn/ocGWBWTkplGinoI93eECtNmltzne/THtQQimtnzyiFGnjV5z3yomLxCDGWNKfiIHH42hXVy
3iV505Hco6WeIXWV4L1vUtXEFvAxWl5S+4oEajd+gcqbZg13ydVnVTA8qx0kb5K+UNQXwYtYxcGM
UKOooYSuO4VWLypDvlvim269RuhQxfRw6+r9SAMv0JpZGYXk5N2OyLdE1Jl1afiKKx2PsNmWv3v7
plnMjUDMaxROFaLGogzS1TqzzeApXVy02u53YnCOdc09oWICazs5N3q2SRB8jr30lhhpI85G0q4g
n/wgV7iL9ek+vW844vgeKt0QtvEbO9zXsReqV/omWdxrfymZbKCJtjYdGGamISudM40RYh0Ac9YI
21EBDaBgGzGCQMzndhWQL/HJj4iAApokw6bVo8abhtJRM0A2pfHd+awloA1fFiCuuvKzZoAERElW
n9kCRy5aXJseDW6Fxl8S3LDoqqrGkejyuRnwp2LQPdysblcX5HEKJ734Nb4K6Hqz97ZHYEXq7iaI
GRlg+G0185KTnMhaB98TEWqkxoy1CxquBnxFnuUEur7lmGtb01FegocqxZHDkcA21YV8UP/iQ75k
Kp53xtX/JmcVoVLb3voHWx+TWXWcx02hQcpZRTbaVH1HGVprZ2pY6ilsYJ8T4stZRCb71zCXnLkA
irh0ckQfLl7I02BPMD5YpOj5aDOD8AfxQnKQxhDdxElgZ6cMg0Eh2o96mTKa1LP9FuHWfBjZoXWi
DL4Qo8n8QkF6VdIXyboqgXAy3g2bl7xlp47SY3TAuwC8rzGCi9QcA58tiqvyKYzJ1NUezWCSn32S
kWZOADUYVvASyQUHKJRUqS48VVM2MpaxndMtRCOMMROtw4OYFcfyPP1uLUn2sgdCoyl2rmVyYwRg
vMFIKVD0uh4z5cbjCu+4+YLLScwcXwBwu2iB1cLjI3GSbylfzk839FFRwslF4wFtPFn1GaZovfMj
LrpZ6ZteYwKgAc1CT2MeYGEVd1qM81tSLVsOXEFyx/L1351pthhKee5ZYnGzFied80sy+dT2iLeb
Bj2A2Nv2uxDxgoSOL6o56x540PDlBmaFN2SWEdLKz8u/7Gayzw8cY5ygMlgeedSe6DNntEG2ZiWk
tJ4SIFWET6psTcG712XUXg0quw3D9rmolvmsbVv5Yog783njQ7sT3j94yWsg8J0b492CSUgCM8kh
m/DFgtk4xScexFfgGc+kzPEwgZe8epRzGpVpudCdSwEVkWhEHaJKwzs/zu4HYUWqN5BlI8v/zCLt
5gKX/UXNRkduIhn4Kls3xTASteyBXW0pSSGMTU+YfGsy4RxJ5Zg22PhEB/8YsF0HXEv2e4If5CtO
Sk4J/5IF8Q9GYtkdfHfxZJV7cPf6pFsO803/2iJR9Jrh4eSyULj7Ek/Lo3RdsMsXAXvp8Kzl1E7p
HefCOqeqFEd7pO0dLLfuf/aecpggJzIr+X4WNiwful7Z2FlXarB5TN8CNB/jOy4oKbWuwHDdwKDZ
gRQjZ5cCEYB3TPEWve9kVSHIxyKyKXp/zh2+7KgyLbX3ppTi7T+w5MdSjwwVFavtqpLY3zCs9/n8
cDGK4TJW0p7yBrc6DdgAB1K4M7tSgI8HSiMZVbAk1ruT5KaCzyhbPm9iokehKJ+M/69dR9PwofWt
Ac3FRZKYaN7E61elRsNlQMKIofv5Jfw2NJo476snhKvI6dzyudeSlXcxW1LY5RQBOuyhQq/mJXeu
XFOr8g7wDsSBgh1bInILfwRiLbuQt+2+w9PQ0LpQ1W4H3gT4LqktDkcyLtCZjjZdUeRDbIB0mOfu
FjT3NPTk2Nxsgm2JsiOe90BvITq5y423VaN7UbVGlj82hKDZCfqRqXALemQrgfFDGFX9Y9SgCNbw
06CrH/wUInhpH9KAIINTW3+7xY0YZNsAFyXFbBSzEFGuSsW9jgpUsvmg92105QRy6dCFdwcg/pr0
7H6PI0hkMgPZqqlNF9SYvEwKuD3jWWVi2sGuGl5xIpS8XuEZs4J2ljCwxb/M9ZXHzHwaWTzyrJBs
wg6Yl8UsAEJVojKUMPG/SqXNz5eK/T17z57RhiOVyiUV1QSACNwXI3YLSGfCJlSjLSU0MK9Ea7Sy
nidlmu5iz1UNHUj8srPywmGhsX2YqqYDMOso7OwgJvW7BC686/vpZd1+2iUejqdeuLwEuf9hovbA
wSJZJoyXZUR6QAeGOCsU0Zc6/X4szUzzdA/HBDKyCvHn1K8/pkjQHh86iTExwDChifqZYh1OX9+7
g7x0boMYpLKMzc+S0cvxqNDlH0VrZpfi02na7/iP89IWK9Ruk3Xs0mc3jLDUS8ugiJoHc6F6ZjXV
1YvPCnsGjEeRE2xPhggqLwwpR8zVD0P6c7ygCSPexPXLSP0MDOeACrc8nwSLDsUtB2bOOLbyMKgy
7FF85+orITEY8FI0+XAIu6JEkxQEWLKsdARpj+DC5uxbnSMICkadYw4axjS8UFV4Xy0xLRdTwdmd
GQlHRM9BWY4itk5RS7g6OOTcRHXFkTukAhEVa6QMRzJcFcwOx4XYrmYjZsisqWOHYqybDVtM8dAV
9k6T3ahSMr5XcPLT9kOa5sTRWU2lQHCxGn6Xfh9IdP2tyN5WnnqKyzWt8SARG1QKWOkOHDAlZlkX
dLx+0vBj2aG+1BC4LISlZzLokMmJHS9NWdiXjxVS/kirPlppyjhfp5fu1X76A+oZTAzC/OB1mdlk
9txAk4lnuxpYHerl28dPJkLT1JIQ8A018lSNJNM7NUy9VukYa4vuiHHBPyzGwrjRlCorBUqKjQRi
kJJFifgElfxgFICHEHUT5Zr+x6hrlxCNAfZByFVcbeTu+Zs1JJ+pzDkhRjXSvNdxHRx9kY9wp9Tn
g81GGm/61SvNfrr3FG2M60WryEys5hasnxrSvhdIDJ5ByxKtwunnIfoyAZSsYhEwtxDIWQrD7kr9
hh7Qm2PpsyjsRcrJIFe6hydLk3vo2KJ4xFzdqiDGe6PmVyuO3d9fXMtRzB1qDyMszqoaV9yUyNj/
jQ7kXOhLTURQy1zXTd8s1zV+vE+lcn5FUD3h1FLkpCtKqXumRc1Tw4Xm0A3R6+N5Fg13Qnzbl68D
lFdTmLFl5AEGUhagOWAaAvnh8OLV/ziIzmeMsqtLTqefxw8yQde3QiU2n4U0neVG9aoDWnPBIWxU
ZJZ4xS01EdslpyieMODqtcAitOGPTXfOSlcC37rH3wGch6efWmSdKTCBwlM6ZdikqxwnS0oZR9zI
d1q0ftJNLnwGDPNonscCm1ULL2Do0Q8ShBj3vcNNSnnuvJz3T2bHiS+MoXjlJAw63ohmtAk2PPAg
cHNJ6whOD5wOB/VihHEtkWDp/LttThFjnRWXulMLyC+dm2iY9wJRJ+1IfmRfNenzGLyYL+CdmISr
jW3O8ir+oUSvIlnnk6vuk1CfjO3DM+rSyovTX4brUNLC92kET2iHZCvczuasKJMqS8/uRvSIaym5
t01WRGVcugalz8vWy7nmgQ78stf+UlftrTWLP78scLLFwylVujcp1ZmR9jwZqJcYE1fV20v6YYAk
8LNu9qLXUN6f3D9Tn8fan0ld9s9zaiTM1vhhfespy5EVCxmcn+x5Q5LdCeQBhII8yHDiz2ueOKTp
rL8flqefSoOObVFKZqyO/JEPNU11CN3hWux8q36csbTtIiZHnylbYNcsRNoJp2YCljs0wgAnseQ1
bdu6LbcwLp5D1SeGRqcxMzKFrrXmENzHrU0WYYuttDC/O2j8Sqn1rbmC4ZkVXnptT+sEV+d/mvzC
hKTOxA9gJCpwCyM3pJfmdNlNRPU1g1mW8QwVeW4M6FYzzdmFss9wITgWEKiVFjfVuGBDVeV8K7sA
f0C0Q20L45M4oWcbnV5Bvoe0+wDKNmegV7DW0ZkH4yDH6A461V+LJSCFoBvegbmA0B9oPtaL+G14
GHu81n+DaMVxFcDXKhRkj+b3sfenr5dz5sixh+Xi5nl9Hz2bJyJnrwzJ+FedYrvMvCQNEvezGfoj
OnhKLzy4W+/E8HFF8z8gpabeM0E92YHMSlAB8wcQY4/Sg14SUATTMQXod8+QBNLxZKWtEcD3noFP
6hrjnIPRIEUn0yWM90WGZxbpe89kGLiqIJcKpwviFg9J8QVAdJ1DXFZxAsI+DPrLR4T7p9iaGJIT
nIB/CzVQlQuc71TYZVB5lz+KNZCykKe8IaiQAohN8cxfUfF+GbAfVjnPsQ5Huqq9it6/saeS9Tu3
Oif7/IGoXAVFx4iy2Y5c32Q01d7scKjApIoibN6NQ645zQhqSImNM8D/NXURyJZdQvMyYpWPTbxS
nluwXa1ntOsgjSnMp1D1nEXDZ0KrVnNKEXiR0ke1Jpl95usrV6teK4DCmK4OSneBuAEoqV2XVNug
6cwYkAjy0iYhVNs/28IRBF5yikDAxDR7RAr+oviDOYu2QdMDxSAbCuqUDy4tPeVDWmFmrMYnyw5a
pMGlDHlp62wamidoeplA9r56xuZSxVJLLRy2l8guymzH0xmRUv5eDaQ5XvsWnBlMFVyqmx8WC0/c
HO6FBRNsvKr8IPfDbuxWzAUKGmnbZ3VDxRTgnF1o3jDz4UAABWkEOnsbcakXI6bxJDF5ZshxDhHB
B5DrsjFFqUWNLsj6pqQaoW8BwZMkab5fIgwmAEN8VCvu75c2uAb/7JL4mlEQheKSVJEF+2JrNwWq
TpaYBxu7Yk5ednFfs8gR78pqzcOjUBnbcIN3382OKHtQ5ysS0A6nSQifVFKYO6+ly3sbaU/JOknq
qNWk1VJPJyxqdK2zaoQSyMrVnExJ86ODXMrJiLhSDpkMUbA0KcGX+S9WtynKsHL9edrI04mF0HST
XCZm05RCyvgh19WiHZ9or5z1bCL7sLbTIM5aX8Ha7JaICxlHt4Vb/+UDCYQx1APG0Dc9cHa45q5J
EeDy2LTpYi1nk2xRP5/Z9Q9klQutoynpUHeDH8IbjClMAV5zSKeTRAzWAE2EKC6/78LtSJlNbCbK
vAWpH540LpouRbUr9wx54dFnulm+WoOiWZ5lF6t986GEUfS2CBPRlLXFbMO7EdASbM6tkth95NbF
2WH3pt2hrDYgmp/1TmDl8/Tu2mjnUHd6mAh/58fvk19oubWHtto3NXBdVkwUfw2vE87oi+Pdlheo
4pZQ5Vi/Hg9U1CdM+RAKn8Uwrq/25QrVpV5hmpAcij5iF0Wa8mYF+kPyeaFkYrywzebH1svDhYv0
l0TPNRFizKIhzD41THM3r4wRGiFPMcDK8iiliM9Dsxqz4rph/SY/OxF3riLbV94yZiB120RXzeIW
Ky0s+Cl2sjtHOSFwVXxaFOfYf/KhATgY37Ioztcy2TRbHsOWO+MJ4NAI0ocPuCz0f1mBRQLopT1y
DFCq3ijaJrFqjy4UrYC5P7FGKp0dqG6rLiWOg0vSA24XvvmH++BMMe6A+Lz2x2BAflJrn0cfv/Ba
+ZiS8eRIyPHnZU2uWhvVx0Wy8wKpwC+9voi3WABESgBr/AkWYFPTqvlxdav7AzmojLyq95UYEFfo
l1i/fI16SLbswSr1EVzpkAemAyGHKG0Hyw3Wwanjx3zbJyw6Fw6cJJj/Are9MYFs/tZSW7pGIh0W
gcjeTw3g6NB8J77wysL3f/cF+nakOPVI2usDXwaoW7Eq39lvRhIi4jdTaPTW6J9ytDuUXKXsFLK2
Nh7OjvfSCI3wKWRXSogTBELondE1cE6kOZFs94x9VqSn5Yjbj3kh5Q7b1MlkHZ/oGV16lhk2obut
lOwSrrcDDOey7JvH4t+BNNACoalPXyG5kRcjaqi0bLLRKfZQiLUzhZ0hy3Q703L6372sdnHKa7L0
/MQb5zTRxJmsaT8gys+IUMbhZd8akDf9wwZOXgM85DRnbMPbYwKTAL58ywJ63WrzcRKmewp2trXN
Yp/8oIycdHtVIFjIuC+dQXFoPD59BscP4oqvhzRm2byIGbDeyudZwSMlMZ3QP/1H2Ykmi3iTRz3X
2MrOym3qJyQQNQQKo38aWhEXM19L+gDrP19gJib4+0D9ktJUBtgIGLlyPCLHAjytWNyLehsTv/I+
NQHNmAl8zIfEwy5aivmv41+bculBg2gohmJqLRy//lV7yVQAmxZbA5WJIXNQYxTxKGTQTkMGcbzi
rDURpARVCyEJ6S8R5L1evwRLqEGDsCDQqseJVaeh+TD0g/eBc4Cd6cYrr9/f56EeqQlKV+AgeuSv
X/uxTMURq+qb3tTZRf6j7O+v2iGrbR4fy8dXg5JA4qMiKr5PLBw2OEXlRnWvy+tpG5O21FRHv0Sf
yZossVAgkFYFaHEorPuEaeRWHaXk41yRk8pNqkuXt67nmxIG3Y5AT/4N2zjYictx/m4QbM1Wc5i4
Tq6YFL4q4pXoYkIZW2YtqfvfayY5MruVmUTC7M5cxd9K/XEcbKU7oyglbgjuFlDfpHxzg92jcKU4
k6bfDmepcORU21o5RJRrZ/UiwDVuhlMh3eZohdJUcdaamHCh9q7PZcipDmPgO1I84fqntBOg0pzs
glduPQ+nU32C9l9e10H1XxWEPVhxYIIzYxW1oQkl+Bj0K8Z3MFQdF4nfNzH1EOdNGPuj0m591kZS
PCtjDz667KwpYK4Zjtr1R0l2xoAeovtCYBLKILS/FSo8Vv3nl5ftHSZN4agniMUvwuzxz7pk9XWk
Xb5Y+zIADD5JNSiSquMHmJhW2LNBwFTLg3hE93aDwPpsuzF3CkMaXkQWWQeyKK1A8cK0LP/H/9xw
u6tOCDGynp4nJiDgj/4B29No0XvJqFoeksEFxSUtOljVfMU6OvzdKAyG8yFn5vqv9KvWzRbM8mCB
An3MpykAw+PjFSYzGIRv0bGhA0bI+2uR+janAa+a8BqY9shXbqn2Du1KIM6ItoaJl2s2N3lEhD8E
0I6QDmulpMcONThA8iGX7SSUsHKzMxtPf2uu6tx1TA4PGlrTPcm1nHaowGSYE5USoTNIf5hp/D1Q
vWyAk3yLLldvbfcuHUOISS1OpU72jgZgdY0t+IE4FRs2Opyqytyw3jCBpRWpSFTO7k/k6r/jkGgZ
eUgGcyynMvBo8u4vW0Y/ANDkXQMeoAa/77kiHPQRIgZbVt3JQ8PFLk6vQ/u6V731Lx10xUpjSR3U
TYklwNy+tuywbsH4QuRkOglhJ6lJSu+Iw2mTtf0V502CWElDOhFMQQp8wNTs2xfwsopi3iJib9pj
78hSbkLpLD4H16YLLoMqNwvdMxFRJUn5swD4AOOsc6WuRt6hyVR1DWCH3lvl4SLJB3rWiQPVGaDr
EtN2RpYqlRgDWZcShT8LbKA4lok1NCFBKerUq2rgN3Js8hCDk3jhZrb4gXLgAsdaVxpWcFy0/OrZ
0OQgu49jd4yJ6U1Dbw+PVKXpYBtGTFLcKpITuNWShfXEmbzTkHSl68s/Vw0ZowKoGtF3WsLU/Qli
lpZIszeK+We1GNUniiwkE8vaklxez9j4jflXBqSD9aYf8wCPvD7DdcCU8U++Zi0Ug/UhHW7bwiuM
bF6A8Hpsw2UHcjO0MccCOjeqXB0HlU+E//A7t1br/EI4z7vyGm2rqIpLhMW2GaAf673Q10IUOfpP
kEEezRix8o7LyPmz5TIZTAc37IzLDpq5Q8MkKKLfrzB647Z/GnZptbX0XPVGJyNaBGqBU6dNtCa1
Wq5fn3ROY9zzfWHRnNRb7GJ7tKOrQczOZQ0qmK3Kv6iRC8uU4xZkqiruVb62H5Vp4OY9MmZipsm0
9LgfIGiCHpTIO0oDgXcBu/UpazI/lZo5hVcAYPFBoFkyH5N7z55kzL+CUhBusmqRuveLEuQxTf8f
4wy51VcGKt0WqITEBf+Ha7uTtEM8bImrH1t1D5if2Eu541+uXWUPZdhEPGhU68kMO95+8ZyBY9mE
fbD0FF73yKSPxC1gwY28Qt6KmWZIRod3GBXaK4HG98IPlGxUmcrmH3ztYOJxU3tnQQJnPLVrjAk8
6tHr1xU/QyqZkjFg7n1iyb22/F7vJzehSp4OGRGn01SkMFb0VaCtUb+3QMUpm806KMsyalZm/piD
Nxgi65UGGJ6AD/UN8Vs0x26pNis2zBKUePTcxJjcrfOHyuL305jGiXhvLR7im4VRFca0NULeeZpI
v8r8a0kbiwcsDf9sC1k8dFxyjoCjyJ+s+z6+lYmYQjmMvuBcQG5en5mwB26gx6MGQRZatC8MmmdR
3tMXz+M1ZCKoBxYdxoVW4STY8On/CnifQzkPH6iLCoH+2E7+RmMiZU7ThUPWl2GjsGOgaG+W16SP
AulcTyOUcVx6gEiveE0kyzEjwpZKr4HUwHYaTmcl6r30VceOFI9ySqpHCdaiLdu46sOS6l0wht0s
iEKbMBDwCaFLUw1HCIF7c4gp494couiQOjIhQRbyVmYnMkX1z7+uyr4kdKfBhn4DwYGGi3scobNL
qFQ6jI41QMSwCaYyZpnEZ9LQTaHvH6/JdC1KpJlzY49tq2N8g3ab7v8Eer+W6IC7zkEoQTCrzreh
EdHamsW1N3mDMGFr1AZofkFOnz6SPZt1/IDz353nfKvClAKVfqeVdkwVHUl8B8ivisVOCtPExwJg
ua6V0/8XlYHo8CZ1NDYJ308o2VN3jQC5A2Vn7BjA+Xo/VcD85WSwaa63Zy5kah3e9fVqXLhQSTfO
o1qtmy9FVB618IMXub1H/bs1HkVOYL0MB67fGVTpNjoPywqKsEs+QN/sf1qIiNXRXAMZ9Ki/Yvwi
MLJSAdKhxnm2wo2rNdDtvviFgoWebkBY8JyVz35PCscdLD6oSKj7Vl2swhfz7hobjZQyAvHTpWbs
rCPpmpp3WHx0u0X6WqLCNmgUnE5f3cyQvO7rKt18SOJli0AAMyIJa68szP7pW6MVEKVgoL//G4Lc
hc+YVA23zkJmq70HvDhJU/J9MiEaXRNXDGfOK3Lb2ImRzmtXHWpBTWag1JeZXpsDFPNhTUp5+X8J
HMz0wVGCtsrSCDo0nQGQaIq2xIo1UihqwsHlwUaWia6l1B+VguqlDDTgm23mtDRMniji+NggBcnz
OvGuvX3sA8LbOAnDg/m2PG9hec/CmCG/vEG1xgCwmxeSP+x4N+WdK/Q/mYb6ehT8fDPRYrr/auVn
OxsvLGrRndJGsa0OiZjx+2J1KL8GTtudg30Zl5l89ZQ+ECtdbwcolpkTzAbSY6+CYTXit8ctNu++
/+qmKfP8EH2ACUea0Nyjwg8VwL/YPT/tfzTI2wOPvHwE+QfxPwePyY00SRUTuO1pLqcyEl3Cz+Ui
aeEtD2RyLVURPgRHE8opfvOSoIN9o6rED/ztKQa1sEJL9S+TGeERh181QCRZ01tbzJ6/vn5YMWkL
wlG3iN2HOWM6Wka1OH6g6WkBYhUaq78J8GIkn79UQrLsVUnfUrSGgyde8Mx6BbMDWxmgk0SpfHBA
mzLmZ/vdMwC5ag1hDyYr6Ge3GF8GiyCd4zCwmUzyTtj4HWTbBzrVxaVdBhEs0mfVqKVnz3ziJJPz
T80hdaAE+FZKND6FKT3MeV9J3wY992kZu5Xnmq/AecEwYE6lem6mVSAx1W8bXemVqFCM+C+vsiv1
EZGD3n5o7B1VpRIKdiebEszTo3miVucxL3/7wE9wwpXXibsaRK2SUNSXtFPJkYTfj9X7Ym+7GT4b
0PBtsrwyIdOlKMwoVeJQobnPfC04EsXc4nH8K8WP7Ll3X+GUn6nR1CrVAR0l7WOmkzS3faoTLHaE
3WX8kAyjZRuxQr92GBlsrsgyXnnZFGn6TdI+fw3lV65jKPGSE6Y7a3gpbJVNtxPJqhsSWGCAWYEi
xyMgzQMsjd+oOvYEwGMboFLVqplETBECsMSRIg2BcI2sQqZ0dytW3Ul6CQLNOll2u+bKpG3kbAJI
dLTrAtDg+aWE3ZhebkqjfZva0lkf2DNEqsO/MduVZoMJzdZxESNcCreqFHd7AYCx12mDYthTLEA+
gooreEOg7btgZtJzQKS9EejLQvJirOmN3T/jmqQhsHdtw7Cp7uDunl7+/y2+oM2ePsnc1vOBaJnK
PCg1e7WD5tkCZ3zvIe4SzwmVCdmdP7HBntCKqh3i4aX+7d3phK+7OEVZ1NwhKntwWa9YV8Cqcqcb
S4oLlk7hMUYtPUan+H1YMmmCO55w40hT3xRdMMJzFUrmFEWBDl8EEzUfXmDkU7AvNsTx6ZqCgHkm
v21f3YYAdYbu8MHdaMEzFNiB9WaeI1Bapo/Y0ti/DTWV+CjI6RBOec3AzSefJIoOab0rI83E42E8
l89UZdltOvcweYiN7PJtugdRD1pHzFW4dPdmnHBu1ikIwZUnBdl2CwLZd6vvdy3IMhKY3FffJxAc
k5OWjPJLspfbM4XdVammyD/4g7HEPQU0EMv2AwIjJEXmQQwsaR3/Ub4VAAUqPhkGkcxHwLU32JFE
CxinLKXfdRZwlw8jZQuySHYkp22EpJRvV9azbWIGGeOzkGArjNAZXqSiCpx00X6Rc7IYheHA2ZcF
1FaW5yH0gt7ja0UuiLCLqd+RbHXnqJBEEJv8foIpjlcy0k1K+lObQNZJt1VXBGggO9WVQ/Vps637
tZK0FgPE6WSlLKi/Wfd3NfD7gEj0IPYsVNRpyTs8aXUgn1ovkh5OythWHyg5Yif7x4weA5JUGSGT
yhbuFE4jsf5Iemprou4avAV9qYL2ovYq73Wdso7nSuBO1EC2kl5ZbxJdZdWjlfijq41YBmWEFCUL
5Uc/YwIXjK5klXON81v/fz7ru8caIqRKzkSIfl19WaDxUlJoiAuu0yxn3ayLhtTFsg6/RQM8hCjo
ujL4+E6AIVfA+Tshb/XGkMfmmB+8cNPdyK4ttbBp+E6kG5RjCtjKhXWwHJVN6QX21WR07O8Nx2vd
WndIpalYP1NgXiRmE9Z9GGiwMZHFNlLarbmyC4Xy4LpvTBz/z+vUPRGZeashnGQ7CUnh1OGjECVQ
Udbm8BOeE7qXdTGE57UE+xzMtsZQXsuPDzwADAfBWHV4uoGOrir7pfN4xnH2YOcYOPHgqrVU7PYN
gOqoj5ZLEQrO/Y3gaftvbTekYkvYr5Q24yDD+ZynlcwFLTvTfAQRc0kJpyeKSmYAuJGzQLTJd2eV
VJYRJ9tlI7AgtI/aczQ4HDApdmOn6lCYMBjylAIPQRC1h2hlqx5MQ2AuXPYpjzK5W5jvxf5ip+GG
oLddeLzrNqwujylbE/tEWPYZBs16o0IjX91x0zvd3sfLJ+s78sOr2CgG4ysFLR/EQrQrGeQl1o2i
B0trwbzWzuSWHPXUgEeq3XtwFzj2116WtPkfOylFgdo6of86y6oJEHNaSGb6qX2gX3FeKV7775CH
LWFzo4BDmECZ7o3eSgU2h8G8EyxFvUld481+TU5phehxhdorJyJ1m7IUl8HhHbwuxiT912/qIcsr
QgWs58OTB0ouwyJs+7sBsA09YR6QcoBdEItUSJVp+N381l+NhKaRq18MS1HeORhTJE7L/wJtCP1P
u33iuwrJtPZHs+4RnM0okkM8QHopRbbAI3DlWzt2ZkxoFzpzyGrpjMAU6OhdIWrOkTlcqF50bo69
sg0CE6tMrisZaUaZ2d0N7Bz61ST0P9WcRHjV1Dto8WrCC8xXzOIJyqoyMKuxppJS0bBbjxcbOv8e
acbgaaJGR2VkVOsM7qHQG4d1Qf0CqTl5cbdIdzdD+k/NXNM6CqXZSe/CKqkxh6mNYLvcksG6lNjb
z+SQhuOFBKy/HCh5OvPW8UScqmLgxcmhLb3nespDN6o1T4PghoD4wf13Z9LEj3l+5RWAXeSipb39
T7EykKvOCW+TZfvPb6dAkAXFaToLZxCqtc7NOgI59g3Yp+XTZR4LdzLjIhwkjTzWIDjxXT49p7QK
TTJfeuKUqChcQSjnNWjzBKgpeIahWcHtpj9RuB9tuyokbn4vg6l5tunp6dKhkvXopMX4CGwMIKyG
Vu5mFodcYq2BBIlAxuM4oZ6Y9FPsa0PAbE1UZGqrXaT8fcjEavRgfm+zlOqtlH8TrBzyUdl9WSQy
GlQk2X8SBQRiPDv9PhHnBSkYziT/eAPNHarYOGsRi0JkREij7bl3Uj/eMjybGXjNMkMbM5dGQpNP
Qjp2Ixv82aT1iKOZTf6RIxs4zjgtjUObNeBKaGiNoa1BYCp9mPLAO6aRAy9qFIiiSrmMNG+oskiX
iLs2XEstNJpHZ5ggkTSiGQnjHayOOoscw0NE95MCoX5X/d3xOfVMasknxTPYhhz9XUvqaYS0+U5P
RpBxPFSJIP59F7w5MDI7kE6YVbdfI1ohZCav85vE57h6NZ2CjP09uD018gWvaE1UJaC9xGVx5mji
eiU3hjvmlmiWcinkaLHLmoDUHKJDvFZGUG9QyAEaCPQoTKKff+vFvebuY1+vUBhL0CUXrak1KD/7
LEjqa7nwGvYV5/wCLKe7qrlJJIZTKPrSCdGl/OBWY+BN4MdKtU3jq989+Gzi9N3PY7XoeasbGWu5
0yMfcRYhU95rgcH6ivvLzU+ZUeivgBJgFtATGH2F6y16c4dmYvFLiSKcuMj0oF9XHf9M4prdRSQX
SB30xaq7thKjzKb5b2X702i+uQoYoji790Fp8TC6Jc4MMXQ9u6nhQRAtUeUm7aWuOqsrBrjEhpsJ
3i12VZIeA+cU5LmxkZSwJI+s/74iSoaRnUBNcGP1Pao1qXGr4xgK9rCz8zH/TlU5BRrH70SNs8Gc
az1to5v9QavE2keWibSXgLjNDNwVRgFqk0c+w6drC7RfCTAwzxY6UFMOf/ObPV4C4HR1/iKMyYA5
rqbkIlKye7mXuCgYHL0QGMiIQXDl/22KPjs8NrpBnBmMmtZLBpyjbQwUN4OWNgLqltnhB46PJIq+
Z8spjEGt0+iE4tDBVhnTSxGGQK4V88WOTf89qhpbW5FV9l2sXqEUCZIQvfXpJnY45KE8+N7vGtxw
kQZatcIopVweO40fs2GM/noPdCAbSZA9ZzaPslDp+K0BAuJWCVaJskEcWzpzDe3INTmpw8uakyvz
TWD+LLU44Xc9++r45vSPe2mllAs1cZsHemQrxZ0AB3QlSjEk/vSz5GLfgs04S161x7FwONewBF8o
T24Z+tdT0N/LKQPMAIEQ3G3J9Xk+zH/gIIUTXRDsObbZvz/VbCfKXmt+0BerFvt+oZurYarM/u2E
WvZg4U34YOHAqNiWfE4ysHHBQtsV+SBzpfhXuLTdJ05UUU3/4oazBr5+bbgJmQidLosdIDuymmlL
eWXQIdpM12xGDhIGkTvrnHxrXkNGnuQ4foaHjGsJAQjyXuLJOnRhDeHowvkSmwP+XiSW9ts7B2LT
I5D9isPt+bXykaOS+/OD5uZkjVNI82NsDjkNygDTsIWIvBMnL1mpSGbPcVGBL87vQRojQ1y0ILFL
HQDrysfZWtn1J9WH2U3+1ng3duCLjUurksVJ8AulJUCvAxr8/kj5ADxEqHxu/IXLLBBpyUUszPUh
DTqDL4rqcLFTMlO01GTmU0yzBM9Yno/ME1DLnSi1anduOLCRzXJpFK90JD+x5hNY+ZXG9ZfmwSx1
OPLqFEjxGiEYIL+nJ9oCoMJDcQDnOe4Dj1TWGfy6YdnxeGgq5MDBqpJdgMfMfXK+scfyB0gPUrgi
3LHK4DnqcFwpfOYoJAb2sjSlbEC+dftXgMeBsnNO7EJKYZxTrlv3PeK9dWQSXG71cmBxykL3eFYh
W0C1TViu/rl4HnYLrCnRY4GiPjuwH6KEhmlbC1QKY+vLTHAxGkEi7vdsXUkY5W7JtAPEPNtd7eH9
gA0+iKDjEgPIRwNoRuLRblOx2qPvoJo0RjjAyQoRLqBRCFc2GOA2zi7j0pdA8Em1gYEwcGFQgKTd
CM0Ex3Ef+O9XyEE2vBD1FUsJnQW1YnMMAeOXq2UaDHq92WVg3EArBpRWkX0MYZX4vp3LBmIeXWLS
0Ojh1wIyQG+yJfOJAwYDsr5x8UXz826jQAE5VZdQ2p1InDM6Y2xmKRnBcigg8W+WZdoulcJF9qAO
82dsxfGWyXP2pBm+0vy+5QCjHObYmL/Bwyuoqj3udWFZnefz5EqVuLsTevCSnLKeL3mWRZcM0yql
C7fWqNYOkNVKyqO2bU8u4D3Vau+IWYKmeXsA09tk1o9p6bD1eYaS6eL5S5M1uMM3USxaKuSXKwfV
BS1haAIyVUpNo1JNnJwKUv38OXyaSzT/i0ro7uZAePz8D2gARXDAH6tRaxdEBdqAz92WsCiB/+LG
9Uc0twwCgL2tkJSbNn6+4r+TPkJwlQSfxXR/9oh1QUG8AuooIuDa4iqSNFSSG1Bi6ZbaH/KBDJsU
dnuloRDi/GOTS7szAblan/4VJeICqdQ8d7Xe/k0Zs9CMyNNvdyZet6LqcbgcukFLY38WHWsNfobC
jbMepJeUl5X4JeAG4trzkUdHlOEwYmANv8O4U1JqzyDv5znTB2IRaNKB5cgREBVGeXmiFVJJiSPV
1h3K4PCRRKvb6tDjqfgOZKy7YeUKUFVCkp65+qt0YASW2Ex7ITToOhTgO4cJqBTByUvyIRvcyINj
ejXfC+wxyedNj32IVt7JTF4KKzEHGThYiMubmmLg0NjpES5nU/FDmGL0ISArVBjAUTNeUE+9UaO7
oKklou3vCQ4Ko/ytOW2IvXlKUoB9k6c6RppbmZMDVk9amNU9eDhzH6jf8Oys10IOqr9q7xLjPilz
J7fBYIJyS0RhK9SFxZLCx1wkH+BpaJIKlrq5YNI5z2BuXz7dmcbsgOTDkf0sEyHH01U4w1qsskVs
NThE8zoIuGxSbJPzLU2rdIzCDCEEl4qn43lZ56itcCoodMDEFxzx8JjgzA0ILLTQrPZXejKHuYka
9iswqAtIGnA4Zs16PYPOXl/HYdR/M4j48EMGfc7hwNHmhfpqEtxtLtuiijOeTLmJAB/sgwglc5xT
U38Ek12dUIqQGU6x+FSThzNDh47R6M2Pou0nEy8UIW39oxS1xNZnem4fs/qs+CRyJ5LPEL1iBsSC
W6DNlVnk0Jpbf8gNycHzaTwkNl5q1Iz/WnHlO2rlE2GSjoUs74yf4DAp+riOX9oxKJfNQAqpojN3
vQA5OBPM66BHBCqkncHacyG6B9B6Kb2KoeS98hMmAHtaDYG68W6P56F05uHf0TT36UCD/UgR9REv
t1VEXOrIOLpOzT2lyav7vK8Ew5FsVZ3v+MwcsPPvzIMTBhB37aWwBAYZDJT6xnPF56r+JNW59oFG
33htPfElzxiLvXWBLzf8bSOj4V8DD4hfRN4XtGWvEKatt6LygVy/O0KNZRuOOsfgiWIhpTdJWo4r
SZ1Ycm3sUccHWmGyO409Ueaa9KHiZnExV80wkAvbYFeQ/X1PjdnB/gBiPAgd/8+V4d61WQr0Zx0/
p+1QaPrUpkAiimtD533HciEy/3zSIgmdt7jYmPs4LpQnUk6EbnguhqWa3KrqIfdOBQVTEzeLrqBh
LwJfI2vMXBYm+AbDbAENzSdoTwUZ7sK/NnBBXWgtkUNpM0CLda3gBxPSmuTkld+ePgF14YC0sM2H
6GlvTY6uMRiHcDZUTsMbP6ieWcRlwxlyr2VQV/SsncSBG5YUz+0uF50fTdT6+beHTHlRrCZKcgXX
Q+0ipyZRMhjTKkobkrOLuaGjrspbHEkjIjZfELVXuu2Rj/QDd5CkntKQ7r1Ghrfrr/56Ty1Z9SSK
JEG10kK1+KvNASwv2P/2w0p/2gXTvMT8gVHSktto2T56g0PCNonTJ/TJGt+SACkUGUAZToQEIg+R
mrr4cGYdLYXlYPalQOVu7jlWOygy5CxS1ANF+KHoYMyzQRo81UZ6PTeZVYETjsdLr+Gnu+6NYKhP
zpTdodkd1nIZNocvfjItcCECmXFOAzFLXjcr1Wx6B1JiTiH2bfaK15SAhE0jC+Z7x/3NOIK19pUg
pZo/GELTqFz/F97rmiZ9Qodzv2uhwYKVBbiOGWlSl0v7RjnVZWBkVnkPdGukOSoBsSnwb/VMkgwE
U7MU43FWQN+ORm2MQS/TkFDrEZdWe+2ozD823d3UEGuRcZS+4YUoh4nfC9PgK/2jk5t8X/i0+7RT
8fGkPYHvSUSNdh1UytPsc5Sc/Rx7PVoGPnSm2H3ICsx6YKe5c7qX4VPUn7U18DfIk1uWNQ6cPuHk
yJYP9YJf3FcAsGjm5aSEM1csEJA1szvljPn1Gj1Q4uW0/a02oOEKUbZgDCmII1DSQUmo8VNRHIsi
x9Ok69jvx48nFfOC8tM5pWRSMewaPaz/Bno+YT9Oq2WV41MW7Fl7ylNiNIbIQOPTZ8DVKFfMkiJ+
x8iP6986E221zXJYS+VxKiigsb/yYJ1ptNMm7aoZckeuMwES73Kv9+e8GCxVznClhi5cdBgUNxYX
YPVC/2kQChj51slXtcJVYkxEAm2DyUcygE/byyyJ44QW58AMeZMmRvFw4bBhK1Eh3Ju6k2MTo9ev
LbKa4ULl0eL+LAPov3PrblaKWtzzSnYET0AkeaiJarY7SXvV8McFMGCE+lm4nhbLkbvH/Z8ftnkJ
RZwsQPvaIs2RjT0CEXVp3v9wGRc5OVrYYCVgoSIw4G2svNU05GRaV3X9jBiBePAysTiHZgDaShu7
8+6muMQYVSJhw6+SAlvCxyrvLG657taESMTAYM4M4JxqZ0oA8nS9PaPexviaMiq1BRjbh9Sz9jJy
4C+VRhEMzwN4MB202QAjW1BpLBP9CKjZCvE1+6zE7FVu1hir+hWfQGiq1v5zo6IfsovR/o1nI5FL
A98rymnPmUPr8iHO2MfYUovwr9IqS4pbPyYzgMQdM+5Aj+27goqayAaIG/t31W/er83HYoHhZRjV
EjIBrw6DDu78kCMr6sHapVbWkz6hoeI8qJr65OPvif4rQGVm7SFKj6OsLpSgAW8ztslWTmOsB5XY
f7fTP+y9j6/fFWpB/vyNbvObdx4PH254qJ1xo3k87miNfVe2mk0k2Z1UdVNhHF/V0BFaNIhpLX4+
7ssO5JLjLEYvWle+v4ZkCJiUJ/M++Z7VJyEox66JxA9S3652wSsakNOk2ub0PNvOEJTGR9/VtuEj
PGmMc/VMGHi3IWbGQspF0P0m2os2wiOToG3eO/WSCYj6i79UrWccx0PK4o+Avt1OACaQHoFK6630
lETkay4pBnBx4breW7n/U30yoH8Mu5JrTWmyyOCI5nMMcOSErkyMmXyJo2yG8sDh56A6XfkIO7PE
UkDF8U9eMwdT/dFxd9oLRZqdqa4/+J1/ebixX4ZqmjYG+pRZLYQw4BwVCbtUFxyI/UPKS44grcqF
z1ad0XSVu7FWckicQWh/ePNwtc/Pb2+WGouWSa+Weh4e7YeSAZC+nV/BXl3vey0sSA00j0G37TvX
CFEmHU3YJY0OfrCQiRpcoqZhiyBVnBe29L9JhxmGAlpoUorf90r8DbCtVvhcAqQ6ZNTcHH8HIuIU
JElm1hRRyG6qN92ejsmDW1MSLB/d5cVqbO7TSRhjX2j5OYo4IKYlV4vRO5O2j+sxm5sN1dWWkDAZ
6P3ivRan3K39A/PtkSj83AB0Uf3RFJvke301LbTmlaGl7KeIjsG7Ti1Ln1T11ngKVZQaX7FKUVbb
yL/OdqIX5iFc1gcA2SFAR692doettL+WF3ehAK0wjvExExV+UR2aEVeQ8/u9BvM7axrw+4KEjYJ1
HmuMYdJEaWhb1kJsMAXTPye1qUao3mxV2mOIPtbwyTnWhIYSHsQR4wrd8zmkw4iUa3l6qHMg9Bkd
GEJl3S1f1JoggzRKEwHilJ9Pe8lFe+xfiLM5GAcPVMwylZzvXSDzxZuOv5zZukJIEV8W+U+7SXx6
eNGtDOVud2b2ReLzFuFtxqDOE8gcSarVYQpvCC9jyG02vnpFg2oJkOJN98DnwQ19Z+Q45wkUuqT4
6+fYsjTsAqlKFqkR2luO83r7Z0yxH+8heJ4QP480QTMSQDyh5oKIQktlPGoxtv+eyiWxgqeKb4Q1
j3pUchi1Ujgk71/XwgNbmN1b5ROvK5P1u+GM2DglgnV+XNTyfpaEbVCwieaPOc54fPD31yt79llX
hSH5fEHU8ShTJXlR4VgHyCtNoVqQ7SaPgSlxXJ/4dFRAeiZ+mYn3T7wYc/idSCoF3DwIptZ0U+eG
9g3WaNMtxtLmW+vrGJz/dUB998ld1n9JiVmwpdqU71L17ebt/bmm3H7JraZOuKoEiXcPwaxTQcjF
jkwmZh1uDVigOuHuVhgMVnJJ22Xiovm6cq7VYS7errB1wvG/Mq12Sf7MvKHNcdGfk41hjum29J3P
OYAVlaAe4uPvmz6ypWzIxQCa9fiX/7WJJiRaHqIuZBLCkESo4/7U/yQD1BUbEvLov6LifhUXmLX4
ckvb+Ypk9MiMXVODuONQBqMjusgPi3xBvFDEdQDlfWtMtaKAmzpC94W4tGIRbdy6jLCgWrN3QiY+
6yiMoPJoko6kEzKF7FQAdLH+aszznbOGIdxsH1XelmR0CewKXczt28cs/R56O1TsQ2FpwEyKo4RW
llUFlmbVg26qMvXfYg0PvbjnkUzPk1leGSYnH1pWxy0kHSH4S9PWRV4S9tURVef1CkkckebJ6/7T
PIQvoitOqQvu8FDJ5kkU8zfuTG7oNHzxDfx26AkzeUJaAp65quUdpsseWGyBhvUCELN6XxUeAKGD
hWDAUyWCgueC7qCPbQBAEgVW8e4e630kRS2HjjiDc+5Bqxj8n9ppqsVAZ6EuTsSSrOSGqh9KalG6
CAa3DAR00uVTCcT/FsQ4QohmWNUIAXX25J3Izvvyx43cw3VcpRd3CQwrY5tAgg1W5xkiKQGZvM20
1GXK7SVnRqkLsfXB+g8q4R0K2RXLtwj4ECnIfPsI5gN3R24alH9AVYkL17N8Gl7NHVAbvm++ltYR
UbgczebmSPtRD0aCzKp65FdkFjQylMmPhJvVqNmbhVMgNfV0hUjROhgmHQW35mM9Yz+ZIAugaaQV
peSPgmkFloj+7oYFktrl+4YUzn69c1GQYMx84YV35biz5cOTrQoN9Bf0QBF1dT5HdxJvigHPVFVw
OjItUUaoaTcYVq5xoaJaGxl2vX3IYKT1qmGi3z3Zw1vvvSk2D1iOBoOrSCb6KnFRd3sI/sAitSqu
FVdp3z9lSmdD9Jdhd3I2Tkt82fdjFMJxdQ1879LEYV2h0SlxlA5qoN4EyxfZsCZiJS+G0kX3NCRf
8t55AGCi1w8qN34ya0C5S9QopD+w0fspItkPk6iTO/SNxr7TNOwspTOp4GPbAia+KHIQhn4CS9i/
4bUIBRa1JYZ52keSZ7Uju0iOfhKBH+JWnHv098j0sjBHWb1MbGAQ2qMhBzl64QupYoxIAMSmbj13
JUsIyL54pxtxJoE/VVsrJZvNoaz3Cf5mArg3aXCSGH0kNjsWnC1Qd7uBF9L3EHp9Fmp9nFlFrd+U
RK2rQ4frM2KxX5fHn1hnbgdOmDjRuOKg7xo65PTqQ+Vje/IF9wwX9dD6FCaHZdKUL07Njg5uemaU
wPsukjcKt+iASTRGcfyQXq/KHUxAmmI2EUVWfUEWT1lg61ODs14MadLJDpV1gFf7tfgijpHYjiCu
VZoNZSo0xXmJY9aQj2axiAt+ROnIAuCNpFCwC5k5sbPTTXbBovlqDa4Lv5pDzjCmz0SE1HnD6fF9
nOI10zEqn6eLHajXaGYB8VDag0L4Y8PLqx/CeEYjsKUaQ9VNk5oTcSBZjHJo5+xPwSrCqXnLLhPS
R00J9/MfEXTHskRa5XsrwJRqysv4/ctTwxqyNJiGDvAKQceWOgF3VEdQ8VIC3fWeTv+rGW6qD70T
KuUfrwIIO6zOpejv1UtOJS1Md02S4JMjlKAk0JgilwfviGMkCEmSScI4BemMxmRnYsyRybP+yCIm
n7EQZYa4GlYmBqY/JYIFAtQMD7ZVQ8pt9yl6V0GzxlqmzMwGVfrzGZSqK4AZp46W+J3NWFWbT1S/
UHSx+PUV9A9oIfbfsfjnEn9JZRD/kWt/CAiAvlNmlr7cy+EwV17R3Ca8QZUTJLeFswnRuck7hIIc
nTIyK8NizxiG/C3SgNo1bVxZtJ31rbN1fIOiv+tb4/w2IgVBt8U6xuZyNdtEPyY9fYEm6nYvv0FP
3CRUvCUe5PA8V3kd3UedHn/dLHEOxA+BoyoSdmosq/Jrp3v5jH1S0KkTau0LOk5TIlXM5pU8S4UD
EWb7INSRa3SqLS9jwlVspCqy6/lzcluymAABCk1b5loEH+5iCjF+9SLujQiv13AEew8Sk/l4VnYn
UStDYWj0Pem1ai70tbFQ/xyXi3U7Gh69XCsqysIiyYMMscwm9Vc7YhQdLsjKmkTr/vibSq2oX2fy
2e9C1nAw0a+HwmQaxBmmy5a2qhXoaL/GdA0H4Xo7rsP9VpjPBCDtiZ2yKJEXvvIaxtWYU9/6xkzw
lO+45tGWnsS312VJ40eiUCOwFThBO6nzJqiGnj9ygGm+sugOh4kHLHrHS8t7EkhBHeLjHSA+whl1
I5SWRYQEfouHj+r6rvdm2U5CkeLHXbipfK2G5WBsaGEaTtYyAfFsqH30QwIBrmAVWg3QQ3L/F+6h
h/43oZZ8FJhN9mSX4d8sy63sQd0F6b1IFVNh7qIZkAfde7Oq2lx38/SffaVz61K3aAnG2pqabNL6
Nt74d+qSZqizCJ33T7F/P1TBkVvFlG5W8wSp0JbJ1WlaLKzdM74RFZNwMPMoqCAEqY3sT/a0Fuvm
JCfaC6YVaZ8LKqoXozTWf3elfJr54XqCB4bqlh2xAhg6c/X0ZhctJvv3qJQNpCjtQcFvvseS5RSV
3k5nPOEphcSdipyS8rVEmqdzeqcfRWWHGiC9WstvJCWqLNdDuHBHFU0uyVmDwOpQS524JXgt51XS
7bKbOaUYqJcO0i/bVMFQrpluHWaAc1BEY2jIgLo7g9ycCCgr4V8WzhWBNynw8V9sv0rh1zjCSC34
h+LPgxV8OSqjaoq8IkN5muvlBA4p59GyvUPmDpgYsOK+S9YMGR+ieZaxNUw84YO4sHK3Z9gpClvr
HOwqQHr7TAOREBO8D+efyvYY/KU0mxgwY5pxMcgJacibFFUU4W1KUbD/M+OEAplsaLin+B1aNeMY
IN9C/VyON81jNTrXKcSAlLcy5zMk5g6aQGo5lX/i1Xwn6K4yYo1muIsIno9QwE5vD/UDy/OFHhff
9xTObpNDzKHqvTRbCtCUDOFeHFm5RNs/ncaCBwJsOCk9Dmc+lHoQ3A+0/sRNIrKJMtuctz3ZNB9j
VXAwCU3dzezVaLbtLp/oS3oWaP+mtF4/ZJJbOA/BMpWKiJ1TJsEujkMpoF0CKFP+IF9x7btxXC9K
RTtHtG3Y0Kq7Z7yJfBy1GpjR2PoZTXQfUAnHUe2svAUxnfQT4jEQHU/imcJTTg6/moSn+/Ys5c0V
dFbvibeW5DJbiArImvQcoMmQCvnk1EDwoKTx7jcEsfGmnVnK+5wombk2Wu0BArMNukc+nBs/Pd4B
hqFVBC0tnwPL4RUT09Tb0OU+LceROKJ8wud/5mOlhW12pTVDC8UsNliTPuBftDXP0r+/r863R1kR
EJMl64UQSuORulUpFAp6ZS74wqJL4G98rBqbZaHffsDsw0CBqqSz8RkdHZypvnAVW8TMwLfiYDXB
5FrzXs6NE/cGCg+AMAfT95Rdbw1k/lZyuG6EWs+e2e3rdfU4k/PMW6TL2n2W6zIoxK/K/vPUGLPm
EMwUHbb8M1+7Y48/vnESKgkg0n7uXtXMbKW4DqDm+/FAvVnwNy5+Q6XHJwQmk4C88vM8iKHHR9ML
SqDLF/bcmwVayk2xYTAHyirvT6RtSP+BuNUVAOG8jpa2RoZ9IYvb2XjdT4bzmKffIddF18WY37mr
tQrG6fH8DjdNMFWlqc5fqjTNRme/m6rRfwPb8/QkPLsKDWdqzROpWl0ppDuGAvxs9eEYYjQH6cH2
ao6rqZZN7tkFlRpfb390UHvR35uyl4kSXftUg/CoUbyxmAn93kD7yjYWfa3E4tvrM3uoyqlF1ie+
Ouc+80Bn7wt3nr8fbZ+mshtUReovUx35UD74ES9z69Wi8Q+mO9bMWsznHYghBNnXoVbtegHIiiHf
2b+7r5vM7QhCgOgb0mTr7xOSczXwCB+fRj94SAvLwjymWBSCQguRPlZfKEBB1L5Jh9XIULnvtg4V
chzFCY6xYB12m7Rt2qefBpy/SmyoH7ODX5/8glsudqBcGBSf5gspKNglTFvjLtKLfna/q5zBoiHs
bVHsoAEeXRkGr38Xpk/EExBWC6AOzLDCfTLUM6d4qmWIIC2gZE6n00HAGgihbjctzC5+DXH1xhZ1
Rw4cs3nQhUxiOU4dmriHw6I4DeQy/3n2L2KlIWEpoJkBl1jG2SL34wrAedlqVlyzzDJCw0A8KnAi
df2EZytA7xMGC7SRIVafxgNeDoBFiEvTTB4rXspPvT4oBCqXYAf5UyJn2I+k47RuB5jhh388fAg7
6S1AO1QdDPjJn0eUOWRleLfk4hsRpiyONBuiDLbtEHv7Pu7vFhnqtP2Mx+SyDu23zPwDO6OA4sEd
sO/pfivDkp+sAd9dbOb6EW31vgUp0n00bj4OMtq+P4Xu/WymQjvWwY8VdX3DCd+w3S4IwjrZfjTR
8h1T4dw7sVR2UAOzKMX1ODMzIZwkB5YoFo8XDZj2vI0KWIZ/ixBiFyyWSoXQO8fIxuZ/+K3aLeZl
l3G8nfm5kRutoWk1s0+HzYdchc2W5AJtiqKoWZHL+5Za7xTRMjNpi+0u4RzpeKkOwi41e5hLqgpI
mNP+AWQXV4wx9FQ/ILZB3tVXAcTFzuQFT7/xFBogeo4P3RDrowYUlYudgHazwsDjT3eBvFEVulJy
0s6sphc7FJpECciM71oWlBvfOSCufROekElPJaQ1RhFyH6Kk/aWP5bDf6hcPll2q6xws9nxyP627
fruYZgVp4xYiIxHQfxV3wpWI7w4PuNrFvehiTh8szE9tCVGV9/MwMyFvi0vTh1Ne65ycBxyginAZ
ZUjIU9GfAci5UxeVz2cm69y58ef3SHXMT2X1yqMFzIvGHvA9Kwd6e7eCdUxSOjzvLOvpMwewRNoB
Ey+7m60SZ92fC+jEJA246wlbPwvYCQiw6+1zcWJdrZYeqcZ4unPJ9Q0y+lwNrt0tAnfwZ+THWQe9
BDvlb522obpFsdrRiIPFt+GqCTaijH7B6v947TyBt8ZByuDoKZ4enoWkv36Ag2Bp7jMgR9kC1532
etbVEqWUnsrjCmM7shkKAvLdkCxm2SJ1suxihnYm3T8zibQfnbrapBF32X9yaxjv3xfYhCg6E2bP
weGjkMn4Z9/FBkqoO4QAfK1RzICnjfais0FlbVuTQwwxJcL6vWsmo2FSdlMxQdRpbFTXM/YQWFEM
52wvOBK5QmGgimTUNSJioI6rK8r2rq9xi8M5RaeL5/n8nm18EVI3hFlMtAumLVBH6AVqoixasJNN
EgMcfMdPJlnsNZ3mDmvk5KJZ+9LIqfhuCx542AnQ+UnmmGrd/VQ0gssd+PzTSYmtEV0pFYx2Sx+K
warBs7bHpnEsAakMq33UL1Cz3fVWXBEn1WkbCEOXIAroxCdrdQLThxcjDF3Q0JYfeb5xeJYmESO/
xTenmVdpu1BG5TbV30+S0zVAKVshNrnyTW/NHBkNI9kvRnKWVD6XeyvpLmwpJTdltQbyhvURelV7
E96Zk0xUJbwsKlSWXlJBeKKJT2qv6HVYYhPQB3zDBtQnSRHU6p0jONvNV9ri1O0BRSFWHhPIDGVN
JaF75l7NUpkJlB546nuym/l8CuT5ejbai0y/3DzcsGq5evBCSyCZL7yFeh85APQhYOBHP1hrQfW3
9NosqJLDMkur/GOY803maP8hw0Gz30bqVKiMeULAeYDIL2Y+Gi4JifNDW4jMfPiAfKoaHU2pyMSr
2zkgLvjX623S6O362AZyEjs3fp8MQnPGffXv89fmC1rLEUataL1VNqo/9c+yUejJepFatBKaIHyu
I9j/p7rZ0Qx3RJDloGiwpmdFpDlGwaOVd5CFBFkufF/wuVuAvZ1FKATmkGytkrvkcIjVFXPCnUxS
BU1xa0EcaqVLcKRzBq78JDYBbbZZu8bamN0biHUhP9++ZdR41SjI5hCEfdulU4pDkw3kqhe+ZW4v
Lf6bSwKC/LBfvbdSMokojq0zvi/XaS+z4nC/P6Z+qgh5EHRA03/XYFk16XZOyO1SxJPoji7N8oHK
R/mzYaIDi1zkF/TimWhzBbJwRBOVGbz2KQzyHrWgF8pL3/B6trwz6aS0c6Jy6fCd0sZW6kLCG1/9
PvG81H1Jm/u41OA73BQrTZg1hmvVFeyVRY3hjTDv4zlaoJNCqhN8ldvRIt4flCEyKcRIFr0MMjc/
qdlFfGvAyWseYcArkOUSwTweDy/SuYDq6UisuJ63bs8QnjmznuegQR5EA596PGgPdqhpEBMyGGmf
fLD1XsW/gP7Htv4ePZNeipK6whYP/mvZm7iwgYhYRPLXJpJa45bLrdIxHgZUOd8cG8OriRgnVevI
u+ol6hckZrKgZShiY0r06zDErXdPOI6ciSZzwurkqMbhP4bN66qI8nkFFRVPb4mfG8QL8OeOE2Zs
rh5cKiRoeyWqB8FRBjS4maFkDGE+QOuEvAA3lq+xLh5qfo984sRAxJV9GvO/Z5A3iN5VYcoKGgPc
WRzH4veT+2JdeVYMJ+TmH+SvYg/0VjxcYtX/iQibqE1qwouqaWZ6V9HESTjcDfmDx5aC5eULfTtr
BOwFp0aTvaSWcUahkEDm9JExlhtg5qnL635wDkGs3J0tVUGxBFDRO2XvZwVTF8bdYyToAFWNlGph
GojNPTQoSB0kGKu/gvn7ZU52b2pzELUAqbXjJdjGJVURONQRd07rhxyJzhD3raICbz2qckyRG6GT
tKyQY9m2leuSVrkslGY6SxyCQRcSNY/MH+MF7s9U+24yy/dSNqhz3lIER4FTyXKLmsdcoKEEF4B6
htosMSDlQSSIEjn4HWhxI572vTVqAFWmmGaLeOD4M14UqfSnIJuxrWvN1ShyZuniS9bsE+cPor4K
VG1OPK1thORerS4F0rzs35QTCjkznCuonh3H4zDFOXUXq/8yPwvmsVP8wm6wiqGW8/Gwja7h38EJ
rgq4INcpwHMDaMxlvbyo6xkKPOqyiKSyMPv4W+saPB/4sCGv7GrOSF5QUUZt4uHLyeVZuG8WLkdK
ExlSoeGpoI1JR6XnBoC308RhQxLXmEGECBSBrsjfRfFaX/csZHze8lNmTdMJ6d3wFmhf66yxXp27
WUeUC0zA0Wz7hzrS5kFxhV5CDm7P7tIcaj4kMCOW9VTjphSQ1S38/zbRwC5AUebeFYQKTyGdIHTN
Sy+GgLTE/YWgzFKmFa+Zqbc17bQF92JCHJ4zGrVvwQKoN3uKAgYooGZ1/fVNIYuq5xE/vpH8Momw
7cmku0TPAU7BpevsiYY0nJ7gCclUkawPwqyOsMTXYwCWtvGTdmjaSuNE0Cql2BOGXpW5lbLFWuyv
JDFFBs5y5OI8gwvp6iPfiRXn63ANVFuObjygWpQJvfThLPyCw0onnt6bAAGFT76bUb36W1+thSq6
va7OcoMDmN3H0Y8xjU3yuo3IcAEu7rApjve6hG2BFA9yeaFMNv0MLQe8No2BLW0SuKccETP91WQs
n75oVYsJTh60IPR5HqYS2Wq7Ipnh67XPdudvAYuzGptu2U2WQhDX2zc1UEga6WfOlYQToEBAl9xI
uT56osomEQcNW1DFU+SDZUrBo7tx9/T/cf7474IdInE9F1cAxoPS2naucNCUmQ2EpwXySya+c8pe
juSegbLpZEMjPeJ/P6P/XvlvQN4MSVqjtdYKHXk2XIPK9NAEpIMLcJSEF4F/sNDAwIo9FRvl2dFi
F4SAKtr/U8/GYD5r7Ts7smvZ/3oS/VJqFW4oP2NPhExs6IhzmCNr+C9dNN4BWfuFxgS/RTtLrwa2
RADJv7NGMrmsQZWW6TYy3KXH5ZKAiYWXPxLT3JICipWFuADGv1F2KQOem6c1qfvRckg8+9erQOay
mzITyVVipiDQS8LwrtJQg1D9IoQ7F94MzBMipzIf53H7njFceLVHhBcXX8hTjjUJ35RW+2Ztmn7T
nRAPyHtCQ30lklj67HWDS8t2WUrqLILryZXsIod2Xjfl+Iz9eiqqiXqIK4axPP1Bojy5qtoTPIGc
LSu55oku84nCIxww/Lp/FHKL6By06AbqtiieXYedKl8bRCWjJ9rsuUE1p0F7in8iuAYv6vGUE5zT
GnQIy7mAP3NDVQq88qPI3bEoQGbpbpN0Kll2Heu3soKg8C4Ow37Syiz2izL4VpNd6J9aAqmRL5gN
me6fVHXCR2becTOQY37RHtQmGw+Lv95JzLTBTag/2zUJ6c60ZEgoX3qELoLFEfXTdgwgn+OJCiBs
p/xGfV++en9WP7sLYAZecA4LazPPAyP3XICNIg7cLEfc+xgbd8FQ4AJbmH25jEO2L9U0pElFRkom
r6m2CyzHniw0laaZRawLLdkipy8Nh6UzETjl6IEW48ImhcwG3SYCsH9bnKzOZA3V4jfaZGlmDsH/
xspZg/tY8U9hphMBeBK4y74Ut9dGJGg7Gylqg9GlJdnLE7az/szW7ubUm3YI4/mDqVHDn97A2bxw
njYGW+DuicZeywt7mfRG0nu9MJcgsaQjEI0RqrkWiBdwmnhulL0ZuPar2IfpuROtbL2Wf1uDUMFZ
5TnxX1TmwgQC1Uhx/UZN+pcR69oTDik+koVjcTUWAvFR6DOUNxtQQWMakix50iAAN+2EiLpAft2o
NKHeTXslOE1BMf52Pgj2Jl6LpE5XE0wFRBVHkOaG6z12zI3VQOiVfBj4DnpS4ZC/AlVAzZqO7v3G
wmMr8+nvktLidPTPj5ePucil8G8tIFoslasEwNelBbQAmiPkcguC67LcqUaXhx3Y8CdV4nf1O3rq
XvfFg6ZHxqbpxDqpHCuk7syVHhimkucyfHS941B6qdsPSj4rYRPVKR9ztZjrEB2JzEXuHFPPhuMo
fqQ2eq+IURyVxQDNBtdiYfKJiufkciKcC1S5txMLWm/4QQY1HTtJlCB2R3ytFzoPnhhMQApDsiw3
dvMzpiVeK1zo0n1wWoejn8d+2A0lW/XKqSrwqZ1kch3RGtJoZj7jPuY71cRGx3rF8trWazjm+WwO
TdwPmH4+7OwRUlPJL5ky6KJklppdB7PtAAewFJTIBY+1xnGrPB7AtwGbjobljnbxWqrqrkXmjbMV
tbTFvExZfA9g7ygOf4y2x4GB1mIPM0L+wbGXqTvTwqupw3BMBWcNVvyDOKLDSJCC+i1aqj1Aak/J
u7dYj01KRwhZp0pl5hUAJnbJodChwf9Sv7xAp8JuEIRzz7iEZ3X2OE9HZTylX3dGFxuwQb3nsixb
V/i+191PpTQFAw109lort9YGlqMYCIzZeIbuuER+NZFdBBKHIoz8JpILH1kSXtQiXW7hJoIruxOT
f+KcivhWBCk2ZsZRfgmEWB9k0SUybY3lL4hoMda4GvaMBhADY8O7zKBem3iyBGxBaHyFnFYwXKcC
Wgf8t725n9oJTFm67omtABdBWe+mKRJDNZHobFAMd9i1Qnqw12l+Yt+rTOxSgcF3zpsOWjnpDqU+
l7V6NVnb13NT804hWrAqDF12ceMw/1s9tvY5IRyNTetPjzxmc41fboA4lZG5vDq+6tRwUL1gAu1x
RM2ALOI12CzYzgj0OGRUSSa1hgIQGDs3eDA5W5K7ep/3xGEOQZPKgsiR7DW7amtZKvmakQzfvdds
6Z0zdTJnLvnE565RU4rz/rBR+O/h/O/vdjQr3s51Rt9c9QzFqJM9ABQJTWCM7ApcChj5o/GtXrR/
n+BKb2jL3UQX1iE06oV+XQr7Ik5S3xXpWwEcc7PYlkmWDv0NA72V5+MrRYZZM+tZL+j85wdw20aH
LO2nZHETc/GEeZV0MvGcpa2ATiZC3utMuJDl/YePXvZnnh8bOdSa/Per8/Gk06UcMuGj4LHU1Mt8
gMj3++N78Ove2Uv2ALzO2V4V5r+1sASWrR49X25VXvp65Eg7YWXbX/4GSu5RSzv1v4oBrDRt1CDE
ac/LS8yT65Og90lCYtETnpI70Oo61pBXugDhm+z+0+cHPFQIQh+y92jEnErtwHKDp8mqdqwiIuyn
dq9maMV8ix2uV35uY/gLEKDoqZezob/uW+WGBnhuuPT/JXjcUTvuUamWgyl9EbEzwYLqOIXiasHC
ApAdh8CukBKYNcF4pRwCDGQiKv/Bp17kHZB42NNiApCEtrtw8GvO9x0It4XSCZ+7gKzec9TUMMpz
gu4QXzyRz2OProYEECYEKfbBjQyFO5FpTJ4AbgEUSjFXX2XveFcBWg3xCO8zscyG+kEGH/cLn7Ss
OQb7YmsGkX52aY5PxzOkoJfNVp2SgorcfNk7HdSdmfqWvTuvgAvcJbfdpm2Rm2rfoa3u7ORaulIB
Xt+jTbdwLuURpFcnqCadllBBm4ljO8Qa48WK6VVVqDhc0UzDEi55XtgQwRlyC3+bHsIdwWasuong
2eJMr2w3QeOdchLcTWJcKGeEYT+7XovxkYkely+QzR1Qoro0PxOjTDzNxloVjdLu4e6iAaFlVbz1
K0kSLXL85LtKUs6OftDQdZxh5ItdkgCoYHVdj+2rU+mXP90ag0rbn2O1A2Feg9Zn+3cXiL1NgaMH
m/sKT+1uzBVyZ6zLVMa6Bxy6MSdBQcHwdKfU3pkliH1ws87Um/NRiOpU6RFmScm5QIEniZKW0PYQ
S+WyqSaXFRgMyo7knOaRcVY7Pnq+xe7ONO6Gt+c/CskNQweEGyT3w5AQxuyrSBgMcV7Yx5ZnAGhK
K2b2sqFqhAddIZueRArymRwZctVWPpuATdqP1FccmnnsZj+5QxOFDK3aI5SrvnRvw0Kb0AmZTSvh
C0x7MUDtM3GBkW+ElzgKWAdk5jk2bUKk9GulJ6Z/MhJXM0YEYbzRYC/MY98nLSkQUKRZn/OO986Q
UW5LXmQ16B0U2x6ghFJbctR6iENK7DZgA9PZmUg+TMclsfE2aYDdAUbv9oYda9IUi1urPuvT8/wO
jbDHlnA1USbKUxYOQBeWAJgDquFbR+m/nonUjGB9d+rqNErS/uxKixBx0AsFC/DMyISkTwqZTR7z
N4F0MKqLU2Zs9vweMZ7xW3dLEFgEHpsgcbnfyebqdr+0GE2k3idlycxxPaiG4t9RZEzyXSiZ/eII
B4RDSLVhLf+wusNDST0Z8/zfppDE+zx6Co1J3xtwKYmVyFzV4YIEFgNZlvxrPRn0afCsVbMJ4and
TCJce3iDdTe2Tey1jaCuxJLRqgCdPhXvM7fehMg7TJ6NGMmzeVvvFmON5xKlNvRL1u9B5/2zWck+
1dAYjKIzx2jMb6Zirbi8yUqnevcTh3SDIf8ZIGsQ5DyUnARKMuPRrNAjawUSzKFNjpqwBt4bhZqu
kUYvZgCoHCnKKY0/mkaQsd9nkHc9SM5AciSbH82Q1xEookvNI1C1YqjL1WWrf7izCAOzdaKuGJYb
fLx8wRhn2G619XsYqr6g5WYScV9OIl9L/JZeegJTPi3A2c6fwi90GVs3GMck/Pk+9fESz5zy+/Gp
7W2ctAKcTabZNuuIcZIcstA1PtwLVPoTmdQ2O/D3IRGKSYUvBBCeFX1oqFed/t22QaZG+5te4uRA
ykyVE3FYic4zm6oKSDW7lxLM9NAI87HkdwyXuS1THXMVmSciVjEI0XJVPWpubcC6jXKgpipTdPNu
r7jlXCrAtkhWkAqWgTmTgwZQN8veMGlZr165FV4nP3+2Wk1RpyVnQ89VvJT588wKXyJ3vLxdQJXK
Ipy6b9F8nZvpz/+xgGGZG56bJK2/0pGUtngnwrPlna8iOTaRD56t8xGr+k9VqCd6LP0jdi1FBUBu
ooSLqHusxvqRV0Lq6OZ5c1LULXcOjG6hXyx2NWLC7Q3+5TQAKOKCYZrfGbC0Q0jtLgzKrDrMKSl6
swkRI2BHj7L5FtghOTVEYE07NfROZuDb+0Z1vbKSR5FZbUHxVtU8retHPwyzvTECm4s6J2Arx+Yb
lqTrBIL4/RFbB+B41aw36jEKJTF9NrnNDAA3kQhD0aU3+WQyWkGVpp67c8M5AW41j/h63Oje8l+0
Dy6jE79bp1LpeE+W+BnpG256LPTD1puthslRzShidr59qpOoEbJDzeKQt15cITk/+S/IK4I7IGrM
azJGlXJrDYDWqwT237ogVn5aQx26OgtafJl33tsY0YLXd1AOqZrEy2lYU0XNNfOfoNoFRkYdelt8
5ZQDB8XcQEVCjYsG4SCbPsIkB8lWCT97kGQtOON2IR+FXajGHtpu94rSXOkOAfhH7hfstXuAcMj1
jGYM+C831J746m2XdOpFRlmQ6PcVGH8DPBdikZIDweBp2VWFnCWWLe9vo50DmNZBLC3hwZ4aTKn5
en/odSYCeCacZj1JvbKyqK+35eONLSx32oiz0DViHwjKyt6lizaz16dFkpKIUAWNxNxtR+5BKu9P
HiG11m4Ui57eISaUhXaqqRSsPJAH4AbYt2/rT6HUGi3p9WaiZwRu/jMKkA1QMoDma0jssWk2v0A6
DBkJVhQkoocUX2keejsisbJM6s+0zPVEBlF9blkfaWfXIhi8oP7SbDObTFEdmb9E+Fm0pIIn8Nsu
VVLAvfK1V1RhHwjXPWvKcVFCjZvawgYkdtuMfvIceBeevx2Nhr4j+zNdtl/DuPOzVZ/TwM9MePkp
9eo2zeXGmZmk8ssrRDhm+6W0AnddmYbsWG7L3E/Zs2paBrMyko1jjlAYhrO3WQlA0MrSdrHOaC3i
AofifOCcu3rTehwSB0+n0rzL9Tz8wEcmdcJQKk5F2mrODdjw4smvwt18Y8ZEFyo96qVhigTSCYvJ
Ig/CEMcN1GDmxVCO3UGA8eHlZ+izGzHmeXEiUhZXyN/JWmPETOokFqbFIU2kaD4hq1bQi0Wq+0Ta
WyZ+X4ai+XNpyvmY3KFG7BJTSuKXJO6tzD3bfxh9Y5wDR03usze7ZNy3PL8dWphpVpUqBadF4Xey
xBa+3P6VR9MiLsdtlLLGbrv8kTz3ceBuoAypFDs7hEsC2HgIej8Ye+EghkHd/6TS+IHY1WIANgDB
sZuhCYHeoyYTXMemmjgcSq006MGw7BPgOS7Hx+1jep5k7sfUjEl+g8kHoAW7GA8lTpEAAbGJjDaJ
L97tFwTIv8kT6IZShfhV94DiykRwbqDzJu2LVmwGdX0q/BwcbC22GVV24Wfq+dQEA1j3Ew1NPPm7
xx0HT+Mjw3hlqe1HXRxdgBBB0zBMyWVkFm60Ppo3EyFYqciy1qkr4iuDqVtatfz8D9kUP+khjfA7
GVTlwMGVmwlacJR+VOQLemdBGu2PxnbvRMaRUza02+AEnAEGRlYI1jqA6FIbYb1gLn0HBsSQfGWc
MFXE/EV56JmynhX4By3p9/05qNrSezZ1hI9dm6vBtFin0ViKiehf4pN6woxpcf2WdIBR005QxGLB
zP2W7K0eY2+RKShkf9xr37Xjy8RXA639cvmpTVkt2NO/0T8G60XNG3y9+r00c4xpbekMkh87RiDf
7b/T1VgStcwBYy5l58Cns4rgXu3P2foCKIFavApox5CyjPruXIseS+lHgdMa0dqrQIkdqICok+MV
Mr1OkkNDHJ7GmOy9lUZ1DXIiCz3YgTU4vp/cyVjaJgutk/AkMCDFTFUE4BDM2d4C5essLrXWhe8o
jUj2640MJmZ+AabwEFOd/6CEUWh0p9KksK5SvveLUfkp9VeiLZnYkjmILVNcXBx+0P3F82muMNwi
iV7wfooJrp1WfrmzFtQDvahc0GP1gFCKOZuBnfktAzngf1o1NmVrwmuFs9nOFr3p1Mo3dFzJLPbn
Al+YUIiOGVUiGT41AG8iB7Wd/FPXdbC687zDVNl3HiykAkrs8GwpS9uZhGg9r4adhEcGkpeqGFfa
2bMsUijzEEQ8GCEGWUJHwKqov+/D+eIbti+sCwfpKYD+8yD/Nt99NirsyUEV0RgJLs19vqTo1WLH
bwwFd6ABHFvKxKbLe4VKhIt2I1idHQx+LLWF6ECUc8hEtoogl9Ukxo+FwpC7QXv17UhWyqAQ2K8G
c4BtE7ButRIqbG+LYlKFP0G5o+UrMFa2wSPahDZ9WYZbZeNZ+afP8xJzLE11yHUiyc+v9h4IjPmg
nTZhAzxYx+f5cTkpz4HCyvYi4pjddilYksa3uGKIg+p4wiU+mkrwcL0t0Y/uVrAcb3x/9FyurKzO
0H4R9+TtK03HQssMT4l6Zc5p9ZWhy5v44WUitki0zEgKuvvla1ZmRgKtALqxzCnkJrQJfyT5D7gJ
Ux3RAxp6sUnlkHl5c4Z69QWqhc53SnTcyAIOlh3Cqq0KiJy5+8xK+vj1PkWEdh3w4IQ7g9ZwMiQ1
rbzGuS2UnNJNRKXmeXO8HGxmQdShLkN1NB0oJMhj02o2cnYp0t7NwdJ/sVDBB/jOogO66N5bR+Ag
hMKpVY0r1RuIXodh0g+tLoGSIe4uvJpxCvH/JIKphKjz8wsAR/hs6dFUQDDavPgqdW+DHMnHEu2O
seQkT/9hYIV/1Hn/WK88LtoMitFzUW7+K94t3inAdIfJmFlOHIs0Q8hVVfsObjHwn8OGJ7ILfAvY
jPmaoX+3qot6He3OC+Qra7wDkiwtRyGpAuFRTWTmX6csSlQm4d8rWBMQhJWIpRNd2wAl331hZfX6
wGBNyxczMTlggU+6okLw/iDYbjqOG7KQ6jyaaOtubD6ejiQnRJIE5+neYls6jkAlBVQOGWrs8ZaB
0H8goDKY171A8ofGo8mvYqcICWOGJvrdwEjrZQxHicuQb/xH1EHzC9pHw3ggq8+JV/WFq9v0CaZQ
KljGGJbLurr0r5iBaUrAgHUYvlnmNWzcAEf2QUJKzKs/95fnRsELSqPAr2ID4nnH96gKhccny5uJ
VTPACxkxrcjZvX49kXMdGH1hOOkIZVpKiFSta9JaEEfXGDfekpeNAH0Vp2+Vst2GIIn8fzk1Pz8U
PUqMD/NPYjyG0PSRuwOtfaXXL6m+bgNL7u4Z0B+lhhGaCz1LEl1LtiEkwKO4m0eLM7r1emVdcxdW
NSl6ZDIAYPh+xMSXQ6ogLRpOMrn9uXCVxiE047DBS3yzQ19lwwAmvIX1fl+2MzXhm/JW0KSwD+Bf
z/o6gHgAKar+kPiX1bgT6Rxeg8qon3OzcSD1S+9XDkxTMTaydV+PhuwnyRrhnXexBOqjaGuco7yO
hjKdraVIhueVeia/2U5jGJ3mo8DigU2UNqwQHKZVlgpTXz4+K32ERVl6YesYMwBjUrpzJeHbTwwN
tE2WYVxAMwgQQL4MLzPZOpsz2rzEfIkDTnfgwJqYgLbXimh0sizzD6KIzVOAYV7GUoZRV4CJRKX6
86FLNYZNfO7+Hov7DFEG6MN6K8jL/UsG/tMrL0vEcNhaKtjamt9UfYwh3Jm3gfMy5zGua26lSvUj
Lxpsiu9OAyOTS00NcT2eBbz5Xjq7sB7+4i+4IfSsUJiTavQTjjIdudNTaHMtB+w2AcLFvHANpr5i
kS9ahSxf5MEXS5dho4T+bnBHpflIIr4Z/rka4gGNBD2FmGX8/5GReWldFEG8IGSdhGK4X50un1o1
G78zaJd1DlJ4uO0FnmoNJ0nlZQzLd1y889uPh8K9VsGIPl7TM7g+p1dtaifDinTVlHj2gz972ta6
bAk+hj6B2LdGhAFvxkhC5ZR6Uy7h39wzbXH1QP5uXhLrcp2nniS9sqe7mxsnu9rMhDo1C2vebDjy
d5cQ7xNd+8rsOsgEpMMF6Jxve1B9F5+/XfEYkRGgqPozLssYBdNaXrh8ueUqgnsfgwgg3NQNYthF
XeufWBgX4FjbOj8fFm5+HnwbLEjMHn/9n2ktrc2/KHtMIgIBOT01mexakOmGpg0WwFR5WwW2SDcb
AycnbNnQN+TfY2ESpWbEfgy7pL4AIRpBmboBvSMgp5vzMTa/v4OnXvvg1sj0j73RSR3SB3eb4exR
QC8u884Xv7MaJMZwGkQ45yhbDMB4Ky4fCnbrjk1zo5fb2sPuhuocmQ0QpxxBz4klztozGfPMvUuj
V1ot1cbUvBUI8m4yuhaxQyWecVyCy5P4+HtbxSV96TsB3GO+hwSba4mMpXdMXQsYqPMvP061Zmtv
Uv1tbod8hH0tEgoiG7yzlsEcwlkYKIBjnepmHKYNXnwYMm2twYfQU7n0eYZGERD5M0jLQT5iH+J8
a3IRhJ5fttjx+42T78g+9zKQYkehTfO4A8Gex0HmWmozLH2/p6owQWR/elZPEr0yvIV69rHjHQZC
2/34rG8Wtvv2sdkNgS4pKBDAlgSb8Udtes46gpGScK1X/NhDrLMk5H/n3QbhtKL15x0LlhNmkzzp
Nxuy/nJHlgqOGntsQ6xQ3BBoZVu0DKwtJpm3/rypVzBej9tlq7T0jQ2dFy3tdKrMELB2mNxJyGHU
JqJiEtM+9abAAiTR+DRWorJA+Q3OzjNIEm4qTHXP6yfVCEuwMkJn2abjIskya9DXeXaL/XfPQAN8
MZgxaWZloODpd7BjopqTz7UfvqXeDZ49pyW/5hhZhg7vya/Avfdub2pLfSCWvKXO9iPAAyd+Uzpy
4rgJ2sDNjHXhGljw30gHdGJsrRcqVIkaf266f4/6+aJlhS0U50LsuTBGDTmqBVk+aov/iKLACTKI
XOabrz15KnW64DQQQ4KAwdwhoo1y7VGIbsWvkFurpQ+DgLa8YhDH8kmkljj/SWfO5NPCFWy86nSH
2kFVKKpse0yu2sHxuc7P9sr4OHdfNWxJGQJZpAytwV0rrmhpuIpJTCJbk0xfQnga782BR4yMss+q
Rp5aqajDc5FCEQcSoqz+jrHHOeMKkkwbQqTr2gHGjxv9VqC8YEjHdjifvvUuKRJGENP9bRs3tPJh
iNPhmV9d3QrWw3ub3Y3to4lP9zG37/JICjgdA6/5Qu4U43Iy1akzwTzgYUPS+QIwrX5PbPDajcSZ
cpqwocxGjEZprV7MDI5/k87mRTW/crFAZv44QqgpkHRXBao53qH8xCvhwCZqcoy+pZPeAaB217al
d3c2MF9R0ttkU46jLiQ8o9KDfCCuQPh1abYUmzxg1s+eKNMLpvYqX8i4qD7uCeBvNOEdMIsvlT0C
LcaN+wJHmqQcuJbGJauFsqzwqTBPhH0RJA4rn4XdkWiIJbMh2gZL/Uw0FnQjrEhjqHW2I8Rs8yi4
WDAhDVphuEkXWzLTclg24ktG2KLhWFlD01sLJ7DXS0IjwPgj98Vd9GKLklYD5PqF2xZr7VW/UeuA
1M0Zyy60oBqGfdAF0ma0SLLveRX5U8DfTAs/+f7uVHeUJ7B0l2P9tXUrQ9c6UB52sMtb0ZNf7qmT
zAAbfWoIUY3qFbTrdD6tkM3+/RMc/09CLj9+55PgqYCHQ1Wp3EE6CKgxeSr1yavwK4UcbptdqlQh
CG1NxBe4SrT/dgWamLYfgYZH2TaDMLKNeD3prI6zcBQS2ZIlsJe1n5VEFUJpgT6eDZFLi7Ad/TRv
pZDygjKUXuIPheeexAhCreteBrKdEiuWynbhxSdr86lCLFpYNCc2PvCZf8XrvVzl/M7o3CadaXv3
zahHgKk1QAnXoyFeFsk0q67RxZZEpSm8lgfG6ivlN+4K5a9I6QihInXcMrQGPMuIS1Qnpgv54dLp
s0haamndRHEXhmQBcdprLsGt/A4lekXtXoJv2uSRo/aiZie3xCv3uDej40Debj5eKEviYLzPjcmX
iGS0juNmHXmJW1PGaFysKTEMyoSHUXSFE2zY8mP5SFt4TIsGMJrA0W2UpQyr9f9+diO4G5cn+/8m
JzMKQaY9ZB//40h8K3RcO7oSwwIQaY0h36QiMBL7NyjLqddIfk6DhyLuxWMSicqw+jcW14G0stKb
btphVwRMwuDUDr6MHoq8gMy1q/V2g9sANMtHkRQNG2Q9cKXGoJco0O7URslqnBhTUSZ+DnSZ/3oe
rhHfEReU2M2HOaj7F9Rw61wExdGcaHKJxf3m7Rux2pk+5wJwUT5l6tZvlhlT1xJ6o0kDvuik3QE2
hBqTFCy9esGwviuQP3ZvCwPPub34hSq0dFRF47WI++tkwzUjT/S1FKIjHfiXNyTRJAMniPTN3BlP
/nIQ04LTpvMa3m8pEv0KJ1W19kjSwHxY8ot3u72KCc0Yq199BHuND9TGR8rVI0mWFVvbfT9v58iZ
5NaFIhuY9z+6KPHmV7yQbPyX6V6vViivXqQqoaxnS+NOXsrBqKf+K+jEMIpa5gV1f/+H5XL9Igxu
iz5kp6YIT6U6oICB3e8ZMCDZ7qAHrfMaApoL7r6EIOt5lLFI5XN6B8XfeoHnnuem331rzhSrQQWK
jB6jg9BPWSPIEcQE0tV4ZzgR9YAZZWGoUNui4hQLIJYJ6A0RyTXHctyUUmrbDEq7jpsvw2Fa8I58
lx2p4UEqmZRhJ6ZV2wMwzVk9k1G7yBGZvHX7NQeKGP6T+0ZJdEFXlIkJUhepZfooxa5Iftq2TNVU
/oI60Ajiux2fcm+bz3bqr5FgscQywVPYVbbg3ZsEWu+AVhhTzhe+T863ZPRWXHVAgx0sZAaTi3O9
ec+EOqdHGRZmOJtPUl9IsaLqQaK94ASci7+W3JVxlT35S3XyePJl9Nm+fXhQtSFJBwA4EsmRZjtP
b4uUtYxkwDlIjc7oD0RPeoUZqyexhm7QiIGJrPtXsqWTU2bbdCFVUu7RjMzI10eWVhfwR/jksqMY
JGsNobTKNjzPJkHHcd4iI4HZ6b6BNE55gSZraK4vJ+LVZl7shYQ4YpO5ASeRuekK3sQyt+SRm/MQ
i0Z+eWT0ukSvXyoiySPxfYBOF6fksKvXAcSvJA+oMT+HOxdqYKt3pqrjZ78wl8c7ywg2ohsES6RK
pCmMyEmh3bmg89dNS3UGsGrcvGAycJUfux6Jky5kgbXfWE/I3beyx8JcpbL6UGycFk1s/ZPrB70+
2mkwnYEDyOcJ2SRBmnJPCXYrJGIcOJkRgjwP/deJlR824w8qPcq3SGgqSvYtUcGeko/rqEtA6edP
1NM2anL6E08VkTL94OoQN3cGUpaq637JT0XRTw4WsFHSiZjF4+87TxxFrnVdTAs00JyaY7N+26hk
ty62diGqrM97m7W8D0sTk6KgUMx/jdG74GD/8iQPXyBrorDwrpZ87sVMkW0LbKncNK9WyQ/NhUEW
LuJmvpF1llO1gb9qbA7QafnsmXyQi+ZeeBEioajJJSmBYbnYO/qbeokw9/xyLeQmd/xoY1KDhZ3K
a3g4oQCwOo9jSbRO8MkIUxAkd3puxgpp21IBXGfkVLWTocvPIk48fCz0c5mpVngvpvs5btm0kbZg
l1oTu+Vyj0aJXzbGOaK/kOEtYNCE6nNvMS0cKPEOq8dW+c87p7kgyZQqthoTIadCiGQV7OJNYIwT
lpFXSMZa3hR06bRZjwzG1aJzfEs14hiHJ/2Ctop5MpMiwaBx48stUINwLDR/qQl6I/1FEcFNlblb
n4wvo7pEQFdrNsALLFhhnCjk4I4sWWpW0tFtmQD/lnolvXjyAnX7EN+rn23yTle5/xpkNWvuLky4
diiMWKfr0f8nzv/mmHDNc7uQUX3g5RZib1hR9wT12ivm7tHSN4KpJU3UpIBrrhmQ1ft4qKCg7grx
1G5D6gcErr3h2VpY6CUAhS/ziiRYqRsBslL+fVY/U6NB4OpEn+vHOVxLnwgK/5m2Zy37LwWwipFW
FU+c42AtsjrpWHGmnqvIbyHMz5jgfaeBKDR23fYvkTJIbDdC4DEhkLpbXE3vTLpH+3FhS+mnqHoD
3dWA/MtH0dfBHE3SU+c6oBGC0710MEAWutlkBMVAJwaQ+dc9mJDiqN/z1/gOovXkWdKGYtgURZPa
06ieW5ZAXwrhUdP1Drk7ZEOyc2cKD58r8Q+t5EGR+xflPK1asemv0kElFng2uPdSVfPY5IqvpUod
EydIvHBhaaqBOERi8KX4L+g5Gom/BgQg6lkJfefLMk4xCGdPwwguxkgcXcm2EIOjB4+LKTNvENNB
ZTgj6SBL+wolKjl59bsmNHHw7KfmDrjOriqLEg6/oEuHaVJL8D2R4IP20jG5GBR4ron/j5MtmgJR
PS++MP8GzFGB/D7JKZbMGeMy5sdPu9LzPOMqrY2coUVOPR6VldvEkuNkKtY5PPbFfNctFG0+CEo4
vCO0RMFe4I7nZsRoSjEdDFf75LgdeJdV9/WKg1idGvjHi2CoRlBBfkNdz3aSUPOkT2UpmDDwOMtg
ht9x+5G+Qv+0LpFM5RkeINkjxcBEiSjFYr2ET+yChz309eJDK9BL/VYojUYeBdK36mlEkZWBWOhT
iaNFnSNCIsli8bNpuImrASHEyW/SjU204iGVMA7nGT/KWeBAro1tiaUJYi7iVwIkuvfFlRBrnjgI
7PvOuqEJ/y8Rd4z1GU6BPk48bJSANuNrtzSA75XnnnZa8CXu3K79hcCceuD4MLuSC/7oJmgRyj1V
1+sP3rJXf+D9VXXRfsC7Yggq43rUK5kqgh5iCEV8DlGephWqfvfw1CKhwiPZUl+9WbfWPZAAB06r
Z9dTbxef6gb/zUKXQ81/hYaroq5V6J7OiMeayZ0mumWpwOI7+klQlhkspfXlBh4owoZRLvRQEOWV
F43SeDIqx8kKUeewiehgsF+K+A8EEyhHKgt/bFyZ9in1Ram+Tuc8ThV9c1qmutOA3E7J3Jfn2Wt6
se3u10tr4DGTVXGChlDcuyc7S5J1CvV9tUJ64FTDUNvH+uvijM3n8BCJyf+0MekqWAqzFj/TLR7a
W0EVyZEqCINQaaqSmZj5fCHhnkFhzFVMd1lgI7bQ2Drb1+4ZI7g7RdGQeaRwRhbl6abr6htOaziu
gIHRWoH7NHkklzEIwBzLO37YryQ0FghKD0AZzImnNflpurUW/YPPqsRjqvE+/odI1NH/KHzKIbOo
DalegLPugJgPygPlH3m+RgzREAOkPh9/MUQGn3CvQyJsJF+O5gdrtf01Ut9FqEgxp0Sp6chIxb/l
cZWOTzCfcfV6e4Jf4/WCqxRS/WFiygpc1AwVVjN0XgN7FUdd5BasgrbylTbg5M+NkIRM9OxWxxkc
aQXFkc6M6bbeomZkFQlZ9W7bgjNJxwhqSnukdA9c0BK8R/7Ylu5wQIIBCFM2Z55VjQ/nwddEmUoW
ok0ynyUtUT9cD2XKCj5akp6W7V08h/js5olfXoWTrVgKEtEg/FXpxK7xcMij/+/3z9oqT+MfShDY
2+rghk4i4YUnT4dJyEX3qn/gxjsHnfp3DgsQmyFry6fShZ/+OPmgRH11bL01cg1UMwpMOWwqeJQD
X8wzOcvT+kDHuq68gG3AV4KTXbRvzyb8ooNJbmISsL6mr8LmGPSm4K2OU20KV6d8KZ5QJ2kgkdWz
rybQvSaHd0HBs9wAQRWgMvER8ktyQyegA2VswGk7dcAu//E59FdDuJmGdv4g2QfQGytf9swILlBH
TNfl0O0cQoZGmwUKI9FDBjL2UOSFhNx3jXqIsiwKDpAVXeGWDTzcbqJyp3JHKNmECG84PEikTaL7
AF/zGr7wvcKU2WZ2WPnC5gHG+jiF0vGhe87tV6OKKC2xeddaJaqAgAccD679fXQHqMZkfegzw8zS
vGcNHwm74D+D5YNeMujRFcgK2aGcC9LSkXzy3jSy3nkhsJedZ5n0DNUshKTZCrJwfXb5DjM0GaBv
3kA5b38wIW8rZ+lCCB6noDzECtXedSgxJWk09/Q9dMfLSJ3FNW2trtlaiwjoIYN758Bk4EbPEYqo
3C5IafERRD4V4MYxkPQS0NbDXeVI8HdQXbEg70YyaFxdmPiYLZCSXQ5Pu+45ukI/ck2c1+sZhPd5
XvUmh5NcmeWCY8/FdIfm3ae7vMNroFsAiCpu4rBCMbTc5urHLm66brll4QhkoV1C7ga8CzHAV1/y
kJrkALa6pzpd3ipv3CM6I4EiZA8T1ZkbHRCV5VdX/xiIkaHkPcYRaGqq8ef+zhBTdsRRswz69B7f
WeAefCPBoiqsdieET6TrYx6CD08HyfVB8hWlpb9TwAx8D/tzkP2qaQDv45/va41vJagSt0LhjF5B
4bxvczHyZmcd857gkPx8bRGs9EUyVpNhE+KLf6ZcgTefMyQAwjchoEM0x0IpH9NfyAGAZBuQgADt
jeYVPAAlpndy5X2NyMNTR36bNWvuDyzVPLv4Tk6GEYYDfA2ihDGNLhUo9FRGeF4EM6olvitCj+iy
Okcso28TIsbbPSIx2T4o/Ox6FnF3thH3XsJaIqrexee4eJ/qMoKwdtsp4lpxV8Yz2/k4Rv55xRTE
Te1R63/BINMJA2hYIJzMECQUbRm1TTj66Wofe446IjP4aldykXDy6XZEbgYibeeF2iaev/vNLSiS
P+oN/IFhXdkLmKxLe3VR7esiTAEAQW0B9fLfMj3VsT1HfQr2wFPPnNLuZTxhsZCUFDAtURXxjn/o
f6VzonDnMzATwrWTypvhF4Hbf34OMIIKdD1owDO5BRgmqf11GHTCh7BNXUX4o8V4Q2PybnOstXFW
CofBr1lL5ZDcBM6qL2LtP1Aeh9JH6TaU7Ye1NGOn0KZ6wmYlcQ84dQ0e/o0+OcgdiuChT5AQEFcJ
2YKykExjFJJyx0jduOND9dP5lL45wrNGdUmD0dAXbDg7qVOKtraHI5R7CxLOAAVcnvrzn4boHzbS
/Xq4RLrOCmDsXMojFUJP6HOn+/+sl/6YPu3LFbwg7UBLYNoLfglp5n1Gw9O/xRNUvpmd1I5DxZS7
HOkoWcq4uo/ELtWn18Wo6BrNED+nPI+/DvC8IF2wALlsjZRgy2rlHuotip1/g6OCkUN/qvnCR+9Q
8oIu+Fwm0X8+C+sQXQJl5svZbfAd3sTf1KdipSfgkVEXE6GFKvBOmn4NahQFYhRxzcOd47gtHFpx
kzEmkrVQw3O3kCwNIMGbB6mXLzCLlo2x/BtCZDi4mDXqNhd94WtUekd8ThLkn2vA+naN3ru9u7cC
jYr6cCMdHluRoHcpz9WAQ/peziy5OHHCUvuStI6bEhxaJhLUVifM12Ycnsw9eKz/mL7EcYN1FSIP
GmJrZ2h23yw1CW2XQGHBgbpQ9rVuajd+zo+upehOeFJdTEju87KAxBWEPrIR+lFxcTl+TouxTygx
OnY2xE1UUa6G3ubN9BGynsNqtqa//F5xtFkW9yOZwiNQILie6Dl8lStJmPMwP07S7POwMrSvrYfs
gNBzvkx+vq3U+W8UYMm5dDACYtj3um/3zF6OoHhWAyiZ/9yVVrsBDJ1NPgROPDOcIZ/fctLLVDfa
JTqBYwiF9knmVI9RBS2Bm4dL9pX/6GSRxDgEsPZMejqKl4FpZzq4tH9BUWEPcFACHX9GMY7dxrAI
9is0y4iQOLrZx9deJ2jbjqkXM02SiME8KzpWvHee5frdWifk8glqdKR9A3Ru7XwcUPRuPuJt1rQz
zllC2eWrylP3+qIo6iZS9v89ipRAo97KLqw/FnD/87xto8BBKcNEXQ9hQv1+05yVfyTp/Xp8LGa3
ekq4OKGh31t1MqHvMF59LZOU5GwCLKVsPMZ45iRE3UFMGzgxtf22L+2787PZFSEkPLVFsP570Rso
bnDCrc6fK7iQzQ64cUkJR3aGm8nzVaMprG0U+PXNMQwbtI+yTQ/ACQeRehAMfN/YhIJ5cc5Bg9hb
GiMOfsTVJgsczt6oz5sAEw7yOSVDQxChnXBClRWMd8BQO3aS+3YkFkAZBsdWFpOwQ95NLARCjlTR
nWNLy0sYRzruAg1IfMA6cwUKsIMPirSbPputStE0QZgmcFTeZ9d4fEIF0a9kz+dPYcgAljCNScIC
7SZElYQTStVaaN5MMLFzUqWTTWNUg+R7r94odF84oEFHASYmwAGkp97Hj4HRz3qO8Cc3bBL9ARvb
don73YIfTH/44R620OGySADqlo03otSkv7CQuPXOGKZrAnSC0u0Aa5DHPTOk5VPKGTtuhLxFggS4
93bXe/Pt/zFt2b+B8Ba48c9FP6Roz989V9qDpP3lYRvGSbQ5AXB+d5001+Agbtf4WzkQKYv9GK6G
/zOx1s6e6ZUtDvUimGtpcLsHInTanWx25Y4MI1VLTBxd0ln9f7IOQlgJ92eQDYtsgr4DK5wgSAtW
xI98GtwoYaKiFEg6lUBs8LrPsckbmJoCXYW9ECKIaS5sbi2/R4VemRN+3jAaqeb/2LDA4vI416wz
emYcIyH/6/zDEo4YG5/iJfJhLbZXstorTXNeYr6tLp587eoIG5ZbJ1z8b/8hh2oO3oSmIJJvETEJ
X9X6AgkWqElB6+cYoNDBIw7517GcECJQzf3DlMmZWZYbCeQViw0eQfqLdU2lPUOnqPGXhExeSrLE
HeX4urRNZbqJhtwJevXdLD7onZN/ksSw1qy4RZIX4Xv5WOATe0upaIGPO4T3SOZyz0LOzVFCESAq
SDAzBGoREnZqiSANjfnOxODLOKlkiQjkLM4/MnWXL8Enn7KuxjZ9QrGsomIor96IQV/BmnEDptCT
V4Is9Jr6dhr0Oq09TWLU1l5wDckWfG2yxxfgJ4UJ3cDOpajU2BjPMF5Ej+PfhvpGzuG03DBIfEfH
Luc29Zpjf+gb1kU99dTPgkK6f5b2aTJ/+3RqXjEDXLBiDqoFyFNaa9NZDjl7WdyS1jSb5w6eBLmi
mdvd+AZWE9G3KOzoYQRzMaZ0HypID9NksQcl5W4NT19FaqLJMOgZTcn/vjY/bbx1xbzZqzi91dOr
FaFGuBsw11YXWp6hzLPyA7jSW7h8mA1tmHS6YPWEkKHK4IBIMX5+QXBgSNARmv3SOlpMdl2+QjHB
EMPjVwcU3+TgVdVfE88kjkEna9pPHMk8uVUb3Toiozg7wyWtE/a2dIrsiZxShZ6j7iMrK/c6lrLr
opRwi1hx5vfgsiSkQrOID3T4B+4eJuN0GNF/XnQk7W88J058SiFLCERzvwO48qp+0qaBkLPkv0fu
MyO0asDvqmdvAN9of3/M1D9EfHh5SzBv+3DtslY1IwkgrfmigsPp6y82iraYy+1iK17fD7Iwhz23
VCqe6YaPqixuTt1Wvnaor94BHN5yjhtnvcrmfGToVeQoa5UFYk8YVqB1oy8QW4ViWftvmH3NtI9d
oNU/nn+iOy2JRiY15+H5u7VVfjRWpNP/0ztjd3HabsD9JJbV5E/zZwWnnhflIiBqjVu479vhmojl
xBobiWQRvxcC+F79keOhgyuwaCQ5AqgvM9X0OWEKNhzWdPqLoKzgC772KvHiPAGKNBiXb4gdoJhW
XQdiGd7fmlUDRNhiLlA2v86USPxpY5zjLrrSJkbBMgvf3sI1mrrq4lda9dLVzAj6IUPUKdlk+ssh
WIVLvWQ4xW3gowwYRi4SzTwbdQdGrcjrSWLbPyHu4wkV4q4WoT08o8/XLT8hfgzPYnQQEOSZAEAC
ARzImRCpAnRr5qvOLZNB97luHRPUeN1pFATCjU8rS9D0NNZ1F0SvtHUnPEXGhc6uc3xb9GTh2qI5
8oREjQnHXRMfJ7fYFj/o/A+dsmf2Grf0kC7TXd0gjqlP7Q+S0UUoKMrRjMwVt4lOzx1g8+Zk2faG
f2cXgoXSmb1RQ4YLouAEqjNgPoFBMfgIblagsmGD6cPcdnlnt6I61JUWFe2HekIknABVMBPHuHEl
G7VTyF+dUzOuaO7fJKj8N3YpWq3WTx/vPdPHOv1zKwRfSeqe5Kl8dzOqRy1GqPK5wTR4X+zC4Tgp
TlBZ/FzBNJrMMxb31Cvq6A3/FhMCe9Tfy3XgVptQMyocPOd9cloowltubiixxHCaQXjF/FFGN2bG
e4Xdnlphp2HrfGjn+DMahYvgJZbTyyRbn+SjaHvVgf+4dZmaHdITtQWOSAFoBFubGGtyxqLQ7GJw
tKhlutgw9Mw/KGQ+cIkGty74rPeeQ5FSglfe0Wl4SzIC0Aive5ozGe/cPKk62O+3wkaA0ygxbMvP
U1FTG8906CuctNl4fNIs8nJcwYoZ1Lu6pwDfgoB3kk61bQo+Wj0am1Ty+DZ+FEDvxUIBAP8lPaqZ
n09OvhN1JTfDYf9o0vDJaK/c7Pmege+ktnPl/3V7af7NZN2tI9Y4kVkDLWwyraVS9MlXRjdPSgEC
1aKr1USqi/DZNYR9C152JQlV/X509fbk/1yGHn1r9J2FTUOHqxzrzdrDmVWAQuD7L3ufEmOXOvpW
2nLa5L2rUOqpfjgbJrxFt7culFoNYXof99H6GIKwnhhF9FSYxXpBlKIzGG99LrduLhkky9ysidY7
rCIEsAPpRSXNadITveMbrJ7bXugk7/wPAac75Mht7/udWQva1gEeREbjKCBLvIHp2GrFthMAFIjz
IS5qTIzV3G7IXugbVRzwpPQpYVLEB4LfJ31OrvoyGxIY/CKDYASm1qxemOzwmxZ+N5hHeXC4vAuL
kwFx5H+RbUVmkICaqRpBAlzxSRyTiwp9MMg6yRLK3ARZnRVGQ+LPrVvoq9AL+2IcRwSmYXwitmVI
EQ294q8L0jcYPA+7z4LT9gSrS3LDY790P3gvlHZ+4KkMG/aS/nSgWQT5cNo4otSrllotdgxuUQKb
1EUkdpTNFz4n0yd/tJlVU1VWzpULqtzsJrGyGt4ciXc7NEO6z8tVVlW3BHjqEOLiqeR+syFjRHuW
Vjr+1nhfZGBbnpV1ZsXxm2kQwoxlyHg/Cs47iHLlyAlKLFT+yRjMQ3lV5bEGX8lnjRpnlGZCFor+
O6pyChTaRAPsC9q6y5upgZvbSng8fOTqFbXHt/oebZBOFAstrt1F2DHtnqySVJv7fw+q/XNA5gsV
e+CWqCfnwXYKtUrCtRVubbjQYELEAi0lTeYHO+Q7P3MdY0xyjwqo85Dxz/JANUXYq596q/lEp5/X
41cdlJnErdI2fhgrvDaKbKlzb6WlBWl04GGgsCxe1MH2uOxYk2lssRRnT6Nvd9jKdO7QAPADH8OO
/qzuUC6hdQVKWSedYnFgOi7C7XGt9t7KwSEwYj8JSjatynQvNzJouNRmGvpcfshTU+2aVR6H76f/
gzaoacXK+CMqY1uPARCVsAmAKX28jFl7xsj+nVi/29LDx+6lGXv2yfDjG9+MzFlaLG9CabsYXJDh
2w2YE3VC8fGCZYQ5xEnmv52s0u2dUaMmdvyIJx5ZQfK/nqnTDxop35hg4xP9br8V6W9RyiJKcmLW
ffwGefmHFjCPitRSYlRnFf6wP9JYnFpUW8amt7ap8VQwmEn6z165myeEpEc7WHXsjjKXHkV7WnwM
WrwIqvKrl21nYbuBu+qzCoDkc0Im5GHo8aQroJKtvlLyI2ZJ89nKjzh65yF/FrS34alfZKPMul8n
CtixsUq/AiSERn5n7Hll+ebh4G0LEJnCB8XMEnhCwpA6iFxVEk/CqoESDQPmZPm3W8P2Cm7F3HWt
MIVA0MccOssj/rmr8ypi/efmh8qOtBv6nDDazRu7eJLpWMTubSAGXm+VFXE8rshBoWooG+fFkXMl
mkLzygzxuEXqpMTegfj1oWNY4KNdCh+sOFWhmy6vzc6JkNu/Bn7msTBlZVvEYDGXyX/WWYZCNADi
1ruphp4ERisvTuz7pHqFB08X+QnXiF+GselLl8+oehMP4Hzm/FJiw9c6CQw3WwosjBze5p+ib0vi
wgR6GzCzeiGTWlRkwwQ73c2RchyCMofBjRkZ17K1dB9XkXoaI3c7UYQmha/L24bHzYd6H3IO4KEP
JNbiFa53yG9CNrJROPFqxQZRMRPvc8nH6KMTYGq2hZHkE3inI47rzNnY6Equ7q/J7+61jLKlr0BL
WOj2i2xoy2hEgf2zhTtR6cK0ELX6C0aPFmtjXe365p1Evn5NuZHN28VeVCG1w5e1gFL4A+kmqNAC
k9VutJbGI0oSBu7aCphmEh2AkYOa5fSJOjMQd7QTn9GmZcVTwkxfKwBNH187AZFrZFjInN0zLQ9I
sSxSXU8p3C66TyzwU/ra4Y1Pzb0YhDPpoUsPOLv++m2VCVStMY1IJtpoGIoEWgIX2h1xvYnLtX9g
wuIGL0O/SBQ5VQTJBcekRX0AMBvbq02yKUNvU1oSM0MopXs7DR2SwelbxGERHrtZdQiNsBm3q6C9
+vTyNdewSO7Gfu9jAixrfnVqtrRxAp973AvCr3RP/JOOk9TQjw3rjaXZ8tl2b3kmwslMpfBT7l3L
kojIho8g8UP9BVzbeZXs73xrDg9IWqGuW9ntNjZaHezI71DRFKeCNAYbsX4XNlzLFZZlfCCjLQie
HG/Ps4pCzZ/WTeRBiV3eKrPsA2tpg1O3jx/CLhYFAKcAPnARtNOdnuERts8nlCMnn5uB9EKPHbdD
EcTjXaKNGggVN2mmM/mFjG0BNxrrQ+MgovPW3tnJnGMbnmRibA22vhyqZDnmQhRkqL2EmtLRYH/N
WxJdu8WxR1Z/ToKPuioGnEWN3w+O3+4YZdwJ5bT6s//MORluaV9Rxb+WZAY81xOJNo4nw+rD9GX2
5vWsBaMTftHDEKM37W0Z+0Ss0epERchcwB55uBs6LaqDSb4VEeQjB8XbaFmIe5bCePmEWAdMdrJ+
uQJV3Qhz7i5E9xmmRpEX7iLZCly+OmgQ/fa+2lFitIFEWNK3fmCMPQVonipjqSiLEAjMQkWaRj1O
HVQIolvUy5QqPWp0vSuq/6nTHyVSe8Y9Z6lTpC69AvLlCo/TA3sSIl+8hIT58ynaD2D3K0SPLKQn
j61eeRmwyXR01YEafHI36a2DoQhP4+3emwdK4km8NO4hkK+SDY0PqIXYFIrB8z6tkKHcqnXII+aZ
dz1oqaLVgZ0xrRts8Te+3OrERYp+2eVkVeeTdkpD7nP2qiJr6j0JjqywIIWlzcqugGbFwbxxYsFX
mRSNIANrB2gwiJpEmJ7N5qaw8Y9K+UeAKXahijinySpo3wMB5ugtUrlmXJuAe2rYELaiXvO84fQD
lLtM5MrQ9RmvTABLKWwiYzMH/INsmzq4fkZv/L+9M+639r3OBAafnCtpWO6lvdOePD2xcChfMJjK
HCVID8g1SC9bykqqmIhulHwDixQspeHitWlKFfE/xhp6I+iDEgnPLO3NvjPXZai0Ft3lK41T45pl
0YGKvkKOU046cXQvRk383WdRlx/DATpojbKbwdfWvVuah3fVcFJDTQHRcSCAWaALXlNv/dacFoJK
4crXjc7TI1srWh4PQFOZHHTTjM9Ti296frWS9cjZxD8Dd3VGvV4xoDUBVvOOcSH/MPn0INeY3dAL
egz38RNRcIxce/U0FquB3lH9l82TKEoAYHP6gQynEVuECCCbcHYs/wsLXpPImzGcWjh7hRIBihFZ
qE7PZX5gOaGWofaEGkGP5Ive72wvizHiX080CBO37rdOOvkrm+2J53ySV1V1la2gVEpYRWrRKbVJ
/pfVvEZzHm26k9K3+GD5+6UpBo0mxX4YqYu2E32BFYGalG2WZQicQTzNLNisDqrmRCtf5p5ECBLA
1nE1PdIIPwbBBnF3VXgPc678fS3lt/OTYTURsRTkwHhAmTCZCMloczdIuUFVSYza2UVkhqUB+Q0i
ftu+bcR3MCUHZoem89zdBRZYs+EH5xAXBO7/POGE/cITt/umPPtmlAPmQto7ntO3SOs2lsq/6qOH
7BFY15siCJKBv5EZgKeO5+887JEOvBus/e19QxChudg1tFhXIgf8eIs1YEKV4bvCpplm3qk+v/KC
niDsXHENTJOm8nB4oasDpdr0T5gQCNDAvxQlZs+/xoqaNNLbxQs3YQcB1AjKU9Yqf5oqdhtsr84S
nH/5gLZUMtAKppT+mjStAOVD7UhROEp9zEvDiyBj0jgogKdrtdVujPz6XC/QaTw4QlH8Dzg50mP0
Ck3ZHuiyov7Wex2KUja6WDkZ4OVUc1PRb52orAWw9PpdgxxALyVtHPHGZavaB3tyl/ASAbiFbo9O
64hBeew3VxM3j5C5JxJwtPUGSmenXmxdpCsQnloPVpSw438DOnRfthNyaOyG+hDx/JPsq97uPF8S
f+F10BAxvawgjAfnbLAipTgzuZ+afmBt4qMTiEaNdn9Izhnzl+LtNmSWMWXF5Lscxxgr0XRX7Izv
Yu5zXjeuwYcloVz4eAdBWJd9KlyPAA7SzOu2hu15/Bu19m+2LeAKN+Jz9Zd2rJJfV6nz/rTe/L4v
SCSXPW2U96zObefaxAgj5jcobVuEoH98xNbKrJyk5QoEBHrOpQFS1oGEM22h2QhR2yLRjte+RVk+
0OyPJYhP7yHeLxPE75R4U+/YB0hcspAZQjwn0CI1rnX7jUWrdLr19IeiTwq0mSDiJjNqrvwDaaMa
eakIP92QwvXqvyD5QhtauWT92pzdRRZUP9CgzuUub2zKsaf3HjStTanWo453E9HU8dqQCrkdmDkD
Et56rQattGIM8mjLeXCLEJe3/p32jiVIqJWA+SwjKBF0KPIuEb5Iix7bSxwmaILkDUnj/5WfoOLb
uMc0my7+o3C/qx8/uvFim3fqxj2VGSEG1cJ/B67Iouk6060wH6aT6B+xh3RGJkbTcNt3HnoLWHhh
qmvZa1HryFvlmrXa28NKGIHeiOxqlqRhd0pOflcMINTAr2PUNJp6+HXeC0GOGNKHiGoadx7Yd+XV
69L3n768onSU6aIeKd5XrJgBThSy8zPSNsFbUFNVQ5dLj/xCVXsnMrIOCPv+y9NPoF8SIAlG28B4
lDjo+PnIAg4TZJXNoB5ZuO1kzx5kq8Kus2crQkEvfbE7DV0efBdX0nmorgthFwdVBCqyQYHvvO+3
xjOjN65XPe67TSZpEuwXHj25Te1uWIhL1HuxIfcUK8WPRwYFAlVzKFOHxMSfEPv1o6zNVvBNVYO3
IJVufHhSHCM0N1RWsnVy4aNyw5JewJcELWwmfJwp9pqAu9DfD75QS8TB5sbqHc276KabDKAYdLVb
tvog+9dkzd6QKaVjF39B75TTcLYSZZElwdS2Pk3Bw21wmUi86Teo0Zrc/GQVNXyg9WOI8Pn+MxJ4
gZ8M4RcipWl02yzzXhOQKCjZwTXI4+wytcFxwYxVehJeFS3V2bNqrX0q0PZNAsy5me0QdhRnn+Gg
bV6KovP6sUfCJj7+M+q8BDtLFhMBoZN68DXn6jojYll7tlekBa8BVUc+httCdWx2Xm1njdz8/8FD
Dz4hJYpjMfY6VAch2gYSOWcBqMqyxZMD7chAro8/UEVLPdv69HmQTvmhkaemw/rPCTemRG5t3jEv
LbRCAegquSCP6FEGYzzt8EgXXC/FIztlxPGbcuv/8RIOFDhp8iwy8UuFUB1vHWHO/HcaQ5d2Gba4
qql3wuRiOms+Vb2bMO+4BvZU3D8y6GpnlmdmoNKE6YBwlYynhUQIUp8IzLmAIhNzFZ5dBt5l3s8s
5bioBCam/kwDJJJwjyN38OTo/9T8WYfg80gVBLKWpLYlsoE9kff/Uvj30ExsIuZwL94GawgYBF5T
j77q5QkDLkT0Tckh40Eowkcb5Oh2yrv3DzEND6v/A5eri4wIKM9XDIku3iGtPHh+euYtXo8Q+DIO
T+xiOLdrEdAzg05pDE94ZUrx81tZ1mTDHhjRdDjy0oiC5vX9enObOc8jxZ0jik6QmKoZr1Y6Odq/
1PMLlcnbv5KpC1CzipcCyWW5wPk7CSoz3nsM+kwmPoEBraCx6gpuh5/UIEcSAUMzl5Th8TzGN5Xo
hm2+/Zev4RaG0TdFGaKhiLl5QPhxOFol/FeB3ekv66vguML0mgofX97cGF54Ue+KUeWIOnOwEGHe
v5FojPYqsbq5XogZRQhPwm3JCFVXqRI3CPMjBRQvbMklRfcSlkMxn2hAok5Mwi13DGwejJkqRmW4
wvNmMuBcChM4M31eyFjZodxX05rHf+KR0KD9DWwMwWtfVWMi+tE+tLiONOB74AEDrhySnaIgcjBk
kumHa3irgEGRdHo8Pvl7XM+NAW8o6YD+GuHxb8/mggPqQlBe5YJf7vz4KfjOYjC6JixFYiE9z6HL
AO0tT4Ar2BBh/EnPhSNsCm7QYMQB0+2DXXfnBP90Uc5UU5YmF0fgKP2KNbWCMb4pUdSRIY9OAeC+
RG8Vze9d1eOGTOhIQepTeMzKWanSLlU6JAxqMGBB6LNtvocjzw5sfNiMocbMpQ/fQ+K6pwUBa5NX
Gura0AiqeJQyHdhT+3ZTMUhJIv7aHkgiWk96Xk6ppv2Nez3m7mI30ERw/Ukqrm/wMPJl3TNriQ68
0rKSm77ARRZhvev3Dd+H+5rv4w9xSd90H/uM0DN43zkNQ4YHU23QTx+2MKpSmu4ti9a5cuOutZ80
pAKuT7zAuF2dsLM/EAaWGW5o+txaNUQTEdAp8xjomqLtdz8ELvLZhq57pwYQl2zrYMCcmPy/Ydbg
v1bHyX5ZlgatqW9lgeVXYqEIyegsh53osSt7tyOF1cCjqL2u3NoNmDtb5/OyW7wBk2xJi5+3JYj+
DFMx7G8upxjT8wU4nHs4z7zzXRqhaLqL2ZK/MUGfJGfdRxJHrPwHKZ1AZXifRfyJx3QHhxvflWS2
52SF9Sd3JsqOxFqBKVPE7RStpqGIQgGnzXJ8533haTh4Ybq7d2d7r3/cx+6RF25mrCAl3dn1Z+Fl
nu+jJL4mEoqN7hn+obThrc0jEb3KX9Kej6fn/gp4rIAItCCuTr4n5vYCwdFiaYn/yWFKHWR1gp4G
5v1uLRdgHRei1lf/6FibEKkA+3Lu4uewiRIytEk9UEsjeHSJL6/7lLS9dsIwsRMetyT/BASV7lfI
/9wUPC9H8T/ZOKdk9CiJR+D7NGHFgPUFR6TRB+INIh4PDda2Tn7VCPrAv8ZLxDxROJnFvqI7D5CD
GFznruHOR1Oju5PxyT2BFeV9mYqRBlsJUKSApZ1bPB0Kw8UjhrxgX0aHTjc7Al+mZVLhqVeG8aQ0
HQ+nexje7nGMmiz02hDrJjLrRdDOXkNF+iRSWJ+sfKKI9eTFGq5XbDjqpAzYwMxfRzwi81vxP0M4
1gqP77DRixfNM5pE6Fi3KaCgjA+a5S8Ayt2nTaBbxkfaUMgefdCbWzFpk85KID4/5Ndiov00sOtr
jwGNrEZdG21WAVlIY3T6of+zw+yCLGdYh2jjR9aKL70qFrAEokkzxLGzNAFxGfVJI4zNpPMFYs6p
PvyPqOH4VjowoHE/p543sVEtBvEAN1JUCcIJVWx8BgP5EDu+2qLc3ZONj3C2xHdqZj9uui+SeLIA
TaCwzFBVEboWqctGV+PMJNEGzhZil2IVThcITQCYVRQdULfr3uMHzFEskoRazEaS1rJJpG0FpZ5S
5D6upwFdgJ2iE2PYN89xFrD6NEu+D9a1qRk7YoN3rWL4FCUOt+keHjHfb0G2IgNGAfnc3g6wCI6x
FdCVHIHSUpnZoyAHGuTHfYyjU4BOdaBwrdPs1SiONj9bIhzF+ouZip2BvGPglyYmKUlZaoMTDNgm
uZXcCNQC5PqiUxUzNOfnao8LuRdHXWs2xfYrbGOCYR4kbWaeQ1kauWQOJzq6IdXpw1EYi9pYhkcV
kmkjaDo/CA6Ea/Xu1cYMu+4TuWiObDQqwlWR+8vzv9uZ2OU8oHnNpuhnjo//mYcEgCjTDAPqyGJg
rJT/MxBz1tn94w9IWnUzZ9bNtCZJvi5xImpFrS0xfCoPrfJSfFq8UteMKdPLnh+szHwSomQzhaKU
kIIUPqkWA/+c1KsuJtLXcQAfBOlDmEzRV9aM0dQxxjPUFOY2Wx+d9RIz7MImOfbYbzt+4tR2H+0J
/X7FExiJO5fsjaPhcOQfv3yi/Y06kJJjS+rOAH3wdw+VL3/wDHDazdGcYB6dUsaztBCfsgJRfB6I
D0t410GnspypUHjmo1gXz4AHhVP/jWJhXOTXThF1MczwHhEfypu2UUgIk8w+NUb8j8l6MT4jYtSW
aSnaJF4uG7rLdpT11hli6DJYMZHgkvaynMdCeEV1/BMWORtSc4TrDFodg6HIPzfR9aUTcR7fomsR
K0GFGJUu5oxSF+DBv5DsatuxqUg6suDt9ACyQuePpFXeAkuTaV7GP2w02OJ61Rl9OuCD6TkQZwRR
vOhKGE7AlycXsTIpaK3PM2hc99YAXy3761bB81LbdVTfyFvtUeaP/qzA6yUAzesVkG3mX+ymA6Vc
7qKPJSb7o4kJ6RzhxV+JXT3fkJqz93smigry8a8P9nZhHDREPonGwLyQnlPnCqf6oA0wCuUXyyid
v8hxFE9FACj1ADq1xonSiPRPjwGEU8J76eFpMh109o9dEQ8dqUXcWxOB2SuNvkfkQz/CBGM6Vxwo
7hcJ9j3ItrG1uWoTauBAb1/Y6WwlN2rwLtfSbDNWqida8Nv7aE6HPKof+hu66uMeULGWWO0JrsIx
0GbF437ZC4rIt01cgeQtxaQWBvlIUws+RfQScInb9gS1FCR1JjWTs8cxxjsPWVSh+4T2hvaVnkCL
cmuSdrZ2wTUErBvntSF+9Q954go8Dlbs6ojwfeslLFMIY1axmUPoncY7Nyv8vrfBf10Rq17cn6vJ
/09FF3EgL+CxgXOSh2pZtrVES5U4CRLIKEvBkbKFGdFIyAHyXPVUrMd5UfH+vqC3xGHa9OdIBBni
wbY3lNBpTGq+2lYINMPVqokApw+wvumsisglT86Xy7+imkl+bEJYoPUSSWdq5QJ84eLUKAWUFfM4
Mw8O/BfyGQQUKh0lhDnEuxdVND8raDFj0//3PbIQC0tFNc1tANYGRLwJvv6ziJ42JggC/ald03OT
IW/oYatTzxhzFzaAb7mmWGUMNmWnPosTzwqbJTLoAaYMEBc31jJw42fR+6zc/6o9cYiV0YcuA6hB
EkimqySJaybicOPcPGykS6WrMmadAaZ3jUxg8CS4XtrlSxq2SehN/cP+ltM6iE3aDPRb0M41wZF+
iD8DcpNCSGf2yy1vrXolBLB9A9qSi/SNiFvmpvJoeuNvRA9Bou+o7aM4KSkhu+VGVxLrhiLa3QzN
QjHOVUBYaXXFkC1S2rtgdJR9c+PsnXe4L5lkgWe7/CyRyL+auAVT9ZZBG8FXqEXhE4WWuK2wJN1J
ufCvLWZN+wBrMGeK/coVi941fJpdBblNNuFMynT8bhrAdhrwN1lx9VY/+O6pkyed0vjEchYX8XRV
ScJlHUPO/ervdKeXN8jXe6vCcNvY7+HYMxQo3PFPy1wILfcmwOzOj6nw7Fe5otYyASJRwCpJHObI
br4G+Wc8HrfJnwv6zDh16vyREmCuw2RQIzRlrT1bgI2TM/2mXKUSF9x/xXi0fF+7Z5SwK1emqwVR
bSOcVC3X//eH2akbmbeD6Uxj5fZKSH4zoDn/PLZ0dD8T1CD5qmtLkXkuF7//xfNf6b/biJ0F45oW
VoBkUe4RGQi14/8zVsg2X22hSS3RpwEjN0f8QbBCnhKJhqNJ3WRNTt5IMUuCCwmVl/ceXJ7RIpgh
Sszw+NW2J2cnQPQXcVdzrmcbgnjUCY8L9nSW4HuIeIkpzD7uJVL+2rJGHbR4ABSPijpQTUP1Q774
E/V81LmxylNGz+BJbdZwptZdE4kYZYuIFt45RRt859oeuR+KRJZSWac00Njf8iqPFtsfktwd2aFV
GQNndmniljYe13otxpvwRoxWP74tUTxrFUsUmdYALEkKFyw9lawAHDBx/NwutcSUE0+jAs7xj2O3
XtURT7e6Yu6iPoSLJBo0u8zzY7SbnsynzPPUVbCWMQWkroQmjZoe1Jn0A9ami/50MtycflZCbVCd
wUByYE1AJed0Kd4+/8oteAwVEHXvwhwAwFup6br+xjbzgBh07/ZF6uTNEetgAArXmrDsp1w3UKTL
/9PDJXgZhUJIN74zh4obik9oefG95K+LORFBWax8Rsjiqjc41CLGcvtRI3FXDmJ1dwl92Afadacr
f8wRDfXEFWo4rJcDklzJK2DMLQXxdPdUl82kdj1UWXAPOi2FIpr65eQde7GfJ5RTUKygfeR3bRk1
6/PWjstlUYFQOezq41c1YqjZ2SFbRfApCgtrw1r5suD9OG6au5RTCesPMY0MoAndYuor1r/vb5+a
wqtwGqevdenzvH4FMwg0JW16IrIpN2pI2IUGiYvYSkbYWUMt9/uOxfstyPN/WmTysvuBVFSaA7A/
r4PTODrXSMIC5Zwzqp2mKUKjeMvWXeqONd1nw9kquWvAGORzpfE4beoPheqxK7O9LeS19Q9ons51
oJiTXj4x9jp0LWMNZ5hH3tv1DppaZpBVBePsNtMKLU4RZ25kmGqyfBqdmL8nssP1yEb3iQivbrsK
qOFC1oOpQ+2sWFa49xAB1O0Oqrr8f2B7WrvUnoJKLQhLe6AKwUz9WGnXUJljrLXUsRJ6DIMLP66h
JAR2wvXmPMNz+ipjctTrA7SJMecT/w/koCBq8MjKJVu9ECGb/sKEo7LjKNMn67YrwpGXKUQPx+xo
F4ucyCioXoJFu/CLyioAX6pT4tyyg0AjoNSbWH1LZFrFe2QE9QBwPlI7BO+rPoCv9SpAAQSy2QML
xRufb6gu3eMDvX4GrXYjWP+7TH0aHlChfOC/WTUGyTr6G+KXuaa9kdHs0S7yhH3GKldpGZB1GgdL
w7o/7aB+9iKLowRJP0TBitcn+hT5ISnzla+hQ5GUHfCn0HKbuYlgFOydrQBhLeY4EH6Xelnbec42
f0sbgHKVTkDOjnWkMuuuhXig9T9zXmSCtfvgHWPgozY250o5ngR53EeTrEJqGCkzBU7tge/wm27u
1m5rxH2dIXWytDVfDrUTmcLYNaLztjf0cySX15j9sRnMy8GS8PE/jbiDvlx1IxTL3HaK2irU3+LK
pqH8GO+P1U9TrLqj6hK/71a8w2pL9BQxUiqHK7LdVz9tsuLj0VpiiPGNsnz3RwE3TAj1ynpbTB6U
AH19NH7PG/NqGHa6tb4wl0lRYMotfetlbiLUiQ9hfy0CDCM6E/EERNL4HpmEg8mDhPx/Uoy/CEJ9
DSQtkx8EeP+WOcU/jjfB3y1857HbpXvpolLYYEKSHaFPmqYB8e0HACtSf7yUrsjts2qf9crIK7h0
sbQGwxHm0//3SVvoRPQ9+g2Lp/DGysucx96U3HeGOdi6T8QtHn4dNLXdLILfVa0S3qEuq/v9HAec
swrEiYiJhCoavOURTheossA+Xw1Vlj8myrijzC4yl3jh6eSugXvTU6sl92vwjuP83NV+n1QfPQor
eHd6gmrWmq6kT2Cw2XmxUPW1ZN45Lq5nXCPZF40z4dVFXWRlZd79fbEkkjud67R5QDF+hbZ8TjI/
/+zMGBEdpTF6TaVZIj4/8veQQF+Zj67k9eTXcbCmqNvGd9+MUTzZz0ZvAFR+WbcL+8g3Mdm2Fo/b
wS+jSEyFI4SDFmtl8vKmBPhhSGIpg966Cp+7ZC0C4WlAHhxpy6nCxpDvr/GSot75NI49aodoa6vp
+k8UbzP+lKCgL5eZBTAdphGLuCWEPHQ6fPgZ/eStreFUlSirGYcg3HiAW1XczzeMwLAnlV90tGDV
mfTPGaF132CrWO9yGnlb2lOnucHUSgU+LORSzw4RyYls2BFdg4jWIPEVRIR55ADgC+EU1m2H60Ou
DlcwYm7xmpttIq+bRf2jCuN5Y7NLCF1GJUZIeVbM+uFpGRrCqkALW2IdVJJ17NdjELlp2iXUBnVA
N4jy81Y9BWlKa6Sg0VvVd12emTVAipid6EcTleGmPN+JQqVNl3n8dcJpShp7K4dyq+JJs5bESLyw
doOkRNqUOaedF3bEHEUV20MH2XlyfHDCImWJNNfqx9QFqQSroLVMRC5/Cm5JYotiQpHmIPV5f62d
x18QTMLp98XarJb0U3JNT56LxlknpFZhKzQSnFNcE02q7+2VcYzy/iFitNlyvSh9Gq5DekJdWhuU
5hTTahPTT31Wv1Na0SuoPqaPRKQUh716Qv1ms2mlWi45Bd8EY9Z9bhG9mtIaXXrWr3IbV89OgmVQ
LoGXQanK5KrmZBB/9MJk6poJTJFh629q+6UNVqee2tbbj008KqCnP6Jek+qzxQ30ww8wJQTspNtc
a6Rln4hhJkkm+T6OrnuSFGle23pJIUiQ7X3nb7mxviV8WFrLzJx4Dq87K8Ur/mwa7sPrvE0kXx29
9tINtZCznoRpq5HEgUipH+jygAK6Pae3R8rMqk+i/XWalY6lqWqpQbh1KeLcgobm3WmuanS8gz6d
Wbzxv6MigE3JdGf2VyCw4S2a2On2hM9yjbZ4ulpK5KWi4TrUKmY96dUVQY6JcgwErIVqHjImm+Yj
kMFc4oAEfpbdoCd6oXg09G/u616vW7wwN6b7Nuclny+duG0ySw7CMNDEPQ6Qpt2zrhvtKZkV869g
Clsqs9x4mHu0+MV4RztORQCJkXfQjvDpvBjIZa3EaZ10GKOyRUdF6eUFq7tl3tl9XDcOD9Qf1h5D
w6fMa+JCR95JlaD/Kg77XK88mrUi3SgIq8Xz4ODBVvPrf1zmEbzo23pnLySTBmyPz9lGL2CoHDzc
2YCt+rTBZEg1fchTQ8WR7O0DRbjSb7g7YgSDPG9orVq4mLIpRqURiGoARJExiC9gozOYetwHJ9jR
uov0b4RBc1GhZm9yVJROUotBDl201ws/18EzJDA+T/29DNlc3jht7+DmW9tRAHCgIicu9ok735lY
NnngtpGrZHw6UQfnGe1QqwrxXcqvf0Y14iFrbyn7HqVZq8b9DEotK48/WwwkFYYuFyGARR6jCRcI
MzUtsWCYxgkz+qUPT8u5heNdhCgzWgQq6M5jQQb7wj5PPm67QQyAvmfzVeku/x2FC61Q9Hs5mz+i
xf2/w6JxbbQBI7ynHGF65wotO5kwQ7Qlil6osahQxAMFUPcyLKvJaPjNhCDIFYDE8HEML2M7Bxay
BWfSu9u3JHAdmQYmpwbPDf2nNJbboMUBqJBUSBuciIPp7h/poIZYyQoNW6D6G6iyInyFd+NtX0j6
XUBiXgXRbrTGfr8xrwYdmCKIZVhfbya0AlLktSlcTmjexsxRV1tpTXdKosdUnom0UPMYFe1JVGaW
PX/vunMRpMNKYH4T0Ca4yn0K7okMW7x1eLHgh2G6aV9llZfiLqFutUT/rYdxOYDG8YZq9jr39fzc
MYyUdX8w3VE0B42hZ9CVQu2/VBD9rJjl3MM13XgF2G7ZqQZS9uUtg8QzcfTcp3oM3tacjA2RCKd+
GdD7daQHZHYMvd5trTxXxRnXjqid4xEYOafZAZRHwj/5C91skb18Lwcc+SF4sXQdgWYl9tRJlaT7
2TMwufnZjji8tFqtDPh+wrm4/OGTlowU0QCtSKLANlgehVxYbkywoGyptz+75y553GJWXi31Ma+z
ejWwJ9F7MJu9hF+F+UUwPdq+95NqOyjWNYiZuTnodhdmvoXYMGAVLlI2jjEFYKzKUOkjCsz1ZkPM
Sx6s/H1RxhsBh0IZIEIatT0D1kDR2bw5zjKvdU5eXtsiYqqWMaYrPawRgOo8zoT/PjuiFffHl69y
s7yhaSGytryRE2WkJVg5q2KkxstFPgQFEquKg4gKJneP+R0En/oKLuQjcqBXiRT31Xcva/eja5wY
V+VhoYKPD9GMOZdarFf3D/3C7PfV48o9MLxCxndPRymbEm+2Q7DBXZ9vCp0IkCgFxUnGdp7CZ5g3
9fkdD7lq5MEZMI/lcPVTkV3V+lBfNM7xfNAhTtZ/kC1NMOlOZH5tq9+T75Wm4ZbdiP9mzmFJfYcD
SRHVzq911IIwxquq9RRKEnWWGuqny4jY972h/s31uXTh/cY5PzeyfFT86tBbrxPI3lWtYl6VinAB
I3Ah0BgVqotxvzRV6uOP1AnqcS9JWWmhFgDSx7421+Tq1hvp1zY3r2XNJ7YsLnIPctSGOLQ1Cqjo
Z2NwRZ/MMTLeTrb8Asn744nD/7CLPNEOMWTsN8XmbjsSUzyiSIp8RDvKd4/vueeaCFJNlPghPH2Z
mKcrkekBjOvevdYPJKDiZVIHf0524kkwJJj199hcfP5pitlwaZc51irBXszzkXKowoun9z3QSa/V
8bhLhVioRZACd/I+RLehdov7wTDq468HRMmmWoVvY2ZEs8rUg+R1M7UyUTMWxL6L0dPtwICFvo7W
o6wtps4Gudm4U1ItKbWGig4D/6fZc+b9Z7+OwLmIxZS1osFmuUzHn2vZ8KqtcLzY4UacTVXBLdYK
2cCdJ092CePUOS3nO5/mGPEIcSxBPom3TRMEzGbvugx/s2g9UEAySLGqwiBvStccp054l2gahLzi
lOhgr2GXcwsP3Sk3VLisgpxYdPoILTEtJ0U8rcGO8NHCkxFxg8LJA6AbFLV+eae3n4YrqzpwpqbV
JpLxUrvfRqoqU70HGhjtAGknE3Ug0LJUHY0Nc0JvEcu5C1bTpMplPBl15Tuamt3y/8JZR3DfLj/L
kG5xd85u3yj+Lyj7UVMHzseZfamgFfoeo95xYWvz6Ii+iTzHWtsFX8chUGCRIHuN8n+p8nLx2gi5
eQfZT6CE6FNSeef9fHJLSEIwKG9tXt1J8arjTI5Xi1fPIgEKJzczPZZAUENBTprHx3A5XrC3Davz
SQNYTwNRz4IfIDWdhZ9ZgzG8yWFHj3wSqrquytdmQ5Axd0dtcS3twgAkreuW8lHlwqP2D0ZugR3i
p2/vYztVcywoKZ9BIsxQUM84SAyaj7onzIJ8w/PNG3WnGA1LENnS2Jk6f0V3+g8glHewuxSPQSkL
S3jfcxaojR6QkNpwElKophNB9ypT7KJRuKUNeL/XDT6nk6j1mQvqxtKD+1ENFMsizmo97x/dygur
7qUM0h7rV30NwQJ+nFimfHg4I6LbJ3aGdlX9FKh/OxNd4/qmrIZST+nFxAK92Boc44TIBlqmwXJi
60/m7T4bYPM8oIqfLTEiyo5N75l3gys4Vk6Uc8s+MRzEdKsWf35uvVNHYPHq7WtHJwwADB1zy/Sb
Z68BgS4H7k6XmvC7JtKKaW8CEpsKOpy341UUiPfVH1iNjEkfGCuXbCTwYu7swsr5A3ACm4v3ZZDv
1OfBox/tqlSckvr/zsnFrKb+D19Fe2wOh/DwMsueFaySDxWmj43zSUbeQ1ULSgHhnUWyof8qSRRZ
kcyy67+RIQwmIhLVS/JsqDtAPfqGf+kBY40yRH0youDT/YNkcOHF2NRJkSgAE9aidx55qmurQbmY
xV5GQOaDHmV3J/LfR1kKo70WB4peSuW9+Am9/kMhdaMrwyu/mYxYhtLTjO5BtMUr7v28usdyuQbN
Zx0gtXb+pJRApfTdAWng6h/FIbuGK8m/ER1eHvpY3jqSUeu45Vl5ihwnPIgO4kXPtz9UrcEuhJlN
JuBeANbYv6d2po2WoPrJa6UgsCzpMz69wfWQJ+DcCGGzj4NPL/5k7Rfd2lPWUCmhTVh2c5q6CJm9
v7TE5iaBRmWYUSITZC0ppNIZ57Z5zcm2VPsRTc+caw+a/QDP7cCs87PyyyGQuwRKnTPAY6Smk9hj
BVuJwrFkFxoxK3ThpURU0ZSFUFJey+HA+AN9woao2DsB0mCp9vShZBUADnOdK2OTKvDwtvyk9Lob
vvd8eOWFQQKp+7+HWJf2VltM3yh+sUlQR723Qpmw2KuLO1lZpk1r5v3eiCnfyv40KguShoDDXpuS
hDBXUkTj+7q7P4yo2rtsgGUklguJh6B3pXz+T5BDxMHi9UqF3vMZHHR9pu4xOWwzyVEv8ElDLJaQ
Vq2N9gBtsipe6Zoz11glPFj6IuY2QFyI1iGbZvohZdtLeQtTdZd+gK9PCcvn+KR+cigLVjYBGifW
LKC3XR1zbC7nxwsAbBgPYfZOa9n5L5ipRD8gWIQ9dx4+qvlIG/3u4IuIP/meMq/qg4m95lEEf+eA
RiVYmv/Nbiil95bO+3eKRGLfLCmYBQ8LbmsiXUVJ8O5mb00qT37QUe/bYM3LTgXnZ5QH35k5jBoK
U0kzH/7kzQTDRF4Y09F4wPq+PXiP1S4a+v8///UVOd7RxQZf7bj8OtCu6SLlB4sV20JYCt8Ew95a
oGT1RsO9FkDgv2EngPJmn5N0Pfcb4AdL5v4pPNbimwXHAS//M0+n7lls6TYRDHZUP2h2odCBmjYx
7uejraA/hgQxV3VGLdvuaXSaLNCFfvX3GsJz0SS+0UlvP9GvIZq1RPxJI82eSYTdEeSZFWNJ8/uY
MWLocN0FLRoaIwy5+SlmdPIWHdRolxtxJNmNkr5DsxbuXogtzGCTl/2m6Ee4d6j9ElgE143MzPNz
o4IeEOowIV9tAhRUPVf3tQJRdgKqvEsYzgOeU44Se3fz6N4W7VL2c+0s58upckypaSuZlRKqGE3h
JljZ8U3bVuiRJNCVrM30VNdc9kEPqMa90xG5iMrybiF/yr9qVH3esk5F+K+K9974vOlhxPgjp6qo
agoFn7RcygLQdDebM5u1laNMa+GT9ZkMmIdHMixZW3vVY8hCQExiS7pSXzW07MPTygb6pPHNH2jN
8Rvbu/WASbcG0hzYRBI8Djyc1Dclvo2IcMcV8r9oGIKOH8B0EJ2ga12thwHX4RN6WLOc4PZu1Zgl
2AY5Y2INXRWHh9+HXo4tX7gqQiG51eDa1/ITzjEBmKn2M9g+db2yoWnHROKIcSK/aFMlV8RO0Qcr
g9mc7aT84dxhzrOyw/dtxkRN+aCWFQrQwQGyaTzezfvKxZzpeKHdex/1RQa2Ynrs5g5PDn48tmJy
TQR41CKkmvazNUb+mtYoEUHVINQezdq4F9Fs7KDF/pz2015HQ9UUrDsJWlQqVIzra3Dz9M6Rj2Cq
QscJIPpf25nqpAGVbPlDizvpmuts4spb+eUt3HybYLrK7/QUNTxR1XTSes1rVYC3CcVHY5/3DEWD
39pS1l9C1J9f3pGMEJU2v8NF8TQ5b2r6v2+7caSQAg38T9BqyrM0rbbFMmyl6hS9Y1W8HigS/P6c
fQjn2LOWN1EO6jbVqEADTBQ7en1YahY+jiPX/zOC+rVDINTQQuXwTn29fbjyaLMxdxOXYKrg1/h/
rhVdjPbaiUXDzhZkB8tmy/noER1e6zPiUpIjCV4XPZkOaFp0zdmXIlbP52srHXzHpVlaS+Ph7KYK
1jA9avuxVCFU50K+DlpYk+4Wv7YNgdD2rZtv4Xd6BWef+U6bdSmn6cucAmKHIvP6TOe9PdOnUU8Z
qrob8iOYdnKGmgnJHO0UmjlfmEHJYZdfDF3i1ljCf0MGF4Fdql7dvKKDewO6dWuC7hMJqVaxyoH6
2yzFTH/GFCakMT1dN/D2FSv4XMph5b7Gq05MRlu+Ra3DK/7T+YhoSMHbJAtymiTL91lPRi3+BdcU
x+UaOU7ri2QqcdO8GfLOGFydosmD9CyJjfgJXJQwuEbpFysHTShhdhJb6KLhH0/oYZOUr5CR6KrG
0oRvN435bdGCPwpG26x9fsttjvqNVlFy2w1nkx39P1cvfUeaKrlOcE2NVAlmyAFXf2ij+vT7ikeA
delL8HLTVfc89S5fm6M8D9bofesVewW66mBn9hz8b6XYMg10O9+NMH7bLpNs4lb0X5E9SqeODmMc
Np/diHl/1eXq60xgzIZTWVVGEHHt1mOknkahLti7gQfhM8m4u95MW3W3Xu3Jz+mA0FT6P2PkLYsj
8slnaUnTvTJPGkWRM31vqtJkCyCdabGgIBLaLz8F9kk0EUVNN6UqtODTb3PFXCsE9hPU/9jlW1oW
B6NEyfJeFIiQpQoBK+ivIj2Ll65JO78SFwgpTxgnlos0hMVj1II97wOKvBzJe/kyNWh3DuYt8vo/
IxgWuKfJ3GVdmFlR4w+yEK90BMy50j4qFZSX2Awj6Dw1aFoFrsuDA7+p9B7D4cjh1Bo6yZL7A7Zv
B/VrBmPvrH2rza40/E7YuT3MBe8+Jg3gYwkPekeh/3CF8aURJABkQXjzrYbJV9dmOV42CLklqbdy
c7WIQa7HAMqgslycelg1nf2fwOW/f34mDQ9UHuPh7SIvl7DCKJn/sIn12USWlIFXGbhkvMff+9Rj
7nJYOjB5OfV3tG75tlSYM/JfEZQyQOP0GNsc8ZeGOftdqXuAGruQqBkubzvXJ+u19kpx2YjEfkVu
YVzed7ZS7utisZmbtKR3rv2XuN6WD+tlcjtA3jVYAu0Y39V4JATDV1qj7RbTFeEh/hT7/29hDU+f
tbsEKWaQ+vMXE0gk7HgNV48dcTmJHn5bJX/yfwuFtX69Cke1nGfNRxR1x9QTGWtK87UhMLtuVww9
HvP73yM4eRGTnuSKiel1dcCXQvsjrjF/7SnyLD+8Wuyq7nz+kdQivhUhcuVJrr13wC9cEDw+pfkr
EKWF+uLWRQEzlfAaln4Xdrz2wNujSYL71CsaLPCwvapfP2R+cVYPGn+5WXD6gv/LRiS2oHb83mhm
3m3t/3UM+W98uzpWNK21UwGMjjU7jn1NgzU/z7s9hX3cMdTyX+YlGPN9q7bASbn290DeJh9U/7iR
fQW2hgydvqI0QQ/+zT48ZaMj8kskhzS6chkstZSdpHhROoG2m36YVj6GhgqXMB/lT77a1nRnr/Vd
XiN9aDvsvqV3n5bfFXob89Oco12odNUOHjf7kxikRdho/Hc9/eO1iWg/2JrIzuOp262a4I6RnKQd
SfFa2V+rP7DGmgqTwYxvneNd0n3Cal9y4XSkVXwlvX3LSaNPNl9SAGWlWTGW4avG0DSPhE5whLJB
cFj5+1rnVRbq4e0Eqabl8Bb1vjSnxHLtgqRg/LFZVGpYZU8a9PU2NDx+9x7Fw5yJhbblaqVKybWe
BOsE3d8fOrPRDW7ZTkBnhH+JcwCIp6rMwV/1wyNesUZLRZFB4hnvitE1YDdxvymoKYTfwuiq6t3+
5aleJ0Fn+GE/2/38ZagkbMSQRQwLS/QFtvF6ZGsg4/Q8RCTGcxQPQQ4VgfmV7EppKdGVTTF3C/T6
HSZ6A05+8zKRDc9hNRoVPJdnlNPsSBpTjOoyZUXInZHbS3rWuD7OdS+TfhNIM5+YMntVqACKmfDB
d1YnxrgUHm6xUE1ch54n3ctoxnntxYyqzu4d1P9hXBJAYp4pzFkBgtwgjSd/kacQ4EfHQx7MBzJR
1joFeFb5ux7d7ICFXKdrV1gtZf7bdUFJhz8KepJsOZeF/zre9e4Ph3QyFFP6wcRAgWThbrGq0HUB
9ZgYCVf1519R/kQEVzT9Ux0QXtsHus8K6pu7AYlg+90pgXhIX8l34wd57lU6aUXqAq67wjiWVvcE
gZm+6sUXC1C8DK8GDKRkksJiRPjlDZBBHey/BwvcpukZSbQvhg9/RelKG62/PeGmpt59s44YDgVK
X5oghWjqklqGQKnnk6F0V5LpfeAH4bcPsBFIcE0RGo2PMrXuzA+Xpulg2bOw6nCGRB4PSDjX7QfR
ivZ6m0csRVINB2N7tVPDqyq2IKtI6lzir9UA6E95uTPNZ+jfdJYSDqiQnZscjhb7VpoddC0PyxgK
XSnjsAHaDTsOMyURl7rHyD1XsaTMId8q6dfKFkSEL/I9Vn8Yj7LYgD43eUBPJ6uMYPI9NrAWT4iS
x2vxJKFkTCmBqfCjsyvMeL9iD6DeDhrZEDSNSXrtP3e44FHzey2ZXv6un6uoa73rIeEJsLBVBoc8
1/p+SL73DjsWW8AQhTdYsKgiJ1JekYvYKu32wL9kIbNFlPbaqB6rTMXDKaJCQXlJJoQfhJ+LqL8/
ih0C7ywDj3c82Nhu9SZ3qKjssXpL9j9JtHgVuG02eLrdWCAMm1nQ4di6FKTJ4NiSVm2VKcpWDhJS
EKrt/kD4MQeIZX4rAy1BjUyfDRfR2os666h7JEeH1u6PC0rhBClQsNIMYp0t35F6D3Jqeq3TvmcZ
grj4/Di//ue1n/d1IGoZto4x/xnVpbiEjtO4txFoMLh7b3CD+++nnSMA99L1m73Id1sTslpyDPOe
dDdD9hbQWKOzg17kv5QD0td+2v+eQtU79Zqk8tVhLO7bZdSCrQYVH75ylITty99YAeS0y1fiNfBX
yGYDtc4ynsMU/6nBU3YqGl7K0Xrar0rNRdIBXmfDIRvVj3nsd0uOpVxu8jAT4XOiSlzPaGypZhu2
TZpPZxjT9eQThe7NdDzZm+k1n5OBoTtB8VfqSh+2TX3JAwwD4JGzSJI5ptkYHj4A5P8Bb7BTYDO0
pE4mqk1QPLA6hlH9EGXlXpiim1XtTqTD3JzOEqwbiSLvOANJxBKcwTDn4tjb/g0MwdmCxhZa8Iyb
RCCqvD8lXhvNN3uYL63yNLbo7mepAXKP6LI4263sXcGVhFznNf05a5XZvtfYx4mqqaSDkkiYSySb
Z4bKbBbaKP4RlPcqYZP5MS1Z7YBBrlee+mUuAVthSDtHbeg+hfNQ+JdbRBU3Nu/Ae89AVMpdgNIv
1B/lNjdxsQggOgQLyTNlR8kOgCobjOSaYZ7Yd5N/Xab62BN+G89MoucPjGaQoMQyfka7PpFym2kI
fGPhZvQTYqo9m4lIGuVRjRcTQiLEGbIst2Iqyf1NLkNnRpKzTcE9MAXB27UI81bDFbahaYaRi76k
P9YC3pzweU0KShMlF7Y12x9wa6OP/5fIXCcJwhEMxSJNp7Kml/4WytY66c4/DTiGcGrhYg3yMqnG
ZU7N96paYc0axzw1jyA5Yk0J4PRKGcssog3NVNnE/z9qVyoPUOuvpeGMvKNucQcvO0Vbkz7Rvl/e
DkAafWyiKSqN+wX4dmh0AxgldxWKB47hr8mF9erH/GUVi7iuuSKBewJ5prHZ/tONjm1zmRf4pZTP
NkIY9t4kGdWqUZ9k2/Ku+VeDgHHI8F7qc8o+g4BXMBrk57Q3pkxX95Olnta9qhyI7rLEOYrGKpI2
rRUSswjXly/OhlNg0D4gOni+cwH2PX7qMhXB93BrSfnX7D7IvsaqBxXoGX9lweB5i9L0IWeTHy6B
ev477Z6xZCBdtHSkF+5SehRgRQea+iAEKUUle5B18K4HcjMWcp6ucyh/GIdQgO94aO5scOoSPj0K
gYR4do6KlcWSyPBZu9lIlK8zF3u2gqYSisNLN8gM4o7soais6TnsvLZv7jKAz3fpso1rYOTljqnn
s9O5BjzTPaYD/v4+X4L+4UJBDGv5dTb8Bxc68wDMsusbz+OgTzDcjM2czf1E6iR9OP22/94NwIqy
2n1y3WBLoZhyB2pWsWDytVFJ22FBUs1DIlUwWSuI1LDBd1xSaF5u1XzvO4SKxQMcm/FUFoulVfWn
KQIo0nPzRqq7J7Wfob5dQLFYYBjCFPcoF2kw3SR4xUoKu6pakrrjX8Qt/MFicdF19c6HpE8njqj+
8kyb7X2uXwCThHr15bPA3lGIjKCC6V7UGCG8j91wgj0DfRdEEqvyQJK2fu4gVbLXekDWBuJAY6FW
GXFdte/CcZ7srkGfNdrW95MDEvsnXTJSEBlSk0h+oe9iUThd/BTyaCc/jG0/Xx4KhjeF72Vwnuzp
gEzdOQq76lRKQ0p+a6MAUo3BkhUCJ5/s0AmzvCWHxQnvmqTFHB4P2MxaNHPE2eRkYtJ8dAx5CFuC
L2eAE6eilH1B/fcnC/R1yemRwGTuE+pU52HEhbE8ScMFQFI3DVLMwACGYeFsqQAEoM00knliwJhi
aScmLeBlUBiWz/pRyyD+m7YDoCx3WYLdCkDP64F1JdPKE08Zu/SwRpCsJIg71g2cl+LKa5t8y9E4
N+DLpHYmlsTr1VKsSksaoRqEtMhtUjq9HVgb1cve7e8ML/XDrj9hueoJm0HhYboUTRtJ575qdYtX
abGq+pkBwdOlVAXmOEvfn/xm4yenXaxUiDHEN51ErJzhlGBoGx4sOU28Ag+cg3yZJAWAQJOOOf5z
eSwShq3crPYIWlvsKm+x/mU7NyFEnmlwVznZ4VpB+OVWzmjvFqH9e+9zqZxp698WYsHCLU7y4cAX
Akd5uQBF5n1viKrO26kNOLUFjd40KXa6IuxUxffyE52xvDVweBBBc9TpSxAJOjIDrei1Bl5EarFl
tTUsdlp7K26/6FeGyXvvlaompbFxQAFZj8HILkh/3cp1yaQLV4hVJZMuJ9my6ctoKfPKpNBm0JiJ
4v/FBBAhFSvyARI+eP13FhligtkuM3JWhxHSkHQr94EGZtGl5I8xA3I7FsrMKGbg796e1r974N4c
SNTe5If1tXp0sPQ5y9AHGZDc3PqoIyHyJyy/6k2Fprz5zjlrOg1bacNJeeo6RcPIQmZxcAKGzpz2
9VRPXFocEIEVxDRziefUyBvZlQoq2grvnPzoQblHNPH2OhAl+Vl3JEf9x3VC+Yl9N1pWAhjP726A
Gozl3aM4MF05BZ7kbrYTNKzGnT3PZKjD9N2LZFFdmETLRtV/87fjZlrxHPddmN1NOyi0FGdOaVWe
yfXyCuO7sygsB53dtWf6NaQ5ThY35EO87K4fmTInLFtVs2UgWuKxM8KYqSiGpLCxt/f0z4gCHg2W
hwo2fuBuSPWwiBuSoA+vDR0i8Oleeig+W/BJ1+Ktjqp9+DsMgJnQ7yZsFsCuXYtcaSTZS7xsD0UG
ZphRHjNg/ju5KWLk0TVEKMX+84817UG2P5tsE7koG0a7ExN8UxtMDLLPU1JybBk1lYX8P11Q5Q7j
acTJVhZgDjf/93VcOuYxtwBwshDif8REpQFW+lMFqp9iD7i3S5kKB8cDDFlUCt8oFtoPUCybKFzU
w6CrWpy66a3WeCPNX7VJP0ygYYXoTCJirFFkmKPfdYknzicF3iurK4ykDZjXt5SaMnc9vndDqWQo
Xbt2UgH0QWMutI32Cq9yfQhpWm31UN4zTapgaFjfp+kSJ2euld6ZTY9o59j0x3iaKNg1wd9CC+QD
fHF+JXybqwRyTHAeaUBqsXu9a9tuTwbI17He2o3gupaR+9rNsU96oCtLCjsywY4hHDmXKTGJ/bje
yZgdQM3KTwrISHUUYOuoxxkpdnZao+Uh+/SOznjC4WnFGYobtxHRe0E/Hoewbf1rz/QMsKOx4tQv
raArjIp54RaYQFrG3bbzUszcjkTcJkFAzNhO2E8YboE68HvW6H5nksLMyqRxwd/TqS+lon7EHzbe
x9+5ZSSJ2cFJg27INBiRzs6WH1efcLwbLm3bHwv3sJBZBiCS8Z8h0Ug97Yq5A+y3+Pckv1A9y2lN
TXAeRz/IrlKsalIit6HKEfmpMpqqsjt+w7Dq5v7tong+Xt/gqdg3LUUqWYGatcqqjVqM/0OpD4jZ
ZIXweoQAIU3hlRK4NTcHynPhabuuS590eSyq8DfY39v7hFDPl/NpB2S1oLNbBHm85YVFGYLEd4qG
5Bdz/IX3POj0SQO35G0TTK9OsFd7oj+RJBEZUBuiXMFAdUG/C+RHGFgdokG85WNcFbS9JJlgY2Ir
IE/1nSflBWEKmPVDg4XGm2Yp1sYVXKVT9CvW5deQSqk6Uy9KU1jxEWoiI0MGI4736d3l/HtxDtWF
M4QmF4GPBXHdIvEjnOcO5+SY7DIdSbeW0rqp7iAXLMmmNX12X8SYIiVgZm3j/vsJKcZEK7FRRSKZ
0hVFdbdcu1mZtO0qm6z8TzL3o66HXQKczvbRkIr+GMHBV1e3NBwfvfzKKREWtHfLosqYxxuOEfbt
rnq0uX9IOcnBz5+AN5FdGrpJQdufmc4vXJgZ4pu5bk4EYqNKr6o1NAwTKF4CKGr8zlO3wbj6dBsx
2y4tri922d1tCiafm/rkJAcQrEx1pB0YK1ZozFhRAzstx3g0OtTf8Kni6B7NTe9VCUWM1BHPZFSq
6OieqvD9Ihr6um4qJJDb7JIiY5m4vg3ZuGg8gASW5qY3fLmz+mD0csL884R1Q5NAY1cWHSXGivQ1
OESmsMmBGrGVIcGTWReHwYO+oj733qsBwEcgBg17IrMmL/eaLaYZip+2FmqH73qLAnJp03MceZDE
vFyGX5Ei30frTYYWpw6dw+CDHDQrtVSbox7EWzuNXh4LFMlkgOT1jVTxXwwWIreJreTzOd7l9GxH
VeZVOswtMVBRs6eY5LcprpO6FV8Mm3ggj7HaFmeG1ChCmRtmFo56mlhTfjfwPyr89webBpQzsWux
iOlgQf/JD4btobR0IWdnBXYG4PqGsJ/1oR6/UPh4wbmfw4GNSbQQQGPcSYmXY0ypb1eM3tT1LTth
YwDJPlQBbeys4b1qLbusJchP4etOtzkI+qPm2CU/TcyaiE5yd/JIP2v+/umvAaXyc11Cyl6k1O0S
ZJ6DxAYaJ6KGDiWgPbgRW1uqjR/SouFqluXSJFxlx+27YrWJWJDekfKLA0HWMLSNynSJp5MGEeUu
1Ct7aoEaM4rVqsWRbGNg3H6sH2crXknAydWOAoi/qlLZOnePkY3rocFR22AbVsNzU0NbZyw0fAXG
VAExBqos6LXjDZZW7jCCi6OnZWiQUxL0gYL1leI6izldLmKFmtYqY+uk9BsE63PUthukm/7R9BNo
Bi5T7EqmoA/WpfIiGeWxPmbgpbt4I9Uo3Jri8Py/cRgTeAddjbDs5jMgcs3rIATRPgvmbCs5PHQB
S+0TGf8+O0mmb8my4TjwZVS5c631+ug9i+Jdyu0kQUojPzX1JRrHvmIzuePj9SBL+xEdw2lGKsT0
TWe4Z/Pg1qiv5OxV6slJSSz2HdidLhk9//rtnUKEJXcbK9kh8+7wLHMdxB2GsYMjQw/FMmTjKQrQ
rOQ/RDesuNHAfGOFTjoxgP24mJTo+z/wYwtRISP+XdM+NnjJYvQUJoa+WhgCvYSc+vIIlvPmnRub
Iw5TZD9rT5Ll8Yv/TNaaaTpKAOi6yos1PH3tcuj+PiI37GNVT3jXcUxy4jDyzwvm8myStuF5aog3
ADeUjb3zgd1067XUFNSaDdC2Wz96gSqaTxqWYiNo/4lFCYiSKtA0fz4VjtCzsXx7BMcaS+fbcmtj
GO3ZRqGgszu0NWyKFdamCiq7HLL0x0UmMVlevjFpTivKl9kDzJcwfDQiA94Z1iWbvAfYQ5fIUKab
cDweLWaWWozf3MKdT84aWR40Od+pXvrLV4MV8582ueQiC2C8Jf3B2OkpFlNuNBydrVSxkeASImB1
QMwmXx/QUc4WyMGrqhtlulxWJpzEHjFjnhQAX3p463aJOXkQolmtDO8xWQ98+0dolVL+UzpUcBf4
CW+l8sRkoSXGW32jO2rIIWhxpTReuRwvUuL1VPGXkRWR1SfM8Kiv1gzDX4dcdfTaeuJa41R0TMLl
JOQkRUrSOG+Z+/545YOwf8TfQieIBDXfVoT/qmjGBQ0QlSuyUtV7DTUOEWQz/RgilFUZdQAtrI74
n6DLtqIVyvswLzsGExVIX2ibpdeUYzYDsocgr69JBrWFpqZV7MLWNndgHHplkxnhU1UEsxJTOqUi
MZEAU4wNVKT1LWh6bl1AXoA7Cm7I6lWMR2zBPm5mgeJ8jhACw03dTKg+4YRHiEDm/xFetpGzJe1S
peyALDxIRobgv/YK8zW8OdtU58ZbYYhqbOt4iFU99WXfjkLMFnNjfqrkWmBWgxX5ctxvOEYH96ok
+8WLlqutaGhczmdDs30Tcgs11c6xtYWJJX+sHt3nnDX667cuT++esNdHdW/qvikpkdiixfSMJ45X
6+I+UQlmv+2ZAa0beyBZIeOEvq9x/IbPABLcRnlnd7cScHWuAYEUos/ICYoIQ6rri4KuPg5xnrfO
lwozEL9xW4I417ig5yRdr/aNC0iZp9c7ZjDEy5QNIbgr8k4WvJpg+GRmlbxiHCmUTNtprJEfGUWH
bLouJVcgaXrPI7R/Eii6xsJyS5IKbBlP6JUCL7N8nhyTZcVpmJ6sPF428/9tFXNm5UknbztFqzTL
fGxAr7R00gv3WQwlJ6R2fDwtW3boD03mzr3r8LDAzi10EbHC2/ljWCZe1Cpu0lvtG2SJudl1+FjS
YQ8Qt9ngXsS3QJrDPibkU3P3Au0k4W89+znNZy3DTYHIjC6X1zZDNlg2Z5ijrdW4fIprPUxd4xCg
Qvgm/jvGulpJoF9lihiXoS9lpw4h1IYKJjCNHQMNF2LcIgStLfSA1mFBOsE71zJV4fp1oj2Til/g
LeI0/UNZgs2bi1vcHLaBQOQrrAZzRSIU3yLMISrOSBvi/H4RgJ43wGWcUUAqv0UvOs06u8D7D3Dt
YtdXFd5x+1qTZ/LhS65faeTEsux+f3lSdtBUfwIaxhp4eIcuRWSOK1w/6tO0nF+aJupwAVbn/2Bl
DGcAQ8NCGmHuRnlw26PIGTxTHMe1bXHTIA2qGMCcxv6OOpHwOQo2yCdIlvmyg9F9hJ77GmfBpLmi
qlyja8U33EaMLQTYa42IUh6HI8SXeestAfWpipshIQkgwS+s4URWtw5W1XtDKaXQe2Teru2vZr2y
mOUr67HEgTA3Q5Nt/dBOrnC5dU5TNu3SBBYKfV0sMEttIMdi4MG/dAd3YyKN5ckKxg04Nxnk1BC7
7STYofxDS2tMlHxzUXMp88AeH+Qa5N2lWdd25CXL005ikJh+i9Gx7zDL6dJslFLQQDSHiTGBc33u
TYssw4enajq6iZqD8Gkckyrrm0v1N5wQAB1FIeOj36sq6Cp/rW0cWadY5dn0AT5ZQTCFmob1povL
MdLtubgNpvr+82WyQivaWKmhzza/COEzTC52EfeR2Xa9DDPCa+DyHFqNrXX8edbILBJBFLtVWr4u
gyBePeiGsCZ0iyyDZELgYk47MCpafAGQy1t+P1wDtDknKoBU//gQGgY10Lix/yLL77hnojphzqK7
3eT7NHavs3hmGwOmP1/9DFkMchPfBLNZP85ANHUDqsGSqoVul9Uh1795jjpS8+mHI97jt4qQikTL
UqCRkZpJd80A60MXQZ6KNAgB7Y9VAA0KaqSiksbQJTveOcwTe/qLI3bwy2JsvMq91D3lC0ejWsmE
4ab4hNl+oK1V7jlJsz9KkptjE5VxXzkIJdqoloUe8eVGHby4kmAv9bIAEjq9SL4VhDe82Dyv7Lgz
/6dWAJHv2WZEdod9a0vAGa3kWJfPcGcrW1ZBf4ptq8KX57qwlw9zWFDZHPWNS7bqjU9M4inqoSBp
kBgD3+FHlc2F5YxZ8nzDUwtuZAxwG9hSxT2ElP58l4cb3QXdz/7ZiTGPW/VILZjoKsBlFALpeqIR
s4cFyLY96hT6PmVryiGuhqCnVDTR3JJvL/jYxyi0MOsYB1lBZESe4JSkuuamCrJLMyaPcQolqXkM
xWD1Yq4KsB+oAilZ4U29Pqq4yiIyltA051hc8Y2k5TD+kt24u3RxZ9Ky9OEb2EYcxBU2MsE/K9/o
1X1kXfL/0w+IBW6h/966nGIsPlWx2MTau+2WcpQ9/BWmBSIDyGm6eQdDZAknoPedXxCYJ8O5atoJ
ped/DXVz0cAgf5DnSy4kHWCyjSj6vzQPGJehExKTwd0GwbyOG3d0MCW3va2rWFcknKO4h/4DN/Ie
v2Wp3Sx6OHNCckv9dJ2qyjKIiFpnrdphaAE+zzzboF16kV67fR7cx1M8mSM5o868FVhr86uU2Xyt
03AB3J9/s1N3f0+oU24uL+qhlLbgYOTyUoZwKHABgLwMZnBOCvvQ0K0+2qYVlzPtN3fAJEmgIRv0
BPa8nl1JYQX6nush0jiL4eOvAD4ZlTm89ym9ylJiC9X9Ngsg3redVaSVbibRfi6V59uafpLm8NDT
ZK9YzUUmiLqVHMF1CfZVnBK4IpfQB5bbUZgp5mPwdcjlgko53WyVSpHpdittLslg9zeaxGe7AluV
Vc6EdP49mBpnq2xv+Zkv7H6Sy7TOLWhWYZ+hlLimrKXFQcOj+R1w4d358UkyBIYawCPUiDowPLfa
RXMOdgwVwG0RITthYC5JY+yViqEjUb2Z7eVfpbeMQgHxoshOoZK4xcKB+vnMdwO1od5LdxgubUt4
bZNK12s1mXn1XyVVOp+eTNs4R9XEyGw6y1ySYz8uC1A+saZ2l6GzljXEtKSqZ3e+S0Gbpx27Vse1
1kSZuZ84JWT473bbzHRmy3wOPpi1oZPfhWiQRTvPrstuxLr2TwTese3s85CwdBy9vzL+6pEPbPA4
C2si719258pIEX47G/c9OW3Dx8f6U80y7FNVmBO34/J7lra7YwJyXstVfheWvdgF8E507HAxNCzD
AFqTCeV8xpzhePDMSGkWMvNf7GDT+ld4kZP+XlzFtmTAW+O20OW5uTeipMWMIg04rDFhqSFMsq7X
RBUYUpzAL7YKZ7rlayDZqa5+JlDypkpvJPewYTfM3VdyYHkNAta8kp/NPEV7NLTJ/yU7kGf6FFLj
ioDvxAnN7+Nvb8y8I/tEHBZcco7N+U+vCsyPf7BTreRrCQDQ6t1dJzEa0aFhe6IyA8quOFGcqerR
Z4o9vbt5gBhFyGGMORnqfQ2ebjZ3ZW+Y1irRa8IOG/bbHFgBkkvFYyI0og947KbWBdnB1VxOM+on
CDEYd6XwDAg7Yrfk9XuJWG5rpn5xWoxmC0p4fQ8JwnN5W34SvZrQqYELeQNXQ88fb4bThvynIklU
NpTZm+UDVjYojVmdZ74bhcAQ4+vwDOWEogkQJSt7VdUBWfV1lZIEgsLeGF2rb0c9+eiQYURA+NUH
+er1nN+Pbalylh+PIXf7TDMxGEiTWG15bA3qsFATU6vO4QmyXAbgO5XDiWBIcSEKl8BSqrsnEEdI
6VR9VMC9RIidAHIr3aV6fpjRdl1chdIljEVze/xEDEyD3YJgryeDRXLrsQJFAlVoCthhOstQbkWN
1+U+Ux99MyFYpRzNvKdpKQYv8IQyNYECgt4tFhyD9L5pPJ2QcPC0Ca/glhxRbWmk0G4hp3QxJUUF
iwhC4fLILXm3P8SU8rSg/nELOG/Rie1p5Zkn9x2toB56FJu/uQ/nA6C6t4GfQHhxKKWqXABtIi13
Gc16J/HoubdlmzyRgmlXxBKBMm5KrsbFC5KD78r2fumc1uLIj+AGmnvh8Z7qxbPzmTWUXoTtZ+n6
E76w/is03DK2tRoFQ1Ail6e9gCkX9j8J+CsjuhDE2xE5fJs2qhIdzWzJ77x6qr6q1WPdgMfy3y7T
Faft46qaUXiAgFxnkOiZarxNG63JHlii9g4o+WUPbSjMzrqspLnM/f44eAT1KeNx4bd2QXEmp2rO
qrRqm4ZW0BWgDEzDq/DX4rr646o9Yl/nmwxTDDXmViUszaaO+TTmskOnImsfaFlRr8ROSmYyZ6xK
joVxODIH2/s3sDeUjzsx/sO9aNocwrbKynsOqtHxSJ2Kueisx8vXdRajFyod5YUxLQCf5lr4k9of
oz4X8O8rygda+D8qewwd9FD4HVP4BE6VjEpSLWsLNEVHO01RhBeLt1LlJnI3oYsW5XPJLk4dSAhC
2XbG+uvMcKAem4C/sv1JOJ9ooUNNRdv6lHCHwcWMytKv6yrfEOSi2Ym84aBE6SbtJyasEAmLlf7b
oBXxROo54DrKKe1P3U0/4S8ZgxKpGFpmQ0RPVC4yZcpbBOUW9ihwXDYnpDfd88CpcyZ4fs6OuOte
uI7FNDSDN+U9vS0opQHaupMg8Ab/lkDmPXjlD7KpgRNFj/XmAnQZtqmwj7GkzU/KzaZaWfflbBS4
kpmq9ntcCe53tqOQ9JsnWwCK3Uu9Wxd4wd8azMfoi4TJQstON6pp8X1DI9HINEYZY4VgTMvyjY1v
H9G2dVOOt57vHSYZjmHXmDXurnZ5gjOb3XygZIKQS4TftZgS81QoryhppHMgSNmjo8FivgTbCt8i
+9ODMmTGOG7c2otmiR6HcD3e7bVz+RgJmJ69aKdckDCJE3Vrd+LCBaymNU5RF5ACoGp2UTmPca2p
UYbtm3tho94I71RvdYb3c65R/IvGHHDPwV8NBHxoBP9O/iCIusXK1sMuPDeHbcTqlGFEWIvSS2HU
z4FMYljyNW9ZOx5+lb9Ah6Qpz4zUNL7XxqM8IqkaFb5ILdaCl0QJa+mL4t8UQGaf2miBGNaSxiHV
/vnsCcBC9gcAV6CQ63xSmfRgOpL74vMeUb5jPT0hHVA4tBw4nihd3GDsudZH0u7Y2QnRPiymlVQq
gfW+CYyOlv/2xgbdf3DAGVuPrZcNnUiMVbAmHiUHBsBFX7YiFe0kNnUPi0ZHKdd5woKMFfKfADVO
Pet8fKG7j+zfSfFV8zIvk2RR8dKlLAtrDLNw6ztD+pkjaRQj+KCXOFkwdl1Fbm6cIhaQxRzbSq+r
4RbWSizxn72MIE16i8fDhWdqeuiMo2KuXdsVMClu0vPeCJCgoIM3u2t3ACWDmS+PSd61g97Ywktu
SQi1VFOTSVNZeeNp1DM//KkgAJrqig142GiUuL/WqptUeDLOOXG9W0M/P4eNYat6p8x6ap9kHXDb
aZ9EV/naZKyVQARORrcQBVZtmGXNfy4DJEWItxPjZ4I1MgEsv0y6p4pAVbNyFWovCadcdxC46/x+
HsuLgfBpTnnhJ4HR25HnjYBBl3ksLG07fqWzhXj6nddF3qPCzCSar4355NCOI3LikDfV+nCWGSgV
mjhlpfrybnob/ZXdSCDzg0oSgKp6w0hklB1VB5hVxI51q/VFqLW7ZOuEVCe+gidVENLKHIggnAhn
dsWgBbLz4NebdzVDY83wM22/aSnqvrJeHQM/7Sm1y7Lf/DmaoZj7uZpSoE13lOiEAhafuYUFPk+Y
DGh4vaJ19RMqqhCfasDN32gwFUtQXPl02jM93ETpkXKkAFZMKZIbJzcEaBZKGVqPPtIeF/lSsdck
wIGJWyYW3VxLUGY6ehocjwjGKB3h7gdbuyis58i/G3iMdyNdIdw/N5w4hEgWe/LsGe7fkEV+f6ip
ddf9J3kuM4ESjAzd0lJrNomqksz9zJL6MrVRwy8A+xGC8Fb4XdQZPhCtUuKQLshy3cFPqGlwCO0i
rGzR02hVKjyJuVHmik7zHn3VKOcyzlcEuihpqEnFD6GR21r0Ku63xJ46yQwvsGmLTer55GVlU1oP
s8t7q7xFvV1dAlac/W0v4UT0TPjOeebN5ygucF2c3H9Ith1bnzlKGDIJrlJDYKdyauuzCC5SeO5a
N4N5JhuhMiT8/3nxSv9wkowTN1Gs5GUonTq3NU+LD+JVWEGAfy5/IzQvlezRExl3e5vTfIo9Rk60
bMjI9NX3EFpfCjsItQLBVKTRv/9gipfZRcnoHLAwH5fBle7UlNLDGbaeOnRAuxrof6VEdxeQcThI
Gu++Gqjaexntuq6Kbzy1BeBJ/6X6/WgEgpQkgEXR/4k6XmVQIABemJ7txqMkiq0hAeW624sewVyP
odFPAmRbvDEgxct5IgUcLjk+OAS150+XxsCk0JBP5tFJifpBuU48y2ZeqEFPaMVDiGDFTxHVkJ4+
leEwdLB6Juhf/5ZURMqQSpynZ6G9IJhdaKxadIjaKsxfSsvFk2SukHbdiOEdXWQG/c1A/G6B0O8y
uqqH+DWcqkPzybUEkhKp50aF/w0koRtAiOrEtRbUZFD2Nu1qxVWCbT4M9z84+YFxp1Iws9Vd63yA
p6B+crV7WfY5RNKqdM8rwbNnCOjd2wUH+qKhPeOFOdo2qsZUNjizoKCnrPs9jGiznFwR6kPpAIhj
YSvOR0Ds8j4aRKZVV12srCbYJQzsYrov3UQ+Bm+5xOA+nC0jZ231L5K8Q5k4yWFUrp0PMPhzwpSk
5mn674ecmXw4jc0TDVj0e6y1o1Uz3+d9FgVFWuQjLWQnqKpw8PZPJBeRf+58hqMaHV9GSQSuDeL9
G0uGMuUeWGYd7hCrVSHKTheHtB6BeO9qYBT1GoJdp9hDrp6ciy0tzA8n+NYDxhiCaG1f7Kwpql1B
rlD8W19o6TeOTvRjUvDwjzi6ez/FcMwxBlY10TdIjhsKcDP5ue9DXEUP0p0+UxV1pELyCcmt4khO
qnFt1V2X+DCZbCFrHPwEP63gH5nsElLdTL0cv1MRPpcfrhTTXznKIa7ayhBez1xUbw9tTOH2HOox
2PS7UToijN97hKYvSzap0Zm3d2g3koWBtPeobX3uO5kmVAgGkytPjYvzr890B+t9pkKcOOaVTnx6
8tpxUzp/AsNLdbwgPhQzrdsnDvknceRNP3eQmMjrEiKG4OuxBUDhVTOoRltlNRhRHO51ewniAtVB
DYQ9Wur3vLy3M9xqC/8mlPfqv0a9krlph6J5t6/mqGK2tPrHaNj/2qsT5p0Zf12WT0Qfadjwb7Hg
r+UVteHZE7GmCq5uPnAzgpotySEOrFoiVEBV8PUYo5163D1g125JDG+wuaLHVjNwSVQGYvbGMuGT
uYJ9ON61Ul0ysb+mU0dQC67omm0wNtTdghYdOvPaAs0g/L/D2ahaqO3chnNmgc7VkSEOLWS4fcMI
p0uu/OnR+5u8H/dY9Y/Fwrfp0Nt9bVM+RSy1obL/CmItY6iFJdgu8KC5qTPcRPoVv+2kPgGZVfWq
XraIQcDOF4NsEmLbkPZiCWQLQBWWxm9fwmB7tlqUnYmVJ95MQbKc14wzaPsggk/Gp2UGjNXVR4LO
GV/79AJMDJaqNU1Z/MBZu2b01GFd7284s5FUnEhI5S2tNldHMmeTtT1Q3Qvo47O+2CBiMF53YQF8
kmMiDFVV6naKfpuLHcLtBUBoolNfLIYDijfiii2rNULTkDvRmAVoZPdtgjZSrkdzmKv7pcRnzEXG
HxmhrtH07d3xqgqxFwtxvRFt76lfSBOyMQPRAv6r+lJkL0h9G03VHd5Ja9Tbf3BwfmUjwaoc7xD4
hXfPfBm3042XM3oMzvVpy4pXQ5cE+PznbvwWzYwBLJ1NFsHjHuQN1ShnVQ1EKLdyodbQbMi6fVLD
l7yiRSJ4dwgqZ36q34TQZxpWhRLB7r2Uy9Qj5/ePb8PZJglhS88ICFhUW43gVneIwe0EawR0arzI
9mhE3+sG9qVubiU8vCKDZkpJWifrqZwOgw5UBZRRiQYVRkTygkMTtxvViVRbly/6HxHzdfmDUMIk
1zw+d8qISWN/wsDYd0VvKNYlM2K3T6ZGFDdvZzU3ehxmN41bxKbul3yMHpkrtBiM0ZQLnTj02XBT
Y7uZw0MccS+yNxEaplnyOvYQhIzhHvd4z7e2M/zVRMfnzcPdUMqjJR8FHZh96rbDfW/kO/zh4o8t
v8RLEduFfbJAQB5HFEn+by/GkTWbuiC5ROXFAvyDMJlXAoj+wq54ZNoUsDPFONl+le+WcHgluu/L
o53cVHvnlO0PgfwBm+FWI88TkBp7qg82srC/JbM3cQMXZD/xak77r5qXoJ2zyxp+FHE0GoFhP5wV
tcs9ShFoiGgeO/7JVUOUIszoOmZC2XD9vcW17A7eE4xllXEsX+fHvonso2AQ1MB7h1MDDw00qrOf
DVWkpfGh3nEr4PdxIqlU+vn47nF6NjHROxsvb2OWvk3PLA2kt2ffLQgepzkIEsf6a/VBKyArInY8
W7j468+D5HjzaCwTbBPauuk8ukvzxudwtRQMX5CotrcAR251SYyY7Pl3v+hDBOT4YVFg1Bm4ChxO
4CKvPW5vDKl9Uww9+T3SwoorYvaf1QpN+ZyoAxQAJ5S+N4vq0LY4mq3PM9EdH/ib3DXa4o8jfy64
gBJe9NYZmVUzCRBjD+cDZlM8bNfNE4/OSHmXix6Y6IrwXvYvaeZVI8vFumK519S7kPJ/eRdYADfX
DHkIf4JMF58INi8gInpDSnuzEOcDFJ9YLx8/nH9FnerIrRBfCLpWujYiDTOdKOusCG69p3W8iulr
VfwTGXznZMAQHqGq6c8GRGGLC41095tw45Z10SfYfpwrCWvkvc8TfUCyle0tNA5XQANV9/Hclqpw
BaQgWJQUGbn1CMakAibsvBaoPGmfWqoiywLiaW1M8WNwboSMbCxR/xw+EF8HRhdCM9sbU3fBQ4Au
pvshFmXNIKF/oDdZYg+p1xRGinLybqjR3EsRcGc+wposJHTgp5beP+MZSNxzsICEc6j/HfWgLirW
DNwUN9ntTvaUq1rnHkTJ3y+X2WOZVQuoteerOJR5SAOGSLMRV98fslErEwE6hxI58p7bkmwkYW5N
pc5IcrSAHee7XSEYQnUplDsz6CQiW2IlQ3rOrNQsyvPmzjMhDXaVFDKDuiEsVbcWLSBXJjNTyAde
UnuYAnqYuUT462xPdkxb9SqlcWtMp8Se994Jk/G7+SQ7SRrNMTuO3xuRT0LbyqDnzEAEMYRCDNfC
i6ldDwHi+jErh6WoUBmR5G8jV4bIqalpbLiPM0xkz5TMpPYf6ncx5cOYtO0olvEpVQAdbPduvLx3
amxBWWgVjzmgjN5ub2JvlJrnrQeICZWwBKJ/5b9zVkSImXAKq+YR2UV1mIYaADDnrqNCQXKUYjHM
AC/nQDwAzDvEc3N/9ZSgSNZ8nYuU9rNqnlwv03uqT8+sA9UbQ9DS8OYm9DxAjhzQK+V7JOwfEkgk
5dSHqgqNl11MoRgo/QLqBabrHk8jndZPp74oIf82b1gGaRVYLlBV0qTVqhua2U2hDuocQyQcE7uI
FbDUxej/R8zO6NiuCtSTM7iGw+Vtr5zDPW6SL8DKyKZRsy11hE5wWJxGO8Z5cxcaFf6jeGbKCA97
sK1G9nJq5SkYs5cQPCG/BQ+XmGY+qFx2icG0nEiUAxFjGqN7dOGRf93Rr+vTxfemiViU7bUxEXfV
Q0sCs95IQ9M67Oqzkp8QkfCdqra3lfYtgd4I4gcu/0HD/8YsaRXUy64KVCHsziuf1SVjFrfu0R7y
U8Zhs3xR0+aoAmbaHGQXLwANfkQb5pa01iGQBtx3L1l9/WYurr+ENGJ8lcOqMSYWyg5pwQM1Bymj
+XC545pKH1SH/b8fjRdO6qY05EmxH6rzVr7IFGRUkVcaB4Cy46AdL6wydacKrzPOY9NEcaHJsmhp
hBDwBa3LF6xbh/bhZAEVMckHP3FVdxafi/wiinHrYd3qyghFfM+Rn0luDIpP0+YpYL39uaGv7IGu
8a9/MCm7oFLAmZBXVUcfkkBnXuJfEKLR4TFg5azLaiZJlZ0tDCmbZvpTOnxzdHAFw8i4550bmZFV
024L59ZmaKoifJREDvBXgPh8y9Bb95tCEXtSwXmiAkUveRHqW9JsB2TaPdYViwdN2vnGJD3A0qZ8
ISdG1jdI5ioMYdM14ZPRQSUd/7eAmEnZfgcQXX4mbCixpLD7llE0eaabvN0v5pChNHVL7EfIiefs
1fWQ+anXxInjFG13qrLk/GqdszBKj3oHN+ML9IL3CfJX96OVU4IY6ObdWie9YmQIiAeNpI8aAF8V
l2IphyJkRococCI00Q4BPjNfnPUx78dmmfRS43wpdTIcelxwOMsqnPDKXBDY0wi8x8AxIfYcUCHz
k728eaMAU9YLngRy8FTpvt+cgEjA96VSjnpt4sDYwXHbn1K6EczkqWsCcLGGm8vsH8BKuvzSEtjS
F+pOHNTTmGbSrg5LfOJcgrkD4JiC69d9xs0pZMkP70y+CH5UnlwEbchOdDMixAEr1vQjggQFt5rS
gSdm+eD0S2yUSgCgT5ujW3FzNoJ+lR/oJAYw/pNoS2aeFn/H5ZxiE8gqHaheyHjE22EpYnt6IdKd
FDRcrUa53tY5AfiMBPbMGG3u6oKPvm1i0fgTdt42L5LQ+/UMhH3u/BF9ksoSFh4pUt6rNwsgadmx
pKcnsKx6Pm3F1JdV5QCSa+UVy97sV0wsixkVaAtGMP+/tFwbQfQ9FH8Fv07EyGRjPB9C4KGPT5nL
unSmlBwAJPYcTFV5BGpV8MdrCxS631jeHlW08+XvTdCJ377LrgAhIRHOxq8wpiBpOaNaHOCBEkVh
M6VbNNG7TYCD9DQ3ukBJfNw3JdybMO71cc72oa6fkRuFSHsxYWgANy1bkpaOqpy4f6XLsmKEeMq0
Wx33JtSrFpRCyuDWMC2hbiaX6/dil6lp6v2qv1FLmr+lv3o/lLsJA074dmAsvPHdWrZPzaNuIevp
wA8z9jWkxmdt5nAez7Fmn+jvfcRjszM5iRdQxCYFIb/HXYFVGT8vejSR4dghHKySmpnGmJ+M9zvY
O89imMz/MAaDtudKPDkP8yBC7FCBhpq/fwqL4d2NoUTslll35Ow7wsnhIIZ5hCL9eaRC5S8XkfWr
kzMd6CtZrESk+eQntCTfCqmBqCh6A8w7g6BkllqM2ZHKnmAJgVAf7tIXgP9lBlBeCNr6czZKzy7X
o17DzCj8urj23iVFfBGZOZ51CaPdZyqIE0hh+e+8x43EpZi+mkhsWkHXXn64BWGPPAY42ry2GNf9
JZhhxkJuV/DoLFaZSdY4s7Bqf2VOQl5eTp+xpGPNe6HhmF7KjD4Cwl/svKaa7HbQ4DZb6V7GXQTQ
NTl/FSrYQZAWzrOmbg+QYnYfYLHngijASaMP15bFQKwFQ/8brW4OhtLbgCH+Ibu+ljU+JfJ6YmU4
hAqOTQY0dWMH+5dIjd4hEBwrQGL00FVDeGdWiI8NaMyVdwUQAHfDdVpmS5c6H6HJExmlZXUHFXMI
p6f23URMhEv0bfd2J/AOXQg9ZmBT2LQyW1rAElO0vHb9FEsMSOwkIyaidRIZcDypkhMGyVc20OH+
EX/byexhNR3h+/SlnCs494UhSNvw7EHowE/rUWui9nN/jJ0NZpH2IXv9lVvp9EDYg4TXUpmUdEQF
OEkASf/SVkrD1t/scGgKIcV4pN/m7s99mYwBWAC6sb+Sfw+ZAWJjsyZd0blxd0KGdGVPb1MWrTMj
KnQW9OELxyENOQ2ho2kifP50eGnJEVg3I0o1q5O5WIRte6d7xIPCSCy3zCPznYVl8WRrY54D43cL
BkArOnquDS7dSm8A7Lk2ccZfBBdPYVgLLT4GP6PvVC6qKFdPTRS6EFDbkpBJTcOy1CGZcbYxnscM
MqeJ6zSRbpqSfHHzBGXC7BRuOXwn5MZc+Aw31aBHi81IpnUl5UwxWEVsFBzl/qTgssWHESOIKQxZ
f/qrs6EALNK2HZxC6/lZcRLSj99nKiWsFtv5mlEJPchfd1CTGWHEm5Mlo1KE75BehkPlMpf0q+yM
GO7BjFbNyivjJixYrk1JVQj4qX31QDTNm3beQ/NcQwXqjBRMEOYICUhTE2AUKt4WxKmbpnWLRJ/x
I62o23oAV8zRGvCblgNGV+p6AMphWZzLTQljITZRlnaShklfStWNXYYTGyxNLQiyoRT6InGKcYRr
KmWegDq0MfOQlZWXTl1LPp8jnk1ApZtfP9yT/q4qAt/jJBjt+JcHHiBd8vH9+G+mcQupiaFTtZVK
UR/2b0QRNgXr2hhR1ts+ubO2Z+yWLNyjj5d7FTNOaFJMl9gKxPb8piUuY3QUWG7ekmidlLOFmD+I
8x/XQ2i2DweOYbR1jlQdU09Etoi/XFuSSnB2UeNah9Wvlfg6uYYLR2WBsazVtdlRz2SL4gCQxrS/
9H3q4PmhGMFUsRdIeYS6xn3GjxWqt+lQ/A23BVA6uW9q62QzX0G4X6Vd9lcNEQ9hnFnSqiKoca/O
YdFxl4fePbkoJ4XiP5bY47LrznzbxtIaCDQmWVt7EJ9hppC3Wc1+G63cJgu7Kvne9YN+3kLp2aFf
AjCvqNAtURqvfC33kfERX9nW3oDD9bqiMAoHCNRS7Xfo1rtrmkLbHXsLmwPysTiZ4oK/rOIh28ln
6zsn4VBdp6Uk6x9TJNMN5JqdLpLx10UXFGqUSQterE2++oBJ+L4ccvU1d9JnsmmE+/rWNVvYxIzx
E8sCAA92qNOxMJ4eFnGTRm9k4cWv6Gyhp8d2923aKfhM+UVEA4Aj0QFr8BBBzv31hbQ13xHt9G+Q
g0fSkIgymJCm2xMrMlgBNZxBidCjnWK1Y51QMzCCf0DndvCYF4zApcI/vjqrG0OaaIjxN4zTIxRj
iE6lFpSCV05QjKXkH4CSH1z+qx2X5q6GU2LcMlk/T+YeMeqBvFDlZlLW36Od89jtguZUWrHlNnh0
THv87PGpLZ9ntRCHIHMSdNSUV2cpbkkVcAoyLxDguZgapQfH4USRAFIIFaE403cWJaRWv9ny+KYw
jkpHhnuJG6wm57zJpzqiwhdqZAm09D9U23O1biT7dctC1kTITXBqV+YrD7TYxTXVk8QN2yMUpWtB
T2UmL3OMTc4XiIMTm765QO51lD9+8TG0qSSPdN7UzZ8iDeWsKX/Ja53w3SqxntB9Skh7nuxYrr+d
uTVIK68y+haBy+Tqvj/d6kQCWZr8KWYv4LTb4mtksh+FimjkAtGr1RmgeYdmIcV8nSc6W3HSCSGa
Rrc6RCFAGYuAvq0q35/F7okKmdarli6CcJAhqI1M+AwjZGjeDxnSiEvmUmX4DF4qe/o8K8qXFnU2
0FigBOUZCbSab9uoREhmQrsHt94lNCGx0VH9EvNY410qXwO1dr4qwYggNs94NgAmjQSpH9NqByj1
NDtO6f48l/Cn+om8xTJkk1GxreihWxPd5cnmbduHX53TK7itDq0jyA1NmrvMxNF7+K1DrGOfrSAB
V0l9jXAGyToy9cBzGWBWUHjK6w9l9cHyHK+E9m3oSVAY0dqph0wLiRcWKu+Ijkm2qxOd/EairrZn
FKmYth1Gd9UhFka8ltBb1RQq/bLPUMLzZr7mFz3WJnQOrRPPV21+YwkcOOE5qDZxR5O0fHuJuTHo
0urq2MKbEjqpK9oUe5wTk43ACgGHu/koNkUj5pGbK5ugdWsW5TnMR3GQOj5F+2oJxMrayYj1wPXk
a0V3I7SON66OArxLhwtEuNNEO1gj0mw5xAElGUi3mcAfxLEwF5XreD+/k29qxnDBxsZkfVXE4krI
LheB977aiNa0LPeWeDVmGBj2ZRmNRDngxzLbbekCGJiC8ZPf4X4x1n3sMZV6iQ6M5FSIe93/oMBB
89Hy/f5dO0yNzVji2hzYZFvLFm4HguBsYuIlFUxvODKoh850yf6bH79V9UwvFRaIpmYTiOBuA4Ye
v0lZcNDfodQYykf95PYD/U23bttD6HVosNVTwumCD+Ub/ffJnrTzVhdBo9VKF9ILAQva7DudPlTB
EzqX9sb32icnvYF7Eio0GGU25QSvIT7zfe40/ySjaGIAfh/XGCGDLHNV3rOR6XDgmn4ty7vTpBGZ
5eiMKwMA+eV/JrD4WcLo/pnKjpd/l8NcnuSBnqi6mjX2a9xAd/R9+3KswNEVfMhihRGUsCVVWI+P
8qsDP5Y+IMo7PY3azQxBs8lr1I/BbUYzGnLX7lHotQ4IZx+O9wNuDvAbRe4gt9HIgS4pa7mV84X1
3XjM6zgQLMyEzYBY7gRKin6bAAahuCMJGkKQ0ZXlyT4lMrmJztszh93dAsyG04J5N8rI5mG35RHw
UlTgHnqo66IoB9mRBQoI4PcjAfnoWqbQqJEelMR4Jw50cqAe4MFZbZYTizvv3O9rj/w6MIZUEsrN
ZqpDh7GLQ1lMpyKzav87T/tuTVd0U+BftRIWPF3gRd0nk6vrPu0zt1u4N5YNb76mIT8liRqKOOf5
cd6EbHZbYhcp5zVNR5XU6GTQjlHuLWOceIgiaEZvTRQrBccpMaifKwgehpCQ6BWHVNl0QUqlGT/J
eRodTS7fAD2SvChVZZBoml31L7QEAZh/ie9w1MKjb8MIkcjuGVglCZPgPVMQXsTenMHT75gNyvFG
g2wMo5QZe3biG2WAO5PsKwH4WUeagiqmmLJnyulYj5U2liYYrgOzwnIx928uBTIf++TYe/L7a22f
Ozbq/gA8gahMLkVpd/PqZAtfU1fyv10asgTgDLYDKKcTlZamziFmSFs5femB3daMSVxBu/BADtSt
enVDuNrOafS8QgeaI2J21RTm8MW9Jbusj8XohtzC9jXyh6VHiUzezmx8rxFlBEMbotZkbRi8RQ7h
47jDQE39cwEZHt9omp4aUACL5sgHUS1RcUTtcnijk/Oo9PKIChEMSg5V1liC1Mu0qedkKyPJKIY8
Z+X50TarPESX8JkdX/vV//Q9xWt2pFKDbcC/cG3eWj/T80T9ADMDYJGNHcGYWyLRs3GCOD8LZycj
ikXpVXU8Leva2ZOjxlI4+4QRZ/frfWsCBKFnr13ruOOfRH7Z+fhAn9pMVjcr/IOfHpsUpV0i5ISe
p+4JDUi1Szcb4SkgHUKEDbPW8o298biIOTcBBucjypcknnl+CbUk1mAG9Hl+3dSLZpOlducpcmuW
yBBfFQN4lqu180E0P6Nrz3xUF4N/Q7eE3jrrhU+yV4Vc/kZE7eubmmS6MaiuCRvN1DWJOhwQyjW9
l2BltMTa4PXL0RjDloVZ9HTVF+55BqMHHYEm5j2Wju0bDSKJmSPxN4sACGutrvRlksZqh0elRWX9
yXeJx8mqCABwBlWB9viLp9hqUYU9WFMt9gXOl52u7zzidrMt1S5njJKBCK3Gr3t5hzUw//qH9+jC
0034s7QOPIxj0vpZsOX0QvxGhV8ZUtwOXICmE4IwYaB8lI7rHya/79PpuZljecv1SeYOkmZaw0NG
gKw2QHyxOzQcROmb/qd26a02hr8fndk9G2IA2fUPw8yHGZz3gTze8+9sCXgfcSgSaYaPKNkjmxfC
q2dQemTAUoKxBp8+wq3ctpwyc0+1VwpYBBRIP6jsBT/sUE0wum9MXh2Iqyx5cQukPeuKTAaxCbX6
5w3D2sYeavkNrkj9VQopP2zGnaA3RtRJXA6We3Rjt6xRSspAOT3HJqJtZmf7hZAbbQGNsW0xYmPt
Q0WY/SQTdMQQSvcnL3oQ0Kt1dFR59UF+oZcBHkTLoNhxd2O+FbXMaAQFDGoLmY608ZBtVlK+8gL6
pFiWoeZEFxPCmBuAv4KCUdmblAAtjNyPOeWFMPs2iOnQcmkYBRX2hynIaYDhZvtwcPKsAS8WjEGp
ve+gpZiY7rbFE3HQ5D3hKv7J2OZLkGKIXZwSG0o84TtZ8pBnSMVNbQYCWDLRY+yobMfcuJrq1rL5
88blu+FvYDIO++njH4NADqUHUSfk8U3ejrzfp/Wj4n47XMc0LRHZhA46AsduheKzVFDWID50qWq0
LzqpeOm7On3sWMGYcWuIYVEJCZxDGG084JfC3Al1v/qoQy+oqzxCp1CKw0fMpm1Y9Yxv75H67JCt
6GiYLlDD1WrCG6YK7c4lzCMfJoTUITs07ZSmZx2MiERNO0lq17tuHb/u+XWR8GlRLQ3Zels5LFBx
E3JZxbvTXrI1aqGkWhBi1/hmsbXkn510nDlZdS9fNCEqXNyiSXHqz2mWBGePKRa/cA+WqsTpi5AB
RgNghtx5bQ0f8/x1ZH2ZSIeSdKpbQe2F4cJ09oGgFvUEFjlBFA+REfY+XUvenqU1wPOt5t7IbHFw
/lJ5VbRmRP795yOLeExHBXIlcJzLLnpWWdUcoDGkoAlSic4usjo+lg07EgaexPhzG9dhnOM6KrGm
rxaICJ0AeJ/GHfNH2uvLJo61zPY+iya/4z3Nb6rypvhOCKlICrwEQP4dmYNEOQOIDk8PCzt/DWj+
BsL5yLQvpco1TekJRu8oBZN4nr4AaYrPFdyVvufFDX5dO6809iEHeQ4ZbYPrC/08fmOCIUJSQdMd
SOHgnnuWvO3rHfr8LgXS2WSurMm1OIpW0TSdh2x6fQv3e0YzDx/ePrfE/gIoApN8DuralJLx2iky
K4cS9RfjysAlj+DufEEOzOVlMzxv1zUyttELmNag2217CnNYDJdB/9FZJ5e71Daoaj/Bqkql6rVA
YJ/8ZajCYxtra10yOfviOL9RLxjID0aYLvMYyf1L+y16V81QTzO3/Gpdh2XNnCBTlPxRNQDYSJI0
kuqOPfwL2Cuh87gRPM+WIk5aW6GiplnLBQwCuOMQYEH/6YfRwkqcrxC5irZYy8/3cZpb2EMhMvVJ
fPLwQQ7KK5/qYXrLSnpMGmLuuV8+4i3dZEfpxTCnzm+M7gpminmY6di4wWGdui8GLzFtkuURVxHa
23MukDAEKWweBFtmtd39JtTDHpetS+Je2uU5RvQ2EQiIXAMkH5S3F7hT+mLeeZTBlLwbSxQZyyy+
STLcZJOblQjXYGFKFiMZ9aBIB6+7d7NjZRlKqWo3FhVoDGltWrVbszHLIWS+6CmSjWF16NYohom8
sAxHNQcdB04tmLKmrp0AtZDzIJfKL35Bt6CJZVlg/IGvN5DeVL7wfYmeAg0ZiSZiflrLvZuhJDHy
aBhuJBrcqHrYQZu/FBgHJfV48HQGjYgGtldowa3U0/tgHMmCOz6S0nnWIMb10ZSqgDmE/fqV5wZc
MG/n5u49n/IBWRFW40+rC2ZokrQZsqmue2L15VEemw/sWIaAP+b4hqSfXkboym52A/ITWiENLa7m
fruZq8s6T2WX6hMa715BKaj2J1otZHxvAjJWaq1FPzLnVqd2hUSguThBv/F9r1LnQwr1dvA02H3P
wVUkbXHe7qICcBCFPW4jUyov9hy2RxxYA8/hoeBg3MY2UeAqetL2s+4yons5MNeqp5EaDbLFt2w6
U2/IclMqhUnwjOXkEW2DNbAPptNAz37CnAOQ5EMLEQ1EK0y3YHo6s97HppvY+uzUhkL/Esal6uI1
6L0k8VJBOb1BpUlAPlE9OMtGTBMhmtjMhON25lI/i8go7c2qeGt7TNCoA1lMRc5Wdbs7UjzzaEUc
Mao55cMGvqlhwhxN7PrP+GjAne6pb1PR1uyRQXi+nPfMytP38tu56nYncu28avFDwqBg8eUBxOyU
YsoUdbtsNWqDF3BUxEgTyuJgvay7DmtRuwqZjKHp5ChJ4npL0s+YIilwQyF6+W42ky086gWdOP62
QLqV7alwHlVj5EkEJVcL2+Zo9p2CPaor2xahF5CBz3NAxqKbssDV1Ls5NqykyQ4iVTT8vYrPSQ8V
dnqcaPW5FasAHV6z6WqckRODf9eg3XJHa7hHH2qqyCXf3TfHmCa5qHszKj03LV5/Tpcz3iT3Abe/
r0GaBuY5kXnYypZvLvrC50kiu9X/kTdvspCjtQQyN+RuemvoLRmhrq6jswF7FduJrIccE+1WQRgk
qd0/NCyB3/Q145uzcJcaf2h8aAN9tIVr1UuFAUWYl3JX/lGFS2OTwKteIUm5jH/TUxu+QMTjZrCB
wqJSi7PdtZ9y1uLFdxjiEzAUx5Jd1Z7ZS2iQYA35wLQenfN7jZDZfTeBM7yw8n5mdXUf7i6KU7Tm
l4toXNpmwBflvwnDU8xYXD2ToYGgSy3mKQGL+n9luDoUGaO83BKcdjVZX21GXJ5hgwlojGYwmunW
xZdE7RetYJAvL6CmvZZG15l1znI8qd6CuytW07Kj2pBhbGwPWjSQIx6h3CqBgMw4tux1leS/T4go
hzPQLDZhhbHpjt8JlWrv8OqGFcuL2+otDc87WHTZdanyenov+6p6+663PKKlDDWu7NEUZxbnKd/L
G43MAoET89MY4D28OPOe5stO3vvuPqTW/wy+xTfi7oAw9MxAKIKmCO6u2UKf0mCWCja+d76V0wzA
7e+VJ8TKqGpOPF71FGNEccCxVHvK8jHuln2iXhbzNTIe7x7iWVS7uMDIZySlxh7jw65R/sQGqaUk
EqhJKz1r4bx5IJ0HPfNxuWUvWbVRNzY3xVX3+Ddj6s3TVdqNlwsV5mIHqsje6oqAzM3/ExlcLQq5
sFNmSae2Low7XAyXq+G0lJvtwMPkym1kbE50hOOvTPaSjP7yyo+FHy7d+LqfRDPBce4BJ7E05z2L
7s+oGOD2FzGMWes1Xbbd7wugUis2U5DfvUr4FNPbb9KAinWCeY4ak2FaZd5kVoKVo7nZiFutQi6S
ZsPso86fhG4DCuYTNfHBSLYSdbG4G8x4+sHIdQTRZglIP9e5Wu5elzunBqt5ums1huPQYTIZ5CLt
8mAPIbcWRSpY+YXyPZPB0zgjBtjkG11LP4AM+3TIyzoXNWerBiFpo8CI8Foybx0E+ZOZOecx8jur
oNBa2XnIusDxMdabuvFhDYE1nNmm85QTZV573LePDS2/zfsPZ8j0yvEZyI+GsmUtXEvRpfO6m+Lq
KtpoB310NAck6B2UXLOv9KNSZWbp4w9IsLSGigiyD8Rr7Rq7JnDioG0LOSTdnhZwhYoNaa3ow9rl
fQG44x3dF+/ybfeyPFOpVitkkrofwejx5AUWhQCCuTI3GPUpt6vehbCK6X5A3Pg2epVywt1CBki4
uCnU9DKIm6JWfbNGtFWSR0Q5HO8Tqn2NKL4ro/0GKHmd6rO/XYF+BJ7/wEcGIocZpALRk4EP6MhM
OQdBEVFPTNgLqL6byeYi/PY2tzpLUbpXBRnTmlr0Q9+nukAg1L4hotQI6yFWrqgIt0uu0oZl5Sdt
46JKXcC3prQfqoagJaN1w3eiWq2jeFTj2WZzuJqnaYCWt/oMNKDlWOZfuy2wEzk3otAT5HhfTQZy
SFbn2tDdPSiLtPm8a9VGP/bNBdnYb2C4G+c9/JbPp8EACcoKx5IswXqe+vviyuU579m9JrkFL8jj
OAerKXFEeWHc3AfzNHnFTkEQS6UB+eNGo41o1wYnWKa27mOkXY+2bSBrMZr5luBvApBP/xeknj1L
HCTiJv83ooCJgie8u2lH/LrtxfOaEFhrRG263KzO+Qbf5SxtPNWb2NzhtyizNJTnTe7vz6Vqy4rl
nIcrEGV9nchAgeA83FFVGn1+umEvv8JaxeCMQwbW/3TlL5/tFTP9hbGjzbwzyMQUSeyasrFaY9lj
Vl3RVWVgIAs0tq9G+OOaxAmlYaKxyStNKUeMt9msrHM0bfVuF0bTKL69FMrcoKo4dVxTWtCNwmFf
Hvkk6/QXExYc3g2/HpktQC1ld9eFgIJQ4AZld1SeUYinbOsdbwWM0JmlT2jf3RXU8Y/iHFNU+y8w
fmi5q6jxkXSYIUNlR3BGLFRaKPYA0wrdBr5v/kT+17GInLd3lFbi+IBUuTCrLm0tvodsqq06MZf7
4+Pkjk9E6wY2eBDvsWjlzTSzsdz4rR7eHSY/QXUJfRzsQnlB5qRllSvn5FtUmRlMBvZbSRvWsZ1E
zEsHV1y4nOG9ivwW7x88paOXQMPOy25N1//D7/alB7c1C7nY7Kvilt2MBowIuCeuMLckbx6by8gQ
wZq2T5c2UR8G3VkZv0Bm3PEpmsudpAUH0XD1cypEwJnaK+ZC03hw/JPktY3HceTuf0vU+dtPBkX2
sGahCClejychTHeicY7+4O/u3J5B2wAW0ab/zYqv7ZWGeBdj9MKBhE3Y+MXwTnSo3OJOFOXBsP4h
G/+Wl5C+Ac/1NfiPh5xvxO9fvQ5hw0kWaf+jcWJrY9zRA4ZxOGm3mhxsGUEzPi0CEGWLuB98vZ7k
rPH68nieF2pb5WklWecOWCAyLWTbszkh9Lsg/5asqJcJYCdn5ygKaJPdNB51mT4nINcC8vCuEvpP
X8sxlcbc+owKqDMdso+gAheaqcWYkQfc5jBlGbK0LoEEp+f2WMPiidTFMreeKQdMAJk6r9Blj+dW
yDqlalEFpLdkwtd4F/lntp4g0CVcPLh0OgIHaby8pwWW0txbiXrcgtLrHy/z1+Q56+2x66Y+TXYt
cjhwg0VKDWIXAPo9XXCuQxYmobTdEu5Ew24EHKeUK656TmlULnuF03UZ+P+m90dCysHUaEpylw44
zl9EM//oeNdYjnvpGvKRuF9p0qzi0jXqRE8D5lFk4OtOKBpFt1HRxLwRd4o/IPBWQFKSYHsFACHe
BqKr3f+UYC9uGnI1yu34Cylq8qIFe2yQ1KDxvOUB5KM+Y4o4Cx0fTeqPM9duP2lMoIGvdmIM4IL0
3cSzzle3QMEYzPb7LqSBjTxK3IMsrE3AnLVCMi25eDZBRwPePWO+vmQ20VJTAGBwYnjTpu50JhnR
Jj2/IjGVV15CT/WaQkuPcGvS4Q+u7cC+mTCQT5Yd2SN1hd5/QoprivrGODcDEUA81yc7Dr13c9PV
G1ePdqoOKX6x59BanVXjSDGZtTz/dExjjG53nPggCS0L7XDGvK/RebUhRw5mnIWBFtPy1SgSmmI+
DtbW8segNXIHuN7KTV44dPV2Ver0k99axbiYgC/Bs/khJ8yx4lWOQcpqWxFhlYg42kzrrhdRb2tW
hWURChvKSyKHoD9XsYk2EEmlYN8AzoBKbE18paEDQK8PwfNnsPp6nU5qoW0WJOfixHV5YH6AxtQf
aw5rrlrVEQLDSpB4/ScY95mk0/UscI+WhmAQFzOaCSinSSpA9bv10tosmH/p8IsKRn5MrY/+cSwk
0Zc/pysQ2KVD7bSa98gAQgTy0fsm4TkD177LO2bkb0uCUYHc3P2/1B9XUCVkdiU9novZkSS+x4lS
ck6v7BOO0K/cjn1GL80yIGgxn5745e2D5HZT2F4enOMZ/BtD3IiJ2+3H99asgb1Z2tPE+mM8X6eo
Ckv8f+u5XpY2RQ9qsXnj2HhKMpA7L4P/4zUpk7Eq8J/2vJ0SDaf8kvwp/KmlcVowMt4pd7KzGq3V
icMDUSl+kqleWssNvgbiGcFfv8+4Nc4laFO72y+UULGV57CDfDPdwL41pL/o+Y0oJxR1JX2EyXkF
qpxWiKv+wsAl87NsecItNKehhc+rP/UAfr8up/BCF8oyNaKciFnVDYcbEOs6TuGJLqzSgW7mhj4J
ODrdhk2AO3KGsLGlVpq98wp+BwBCnoBt6bRaz45iu5yntTk+qRHKlOkk4EoXeUtfS4Id9WOWVmY4
irl7CbztoQI450zNF0G5r1+2IffLQVgtrmaDZvjD5LmG9qDSjleQspkyDX6AYdsZ12enKygj2mNx
ggdAGDFEK5y7mouB2B5w6mvnqzRFPC+cgItuE/XpkpbAuoizD9+e8J11qGA3qY4ZkdgbX9tY1wHN
dI56qtMvul6MvKHBE5g9szqEJVbScXt+IfmlFeWCbwpnD/pYmIGHppGMbLHrSlgztXRYCExCVawQ
hqEp19LNb1ZwoBZqVoxeVpxXzsTwJ7wN5Av0rkUL/Gl1zp3ZtcJZIDk/B8zaq3/KyzO9bOBclHlw
H3i98YJOfZgRecsles6VSh1iFAfeupKPGK89HG+KV3u/k2n5rvpvZS1gB4Dq1sv2eck8WnLKlqWe
tw8yvDq52xceB2E0WFjGeStdRqCllldgKxMbCPN6l+4W3Eg/kU7RAXYtZpqX/gxsHQZ5+IKpUHXT
Txw24fAzAApUbuH/Kb1G3qrtDiq8A0iKjy74YohNSq9Ta2ghJyEDS8FpRHqHgYtd9eB5Xt0uoWrw
QmM79KBdKtyxtGt1cdQ54nVviZEcDbSHklKclMSiOsE2NoQ3O19VE8DekMvD/1NglieTnh5zY4sf
I7A969ewsMLxdsj0Vi82ojoB8vhIGraolvJfBA+FxjZr1QlxNMh1eijz0Cn6Zfi1sTYHbKSVymCG
1+p03rbGxUQVtv4djUpRvvj4POAn3dA4Cl3wTDg0yflxs8HI/JLeRD4OaCHH2NWGNeqNVWCRCaLP
WRJvBgmDvQWrtffGrzf8WerjSodxbswDCl9ex2Bpejz4EMlu84JXjzUUJbPtLW5evf6+aPtI01oa
wuwe2z211Eaorq2DjcyS27Ovl2AryD57avjD80mq3aXaHjeRbeL5hNcQO05n6nPpmiSERZV07xwW
FKnKVHlNJo4Mq39VntKKEU8ZG4hryhqaSkAv2XANHkoRp2Sd1Q9oxEoWTK0U6zJpBLztW6g4vGMJ
zFjiS0mhEDXyaWYT+jK3CMyEENPAjkQN91m1DNLb6ykQcttkRbpSdcIO2Hn8RsLLyjPi15IEUfZP
VV7CPFa5Uh3JXWn2/ZnCDARbAdkoPrW9YKnH0fMTU2iAZFMDvia4P5897vSj19S2fdW/XCGkjeT9
RgRL5+XF7n9pCIbbyrXxiGdDFBtLsoNG7quMxkAYA2iQ4lEcltw+foY8gfVpipc9V+hhcRbiEqfI
JFc3q29anfzKiVXl0D6FQDnhpeF08mU9s6buHUvJ5rjoiDWzPjTxMFt9c3MKmnE2Nfq0Qn15RALG
aVhYav3CDuJtwMHu0x/GbnGh1pBL7oy1+jt57GFn8uCZdMa3WmwIt0c8esizWKGXEbD1JlwxVjOy
JWM9A3fmusXyTNkVCgNBl8CBlBP4ZoSvBzCnQRnS66u5dsyDLs7bxABZq6/ovxuWP9PheRo4DkFe
NwPvOzU/DzmAT0iOXyssEqmWsb6hrajslwa1Q0NJN7KrwXyh4tJXi/Xi+EflaV3bRnk8j6ULrkBS
8ZV5UoBPGPYpsLF7MQU6+5AYSFQGYIOdLH57sdCDjLbdVKTU2gapKudenEsOoPIDaOAuZU9ira8W
JvjnKUc5vGeG7OUXuSIPjwqr3Iu4XJOASmpoRtU2dNo7sMB5qgvIpSc9cQ3GMCopoIvm7RmregHc
ql1A27Mf3p1SIGgVKCTvalKuXcugAB80KAmKP7nNZT57Q+ewYsz+82sOq+eDbQ7JhZaOn2M5Ekgh
ManVy0NDfOlWFARjUSlm903ACTgXe06re7BoQmj8JSozqIKbN6txdK0wj+Oim886QxyfxUWhlOIO
InajQbj+ws5+ps3Lq1EbAl2yvW7tZW5wCcEbIfMC6TpRKjlaBPh+dQRm6n4b9sAkTbtkkwlXuGru
CtfobRpMOw+B3MLwzPkt5uS/RlP8AtVC+KbMzsOhEOqAcXljqJQKfkGMGG7lzNuYEpZ/p+Fq6PPq
NG4eVI9ksuMPPAA6IOC27KQ94uwB0debsKsmwfV1k8SfJj7/1yEFpQ19Soh8FJvfT+1IvaBux8v7
6OGMtE1Bm/LbF4AP7S/JLfZjs6AarkG5wdnH9wMlUCgd9VboxShCCpU1k6G5vCrZiTLHq6sL1qa1
2MdPEa/yViqbC93Ez9CgI1BRLqjrUUJnIEmHVEIPIoWpNBNezrxaAyLGO4LvoDB+B1TAtVhvLVh6
e5Mwvq+2eLyLdLk77zq4n1JgcijhxVwXyTjoJu+QLCFATKMU9lTjMpD9IqQLEnOIk/NgE+U95TKb
q/5W42f58h/qfDNv91Du6BBAG9ezn7xSFeVZ1jV/1zXK6neR5aSmt5Lkz0r89TeyRvVQrMeohmNm
hzRK+njOnaLtSLJt/kUfpznjvU2nGBZp4TWmyQhyvC0thKzUr05WKkL26r/g/dDWS/kCgP2ELvKu
sQ3id9x7C48/7jmKovnaK71ikCZi+ey87QhZbcJKE4n7r8hK2JUB68j4Ktuk6FuEwzqLhT/KRk+W
pQ4iPwm6ZH7p77/iXHd6h4zKo2uePr7VSePT1EPKRt+ZYXSwVLTjG4eYVQRjpfOb/8UixWvw1Kk2
bAZ1TNYsGBFjJglkzHLtvFaKZMtDxPqw6fRsjc/PpNwz/jVGd7GEPfyuHsWJ3VORt3TX07Nl9uvT
e2uDyoQTjlB8vI1hkIISSZ5M0iGZWafY9jeySHbOv0BwJWmol+az9txrrjB1uT08TeiiOfEoViA8
LohB2MEsYJ5Bulao2HD8Uw4XhalCtbN16rIji4ZSLxgStxyRrAnyXmQIj7x3DoIMRjKlRh5SUi5a
3XemL0EJA8AInHH4Rr7UfTixI/KIczMmXjEmmtFHP4qg02yPXkm4llwMFRJCpsOhiLPXRBWPAgEn
d3NDrChfCBJzAmruCMweYY8ZpaAyFRwPw9vs9qwcRHFwHzNlr1GoXnJfoYN+u60M3qsThpsfRxt3
O/fXzVDHsRBLGzB3/EjeFnUF6XfoKmnTo0QXCfqbTOM5U5KGL64WQ7QnYK3oug3Je9G2MEjYprX+
7LYu9ODjamAxBSZxlM3pR7BXPdxAQlYdvffIsP6p/J1K4Sfn0GltUbYX9v+qCeK5M4w4Cydx4Sgg
tkAqjHm2qg4I37z4O1q8F5vVZ10WtNwCpgOnHxb5Lxpm7JDSlqPyxwUx/64idXJL7A00/6fr7z/0
pV0mFfpJQZSbPE34CP/utku4ux3wziQAt+BbAUPtHGelw5YmcSy41gphUDLRJyWNtDCssow4a4iF
o/lDbY3jD7FmTc5kD1SjdhwLkzRZIkVFDhgUQ1Q8UHAwnFp8g60L6+fET0ORL81tq+JXVLgmvjHk
fLU87QGwjX7dqiXQI/C+rGX/oAXu5Ox1mBv8wBUfEzi7kXjouUtrV14nZkN9NbM6Tg9ifTrGBmgG
QXIOl7XmetYQdHQ5om+z38J2MUg2dZ2xa6NtkeU7D/sp67xkvCLgPToNOscidCRNQu+snalliKb/
KWYjtkpKaoJJsZmvD7HUqw/bSB8gkXV1MLiDVhYRHkDnOXPJlhk+d8Wu1LAG/1Gtqb6XNKV4cY6F
6U2x9fjsBe9HNax7soevDpVTxCWQdufp/1ytSC/BZUx/Tj56AfmUIkmMgk7G4DWTjOUdjrQfqiK2
RZTqCoUuQWuBaEc3OlJ28/wUvhVfYuav01GNDa5QiDL2AU4Hwnm0Il6jP7i+G6mxhOTm+6onQjR9
7VPv0ZeTrlosU/sf4CIoonkOWZrYA0pt72NYMoA1iuvbYrX/havVptbvUW5pIeQYVPOh6kkWDKnO
PXN6zNuewCDiwsX28rUrC+CkaQhCe6k+Y23qXLnCeyZM9V8RSx/TNc083e1FjHD0n/AkuTSPU5F9
yPaHPJ2h8N9h9WMVmRTc/byc/b59QGE8U6O3mv0HqJg+RSJEXn8J7AjI3O0NkhfY8P0okh9VHGCe
sSsxdpSPxLeWJZnrD/t7YVC6U/n8S1dWAYS9PmPLYou2Zouc6mRqVVItp4k9AjF66/r7hJSRKW7r
eor4qqTcrUe5EuzShRg2K6c3pAb2+PaYa/SahMZ571rCQuQL/Yc2MGBtThQ3PjshssuzpyqfTafz
pk0CrDZfuxfu3mxheAHDVcLLR+S8hF5Z70m6GqXWsEGX17HRvhU+D2YWZpVTrNIi9EZvv+qStgtJ
dXAL0R08+b/DE8R2EvHLomf52QqPyIh+VvzXvN31YYg9+ENM83D/CPL54spXTFGhNZ41UBzedCb3
g3dzo+JIR+ROGNHE040lKyDFFN4TOhTHPRxf9UI4MOdWijh1+ZBhnlUb7k65KPrxX8/NEgsKfaUV
J8Zs3ZIBqqRzD7EkZWR7KOUwwn+VTJ1C+BBpwIDy0Aww/as8RFuIWezi5kogliE4Mew9Mf/CrXuw
McROjNW+KZIp4N+lWF+dzCJI7bk43zeoloiTW/6JB/pjoNb8PbGsuyx+FzJv8cd35evhbGLcVaiF
yS+pfEHRdayeCrK/inWT5z5hBwFMb42+PPnRMSRz7gSaK+dE71l4YqN8iaYFdf14FZiW6qUp5wWg
a0MpqXzbmWyV83evd/UhfgvcqgZN8mHJ49C00cgoEUF8vtAJUMip1CgjcAOP51Hhhcf2I9wn2hNf
w2lZoTCnjjZq3F1kU1piwJmFBgM0CBRIGa/CanIfcEWEh9JtS4+ocM7FnmmMexpB3Yt2HNuNzP8r
rESoNDHef6gKnlxDRzQwRMGw7TagvLUJnR9A8NlvzoViI2iRincGWCufrhXOoQ0AxXZLCkQvzMA2
RKqjPTb/vs7M+Yv6k0BykTEkWbjJEGIMrjqRUnqV5vsU9+EM6ybf1/lyGVSB2B1JQpH6lDxPpMUB
5YPk50JDnfYsptz9UY9bUGCwEXiVx9EVyHQF0B794KhZrjZDe/8zF9KO978/pd/CgynNPNLK1L6T
vQM73DlHW/PgSUrPzc3EU99xPWobgKVDl1gcp4KWwoXLv2jHizOearse7iTzdvihDTFT991wBN2m
FrPK7qBeDI1+Kf6+GwGYZcHkwEZJYwbR3oeW8UsL8N9LSzPPcMUzNIsFnGvma98uywoUT5pfMC51
/aVcXHx7HnxlHYs9p9lzZ8wC0s5XsOa4Y0P++n/1XgFOkNtqyQ2j8Pyt5/19ty2uqB/vxkn3hUdn
e1vTS1YruroKqM3BgwVGidYi5LMn6/rb8UgBCzCfB2mJGjr2Tjrg26aHrZ3gm7qGgvxaePHqIBNw
vIyyjEZ+FM5HflW+qTmoPtkyE01CCJHoot9FWY/FCaViK9P2+OU1ebXL53JgDv9UHX/T32VNaZ9E
YWFUPf7yP/lBrsAmoVdVe98eng5qw9N/O/WUD0nq19sByDj1PcQfmSXkr+bAu0eSTN28+qJP5+7h
qKmJYMCXpjiE1lTkeZV7Xz0W0JT22deUFQzb98udf5oTumZyKkyAB/dDADh94wPBjShilJGlDZAB
WiTOUTNT/QK/a621TR6n+0I/yDJcbYZYj00cty0bkUILHTHAJD0S2Uz57LYZTrppgmCOrwUKI4jh
n8TwSACldGYEuIcLv7C99M5p3p9Wh1Nat+4qK/Kw5eyqDQ5nLbfGR3+UYqiRwRMEN1hWcFPsjtGI
WuaznGnyG8f3Pn8Pv4+wzAGMNZNp6QFU83Tf7gdeL2ckApocSSDldpKQmcNRn2ahURKUItI1X3OP
mxBL1izprouNhSigHvbPbqo83TvGKvm7Bc6Y2VyYkY8E1nGHW5+zOAN+pGy0q/444HWCU7A1iMrw
R1XclfihlNhykpsG0dEF6Enet2fF3OoPPejzWwWZ9AwTx1Ay7+wXAWnoNw1Mdq70lTdkYGCoBvrj
vJNBq4iuDTrCXydU0FgvQZd/KYx11CiNP1+XcKBQkMuwGuRc/SyZrb51HyFCI6t0uKeMI5jYQeb5
p2YyhdZjUn99UrShUL5s+21RmW7EaC+KHAshvKhl0WmVzoBJfHrC8sEOGqrpQKTO1lVq0I7VMo2Q
hC5eJzjzVr1Kk84qx7JT9BRGkzIrZC44gqj9mbGnyIgcCcjZuhZT6AR8Li8fVzNabqPn7nYr8m7F
iifYEeDpzUZVdnnZjvOLk7E4vszO0pRrMXG+HfwuBIQYPgnRrxFr6OCZjjfNDFeQcbgmOT39KdQ/
5LmoJ/jtjLOHYa0DaKElHsX/fLUP4LJr1OA3cLH5ijk9hpCt9nppnryTQYkUaUDmTSBd0aVKgOFb
q+DEbkDveU+B2aWNscileao9/gIg+/2BXY2cPOe0nL+2HHfTZy7Sv1sP2XZKFhcZHjZi2ij2kZJl
E0W5msUtceW9rUxvD9ZMqmy/TUsESV6sxfoxQMgxRg3x5EYgUzsbO6935j7UL0JPCRk4rpTZhYX0
ncUlUzMiiGDrY6ULZGqUTi6hSXdXbeVWI6Uz9SZmBTdoUp75JdNWQEhzi9xSC/cJRvxF2Y4e4SwX
mlKJOPbBiSxVdd090qsKl7XL1EMAwHzZD4Tp6ygPsrfb9il2GJlrKVlwAFic674MQhhWnwmFKam0
ge/Hr+kWB9E0jhCR7pnS8rLxhD3+syxxommUPddoc7yEWj66tvwbulMaC4Ud5Hm2VgknRRBBsPG4
Fpx5sx+jYTd8MBNB/lmX+Lep+Ua+mzOOLTlAbrfmgU7ynswcSe2+6e1qfksTY2/5B621tBrUUDV6
jLpx5J6VkcsVxqfoTFtyDM8XOhOjAM5ijwie8rTdZM3Pe2+0Q+dkvcqfRqwfk1I3fUrawob0/mUB
8Z5GmnyjKlNDMajBlwkqvyHqGOIjIJd515E/97KEGqQJ6Q3NpZNvJ3P3Bw3raXB195nvSeo09DnH
PdO+awIlft+TntYt0+0X4e2QuZTinwQBg3NGeSxTBpsJDClBua4/czj+idZRjKLRMUfDPmyQoWEc
ArqHf+YFL+g5Z0GzyrhYjKm0ITIROZ3PPKJCGKAmuTNRJPUIudtRU+8T2iMntEI44A9rBsdRXyZe
0eejz5T6he8FpzmkJy1Jm0KaUQ/HThtm5wBTpC8+nqrkhfEQoL6/bfDP/JJlMk0Vd/dM8vb/vyii
t8r+JdA+GzNNfkHyjWYxdL8BUc6OfBE1uLbhK+mCX6lpXS28g6JUXmejSECD3jwPehO87RKNvzSk
07wQw+V1V09Ly4xGKHdikgp6EXfWEHZNEexn8Ps0p1y4zml9l8dEMRUPZ3GklllugJpXzq8jxfSs
1+cBgW3++LRP44IBnytoDdDeVgEOq3Uncy59gY+/wV9XiOLkigTH95Az95I+7SHtWM6uvKMrO0Wl
KZ4fOoNsSwQzenT3wqUUJIlp32i+zUrLZZsqyxr+5SBa7OsOfXl+dHmszSVLhlDfmEQkh5vEmcwB
LSjNetr1hJnNmTD3lyu1BMsoD+foCiTgQSe0BCAekEaaL723C7TxzMilx4AbJ5nJaYxJpkIBMYdr
ykT0sw4RvR27DgDJGMxWpnckZjw8vsl1f9ZBeg/Zi+SgVPM8tSIEJERWJzxiADohxB2N2V6Sw0YS
o7DmAmtWL7zjjgWXJV/CkRujZJmlyez3y2uoqV7lJ1LiNfVXAaIl85KmH/f6Wf7ESCZTrX3mTeqx
YfDgisxRawzhY+YHeuTF9FI8K551iwMXyf7pPOwJZJOgZaudcM6ubjOzuvWN1JVVBWuLFaQXvh4F
y5LdSF7CtAev9Mvc7KaWN/UhcayGqbkwUyEm1szw4PGMO1aP0PbuB6+38Eku/+Vm/Z7HabLgINsP
0MjK/GyjacmH3Ee6MWsly2mxBw3Ex4MXCPs4EevXw3C1T5ymn1n5jO0dwounVUOtV3CXfkMWOE5I
Vph/gEY/kAUm3Pujd2pE7tktN+uBCMkPuUew7aN//Kl7blDwnNUqtmHJqOvdV8fiJ8Rli0bFgJ8l
0rw0QxIsWghC6VuQEq26y+F33zviAeLBSt1wr961B4W1mQI2ffBUiwwUXo4yU6uMGOwHefly6vW/
sytt/RcBLhN8QkFovigQmvfOS+e946SdMmMQni7dM/edbaQxPZKj2AGEg6w1W/V4MSgmxx5b0yi/
8xC1s4gLkiiBfh3A4mpnikC9bLB8nUKq1G6MILuf8gqn2To/l+CRfxmeSylLxaR33p9bvql3Hgz5
wp6I1Ru59IjHMJfVEEON7X2mTZFPUm3s5hDVP3nr95c1+OXU+n6gxj5f59StDSsvlHACCiNAOQpM
DBctgwGF4yt7dikI/kuZV7T7/CX5fexxvt2rqKjorncvX9nDJdRTyT7xLExqVJV0nwfRpHJ79D/1
sRQtv8dF7kw0lUCuFslafvG9ka0f+emSUbNmQyE+z84d0HucVpfFiZ46xqXLZp9tFuLfOtywPTlh
no2t4yp+mWas+8R6SgGxJUBcJlS47yX6Ffo4oBM1hUuS4mdntruc8LGZePb5i3E/mVNlYl2/YVQa
Zwh9cYYCbOduZW2jILqKPHrLdVMhIv4+JDeafIqxdcfvGiCnjh3Qk2g0WjGmJdAkYyZdplCb68Ya
jP5lnCUJMSRqwHAkPNtchKlrafpYGE8+i4CvLptkvBzMXqn8QO8OUmdTBb+fbNvksKrrdVn0bzwP
C7ykJ3PI1q6xNYlkOalcOs5NTqXaT0UKiSYN3zlsOg1AQ+G0MjiCrSZ2N+WOjSDlHbW9U6BoRtuL
rAkn9A8MomFEAzF+ywotnwhgkgykk40CLKKWQzRPBI+wn848XzaIJjGvrZWC7X42jDoU1gFETeJn
1mVvnXavU8yO883BMM+u2d3VPebenmOwc9RbdVUvvOopVAO4iagAxdy9UfG9gQw/TghWxcBBB+LW
C3R013+JHzPdSsFuyEQ1en0Tja+NRJpWKPgeJBkKes+q2IQe8ggKLN7ZXYYQDKqYghZK1C6kOYgV
gfX0Ds4NSMC+UtAsJW0JogpTS3Bbk6EAJx0IX0qxog53WMCsHVB9cJyYfxtImrAIXJ0/GSTutkag
OygMFKQRfsNa/pDw0QgmX9pt6AA2K4zFYGArI4qiSKM5mSE75m81iCDU1Iu3gx5FlZHYNSOq7VoK
VBqCdUhqnfbIAT6Bwvh+z8w/m3FVM9Qg8WoRdUdHo4Wmw+oLUi9RdvDS+8wyb6LX9M6zwP/krd4Z
Q+B6O7oMX1WTdxQeuwnx5X/e0awGV9NCm1NllnrTgVFPzPUAJgInsfhweY8KFDlbfjwmD++IlhBM
ljnftwQesr7l/XkXeWprUEqFITIXWFOajCM8dnx3Mp4r2zh7cueURLnE33KZ9nF6NDL/ZhbWH0Tj
rmAr5pyD2N0EY4LJzYbh4GPXygPbx2e7d//w9nChRyB/uYrgZq1B3rfxt1cKuWLeVdAVQsXYdmFr
FAxiZooV6TCkn7JKsWfbf3n/RUre1p+idMWe+I6yICFg23aRn7oRzackHflsuVFDyNOXjwWjDPs5
1UaxH5aS+twz3TjDMoUnSBNAMeEVdoLeQ6qd9wVUmLRrsD+VWFW6z1IVojniuO+q6OlghDh4sNub
MNv9E8zH4xJJ10x/lR6ef/vgyMbuxjApng+IG6eqKfbFF7ujlhfuz4Kivqu/pTxgTJiB0qe8hEA/
fSkNBRUNbnYjlXobVLsY1FGGy3mtkW0tYMLTuihw5XWvSIVkbVrdbVcHj2o/zgXzCWfmeicKTd6P
SfIncZE5ccL/6WbTECJieLTq8cu8jRD9+6PGwPRVISJE5Nyf+Sx/DPVtdTKwZ9d1UWZSD9DJIiFY
Hm81GfzG9cmf/vcekfPgYdoGq+3pPRTu9mObKPRx3G0q+inVI7mb10OagOXGFIGBoqdPsfrCcdTm
Y985E/xJWB+cSK6tUzUYnensfMr8MEfGvNp1EO6eSScx1DS5v3UIpvUdObF91nF0bcDgflTggkCt
d+5tJOFUnCaCioSKi335P5HgS4nPGb4hKnqLS/FUxGFv+20XFUUjabvYEBNAuIJKU9PaAbqV+iQV
NOGCBs+kHi/V3i/7l97CF8Ev+bK5Y7M524z6hDcOQBby8y52VO+29QhLcp+1xjkb2plRgtOyrVuY
9JFnLfwUHVOt0Kj4SESf1ldqm4q8znk9kFg9uCXkJQgxIyUNeCkqileHjXvzJkE6lZvhxXKdKgAl
Sp62b7XLQ1TRhyPzDUDkzYAE5qFks7rMK/CE+eIiFoJhqMosUWHQSIFWhuagq/H9Nz5b/3xpgG8g
mahUcVU55N82VteRDjM24INVK8s39RyTDPTJz+OQJBNm7RxgHjEyMXAntStUYTjH64eW0v3PWsvQ
S5Bur4y2Fjm14+vk4i/jKyeaXQNx7qlLJyyj1HhDiHLOjcQ0BYq48XW6vZjDKrECvQyrd26G3NLT
5hPMVyatoscouPutOatoi4t7lzbEOxmcqHTSqoLtxcXG6PP/TWFq+7d8UG5doLbDr/VVzDvKZn7J
tjTM779ZDRB/xLNTy+92KrKKlB+RXqOlokb5xVQVpDfflVru65D/3hSUWvGHvz4MLn/S5HmeRUDc
iWI2tyAbQc1DiflfoRJ4rYoLf1vUa9FNAxsOg5Oj98nOYExFNX+BW33XznZI7orgNim0x+iAXMBQ
379rDwHp90eP1pv0DfQwF9zyiB1u4TVJIUgY9Jx2k9J+0oHSnZGc0ryq1pBk1XNl1Lw+q7cOLt9n
hv6zYla0xLTiBS64ZyhK8KzlX5sOW2Mxpoy8+N7n61IJMHTJUWyPoLCcPgGLmCGMeIQ+WqOGkO9M
j/Qh3IsTGW6P3Pg+My0LIhGqY9mUXAM3BgPYXVTulz180/N45TYxLrnZqJUuosD/J3hyFDq+Kpsg
Gw2XO2oEz4P2KQ+16LXaWfocai3yA1Ded7Pc5xAd8fntBAXFGMfcEQTK+yCijuD6uBkPMcqLxejC
/pCUuftpPaxBX/jTM2fkejddBhrLGWAeDw0MQsYbQSwwJe2Gg4dN4bOaGzO9f2eLk8FuGy7cwYtU
wx1Rcf2WEjgqgef/mx/xFo+LuNdLg7WSL5wgO+NS566RO3jyP+NK0J7tZHNM879zgrYLfEz9jaPI
2uZr7F/3tSK/p9DuwOPK4ZxVzihV3a1qvU1MjhBrPR+cJ89ni+dmM6sNsKnUiX/lVkrVVEFxnaIk
yr/9QIKZCSRQhWF8zPFTQ6V/QT4tg/knuX8QPqVLATRAT7uJ4YUscPMaZ3WJUGrbABnvp1qI5GBN
pOy4nq6KoE7urlBjXiwmh/yqw1O41/AX4Uh6N7jRAojRAHKzjchQurTD2GxEspyX0qXBy7lpr3q5
hrskfjkIBMiYp/zFzT2kbtFCHR22pHHeiJMUU7+iebfc9OpGKbilL2mjZ0QQYbtRCnC4BFz/9l/U
wPNHOOydiYssRKoPZ/mcVq1OMHfcDzXqjBswArs22BQmda573/Yy5H5slOb6nf+swOykw4AYvWlp
9mVuvPnB4OwfkhPDAyKNxrRfEl4eMIU25BA+x05MQlcVLJD0jShD4JgjZ46UdcvW/zEBAP9ydSin
8nHc5WXpMUNp0eOhaeJVvgjMOAuJ/Ta5uVQs/IGq/q6zgp1JwWOKVHFxSTCdDglnVOZEOiQfyj2Y
fZlZcYVc21yF8KhPlJo5KdwwjV+yT6SRYLVcsEiUg3X4zqP2kGtdmtX9arUbl7StrRZlq39kJ22K
yULuLFQZKKA0Ig01L5Syh5CGphI2c9OUs/TfTixnxGTqhHOcRDPHdllew2iDhzzfMjZB4FWIS6oz
PpdafYBWH2wSqV3IzrQqc27+deuy+TzYVS/laguAqgl7nb2886ljg1vUApdn4gJV811yMrgQ2v3A
D6ZP051QOger4qmV6Nhk1R/Klo5SJIEpQfuQf9OfH70mXsPRBr/hABOCmQW7cMdUT7g4BZB+bGX4
ucFobEd696p354p0Lw3NaqNV8quvoChUuc9NpIYyQ+QuzOqEalNKiV/qS/BrRnxNlk8wwiatXBou
BjyBxKgLxWCALj+bte8Xe/nIEjWoNhq4q1nB95Y/sfOpHegsxX7Qqqn/VU5o+ZWpv9uOZXRovcUq
SLlTnR0r13AODmjyPbK+Bho28UlNax1Tl4fVzxtn+KTw2FxBTFAq83qPoDwNPb7y3u9WyotF6m7i
wFZ9T3NaazE1HXi0WrDAovpFMV+ypEihU/JHQovwXPbfa++w3BbgPzAi84HURm8nMYrZpm5niy+o
bUU/3MlfYzXoZEeckwerOwwfTEoxDckH784l4LpVHGOpcK9tUUqEfh+6wOtiXF76X4OsgFrTgoZV
hX/ysgKITlNDbCtANI12J8qDDGk0HC0Td124LP8lJcLRJQagtzKjJFgnD96up9yQuTDrT9FwKVQi
85mzNTvwNKagVwQzShAtsYN9hJ5lmB9zTfPcp/ededggsNeE9Wp669SxOExpAvl8cPNzK1J7Qf2l
G1OkGc0FHdtrrA2HUqyECyaf1DCPNVwZuqKUpXVErRDawrCQbLJXhF3gGn4Oqh/6XlkNTWrtY3Rw
e83TA2QOYMvHeF7xs1h97vjf6goO0uPb6tlOpnjZW+RzBDv+o5SrANVsZvBom3fOXakgbmkDTAVU
t5QN20/3lIJxE73+MznhUxmJoJGkNUDMlpiGb9jyDhmcS36qqNyTpqaa0cYxYdM3Wnr+cPJE54tI
W+QkW1+hOtgpXhR94y6C2PD0ZaE0//lH6au7V2n2TSkJ6I6rOil07QfmU6I2tM1GtgDUvaLY1iv3
J7TocRWWZsffzzNb2BSVXGs/A3G62NFPPHCHdyGgeAzHC95o4g7QeQKHGA7l+y7y+rnJlvXeUEM3
a8Ns+qHb1pCpFLWBaeD6AMIZxJ44OJ5flIty2WvTzh/4Ar8RPkRDCQskU75GP2OmY2vuujeftxuu
fg3CMMJv/R2sjk8BxX5SRtgtDWmzngMRQyrp1BoRC2bnEs+sDrj/aEuBTmmArqWb+FC3YKjby6KD
dzVQkPQmtbZfHVsPS02QJwfvSgs3CkMFzgx1sl8fVjvXXAut4as9dzYFBbtGsDXxRZ22Op2i3GV7
TlR4a+Inbn/QoL2zutgYXNoukAOv6pxy+pOllpRpP5m+OlFLNKX1UVU+aHVZYdmnH72MZN9+JHVR
Rni8AsgoTQa5/4+KPp/zXabip8dC69xi1NHTMa1E4eT76iZjOJMm05IhC+esUJcxRYjEfXlOEiv0
C6iwceIO/7uhmVP9kH4Jv9T2zTcMFFcddEpGcXav0wQ+WxanVQ0lI32N5TcLqWhbdf+kNiuZMh+I
ifRH5pQoaPJoAWW/IuOoijoV8OAa6pAvDsh70ZBMdelk3RcvPo/GKl+aL9Ip6C8lqPHivycU/JNc
PhKkrgzumO2ZHEJgwghqz2UyIZas8ZqJk6Li5bLALJJIhZe9fv7BlFdtsDkFbfvLQkLI+q0kI08N
GH7eGbdU9+4YWjRXeReUciV+F3Yy/wjzJvu5KDI6/2KmnfJzs0gKnvTeyAyzQ8rob5xhLHnlRyJm
kLX18/Yr+D2wiLDLD3/8gb70dXmm9S/RVcZ7YcdCaECn6/lFrIWyjqDDC73K+twVJfrOLUjo3OTb
Il5lZ0dpAGhu5Q2W+e2qJ3MZ4w4TsDbfUasvmNDo4qRsrxEgE4j9P+m2YlEohZYDu8McKAWoRFsw
xjsLb1MkYHqy1tezpV32sXSr0bcr5bxseDQ8pn4503EZ/WXZwX+bc/L0ZmMeggqozfm108qSnu6c
F88hUukYcXQZCGo0qg/sFTz96x0w5bxP9uMtzVFDQ8BcISOIURYWN16+3lJho2lfRv28wuAefkky
Dz88w43RDnYLWcNRRzIaxpPtZ52IldKoGZ+C2s827PIp6GvhAb9wHjcpZfDnfe68MZ/KpZJOoYPX
3MZYR8QmUMMFmIu7+4Fs33rjNLGkd9yvRH6bV7lT+VxolE82lLtr5LSsCJreGlutHPZuWobgp45+
n2s90T4CR7ru/KuntJ0tkUlRdGLbjOdHT8LaasF80cXBCalFq6EXU+AySqh2dPDjl11I3PRAXaNS
WwmOE306/CMxkKkxXcQNOQ/Sw55gKr7EvVW0NMQnZBQtG+0lyGrvY06APqy0im8dvUDf6W6FUvN/
OEUu2Xffl52Aorm845bkPACbfBWEv0k5rInnpr60Enpl5nbTZaZWmrcpSp2YRftHvJzTYEsyIFUk
cJtR40b/Jsmhvp5w+gdz8tEd1qQSU6JarvhcnccibI7zHDYsxCzqbB/DWZl7b1A/3x3KF+9zN10l
tPEyx/xPZ9C+vJhgzzT8uqKwKaMzcY5MJZSZzgqPcRkkpMAqce1qf4K9+vsByfkXSQDe4bnse8UJ
ULxSfeMVOTr0kwaK6GwlBBSiXg3z2iD6fBNDpR4ko9EDqENmZ8nCADWP2SBZBlorXk+LlPB/Rml/
/2QRd4rwVbZg+UkT134MbM11iUjer6FYWs7WWQUhBQIOx4C04gJNe+/9Ebcr6QrL+1OgZ0AXTsYI
zBUcFyOw3hPCulIu34vz70YqtrnwJbIS1/dGHHM5IoPJOE1XTACw2vyRQ4ogH1hq/Asgkk5EamLb
YR+UWtOBj8O0fA4fUR9y+pgHUNdVVyu9Q26dphQ2k39a4M/c29IOy0EhpmGmjPowQ1GHMNTPtgx/
SIMq5YcqCdNE+QrsTaai7Ys0qVbKZhlzOR+58KWpbjltDUrUofQHFSEb8xUUqQlabkn3EbkefrKt
uu6u3T8XNEIYlLZjDgGjN2n8QhaWOL9SAQIlqrFMPd5oJdmYg8hBG5z0honJgKZGfKhJduIcHYv7
oD/ExD4Buhc2WVrbcAZXUeQWsIQ+kGKYeNbRcevFhsdIIfM9vi8W0XppUYmFqjJR+02WyVyFC8Ch
VJ+iz8UzphS/T9lxLwgRYi2PojuWibb8bM3gk7BGn7D1L8LnNG6czhWCalEMK/OXlsqCLgjFzu4q
/R/hPyhW29WjrBoJH0HhfRHY4gzMjaRSxIoc7esy5AEZ91W1nuNMKBXgZtbYplNk1s4AuKnp1mqv
+yFMY+N793xvly8ycrcib1Y1lHI5yrX1X9cZ2mEK/5SDqPMY3E1FMj6FI1scWLYHyFa/4uHwtS6k
EH4lhpq9iQMcTKh4rER0BtelqS5AqrBs/hp0kbkjSNzCu6/maE0kwVh5GWZs+02+yprQlJYzw9En
dpRLkdSp9UGHrFOx1oqu1bqZKQhJaKfM6INm5ET9wxYZVYzEdiSuCu8LMP6y/9W41sTTHeZ+9nTd
iXA76/pQsmoAVcHHno07IPvXY46viRPIUGEtI7KKLOa2dM2ojRNxDVWvy1pFGTqGNVqqelPtlizW
R84TJpJ0tzT8EMCcuwQwExTMSbPNctbNi1hIII/mcCSS0xp7ugmyaXltG+cYB+xOcf6y5HDfDJo+
qOJa/RsH2cZ6cCKwE3neVkJEVYryoik7WN9qkubqopAvma3zh8aY7yt91qIL+dkaYMB+PSdZipYa
3acC4zTIpD6CuiUMnGj+o/N7TvkFsydOG0WJ2V2tCNlbUia7OH0SoaIakQbI5L5lIdhXrIOvS2JR
e+E5r1lRgTTbBbJXmKrxxefs0Dd54mbOO/bWFr+UxkrYCz2zVnNMrMjfNtL3wEq2DB+A1ENgbft3
qu7hLzw4jVYziLAnVMRECHudHaCaQAXE/EwvvI+62Gs8I3GrBoDMMwotz3AJk2CgTUd0Wdb82Ckr
rFNUy3JZ+3Bt3ihwE4mjh0FAufsyrdSNTJVXthy13A2o2QVoizH/zcBmtR5hIM52rf8TKc0YSLL3
6TS/1OfLxcoBDHENhem6T8Z4kQ6u/Wf0NXnuPjdsRspLIO8StTQ6AwxF0TbuDkHO2hXLKBOJQN9q
bM+Xm8P7IsQlmf3Xb1ygAa3D5BjoR9aZ6lbtDRUa7iucuQ/yOiE8129b53IXcwO88lXtrgx4sygA
PbeCsVeFwsAhT489WMuGnTsaqyXZDjT7K+pDGc7Gv+p5c5huTk5PBaxVd3ADLb6TzVTWMNS0vSjy
Tx0mLdPH7WtRm6tcZJ2QiRng04QisHcGRMT3q0GDgZOQJFqpUvfJmWMIS1UnZwSsDFFgDvI8brM+
H1nLPydnEFFo9ZXrhJxa2B4+qaxDOtb/vyEdL60f8GpkuiQ6n0Cv5mN+pP4zYm3ihZZgAbj+BixN
aiCmprtPBGQe/1NSCiahKIaOiQRGlywkDAr6Rcr1uu/ghYie1KOs+VOyTjtyFe8EfEZu1xGHZwVu
wMxcMsnnhH1dXOXbJQ0KbU7GRlkKuVZQlozYX4JFlteiEaYhzWuC7ovc3L4fGuP6qJPwY6M/7sXT
PJ9NLVpnCF18d2wP2g0RuFLYaJn/frEAJyFXi9Q6a+rHpVJawTAH3A8WmhFUhYr++Oq73Id+gPhC
fNJzGTWW3qe9xy6AyvQXshebeSHgg8jHAutLxupkFZSYUe0xHK3DLbt4VkU7MfU+NWbi4KyujOY4
WCHEsZZUDNvrvRVm5/VX1WauSEh0mMv5C0ci3FOvHtrs4LNsYD6Fbwn317tlKq0OkcoGKdSDdcfE
9ia5N3vdH7Wy9a0Z9kjAtPo3PyonY8OAD04IHNgPG0lZl2RStjKVHKDrGY+I+ssQGD/Xb2aaT9hk
eb0gru9VcIcpYe5RTa3h7Wl6WSCFjowF4PixYX5jn/L4+2t8dJ4k69rQqxDSv6KnIgWAv7bTc8UH
KdK1Lq5Am3I1sPMYXj/mbXtbOA+bAt78jH9mXhzXklPIvgLYSEw9w0XUcX/P9ft3HRQFtlcpQBSe
Y9Jy4El1aDpAlz+VDYoxTdswXodZkhJ/P9zkFfZlcBXsh1adiR9RPLs2CsqJ+7OtpTi912Iu7K4C
r9O+AJ4bua2ZJ0lcHfKbCrYZU0JOwrj8tpHyfinHPo2vaSwE5EJGoiaka9nis6MaxHH4b/PRAI+C
Vh7WD2RFFjWah3hVXLqvQtWpwxqW9nEH064e/aho5fqvKvXTlKGa7iQx/WxpptyccD/gMgqAtbPy
3pZLyyNy+Ctkqwdc5qVAMJaxUNyramdaTmDz5IzTcOht/DE4ItN8p4WNrU7XtcIqaJris78Pg97V
dZ8FUOddB3clAJ+jXMw7CPpy23Yy9pfdtODt6KhEP19UgpNUE55To7nZhCd4SzLyQvn8lHnxufFf
XKH5OtQVlUsiAOAguLBqtatYA9kN1X8mcQfEfZw9/ADjWKMCYfYBXUqBHHSxcjHv139h7quE4+DM
ktHcOZo4nS8WWMAsfyjxn4z5qzemIuVS1OH5pOu+jnkQsKx2GCVAJoQHysZG0DvRikxxU8K7MUBz
dLKQG51Okl1BdhAkBvEG8coo2i0Khy1w1k8cCh1eSNf7FcKBGeP7K0o7EaCeyZDejXbC749HVJwa
xQLjrDZtBGaGdP6HccazAqBMYzVQ5zWi1fbWiWwhrmiin+TZWqK1EOZh361GoBihOx6zZ9M8hxsb
rz/d3xGNaTdotj6hLvKuPVLeIozXFISmhre0axv7JO/TaXcvPdlvynmdw9C9E+08d6UibTj021fm
7kBMkXWgDeJSCr2s4lNBNHSHu7WFun34uBU6aKnwytFMezPQeSXmVpliXkfaWwYJVXAJfZiWj3HV
QM3MpTdLzaq1xtodluXfdpS8HCTIHt2NsZfq0Bbg66grhjXGi766bT+a+VCDewsqwNEEcHCMU0yF
9+COBuwrksvWEEpnzxnq46LpCAyc/XmqIIGp8s9iHyCJPdI0WWWHiXx8RmRtW3+oU3NkAPupvCv8
wRkzQ+zAip5epla0ZMm4wYoUVvsFu0+Lmj8PNt2JzusV4yBRSx4YbrevNtCqS83fyrMFftqjdyvE
CGAdXWFzxebwTBYSWxaiNNjqNBAGZmzQP8BUHwCpFMWoEtFmMgWb2uG3tbsB8YHwwI0LxSPfMVxM
qrzPZxxCGXY2MBhUDEdtevTJNLnfLxYxUo7BJrAJiHT1e86hULXN1Q/HtzTuLd3uydni7F2ELDPw
LM/WYflwt8ohCuGjcUe4xBzzdeC6BKTBBFeHzgNV9neFrHHx/iTATaC/xpm1Urd1qBiYMg89/MkA
Xlptrom8RF2nMy4DND/r+lARLYSJs9krJ/C3eygtqer8Rtr+spB67Hkd0uVzEXwpyCjKtpbheiie
vvUAL0yTj4oI7vWqzJ+tBmjraGuQYIGHtFuy+5Ixu/vs8y9OgQE8+K8cx8aEdJQhIJWtwrvb7ytS
1exvkn7JL6/dUQfKBLv11h/RNHKHU4ZxmSuSHta3woGimbfdlWoqIb9zwAeMKvlTUsTtVrSU2ThH
eAMZOtEeFZY5wbA122w71uEU+spEch0rfEptxaay+X/VoIwqLKMTKTZF8jIoMUklFbJjAQhn5ofV
VvuJvO0a4mdWlnHUKncmwDn+0fhNpBHr3RV2WB0+Lz1IAnITHHxy8+P4ve7US2L121L/8ubRH0iu
wdxWfw0KPpr20eelXXu/XxEPopWXk7aFHErUUvjt9epS2IQNSwaQKgEfSK3w5v+OM8rDrD37sf80
5aDUxJx2MOdqzadUgn2WxjC8gm6DUs+gqPIEl7bR6zn3xFyKfEvkYrjV7VtEiSFueWgqBS9Knc5L
/yp3TMs2KWsAvw7WlON/5T/Lhf7NKYr64bVVkTp1z19ZFd8I/cpES2ChUYbzwTszBynL1om7/Fxd
gkQucrCbmnIL5ZqapZWWtngeZe8lpgEWfkkz5FP33vUyG32fCiJXvTwKQa8EHxjG1Sygs2dOevvm
cmk4213vlaM14ABCQTE29PWTMGsdzBUmP+WWhdMsA9wYQgWbHa+zoE013cecWyFcF4IBy4qnjVwB
WnXfw+W5wq5yf2WcKgf6/Av7G0nPrbL8IuyGLeGLL5bVZTmEAfLFecSVa5w0AVZXIo5w4hJtwdwf
C8Z8FMBxhBnwrkaSFGpt5YiahF9DYoYIdSmD20JGuQ7VkZ+zaywwIpJukjCJc9spZBnqzS8x7cWr
fbEK1dpvJIsrNHSCdAy/kstMGn/P15Dzh2fyM9XHEk+g81ydPUHycCLB9HMvngGuuV7S8wKc+fHn
zOhkMi3zpniLmiO27ikYVxFhtuW73MmDm1qNPliiAjsVcn7ZVcJjYHjX/tiRUlmZgzyNnLo9ADBs
Ttl3kH6k4krbeaXbdPOfFicMaWWdrZTGQDKSGTQukxu44nhOzBaLUeEpdAP1otDBWaqMVAw1fYZH
8Hex3tIeev1xp5s7nXDcqfdmHF5QU1tWwhxH4YoMdP4wBxvrRWstKFy4tFh7HMXyg2EJ7ISQY9dM
ZCRHgOsNifd/+DcRxL8RcQIfGz8o+9CPwJ2yRRmRHbsbAFKsvJFucDEZ/QwEvYdDARD9AQr+K8oc
lIEc2JUd4M82CQ4xfTlRVYejYRgYQkennkrVWX51asqgkYHqUYFmjI9um4i0D7ju0R7V7kLtyQ0i
qVw5ITtEge7nwXv/EuYrDKXi9sZmjuI2I65lzfFEDTgLt6SMecJVCQB/XfEctI0HRMr8abRvNRFi
HtjZ/RT98sGF23KA5MKTz9UuoXafU6w84n8cje275NRgsSgyLHcAZ5AOBgctkmd82wOTRzoHpMxs
lsOo0IWCvZdHLDoWUUi6HFIwYSfuDGNa2iXDpTH3s8Sb6cNIbIaOcjgUWXbXc95DOxLJ62yTMZRD
cUf00gTiOsK59uWbCeYCWARXfw01/CdpYhyslnybZRxpgcYz7IcvDTcon3MfBl5SuMDCxw/VaQjP
ilBp6QQW6L+bIABwiCJ6ZxNtETYNdo0ipcUgqqftrnuIVi5kFl+3luBtGsorsocU2wh2/CjX0Aoi
S1JBQHSO8e7ONnRLyALv7hJLPsiSSzLewOASm8v72VTml7F31e6u0M5QxDcZR5DURjOM0iZclk6q
IpYl5BlAH2eHNGL+C45iSzvZu04+xA++jXG6U6NeWAt4bzOBZrTJgMP0b8ZyUEkvgl51qynqfBDn
bDuL+XADX3CI7HjYvmMa7QZQ+s/cAJVHOJrwqldEJ24f757rB5uqU2kyMVQ+iXmREW7PrfINGM9w
rRVULRIMwlscr03vuWtc1OjggmGAwOy6tCKcPhsyrlqqRvo05dfEPWKWRvBytI9XFQxWhcKiAlHr
hqph7o2IYOScN7g9QoA8OKo5R6b4eb1SYfIpMMLuqMeWMWuOKLGN1rPFGhK9D+XtQt46Np0SisSP
O9Pu0SKzfVC/N+w4j/bcKWFFeWAoXq59IDro4VtcWuhREYzut5+wfNwYCz+gWN7/So+9wkI5TvVx
tvVqQyXmtshIygOQ69dePPzKF2yArDeF54kHRtZHBuQu1glEcEEnJHhA4olPYwPl1yknrWpOud2a
ZlBQ2WZ4tSgiIu94OETSJWXLMJEDHNsMfdH3dpv2weuD11GTQp7IwfDYTb4xPziNKFAlTcWZGDm0
AmiXmnESrx4BqdkM4wXHhzZx2/dViML4r1jjyjC0CuS64AHaRZLBOzv13HLsQhB6n+6E76apqX7h
G5qGYZqlv5+DfCyucjnDFiGEiUrG7IyLlTn790e4IoY40Xw+NDemOTDDxINN3fvh7Mv9H1Zu7ut/
GF0ELwh1mKEoUToUYkpMK/SEu4gnjrgethcBpZj6e4l/AGyJWpHaiNh1TD/p2DkJlEA+U1qQrRBg
xaJDepw825IQ3IZZh7gyMQyrGgcgHyhrXL1oIKGJ27ph0faAVTc6W4WyFZaej1TV4CvQ7WZ1qUCl
78vmvPFxtwEfQ1Ur9+p04LVVqC38VsztGEGkbBcMgDu27pEfvlOjn1IgQ+tyCi3f4OlsKRuIPTxl
B/PCGLrOvygiL6hBXeUyYlNqjNLyL03MD1jNeVSJZr2yZeoR/IRYjNBnTnr838/X+uHgCHP/uxkG
uSBu6lvcw0VUCufx7vLSunVgQxf6OXTAJU1HvaW/e0pDIWedV6RsZZP/LqrPHvuRj45J4MSXPylo
8rOWUt8tfqkEnnOqcp9Iaql9xCBE10GdwPxbc6DNSjbpU70Xuuk4WlSCReGvR10aebBGyXRtS9Lz
TGvyQLtEi75T6yzGzsZKEP5OTMIaXRZP6IwldwiXPeQ9bdb45uhxs3fLk2Os1/hl4dRzKHQgLRt4
bZXilhFBdtTszItjqXoWYbIDxdicG/YC67pT2vYIC3weBXiKdAPeUS5ari7kIOumlLtHJZuYSunZ
MJO8Kt0ia0cWSQxwlnsHFMbe8Ad3kFCxLkbOLZ7lpC+vYYktqLUNZ/ua2EyF0zRobxuORdngraQx
BQvEI+60o2PmsaF2DjUd9qtplDvvLmMINKduQ7aO9UuPaMLl/VpxeKcdHUJNAdzP9kFx9cDiALuy
wES18OQamqYOu+rDX7LX4uHN+bomSbGsKELVZagljRau7z5w5c+jA4J54+3utIopfVlixew9NvOV
I90IX7haxMGoRfO+kHtO8ldFNfbFQr56TuhDMbHt1coGZM7Qc8c+hQ8ckAR+YfdO3wPZGmCSW7kr
ot4KU+WMdmaaTj7wK+mBSYlVd5F6RZfZCOT6KwGp+vF5P42URj/Dm8go7VJ2TYRq1NGqM2bVTbON
rhohdhJ77BICqe2nTuGaZrw9jai/IbvCYaC4/PXc7eGHsB9AcG52qt3jbO3R0zAd2Rg8qin/u8y1
enzIf/IbslWTJbFwcASuQ7x3wAYhwcL/KskgECHpzqsH+VsBijPhOmemUKqBGRmEeqpD4BavVLD3
objIltQknqrXknL51KzTuxcfRXsp0u3dhnaIRTQdItw9nMm8WFZzBN4dl0Z3LpcuUsGFbpEzaqAr
7vM0LwHVTvXCyW1Djp95HaP3OBQbQV5kao5JaCk//uB3B6hGA/izs+WANC77OxPKuIvilfYSyS8z
IidWAip/3CqgQ2Ypj0uwlGMijaaYflNdLH1QMpfRNCZVsWAwxLtpmIF9kefmV9tQx3A0TosLU87Z
QQS8bhzNBB1R8/myLDHEkWPXPlYBjccV8fUFT0h48JnJ6F9Q5j65rC/lISx/aF9DGsFTTBF6cweV
X4V+Fbxa8R58lHGUpW+jQL+jrqqENtIPh04vfhULv2vciSYDiXXtQMeUIMXhRADiadwHOj+1HNms
wWahqFimWdcvrfl5DO70DiStZNSQzr2pP/bRUsAU0YkrmpJCJJkFEdtNha4hG8w0E54Qhujx8YWQ
r6LF1jsjv3Zwv031dZIvWN9rqKQXeHeyR2N4LDFD0ciut0a0eYXAwZKSDTCopxldOiau6k5nyAD7
5PKgK/oda/rD4naRiiQzgpF1Z7++QQNqiipJBp81sRlmYVq0DF23DGOU0CYRH8o1H7LsPlKpukYt
WJwWfBFoEx91xCfHMnjEH9O0/QWpAkLPiqUz2PPKZsHG2FwwtaW9oBRb1xI4xDfzF3yu61a72rJg
MMPIIDxTgozv8/Of6kXfhj32K/7uqWOIZaK7VSnSn99OTZV1pobsWWLYgPsxGG4HWO6/HdPEEWIw
EkWkJgU8Lad1I1xKEjtx9xuy5eLY2iMQar7f/Gh5YF1hjx9sTDk0Vqrj9IJXV2de3/1IZFqFDM13
f6ah40Z9kOj4LkRedIMATv8RwS8d7bl+4iKbHQeYCLf+2nfEjyJoiFjRxPFlHNXAVXnbSep2delB
fur+celUsiGSNS0zAiC4KdN7k2ZmZFjg41nrV21+JaNL9gPiSYu7J9pinkw6o63r043h+um1y8TI
9PxfgPHfy7U2EOb7JnPZ0jIQYSvD8gt0+1yPBpO0hBj/EUBNT3/i/thd0FEh4GmKDNoUJDeXpIc0
WlyaFI7uypgjr4dfA7Qbe9zlD6Zb4dv9wSEffEnjEhv3dbXed/NKA6rotz0sg6ITpEMiJXpv8bqh
GRORVoZ9EgVXP3O9w/f4HnG/gSdmleWDvs2nb1k0LlsbBUt70LOqnHk04T4KigYWgsfCpxt/gTmE
LToprC1KLP/cEKgImxg+gVClGEfWvmiQs7RNBrS8m6LIjOyuLZ1k0QgcMrnBXhTHunCADDrojmM6
EMrSzyhIWxUWjV3FcqFS3OjTz0Z5zhkBc+0/1uJo/NN2DDZt7X7MaeZXUi0NYP1G72pzeQddJErJ
GzRmfN94w6JHOQjHAZDIjST0XCzZ7o3cCwT2jC0/NaVOugXZcjnDUVFxH51+Jtd4j60OWhJdS1x6
Bpz754t7MiQ+FDlBB4lbRlUtk4/6gdK8HSlHe8oGX1RpxsXAK06rkucrsFj0SnyEfUytoCGpph2g
PcnCrhY0iQG8MlYXKxLXV/3zi2WRvPbDQwjj/NFvzbuMDxejlkET1qcslO+xspybtdkwQWRltBQj
BYzRKu41apwHvr9xrsPgL2RQ5q9gNNPyOxatBTx7T3cciMCmHJRpVzqhKja9b9TWqKusbYxsxXD4
wPOx3SB8zmPQqikDhXdqmTZu2a8ily5iljl+OMeoYo55K3lmOoIaU8d05E+oj3pV8J/3zHZVAXfN
DbsBALuRhVjAhLmTpSXO7jYOQlyKPmdenRA0B2v9sUcDpum5wdYfcPezrlifbR9jdXz6FsHSMBev
DTUEvQ1KPP+bAijjPvov96OZ9tt135qYQDmj2NKRDDGlW4GpRFKdlletB9rhNUf54nuJ35Nz4NQN
g6e1Z4k5v/8ABiGfqIsFfMQGKa/cqUvPlaUG0O5TL+vEuNsUzrXIoNJzg0P9RA95AvfesRxkHm9Z
I0BGEJ6pJK7EfT+VWYeitfsO6nqSR2p7Q7lTQ2EeGFy/TqSJNKmVvyN6p17R0zx+xuIpLWGHdp+0
b92RC4vGKR9tRCHAqN+pdz/Njj8rLf7P6C996y2iwk3dGJuCip8A70/WcZpzwn8DQvTQ6s2X7TPK
d2mpC7/n8ocxGI4Ii4L1ZF7NpdRus3J0G293Pvq7FG36PTNByFgyMl+8jhGDnktY42cN6kY0D3Bm
8B7Ixoik/bxYI2UaMxELnOnWcPy2ll2lwNSkpoBnfC9aZwWkUJRcxZ0rlX1cp9qVg+Gz98PzkrUQ
GxPeV8dZadSiMw1y5cDpxxvIa1mJxSyUEEv4JQPiGCmsSM93piZDWYci952CVPWUJp2tv0EihNe9
yzWxcO2nVpG/esYZPHF2LIEMXiGMEKwP3nUAE/p537hZO0WIO+NWU0dYlYvRW0QbPf+j1I2qhBrI
UbUB5t6Qq9XvTbsaQfTRC5eot7o7hC3l2kQyQiGiXCKjaWslc7tTOTiIe/qgCEjHnGj9uKXvOfsm
ZDj5j3i5Z7eCqTfufBUWwNt5qBJ8G34kAR9pDzN7Rozq+ErWtau+dqtaNNyWeEE2REYv628sZz4D
XeW2MmqxC7UwmbICXvwiOhWJHt1rH/KeyDX/riiyChsCReSg5+h7V9obLV16weWz3BJ7ZCDqusxz
v0tGSYFQ6c9wFo2RHq96nuXjiTnDUilxuD0lqbIhVBNY1GuX29Ok9qDqR00WfTLLootXeD/uuY1o
/LSFj3YyzL+3mRYvGUqrQ91moSGmgGQF0y1fbH6XBSPGT467Tmn/8ELmOLouE5mn+Rt6MpCyUos0
uP266irlrL59N98U2KBsME6Qcbh0ZiZ9fggAfb7sYMpDGaTwJoasMCsNzEwf5zdbDEqMy6FJA1Qv
esdL6TLOnzKtcQ0dyM2nQFP0Q5B+2hTO5f73Zih2wFFsgg4dbRHgheYIkCtCac+JzczFpEmxQlgs
JCeqZOrIJuAMSwUO4CYD1htjV2aBmRMQqFMvy3K7FXiNPcMv8IgGzZwciz2cAj7NX6dhy7sSkxi1
CZLGkUzjz9S9N/zXzcrty6Ox68BUdEZuXt5fZWtg/W9UEnQnLni0rkSc3DNUjPaS/ioYnggDPwtV
NLSSE9AI/2R/yBJIhRhkgG6yZ0y+kyJc2+kl8pWOxst/OdOGGuotgyvLmQsOkM02lUGms7Y6UlaA
U6/6LQ+tUNv9/KHr7Vl3nDA6k8Tk2z7CSj0YTrdyXlwLbdOCboXSUoK5Q4iPkI5r/PrwhUw8I0Tw
APfTowlmMyiMGlbHdjq07ff5wmmSEhB7FWp8H1Zz9mNA2tGKF6WZiCrnFzTgNuq2cRnqF1af9ezd
LT546o8VD5CnWgHm+pxUwT3kiQlz2a94Qa9R4mJdj9AIYwfyo0qil7RBiJQEGYGtfxzupkFEN6cv
SfFReFCsdodVn6PN7MdYyxGyWTxPZ23fGcb/SDGegC/sY+EP6ciSvpyP3HD/Uxr1p1elNso8XBU8
IJxn6NMsDSUhvCf0kyQFf9Abzao5yjP7kCI7uZ8w23smDkorQJHiRjm7DJO+z8Fm/rRKrYSsm6gj
1dYcREk/mLlEqM/2YedqUJejHVXa1DIlB3FKj/ZslD8q48NTdDJRJxD345bMq2GfI8DPzAyJ0C/9
H7iqyoYsN8G6I0VbbDx/Cu1zjIeMJbj2j3zc5iiL+TEXQ0QlShq4PIE2jlCT78h47XSi3cQtgoCR
3t0lo+fAFBt883fTOyTFZeOZE4kJSOqtRQsA9VfNJ4cVXg+4RCSZjMf/CVPLS1dQSY/WcPZVqImL
0fpdrYh/lwlhpaG5qapifULoM/+F8oroPkwPjvHSQaKVCCwtiF7yxi/YIMbSlaoYv07Xn0fpERPV
xWTDcTTSo/vseq9O5dvT/VBSnKiejgPMZ0OAvm13gQHmfR0rfrA3Nn1gvvibGEvCFc4AtI6pMq9j
JzEVwTprx2UJD1Xbx6zJi2QVynJlLidjO75Ci0PpRT3pVDVbiRk9Sdz9fZ0aO/gDTVICiqF9diVP
+TVP2ywueUd1g8P3T5MLE/O7qJGviQ1kF9vRhbYFJDE9N/d2l/JDS1px7rDxKxi2imOjEnJyQJvb
sqG1pp0aw6UfbUq9wATWXzHWIz6UHD9Hir7cvWVAnMAJ6Z/js2u8Jr5lzglTUHfzh+EwXaGNjCTc
wzWhemaShkpRbOhWoc8Cke5I/DTddpBxDcXM/IHN9WINbShe3JyLJFn2HLhdwr8TXWjOA/UemBoB
tyQaixxikpeP/PGjo3E/rbEUq6Wd05dIMqtuYgPpmNg5+6o/purwdDtfTINLFjTSSRI6t5IVhg7U
pC3HLe1XdxShE/Ly00A8UdpECKpcWktQVLmGdivHsOYpycXwOnAe3ZXEFvMyRhaNLi5lTApXaM9Y
OrF25iufgxawSsvNF32HikfWZ9+izW39buU7fQHgcXC1CtgBWAKC8k8zZAkpUKXxn3/u2pVsKeT6
RjdTlap2Nm5LQodSXfTddIhauG89MYoAKDBuKS6+Ez07FFzahZFEXGE+6fZ3SkK65EAjGimYIvKQ
M9fsdL4XxfVUgv80RjORwHQqzyIULAvnMZyEt70s3WHXtMcLLT3lt1sUqwF0k5pRpeyo56tQzEuF
mdTRNtP210oQGvOKUt7Ot/rl7Fkt87uUTUVWEDQys5G9Cfm1b0LJ3hY/HnAMt/R2ThL/gPfbN1Xb
uTOxb4Ro1idwh52iz8v8kZ+2HNQx2ZH1V8bJ1fsxVE56SqJI9xWZo7nqL0IatY8STDi0gSMgArHk
jKmt5X+g6i0TUtro8QFLeEKVoXKeQk8O4qEPaBdr5740oeLas8PbDFTkBmREcCiXAh60Vb1S8u5y
sD/IW5D92QxEdsJReNd0t6h422miSH6dCkYa+l5tZ/egmSMmDWrRC98yHzYIZsjNNEKVy+gfGvwv
p0pn308DUR4sHRw9puhZhUPSoX/SzKrEELsgmnX0wCC2bnmRqFb+W5Z3iwmIKgZE7bdTtfBajxnn
ZGNF5G+om4gDCBVn1N7w25C+gSTK5MYkRkGZoJYt+9XBiACsK+/HrWCigArKK8pINbSnwvNxjHv5
s3TlWE7nDmERucsbumZ85ISvvI1qZz8st3TItfAFePPfRiV5/Qzs3b4zDta/Kloz7M2naPFJ15De
jXQLFU/d1BwYOZmv9mTGEaRKExDOB6sVtz5BfXK54D1hehttdtdzzaAZnk+z9nq/S9ChcdIizCRZ
Wr7/vkxAdqeJCcKqAhKn480p2Pot0+dhJDRvKmyAIT32nBgWlZpGuCMCWG9IImfKOXA7Bx/TxCME
93iFssDr3cGloZFcoNxegDqbbJNH+8TwpyA6QXAfMIl325cnpFVuVuDln7PYgVnLKDnAYIkl91nD
4MxmFP4gx4YjbWHebMncs8DhlQKvSec4HI62V55EFH2E7psnNpL9im8DnOsutNwmNRhV3aYHwaOR
G4AstsWzCv5oJh+d+uNdYgybqUStpZGoVLDFdQOtSPOeLHM1rSJqukXMRrnui1o0TZj9+2MFFlfI
ZFDFTWzZDQ43swrs1Aup4/RVL1woL1x7vrCJ88L3PqIDe47PeLq2lwMGhTmz3RnOvCNhp24Wj5bn
0UoM/WHopO7WZB/Ary+7eGL9AawfT51nUhJepPLyE3vHWiWlRVdAN/3Gwun++TjIH4M21tisNkHX
18c9tA5OeHf3DvVdQ7c3hJL42S32l3+Dsg6Eslb133yNSfJbGOV3TRd1EyuCElvQHkhXoerMAU/5
ngWEt8+KFUWmGpqRsRBFfPcXKwPxNDLRYnT0EC0p0JV0S4vcYtoKkqc0ZO2uLUJ2AeFpiJX69nVT
A7hijL6ywdAomu/xN7mTk+1HT2D23XgfORKITiXrFcWKSMBMv47QAHrodGlInBUAFtmjYIE8be2s
cVSjbKsto5uuChi82E7B5h45udP3U1vJ68gkBB9QtFwpntFXxB3iHrpmWlIKM/Z8FCoMfHgynPOg
z9ZmKYGOFZXYhgKcpXBQxHM9DhyLWabmP/GA06GTGXlB6Ri5W43Bc1HG7t2f4FVmRhcE2CqLbOnV
x3vMRmjXAzyDZ08Arsmvi8EcBsFCLuCFml7KbXALe35ou29Di+S0cxLD98VwcYbQr/mc2Bkwcb25
YRUcyQDM8kGkoslzJWJ/3CqqwB/aEK4Dl3smg+m14WY+BJD4LE3/k74+J2qe8knl9MPUhmiFS82z
JfPgkAJ0VI8h35OK+c/LaD28g1RjTMuNiIo3FnApMlXiSYayvgxftfC6yfo9R8TcRRql3NXpnSgh
SmYEqsZnSOmvYteccBIXYhHwQ0+1qmjk9zIJ5dKeTweXA5C4n9+1VOL+l72tGrzCe9nDsZ1uJbHr
6AaxXpVwhfnWrtQmCMmyRZ/pMsKogW0xbVQQyIRwn96bF2FxXPqM3NPrMS8hbG/+g1Mh+lJ6w+YT
EkktCM1SRUZVA0/im91SSZt90JwMfH9GBjYlyBjQJzsVZ1Kndu/hoRkU9EQkXPqqwrowsMs5V2yI
uI36bIgwFsyXosTsoICpYj3Q+mAuVU7a7STPeKfzSHbn43obZOtBDwxKJqrHug7MPoulhfqCMHNP
KAnfDj+ZWQ1gjNkVEOzfv8IIK0SRGwmaNsNlD+E5Av5rIExGs/FXe0GNn+c12BpQCglSx5FuEvvU
7nd8628asRSHE+GOd/MGy6a9Qx8HeMMINMV0UhMsW+h50ey15z6QBsV97CPB9M7S0y/PrQ5XINsc
8FfU2tFqcdA8DtMCwiUXeUKAZWiCmEy84Ra/prZ/4gCYIYKL4cFihhHu6xuN7FHlZGadn4/5v957
EDi7jMnnxUcVRpgzUSujmqetZmX+8X47cd0VW5ka+TWYizvZXSOu6rcRcJMo1fCTljVQuJZixyjy
i9gFoXL1cN2T0i2RJR69d6/ZZGYY+0b28RABh8PXr00Cop0VwPZW5RLaw2Chp981A9K7dsB93/tD
dI0Ku9fFZZMjBbE/bQuvrlYHgecJyc+qe4BMq7q4qawhGWLpHv8v0BPPJ32eZ4fGVT49Ywihe1Vw
pkpqg48aYGLXhHvX5mUDdu+oTQ4SrvM54Tlyt/zWGI7KjdCYAc1I11YAicGSdnjER9NbNjuD+K4p
AWJ76P3cBjrEgVKObPij3sdVwoVLzMUlEeAwxTZe1I3spYiC0AeUucs5xv0Djd/pdjGgWvg8zUw1
5F3keLrEswCcffjAG0Vaq2jOHvRsETSqYf6D4BJM2HbAyOvdnHRJJqEejIB8S6fDvpSYNztIkPTl
PbficgJuLauWKodq9d85Mx6WRdo4qsooMLxjjCV9SCHtsSNRl7J7P7hZd7cMQOibJNNFD+hjL2ZS
soroyxVvBbzM3tFR2QAPze30NOCRyq51eMxulGk8aVCUyVIAheeRrxe8MwfJz1TixrWjgxMGmWUm
0CZ3NDBMg/2cifCsgfq99TAiQYTE6FfJ8FvcC7qMjoFOL4JvhFd019R/r8zpiMCd9fzQbYvNGi2S
glPlUgqZVP66fXpUhJ+XnNZVV6NXIOMUxz9SQm3RuKebvOk5SPir0KbTzYPsdx6ifzdekD7/FaFn
ZYxBNYvoQXclfKNN7wqKzTNlo/Y66sop8RJSC4ZUv4mslPqOyKZKrN3XgohbjoM31QnzGd7xEeyT
44jlsG2igCAGm+wADH2E1MOUgtRx0DUuvebtE7AE6tNCruvu31R68y1GlZAvkkky/CThYdAmBWhd
MPAK58TMb2X8NswfTQDHU+uTtyr++6tA8mI4ylfKyVfuTRmmSzAPDe6lfhcAgG6Pcle8QUqOGp0y
luG5MUtsZRVVIagIU545MX0rawoGWgUMzfDGFGweD+vdHG0/EAD+C03lriznJcXL3L8U58e/Qn/U
8Uof95lficRoObaLMu7UNdQFlei/nlXXkFtWleh+KyimnvwwtqNZb48nJxMi24WD7sxAGvEkJT71
aB49YtBHiuFlsB72vj3aLMKSBAVQ1HX7izUgj/Cz8fBI+O+2CbHMF0mddc8ro/lxoBx8g/bC9ubf
GLXfagsLiXOR9G94tW5/ahDoU07++4D0HahCMxFJNgJfedwLFNToXqvXPNgYV1SLoQqy4xhzRB1c
ZY3/KrOcHI4PO1eWkuQrLDVeYAj6w1lKdZ6eQxjnrOR5eAVXEO0rs7eVnJQLkRSuKVwjXXzEnXjS
HKQytf+9D3310BP0vl7lEk2r/pYTFU1GrIbW78WNUInxWEdZg47cZgY0b79j/rdm2zlwfIk1sE71
6sgmmEbvSG+MZL3iW4Y+VUSejhmj16t6AAhLA2L1VzomR7/SxonuXvXo3YAbEf6htXxkAhdRe8po
qkFCNIE7kn/tmH1d3FnQIeK9VXxq1OZjnpeZbNrtFCa8UlkhJxB0WLrEXQ98VWMvrh36LhewsLf8
TU4oheAGLrwQZoKrDzFUDO97gct68z2vShx8nKI2DYCaBKjGu8B6bs+LUV1vmvR2QCwwTJ6FKSq0
DwWtaRMWnuYX8AV/TTl4bV6pI7MOzRs0Sa+AUg1uVWku/yJ2WIxIqVBJDTULvvCQzV4QwSzc278b
i8RTc2OJdxVwsas1XB9UpQMz6k4EePcBb2zQKDoVH65W1w1S5ujPhp5B/u2nuN4X1ugYM4NEVzAb
X82O0zZZHQMLDsZR2JbAsmTCGEpm/ZS9gpXcWtxIvphCBhmxj6HyHqe5JWoPuvJE76DAz0hIxIQc
oM3BMA4zHlu9K964b97ivRjDzIVUTjiFABRI5SBvfPtD5YcaUBB1iBk8XRHHpTnXlzKWaaAdincY
Eup5XmLXQxG43E0HA7PrVab056fDAG0RXLeC73NiIBhBIGWDdH52gFYTAGKRam/GdiTJsOxy4QFK
THXdIHbRz0v1sSaj0VaY8Ah4pWHZfTHdN+6IKk76Xdb81kXmm125ir5+OmX7tkSEbWhfQ29mPssv
TEFPY3RIF3W/N65glDVIkMoLz7/2K3W13b26ulgf+54AErXb8SDlLk8sw5WMNuhMYCwDDIvL/ej0
B+vORq2LRm+SP4LSgXKMSokFakbSaegk9YyVHdf3yoAObgyIrNhdHlECDlqM+UaTZRfP4nCRLZNt
sqoN07C2l8jVMJPn7sLpVS4/b2EjLccfEE8+3inCPacYk2RdkLNgNtdLT8Nwhh/SSKrR2QbuognI
TwpyfILedPUXqC/e4+AFMf4V5Mb+Ags3a3Afu7QCWgB8fmX+JBHsafd5YdpWVg8OXt45Weu4HawC
EU5LhX/UXOWwDTMpQCtFpgt9wXYZXQUpeolfG6kaJNIV3kEYRQrsS5ISOSmHdXAYeLNZOz90D65y
xze0czULAbFrwrSyCWUm2narqu8LO7UX/BeWuqqiS9yCVsIIBtsFgBtOo9o5htPv6VU1jcuzbrb+
IrSmTZW54v3j1EBuryRDDqxwD343qT1dNO9Nkgp/7L4Lj2venzIODAzuzyLpRAZGmN8FnlHpi+nr
iEA7onS+A8Bgboykf50QLCKkjuTRs8X36JJ7/BtqJCI8o7GmEQo5t/ww48Cg4EIaz/LaZZcHdRP/
J4XYh2k9p51piGd5CIVX1QfXxIkE7L27GcXhjaYH5paKA5jjfmoyKoNZL4GscJJLlH489PWLRAxk
Xby5uWVWapJhmu0E9qM4yS6mbPB0p3dNbP848afuQhFvM5M4ok+pIg57GwMiSnPA2fF8p8UcM+jJ
YGGdTSWU30QYrhO0vUM1kBf+iPee2sIBTAXJKzeA6KWqg9B1R/OTkC0mFHWfqKuN39v9y5tkZu+E
WfTpqqCTYLTuohFkIxvJe2MVjc77U84lla0tTdswX3tFk/rAsv1Sj7lo/TC94kIzbWo1wnH0s/Uw
diOsxPxZgu0tu9XaR2A7XZbCSlXnHN1Im7IoMi6siSWy/vtHYTDF/8lXU2EmOCIGnwEXe8ODOu1A
5X9W6wg5fr/vk/ACY2PpvRQbzm6xIMVh4QJgLQvxQzgr9MfQztleoR/GH+Mbvo0/EXeVhfJXAJL3
QyRPJ2luSIPfYEzuTGROrMUGcOtSInqZx0cHh0EOamBMzvwisDv2Veh6z1bhabpEHAIp2ucrEAiw
fqSs7eic9P+Y+ukgDhFrAVLdgbrpz/4Cp6FpG9BaR4YnsULGqjX3T+cC/qzPpqzR3UnHXoSdC+x9
LTnZxN6z/jLOTCJ1BMNU16oI5NAsvKoR9t56xofcjNXV50UjcCYcfdQxSTvfzL9YXMxmSPMDURvF
mNOyKym7xAr9PX/sFgUTmONa9AIbE2tJYMNNjLLlhlrZTYbSFYOwBIR0W4tCWEb6zfsfm6fKcmII
kjx8z4z4rlVKn20TiDRs1AKluT5nPPa2OKqyh/iUxFkCMuCe75SQ74AEzEXfwT8GYfIrh/5WUMKn
e7hsPhWaTNUe7TNoBZTz0OFdf4/f17oZYT8eiMZTD0jrbCeKNRaQkLqA2lLmgTga3oH687p1q2Tm
qKb4IcNEhZZENEz675Feuddoq682/X5xJMk+oxO2OdLcdN+i9Ed8VQqAWpBZmNSggjEC+3j4sDd3
hoKJ/p+y0wJq5m/VgojdLgcQKLW4n1xOMZhdIJqSaqq5zz4sPpApbRsIHHhBSwJ+OwuIl2pUfvhF
AInnaFK8ENZ0+MUU27Ju+U860OVt5Jnnk548zJ6q1pMEOxt4kBblpB7b1soIVu2+vJBLnUq50amS
GcP5RMR1v3jaVLjXlyd5cf0XwttVrCtMTfn7L7UKHZ0mu1rZo74EOASnMsFfA46c8fkfFNM0hwa+
IkkKQwL7/Hn/M7Zkkpq7pSJY/fmtwK8Ao5AzKbZDULt1D7mM12hcW08aP/Cf/S/e0IklA+TkVSvt
kTBO1GjTo6i1kxSIoPHs4M6i5Ii6WYQdmftYb0XHw573AnOMU0svFx5ivw5aKiJmrzDTt7JCk4zD
6Hxm9+Ypy2tbgmCNTJdrjtnb9wcHPWui37MpKVRmVY/Elio/X9FOzKgLEGVOrsIFV70K12z/vxqz
KoD/8GwMTkBHjl+gHrIC3F3ZLpO6jiadmqWtsaxz9n1Zwl9SBof+H1Eo7u1sHa4CPW69waW8JHW7
AiQ9St19fCgIlT3ek0UozIQWlENWgdw0xU1a49F/vcDryv3H3lbAj3vswUaqNwwAzem05SejfDyl
GYPb2t8dta20WtG19HoPw2ozFWps76cU+nHftfxjuK44/C1e+9rDPYLWER8w4PNA8Rcx/surd4JF
p+UBGvQrsGc0FZtlHEnML5K45nk8WJifl1TOjXaXGj5iVi6E2f6SvPk3EBBeeOVhIzch22kL/s5a
juwjYCUjwXi3S/1lJNSoEvTrXXG+P7lrZHLTd3sQJztw/jm2xGzSFmaVfSi0BmG0ulxJcjWHz/Hz
YY8W5W2J8jYY5DZPXw0C/vNmb1rk7P5jZmt3rnafJjd/rGP78vfkq6eY3jTEhT1PzXhFeMN4ceCY
xAS2eZInowrSB31qykg3YBiWYEkiWP+Caygu4glH9WEOiRK0B9uDg6sVF0bIaMDLLFi507MJPOU3
fzaYTkaPWH7FxCiu5rvok0AtUEtPY5VeXAgd6BI9+oQkCAqVt6Bgpc2VdSH+YnlkbW0TspXUi5qw
eQodigt8dBWybVaByFz2+LP60KWNQpUPlL29BiuiG8eRMtDmbagmx3BACXmdjBHxn6Cki85K9KGd
LLke1QkPx+egKW9VVSdvqkwWjaqLLoZecffnkaDLBjG9tmXKEtZ4OSMHf0/nDEuFSnZ/pB+/w54v
dM2eZl2+qIXcPVDhUh1cRCoyoajSG9uu0m51LSIHy3kuxP8OmwhDSk2+Fbh4Zhj8MGANuN43IHD7
E9EZsv58LZfhiYlC9WKmKtVXmEIBFt9miUTy+mWdY/EY9uJ0T27121aHgsQMO1R3eUoR7wDY3RtP
UXZpKarjGBNBebvAyDHlXDwPhBXbX8bi2FCkWf4O6GpWUYrR90YGXl4KaOz7ClMtsSSKZXK9m01O
JPa8ytE67uZ+UsXPX+Yuk5vfbJVMFlvZvKf7B4nj4Ugvbld+eWZ+PrTWWfzLYoFlvC/4ftWu1mdx
IMs+rrjlk+Fakngo8g2298ppCJvZxyavpAylSkw8Ksk6wGBq/HocX+bgOYAxSaU14MfPh9Y+em1t
0+s3r3nMOx5VbdCXjxyXvcKQa4Zrvr3j6DmkcyUYcHfUHbxjOdOdKC5TXN1+EBgEargISqOuZyOO
LO86jWJoPSHLjZ99teasQiXqOPoHKORQvRGJ/w0Jgnrc/7DtNiWFC5P/oQuy1HbYGUYR+k2TQp8H
jybjmZAf34hhg0NiqONiqxElK0aI5diBOPhH5x5AQilqSCu1XRrkuP+wigWCffUm8hIZcIQX43Qa
FP9KSjeXlYuYul4/TIunudaG0lmwhz+zyaP5ml/eV/PxI+cJTYP3tfNPtBGuEdPPog6IBGrcm71q
Q3lOVHZSqDPrf2Gwm2HCeoB+roLW31xdSaBXY/sLhb23djHo0Xahkd/AxqXlJAn6//fkfQPLRtP+
F6UplkLsCsAg3BlLCWa+QrsbgK8B6qO7FupuWtLtRMBZ7i2P6hyfogj1fmJG6ub7ReUXN8+8SaRJ
htuamuVoYamf2nNo44SR1OmaaKCNSWmGS96SYfL3qhZXTXRIFuBb9nnI8nMs+DJazlTjtgDjF8Gg
QnepI0HQK7efNkeKYyU8fxj82Z3FuBA7g+QAwjw/AfYg9+g174l+3wm98j73u2Hj7sCKnDSGy7CH
tST3zlokZ4FhU5BRbyKdcM2XYz09eQQL4QUd6n0kLlUZsPXqSzpa4LNq2E7QXUYgyiDom49927qJ
Tdy9OR5omTVsIY7EZJCymhMht5gUJSrlGoNzX9sQX6pGL3X/GgjPraEt62qOCLqmBybdZiieKhdw
Njq9YjWCPfdz+M2bEpUoP7zYvhmBvqWRRFmAtl/gvihEGPsPYeU3oqqewc45167R7otD4BszS35E
kDo0fXCFlL5U3UMDOxK6XqUFLUIcz+46/yxsDP4xyPFLEX0c63/nOp9WqvBDstcj+ralfFRavOab
KgjyMn5wfrBtPyPOHEB4APku5+gzHFXvojh3x4tAVxtQXY7dVIrlmtWMjydvSrIpHq529xKh83F2
Sed/tfZpwAN6u3ZUm97SNrQLwIeRSLT2RnVLRWyTHgbhFbnhC1hGfTQ3+f99LfPNpGbA9kqBNoGn
lxWaVfw895u1NvDfhCiUucrVkHfMCQSIJs0QECUByOq/zUzzGLKPlCJe4yRpk8SgGcM//h+ykK1a
nd8ijHZHlhch7g2bKlLcY1e5J++ePJTrWsh9M+qAFSNPJfNOBaaSywylEckxmftY9tq0oj+pEFeR
5svXgy1k3VTpcmf1SUkaxiQE89SAG4hol8F195EFRVqU6T5hWtP2RFhcnW7VmFAmpfQq8AK48pdM
a393eyvbpukwPoSO2IEqOAQbaJl5ZQwu/qdeN5CyThrvB+f92RxzkG+p0XNnVXB1JatLcl+SnsyK
vIX2V6OmEH/HSFen1OZBvEyo7P0hyyW4vC/+vJtbiu9cIsDceDBuGq1bX3nSQ+7VqA9SYnQAciug
kjjv/g6wslvqCLrbIhwY/OMg7Np9u/zPXF0PgVL9+QVoZ4IxuJqWJ33tAuaZxoywHliyfjLzfzho
cYLJ8RHNHA7iSnPtxQzxKLmCgJ5e3oepkwCTTYzR3ODEkX+70UE1PCzPNbPaZwAHYuaLUQtu+Eq1
lxpsdZUYR5cP8uKtl7vsi4Vlz49h2jVaUCtuFmeDnkt7WezAD5qRNmNqL3L07yImVGiWA2KeBl/N
UAu7yWIBb4K3fk9PdmyFEOHEHysyOzsSr2udSWvADh1AspAx/rSorba7ErbcA3r7T45gbyF9e/i8
zFGVXi27oAqAmOzRAo+RxrRODvj0nXp+H0LMtQyvT41cvwhbeGrwBAan019yq3NcbXNShlD0dMia
ArHnnBjXHf8Y3m1MQIokIX+WQQdXCTyk9tWVIbduuaxS6WWaZGAiML/qwxJDxbC0QWvUrbKKzSh3
pdCIb/AW5GNhFrkpAH0USXJZKhha2vruZBWzowHbYe4Qt2muCAPCESA9pr1fwBvgifiugoKiSuKg
uNeA0wQY2Wnu76YI4qiKovsPGWHqfCYz1cWbDcCXYUYrtrOhCnCgtA/eGjIJfeupPtJUpUsrDIK8
j5CIObc67SqLlN7Xk+5/gKUrzGcUTVvcXx3+2kTCSdsfVln52m4l07po4Nl2ua6Xx+pt0HARu2Xy
leEt8dzXumqzLQssVKnFS9JG/PEN9DGvdq/nSS8scp7HFGOYTyJgAbkd+898bkmHc9k5Bwhk3aiQ
gDF8MCSbF7ms4WhjSPC9AQvEvDxDEtc9zqi3JRsc6pGrT1y6EgDnscV+WO3qwciRisvK8Hg5/bO0
bKwj58iSNjSqzB05E748dttMayKJoni0oazu7edAIA8QfGB72R4svvRy1zkkAo5HIo5hzV4kWdTW
f8SV3O3Xt4Q5IVINIS5qO5Iw+tmzSJT/V9ziRq347cyUgFgz1Ue6ap7dGqhNIOXvzCpj0CefJu4u
vVmjxg3i6uO5pGK3LZ4B6OjNDAkgnxbk2nYBSSq6R2f3eQ4IbUpmhqbsaWoLgyg7rnh9kyneNogC
MVF2Yj7mxjYr4X68ygVsg7SXjpa/STPKUTejKe0Yg4kTqRnTaJ4qjETQnCr2J72Wi/6+IJX/VGZF
NKM5j4OtNu63E+fX9ZhaNEeBVgr5U1poCrzNmMm/z5an8njLudD82kwxiM5rhnjkqfD3xR8pz86E
PPg9NMQ1ZDGOOZ5RpAY5ZZ/SuYXvgwMEPJM/vK1/PM9OwNkWcVmx5Hhd+Mw4IrwvcL7R3dr4iRaF
JbvAOws15VdRyeYIrWyLtdpaPGB/u+aXOHaIWQMF8zft+X3yy+p5bDw4Wmp1qoWLsfJ2hgXkm9G9
zHnzajkNu/I+sH68TBY/AA13ig8PHTIfV9gWF4J5jXCzT7bvUzHNg6KaZeNRDwuf6Hzhm1TbT2H1
hOfA3q9X13k7ffr6ramOwS7ASOnL9Xe7xRBOSzIk4g9EGAcEgvCGylJ2FsMH21Nb9UGA5ItCKIXe
dtbJlr1qL3sv42YslRkwrVTbhRcUuC8j8Ti6m8+P5qwABSlaqGfM222GM/xBshliM2KeVoZ/h3EA
M/HkbRhIplGsmsaFAqk2G3jk+bNmoHxb06hfY3YQelX6BbOzmpB9GR9nH37Ku6Z9SCm7kPrsMchT
JYs/GWbkKnmgnM3qwE6BtcBcREjEo4RlLa7QqTQrgRgWJi2UNznevW0MiKuFS1CG19eqIJJkB0AU
C6eK8VuP5xFoWx7iTrX6jQOTqEwY9CXD2Xq7m3NrtkDvIUt6U1COnxSqkLnyClfrC+2iLKWTBNa9
g7ir67PbGQP0Lb7Unwq/csJM/abcp4Wm66cLspdMNW6nYxoVdnU7Ap5tyMCl7WcE73tAbNY4umNT
kMN3JIAziThYeIzpOCK2hlEI+ncGJDOxzDjbWFqu5VLqI6InLG7ikmkqWGxHgJqyPLTG5fGucqTI
4RVXpX+cQK21LRWMBKki8W9+Z/Ets2CCEhfElJbEj1vXtT2lzJtnYJ/ZOAzO2a1cgkpHcV5dVSs7
nk4GUOYAD8qtbX4i/nmuil6ilqUlVNRJTlbJFjPuYULkXS6rzR2WfAdzmTsf+GZII5OJoMgxk6Ov
p6BpOZ6UaYCC+/VeVj+Mg4dpxIRjdT0ZgyaP+LHxpcWGhdpSmjf9n1isNvbdcN+7Wun8Ok0enBgw
Womx5uL3S5S0IQdACwdakkthYOpKWx6PmDmwG+XjfrG7xX/c/S+fXKnzwf7635Go7fudBm/jsVe0
FB1C4gncwb9I44qFjMp2GypwSddjZj4fZ3kh1+SH3jHuzM+YSC2h3DYN9uzYvPNp3zjldcIH4wSB
Nb3DvAH+KDpvRSjgmtqmgBAUYJpd2tIP9m9pXONoiWwWKxzopqjCLSq+zDVBn0SquByQeGM7rVpL
LZ28IzPTQ1dkPtDYACgRAItsS2yUK6sNCTb87klArHuYic/7cYLUMbyeiGJwT2Yn+17AGYk8WkIO
Up81ztE0uKeky35mTZAK1UMI1TRoqTKbZ6xjEMxoij3E/UQJQGiYCxSj+aBlhNbIMDEAAgZDOZHu
+W8Ak+3+07eafMRfbUgEewAUKyoArXS649K+KrN3CUKZTmb4TDPNDFQrRveU2/FgXDCABVB8ovEs
IS8shzBE/D5nPrFzlBwYyiyr8alB54ncQiv66uQcBGZiPBjVADPE4GCNnn5Vqt/u1X+LDmeG9DbA
ouG7ruDqL9h3qLDJAaSwiC6+FuW2Zsi7VgkB7xMfh1PVHCEVW8Wfl4ghBZcJoVPV+/GcWYLxISWM
vdvJlv0y/CYRPVCkyIecyeCmWDAOhAjwuFdvJX+n5JjcZDJeyBG46RP9cL3dh4DSCudefvVD2uqr
0lho7y6iHydSsfm6T+GOR7kwZfYgNUL9zk88t1b+bC7DIkAnLQSjJ8IexspgyswLMVF0yMuVAj6g
578Pn4lYsaTXAYBJnnXR3rGh29X0dIB21X5FaigBuT4JqgfSNVrULMqO9FoWVnIMQLYYjWDGYflz
p3UGBksUl8MNI37HCHj2a0zI8f7GdEfhPwpCQfL6VKYRSBvvHUB8IUyjZs19C6lTwPn7Kvd+byC3
poHmgENqcmuGtGdGEjUNKd9sQi0HUGGVUOpsK5i73muNJn41Nm+xB2aYB1G94L2sANIzqgmrw2mZ
5QTm7P8+eS26W8dw4VsMUGa/hgO+e1iMmqylfuiEZhfoGqRRKurn3fP2gD68H4CfwnGzCwuB8wiv
tEehaP0+E64K3hro90OYBDJWo2Fw6SfOiuoy0wR/9pVQnM6gfWcNrmqzER/BMO+R1RWgAwjgc/rV
VQJX/+nTXJdr8rzZ4va1PRgkDyxhrbFc7zHDXiERqpb1gTa8NZN+a6zw+AuMhk+HNm/9/wYjmvEa
jBuZNMAXj14hQXNqvCm/GVxF0I+T0Q5eHEmC9xYqjzE4CMMnQ+SuL0rfZbqjDW7748k6X2QP9EpG
xYBRZZ57+sDQhg6wd6p+BvSrRLnUKbHNMsNd0/hRVHI8McaMoJlSkf5C5Yav34pyo4mT9Ma+IIY/
YmzIua9yD6h8y1IafKLmAsA5yiXXQ4zZrpqnN2ROS6j3y6vwU2LQPkhz117fZG2ONcYgdaKDviCc
C8eKjln+ODVEY34dn7jaUGRZtBhR3ljijqynGe2IOO8SWSFY3OnQaIWqoCctnUParBxwJ8mp/6So
f3rMNWypVMNUL/bdkYOqn8M7alFy5FUTqU5BJTbd5SGBvNYruNsmwdhnqrgjzZCHY2A8q/K9vqcZ
uRH0WM0iwVY105yhC3DwZ2/nFtEI/WnxIAnxFSaKCuUZXv3RZ2vAlDHjtaT9ej06oV+nvRrRij7u
wLKn3Ceeyukgg6AB6Khjl9eoJrYZMBV3LHOG5vJLY+k/HvPF1Bp2+zFReNdDDdYXSH2K+1unZxLW
bx/syT87gNi/KUIUTvM73p+BEA5UL1ZXqQ57ENY16o47cKNaklwVxzXkN+wi0ZkT0IUTuNUQHU5O
4VPlVcb5R53Ws/m8M0c88JHjwtARqzq1BhBGBbcowf4UyIdKijO3zzEOIZn763UId0hEd15Pbyk4
/c/xZtKQxfC2Bol9DL82VgSlm+C0BYAVdKyVHJ12STKKsIV0ZxRKZ8HTAJbzlcoM5ik25oJdDOd6
Ky1LhcQFyupRWHd9C3MePdufJl8/LhCIMBXk8AgcT2nulUJwBWdbcO6Y3ctiTI5aCLo9Ir/0mu+F
ASFmOQqR47Jw/5dnA4evI/5QAGtuVSQbAj250Fs8u8XsQyf9MQhZkIBG5YBckBWDUhNuW7KIB+uz
EA1okDRHV3fzEoX9wYnbcVBZvDxW/7ZdmapX7wgMMCF9ecEvNDN2PvuL+es0Fy9HDFbrqP/HZDYn
+6PwnLy7dLqRq+kc/UuALojZJq0BniBIWcGORUwr3aIdWtpNFOxXMq6VIyHZQlbDmWfg2Wz8qiTK
3Cmw/Xm3jDAgOPeZqGHIfJ7CDvra29NDzSMURljArn7fVuxoppUzgYsRR9zaZM0Pj0HF2n/yi4gj
p/Ifq0TbuUkuhttWlDUXwudpdMGCJkJDMPlKcRbLQhutykvSfCWKQAHPe77HCwPicBBlgwyyCouT
1EoNQYQKQsVO9wFzy8olTDaXZk8q/jz1oIMz6eEb0axu9R1gFPKgQ+U1S2BprNwcvv6H4MQzzRpZ
J+tilZRv3vujR4sjnzAnfgaBj/gIG4RCNxDt2xLxpzxoVURGlYcty4hG5dLtdpXWgESDKfDChmyT
swB6adZvGKWSKpu5D2Bd7qS0LC8lcWJhsVGjGxrAXQJamQSlxPHGqSQuQRdVqHQvRV/UTqmTvNgF
+IyHLsCYJ4s47E65hH9W/9quHTIcP7tGiqVgOt55FgIK3wpV6MRE5U8JYvmnFTcL0rvyejqpV50o
Qy+Lm8RKYrLsDReBnG+xV2r7LaP5pG+//wR2fThjNcWUsqJ05IeYi4upD6BW1+wF2gvz3PQmm6cx
pYaveXhMmqEgPAy6Vv+0P5R3NxOSNVv5r+0jTo8bnWT/HweebeG+El1Oq6pSD9Nad5smAW4Tn0VZ
9SdAXDRhQvGZjXBIgTpB5wtOIxIfGT8ysIRl9jeTjkD5k5hKwMQ+Qt3dG/0pSsrOocn5hQ6HNQBF
hK6nxAKIU4pXKqSCivLI5qxiyVOxQBwYptT+Y4a0hOKoXLTqEp542HkD30hycYKvlB8BEZHaqRmi
vPH4L/p1KbtDpmUTfOKBtSiREgqmOcakbiV/aH18vU3IzBxFKUp7uKoqYp69BL4kw2nPAamY/0M6
HVAniOxSMNROlkbuHc3reHiPzjCYFgQrr1KktTGCtT6vw40sXlkTBjg6VKTwMtDDDD5FIv47TYK+
2cZZ38nw34SHJwURr6RFVNFGl5tkIpj7GEUvCNyJaWdx4zjlqnu1CrMncmgpo97/WqWbQ5TeGGpf
rm1l1xg0MZJbbR0r5SD7tQS6jOpIxrrSgG/USJT1ycfsYEW55HRnJGQKAZNl7ebtdcxbGNjBvpXV
to0Q23bSHX79QtO1LtXWZQsoWTVnq8OHsQxl9KyUeIJAbdGU2y+/H0tBn00z9LGP/hAZLmJbPqvW
TDQGoC1M6VRvB7Pt559qInPREICxKjOaZ71W0ZX9Qds835+aCjDcw/CEAEqxReR6zpny2SuiNZtl
m27L1cCcFHCniskXwmEqwaS7fYM4INUgVCJojez4Qc4ZObKEtbFA1QkS+/5lVfCaD+Zo7yNwbg0C
hF0nhbErRMK4Fy9i56bpzb5DnNxojCMfDfVcS+C0hPNt1LXKsayjh7n3i4IOCRA2KYRgo7yJWsk0
vRGtmSi4DL83hNCMM2Vq3DmA0u1uB659RFBYfpT2hMyDDjPkGbt+hEIDhwBzMo8pBp1PDBZBaR9C
BZu9uIWcjIBGH62KFmwCssNKrhCESZ4UxPa1dvUN9Yc7Oac5mcSEYU5FyU4/0DtjrL6eV3wpyJ1I
HPrmKdJoaowlptHBX5aFvF4xo1SjMZoVFlmod5R2R2SagyWtX9yNN22r1/DBZacYWhuBC+NhtOxX
f+NpPuwqYYhdSCNUdkGDwNgM1infqPI9l1CuLbpqt9Jfnw7VX2ylUCbTTZkLcinzLlFKOdcq+7r4
5ULBD06c2ByneGbfg82UH0wnrYWPbjTBmMs6J7Cv9iW7fq74UJyeOE89ogf5qETz/8hUnmn0CsPU
lk759Qss26e4H4jDt5MQpDAaeWL2Qw/sQRlXgJFa20FM6sq8Q++cpRjcY0Aeg8pyu4PHk72oTIAu
Ofed09cdgql2u+B4VPyk+RC8qGeFsapk2NACP4vw5cETCKJRYlyn3eFiMOe1L2fNCHAuDKf59D7X
A+kvROcrJKaSYLS2+NzYri0hC/a1R1TXKHDDTThxKRIM1e6xPFpf9AiSCqyDFelbuSXPceU+YsY+
76TwJFzGdoeMTXbt8Nh5ht9UsAKpFbkgm1Zru5zvgCZKRkC1xC/BdnYp5WlqfEzcPwUADbFyZfjq
+8CwEznaOeWuK01YlzUqkWus8e/WlDh5C3g8zT7dFubDSAuVwoZxk5g6DPCUWvyg8vNW4MDUNOit
rlZj0eroQSoDZoCj1kISqXqAGBgihnDJpbx2yC1TPR8QYiWlbv59gA0yqFa5cOBe5pMBaV4FmFOW
WVFv+Q73kRYD+hb+edoLB4tsOm69TvC0kSfHikRBTHaIJlohGXa6NnOH5AChKsNc8/UnUFYoBvaT
WlcF1km212A96JpUYmKSbp0jhU89mWf/iYdxMXzJ9d8VOKxpcguEzraFv6CdDbxH94MmFNhk7A7h
UFCmkhN2lKnnrIT1Z6Cq0sJXTlktvNAUdfVBeftS8eGRyehL6fP2dpKQLkADWtGJOociesf44t8T
v5p0Z81U/t0mrZzLeIvxW+tsPtZt7MHD4QGROLLQW78CpZ7nr21JBlVaZVPG6NQDko54VfDPnBDn
niwnIH6wqwsKA6ucHyd445ZL+c3IpcnyL3OGYTZ1Ht/fuAq01i+tbWCtbrvNyMOnO4mqjZO/+uTL
6xIaD8wq0HgK6sOLHtkut8uYCFdRvvh6nfV+cGFJq66Rcr+nzveX1OCxgvASshWHMGEO/3jqm0sB
+idTudCzNGiUwY3mdy2d5pPiwIP/lPiYstMuX4zJ5Jx3lGDUBs46N8VMRu/I31LOpGP5jTZmY4nc
Ms97xpkkMJXIDMDW9EXx63sl89yNxulBGBRL/OgxekVDsCwPhIEOOPw35aCOzvmkwzq6GS4aJ4KO
0WBNiHAGEoNfAveMxhOLp+7e57USmTJ4fEC9WZnVN3TcgiPgS6IfEXIzMtjDU6kFJNlTevV41kiP
x1IJ8FM8vlqKiDv0NN7bKv8sG3TIVvJu6rY6/TsvCZPp4n0EO46tZ/k/3/BteV5OZKNC2TXPRYqK
QB81P37xIKu8+5rnu3Pucexm7k480TpVYXQtlj+Igmkznr6JPpkTM9wBeBDGqn26RaD9zqxoNFhI
W0Qg7sdtEldZbCOpErTZmjf/54oVF3BGgSHb7BDf+EG2hKrV0LRyI9UyDxVyZLS9q7EtUWORso9D
qb3choCSoxSjWpikjq9bjpydBKUI4b/NPAFvvRZBUkzLkF1VRHbJKiU+Q8g4mjrqUk+7baAo68q1
0dAQ+T5X8lq1Z+O9EG9szyKxMDG4v3bWxjI6d3TH5y3ffpKUOvXjXcfvw0m35LFDte1O0y17LZgW
DTVwE6h2Mjrz8cxiG1vx5J8yngMMONR6b+HMm8yT9nVK+EjPSzgMyaIcncQXlWLGlJsv0pFa68z2
U5NBzh/0H+DIx02buQeaE1sxF6grm5oxd319w4Ea7dsl01uqyyhrvyV92TJa17PAPD85diP548Gs
3ZQavE5pLLhXXTiZLVIyeKK9/URI2edx3ZnuiSHJfowzYcS6Fgl8naC8g6iXiVT0Inl/l7mEu0WK
w6sBYxd5usnfiz0T3IhUD1QLZMA6sp/on6BQtwHKkDKrljHO4v8+BM6NAu02i9qTe0GJbpJqoF8d
sVcYIa66gGqd0/hiPbJHHhiBReYMuQADG+zAERRVP92I9wQVD4fnxyBgnTruRwIAELyCUmJVj7PW
P8qz8uK5i0rZpoI/GQxAcUr9uAGXulrnTJh2c5tThfvFRRQx8ZrudQskwxl4OHXUXX5wH07SkKJk
lMVkt+31Eiu2NEChd/wbVOb2am2+GcjdROAt/s5QFkapgbB2w8iEwLzu+epgpiPGk/CEojWBhyMZ
qrE9ncs10pOmWhfq2nmWQhc8C93uC7xRWauhg6azfin+spZ4e1l4AP9aACvPS8NYXPoaGlCfyTKh
SGXVLedkgIeHD+Dmse/QJ3jgpD6h2L2jpV1PMNlBqdOQKTYo4RAyfFPb0PyzacKqCWWdNxoCSnd1
fiA+LGwcMsfczyViVstdce70fwlhTqfYMcNawRqfs5M2U+WR4E/iJVUf4ipAVu6YOwLexfW4ysVO
h+1dCVeT22Ck5nBwwEcYZOInqEDbloRqbdzeOBjygdway0cPsfCtHaUfnSAXneTzYzvx9IvZPDKa
B1dpX8TARNQCNDJBauxjzrvR0WrTDD/0ZjI/6znLCAqWp/KMT0OxjiiVIU+dt3UA8dzWQrxdlviz
EdKNCMsDUWXojyEN6jMQ5NCjvHLe4PLvW6tpcczqBIiNg1XNTkBrqbaL4UsBGnbhVuDlL0AW8Qo/
9gKOQgiKlD45AHWm/lRuMxhQJsYuFKQNQhA91V+xfCot5MI3HJnINBDiKUNDArgBvk2qextUEV8E
gQ19tl3v2IyP2xNacpOcnWM6LoT+r1TSrNgxLDy8vz1Mqp6Xyjr7WVd8aO7TxBb+zy3CpJKlw3pQ
zsDmVbNEP+2X3OsBi9yhpdp1Hn6lRbYEh1Z9eHPDIePt4/mDQnTyLtL+lBYu7GJCPsDNz7uAHnr5
yxgPyzqWFwfan36vggYSt1x75OQGZaqfrC8dlhcUUoTuEaOcQOobttmOs36UP2jkKjf5XppqWVJz
of/QKtJC5RpMLsxtavFU29csHp4mOI1HsLlLVkqqD3bAbeuaQBxq5ksyOeeFK7aIj0b9hk61Tn+O
5n1+Hiu73SVuqM5yux17XATP9yheTgZL46noErjtj2NtaduZMjfz0QN94IRzb/Ezms5MJA11Ncy9
p7cqX3aBnsu266BCjfzoDYJlO5V/Pu7UDvfzzgBN0WfQJwCazCq4vqqArKeYxDnMBS4MZIZ3vtF6
Smt2e4C1a7UgU1e59/CtGQxmaMX7Y4n9+qv5m4kd9+EeUs6RyNc+H8bnq1UFu4w57IPmnFwuj/zL
/k+955DcDMzsoZI+szQUinNnX92VQE8lCrRkqCqZxiiQjG9ZNybr3l0F32hb3+5fDfiGgPmzaEpg
HW9IBDALfmqW1hSdotfnY4L5+ITY80auVddiS1OFUysGVuC/zftGtGrMMuqXxBgpZHvCSbCuqxgf
npYSSlkN8pTxak9NKQK8n0/xvhNPJho+6Uact9d35xlT/JD3Tz/NwlrwIhXaUeYRzCj2QIqUf7BO
Nz6Ot0ufWMprKhKtsyAtA4OtYslqtl2Y5iHi3J5R0tMpBbDHyR3c7k61/uVAPML2xk5uy3mNUMPT
Hu/8Wnh0vQpRfQgsZhNs3YaTCbTpFkS9ce2aect4KgpR8JW2rqsbRjiCxEQbI/DVt0Jg/FM/wiHt
zDPpfLlRJ/UXK1IOoHg8KNlFGCRijtADmvTyzAXdOGVsXezT2/1FvjFg4JnJFmaS4pBkTbhvbrg0
lWb20dDr3tlfNHScA77lTCyX5VxpcaH/w4PK9ozrNkzlboW/YW9XCaWjEG1muuJz9Alk5B473mJW
t2f7knDcWTHR3uxj+pUyLC5Fu5d8OjZ6jhy8Nrv9DxAmNvZjn0M2Vdk78YeJV70q4HeXrZNGiOYa
BVglvuYYRu9okR56IoTAsVBYqa8JRY1F3zw9l7jPgvE0eblFt3UjVV1hhfJyungciw9i9EmRN4Wg
2U2+b2x7AdMvzcFDvMfYwrXLejwhXbr34/aS9Lm4NwP9RygZ6SRlJqNIJIs5vUaRrYDBrRNdN8pZ
Yp0jL9+593Vt1R/AXEfnc2HLCG+t76zzIDERAqaeh1JbOQzOoIc62EhBmDOKo/HojSF96jFlZzvj
cTzfzGLsbtAmFsirKnJfst3HFfCTaj1JwWYVMIOL59dqiQNuW+6lGBKZFGoV4yVypjhqbf5ZfOmx
E/KdBE80pOK5H7D63STG9L7jGpsfcL70WGw2SsLo5ZBetUUvaSbTRW3OU0Y2c4HfanP4rnKFMgLt
KviyELxqaSeXqagXL0gR1qjSbyNMyzWiC3amtO6ubYFe16YUF1OQMA2Uqo37NxduIhHwKNZ9hEEs
CsOssplV62I8HCR7W+nEXH1UXaIV+XDWlbvCffAl5LtWRoexoIGEigDOCqOFndbqUJr6ky8tVUV/
KCEdcK1k6ZtgR8527apJgLWuapyuB8KbaqKJrgBa5BE8Dm5H/zOU2cwQJHJOzFc2qgyqIBe3XQ3V
XnakVLiZVJjOqgKoTrrRHoTxoSoDllikgw1aLoh+K7heZVnXOe4CMUmj7nAzM8GIl8SU5cioXiDP
zG71JZ9cLKri1SBdfc29xbQVzX3rgbtwuHrwWIXv9ClLKOoHeRIZH/6ssFv/AVsikgYQKZ0zqA3E
7dCWenQg9kAaUHEZYSY/Qf8+XNLHe4n++OYNXLvVVyY8tdz/fTIxNJ3pRuSg9ccteaerX371d3X8
MaNUvH3+MS6WGE9Is9tGZNF5eYc5zB17Yw13vNaIDIhs2NMFelxaDAiBij5dULY5JPC79i+TinRu
rOGXcKPj+t0r/SUMIWNrmmDFhvOHdpmjpxcg2ds4A8Q2jIZrVHNUEVXDK6hMYQKi5avsUqyFLPMC
R+6EAgvtYfLSoBX8EdL7n+FGpThKDDtYvfGrD3TvgM87HfY/zi8TbCOTdN0Vy/ayl8Qpo6Zuk29j
OGbDiFsugicIA+AhjCly/5aGUfstnXGryww28AabZSampSFBI4k7nZXeVjSkwha6dAYyg1aCJPYB
rn1Pzl06BGJeGIiIaW86dh79eIOm1cIanuv7h9SIWsLHMJvVSKKfDofr7LRqo8/yyMMSqZVD/FaB
t/i8KHnceGVVCX6CI/BlVLt/3eAE72hUB+bAcvziVwldwLVyLqIdsS3ikjhfEX5G5SvTJBsyEpea
MwK2eNGKaJAXcRGOjHmzbRmxutr8MNatQZEQlAjgHzJV2XndI9kQRA9GZTUU7Jwh8igZkmyR0s9U
N7O9h9Dof+SNwmlGq9b9ZHDx3bnje/wJ0jPI5/eAfSz76+SWROUmtnI6Zpp9VLy+6Pd1jtOwS+QP
9mS+14odgtQnGkeKl+INXQq8iQvmuCGEDyoHBr9m+RgAE3GXRdx0KdOYXfIKdRoYvMOGWAUkqQY1
H12AjbO5W/LHfSacxydRK/660Ng0pcUNdb0VBqhSSMuI2BzrNPSf4Mk/j1P7a9+U+IRNh2pmAAo/
pRlt9kBbTYnsDwObxVb4WKx72zJxNtULRKUWEtclfdk5nFLNd/eq9iTzQofLAyN8yFyQZIHngZZ9
OdjRhW3uuHG2ZkCVQEnEvzQnO5M16uCG8MncFWFdzjySsOjjByP0yEnSLd8Hr6frk8pIcTx8Lq5K
eLuo8qyIicSrAU3c7FXe2mpPWyTw151bFhzUI/U/Hj1y8dk1zliLZX/WRYaMvaYSH6DP1SkC4bd/
PrWsXfntoKBU1d7qYXdaOo97JS4CKv6rRUhPNMyyMsgCOUYubtWFGNMbyqEw2ghzTZK1P2LXKRaP
wGPi/3uR9e5QzxMXO42tdhl3Ds+azBOhacVenp9SvSIJFTmG7LjhWhyjkIaNhGayWO9e9fO0hk0o
oxN/4tAH3gN2vjUItvYwZ3aNVoI0jXWvtih4nqWxsQC4S7FFuhRflcK+Cs5gFkDvsDJecCIC2XLd
rOBbt/UHXpRiGCSrcCiyLTma+Hrcnj8F+IrGC5Em6f9pHbX39hcx9OTg3KvyEvPkyp+b1CD8VToj
eb+H/NWAjLc85FPffLKNrExcPxrOtQZhIGlft5GQfeJu9xRM7oKqqXA0VhLPSEzZp2ziNEs9SFBb
/Jj+8J3kfjYBDbM5hFPDQiFEb7pE7hymyF5ykTBNtcdvfQUIcGBHF6+qK2T1SZTAGDvdBTnvk/Yb
nWW+Jtv6xK1tVvQCqy8awzcn15fcnExAwBlT8ftgrTeBjQhyszrE62gF8wvf8E5vSwKY6YmP/Uex
RbXhizYhUtO8mASGvZ/MJKK3tW9wlkWQBcHz9xJhshoNUVi2ik84yTyTHyBk/tRGvbD2K075V5ei
TvyxUnbfwmUxk7zxcYE8wNxG3upy+yuVWRSjGWb19pz6ykgO2cqQpF6aRCsZYsWgPbN3YLhYWh63
mh7POn/U2l3TSVZiXSzr42TjDRhL/sjxMUcUbfKp31PDdWRO+xyVUyw6VKh3d2rMsCZvp5mFiGYg
wuraVvyNrSIbeZ0hd4rxwhcr9Pt3OPmgxqloiJkEFpXHpTG8ooo1/k4jrUquYvKoP8hcQn1YWOhc
vbrFQyVHvQGJ87U+76CLN5HUBpYjPRKy7Qy2+BO9vsH2XILVs7q+EPMXfJsWZXKDMw1yrXAMrpnX
rSk1prdxbV/VIDiflzIP7ZciBR757me6ArTCvsWeoppEDNwjqq31vGY61v4iVwpkUBFQc4X336o5
bq04Tix+x3ekqIXeU/55tDmGQNCPn+uvRg74/rvo9j5bgFa1QYZz0b/oF0kWV4TXFWM+8l87i4Ks
FxLWK9fsI/qqFY2689B+b1QPpB4M49OyPNese7VnHTIpzuvo+OM4rnDxojfBzCuoxtIXvljH+Y8l
4eB7ljNTDdryEaK1gf7QmLiXEzj6lca+KuHgldodFGeSJsSoSOLSrV0k+QBNZe17Wg26RJdVg+SD
GkHruTKj0MVB85RYz7isjRcdb/EiFRC692aRqeRLahA8g2wBAD1VoSH/HYKUWWepEDCV0oVJRcU1
b9bxkhEJfM/hwsVE9Yx3V4V3WcQ4kW898ClBi15ZfccoPU+T3fEaCaLFTNoiSM9ep2nZpqjSaTom
cPNdOs8pF7RquPRC6IR6w2eTYVzg43ceZAgQbFrmcdMuGabgm9zpfpX217yr/bFpVYHbTPYiLSs1
fkmLIPEqLOTXGREpYLuUb8ELMQ1yrqYA8v9TGrTCEXpzfX2dhLcuN86bJfHTAbPPpipHTYyFL6ja
WTDBBA40GqQynsgP4pb8EKEJaPffj0wmTLm7jUufaaTWdLxjawgI7Ld1iRbMNheS+b9G+3ZAFKlF
FEETaRRcFaUugRE+jc0sXvNfxCckiNls5BA3PyRVBA3VUqBUMcWpm2lSN/nLxRkYpF1JuzUEUaL0
LTS56W2XAmzAyQUBgZ0GIxr5CKdNuHTLYlh97PsjFkbDf7hTjJU+m7ZXRxSxr1rgEIy7CfSyNAKY
uCj3WuLKg4Uq4JoGuBrUNYRT6i56qJ5nshS0W0+6Ez/O5JmEmxiUGBNYE3sMz+xLYV7gpPnpIMiP
ucLNdqOgeznmCH9i3YaSZ1aBoJdeVNS0UYb/DaY0N3sa0AV5QVr5DQ+pQqhvWysThbpHZQaFbZQf
556uYAmoBcL3iPbqoEKsjRB7IehCCCZhVJRlRocjsqXrLckkOaXc/IOVZS5fzTWpNCL+HeZKCLto
xjyr8wabeRrvY1E8kqMQwzzMV7dZasx6zt3e1e+e9169apkew7r0J22a9TLdn1l1F+PZYLJfpS+4
XDoo239fBECEOdyoVoBvIf8KGVJQqz0/ktxlPR0zw93SHXb52nsbzQMF/0dlzNWBaR7/gbZhN9lE
3dYqHtXzy1sUt6GxgO58aCZ3fiSbJf3218qXoA7/nK2bKWxNYHFA/WQyb+sMSPu0mbUP6DbkCu3T
/9yhfVwnqLPBIFolCsvwdn2lArvqW3JtXUcmPiKveZqiY3jl/G3O1NLxbMGqYJxHYBQsyPEhXln3
lKyLQLDgiQuIPpftrUTNx4va59lwkkjNjcOnFBtCs/+bpbtAOBfnHsyQXuiL7rlt5HdLGGUWYQx4
WArCVJ9T5K5CFFAyW+o4wuJAnxNhLK3U57z3DfN9be24zZCpq/xFIyfhnWnbJkm1YxN6crdAP1mN
pglij5h6icQK0xNQAXqHlGOMCqJMVemmvINlVCzFUsIuSmMsORBeZjcXgghxb9cc/PxCSwLMP3mI
8TgTLhI8jzwQ/SPSrzbpHrH5MWLzYPoIwFkkZ1w1CBn8p5KXpmexY82xqqZxT8snqxi//lZEeHGh
ZsEk3bsgpOtlhgnH+rptCGM1kQWlRkKAmFnlNLz2Zhj37HwE4GIqbtP0lbOLKpPJ520T7Byl0DwE
rwIiEUc2g4wyZTsFR3AMsEqlSXz6RFII8WJiB1Cj857s9j5x6d+fnxZdfXOCD/qOUzi+uQpg/+r+
GyNYWKHUKQIDVsWWm050eUQJbGHePXf/+uV6QkA1876GWhtkQUp4l4ibOSOK2BzChrTZQYCI3/dn
zIrLjEGwMxWBykdAvbeqdolXo8f159iaDLEv3bDaXmpehObnbCOziVj5qbgXbsbC32ZXT92OrnSM
GX/1RZxcgqyA6mCXqt3mST2F09WrVMsO1KidkPE95Q2GvFWrcd1qtrAufELDA7RIFrwAprsaQ+AR
sktIMQOd5ml4t+3lT4dMsqnlGp3WY6AMsxn2WTPnV2ySosslNvg2QSEmurOY8IkjHmlng20kGIfF
KxSyxC09s/mKzitsfY2BparGW/7Cjxz/9UxoGr0SMEBRACwT8e7iAr8tetcwB86m6j6UKxrSyJLg
BDcX61xeg3MZd2ntebL9PYYFYC7nnStt3Sr/I8Ee18P1SU2KMaUspeyd2ddTqHacGm56w8abXict
6YebqjnrbNZjy4gEIb6IfxyeNPt6sRloUayq+3TLDs8HB8Q+OBZ+xqX0h+zYX0emNntF/fJ81ncA
rDpQCFFNueY9eQAy44fYxEymr5ggZMTkiqC2R9HlnNT/wX+HyYZB7zf8tgENmRPIn1u7ChhiVahI
la3hp3A3DudzBZB7Khkc/yLyH7Wz1R4kh76zL1JUWpa024T31ruvZUvrmxt4UuUxAhJJgt56e1BO
Ejax8CnUqjiP+5t7SqoreYhATr/5TCX4XU/7gGGQtjgDuQ2S0D6j/IF5yLrYLnV+x8rkefo0wIKA
0AkQa79gs1z11ZG/z8ZM03jvt3ZEaM9wJmSybhaAf0xN5zcJJE+HJjG67svKNwJWahQWK38OCOA3
+pCPpCHNLNK6/6KkZ1Vljluv7M1hLz6K4WrpDSYzOcjXZrCr4g32ny/kUXiw7eqbk7Enid/ql272
2KlZmwcn7b0nDLzXYas87iOStooVe3ynPEOJi+AyuTsVW/LIn6ZJGeuj4olCNfM9l8Q+NKELs2g5
mN/nkQKmHw52uQlRC9Bsvciz8OVyPwE/wRTW51jClGSGjG/sXSRuZi/kN/efddUI7DET1pAZkz2d
H/QJt3m1LZCZvS/zntX88o+ITRK+JdR3nTZILgF7YiFlIif0usjflkWgFbkqHPay+616QMZc1vij
BhQJiU/JuPT8vsb1dpYIGwLBFwAaPdxxHvKpSW+BC/8Sh/uQOgwoObeE5c01aWvLc7BUcXBBJv2b
2f1g7+fpP/oHUuIQueH4HaMa5oNHRWr8QbkVbkmNB2TsbfqN83+DhAYWdBciLffKacDAQEMDhnho
daMdE8jisvOdzY+Zg+JVYALR3e5COgqH78rePhMGRS3r8YabpL306Uk+2eETreDdW3TEMO6Xk4GG
Fwx38iRbFWTsXIsfzNT5ipGH5ZjmjmEk5Ne/3YSAWeAz9G+rjBJNrfnu4nJKr0slLm214+LlHpkH
pWLfJ0w9oUIlM2apEPR6jlQXcfD8pSDqzuAwVEVHkO6wONbk7xK7+v2amCHblELZzC26yZaU70ew
NIaqpHOQGSrlP9MUFB8/3gssL+zqPqVkUBEVcURFiFsj2+Z58Z2rh9tm/Ja/sAJqzMQqSD12V0ra
llik5DdE1vgVMidu8EMx4BzJdA/CEHEexakLYYDvNB+9ZQ/XQrVDEfRNa0Hkx2LY8lOD+K4dEDbV
egQe1esuzmNJNlBKGSCa7+EG8YQmNlNvqbCQnLK+Kd7vJD1OSskV0Gjaont1RNgZ63ZigP5SR8Yh
jEsb09pT+HOZmCk/KvCW9gwDFXqwrXw7FScBGE8P+tcpTDuKgUwIz4JrT5o8uDUtaGf/CkhHBcs1
UoHmjo/bPB0T787T6LQGym0QNL+kACum3ikqk6LyebEHdIEmzxrkj/09i64uKriwkZPTbEUD0182
FOlvMxqQ/BJ0eX2tx1zeXeh3rAAMOUJ5bzU473XAYiF/R2yi0y+xZQaf3aszidHq+tmJ6ShtGt1b
C1x9RNsgMfGR9MsSDYLlCYBhnFyLuoaxdVyWt2y8+4968Pw7qjlkcA27X2ISafAvsr+IBzIQgaOB
ssmv+HRT/QvO8A3e9MGkdy9uM4IC+G1zVB8wsN/BqOMtaBhrQUr5Aqkbb2QiHG/UN6yiTS1jORlX
Dgmvxkqo5Y3TAOa1+IZqwb3qZUmjamMePrpe33UrmbtI6sG3tF5XbFMcMWA4QXK5flVwmFc5prVv
XBHSEyjJWcpAss0QIPKjiZ73vpDT5aywSvCj0r9fTGyToq+2VivA1uwRx5sDMFswEVODC6dm5ggE
TT7ROboQaaPzB8AXC9ThEHGFB30lZxQMlCSPFLtNMeBDjDfg6+lBg4cdcDNbPS3ewtQghQM+DHjf
w6tnPVZJhiN34BbILkVtG7Bl+38zv3jFysBPqi5TFnBoess2IqUZkMSGt2spsv5bpXi5x9Wvmyx+
QqCD3YScWM2FLiZjaSntJvdvAw8+c4l2ilrZpqH4VGrIqjOHXoQSJcmnEvUHH4jgDHcohJ0ZGQaG
HLstvvVb8Zql+O4L1qd/LwVn53XZ1V2WI1U/psKY3BaQC8RVAPTPTduzhmv/e0rL2mh/KWNF3Yjz
ZeMDjuoQvAyin6AXsu3ZHSfWt/nmyjaaYR0GDVTd4a5zlf7CKJHMjaQnPu0kXg93lPB4iuO4Yqyo
1mwuKI9Ig8uxoWsRdFlAiEgdVPUYGM4mXUzIz1xPcJZ0HiKsDq1DxPJS7COxcDzQvr/G9em1UGkR
Y5uxN0hSdksaFe/gtt+yE8pt/tQ0/+lqNVdSrP6cuF1wxWZyGDqzidLm9DzSRHngVeKQGWbvrYU0
OPpVzhSuI+ryk8wEnSgOBS+CWjwCPckbbnACUVJwzqkjI+VW8jUjpwJ+uZJF3x2jeI7TYX6ghLCp
ZuI8MFCp+c6TUjFWCP+tMo3piZjFvRgzfRI9nZOEBhHiUt2UEuSce3ebk/Hjc1+by9+1/7lR8jIF
LX1a0PZ5CSOc5rpZzgKffyDVsfjcwHSgSHAZZtQ0hIbJ+p65h2dzZA+tzXqu+B3dyIpk9Mc9aecT
2Zrr+0g0mFz8jfxDKENms+WNG2npGw8qf1rmkHIH7B1Fa7/GCukNQJanJ9YBwKsFULnz48bxvJvK
26ua5LuUfhmIbVjFhePxo7KRBlCRvaAh6oXVwtzWgVlCgd0R9HYj6J5GA2yXz5zc/gty569a3deZ
zAvZX2b6Ve3OdlYtRSCO/idmJCGolUzphXGB0I2ACo56PB1QTUgiVfzmq5E/lXUrbkY+r672EJnj
k48NbCbWPSnoPVMPC0Hhgs+JDAFxuG/XF+HGAH3TM9zy38K9WwI5evzjDZu+MPV134LYOwv1ZaE3
gV4L73O7yS5q7vxrMiIH1X5bQXB+cyWj1MVXxNw8LGadIIPAz3tL6xb80iG1KvEB0MaYs//im9gY
XwU0XNTpLhKVpL717A4ZnaSSR1LbQ0iO4fVmze1AAVRiR+/VhbUZcm+ehMJsdH/rTUkHu0HkA5no
tMd+vJG4DB+xEB7IrB+Dl8iA/s7TcWlIB8qWreelcDyIOglYDCW4kK1odd+vu4U+z2zd0CMaimEP
8bXZQuth3mDL0Fi3ixLK7rXH6VmB0/ZNGdk7Vy3yZEKIkf0fhmA9NJDMSOxMeLBwqmGKFGHohsny
zxe3WDCQPaUgF7OmYDPQwrXAwaB34VWVJUFjGHfnoJEmeQ6n/TCY1KbyYNIVyyBxJ0nPZamU5amk
c4RoebjfsCR9JBe0heOG7j4IeetiBYCqnnhuiXsQN0DKMyovHKRbCjSKwW5Hd6Yx529QourZeJgm
uy9+rO8/2RlkTByTIJk7Q9Yw+pWlSmpFBtBi6iywjixsWukxoMqO7ghexhOAPHQB+LO9Fmb/3fgf
jLOfPH4xgAF96LhPi+9EQnLIYkoOmKjo52cwdXJ+4/vZblBukH4WQWlusE57w+HWByb5KsY54JZW
tb+oOodByXhKgNBOvIf3MHyW0MYq9eoNVuJR8XT+5+nFsJQFUl74GFBES6JMk04yz4EzXiakFMVR
/Jk61nN6AcVm6M9ZDgq+5tT23YZKAkVeFxq8BG77oSVPcBnV5T7zTTYM/85C/6Lpk8lCRoPHpcti
qh6C5aJsc2TFlihmZZKa6s85YwwzIx4RV6XRy5exTiA1OzxPVlsOiFr/9DoHOkujRvoQBMVNKSuz
i3Pj6HuBtUVni2kVGVSWI0bcDBny7zERSQQ8wVWnIrayj2iUsX4uVIFX9sb2VF6byPZmshUKyiKK
0cXlYhAuKdV8RFDuJOQasbDLoKIvPLzu+/ZSFC2di6SfdIAy6HAPO2X7hWuEc9emdaJe3yUJFAMB
gp2bP5i9x2+RtCDfGgb2axE3syKs4RhkTi8bu6UY6KH+r6o1DFUWoiGwkbRdFUUszu3GGU49QKM6
wFCov5CV/WX1Z70KGktiO6RL/abmUwBQTqMMeiAwb4KrKxvZ+3JKKRyMD5XU1FrJJTKrghorlJR/
RYCAb9yLLIpN8+0tQOJ7EknPCFsm7V01sX68VgprCQCGgZl+ObffZf+mXQimcSXjpareE2H5EPAs
Cvh0t8yatseo7nLVZmv8rsBo6Q9Brd0aXT7ybktcVp5x3C4By3eDjrYvYBE8fB9BbgOxy5ZGuV8e
TDBaDc8ZLRt1yeDeQhgWOgSwSdD0PCbgAQNjbsRp6QI/FchX2flStwPEi17Zq0e1WS5YKM+f+xn0
ws5ZvmdVWvX83wqfrFy1Hl3wpkECsu9GnlDrnjw7vRPGZNiF3xGmbnT5IT6F0oWiDxco8H742qPQ
kZiBMYBHNNFGZjWlB/h+fsAZJ8Wa9m44X0GrkVJNkWwj86gol1DUf+ELkQjmz1Ad3df4bqvkqm91
OZib5xYEtd0nfsBx58kyUsm/19P3UGmoBzsPzkXiJlLZ8K1SrkFUcP/YDg/45rmvUwuXwRgSqCst
csnLsuOaB1eak9vhR20UOZuVLk9VvkTFouVABvl5wvuEaFFAjeFIKkojs8FNEjfo3pQNvTUp87xD
fQDXBS7QZdDc9yfc2bv3zMbo2ycgNb5/ySh7NndqJnWMqCr3TagvLPdRz5lR5Tmf1cS31hUk+F2m
NR3feUDAgS9VyJmKch+9BwkINI+i3K7DqQuqtwq8YqSpWLww7h6afuvI/IOkDOMj+Kfwus2mBeRj
EP2GCRruw97HdZJc35UvwrgCk6pEajvh3bewlnOYuGRaE2pc7XbttQLnkrV+IHP1xZ4wyQju1ete
dkEN8hMYjf0g9Dny4MFAIwZBBiefG8123mnUXPrKv7TA5AEpju9r3cCGN5qWLxa0E8WMnuNQbffH
9d+pqasY56eOwV0jCSVSEB4hk+58sJUW22J+u2NdnzESRAZXFcYwI2wGXq3VbCYpN0Cz/OC+9S8X
KevZwXV2mRW2VPaA0nwAIFHMBzwhxQTaHrzw5Ic6aRDA53jQYkr5LP02LP94UMfmiFMD9GBab/GZ
9Hcbl76ey0b+4owQ3Lx1GYCV474nc8/5kCYd9RQhkiku9ejZ0rCp/vWXQjvlfBR5VXHuyb/MB/87
l/uNWtO0sEzNjdLdApcMeO0VCvmQIyfyVVN08ypMQ0SOzSM8Qe5He4ybsXhKhVnT4EAXC7lIPA79
C6xE9RzCR6ISdqbwz1qf/TbQ5P0H4IU4AzYCD6FDfgdvP4FrRohX/ZyMi8kn/fSb5Nd4L7mBHGY6
4k4C/407Ldbj4dR+fBK52hy8hjqmDB09VFI0x7HCIez/We4/flJlFQksMNnahEthfZT4V0wL5m8U
rI/42H4duYLayF1nQfFwpbJ7/hYvi/kyvgTGf6g1VBOwdWYWkr8bIotMLBDxVCa4c22dnkAco04z
beqFI9YqCEfCMYLYL0OLxRd0sID6f4Rtkp+2cMl1Czu3OTzgL5xbV0mQDvLVWRD8htJIAR2niIZj
I94Xljzk5/QEqJGMSdPlP2WwSTI0FxkOPxYVEM3Hi7TqMRg8Mb9MZPFLd9BFEKspOT9YpzDJ2MXB
QPopZdg78VHtCxHt7nNndfWBQheWm/lKgjjGZH4MX367NezDCyc2skWDDhtWn1OuVqiodvfRVKoi
xlrc5to+ghrIvgIOjbEBWNI7vKVLbrR54JJ3cGmBTDWYlX3s01WLE7GmMkwkP4UdQnB0Xn/P72qh
mXvcBYvXip+29VsXaqkL/qi7/j+OU+ceRxktYWXiLBtEYn3yJzjuQDsdnG4A+b5ACxyLTxcFe37s
HF+kxvv6pddw6S6IHbCwDzJLOLFx/je4CS8VUdt/r/bTCxRCAdEGTwv3LMstSu37BQTBgYXfDT5h
AbeFvzExlOVOxhhOUo7SMc9LtM8oCujiyr4UStbGlsgRvXDvfcM1zfRmskdhAaJ3c7mY4n1UfyAc
P+XPeXc8hYQqEAnuFcocUdZcmYmkefs74Y+M7g8YzpYZRuH4xb4rJgo+zAtogkrnAsVFMXrxiJge
7dBuDYm/242B5HrbNri05b3asrUlJ7Ne8IDYZ0i6xm0i3qPNlYJBS7d2Vh5ndYIcCDP6nhae5gq1
yce/7ghX26B1yaSwCgy0EFNvv4iV+GshkEy89+N1LN0iakGMswRIyUMx5MSiW35AcIXmaCDFmgXm
bgPOo7a8iWDhvYBlap+JaYrefwVjaNCnuIw3IoohjVO7sXazkBqWXLQd9hLZJUXUzlZDQGVfNuQG
UITESK08hDGZkgyEDdXS6tav0FqJjxknAxXAXb86OdW/N2QvDZ+5FJ7L6cWpSfrtGqmenZ7UtY5O
N3Ljq9wkCi5TJ7Ue0KUC+zk2TwVTkoIr5DpBTGgs8C4MLbH3CmSCkPCz1b4ETGlfw8M20vH79Dqs
PUqsE7wvxCR/qlrANDGm/nQ0upwJbmAF7lm1jQsyy8EiI0qTTdHbEDRtq5OeGmqysSzcj9rfxAFu
bSD93ojm9Vpl3xYKP0q4NnETQaMWv0pU6iSz45HlxpN+kBqmIZiWW9hrgsU1lCJMauariqFP2/m9
yd+DkENJkOIz5P7lzP94PMvVYn9v+4ak3b3eQwQ43+5/soGRnRA2rdGMlvsznMVEAarS3xkPnfHu
8VeeCTm9SRtsOobrG8dT5YqOXcvw6DUZ37yXFGA5cTdjP8MdoRfkouYpcE/gliidEdvJ+XRiCKKa
8sqvt2YtgzGaSLCMV9c+/SB5CAxJIUMzhqhWAuj04j9hf5xD4kWSWBgJQcY/4PszfHntDvuBSCwF
bIrTS4fJR6z3vtgRQN6GLAJwuyZJMu6ZZ/WdP6Bd46OebMMFsrXbNavNrpx/8lrSbjfs8JDu/X0q
LuK09TRo2/ZhiOk2eHRZFTlNQSNmmseB62HvT875JOwldRq+2nCRqG8UdpJjSMrmKn+So1f17OC0
F/5K1unyHSfccA4KNhxXiw3S42YmSDlOyFN0fEhswZcFIre3H0brt8OOGyauacxu4VV1Al8V5OWe
70JtSyOCUJetIK7mMZO5cYKERzXt9BoP5Dk573jqe3P1+eIdiPEiK1GuX/z1kDpZRgzfLeP9F+8S
qogkq/RYHAFnGMVN6wYyTJxSS6iPKm1B4BteGHYzPv9ksdmP61xOQnizbvOA0taosHqlAK/IFBhZ
Kz713t+P0irf8uO+1+8Md1eBCyLG6Zywulg6jsmqhEIuJjhbEK6l8P5iLzwsal/ryFYtxgzUKOcU
j9XPEQ4qP+96/K+VKpVnx7fs27OHUr96wiqbKQ6bKdyNGZwEZwAYX/gcVEqA7hsVLgO1MEZqEBlU
NL0j8KMqz/qoCgHvIqJ9IreX1AMqV3kDxl7b52FJzkcqar/cnHqZpT6haVUyKCnjtnvA3seTCySP
rOb8/t2q4r0Fzs12gUgc7TlONIw9L3oLa1oZqbqo2EDhdRSn8UmFhyZRnrS0qeTaRMFEr58KFcHu
GSHBrWYb5eNIkz51UAZA7n1LBWXBZvBVwJPv1Tq2Q4Gfxzt/jR3qN/VNCWc8ztcwTKVL8In8bW1b
97gl5OP6jcLJTV3vvaacGrMPVXkX1P6PUS6xCrMsi9kpo3h9Ds9Cb0TcTZy8pEhxwOewJXmfoZaC
umuNzWaEImAUxlwERXsLNTkBw2vtSmYmoerU3I6SDMsGtui8l7JRF/MZBAVqKAu75zLi8f8CRqBC
dHcivwLxHzjkPx6gRuhNpG+fxAf/v02xVV+X2q5e0gbq6/ujE9k8nHjiC/q5LzvlXCdeInRfO+BO
3j96bQ6mjV+laeOVlkSOPH1Wvyk8Xg4KgUYbfjWgxyOZ+fne9lGWxHvpwfl5iKj+TOX97ROELeYh
FyIPxXwX/Oc/AVaBFhlWwnfJnorh/s5hIDSD7FOSQbgwIGX0S8hTVgqvc6neyELRA2xpyPvutnRi
TmEWVeN2PWc7s9oal2kQdE3uwhxUck0uxg5KRTs+Q3D+9FLuR5N+l4V05GjawBbtri8FZ4YH9MlH
cB5QAt2vznc0EwEipjTbMqik8f74OjEG1P96rMjc8LDGQ0Q5s9UWoTyCKN3TWD/hy6Zr5x0kyxdp
Xzuj32YuBQ16D+0TNaXgEuHV63mjhrJ8hlBIOB/P0ZUK+FvnBuKIpy9mzfgyNPcbU3WJGAgsUIrs
+ZrwH4PHyDYqUQNLDkALJOBipIIZiLJEvypMA+Go6JmIoPC/woDq6vvTV04okAqlM9shnu0yRsvQ
pkstogxaZi12QZvP3g91/bJ7RCLQ03HSmlIvxIZ/rsCV8aBuxjDLNeQfV5Y0GSvb1R/dcJh7WnbZ
YiAIMTC8tx9+EWjzdyJWlNwjMjMIDGptKkWgee0Z0DuQWBzdJntqscu90SZH+0KW72Ypf7wVzN78
V6a0RplQlzFZx3D+s8vtIpbVl2NMsNzUP5QFUuAIEAM+52FifXxybvjfPXk1WB4v1F6PdjdOGaId
qDRk7HmJaznCNzBiB1axVmvCxFVeR8Sc3KOo2X1HlNUG5dqv2zM2bRxpJI/4ss1JqLQd91W/qr5x
wGlwWPrX3tV0YFz7bH2uC43PBQmER4b3r/WtwwEeWQPjoLBjMoyPxxG5lr0HTKo0QvCOKxKn3Yac
fjDUBHvcjctVLvkmkkLguvLnVQVjVh41KYY08/H0KPA76lPSDfw3WU1ucdYR4nz70HhbDRSCsydy
AsjwXGz7eTilOb7gP9i1imKxBU74ef8XtHykqO4vear0+tXRn6DqMq9Cl/W8pg86jMj/eHiLImTp
ta5DkavPRwVj9etxZ5bK1Vk+h5G9QvI6DwJYs6gOuN7TkK88WC8mmwLxwQUXNyNlOvAiR7fEH3tm
+DP1AGpsqjUiOXk9tdEP3TM/METSqzldXVt0s4JIv2v/RNvk4CUafw8Ua88zZq+RZNsx5WjLpEza
Rj9O7V2Km3zYccFuI48hRL98DGlNsQ74Gih5+pjP9FrDkpsWpZWpULEJ4Gx7sHl8fzw58EOcfypF
RBiQdF5u04bWUUW6NXTljbBmXfv5BYpvqYaPwDM1mPRhKIMf8d9KJLloyzbQiFIH9zFy5rQC3JwF
4y79YyX64cvTay1vIgozzNomLu+ouJXGAx2bYHwHrcWucIEgMKxDIpsA4dAlnLj6KHVHnedS+D4X
abYLBOyhbsEwqP8h6sr4Sb7o8SQUXURFpdn1FToeMNigY1ba0YpP1UnV//Y1krzU2TXioGNJPh1s
Va/wHvOzGkpjSIXN9b8Nb91Z5u4PvbVXq0qxtpVJvNplnFTPTn6qUjYcMJwzkrB3AFB8CiFo5ZSb
OgWITwLswmrd+AjWBSVvPZQHdXZq2kizrPo7abiB7wxo4hnW2M6MysizGogs/Hbot5BoIjtCDwtx
CcIyEZrzCCzm6/R9cOIrtrVO82llpGrFIyvTy1FlxyYR7Gk2PTwtAV2D6TD/bWGqJY7b7VfNkZJg
2TG0MihEoUYbIlJE+btxSkwy1uWtufyruecXkO31nN/XSvnGt2XofS2ZEIiSYSeI+mXWiFzabisM
o+VdjHGC2CnM3WfnTev+zDVak6w87TMfTLpn06FgDDZ5ERB3uflNzH8d1Z/9J/5RHn/kwvn27PXE
t/t7fS13BDtlfla0fbV5f4B3pwdXawudoRT5fz6VsHEtLXpjNZvbJulH1lkugt8mzpos4C/imImZ
gSLSO48gle5B5nljqLwPd825LHCO/nFeZlV13Qbg3t6YUbC1RQt9I1lYIOz2ZYuVqO1YR+Qp/fjo
uC/g1ENos1Y8oGrMtuGT2kcWM73pv8AqayJBJZKQyiqBOfSwqjC10lpoRO29wPUE2m5S5DT5r9R7
zWIoErC/t9FDcct8wdmd8xciXyy4P59N0Xt1oot4wVPPpwRISrSSBGAqPO+KrXFSgv5mXPNaaWDn
lBYsw5EccP9RLApjhxzw3wETf29mZdWcnMFJkgm+QDK/116aBBDqxtSRRyK19CoZrO4Q9EVg1SqA
gl/csCAHcI4qG8PAMojmN1o9zZKf81dnQKJLXx7PJManxCZUrJbj/53ZFVYn4AMRE3B+JzYFrV75
SYe9LeDi/SRWcLVyNKBD3582ev1aDzexcV1y2zFpkKkTiIgSVpryeIgLCCUYqezj7W9uWGJ34MbH
lFJXVMXbyRlQmTWYQrTCtm4sAAi/XLMNkweZQBjIVeq2j/U+a7jhkKNaIQfgJI15NTpKZnINJJgx
GZ2P8+AfKm8gD66o3uVqh/rbrnMvB60CaIH49pIPlV9ZzFDg9Iec1vB2sdmsL8CM0j6dELxVyKQy
FwlSU0Dz3eXTqwdPMqwJP0j0y+1kFpGq7402dj/Ih+Ohkm1MrQT5yShAf4U6bkWP3cX3vEZqBKBj
Cn+3IqQ5LRNzH55NaDJdO2Fr6TlQL3WFEXclYVZLE0Afcqh7DKlr8Q9QKPU2EVWKZ8L3JKVjN1Fu
a+F1bjpNUKrj4hw8JeYw7BVrXlJ5UJ45+cQoDzSaUa6rtvggT9VPEQpC3VvNN28LKzOKOn/3rC98
3egUml6POhjyuGa014V/5sUS/wirVKhWAIwzTRPmHSpUZ5HqnYwOFaegvTiSHh3PI+kSztPgqsmt
JMOCi83bX13N9NYI/e4bkL3/rjJMCrexWFm0UT0GK6qb6zevNpc0C0LC7Ct98la+JjQHnIbItJaq
5Y8cmH1lzL7rqbZryiJLKojBiWlvgHOaOE+EtnePpsCowd//3ia6bqa7My1Y3Vbl6nN83fcqNnTn
Ub3akbWVcTWqTeRVaWHMdQIFVK3I9IWYFxqMmeqljiXJCsI9GpPzLqABflGX7PKD+pHADr96T2vF
SDiIgvyxxniAf7iXX/YIAtRIjTXYH+NfQXBJm2xTJtjptlN2vVit/4fZ5hVOrdWF4ecEGkPfdv/Z
zhQgqwUDDuLuaBz8Q4P9UifPTabsAt2wuaKvS+/Qt39e5Hclz8wZs7mlJ8hoTGZ1199NKXTaPwEw
pxQG+DMOT/go9IEy75Qr6uPMPtD9TXBeT13LKZBasZYk3T++f8sV7xIpf6xeBwej9t7jD/UR7GsB
oTnSqq5FbBb3DB0GjZM63qRxtbfC+ngpGgUy4hkSeBW8Z4+l17Z3pqPWF19e2yZLegOdttBKvgoJ
pIjRyvnj7ZLal85Ty0ISnxTjwlu0YigupLl3vF7hOFsjtVB3lsWdEWAJN9Sxy/3a16onVc97v4+I
XdlT3kBv67tQHEXDN9CRL+hD2Jt+lx9LiQoc14UT0m/Dp3rnNtydTptEwwZbtwHqw6JswKEU36TH
zwozkhml2OS6bwJGvFy4qddaO/tEdl4YbcvkWjcXUHPjwZNVXtisMbcFuwPkmhAuyau/PHI7XSx/
q/t0lk+Yt/kvA2Xqcuv1GE+aZYHDnNyjAs7CJ5zcsVzxEqEYNOFDLlyrP9WrBiChdgxX3tvdqrBW
pbx5kf14EwzN3wp3qfc9J5wrZPxZzEn2+JpOVh6yq/bSyPoo5qUkw8ed6XNYvChSsmOzGbgOPeXq
EbARzrEWqhUuqBOMM4F27YTPP6NOURKhYpHbhsRx/jwRUZiCSJmMe9J2CarBdo5rJeA7u1CDvnfm
iRfDuguT9ZaQzQumnynN6rFjGMmozr65TAOlZe+81vYD9vpJgNUaPcF3WelO/uoGoCe9DmMbmc6a
b5yd8Rk1uTFaoMigOvp0dVWzLVyG8VQoe1m52GJNBwm9YlQF6PQuBeNspmuiSSuDrIwOOvwqVQ1G
Iie1s/A0zVY1MthA/dhF6tPmDUwrUhGKRXaWPyHZ1S7FboQumK5OCJ9MM3XFvmKgygsJPidpoEyg
DVGbaWvivM4FniLVZuLvLPtJN9kOX4p3XBdkesk/WZ/l9+Q+nbdWIP8OKiAth94EwN9qaIzsbRmm
IJ1QE+rWSD8TCaro4xEQtFeh5cxfUV6fkyk6RgDH2vnAXKP6vq4s671I2iqY4EzCGqvOrGAD9cVW
p241AfX2QgnQBLJf+pxpI8V2IlQ/cR2O4LfqZeCmHJQhbZdDSdhE7aclbcgeC1wRF+6KbdiWO/jt
3s9AnayTDQHsgswZRF8ZuKz9bDq/AvDPZWFULsttOhuAUHn6s6TYa4jprOv8TSa+yl4yHrNJG0XH
Iu6N/jYjOZjI9yiNH9UGxH7wtnb4e2wfMQE5W1i70xunGKIocItodLmwd6GHbq7Vnx4Dhj1XGXUn
dJYxdUi6asufKV7UjXGjX9MetZ7qyj2FBs5Gi27dFun8Bt6FnYKTGZZxe432xHe5me0Ulx92rYFu
eUIdLBFYH3jYvveiUTfzHLsd9NgNRYox/QmTfTHfdKBJE00OFMHFLCGd5H/fULtB5yzzAisfinqW
TfWnsLE+qoZIrAjHB/Q+7ulODQxJZgHB1KgA0HMWWyl6mhe5Cbdeem4pAE2pjw+3gAQVkZlzsB7Q
2knlk4m/IMIiHyqEodFhCEh8dj/JUnXsexsdusOiq2pXpgL48OqevcA5kV8MqAZgJ/B3QdGRKOEf
leSZ/DAhr1zXZO+U17RgddWBRiGkOfEn/7UBGJFfXY5QTcbNaQwbuaXCsNkU3L79ViDWSUBtLvQK
JIJNhXbKADbhUprcm4dm+rQFY7jSflA7Af5SqOCrKRf2h/DPGRGFQ7mpRIytwizm6Ua2lN6BB72Q
l64XCsNCcdaLiSqXm97XEMVOXTIvav48scWUXzR654zJBn+auV2JosNqZTBhmlCK21XFhARD1k3J
Y8Q77umyoPYy8t0gEjEFfqcoow0Wy65i1okBHhgR7r4Hnj3XU9NIj2vmbJPkI4t7uzzLFEW9/Zvr
u+V8V8fiH9Rooe0kSusQX9WSOn49Y0dSEcP1ZLj3N//LZiU7eOSLckMpSO2FXkIBLEp7w7YKLonI
l0kh6tdSD2RNZ7JmM3EiSwbsqyQcmkrV+NbLmtbQL1ue5Vy2v/TUCqkhywx1o40JIqRxVkWTkFtI
WAgoOOFv/JNFjWXtH65K5YJ/6UdKtBits8FFq3M/QhSaxpjmaub8M05AJt1br/lErLuGyMejNBbe
g3DthcGNEakNcGn5HERwELMwccu4AcQfUoW12HYDiwZahYVxHvZQo0sGN1PlNOvuBZdgTHBzjCIV
hGQolLGQJ/uBICuWkxbQiVPFNrPEPVBTtDkHC9KTL8EuW8uCG8oQ987dOBOhnb8iop66OPWQccKR
joC5rxpkIsrU4gEGmAyL0ky7//QMvtD2diDSusjujmspwieepiuvmvD1I1sRNFeNnjufqjlC6+K0
bwX6gfzZMQryco/H5bGxkitC/IiEgnnm3tCRcPKYS3j4IvheL+1trJf51A0JJhUrPRnoB0UFw/qI
8l4nArUzdFvdY8cle3ZnCwd4G08AzWPHaRnPfkWlIbNLKWtV31pX1D0NvZIiRBh5Inmo/Yp0o4E/
ouMjxSzslip+sA1QPkp+/KEbHZ5u6/OVw4hv4DOAzM+LrJrIE7x+xXNsNJcyQ4VQlFUlzeeL1F2q
GCFf4EeS3N80K5kWISuQ13J4uwFfmTPYrJwTTeNQzHmaSAT5QjRg7vjWUDhUs/Jte5wYfpepOs4W
KO5X3q0c4nurFSZSp0VDYkEWBJnUj/Dh+jt7xiIohreh0o7Hu6JhEbozNooSqIvmB+qCEMazhuBe
Y0ZglT1rtSNdmlb0FshshDcl9QT8MPNw31iUdcihcKD+HWwJkcNMqhK4p883louunBgHQH4+TkTs
BsmHLnMgjhhPmon6jiCYjRt/HH/xvHh0UfJdf2oKeFbtEOm4TF1Uw6Htajp/bAAxL3tI7fb4KsXM
hwNU6YKZDm/4GSG4CGeBcN4lXLqDBTdLgMCBSB29jhFdG+P83qWOkexKw0QoliPNskZFTtOd5ABN
mbRsiBGYn8+8GG+oQyQjb0awIb/n4C1SXRm7s0IEeX5GU/eFxgC65BPdUYQBEhKGkepHJGmgx7j6
sa/YhKJliefqqsVLzL4bdowcLSUr02cDGPfGu4W2iMLqscDETrrKX40OIV+m/E1l9ad8pV9H4biS
Mp7K4jXvHrZJhXoBT0dS5JnYhnaWIdBZkoUIdWyeic+ndT5rpYtHV2d6Heg5oIfXBWDWxjreBHq5
7REwNwfTvNSMYGerMxtMC60o1UTo+BoxQlGZJoAmyTIcGvAus1AQdTMB8n//1cweTHWbMmjxHYlv
/3k9azoMtfcAf4AyrrqALPq0QcEbIMAlztuCboulqbt7l7hSM6Rq943/yRjgrjpNavoCOp3GqTe1
5BaBIiw86Tnw2af7nZfyMuU6sRob5nmZtrv7VXuPJ9OOcrJJFjMV3Rj6OrM8kPkNHJ24oD+mrVFt
TNoVp+fe33FMNWAFyKJJnpHeTnCIbqH2Ryrd878nqXKZqlhCiyfyIEAPBYqPSDk2jfyoodYgntoX
cJQiW1oWUNecnolKd6JS7NtB8oloaN8WGWYQ5Tq2UM2Gl8wR7QtcTPW/nDvDs9wNP65Rybar1m7r
0Q/duFNwOi58zI0IajDnEA39yh5sUyRxfy7QziJFVHqjMn3vWRWSwKCAl13ichYKgQdzAMtJX9Vf
yAiI19Jr+i/Mpv0wOkFAW/Pciy1uk5AKtdM+69MadJmWzrcXDEOwUQJ88ipfHGbiQyiGe8dibcjQ
CHO2163iCU8vkHWhBID11fo87aWpOqRlJ2QD3KY9/CA/Yqkun08YwEX4QghVnHU/PxekZM9Bab4N
8JiE9z4lndIJt2SPrVMgooF8DdSMGvmQFtHISULcl27onyLNcD/wOyDnx5ntIrWVOH1XefbPvb0i
e6jWI8pfTZ5PcwV88rI1H507sxUW/+AmhmxWBI7AACpA5Eqyx5w6y1SYX/eM/eeWNZyag34f1Ugn
gK0AWN9c9Sj+QLEgS9mOP/bG8JxyCh6MBj7py8aW3gqiFAoAZYSV6AtigC6l/XT3aZ42n0oVYHOu
bnyNb04HcmesZ2+EKiwAeUEUW+dWVFo0PkdmS7sOitFYsZ2/tuqHQKYFDi7R7YZmFeSFQXcceaIh
CWInR2WCagCFg+Fv8y6+6isHWRbhU8jGlC/xYpCzcuX4z8lYBwDof1v53RdsXH97Dg0SvB3ncf49
Cemxdpq4l29aat/899H8hMzueYVj9NJfeqy8ORf4HntLvUOtzaAW/SUhXS5Y5L0DkptjXMQgfBRS
dbhcJCbub7AJis0k72VDU+V2Wcpo8bTolyIG9kd0ZwSsHscLbdssbr05JM5RKV9kNxkVJbPnfgvt
QeUFSmktsTLVZgr2OV/4YV29fMpX20QPu73efT1PqnctFXQWbsTIsvCoUqznSb5YxJtE0KSHbFxA
V1E0nppSyvAUbBniH4qCh6MmAe7IU3/fvnm+YqxpXwiq1GIo1272/Nr2yvyDfONYaIes9fv1pZfo
wCqoVPFGY3dEz6Z3arzQV1NCgnn4C4TDPYKqOWxSmzTGNKTVGLen+Agp80DcNOFZv47YRxNp/dGW
mpGI20oNK1ViG4LSaDWIP2LAs0gtNuoFA7lfkoe2MsaLJBE5H+mnXRppINV+6goNG0fFk521C6sw
lxWlzbXvCeaimDvD8+MdciS4zLAdzyws9nlmC1B/j37o7uYQYYU/MtTOSQHqFdGGKKDYydyf3CeM
LN1don4mc9H94scQd4759SYCpFE5Wc/iqPhO7ngrkSI8VpeEZ9ma9WRZU+KYZ8wX4bgaDp+WN1Yh
B96VwBhiXooPGghU+P6FNUqC8jF39Gh1giuc/PRoJ1coduncTxiJTxnYyAmzXuDL5CWzlW4cGW0s
4HuyMKASc94nGFQYB9nnLdtKm6KEizWWekK/5EbtDoC4w/H+71cIu5NP99mcsssEWaJ5FcGpVs6Y
RInAQd+CqMICLnvs9IZdebymrfue4HsV8Ag2t29i4BQz5GU0bOF4T415qWzT3j6K3CXxQssrHCLP
dcJwmhP82jmqaPPkLIxhQHQD2DNPkzfgqSVZ1k+tyDf2RUOD+ksC7eDYdCtIrogSNit2ZrrJa5sd
CuMHIfXvJoKtxXM90MWZSK2Ba39Eq/yeF2cv2/ys9EEaPWmPXiflVfEDKvmCNabsL5Yu1xfJQl91
ojh+Ef7MeBsgK3iARJIUWjn9cyzz8IDEPrmZR5+IToL4aLkMmSfrA61PpGaQRc/XlE9ETqvXRB78
sEv6EKd+dr5ci+DjXur9yrQ3truXOvEpwByxhESvjwCntox8tViCCuVpnLIlXIIxvI+UKUS2QaHf
fCD5I/IW6NbKT6y2TAAq5+H02mFngNu9bsT7VeUuq9gXrvSqAQXUEEHCuOL+ZmHQNF6ZkPLs108z
mGB/ZYuL7YN4Ulc6/xhc5Ise4jNHUGimuK7MY19VNaxy81Dtz9B58l7FoYsNEoiDFONziIwJbJpX
IPrjxVNoGtdkxgaHGDMHhsGSu/uELAwPZb86UfdImDS8Zjr7rRYbN7iG0LCsjnaRT8Bb6fam4J3n
oiuTYT3wmJROAcKNVsrvM/6ucLjv+i0f0V7vIj9IXtMR8mM/ESRNEOhL6YP40smxgMq5cbDsXB6M
V4JVYC7/zZpEewy+of/ydDm+7wkniB1q9q+ODkv3k0nkVEGxzcmt+if+PubVKgPbQnHHoYd1gLTR
eIa6CroOn2AdhG87nRu1dIe+L/QlEnyQSs8utAqAhs1Y/Uge9ExqWoH6G+6gzzlZPUJ4fuF5z2mU
ac4YllZlCWU/mHYaDBr7Ra8vlDmfKsTXPhTcllo1s9osGnG2dbWJoIOKv/6rueGRKJ+kEZnZ67CD
rQI0zSrcmwnczt0YPojrfZnkHJs0CkjT2tRO+9R2fd1swAaDyGf9nHk0X4PiLZK1PJC79LGSeH4t
u+oXUtgI4lRcOyFonolj/CvH5/FgJ32GT7knpG4In+GDuX+uCPpK7Apdwf9WdjDmrXNsXecUZnjf
ekMdJ879xVR7qO6TDiEObrZN/W+EuK58ASNdfcBp5MIA2G7rZKx5olVxDZbEjE3YdRI6JoM9ZNPj
5Qx+FQVnwtNGN94pKG7TIOGQc4fAt2zgY+J1KJnaQNX6HixZs13laRs5daYusW6+2LsdI20fngoj
N6bCw7JUL3YPe/PBT24BYJDVVo7dTLhhDaNB0lbmhSjlKCF3H/G1IQXT6I6ArEd1d1Y9zlPBjHt3
OPROa3tCjyD67hGw9qBxpFuZZydcFRsWDSzOFnnywc40qTRF2HS4n0iX/LQTAcRAglBDZtdrVm/K
EmIfOo727zWfaNPsBFEwCoQiVjJrDwNnfBOt3YphKaiw9n4Q2daNWPHklhZ7tBsN7dSRMPmjc8/i
xx1BvHsnBGFedqqAw4ILp+pnbY87C8hXxmL9aW7mZBnH/KYbvA04GY3m6+0VXx5iNpT3bNaFiGC5
o9T4HSbGCZg2sPk3y54/aTEnNLgAsnUidhPHMOLqgewETVr96rgKJ0IGWw58NKvX3lJ6OD8JF2fP
qhbPn9Ev3mMmfpeaF/DzgvMAGxgU3iYk6bgHM15VO+LLCFnZgiyDdXIq9nru3cpkvslKlUK91HX/
YDF4tfeuJ0mH8yrk1FI6aIPM/zTG9wh6/yANEZPDDKD0ZkMuIv3Eb+cvSKEhA3B0dXXT+SkkIzB5
/TgJIBqqitLQz9NkNuSfnUXO7vBvcscGjEkGcESuBgRsWeL3BMrGRm+r1L/DCsXH/6xAXjTgraNO
K5o++4UyM9ZLiU9BQ46E+jcW4uPDXOwwWZtDMcXwXIvEbk7GG0KP19RpHfAfdFfy2UDHRo0p7mof
hsspdmeM0qgcz2rYTPKPOrjpyEIhUjNZC1aRvJpmPjaI3Ad66wfLVVs3MEKsKdMtlj5SSCrS3GtW
La5pJbMoHlGRuoj7vcwDU9yBduSFpAlNfmAmBB+WKLGRFFGQQKBYLvqalSDHRrK7R6b37AWg6KFQ
fnhyl9p2Un0eQTndt6DkNo1fYwrl/sH1Itz7gxa+HyjDIuVsq5T8KgFJjsQK9XQryEDLQFAOKLZZ
ieC9IVW+VBKG2C8ddWQI4kdomw03Y6jc9gX/jsRc2aJZon3Zld3i+0r9IkhfYNLc4OAYIw9UDJia
ACakYhlOfQl5HRSuqiYW/S2xggNq2J7QWdfiC7GlruY3mAPKZHaGmA0b6mF8pyinK+o6gWb7pSC3
pHTvJYo/3xZh1ud78CEg2MN4NWt6ahazgheXqM2SOgpcYBk9Ufnju/kkdGucwXumFYN4LHSnVacJ
qT0ogxj2T7KF9Mbm8JvaqrEr7alP9mB+RPsZJJjjw9wJKOwr+3iPYAov3XTFJPefxQFTdqvT8x60
p7OzZHENBiNeo6W9e/G6WTJlwmI33Pa1lziZSfdpkvKXdwAKgtslWpzF7KCHLzDa20nCHnRzv6Cw
sUZRVscVYNDPomJk8SKFAyDbyVhfQgTk9JnYPrzsERa3W7EfzRCi7hZT1HhWqvuxkvjB6O9/apIe
PBiyOQ/vXGnQ2AqCJ5A1+LK4uX7pf5dvhD+hyK4YzMLy1mbeVhMfzMBC9zAqIK5BQpHvq+Ft6s9Z
6ZlxlIYTjWFK/S3qu22FLONAF2qVtrWCEJ80eh91nhiXsr/UyjBjn7KYuIXxMC6tdiFil0dHgRnL
ZAJko6YHPJtpFo35YOnVjMqRqG1gqc7guiVVa3DFPwPn65XzYw8FrRVLRF+aPzTmpIIJwllC9U08
iq/pPY31kq0NiXwKyRsJY0kzEu8jdBhV1vwWnTW1PXX7jlUsXZLnzq/PYx2to6Bh7Cay+OKXX7fj
OQaTxeMFS/6p1kfS7r4ynr6NO2uE6oqXFa+DHBwMqUbT0O40tI8Cfem5DFvDdC1jByZ50+wmy59o
EMQ2hwtKFWQlyT40Rut9irWVfUCz5lDczdjTEH46VR+IU0BlNyDXmJZD8RVngvnfc+uNTXL2OSDY
Z8/GrGMCWNINMF33k40Dx9sn9XAX5uVZRX6w6yquF1r9Dpt08DfiY00pITepGg4Ow4jtD9kfKYkb
JGeofp1CjAG1w4sINfUcV8vwRtqGxNgofEDnHuEN54CT+V3UlIeZYo6BoQfzmrdPrEj+3+Yech1R
e2XURfsbpiYChXSiGxtnhVUlE0p97o6hbOqh0u0Gy/8+aO9qsf//bPZm0nl42UYg8CV4eLIr0gzq
b1fqlNjzeAljYCGj45J3gJj/hEv7mVgBmdlbSE78eSLNQMUTpf6UEyAimI9aGPfw3vbo7ssLedfV
OaSNopTyCMPxKFsLT7CwSixYS20aOSk1NLIueczOr+Lpg3Ql/C9X2fBUCnw2bjWVsqydDGRvqaNG
eAy/FPoQQGj2o90gfP8QkPEB5GAGYr6ubSduKCboja372Yrr9N4AAINHLw1qlDgw9rB0i4w1kpfB
mNQZ932f0Q61FfpGs0X2I/QAFhSP5fBM+FTH3SZ0KKT+HfgtSSuJvLAhh1YG9XMSa63ffnlTY5IU
frK4F/MS9EQRgW2RD3cYYncmQSH79euQ36/lJds+yX6Rq2DmmknUSueMTx2i0w+YhoT71iiWonaF
TPINV/7xw8IwhywS2Eg1xyM7VIdJWMNa0AqMFurFHR9cbzc+wuiPq5/isZ2BzeQBmMOO2Ul0U0qH
QoIGjQV9qm23UAgmCxhJO2/759GgdUj+KonlpDNAwSFNGR1RxfuE5PNfMVuaX4q7RgK6F/jClEZo
tQcAKQNEOadxMkMSTVjRalEKGoFpNm1yO+13eq9ZEnhyC/2TtZtmbkasQ6mgazkDgqkgjAlIHusK
OJ0afJeGa+sqZb2XOJWqfwlmfA6o7z2DZ8cDM4I8ViPL/Rlw4ZIYdJUWL5ahxqukge4frOHyDsnA
oNq1+QwOWbbCNFSuIg0T35PRsVWAr6OkVsFnVOtiTpP0an+N635e1zOR+bh07bULXBuHq+z+gzMA
gWWLgljahB/zZIRtqr0kUs1ctuXhyDObCr/HMOB+iDKa76ShurHlCjHpoN/7TgGZH2dMxzy2L70F
Wync+GJIYngYMNRy6u0qZDy9eGtFc26cxttoYSHK1BrccjKBLhdI/Y75JkAxfTsTUSEwtPS1H7my
jjQg4DOv0cnh6iyarQACf+rjMXpKN+g51xFxUiFzw2AovnDALjY7fdnE8wY9vK7Yd8qNfhIbmCdw
7xqj7ys5GRZmudufDz6XzwcPetyLLPWljje5qYntIq1f0UAq3NK30kGcb81zq4hfy2jAVJdfNJAT
iYIKsIaMTOBZhN126G6IZF9rltzbaoCfq6McChnZttWXycYKqqLfIWxnviveLClubEr2UpH4uxtz
Qm0LzbWZPzMIjEa2H2CQs2Mc2g9Jp44u7B4BENTmJS6LYJRFryGgqhLzw7WA/VHA5I8NIodhUT10
0abcX4Hf6xUn+Ikwn8cVh0GoYswZWGOUx0yNiUxjaxrs5wjJLljlQXBgPb1M2hXOciYQYM5MlGKg
gyswU2qlGe5y1JHRMuVkB2G+faQRZveaZwYeWP2pC8uFcBgf3ChAvoOcUSRWx23AA7EG5hBW2G/Y
CXot1RneGEhhk5sHI5iwBou1yLAKNJm3fCkQb02fzBQS/LyS2bmHzDfaKo1nHrH48ErIX6o6XLbc
BcYyrFxOMLqij49giWJIcUmA4AX7GVEOhs9MoKpoApAOCfxWfzqaLORq75gm8SIr1kKxRVTOzVJ2
ye688xwz4Pmzf7QMG6LYbmHYfz3bPlwg1Is8B4WKeBAKswUbLQXn99FXTpTwH0pFszB5bqkXL8ac
PX8zNOHlurp77h+xDwZ+LUASNqZQOPnq0UME+IxaVN738D+DRnuH54L/k5rsyXjCwS7U19bx1JiQ
cABnl7xcp2yK9ZauXMcdzmECJZwNG2EM/safiDdwyq94uYm64hDE3oNhIZucTaiiRv7suRtHZXDE
XI4dtbfmeluLB9omERsjz2HcAph8qteTP7Oek9BN/RmmVG0pAA7NW9xDXWSbENwC43ZvvdAWZ29j
0ObGdSVRU8OsOB1Bq3mxnFjQplK9I7ADKmuLK+tLqUlU19E+gxizB37f89pkYSMHVOFCdLwKogxn
bn8jNKZ2X04tLOwUoF6t6mhb//ZNHAj+pu/RQjmy+Zbb/f58x557oekPqVYhEaB0N0WuLsYHUFPS
bPyU8Kx5KUBB60oOkH6uNnnXEZmyZnGdtY4Ua/Z/TOR6Hapn+LtoPZT6A86Out7ae6EniJVDSaN9
vGSk4eid6RCzU2aqamCCwODNOi2IXtJwQVICRL5MXBNLKtEwsBqCJH8KBA/TlbLzyi5XQKZeKBBc
zrAqf0WkmDqbirdQ2rU0WosR5RqgHqVqjEtLvP6ymAza+iglG6DX0D982rrsW7U1s+3NwDGeB4HD
kSGFNPWLtxWc+vrXBCNpaPKltX0EC8ARlG6EsWlX7TubBmjz+uu/tDiuwIbH+XRLms0VWVk7GVQW
+1xgOiykcnn+sYfE3wfO3zgKrDecoAsT1DwVgxo9CUYAhy2IvKYS5y7REpKC9YcVH1/sHMydG7Ew
vD3s0g/AIG72a993NQPRpOervlzGW8C4o6hSMUIQQ6ZbklDlAw/CU/rHD2y5njFTLyRdGBDB8yK8
GliAxk991ic/4jlv0I2RpVlLnRHBWeMGf4CtSbgXI2eYiXFy3y8kTtQj7JQBxEKClwNKP1g/7LJL
N2HAYYqM7tjhC330lswO0fU0rg/XxzJBXZIbEs8z1RZ388O3FCDdRYsS0e6f5IYSypp8pzewynY4
SZZL8wt6RgLUUebSITu5AfJ2KHX/FhZN9ux/SqO47oAif3Kzc1r+YLHk6fWjym8N7+ydw2/le9R7
g93+pAAFU4mFbWg76s+4icyJ3gQjMJIvQ9fn1wEt6v50tayMERNXySpT6thPNW+q80688nkIqdQv
sD9tVBi5eDO0I7gZ/I5s4xDRC9dtoYvErKFFQeR2VZjjshrd+IMn/5jF9+5Lwmi4gJmPRI54CurG
g941tzgWqBc/SIVyufeLQ8lwYPxunW5N3JTi+XbT38tugZrsWB0bbbqLEQTToFG7Hf3+iXmwnWxt
SFDJNtgO3g5BOScCqORkPPpyr8988NGWB0K715m4CDnL04KCYxZI4j9mneRmWXKashFiuPRnQ1h8
nRf5wRH7sBatbHg670ZwdaGvjZE/7KdB1OMKerD3qCBBhNyU1cQS9PtCuRQrZo4CGyBKgaDAWUwt
JWxJpf/CWXHjVPv2x6ZhxanXZ866anFDvZEvs4BAB9TLsUIN7af45MkJK35plQ+RHP3TbRysIpoo
R8e9lo+vjTNqVL+tk88hAoWPy4Nr4BVwOG5NjoTclF8EBF6/VOT+LHp2hjM84bjI2jY97TRm1weJ
T6mUKPVpLoeQecjagECanHZZZ/y5C/7JHHrRzPLZd2h8KcgezQbcicuHf5Ud4ge2DGlasg6Euw/a
BilHYQvM2v0wY5haYrHU1gPwBfbUuUQVuTZ/jjjSTKo+/LrMg0u6n78lRNWLoh7qZSc0O10fBXfa
tTen30d/G6K/bB74CyCLHBxouKFbKkeMcV1iXaZKt0nnpzwB8lURXdKMJdPRqI/OflsOpfplvRzt
QlDnyr+5imJu/bCAP7y5eilS7+/Damp1WyWCK19VGCxjmzTj+Pr9Ps0pjJ/WtaQCxT3FklCdrNJm
4T/imS1Nw8b/uLDnwPv+FK5q0DbKkCUa78NxGPF7r/4dxw7HYhy7juJOgsbPQgwU+6r10UBbN0Bi
Q8TmUmXUUL5Z5iFXJK9ggndqT/UHS/bi5DZ5haDg3ehTmEwRmMZFFBM+5u4EmXq5Ob8G76zb42Xt
UnEFizyUbVZx+TCzivH1xRh4V1pmhZisolKiu91Xe7gjssJC5fC447rbAFXc4bdTztFBYD7BDSwN
rXbNPnWxDQD11YcIY8rnSxnIbp7em3f8jRAw8W9heXX9yAXWc3/67rumnDL0OP9VKf62FoKh3vkS
+4sYB7vpYE+6E3mPQ9KLIFY1ur8EzqTGBgTOtPqJGQppMV0BqpvgRLrUOIhVGIrKs1V2DeYhpDkE
HJjCjGqpngsLeiNd/2j9Mx/kodZ/Y4szpWK6UOxcmv+2rhuURgHxCUNcwKsXLxc2Wuo+X46UxyZ1
RdhphNQGxAD/LA5Xl7cqpmD4J3szgOgeH9jStSW3WfwtyylcvIGz2bPFJ3nSEp7OnDs91iHyN8/I
SzWpAgkzYGXOrn74fsqv3ESI+xuI/Q8GsKto2UZxurj6amvM8XwyEKosA2JI8FczlEhYGn1bxPqO
pl5BPp8XaYe7HAw9nuTJQ2RJ4BtmvhRT1ebyIK2iHxIf53HS/kefgBwNe0yzM0kngMykqdA9u4ot
PpcZx4Q0Hv+GE6eMcBBIGHPjz/m2WHiXThrCBiYe2LTL8CSuxANpeJPuUCycK4VZnpjz92dqzyBZ
PnOYClGLeyvxaVLoxts4ZZd5yXx5dg5tbncpxKhPhhCyGzRGjj9jfds1hXnSIKij24WuGBl+hWeK
b89DrJiH4NFoyXsEtvoNgTrSK0242sGKEuqYplePFMLPmvV7xvEMCmEPq8buoGrCcd7r3pl+dEQw
3Rs1jR/W3e6akHAs/sb7Kukktqh79diyfs7RZqp1Dxb/fd0hk1FjS3Fi6+CSC+yhmat0ZSogKSzD
Mv5r4Z+oU8OpwLgx5Ejp83PEFxW2fHgE66cBsFxe0kmPb59KtUIwATIkkCRO1i3yZ65up9cbrWVw
KH/hS1hQBOq1uSCNv8hgWJOJQSkKDnfzLat355Qx737Nyl+GWRCweU/7+x2HwJ8dz4tcmN8VTBvQ
7vxUvM5aMoJaiEB1wbfEZmZx1NdwWzVzazQhws1tMQvHngRije/EzECm+/s+EFxGCutpJr45fd++
Z0BVEnWZFQi7i0WbkQtFxc7asfG8YlJz+q1uHst2g8oj8DeP64smzuy1smYie4FLGcMgovA85UNI
Kop85oAupb28uDMsv96k8AApFbVZBp/diGaMmHxApxRor+QCKstIRPWPFtypVmpDGFiWrmS07gO9
Aa9ecCynIYNfcC00fdwM1A/A40rZgkawhO0XwBhUKAb6XdnfH2gt0mzMZ/sNo/cAreIOcS1ZF0jv
V0v9uAlPsjfMxs4RSsHGpPc5hKqTcn2kYB/bLKQaC6vyrqXJ0VtUNe/DA+yHO5iK/T0lCMUzUj21
hjkOp1QaT2t3kMLT8WIxpxGS7/O26y53Ur1kEFkrxQYajltwuHwV0AqHVFG65wYpTAqc08BgmVop
s6t4/aNGEOR/shc8uVthEW3vSNWz5sR7DMs0ROZ0SOVNK66d6vhKBTDGkGacSe2GFTtKYwgpl+9v
uphizCchBXatdnlvmaiU+xp9oS/iIkyDRV5XjLv11umNZGABGmu8pCPz45oVl72SdT09HfjLKkIf
molm8BlIOkBRL/atidGbj8P5h2mOL7OLE8EYB0KgMi1cNmLtUECMUmNUqBuFHLpIt1IDTnwVf8fh
vFy6CrcbOt+ZalbBG2GqetR3tEe5EamK1Z/hTdCEcdkkoZaOH1GirST1PFUuWjWY1IDzjCrpCWAp
tSBiKSxDhKl47Wfpf9dKJNKUGHDwxWPJ57gZO/jYwcCHfHBsn7IzToW67dymAdz6slAEGlmv7CXc
rez8u/XbRfzpBk2ip5XL4HEn9e8larQR2qlkJGS4HZkOVDBEew5hvEzinHPG0jKsIq/o1soWw0MP
r5QVsN3OLDhcBB/djU5ZFjLDmnntbEfI5h4g3wGHyOrpO9dSkoSpvdi/Vj08m/j6tFZl0qvfvsls
kB/kiVFXzXr9PCOFTonTAxzha9KRasLBYtbFjRfrQ9/J7SLpQ40DWP10fCssBWb+zORWJ9ss8emH
wZ6tBlhbeka3+HZosgaXckfOfdVT2MU2wmbCqYCvIuMrXrAyE7wZTJ3O6wK5s2hIWdqtX8QHRPLJ
bAdTWVNkxWG7Yz91fgNvcR9eM+cMnMR6stjd4RO5YpkuFN4fR2B5kbgdbxsAML1379U3BXkvuU1w
IorI8B+2VdNnSbYyk4WWWttWbKkxBjvt03nmueO6G1NrgFA/rxtv9M7NIF+LhsyJQ5jfn5jIOCmH
FVrgNoPCDJ4pxvWIZjxfVUDSTjn2q5IDuZZNyH0nazJeV+qubnzP8X24C6nyy4K++zTWb5MfTQet
kmN13tE3NqrGoE4X+ziswTmZzlj8P8xwK1s+LEq5lxeJIgc/55qRB3MtP0k24EMq7EV+7AEUBxoj
swnZ6/LmR4fsx50xK4qPB9qVxabtLGmdRWTfXDDxEjtOHhfPOtUG9ydn7+S3lcyyU2h/EubrxxwY
u0ONbAoSfEUlnHPrIjrBKCrUh7YUCneRPImmBJnKqzqoJbofv5AfcfWvejBEpT0kyGXR9ZV/+FTX
K7lMJz8oDjoQC5tIZx7zxApU9CoxqFqmsTqqQmVkYJGxvSKa5oi+rojF/D3blrdfcxDFNNnjH7Y7
tQokHV/BLcbIv+7ZsXBA94dMmJ2YPXJYht91wZHUYy/QsMv/GEYJvjzBzvJDXXxWssUWMZW5daTE
oZAezPBe9XB6eMRFoaj/qyYWQb3auuZYD85DELeWHt6ewPpBhqQqcGilhvkCeCFLGKZ0PZ60Qixn
RLRbCLqcm/E2y1tXIpzyal4aP4m3DqxpMauOiDp3d+NOghp/3BD2Awl00U/AoNmyzuqUKodZDAKw
H1EJWzWZ23nnU8J7JHRhc8j2i8ALSZoWuKCk1Bm4gQ9Qggddi9Cv0h3Ugb6UIwqaHAOHFq1Pdkqp
IIiVvhwpBeJopm1gJbsIATvMurkwc0fPfZLnGDu1n41BawdMxZeIHeP8JhDem6EF8jYFLtK/fgok
BkQfWgrm7HfzWMKuJ7n+lr8swWQ+cRgZK+SkUry21anVyKbTqZUUQYEiFC6UIT+lLCopo2XVugct
bJAlkPjJoJyYSmzaTbm8Z7/77aSfXqoUTzHdQq7Vo6Z2Bgylw52Dr0qwgF1KhxaPs+D0KIFh+aB8
N/ERTpa8lW3iRt3HY1qz5BBXeWDJcz2ss0zohimdoSyBr2sT7pR9wdDF/+hDgewfXNRwcBeA9bkn
1jhn9CGF6zzxbiCn+6W7yQDH3dkFHQfsAbK1F69tKWGH1yJhKCIS+XqiMZROfmGNH2JHip/y1zGt
AHnOWzJZqkyWJVuRT77wBNrhYP6rTR+TagiZX6YG6GO6uhAXTajg8RaK2Y/QPWrxvPCKghQ9HnI0
7PY6RxanTv4KTTu98tDakVJywF0BI3w/JruzQMyF1jAmtQ+bBTI0qqrX9MohVF927tmtJ2j+316V
qmCzpJUGs3UI3jBD6KSBTdGqRnoZ5O37BTOGVIq8opCLhIqtYJTs2q03AKWGAGvc5yaTDi8fpJjb
UA3hgC1fBSEJlkO7Mm+PxZd4K8g/do5qM4F7O4Djz5P8uYAQ/sAEgy0yLO61zv4w55m6zDy4gsyT
n3D4rqGMX36y1N/nC3TRLDHFo3+qcHZsNx9TOkefJbiWAivWPWz3R8pjeho1Wz+2dB15VBvupz4s
tNS/dEG7T0KrmTyZJFxNZvaI4sjlEf07mSe2DBRZsQ128xHo6m2fPoQuYIYrqBs5tX1dCueLMy3P
GSHsr0/+MbIWn+2jMQAf3pnYFHnScmbNri/UgJahTAMG2vuwtf1Ut0Wx57Sl6BjFEOx/2a+KAoNR
LJAI3GuX0CTAeVNNwtSK4GboVX4ayfozRjG2OPln9baQIdkQ+Ru63O6MynOT320PgsvTRzXI+Vj5
WZAgvUsi17wb3/2qnEln/ts2rCeX2mIj06gV7C7oKgtoadM1VyDzRwpspl9izNR4Xdf+GTz5+3S+
kaDCE+6veQ99Kpd0zU61nXznKdYsUnWQBcsXa1sMWgzktt+kR4I5MpxRTaExdW4bCqzwpYorT2gU
oRNiFqjZpxnsoEWRatWTJhBtxPb21o/nxDwU2hpOo+x46b9lwnrOeYMCUCGM93nwAy1KPmLXUUrt
qVIruwcuMU8DZWkBwhF6BWrB9u+fL0UajNHISB98LjZZ73h0s3+867QVq+RsFZrUv1/xAOqcY8RJ
A1TqB8BOjbwnG9bEvPzZ08VxdmLiuv/rr0f4SZ94QopaHUt/f7bZQ/v6H1OOS7i0NXGJJg5vlifn
+Qdt4hsJoqYcCpTrUdNHpnOIxVOQrHN1l2n2mu/namqZNo4XzfUbmlOOgMh0yvdYONes7hQoYvxp
qphaa+kX8xcaH3yfKAKpiqxD/JvDA8QSspWVghmJlibroumk8f0ygZbzfwlySQZ6RsOyysiU1Nlp
8xMCt2g7bAdlqLObaDY5jEmVs9DERkgR/gMNv4ZXt4iLoofag1viXu+u99LoCHMjPZBwkipWaWAe
TWplidFXzHFV+WkxbdK8a4vJjJrhmOFfnCcDt9Z4mkLxH6sUjYhbfXPtX1D9ldaLnnTftdekHE7d
xKi/XYtj8DqYhXc6jAU+jVscqmwoEEplL0CrnEE03DfeJSyQ/S8bbkxQr6PBy8HABxFAlkwekFCP
yeIs6ahAciQCs58XuA4d3mb8+/CXzTyXgky7eP28ES97EY6VPIGjekfecO2ZxSrcb39XXomx+GmB
M5/+3DH7IEcEc6CZtK32c0Gs+r6Ihk1Hco1f2FY9gS2n23y7QO2GsYgbLEn+HlsUfyXPIrBsv3in
riL+rWomw2Yku7gszWE69a7lErr9I1YiASjR8hj4GHIjW8IUVn4MS3Lvn+vwUDT2Xof2PjihKSZK
JYNVLa4hr9zGaSLiVI53hk1qq6IpHFgtI+kM8WvinwByg5OHlflUA4SaTcQZ4I3vCiFN2FnmWAkG
Vc2krehzVthCu8DuNrzJj8od4NqKL9CRyefL58SiBneQ5lOhZ1VibgcBvoNggU454alvDe3Bv3Q3
QuK2clJV1vW+uPczx8ZV9tBSPaSvdelS4Oro7KbTMLrcT4RZfJyqrkjZSheE+Rd955GbnWjNk1kr
OZcnb0rdKdy9PeoHfi/B8y2831DP7GXgiBkU5CCm0SrchBpXgio5OIfllJjdwIVZcJQpyWm/NKWW
oiPwwMpOO8Gf9YAkSA74QFMw+K7f7c/ZK5eDxvQ9LS1zVNuak+dZNoLW8sgi66gkXkk0Cr27eMVc
r82kfahTRi9T+zfBJDQXusHAQ+/cCXW4hXd5TJ7sgVyyuchJC6LirQ24ANiGZGO9/shFGbIoZmY5
IFAXCoWFvHHrTvdR2d6cVo/jZLiNkGuoVrhXes9X4ZyBF4OCbNYg30DrJSmkN1LRfHgNvqnezfo9
3aKOusJo2rmLLRLBP/39CFZMHOe6/o+RS5AIMM5+Pyu8yGYnSv/gRLveWKOL4jlDm/KwOPYjoFWY
DQS0h7bhNuj6SVjQOGN4440rIXaoCQM7OQUGk8rnY51enpqOXftHH+zs9xdk16B+DH14epD9jfaW
jcRSsVHgP9VuM7kdamKK5Kl0e2Tu2VvoP3y0AMatSlTSG8QC/39UwXLEDW4OYyiG6gLJBX89zw+H
9cj9LSnW9ml7R0ag3A8lTXxNNyvrCcrzT9dman5osrBwDil/D/SDKj7bbdlB9SWVjYt3KcHejd4V
n1aYVkFozJGPq+9Jk70KUdCBMY9/im7cQ5yA04evb/7qn08YZrToaYqIve9AofGoty1M64j/kAN3
/5Kshl8L/OokSKbbN1ojNhW46d89qLpBVyoZ41ZMGqA0He5AwSlCizZvzxM37acbObdqUV8U3Nmk
aMRHHLfkWxKTrbiqxajMVamrpykXWL9TY21CvyJa36OuX1bnweGXJ16IWXI7McGcFioqHo7OU0lv
KyjN/XiL0cYY3UkoeSRJu3AR3URWyTfObeXdnkkK0LW2RCpb6Ip+3UnxZL0Va+JPp2cQlHzZjrVP
2awz3hAl/Zi5QoVucCfQBYh8NY777KSXi1P3TF8wDh7k7ZYLae7z5m1eUEB8GsK3V2JtbF4FBd/H
w5k5lsDiNheIPTnXQqff8pY8ly+wKKbELFJqzwlWWC5NjqZGbapEdLUAQ+Ft+xboxTSzG292EuPC
6oOv0wEKZb8Rx5Cct6mNCcDl37LjTiuEhOAXfsJ+QVx1YcXvS1m0l8pdD/vjIwvZQcFvA5KZhvtl
d9D7+7BsETvXxLqgaLIKxWJQR1Ay0BNgf+p4eRmE8UZ4LI0yySKmh83oebCI4FLXM1PXgECuHZVE
Wt/+d0N9kgiwsGcow41PJ2MgvIafvNomRB/LrtGp3DaoWR+PZBdvF+1dF3EMNSGce6RTeeMIFwq8
husE7WAurKwannQ3A9OGLPDggAoBzXC1zZIhZ+7U6eOY59jWU1KnZUO8YAtYHemz0jYzWHAs2A4p
V+ZcyLrj0fE/xSnEfzVP8EM8qVPNXD1THK/VJxZMW/rLgFYbwmXZ6kXZgGkpYc7A/d0L0hfPKguc
nYohN545PILccua4VZLO201uDGyYRtGd2dz0VfBIgW8ozeADVikCLv2p4pqAD55Sn2K0+jGg5vxz
N3j+e6HHCBf8AvAR030FJOzaIqBFXmFmyumCM9UXZYTh5HM5Jkor7lnnpuViTdiEzIphgGhcyC9Y
Uyk1eRBjmU2utp+9n2Vozli5ut4Q5b6UcyKJEkGlG7680ytCaxK1ndTEwD82FtjHRX3Qrs6UI5PZ
f3LMJC6KjYp8NUrplfSYYTJdIvxJPU6ZK8tvD9iOo0czpnDHk8GP6isojRnr7zKHYKVDxCL+tx6I
rYqN3oAsIlP/22dp9JFvePh3kmpzCJg780+Q1VVkpejV1chvYNvhJQq+eiz1VPjgJIw9npqm2mxY
BnAK+QTawuWK16K1D4qZqnjRAZDNOMQN0j9s726nf/XAXAmrbrzq9UuMEN1CRy3mo+1lU9heh7qZ
C0i7rf0kX6z9OiSYyQTUT4B6jzbDuy0Q1ewYhla1PIOQgq72zMMhtRgFQtBvCR5dIJVoznCmp50r
9ehrEDF4o1PlWfW2QvzMin77MY/VxD9dbwgm6FV/aRVE31OYfrxnVjvhwpraqPhadRp3Y2CkbjkM
SNX3YrQKc1MAnStRIl1pPzc96SrouFvamoTeG4Tny3Zza+FZ7v7YmmvUzLMbPhN5fRUo9Al8pGal
7XAOg/BWck26s+vqamepfLA63mWTPhi3c/z9+YHcJQwtlNZfe3KL8DxG2ne2bPp0R7zfdD9bCtzb
uQueFam4Qz35ZBzyvoTiIEHUw9QUuF+vuzF/Em5s9Ii+HJ8AIbwt597aGmoAhlng5RMaTeFJ+xC7
zmO444E1DjcDPAlifgDkSy4Zu23iEnxYIcMKylwaQ8EJgFUMKRDNF9KnsLe7kOi+2AOTP9t4rkAW
a05qcPivOrc5k1SqREmGXNjFX9clYt+EEIUY+C5YyvARPVXo9zhPXvNs+2fHDxqdC9TYTCcmfg+m
yjm+8hAiNaPC2A26Pm3MLlvkFn7GmMOsXpJR+LsknsCB4HcVDr5AGc7xiI765+qkD0t84/k0eZGD
YtAuXOt5lChA28p15reWeh2p6KT8WNAPkDg2tLxj0tpR/0K97kTFDAGiO5+QMSGuf5X8fXXVS21c
WguA95u4L2/AoxvhEu1gink7UYarRiHMak54c/WwN28s86PxNWf/oyyke9Lop6cdgbK+X9WTfH+a
LtwP1bO+R2uzgQP21LizJqbaAbcj90P1cLzIZXMh6rIdf/2qwInkmKB4Mjxh7Ic+Vzoc7eB1ywJF
m4XYkDaq5ZzSPEcR5wMtsTop242iJvbt5WSf9KEH5efIWfsfG5Kc4n33Q+ifm9bljOK8YjpO5bZi
OwsTzwCTbqoNMlWoodjjrJVcyiKBxVYAwXPsiv0qyPlJF9HUCXNGrPm16tXmPQNnk0YXmjpOvJNR
/8159N3rT1cLs1Nz0sUPP+LSbUCQu7dIKNMHG3pMPWhPDNNyI5v3JkkU11636ctn2mRkCBrQ5NLH
jO2jS4k2HlFe5k7kQxBuRRFyWANXnOHZajmFc0zLdTEROfTMEejRlkOvbumhtlofW0tnjG0VAZRa
O1OLlbHBEOh5F5dV737B4uSmkL+ugfHiwZiFl3r/DYAZknTb6/fNDmzUzW+qezDFf0hTAErCSQ+f
6knCd8ftWHs44hDQKi1qH2kQUzHUvX+nYQBJbuFr6PXhru/gmZFD6Mo8WmCcTjLGSqngOaHLGPn5
1Y7wlZE+OUFLMyD0OCPmPi56T2euLe3wNKUqS472NMhmr4/Oavq5myBMNNF4Say6laP34pEBqHTl
ZpXv+FbA2fFszSOLGfv/UTvwTN6/RzTbQ7V3BKixlxTDfWjiC8iZFEmrSk51/NzkWrBJC2r1xtMU
6xOelrTccWpOW2p8BCYRmmHoWffvxREK4v8GULjkzOIUUxePNW7EEbHmGijnvlYE9MI8RGl8y103
FQxoQqjEIng32EixohGwrtWkvWvPDogyGoteVgzuzLC2VbpOU5eXK+ugzCwtH8NaFRS1iNqW8L1E
ZApLgHnwRMU8zs9mdAUb4KQgB8VUK67RJlCOGNiZf/Ph2wxfQyQ8ghXs6IzzUeK3jocjuUtDUU82
e4JXyu4vE65OaEppbi+TNbT39Y2JxuELcPm4sVJJ/2PSg5IY1ODfScDY2sxM6aUyEcuoPOO+xjbY
pJuETcnqPJSsB+FXE0Mk2nyhP/nngAOaIy8NCRiB4wtlSjH3Rp5RmPY0452X+bnqlvRywmVLOme9
ZLqWWrG69RLXjZlybL80Hx5JHCoIe0xnp+tKeNMqzaoA0I4KadZ4WvF7R1B601iDA5kK3ToOkchJ
D+NUY5a3GvWeTdbRV2zl0cArNlWhqYRbvaaRYuYkGZ9kSSABmHcpovkU+jpQOcFnTmAsC5OWuJoK
w/E1lgIA/oLEG+x5vW5R4Hio7KyTbV5eSpuTWUFDan2R/rjLV+KeOFIoiez4KxNNtwVKSnqRwSnq
l7YUgAMxRn0QAmvd9e1315y2DqZ2hPc5wFG5o6lDFUN38iqNbfbx+tQQsE529e8pBbFWojTOYL9K
OtyasoruEY1ssbeephroCgHv3XWqGEdCLCua7OkPlxd58Is6bt6zucGMqDl6wXlK4lJGMqPXUJjM
QqD5wRtMrJtOGTPaNKvdVRn6UL0xu+dm65MAKmH+QCQwwTmohxbGpzyxaliDfzUY3Uv/tC6EWttz
UWxfftaudNpl8F6+6ZnQS7mjhBXycdwvpfQyl/pFku0j7roKKk6YJMqccRh57hhZTABSy/joxnVX
28k4nDa9Q8ABg5PkQEPBOmbI76OXwgK/3o9Jn6R+hnuJByOPtXZw6OP/JK0XW/HsW5fIfLOqSGQl
Ui+zPw2AVNbCsmeZ1y9kwaP+AKAozoIQ8r0xJMsNIqb43jFIIxX5I1ZPFJXFPTu9p3B2dbSP5R0l
XAUOKb5Qks5/v8jKey+Dc8VmTPYn3I8Tn4f0daFVHut/+0fZPc4RoT+lRucuCH1V1tWM8S7e9bhN
9QgxY1iAM9BqdhEmqJGx1WtgonY1e+2fdhwXHeonXbvSqCA9BVzh3FWm9OER1O2dtSXfdbkpbbIJ
B1a+5X52Ad6bd3eFuGTncl5JpnwEWBVlpwW8KY5RNJ1oGr5MXj9xWfa030BVHtMiGRjKYkzYkqQV
qKH6WxobcaDjWeGEDcjWifLRc1dvxlqSImW7zPUIl5AQ/iKK0asKMIJ/bfR1Wx+twNb+zkPa2LHf
rFBJ4mRL9i92uoB1s5Lp83pZBgfas3uM7qGadTIP0H/YcNxA/g70U1qRvbdnVph51CEhERTGmckf
oOOiA0joy1xviKOpwRvj6AvDUgAROAxMa7WcQsk9ghFtiw8ZsWX2MpYE5j5nFz6/L1ESadH4QwfG
zZ+w387UlnYUf4WauOJhPmBsegtf1IWnOLgCPFMA0ngrYAFoOmBGdYpnmDc7BB/M1pDicY5rruel
L4hEMIIq3pTw9C496pAuN/46pTPN6jfZJF21O3uvFqbq5BDMp8ye8/NmSvkvs9GoeBo/OToe6Yx8
QFPJgyDK+ADntEpC1pkBabCDBbxofgOjao3lBPnykg0ssgVnkjPXD+AY4qonmzf36dTMM9jkXY+U
s3ATJIx6LVoAMWmEE2cyzU1efHZ4cQP8AxH6c2Oi/tED0oOJs5kojeLHwZilIV3HOtbom3DjLGYt
KcnANjyYjMMAQ10zhLzlq5eCsmfiqIhdxTB0T5jWor5DZL/4IT0a+z1FaPwdWvGSRvXrVMT7cOcA
X3PSn6mFTyNzwRp8muu4TiNo89nH63y9jaRbm4ruvXdag4lHd15hOIo6+omaTgLvKpEYte+QX99y
AdAITs0jCX3AdxUTYqPB1vtZERW4dk8X8FFb01VU5oZMqmCcUKYwhtSZCOWVxNTjF2kcEZUf7gHR
jKvhEhLK3pG4bOjtEea1MwLsa8yz37V4EVED4W3a19INp4OOYrDOE6Evd25UvzH6r+XAxiViFTAj
WZ5/leUu3Orre+TcnToTegiBVOSDEE5yx5OVfPaUnrZXlRw3upXBRnLn9nI+hTL0fF2cHBhfqv7H
ewr9tWRvRVrfd5GOBaNfNvz+k7ZfD778GswmohT4YeYaPEMK9NR67WDDuN0sbBNDrpnMnWO032qw
agOUP54XZz3LrZEG3+nXjOl2ZONN1ewdDwDzvyc6Y8jj4F9A6lPPXvoHFR/O9slXGdxFY+jFkvCa
M8eOSLd3iSSnBo+NgPHLCa6XeQRZDuAMFri3pBsNa7uw79Uq+TqF1HCjA+CxyncUIKYtBXwZUySL
yOEywLFHJQyK73LS74x4EEHHWqZKeWxxVM1sVfuFRH79v4S2z40ew9amEHDAnFeopMyVRivH5E4p
dIW6TMYCB1fF/odkf9B8DTtew9wiKveFMSWai2WZq3Cc5IZtPLAVg/fqJFsaiklGDDUjO1VI/ywO
BSpdnW0EyNY8KG0c763KhymDFdzTgqAuF5reAMvOowUEBd5rftFssfB5CUiXfr2NHkYMyIWYbQGO
NwBb+B/+7xeUPZ1vZFk7Isx/pCuxuhcnidPYJWX+Prn0+EAZV57uAbJ7kmC3jYJ7wGwvenPJPPG0
/q/L1Vk+8k4aUItDwj5YYIGrkM6IoiX/GOvaQ9UT+IHY0wULia7hZXHa51oW9uDLd1i2FJJBWIPr
YUw3iB6ZoqtHwybeJ/njsAABaXdSJyPj4DxQfPFXCA0NvOZhGdYTDWnd+6tBeCUoQiYGcINSu4eM
EnT1HlXujLqQsKoGntZxcZL5MGcUfcdQmX9dlwkL7OldroZjeEmz5DClVRcZ7Jnte3gNh/63dbMx
oChr0aHaJfyxFA+pikgvObjevAnZk85EcNzluv4BQf3tbg2OFXdEYs0aSpfH3eFKBrjBf1K4/S3C
8mAeVQeYYt+y+ZS1qWKvsTHpAQ2DB8NCHeEKJyWjPoS+I63sNEHIL8OLmFSXu7gkpcHx0K8iziHC
CEtbcSMkq1mf7ZiCgq4ZBzMgca4Oa9tVl1Gr7VaY6OEyZAkh72sw7tyIBLNIDv4hbe4wZsRb7smX
1hkl+Cq9zcYCg2QWR5DexGTgZRzUCd6jDCIDd9bG+Duu+Osj8drq4/r02TH0d9gbUHpvZ1jqlZhA
mzG9LZu4DZzdJUlIkFTiHFWbavtSP8WHdvle3VVROROEePPl6Nprmc6fYin4Y00eVQwo1Ghg378q
EwSSnlJDK9l47AOby5D+kKfbUucb43YWpM29dM1CV4T7V5AZaNJqwQQYEjXP+iA36AVvLA2a6PvT
rGkJLxknpafXDrNxfrBHx8VpBymbqooeo45oMl7UeyCFuFFcnTq8j4AK6Zl2JGOpzY3zqspCXYNg
WSLbVAuY4bvIPNAgLag5v2r8+YXWU5uxGj78mbdi8Yo3XJDz5OZHEGaypbxlRQ/lllbMbljhx81C
D8v1P1/fJal1kFoTrY9qD//g9nwKG2dJoMvsHBTC0ksgtkG5tzNdEOywaUhwtysO/yD3X6tT/00D
rnrNixl+FPC8ot2NmG1ZtCrAbIuAY2/vKsZ6vhnSiXpSSUm9pjEYt66OPpduh+bAyX2Mw126J52+
xyFJYi/KVeryJZbrct8bnhCxWQ3yliUVEwhtTr7vGmpRWlMIaVwDBh/w6s49OqJEW2ozUMvgbPgx
MgUS7Aop0Xm2lA74Nh/BG1E0dbvmaRWk9yOaLpXpHpIAiJ2uyAFRJsbIvF2/ofZvnKAef5jB+oTC
ogtgnFY2rYmSitNrg9mk74QdT8FtidAKCODM2Lssa4xc7RSIT+u1X8I8yj583Iubj8UjbZoPyE1N
4m12V+LcNA4jaJz5cO1MSnyCCz6w8Xvj7g2xXIyoqFu2uttmqLAR12vOEIKZPZPqTuOMeAFds0jF
4PjwxYHhmFJgALoVV4OipPi0xMGmJf3HEWMx31loryIiJh7F5uN6cHJoES56qjtpQa/5PrL3rEHF
GGmXtYAiYKT+lZ+YZDeNVW2Fp1IKRZfeRMQ9ht6wsBZT9q6pmF5ktgqS5q9/q5HVEmo8oivq0gGn
rb6O3/mcaG/F0EzctS0+8YzgAIII56n2WUKeRdgY84tNh8uZm6y52Fd6Kehoghwfzxt01nSu11sj
NLuKCL/n4H8ZcofaEkhyUOoRJn6t3U0iuuvWdcbvNqyAWC0RiQeZL7qdjKyNyj2dJgcpOOko++Jh
caB2VZEQe4zr2zUH9xoFY2s6kC7HdHJQ25pFRZBKmWuc8Ln7+G4rhi12A9L4Nct/1Yr4s1B9/HQo
JMbw5O9MBhhrKRw7it2P8S02YLtvmVUA0xsM+PdzhkjUGXwUanPSsXr/brMCu46w5Cz8e1IjinBt
/Tr5pm1gFzDSctAVRYic2RkXnua+FCx0jy/1XfgP0K5E4olfQErsRwrHuRgeMXeG/YwM3af55sfo
F3Sk160t3wbks9KcAgmSnGHx1xXSdd2s2jVach1SlA5kCwcMNuMqwzaXyvroXVaLJT1XK9t6IR9W
PgWn1StjBnK5umrcLqVc5ge0YEg8Gmy+ht17dzcHn96cr++QQgtK101aQrPUh4LBURPLiVBz7KLv
WclVVVGAVTRihAMY8GA6ZKYQGDAeUhKQw5hS4PvhVEMWWGvEL2+SAKNP+svoeEwyslAUwc4hO2aB
nKSDrLLUy+d/UOngdBOuZWOm5L6afUHDtEqVmVzEyu4U15kY6GOgqYWpaSnRgfNFVijBNbPrYaBP
QFaA2JWGJla/wLZgCrmOTfy3AyJY3DoULw6h2suojQUyx74zhQ9C7sGBpTKcsGX5Q6ARtV/KCvso
MQoTPJLYOO1dSCpz+QFjxaovXpBOU42ZpilElZqGuMUTdpz6isQPh5BDntmf9hD7JNZO8hfH7xlM
huA6DxOBP9icHjvyFz7aSSEavYr+simaAS4r3n+kBwU4Yn/3Hmz/XlLwesq7V90IE7iXsOW90H+U
tbougOqXVFDhC5I7sYsxAwS5e52LmPLxAta+YiBWrFCrvJu3oJUUUEEF8LECYmWkhoiiuXGyX62I
+shjKWxmRc8z+tUcx2HgptWwAL5Z8Hb4p7FgFJ3zIBNYD7IfOyK22AfaMo3R/qh1ZnMHoFQA9F/Q
AJzgVi9V54dTviNgYddvslrxcUiumy8kQ/aHCx96RwyN14xcfyE/XgKKYdlnmQnyJCU/KD9blJ+Y
CNbnPiqRGKAdfbbG/2yqGg+y40FIM80HyoHfG8VOHW9Imu77Hw7ISryG5vg9kTGoQ4S93+ALOv0r
7/HufV8rtNq8+G8wEXjr3jvrSIZW3ESdDvVsAhBY+Peg+hfpTzB+g+09kj0S8zdbzkz7/bwgFMJu
5c3GMhklKbUzNk8pT2CLULaYnLSGc3h/hz3KI7SC4yTtP/Xko3RnvAgoZ0rQ5r+QktmqVs9CCRKg
LWjGzIzaCl/n/JOGblWY+6OchUuCErSUZbsr5TukLVguWF2ashZXNN+44Q5QSD2bDY7oFRCAYEyK
WAyqBVqJ7IHfRfjijw7L6bPFMo1DO/DTEY391JF5so5zhARW1mHFq5kvXqPhAaWFCmDN48IEMpKs
6SoVfhmRv67h7OYZBtEUAtproyQAQqk8MDdstYNqF6Der1gpL4q14wZejaIpX953ejphZ3V1olKF
iDHpTWLA9eUvJc/f8BkQHSeFrZL3ZahDPJUHTuL61myz6zPQfvKgIOtsyMe+55RZdIxYkfTjTQQv
UGeqNroog0w+3olbxWdgV/S4d6bwCJAOhWeyv2jehzWS8Jty0XC6AjIgTbHdYdu8W6oaUoSKf00b
vWsUQp7ZIadtm0flG6WwgqfYKzmb++pXPtpd8a27UGDgqTBSSMwpo22ofG7sVIyg3SvrTCwWcppj
ETxRXcBf+VtfYFsmkvp5t9HAQ25zu5frMWM9CpJ7TCVSLyYz728XY/w+CHHsohkMTnxWg2myv2bd
KJuKu0xwslBxC1D/fUIePUfW4FxOdZx+8hlRGOccJBpUhKKNFWLl8puZ2feZsJkYp3s8265w8SSO
oq2uc9Fb8e56vDGkRXTbRXWtLn2q35B6z3+IbdtzmJbEFnWmcpcOiQtRxbImrEA1mObx4SBymoND
FdIprduM+8aQmB8U0+2g8phidf8XzviLjy+7mVFkM4hpiQmDR+Q+MRJ6TTAA29R4EtZuk8KCaPxd
r6qQCe7e7/O4ctD+sWImLXmmQR8fLHNWtTyBthmxpNOfy+Kha7QlYSBNd72Nb5eNHtYMZAA/5kLM
1PPOQrT/vb0SaGXezdu17wkjVbcUVqnKI+z8trXcJL4dcED6uMX03IVIBVd+u1RX5wypk3r/hznE
K440Tz6mg+2pALJPLYIpmk6jWA5/G0rO1S5w4mVqq9GDWNQWMA9D6P5JKhUjf44w54LMg8kpRv9D
dfNUUJb6nlcSgF/QWqfiKbwDe8FEpP+AoK8G1+ZR8EavrzNM7QI/dWiBq6L0ztCDdaXSeeXx7Dgs
NABw9LRSWEaUtb3KKMv0xywzkpIXrin2NBctnFV7RUeQt5YwuB0GwySb+dAZmYpwE4wyvEWlX4+T
UG/BztXwPpC4Xv/lLNUyPOiZBLHbKtYW61VKEapyHuYhfqqyjLikYIv84OhKONMN9GA4v+wK/W7u
RHICsbxabFd54zx9ufbAiOq7aO1UmQZnLoqWhB2lnTcZH8G8LR3Wg55ZwuLVTQHqY+cL3snGmeny
yLwzL9+tEM/kN9JRWUcF67haaY91rids0h393nuUKNNHZ58q5p9VlVNzta8CcbyGL/6MInl+qPYe
4pPvufI4gZVzxBF9yWwlCrC0YWysymhCa0+4dco04HSVfxUytL6Q5UctiI5BzrpcfIbBKu+k4/Jj
XtGtKZOqqsVEe7fA27FlyIY3Qywb64xn+7IzROtphjDzBMIyQHXXsWFAvuUInAF5JGLO1dyWTue0
QJC2WK2ZolBH/MjO3XvZlJWX2nE+rmQYyVvz+y8heOtrMaVS9ZBQnd2bw8l25QismG/0+MJbJrNV
BCy78wMzvrBOOk2VsGI0WaQ4bLT/6kd8pvNGHpeUyuX2DxMsZ7GOdUxWciCuEznHI39rLg8lg2l+
WCRcOtINT4/ALbX8x2OgVuSkHWz6JCH7nXz84ILuoC+FGLXgf42fMcb/tbjATQyiLDPdLeBKxHZh
rZmC52Smpa/aL6HR8rPdZ5klHDef9rOcHgIaJ6orI/qfZUGfwm6mtMjACvDq+tkKIrJnumI69D7/
Xo32hVjMvONt6kHFPauo0a3wiqxx+0Quy82GPbf7TdgqS8dnaUOE3A91V+kMBK4S1IFBgYfct9nT
zsDi/vJPVxH6/xcUuvwXmtpI7SiYlTjSfVB8XU5/ueQKgY8O3HSKj6JFCWSgAj6sM5vnMxlSexum
1884urm2Qzt7rZ4uv/b39/dMvWRi8s6Ax6hifvlJ7of4Z1FPYLkBdl+Fi5XSb5v5qkyz7OoOYLDj
fr6fBFXKU4+ATJ8fu3qU8XvUZRBc9Y4yox0jArwTxtxyOsdSAF094MIY1IVVpGcz4J6eXDMddk2v
AyPQM4THoFGkfuBGGBW5081XJXd3y9Fz4LzmuMxrDBVTRlQYFHeT2GlRbvPNpXNoyoTt1rnwtZyM
UVnD2Gjehda/EVwnFdnI7uXx5oFoH8Oij4Sizzu4ikZQFfBuWv7mBzYbpLa2svO5jArGWlFZatf7
rFSUv6ebRHY/VY+MZ1wz75p43VEEoS6PWdXwbNjNqmMjTu6+/pPiIBhauV0vSBvFjgko1XB0udnv
IiLr8Hbb76dUipUqwpEJlpfs4pj1iq0c4YQ2/7+pQDlsj/l2Bw5Xs7rQ8JX+ZDcSt4PaQUBmVXem
rNd5fgIOVatarFJEeV663b3SS6RapPSdGMWcGLNot2bHB5oplCwXjzZJjmHeKfUrdNN0rpEvjoMK
cvwZogxUY69oGB9QM+Jvx4nya3l8xY6ifb3wpUytb1k/SQ67QGl5lsj6IMXcgLkalpaa25u0R96l
pgfh+cDsTuUA8Nz5HfHvHUp64UQv2T0Lg5nyiVUh3cuNrrnkNuKcgGaxmEioPJOhki/sKuhm6qvd
R89UOS7oBdqwBGy8uMpgaY82T2xhC38SL7poP+Wb449AII7TyB4WrtBpbPU1Ur9V2eyCxN/2u+IP
bu+3u1C3aZ6S3uNkv8vcgQyJ6A/B/PKL8kPKlFbxyf2CzV/fh5O69czwbCypf3n3LbbMqkdgFmoW
htijnAE6/u+wPF27s4hflh6knkefEx0V9mUycvbTLNVpVoy0WdPG+awA6qfdyyaD12FTlLnmLytg
5Iv5KUONZnssQVlosecXvjBAzdVmhc3WtyWc3fFlHasAYH87Duzhq7qH1KeZ25l/7/eAgDXXzaOs
zUXu24MEt1AWHNQrpCgcR2MMqhStgq87qY0CcUksu/SE077P4/fZ2f4/RY6L4+Yj5fBkI6EGeiFf
vo2qI+/Rv3XO3FBzuJdBcUI8FVjN3htLaVWxD+kgNnJZsOsw+JI4a85pf3T1ebxyV9Bgn0h5dEuo
Q3pTQFByvWUQE9tb7bjCCfJDtmLOotcsw6t3ZM1llYBkbCkzQPe1xBNoQkzK0NX+cHOBroGVKhjo
A6GNjxMouCt5FSPg8xWVXLDYu7kyR1RgHMk0aULX3JNcfmn9CvvtDhuvaTNmWjmgYGWi0tHHhjvL
dFumuK9x/4NZ4/LRYozYobuJXoXzbghjpPtOy3lgpC5+n5qc/gSIa4fuhTs0B4/9EWA5aKJjUoXM
ss+SzuitIRsAIFoe0T+E++o4hq12inLMoCZu7KDVb6rFvQuMIAJJf5hMqXsta5bv618p+JrediQB
pvdKIF4M4X+giv1bnl4pFKTUKqi0jtKFDk5sq3JucjwI3scQVFFyMmpppaq2Kuop2SlXXeTwwoq2
6pgWCAmej7aqY99eFQ4t1Kn8sx8es8c2HO+yP4hnLzMOsNnHj2obpiiIpRsQtAWu36wdY78Sl+3Z
sq8la7DjeCyvT+9wB+RKFYrfnSi0zTjtWVqslTYhb5Vv9UuixLkFHfedurFMpf4qGoYaYAZJ7WQ7
vebVsIHvuZhcrjib/xFpDQs2YCcgGbQyXGxvkMlabVR99X6DQD2H2OeYsBN/qLp82yUIYEaP2Oqw
DS6YiFh37dq4mARIYti34/7g0GelWuNTY1m7V55s0OS5IqChAxVIZFipJVfi98tL+NZIQewKPNyQ
G9GjlZ1ol5Q21NddDiXs1vF6txws1Rc01P6znCBwjKoNytg4QbbU4Ibp8ydQXLysnABq5fdj87Vo
tx5/SFbJzefE2I2xAAk4xXwPjRHF//CbpVxXyfJEA1FRHu6XY9aXfWGECS53VdO4vOnpHduO9jTv
sPbuNbHQXVN5AciY9kgGkepiHvrN/uZDESDjCtbECSux3l+vmgB0OLjKVjiONO7jdzE22kChUulr
bq9s7NAjib2reiqb3q96UiLv1WkKklsuIakkKgOwaqGkb8hJzv5DDqDrd9rUdiWwQAJVhOn1Ub37
kX1z3qNNmOwsKO0r/AJf7s8IDcLnQYQbvC1DfHFZCliL5KnVwiusw7i5VokIHl/PzcMf639KiZUJ
Zi88Xr/t9Qu5zLUXoiAy6/vqpGocE8zN2WKZmfjuZwP1Yvsz97oFh3/wo7Rn4QAAK2rZrppRikTP
QH6u0W78847KP/lZT09ShVg3CX3juX/kkkjCIs9wqNvNJb/SXBMWV2q+wEqP60Fh7E0aAmQY+isM
NxWkjnP+pEF8HL0to5htsKd/8TCO9XJGobJ51m08pA3PTgV+w6gqL0D+l3i8H2quqI7VXkgdqX63
dh5FZTijn7ANdrPTLvwpOnE+qAQUmU/ELE/qlYQHn+YK0TGQ8M4SzWXlVkTpVUGf+Fo31mH71JQB
LVFS2hre/YH3ZtfMUFC6TIpuIk4lA7EZnDyiU4GVr6sq5LqiKN/Nh6TUJLkL8Njw/mtAsaGzjjdX
ia89mJzYjxJnNofW/wOmd9oKt3nhva884yWlRSErJgn+RMkHGuFJOShbmPApSppYkxF+CyhyMh2w
1M7AJ3YvJU2n+ZryF2rckPVrH2l9y1ictb5oBvra22mfWJuWdkK1sNKJmfGDUqQCqd34bhiNd1Tf
Xk+VwuybhG8AAkT6bTP7557LyhYzdmWltzaaQ3HU+eJGZQZY3rImShMzfyDtHDUJCqSM7ilnl1NM
HfcAt5Tym6dYQ18J0ci03NmXfBQFKvbHTylz4Vb/5WEdp492BBs9hp3SDgjEab4u8lADdEa9jM34
5808RYVa3tv8DWr+nuwuvxnLXIH2NNec5Frl1FPEFC6pDvWTAeHHz5kh4SrCmnAMftH19dfk34Cs
Cn6h/J8Hgo6Q41tUbe6BM8lJ6NJIWeou+JunIsMbz76ixIIQU83LVtR+OaYxcTWLAY+S/qBXmVL7
x1u6lQViOr+jjPL1i8MdCyunRyWlG8DsXkpXsc+yd/7Z0vynUzIB9919k8x6jux9F0KZuqe1eznp
yFwyav42hjBWhHcOAtQyPKMq3Fr3UtFzA0uZMB9BsOUPCOBmdiJWzB2iQ497H2MfCDJH6gxBVT59
+n2LiHsXWwz/LuFoF3D4gicTeFia07NcAndLvVQ8Vd4Ct/QnWQ/rct5QCIBkg4hcc3apgMLhlhDY
gnXtwsYrSu6I+0YZejSXETc2fP0ct0fiy9Zwu5h4xbtvhLbzJPp+l9nMI9pLd1XQTxEYRi2SqAAm
E0QE3FKDhNsNv1hFk7l2vkDHGtvSM9rucFdluly5G9xld/GHpMCXSTPi/0UsAOcOmmlkINq+I3Hy
7NdIi7nHsIQ2CmsYFYh+7SoUa6sgIMxflawytjEuogTpywFEsRS8w9PXhdz7pS1ZrjJUp1Bvwtaz
ItWbh+hVyOJWTBHZvlWsaoJ4YR+yITnD8pk1KUkqLYWBdldTuGI3IUepMZDeUlVDvaiM7TUv3Rre
dz0IWFqOReIICqNNccHrr0MZyBbRv5XZ7bMy/IcQEB9AOxd4uXghxMdr8wH1ohPggd7MmL3I+2F7
0HkgGyqg2iJvQMMEvQsYowyoPYog3OxJI8nrB68ZIEwLEhRJCDz62P5Es5CL5njNwGmQVlmwXMgN
RXfLsyNhq/fr2L7fyyuh7oTJirdMP6bZjcGvYVeQJX3mVavQG5J1ZYVnLP5HN99XMx5xS/gLMEAd
7N4Gjxnx+QNP4Jb6njXnqjyinqPWMewdMGYmXwYV+3YP8Yknt13Dvj84RaiIEiuY7eBW7l1UFNRj
vL68V9Yt4uwRE+u0FFaHARZWWeuSzQo5etMobuWKW1K1yCbZf6eRhjGtYLeCRbYVopQOjgwv6BFc
x3Tvgm2x6G1q8+V2rSleuK4eN30rLxTJsmyM2/1aPkXm2hA5/pGCtjkVDhh3SSFtdWhgWwkrs2OG
5kmRiVOyzWrS3JTvqYSjpLKKLB0sVDVKVKv5RT6L2yk6dNNe6Qlq30Z9O+Q+isHhkANzO+1MZq+j
gwMZPT1WCme9E8Kka/+2qLCaPJ1CKJbhdhyn/UAtlbfJWDF2wERw8zhpJnKhfW9jOqK0tmJcTcbV
qb4HHQbDvpNcBlxNyr67HzU2tZu3mEizplUWIMAdC3zFmBRV3TAE6nC+d8VfUzXoKvmg2VQ35vbx
BRW6w0tIDbBdPkWjNicUIcC1hnmivwGTp2fVXladBWewLD7c4mGULEKSqBXsSHCLIeW3kk5o6JGa
TiwZfRfVVuqUHfXk/JpCmuLeKl6xja6pmrv/UhIrDgyiQLjU27C8eBY2TMPWKlX3RQz6OamNuxSl
WWZtXFGc3W0UXwtvUiDcN8GMthUkED+H16TBtPG13zTvP9C1BLc+sz0oI67FgKwJmrL3keS2XMWl
stnXlUsbLBvBII+0xVuzpWxCx/FPATU8ltjfY1Lz4uexmUzGVRwQTK9G9vd+FGLFXMw0aYZ2HTqW
kftUGMja8xqMyhBG+iBNTCtv04InwLaU2L18UAv3H3YJ3A++bcMmwcpIHCvC4fkyitwRjwmQmI9w
S/LhRXyE9T6itzQ75624OW5Z2mNU/dP1WHeNXQgFWyyhxQMW1yHi8X6DxPd2nT6M76/HdzldXtb3
IRABGOAnITrFvLq8lMPrbQ9CIg19IWPfAhCsRW/TXU0UJadKcESP7ZyvoSBJlM1XZZ2xxQFRP4qo
9G+wtHGhQiR7LvAF9xsvqiUnTcrFx7CkM62pG6lj4PEra9cgXAzisI9Afb/4jmi6TIBPlnxV9eEK
U1PnSFxDh20qwgupyXDKV848vnojV3j2DW1DVMj2VDjxPm44zPZ8Kf23z24ZlLlbvDySTT95cifY
eBwSWJzFNZLkhm/8SbOaoarcsQEXtWRPXJt13KrrdGtty9JQi03ge8ylIr87WmQUAVw2r6HWDUIB
2LIft372SfdZYxlfoj2JA8SBHnKBH7+O68pYb0aKwUtUA3vG7kzBiaKobHIZAHh3MAHDdDjvQ1z6
KQyhEHwuKyIxNnbXwRN0eUUHG+H3NYxcuxLrRCFlvJswnC55lW1YFAjFQPMumyRijse3tK8x6jC7
WDzpwsOrp4jlN/MO9nYBjZ4L4e/PlOhlYOSasgLSfn/LJq4s/s0k8KOF9gfw06C1VaG2PFYq7A9O
lP9qfyUM5vN42vJdOl8D1BZh1aMFKjgawgTrCcmevLgJnI6y7h2ZuS6HBFv6cozKNfQghO6aZoEx
FpZqR/voP+wjNB7ecXs8joVLV06NojRbwfmmZubm3EtATU/DzwH5hJ4dWJTyZMeluIccSVS0EnSv
3pMy9pPCpMsIyv7e927tTXg1TMEPh17vB3odQXcd8kN9QuiyJYyuS6xBY3RChF5HSMxIgjnaIe+q
BrNCWB8Tg/ab6huRugBRXQCncNFq2jHZpDv5MCObX1IXQdHmOqoTuP+TgFKYNNgWreSD64rc2y7K
SKC1SfCxd55Olqh4rXQqPzTyZR+vbo9UQ+xFAawmRX4qz7nQa8s0jxArKRjuVpRkD/RboaNUtpv7
6kg5CQ7l5n17emigzFFsiJr+PQe6gh5w+8Nu7kaTgFEYWXjEQhIvnxmQMK5ZRr5Cy/HWwfzWlF12
ySk9em4odf3XVZvNf0dDPM+gCYWEpzuKkQ+unnvmHQ20T7YhJvzswA5LI4eUhLfefKmfk6HsHxW3
7n2w2RKYm4r7R/1GrF+gdXk9QPmRwZcAKkRu1RezwM1f5M9bv1XMpBSK6YnQQihjcIh5uqxh8aBz
9oB7W/BXRupuh8QJSjAlYl2UsI/IwVw0iG6/P10n03CkDO6D8Pwrly4qNyE0WoOD845phPNjVZoz
V79q7AWEGJgzjJEAHlA0XySAFIespzMYk+73NrqQR/XHeAD4Pp9+Nc1hSQdv1Oez9fze0F4z9x1X
3errpNS8zwahCpzLKzesi2OfyT1k6qIMy/AOrRoDqzZZlwfl4i0T68pt47Nh38AQKzyvNVpdsh0B
IwOEupwmn1EiBpGIrN4v7WImgG1DqvjHMdn7XtLdrEqYPD31dF9iLBZAYN+SvR205jzOYkp6deNA
nMsCwgAjSw2zYGhGGoKs6WdKXq+IFwHeaiYY8kUHFbkOCNvPA6R9i0G3WssRwc1TzgBFj1UOjNfP
JERBfwmODe8sJZzXhonitBV5pSyOMi6kga6v7bhiZGt2EScnjkQJHLcPWmqkTbc0wyFYgcHkqATK
wkQ9WhoP268U0oLLnxFXuODJ9frOWh+CvgtMTqJD5CD89Zck0/Ngmv5HfwAPAaPRZrelw64G7DDb
TMtXv4JbVyrcaJrkL9cpxbOb+m5GC4jrtWzJL43wAr7jSpH2aEecPQdjxueIoiWFB08zB9wV8dzr
lWp5Tc43l/fiHt3RfjTA2rY69rwFrUA+03Vn0HH+SpEviUD3F+xQP4zmFGxE68hgwhpXnh8NqUrB
7SBP/Hv3lmWRMITom/NhUw5E+yX2dnmHE5dQe9JGu8kdXf5GtJdZvwpnNu87n4ew8B0/lK7MAHfa
ISW2Ygqkj5PDg4LwciUuf8w+sM1twnwWMNJTZ8bTp3L4wKwxuObW7Eybq80yENhbQjp+Uejo8b+0
rTOk9QVUb27DUBbEu1VmcVVjeuhS6UPrK4PMaoJESE4xrYSDrFPz0acCHyV4Ar7g1zWIjrsPa5wG
bqtvuKyxFiygGpPu2bcxd0bb1JVUUX4285kDmWqRQDKs6giC0UWshdWHfb5ud3G3aUINzDhxYEjQ
+vk9cd3LmSMu4Jnu/GEfTDaPZKTMwsHufRYU98+PLJk42nCgVnrWgMU+fKHJEA0gg78KIThrcURl
7CJ+XHK3EXrwwuGk4R2dobzVVojudqqi5zh3lYzUhn4k53RWp8nb/MTnMuezxW5GM4vPqVnKU5kv
t/7ETHcqT8rmCyTD7Bz2vsN8ruW4rjb3LNMofDcnIIHmTw+vQN/VTC/Q1aUajWuYHY6cfpGms7Ju
cLp4F1XlXQcN8U22hDLHOUgM7VV4PVbSX8UY+dG5UuZ5A/N1F+Mz/kqbdw2iWcqlszDNA24EuL2C
8oEgg/BetzKiNoD6sZ5mDjgL8yQP/Vzz7d/9LVzTdhcq8sta0jHMTqR9K3ZhNgdDCbLcgdrBsEnd
ahUW/yVl046ILDnIGR6Z4yLfDRGtZo7aMheUE+Qj3S9tXNdt7kQkwrSZht6qB7y4SCSGBsOdyeuu
w4oWFxHhO+/MBgCoUxdD+k50X1GgjUKU9YL5Gy7g7Yu29ISG7QnQnVVe/+KKit5B5mcp01k4MLpZ
OiQN9q0Ca4Z4ArB798/f3eyZz+f9fhSd08k9tye7swyABhWGW6tEBEpepR4IbuNdhR3NopLXT64k
0LWxl5Wmp5kuZr0FvIiqvMhk8ykYhJGKXJd56h8C6kFEE1rdx/FM8y5O1Z+dlxiof35WaAMNJ6F8
ZwpWUgHnFjVC1lXKTMMyYSYXVh5ZSqJlFdvg4wz4s+9tuwCf9mh/5xaTR5RzqHhdBAGahvGV6rTF
Pct9q30d6LXg9SuDbK1lVNiqh8Zr7xIUEEutW/jWGw3NdzZlFQzKgf0HqfZefkCWNmbLEw/Az5LG
K37qFUhySrNVMjJaGgFeAulw4iP99XQKCqcxaPI7bJmiBumquIEKxLhYxJK76Q/HOvvWdgN0gli6
cB1O12DpdtEpgJX4pgLCrNhBXTS2GiYl/3y9xWdRi1NjA9mfqOo812oooxV03CySex4BEimG2UXJ
GVJR0bXVvY6ros06y9++TH48LFMUwLf0nmpABVry9sli5MGNocqfVbaB/EIykrrpMaqT9ZOAqC6U
WP9XjWmGJL7V9Gj+PHsaEb0z6tdlOtWHU+QQUDzV9ne7SKmTm+6l2oFdeINZW8/DfMkGKSpkf4Mr
jjbrYgRdiIFr+ChnPt2Rs19xwHe/z8zdm/i8rLOVWFM0haQRretf6R4PHjLSoOl3wb319YEHrvkB
Spsvndr6RrgyT1M5jatOaWA03W+Nlj1qFWdXtdlDGU6YqtE//LJjs3e61J+KeQTnqIus2pdVv/1i
S93TFQOZHcbekKfrdyOVQxMr8T5uyuNxVyRZk9O5f9xt8SHTI5hj+QV2vCqTSYC00kOCxKUduW4a
abuwUWt7SaikKsOHws4krE7p9qw5AS/oJVhoASkVaJnNcM1SagXUKq7yTEMqcP6G3/PY2Kkugo+V
RDE5WUwH2z11+v+Dlte8EUxKZ1UE4eXdR+sfidOkSNlota69DM7BtDOcocfmW8QEVo+nwcaUFsuv
miUCVziLftjBCc49lGKHvOM2mdR4Bntx1uAPLmNPDLJ8BvvrPrsRf3RBJ2npdcJP2tqlErQXRcXk
PYR85WdWpplRjbpgYajtIOj1N7mNhxIUY+UCRFy/bylkLq14ZSPFwMCCy1qs7pxKo4I28A5yWmAK
sGDUiS+lZaLLTgQqJdByQQR8SeBhDKsn77d4B27qrfLcLFSiyN8CbF2Ev0+jcNFOzyLX3YxRbuuc
dI3eF7T5My8vIwmAsPu5NiGLvhkbTdEexlR0jiTwMTC8+RgQ9zMQbcW56NaMKfpT1j+JdwsJQurP
TigWC5aGpVguvwclj1JjEvmOR7mDpRBZwq3WoO7OBwjnEd4XZUP3yMwM9SKc6d/ehl6o1ynacDeL
UE/dsyz+ExkJeKFkA7dCCp83BtMUrJKf76x0k0Eon2GyV9IaO7FZ86BretWHW5zXJtwt+Xus5C5O
COjO9EpXopc9LuGwcwCWn6kPZiNGZtYnStNw0pjAo0G25ofqkaCUSuEXZ9CBDrs0/Fna8UXQ2BYI
hL66xQRFrWc6cR2gtjkr6sT1fmhHLfSbSoouFf84JuF9srDUk84PsWXAI7DNEvNUf4TCDDNy1IHR
9ckGp5SLhD4eCn3tgfytG3c43ieMnsQ+2ZWCpkEv5kFNwDcP285AVz5VgF5cl+Wa4T1qy7NzOpL1
r/fOH38tHtpl4DUjzOYAp7MJr/0SSvUsjkQF+G11IZodEh7Ha9mDO+YBO5A3EpstTUFOhP4Z5bfb
/RA8BeaBBOYLqd0XxJFFu4eE29EmC6Rbn2uXHHI3o6155cpM97XM334MXvfE0A73vrjBLGy7u5xy
lou6zur+Vnp57Q/ovKO6W48BtZBOuSa3xgpXwphz6uCdNBbEldb72M+9OJUMQvfYcTHcJuXu9LdN
cM6t03nBd0RSD4TIi/fgT1qVGWiw4ayiGmtx/UWokNCaCNioHS3XWD/159HRxvkRDMY1wpkmI4H8
Km8b046AN0jWjX2/3dKY1dALdYWz/DQ4DwSqhogscESWc57pQwaRL2yjDGSKoK4Lf69lAh0J3fYc
60wya6tyMnENWRo2xuzOCy3vskGokcZa4JxzYqgMHd6sKhZfiya0JCNOk09gZQvhMgLxTtKYp1et
AvPMUqekPP2/rNAIyhbUg7+NMlGdFfx7igVjBE51UdJ1CWcLlPCrOk0y2rEcvOILheE5MaEJagl+
TF3DMJC/r4NFx2N2fWyuNEr//DRbyIGz6Bn9YcKtKR9ybZqV0VZuLEX26u1tK4UuRewdvaL34OWF
zxVxbPNS/7UYYuTms9j4Oy7bNsnSnPFYhKeGK+/vJjNo9O6MVATpJuU5KYUwY1VKxn6J1QgH1KrV
s68r4GeVj3LLSSGKA32V8QkjRbmUDPYIeXFwmaJoLI0x7KDdvZ7iyGwhr9CEcR8uHh8HXS7VZXH/
78W1u74x57wQnJJ6QB6CcOGz8ZMrqrkRAbNuYAVAHV+VC2By8kD3zutUhbqEj1qPxTr6sPli6TvV
siOE8/Ms9qSVMYd0ff9SQclbzCL1IFfjLs1xaYJs/qcySpVtz0yXHyoNObKsMPYQ6kYI6YVj1F3U
wLAJ2Vz6qxiootbtoUhe9a9ldXBhK30ubUoV8DDy1SovXy7t1V1T5NkOW3UxxqyJ66YtgI8rcoNI
zoWBcA7DALBXyMw8E9MS2HmPxT3/94VSrP/rCNb8uSOpDt7m37ZIRO6SQau7QKFvN/6mIQFHl5in
NOXjzagLkqEN8XYOmjflLTq9LC0fBdXL+olBDNGXHopyD9Sz8shlLIzdLRTs4sBhCmGId8QMsB5r
tdPH792EdIUFRC58l2bqt0ZGApaIaexjWp4FeSAqpNjG+EKJgPEd3n27zvkflh8txJ59oPnIT/Xl
Tk1eEwL9nIarWcScBqXPCK2LrB7VraJxcIu5B7ebe/JfiCeHuoRxXEG3KAWpcT6I/YDjtCkTVNOT
qb/SRdhifs1qfF0hENoU0BbX815cpK9kbyNpJJLmPD4KIBiw9DtR5XvZ08dYWO3nIk42g0F5ELas
tXNQFP1h78ycK4eVwd851qK+5EMhWQUbaE5Jf0kaGEuLDvl1PoDHsPsJa9V24AXUQ+n+Nu0Rv1om
zdvJ9aaAkc4GUgfPXtBXYWje8TsnBCb29bf2w2HMyvOijatejZuhgNZEWLnuFTKKNLWelx/vE8Pu
IPWRVhAGiTBlyPb3m7UVHlzxNlfiJWUy2ZJGVeFk0W4vqKU8PuoE+e4RGhdzJzMs4g4B3MKiC4JQ
AiLqoxBQtC2UEDtWS4SNRRH1ibhQocKUXnnte2EYU8/u20Yo0YF0KklK6ev6IybFK1ue8J9RLRn0
K57fzjP/Q8Xe4CHKtPnhcp9oCLpjzQ3TRH8CPjaY+HDwxuZDi8Z8RpLzeDvGtbey3rwJ8xVXwqwy
1nmi2k8F2fLDG2wnifSSEwa3FOlcD5S1TA6HUgn72SxRS8qX7/6pm8oJL/sXu6e9xSPqekhOekHW
YAktrkT7FgFk4lYnh6VSsyVTzr8ucBB4YOj2qDivG8ACW0xtQ60zzPnuGBfAXoSNndgfDuu5GN2S
aLZpQ++sYR4BxKTAYdfWI7q5gA0LBV9WqDHdvoixpiQf96KplAjtyeA6mqzFrBfNhBmdh6w7XXh1
tC8TQhXZORGgdsHorGNTdYwf52WVDQzEZfJzOAVCkTUyR4DOI5vyWaWk2epjfcb00XbIRnJgddBH
QeQYrMHYuzZ050DsS2+VvP9cF+b3AzkJY5Xse1oeqW6TsNECqfflDraLkkGKnsHifD4fQ58fsi4/
Hy0KPhug4hgpuLmpnDso7ozrroejaIRAlilApsbI/b4uM3X+atcA55bymbEXMsJycUd6Cn0pDCZ7
pwZP/WGYX0fNBiiJEoPePc19iN2cY0qkkOiRE4gExWpn6cQu3HC2PkS1TQ5ABkVMnRaaDIzFkvSp
8fHh9IcY5CQ2Lg8J3gG9TmkwQCLcyXgq+bxMmIrSuyfbJTXF0EDBglG6CS5VapKesO/wf4ffd4Op
txwii+cs5IQX61TcxFqq+xfWAxb1aJRPTW89XE6A/SVLpuvKRmWo7b5UABoaPwGiU8jokmRq41Rn
ATplHpCPDXxH8MTxA0nKa9Tw3loa6sF2Xrhw7yz+KWTtL/AIL/qSFL8quUcgHq9A0syfqK6VymKX
FV5buVBl0q2d7He3039PV7PvALaJFMRG3Ww2Xq+Mj+jWkzNQc18JnkDdP2Ex2yEHKkc0peVvDzlS
9OOw09kCWvbRypUYONm+dHgZI9dVMZYnGIqnIFY1UAEbn2iPguv1v/jGcsT9oaiColS3o5Lv5LZT
tVjEdMWP+X16QfKCENgZnqVHfa51CmxkVVm/INXwxhSyfZ+U+WFSkSLLZnTmnX1oNNreZcEwc10U
h6yilg3QMz/SiSUbxf2RZN550oKIVHN3/adgsjYDVmQRO08uQkEyTkO2c1YWW9nYzCKfgv665366
vQgrzr0QwRUwmjwGXcxB7BYPAtENSk1CHbW912z/z63VsB72Zv3ItnrPlKP1WWUSnoUY4QfHBMUh
TaP/tZIu0wrUtl+CGH5/TjwcDYzqaK2ZE5DC77k8uL3UJGZtcfu+xt6D42gJnzuWqqu2/enoGO/3
IK+IWSyAvlYRYM3SbjrCJWY3/I3vGYSEhQA8rBs7m0Kozz6YqD27+YpJqR3DmeCauBMUOKFwjELe
0qVkNtegBBh9yUuHooD1aQYrTXGhUZnOIvichuCVBNs67R93uZJ0ZjFT1h/UGf+PaUpjRhvE/8Pn
pB1Ic6wFEZ1hyKauKuyPkekylUkt731WnkG/5IWeqK/ORHsVsnesMtO4jcCqTuZgw50f/t85ulZP
YxV85XU9wrlxGt9ZJgaNeRc+UNsbjDEIKTQ3+NlbLeq7N3ikumyGu63i4bhGGMoAYGJ14a7E0X8e
khJL6LEaZ+XbxvnDiQFdCVjxkuzRYBKy81YS2yJJt/UXSJ/gqzu+Dz98XidDrc8m45CGeP8SiDu1
F+e8KKjUXuZ/Qte2hMGVB4QJZyNfCAoGHFzrNFI02TYXSYNDOCHlQOu0ZO4ya/nSC/3nlTQ/8qAy
sPiQjVmjkDANgYkxKRstdhtgsAvq/Xv0YnPH4aO7BmuLzMpuEVYnlVsAVkC0GxZMhO1BHF1a0pYr
yz0rwTumA1x+1JqGUu5x0g5gmFLWZsV5gRG/0WMueJhIuJ4PKKd/i+gygECuc4PGvXXWcB8IaIHQ
PaOpZpSeyVWnnmRoCftr7y/WVEfmOfVE0kHpebx7rgFajLIN+il0nyaXFkbcBGMIY6xtPQmNv+rC
x9OWv7cpRm/OpOkK1F8gHjvUxJwuA8DclBlfwgzwm6VLAKuAAp3vI7Ny2AVz4HcBXlg3GmAsJ4+s
WyfhIW8HDyidOR+j4QoW4umou6UeYZpKDGYJ015X/NOtkCF9GLkAZdn4fPQYfXhAykbkAu17vpoY
52pXMTl38czzg37ZM4GwAguOP1m3i6VV7K6Ec0EbbIr4pbkrroXAMVP7oLjvwLrGUibnip6jFZcv
Y4x4ZMjXoEhCwPDCI+d71tDJbb0ZNslADE4evs7ey9RNEpwhk/PtinNCZPF7oDZifar8UfNS53uu
TYfCyoAwgflnvX5sA5g1pQlaamWEPUp6vhMEOKH7kfDz9sxL46z97tXmY2GI7CGkzOCgzw7OcgRf
A/lKEBTYhQyv9ePcoG4iSCrjVzhf+VqCY1DwbCBiTe5gC7j2NBD2nVH+PXYHILJgasKcBIGKy2YV
hToIhbSCzeabdACs5TL4TcG64oU0gcWM8Bqrmgv99v+HBbcoWL/IBp6Lhi1b0qwOm3mU6/1DoGbs
MN23yuREBIWAydDbYYmV7YYAFlXWpynDEodIIGg/LbhOD3ZOVzKb07K9BcH/6lexX0iAt4UfqsFj
F3zXfDk8WWU7gPBdqIvkc3wyv8+KolQp82vwjEG8uUqwKPVvNHjexDvXm9CicLPN3fqCur+5Li5H
TOIAUkSUO647wvtnRoC5fkhUXqT0HEYT5tQL4HUUtAoVLO+pmLOALabWY3nHH8r84r9r4T8um06G
2o9311qZj6PYEF1o8pCwGIXug7iMUIHSsGJhvwoNPYtH8sDRSZs1O08y9DPJjZw53ZzBUQddPoZH
KQ8VRilCymXO3Ei92RNHBtsBXAOU9Ph7w8r6C33Rl24t7wAcOZroiDuv6ykymVmCp0U+FYt2sZh1
DgpFLc4khBGEN+S9pCan5EY7dMLWmboFZArE0eoopdr7Wj0VSm+yKfj2/ugusQQrwUIfVdCUQu8T
LUt+cbhBfvts9WebfV5TFltUlSgBeVBA2qGCWUpwlgNPKnFISgNobcUrOt4skEhl742RfugQrxqw
hQ6ITqALNtan+4DeJQjKXjMe6moMfdXDh/CsaQq0z2eWe/kMuhkh0KbaoTApGEeO03pXeCT7gb/F
IsZeTD+NwDSXDJFPjBsNsiV2IkEUuyEUdIley8QN8ZOvkxZVEtj56o/YSgkzn7stggLUnTEwcqLD
JgGOMAt11vzXSRl+mkxR/0XXg78k/gL9cK0Az6jD8e6P5FdwOqpzeBeyYb0LRR3BhQLz8PlEEMLW
cgXQX14deffvE++Dn5jmIcp4or6lmKlMnhvwePIj0+RVu3WHpbDwPJj98GkOi5RmH3tJvatK5gVQ
wD4p8fCh+TADdlud+3WvkryiwoeYz5fCAoZpa1oPQwkrfFmWJgdIu8RwaPgvqimbmm3v//OVdeVL
tknKmRHit/YGbQ4Gy4TCotz2uTnZ1K51UlF8UNrnUPTWHMXSk60JLDRsXqcx0tsPqQlP0AuGg/5D
wIzXWaiQiK1IWmLl9zw84/vVn6HJ2s+OE9vF5zRR4L84XuQpGVGlS/IUUEX7HDyS3Hd+03xTz1Xt
oa9jxTaqXvxbqT0QAFz9HEDamz98HHBRvBREKrDNu/xlueiWykDUFnT9CMsxY4pxhDFJkWpUzCje
Cc6UYtszM+nb40gOqlRvjSLu1EMh12a/JWvtVX+i9fVwY5H1ILXyRztHEt/iTwXofJwtR76B7idn
godCBCQgegSppPLMpmB2gXBE7kCkHeVLOjVgcV/ZcW5PlZ4UOm6JzzpkUIyeVfm+wqrhYWBbwll8
uSbLqqCjTcoYQPdn0heuTwOKbFo5UIzd4Q4Td+Nil5HhmxAfS2Yba1sqbtLi5wcMp2jzrMqUWeU8
XKza+lZyWI8XH1OVtYeFKWxoeBMbFruiThwgK+ZgeQRfeeXYSsGBJeFbb17EHyxSPi5v5XDDITZv
Pkd45oc6+ZcMSImD1+k+QnKsL00MK4XLH4r19kvSgtALGp3HhNzlvIvLu3U9UI6oqQVgU9VJOl8T
DlhD0tgf3OnHrkJQil9EQybBeTO+Y9z19uiZhi1IoE/kEjAsziRBpBOwFCoOjJe51De5Rw3gBMr6
7qzpK9gB6Y7wnF4Mt/o1WurB4Mvos8ClM5zm6wgVtGQ3PhLV1B/n0zPL1aLd+IF5MOox8OmdTV5K
YlbTuoKYf8IED94APBXrrWnPUhm9gMNnH25bzxynMIJk9rCSxmt9yu2954v8TOH6Ppo/8Lo4fT0w
aHvK9//xxrd7/UixgNqPHevHauvSLIQPDjl6su1bl8h1Fd2Skjm0cz+ASDGDYr85C8Wf0XPlBFbH
tmwGpWFSS7H67Z0lM7/kf2rMasUQ3ZtrpOxRb8yKnMK3P/vhLUINwXaLh3+cPSnmVCO/Ned5so/q
az1tPjy0FS1w0MOtecoEKNzV0EtSW5a6xMB0hrdtsM1MFhf+6zR5SHhhp+sP4P1XO8yubjirL30t
LCrJXl+7b8ZnlDsRZsGa3KTYyUBSc2qPYR45rVOz6tsH8+nytHF4rgP6ZrMu4nlqZ29aCt2CQHU+
x611gaPWcwB96GGM20BcDTwsEoTAWkivSNTaOpNL1ddj4pc3HCIlJQJnjkUyjQZonxWBrO8Xp6kx
eceOY4D1FUSnKi+lFbWipMD3ttZ733RYzoRIWBTxVM+isMjtSQruK73U4gOo3ep9ZFJpq7bpCkRP
Ngj/UeEDw4P4nanQfVeJgoZv7+kgvWGU7HEj8pQDlomf6ToPOrfjz9WdZrQFeV6jeGFR/5jUC71L
Ih2/5G90HxmxOvJhxmtDMdmm2US93KFRgGIVhHGTN0mfiC2u3Ld0cl1398mQTSZcBnaTJBu8FB+z
kNPlQvEPSpOq8h4hXTpuei+GvtGHcfLisEC/xuGDlic1EUGvgcxMFGE1DWSIb6gtOX4ZR3S6ipg3
H3DeJk4AHcSWdAmQ2e7UpDbHtraf80muiDQ3KrrZO35IOEfua8XdzWmWIBsbID5eLUcCkDebHurp
9EekLCwwg4m1A0SkhjvlgD2UzXYw3q9qpsO8VY0Tan6+3//N+F2i/hk2/7LVe4AeSXoBw04ckko4
kCPzzxYGhr7FUCvyB9ZqoXiHma8lMftN03JI4l/K6h6J67VR9HGvTkfSx065GRHNWuRb2/UKNAAb
bxJ+BVMEyWfHdBNqYfb1Frn92439iXj0deZS6RItGAFAAVX6fbBq7kDWmAnG6tasDSCmF8kUEsK7
vgNkI11XxsY8Q14jOPcoqfonoieTAGWB/KL+jz0380imqhtwoxs3Qqmad1Inrm0tYNC5fxRLaqnY
oZfRiifDkVUBAH5bq4JQP35RWqAwVidxAGgjz5UKbCUgZ3rHubjfAShwAUCKstcmcDL0Rj5asbWK
cJ6CjzOVxZWi7VfaaYK7zrX76BQDRbH6e66RrrRklhwjd9hnXcvXbiyoo+LaDThPLfLvE85Aw6kB
Qk/d329NC8LzcrZ6rjzAtFqT7TciTPSSyO2arBQrj4tH/AjIxjf4VAOaoHEMmfewviZ9J0kn5sY1
HIK2ccfEGCPcMOQTv2NwcQlW9mVfxSSrOI3K0jJCbIR3Bp4MWOhdC1z/Ru5xX+HVIWKCE+bma/wE
NtX0dEdhTC8GQxllzyb2WDRgXfAvM05t5Wl8ls/UKUXG3AkGaF5GruldFGzM3hmwG/cjEH+Pj8kw
b4ks97MhlfBseAUo2V7aB2mAIrtZ8aj2praen2lof8FokN/dpMdjF0qYRHiRATRrUy41GpdARohK
84xrO8Ym1HiDbal51G/A7qgFhmRzoM6UQ1a7hOveINLS8Bnc/2J5r2fDS/SywhEyckKzUG8dewYW
yw37JsEzESk519QpwWQseG6li5/6XLjGBzIvYdeaIBYyBlKWfrkwI14alIFRsgKUR3bsMqVQ1mhD
xQx3Qzzl9WPt8Rffs2i0nJn0644FUnTLeQdSO7z7ongAgkvWWhr00kl3Gz5B+6P3RFV/6PuMwLrE
prX1d5TiW76X1+QA0e42w6n5ly+SIHaFz38jL2WGBQqf3HSbQGa7FwPgvnFvUghc4Z1QsrHCsdty
gCwaRvbmZX6LMPXy03JFM+s6Q5LEToSgffYIz++dhptJNxbRuBP60SBcm5TWiWyOM3I6U3kGBSpx
GU0TAnQXC4jSq0aQwWD/6SZz95qg/GDmfAS9XI1tUYcdx/RfhjmFuDhvDzFO8iifIZUsc1B3er1t
n5+Qg8qQfpoXEhwCjFNSc15d3838Chmt/TRX8hukkBAasXKhd4Mg/Yrzt1ZRxXPX4e968Dj5bNGO
n8ywmCF2kpYlW+fw9Qi8w8j+kn9Ql9Wh1efGjYVvqyzF7nEmG2ZTyECU/bRtc0orP2mOfHSbShYu
rbJCMWkGtGvfjM4PDqHY1pkxYZwKX9RPwffi7H9DOuQE/mifCM2MVcQKciSmNITbCYwE0CHAridW
WYTm6h6gU5ZmesbvaSgn/9he62ho/LsfXjyNZ2HPxaCOxp2DRQ0I/vO/17ueb3Qd26mRP7MJf7h1
1HRY5F7EWB10Jd4yM3Or7P27JyXj6fIY3cl4yWeQ6r8dSvq/Oy38vT0/r7fm3ZtSX71MSSDPYBGA
po5DttDObv5+l3nDG177z5hnEaDmnjgNBECwdpd8aVSNnpr61SC9mT1Ureb0SFUoydyIfMWscxOQ
tudqcPasQ+g3frxzVNuzjq2ftBZSEtg+2SRCI0RdZobFdai98iTW7qX+nBYYNptXeKl6f9x/DnpY
0i2DNiOqyhcCUy8M9eymTzMAFByU8koCmQ8xoTBE+esSqOpmn3cSrLjYjUl0VkKIdnCb7l5h9nXT
NQKfLBNh8sNC+vOOb7+FD8wyQZ8awAZeJLc77/RUGysqmLZM2I9JmKy1Pc0Y2eD6IrNS732/LdIM
265ynt4vo+vl2eEZwiav9NAWZeGIu/pbOUprzLyLw21QSIAcAUaXTw06lEnjDJmHFY/Y8xvMJXlC
hs9eUdf1I6uYwNtEFUZ58wXV0HfGPYxikTbhdI3VK+Ma5KVfBj3dXhlPPhUlf2sYAfduEqqp/6bm
YQOETYLKmnMgO6AoLQN5fR4VLwQ/oCtpmLvPlV4ANev5NF7Yg3VKtB7wN1fzh4x9/9P3jxbxFKg0
T8nSr9ObB5SuwMReHnBud5LRt1tEiqIKYXzFKtgIlJ4Qv+Wu/7usGvNbYJCs+tEbi1zxA8cFgPfe
Ik99MTB6fG+q0XmXY/AUslkY5D26gDq1fza5kFgDEFbivbyE4Xfk5VyRRD4fu0m9QP1Nv+ddK7Rs
YmbLe0dBVNwd+kDpoDUU3pFnlYVKXne63rVxW700oExGChRqArlINFGufyOuAgDkMgZZiccXnjKD
ico99aUY6DVaS8VAfFiY3e51453lL85hwBTTyyx0W6kFZfZzS8nNjp2bOA2y3VPdYPv+KtwvfnK2
KirOzJuEjazPTyaG9YUwt/ZH7zk9TKBU4+apPVb8PR9LrOl3j+A2fDYFGFabSPp0+L1zBt+TEiHe
5FnlyQC3D5qIfFpheC/diki+cmD9VSHmixGkhfakYl1qKA6t2PZGXjTiSN8MiHefE1Zi+Rt0z9sm
unb2ha281G55BuACQNYt5b6WdQzAHHByKWi8OtBcgVOp2TTaSJDz0hpLq720Ylh3W8/oqL48YJyB
o7Wg9dgxFUEM4AN1NP9zujSmBX4DD/7q6Sy7PEeivchBoULZIMkWzYaLcPdcl8HMZwTf2t5QLUcb
jWN2icbtggZuCGS5Wfb3sAx+Af1Zt46ieR/GDD1JeCLW2ZrLJcWAfPiKgfW0NG1VOQRls//Y3js1
nsZkDJxu/ksfjFesSDVAExbQ/b6FdwCKrks9q7BlVCciLMPhlxY5pjOy9nvjuLuG9pg2XlVXeElX
V0z9II/0et4ta1OC05BFNO/hQ8XCVrxVbPnf4OvFm7kYBowoD/dZaHG5rj+x9NxWi/HzG/9goElu
eEy+jOZq6iqlQREDd0SF6TGCayjsqRuEAj6ZKJ8k2MtMgPUXOkVpnTpm5iQDthh2UxRKUBscMPWn
Z2l9yf2CjZH8avzV+i1qOvtdYDLOs3FrFCnCxb/6oS9A8b2fjgmu2+ZcXteXqOqxw4YuGLgSL5cR
q0iJxLhIIzwOyRnqryCS3tQuLzBf4Oe0p9X18yRIrFNVJNDAML8xNIWb6t8rUVNCAMvagB+bufXw
SU+/IyYXKR0ilock2WHWOMWNhr9VD3o9TedgiOgdTR8vxg96Q7d0lGRgneWXZx8NvOpzL7E+Cv4U
Zem13cpLWaC78IVLrjGyekse1rdKd6uu1/vBOudkxDAb/KlkLjF4hlogk7dd1Nnqvi37DBUWDt9x
x2cTQY9eOfDPzloabNtt+tus8wU/9xaJMmrgn48nLAsilLllpXA7E9ElyG9LcXZNyZ3BNu+T7mPw
XHaPRoMWqa9UKndDpPKoXosXzJvsqZgWiVYF3zkcJWON/ts3BDDh52J0KiW2zjQpkZEOTqymhu23
AkOmLFbhx7GPaSFDyEuVMLKklSqlnoCQPh7cphvEJ0E6k9jLMB7ysPbRdfgxFE1YDx/0+AD+tQ6W
iGl43SX8zqXWemGPnlwmn3/+vae6mzLIoWQzG+swEnRocVEsZLRP8/7+miySnEBROX7Y6exFD4Bv
xfTv0SKjsbU49xYxtljTZa0Xu748OLL2pSqRzmNPWPRU7BOhE7maGib86epC7Qbj/ztJqiVwnZDs
jB7X5/1W5UAg6ZAkxO50IsI37UplE3XVH9olS68fb3AmNURktja9feBn1M1RGnlRUKwIWYb4gDTs
jId6U0fROhpNXZkG4NaiX8+cK41NdCWZgAdT1WSK8VzP+DZ0RKiUBqOcVD0VLde00FbmbZ3BraS6
IOjt8+hnJ7rWMALNkJtcVbvV0GEwaPL+HBiIur/hLMr/iohxNezT5LT99gCvYss85xwILsp7BLa/
r3y9puWLJI9uqsvRWpYmHTPK3xvILEG2Rd/bZ4aC9/1LvA4a/MfhHQuGYcJcuZ53toIQiP0X/NyA
VtaFebKK1/dxTyoSr6oBXcdvcQcYO4dxeDemirk9DMCVUc97fNVyRwHPNPwyT4sed/45V+8KwZNQ
/zA47CNAQzlUpMtUw8N+/dCGkrk9jYTOpFnJjsuV7KNmbiOsJIzUCiXStZNUeM59olzP/pezmYQG
f5NpoQc4CFIUAfyzuSxectopygb3WDNcQHFf5gTGtVlAB2ZEBfIj8tP+uV7EENjbsdTpFzrpuSVs
Uy4XUYCnFpzMiw1QpssBM2iLfY+0hJvBUi/WF9Cfv03h6ktISwojZT5uS4RbPHa8AKoVfjoSyB+D
LxKfmqivAt7LRW+0yTA3Y/oQ5b4TX72QhdeVhN4HxoKbiBtCz5iuSm90zdgE9NQz9ZfoAHobFi1p
lFnpiqQs3++ubd2by5O1pL6D51iWh/a3smledQ4NL06wVoPFVosP9dTUCdn6HDZwPPOnTj7PJ9d8
DrAq/b3nG3o8y74XnwwK9sH3+kqAz7xtDhNy5MWREdF7g9JkNHjHZ/S3UM+TSESymMBzGjJZgJBv
qstNHVF8UQa5CQ6ua7Smb+jicsEfd161qBMnqiHhLTP7hRXFszhHdXTTC71OvngQJWKdaOLsYYE0
S2A59W5hBiwMnjXpuVRfz+e0JP8C9H1Rsfr6NjkT7xFZ4n21EwXt0wjs8WBjB9MHvfZUL2MYSf8D
1loitIiIVe3D6+Tn78+Fv6YwGnnqfv4dyLlTiDz91zIGWIM1o7FoUOW/kuXVVpWY95XPGUa4CCtf
klL1xb3F/AsW8pvRqgVws+d20UDAXXmFj4a9iDDPCLv65hhHtznyfBtCORu7S6I40f7mOrNuQ9m+
t7/e8p3iI09BPSK9xQ9ihhFvAJIh4mD0X5SXF32M++j2re1pRNIo0mNQmpR7/BxgqXfAK/iotqha
/VdankkGtq+Xu/iPgCyLfMOQ1QXMKSCVkz48XQSdNeM4tevPW0rEsGnNsLLvdl9KRiwqCkHIcHV7
i6F7/hopt+A8onIq60SdYV4lf8+KUy1azWpmsWaHz30fhxe9oVaWmDBq83BS4n7wQFQ8xEv5ktpk
ijP3jo+n3dbgpVlWsRHJC3O2TGry7ekJJVHp7uTBmtlkz2RM4Lwp8zBIHQDcnj6GLv63/gVsWBSl
Clc6K0jtJAnSWgoPj/qXYhv6INhCfdodbLSJJtZUf1lGkoj0s4Wdz7D2dtGqo/SgAJY/rAnloNtG
5a2o0xZQKjoEuLN7rxXxerCo19GhF5swYszGGJI9EgcbbzDnaG4QI3oKZDPQ/qx6nWE/k1jD4HZF
2IQBtVKIcZ5fSpQhbVj+azGfF9Qy4Q3DXnkaMM41VSGsJvCHK7TKafDn0epbHPZk275Y4jgWTVmx
De1INCiTTP2lhAhvH/1c6k7OBE1AmpHnXHbN/VMahujjsZ11ZukqkOFXNB2tBO83Chtk9EMGgh3I
n9jyRqfuZ+NOFJDNHwGvKgKWN6VlygQa7g0fmO/Epq96CXTP2p703b2/OIi/GUe6uW7HNDXO6EAO
wz6TaGQb+jRxwZJ1Kwtphi/Zga1s8Yh25M44m14S/BUu0eHDN6FItHH5ID5STdD1FrN4Z1V8M/4f
CZ62tRY0d2R6SC+qhrliEQwD5fW8nkZMko4d5rAanOzK/qmVC2V4TnYNhGM7w6z5tRl5zSVwOtO3
dyMEGKWN4Hm8ootAZILKSPKBp/c/7RvPAKJ1+wL3d+VKZLgCoJE95MOe8182oiq2zoaaTPbDwV8l
keLGt0h6jQ0KVS6+9Q0lEF0xmaq3vY4XMIvVKxtghGAl28OwLGi6Wus8M06L0crj3icx2sFPvQf2
bq6eBh0yEpqQvzEBQkABa2NfW4EQ6MGfzUUslBvVXj6GoT8rhKzOWdD+3tmaSS12RF6X4AzUd1D7
UCwA+fm6opOgKWEvwHUdtco2EDUhTHrHXjsS96NA9yFrLJO55f8rgr+P8VXwxNaGYwXdOxd73wXZ
cZAZgodRes5k5dQaPGpXciZDSKgCdWTpUg5UomXPBPsQ5ZE70UiGUTBPMDSOuj2H/mThdjyvXT+6
UQsPvszyLfvf59+f0Alwdegw3aNUd/NA0gLEDf1pXYPkrP4oqJEqehKvJsWAsAWHtX1elmy/fj8S
pQB9D4ltd8TTcDzV84GrjLX+eaEaAPVyYKiUMRh/fnRrSzpjpkUkkkR+AX2ht/voY5IoOE/bsnfP
I/YTeyZKXU5aqVh1M2eeUSHVF5y/bbmXn306XhVYlf35EuqxA5PbIyxvfQ7rOyGXERMWdXoCV2II
slbdG/vtwst1pOC6U5XU5ym6MjD+jH00jCrLkD6ZATiChZXFhG+XVdKo8FLYzZB72UFs1nfo1sOr
Nw1J1iqiRYwnIcQ1yYuzwOop+CJ5/qUIB4tbEhSt7gLhv303DD+VTfS5oedidQl1IEyLShFQfNOW
YYrAyfON6P+7OJw8vFJGkmyxj/42J66lm5WqcQMGwzwM37yW4V9yd7lN54MW4T1LBG7b1ycOs+9a
R18iT5VmofgDpdy2vblZyv0Gg/BVPEwV3bN9O7OoXIgC/AgGuUxa1qGy8P34WNkmMBlIkH3YFkbJ
OrwGLZB2ggH3tCJUs1iHA3ORvfdy5ULEHWJCHuQIDQxzFYtgo8Q0oACRBOgf4NBTkuolSNKFaM28
VT4jZwY6XUg5hDaTsU0BtJVYr0z6CLSv/O/FVj3zs4cAqQI0KlPyfRA7zaoZG9OQV7E3tUl5cuxH
Z8SbHHma2SujWtr0SMyXda7fJ1W8SO2u63ybg8uQF48OBwWhwqCyM6EXsWvVTgDQkwSsReZuM6N0
/j4vZSWvABJ70AXJGUfrkX1oifT0VCMqLydvJqe4U7SWtLEJGLo3R2ooxRVVp0/D6KAAL83w1jPU
/w+gnQtASLzbuNJPktP+SOi28IasG7b0FqWus/402jiXQWL+21GEWPGFU4xodIIbyiVqFhkY/MG6
Xx0d3fa55V/HxW5bbFHbBXkeLb1NUm0VMiVM73j/s+3atyiWHeEV+52uQDwNCq3s8JogYmFULSvx
+sniATQmXjxKdbv3xnEUDDJxCuph4SEAEl/gqnwpG8r1XLNftKJMNNkKQRPLMsiMnp2LpK2WqlUs
7EzKHlp41HXxmhYgo2xv7vb9Qvs7NWFjGBujqMIrBG7l7x9Vsd+R3yXiSPU0LGJgtYywA5BTLdwQ
8bfBvyFqQVdm5QTSs7DjZwWaUQD7hgi8aCco5hY0JfnGhcSGOCoO+TqGNW5nB0wojQeZbxQF74EI
Nt+bUeFchbQonD0QFxAZ0qVIPJNC1j9O9ylUOrQnxwAxtHz+Mk0ND0f6xBCla95OIU542Hz/3Acj
U8hfZ0sTeJxocXQKXkVDHjXD35uLsvWDjK4Z51QffSvg/Crzu4jwpwSDRHwdZpBg4/LBba4rlf92
FkJQP0uaxDgjE5Z/U3158gV13pswaHQOnYuWWZ+cI2MDun5oRInzB3zxOMgo8oLA9ViWFJyQYyWY
CAupqq+bZ9qrQgolrREIYl9C/Tbn/044Pe+SLrobloqme1289LrrFYr0JyZFUFeOc3AyzON9YhhH
rPSOOimM7UCc0A4oQ0m4k78saVJ1ZgpFxzZhE2XmbYhWovj8dGy8NnEW7oJMR/jQAVlo5crJ24T6
yAhxrWWMNB1OdwmG9MQSKeXenOgsCt3Vo3XdVRnsZsYmRm8Kx5LL+W4KT4/NSGQ9JEuLSp+YAM20
WR2KXrwUhTUMbjPfbJeKQP0PZFlji/cmQG275JzRB63dUThVYAwePzWUag3VjQ3ONMXvL7OOHprQ
UKBcQIDTs1Op/jmL4pSC6M0z0d9CoeToaebp7ywcYvHnjBG7KxFk7g2uBNtHOSsrQuoays668yFp
Nyokm5U5RCfjY+Equ/7Qq9K+f9DOVOBw3hXyCeKMMKcMPquJ4Y04SiyyIMJ8tq26P6ayK8C11b8R
TsNCiahno0Z8VgnriQzfT+laqUiepb9sfoWmZnocQiv1oNEJhCrSIfXUZRvM9/GlRZZpwc8SDBeC
e2Hc6SmI3MYm9g5BD3z17umiei244wJqqRSF4onZ1i1cR7S/lM9GRkKYeaedAMDwRh6B+vZzIpO4
DwXK3S6clSkhfMJYvZEf39MTZLl5U8lyPGu1Mqji4l3GZC9Rauh7SGHOtmAu2kWG8pYM3ZmgtCKB
BPprD8UmHp0az8JQ2Ke69CA4/xY5RPA0/6vH+dcPw/U27eAC1Bul6b8/6I+jvJ19zycaeXvd0h0M
0MMi1P9EnWZcMXKKwreWYMSejJEJglofD6SPhyAZ3TeC0tUv45seDe1goND0KvQg/aJn0cf5Zgce
oEAXWWX4spik1BPoZYzGsLFKEbv5tT7/B6ykj2Pp06j+Ley6SUjlfi0uD5f+7aUHspfdRYSKWNdY
cR0enBo6J5/EpXzVVobpUzW6ONVnDAU2MtFtmmBzaVfUx25Zb1QYKyNWTEzPYCprtFAyo35Doikk
6sUgxXt0QYOmlznxxXwQU6ejdg7iCO31d+klQ0QbH181eie6ufKNcALz4m3IFy7i0lsrVGrsYgoU
WkEjkVYsAESBb7Tr0skBVwzWgietjuUF7bjAQMAZfBAavFoTX30ffeSe/dqjXBT1zfnPCigcQwOY
HYyUSkelrmoORU1EBbFUsxUwM9a3EznL3lFFl6aivG9JKK1+lPXcBpnkdt8UEHNZz48nzmGn0yfH
bJhNDdr8aqJNDBnW23vXmK99YRR78Vpt5JNne+D0r98gRtwoLyMOpGgTTu3qXIAtVY+C/fXclHQM
VuYSk3sx71lB6hxbX15gBBn9Uk0P91doTNwU1UwelWn0tNHn3vGKNX9hFLAJUwsBHCFvB9UUviGD
z8tPo1O/YsjczGTd7uYYvaBBruWuhPbk9ynwsSU9D67+jtRRJUqJHCLOT+kLP6zePokn3mKQorYt
B+w0iCUXqC8Uwxs1e2uJCmzGLZwDBALjPkUKccUOWG6CQKEYVlVwEQi7MXPgN7hZl9FDQPJcJJeP
OXvXV4dB4OxS2jKM/mJbJzZn2qokQUov+n3Gt+aIISD/RIy5NIGZVFC3XbmC+zRdm5pxLC8Px9Z4
1+iyl3w9eM9uZqvOTmfSIm3PHvg2x8HlfydD2ZBIQik+bNjTVoiu+nY34RvwUoYOr0jqLEPoWqib
WuoTDMG9j6c2NRYHycZRuE+9d2ED0wiFxaBJf1YIzfVPz8M45v2wherdD6AHianf2MRNGRAOC0RP
eVG4vzK6C4wBcI6wICt7XIw6/kggDduhOVagAMuC9iNS9wwaj4AT/uFLHZwj8sZctyyJph66R9ji
lJwHPgNNyVp14jpWWgL7zEWxZu8FV2oWPITBE+Gpo8OcYNVFG56/BgmnzHJF7F8C/41k2MsTD3Fm
yfltYTxynnD0jypzYZcZSRCP9WSChLaWkPcleHb4Ajc+yNK3UUTpSAVMHTKv6dNeUY8UEYyinXva
IoxxREDWbLP2TBXH9IsdN9QV+NjIhh/aJI+FECVlZ8sz0SGIePq1unImD3gMYZcL2N6vlh3bKViH
zBTp+DLBVJ91w4sHik4hQZ1Z8+ThgCqLd7SFZ++FpY8WHcyIyzCTgRTaZoVSW1a7uaiaLLJ1/LNE
tVZtASD5iEGYEUsYQOHmcNs7ojmA6LZYKS2T3/21yBouDO36iTMS46JopCR2JNiLj7tF5Th55wIc
pn2uAguL6EJkesy+PSkXA661biGnN5ygTCotuowEqCZakUCjsdP2D8C3ePc+n4dK+dkOkxeU2mkI
v/PTLMSUunzwBlFwuw7gxHzE34nUQn3YyFRz/vM0swZorGnZKqKpyTbOzIJBatp3LUwD3XKu+pR7
xydhBFfyCNlWD/t+vGebbE0FJCiYK0RXsWjrZTaqv38ckyymjZsIjix2vXCucAx+x7H6M916GlCS
rORpDrK/LSY+pYzYMlxECMUHFMd0Bfds7yqz25sdSUnRn1/T5kDB5Cupmofv+wDn4Nl4iqYeIs0Y
GKr1ALxbA3HmN4TgB3797KyXQQm3HHNxC5RPrAHyC6Cn74yzrFqEiZFF8rT0MRrK0L/JNpeA9k+2
EFRianEsmda32gdWyXhUE3WAGqTZI8FM7Wkfh6Ld1kAp16tnhmU8l/2+7keTCy82s5oXICaEDOKC
xxiCybO4tjOokS9IJcoZTM5o8xZOpxzyo+ah9CRf1JRUUeDH55w4mq88SRAxFES40iQlZqa3rjUO
5SB/xHWLp4+hpK5YuQR6xJTAP/Q/eJkTdgDwFfhqq59Yxh9djdCSaeqs7/KwsmQsVnHzhewEjdnx
eCKrwuFyELIhfPoDfVsgp3QIcw7upxTdevmuaj7A1D00k8/nHI2AEG4uVt7YYO/l0BvbuRhsos9O
u0e8vV2oL5kYS2866T9w+kx2cZbGAHQWtAl1GLHU++Ji26IsVCtM8ctpLjzCdVdbh+5fGNcANmXY
zQ6hLgXt94OM3z9M9WBZNmfEm7GERmOT5TGxeiwBDBnx5k2dpkRXbq/7teiECBAHgZz5po3ERTi5
Uevj5BFgRPg0sl6fPZkVee83ATyzd7znZZNyUn8N0m63uSnK64dwOdD3bEec9B7ru0z0rejWW7l9
v/RXgu97A7eYnrIs01F7Gb6oIincKhhMB94Uc0x/yT+6xLiiOteYrscwTq4nllbqNWmxdLSAdoq0
+RzkLauF9gIzFegHIz09bW+tdYGF/K10QloXxPbT/WoYvgULgNdaAaeIPDYxSHE6McImdURuJRjZ
H/Fs6l12CAunhbMGIuFjkCbnDA06cKkf16Epy5enJbqb5jW6j1fPBC/H9a3M3pUHn6B2I7Atr8NL
vl/0h5Av3vICCrUh0yGRDmYIZJSiuA9sWHcNTklPMp/+qeDhDM5kW6i9T1cachitGUiLBPUBEReQ
3Od2oi7KSVaS+drK/jRjabdlNIWZmB9GXezx+BqfI3Kh5qJhVRLseYwibtt1uz+KWoT3CzezUE1+
n7bXtjhY+7ySdrnkrSkueaVWcE8Yw26jhFJ3PMN9svRPw69pFK81Qp1RyD9pmGqo3UNrNfj+l6fG
jQi2lTTwkv3A5pfunOY4K9N1iifcHg+ru/2NLNNWG8vSHwVlG8vD+NpC5n3GY8zSgAAWdK+ao24p
VGSPcXbriLb0Mpw2fxsCZmtXwDv6D8q5Zwpu2eEkCV1HxQ7H5sY5nY4/69R2DO1IuRHjQj33myjE
56AFRwiW+fU3T+nRV0hhVbZ7foZ4pbFahj8FbnUjIj5jz/MK3VUycpo/qgQDYdxZz3BUPRLHSz36
bhZThOJa4WW7jQX07cAWU86nkdom/E6s9quLGFFZDP8m6lML13uKtPw4b/6QkFwb+SgNsZXB+diH
sdIyrDoAdbh8Rrj2jPGkRoLtzSaE1bwyzwp0XiIAJxscZ+O/ipF+TQGlvx813dgpJf/GXaZZHnmm
+hd3O5u+2oZo7od5kS8aqAasgTDLl1Pp8YPtajDm1IoYzc0vxAKjdMSUEDQsXjc41d/8SamAQXA9
fb55aQpdDWvcwKK3t2JtEqiqnx4pkn6kPc0rxGqXe8U3EfhKMdA3Q2zur/FjXFgpL8Ozvf1u9Zdu
DK9LaGsYZ9tgVXHq++ruAJuqz51KdPpYMy6MeKQNb/TQ+KNwq/2onGeTMD1LGUDpiezDrQ1gFNRW
/i/290FOyrM3meYCpgyxJNuukddIDX1cszFrEArQtduAqIHO0wsb3TfB5s2JCOAtjzl0m1u9VVZF
J6CN8WNRoiKJtMyL6lsAkun7SUa5PSOgYYsi1AQgD4FsXHnlwiF2P7pjIdn43HYK09KLlWYAuyLZ
88bUX6xdD9Q4jfYJMw9Bm280cbqYx9RzWmuhPUrU7uZgphUzvGzevBo1QEQCYuMfM6b5iee+1SbI
p5mQX52QPjoQTcZYEribkn+fIfOf8+XJkylLTFYFyoAfvq9QbZs3mSsjYJdJ2ElRtkWT/rDymAIF
1T99LgNj+XD64NFzH5Syi+PVdEGknWNE6trpZL2U434pqmmQR3Mlu1S2yV5JccqafChKS/rNIJgl
51F6wMaVQX9WLQml+pT3pgCHDV1wWafKBPY+yAlLuBgpKgnVcan7BLC2IszhVvA7nUsmi0BwDUyv
fzSfxlB25z1CLLNetgOErIzoevHJpZltoxWkVzhRm3qXWi0mtIk3Waoix2YecN2WujfkWXanqsTJ
bHC5rEuwORzP9xN5snVg/Etg2cx23tZdmV5R9O5nSkeu94i+pfhBH+81x15wjs4uy40lnct8zR8r
38nbNeNO/DAhnefbVc3/Wr22CxkKD1qYzwAlSTUmvBklstAj/WZJ/bCJ6cSKiwcwsULcESF+Kq+t
ZR0Rd+SpAlBK2U45n1Hc/92BLMiHl9KaRFgp0fnVWb+aBU67B+RwB4SYPiRbtUWcdkXmZA8EZ+XS
gT5bpbQk4+13MXAXOQYD7xtMEwsc6ZlX7YmDzFD8D35VgMO54lQ37ddxy/mYgSQFqfHgP22Kd0xM
Oijzf0uqT7HbeyZHf8p6CqaxoFI/KqUcsxi6glZWocIA66/fhdAXzAv8bWBf2uIP0LzBLJbDFJa/
lGnDECu6oGDA6jWrUB9DHKsuciWWpMTXphCYSMpDELZDuYKnnYXkVcaCsLOgAXZIb8FjyEhPlxlt
o2pEmWYNUHpPDu76YxNJDG+ChcxSS5VmKW7+J4GjLvoGWlsEwFUEFyZ42xUZ+VfvHvJ8/jK4IMkk
Fx2N0WfCl8IRjjeoHVxD9wQOgBZ6aps5gMXJhEVG/7/cZYJiE6iLM4/7TS/zqTQD6DcyqayWk6Kp
MsKcr90xGlnlaD1b+psx9RTHbqEQJOuxHPkdRdcWDnxy3gGkRuLG3AS3PPwU3+hXjwfB2GJD2oUT
eqliJZ+k6j3h5PCs/27FaClgJE+whCV5/4ByrjtZW8qSsCEizbiAIxOXG6OPAQ5wHjzZzvUVJjx2
uvgBGkspUCGNMiszKNIEJiG1jd5xSIHZGptKsTpUncGnPkircM6nvGlvKbH4CNkZooG/fwdcuLz/
t0GuFCzGWMtnmYNxe6Qobn01aw9tX8cJ/GRVDx6HLH2QcHctb5qQA1PvFTEejhFVcVoDHLUOEKX+
3GJ9Gt0z63YDiWgYbTbev0EH+I5j28QjFHIgwVJQ6h0rzXy9IjiEgjxOJSzK5i+IGqmYoyzR9H8L
dKlowZTf/TryGjLGB5JiG0Q6QK5dB3t19IhmMF8m6P13/aPwUhNeHZZt94KaV+EnJaQXHwBy1Btt
YK8oDHeO0Idb94n72QA3tuPOopVNrQknbV0lrWXju7Bh+5gXa/uUaO8v+pshVnrUbGjadgU0vXqv
+NPvE8iwaPFOjAzyMtoxZnvOP9kL7BAFOLqjcvRtrKqSnSH1otDl/bqSP3KRGcjm68FxT0XGGjwM
mgdnDC7/XT7UyFl8PdrCbVCLG2+zcUNGH+ClX2l584zD9NXMNLZOG6PKzb9QCpYgyY3sFRsUt4vg
9MggMpqdn71/PQ3UmixsGQ+ZLWkB7I/r9x5geQqYPvnet+++MMX1PoCBrGc4f/+zZ9b43sDLFyHq
hPTf3vI0P0knZhQgi8ZjsiqzOf+thRnzZLOPlKtPTpnsrlxHAwevSrch/ZFoAZL7bbPXDQPuBtrh
0n5ORh9ugN2sPdzvFidY0U6Qgwvkjyx3V5Y8d7xLcBm0jbRgIx7P6XKw3RV4WckIpzYB9/6KHHok
c1RTIdgUbuluawp/AgPifOZm/KC/v6r0mEsI6ON/tIRplv3stqc8+79hj+k8OMxj3AUdJYFpucOA
X1W4C7O5OuGjZuA8zS8zYLq7UNROJ7pgHWibrKu60Wrm7dBsF1lYOcGM+d4r2Fq5ThPKcPx4S/cM
PJq7B2MWk7o7nDEr4EbsMgh0uNr49Xhf14CVDpztB/8yPEXPFP3aua3WrTKN5z0qrD7QKwveqbbm
kg6Y1tJbxTu0pvRm8neQa4Sey9xs4SdDYtaIk2SP7pD1gYHOhClJ/NV1mTLXO8ByiAWIU3HDliPi
qv051Q9R1CXl6uWjQ719yaebS+NNcpcaXdtt/eTvrBFmZbDVhHes9n5Y4gFjkCZ8b3kWSBwfpoAy
Ha/snuCZJc1poXdOq0nFjenrXGkMYxcILcqRdbLcT+vm+g3Xu2SIzBmNomgba18A29SDmdf+I2MY
XmrOghYv4ht1JdGCdtpEWUPBBU5djdKv6k8AbfFmvyZ+k57Vhpa7eSpDW6Itn6N31Qx80/XjZYfY
QQewKhM/nGK3PDhp3ZdhvJDMpU9d5r1sErEBftVXKkDxAS8yEWKtXbQQPkG2hIdH6NjtTaeKiSiy
zSpfBV3/xUIBuR0rK6opK4u7ctCDshKH0kgjzdObmfoSsoQvr3nBL3V7UTCSg4DmtOjRKo/1Wgyg
sscGY5BvjFg61UdKy9KkebwJmEh3RKCjCZDpzXJJ+VHqTMnpnNqjuXhl+fERyTGOF+7PiE/Rn2I2
VGCf4wCnrCsiEfr7DsynGBp0MmNTeBRbsUCQVwO2EbVmWLF2Hn0HkrGgmsn45KmJzdEVw0+FBLIK
tIjdZ2jh9RGVHPMV9OrZ07HPaU4u658HvL3G3iiAaRT6L636n6Xxl0Wc+odg/7HUguga6nWUo+NT
ZZD9oivSRIU/2yY8wm0DUZnJBX7lVU8FXotiB+LC3ofY1jHul/JJNqYU2fvSHZ+awpEqB8KZgLav
rmQoLiU6ninWQNmw4dsGIeemL/NDPFD88IDP1aa7k0WlsZEJnwcmHwbTnM8GxsVQhebfBbKDxQM0
4JfbdMlfiw6EBVDpZ+9artYGkINqyirovqYIYeObRPEy7jTAXJBdMb+xwpFOKXP/g7qpZZaNZSHY
bRj2Y9qZwVRB+v1W+Gh80QLKiQPhuK+wW3a5sAgBFP6LrYWkoIfkKsWbb0z7pZjm+QKAG1gP7gWM
A9qcibNv6sN8ItiHqFuj1/J+ixV6oJMRoLdjIOUI/cPJP7XLOhETCWuWmPWuoZQLpflp1CwNehZk
S/INejyAT/FmYRaEVCSy94TCRfySbJaAFfshvqvScWfK3U4pCfjop9tblex8T34kr/4NRYIRAXn0
snAP/GRJhIBx5eCUaGCyl+sFMOSLAgcdSJ2Bl6Xf3VtPehQulnmr1+PKbW/izN6h5DHF0JGyTI7R
m+d6R5FbcZnF6mf0HOFqDmYJqtljafC/EN2luX52MEs4PqgdH0bBK0oMmqEoJYUVFDrGbHcsG+12
L4BPH2W77hQbLXll1JCSswAgZmiNMVNtdCPJsX7WCGa37Sg9q/aq9KMcvd7Ml35XnigEdOG+Wjyn
TG0FTaK8LH8BiUUDAqXKvlpOJKDz7apDlcUfdG2A9tbFeGhU2hgv7mV0RsQhHCeDsFAhsR9Mrr7s
JejEel8XAFhJm8DwTLhBYVwv449BlM3zm5yPqf7btOhQ1yiUk9dDOSDcBi30cNhXhZi+DtK6AD8x
1IZns9NUFbisPHXfcoXIxjLXw4vblFQBb1vtvS6H1m2j6JIWQndy0PzaN10dL9Rh1BZysFqTaQHf
0MFwjUa23ayMi6dnCvAjWfKVCz2co9U+GOtUrL+5ksIEVkWAhj5Xd0pLknukyZiPSr5iMxELlAK1
1v+MMoPIjUWgVL6cYt6W7QPgaM+OeAJ/MPmarho4fHza8doLtJKRsV9zLA4JUZ1HNRkG1pUFyBUX
e27QE9y+oi0s0VmhfWKnVUK4dxIAcvV3vy6F4lDZwEJ6NTFC047K8mlqvz9DVP+UylW4jSWSniMM
uqTCOSonvm8Oc1HufM5j+1iqTfTku0Y6NUy3MKhK2JH7K1mJKe3wK/qVhRtG/BF2huTfPxxsNdFA
0LgRVKfmfpiDMN/evoOxtQggplykqs2HNUDrFHIJw+QvNrFiNkUBc93m9cUkFhFhYQ4TjSS84WG1
WqBXry9r7gAfNIgPKQz4l50c6YWEz1QJpeCFrlUGiWFuXhJEjKE/CR60Q8UwYz83S/3vA3IiaCzS
K2sPJQUOTcuqaOQPzMHNKkErZSxvgzgxlQz5jpHQ/CNcaznkG/31uZsQpeDmogZ3hma8+wwYjzM3
skewQirYyMnnF/6PyaBgESR/1eQ48HEKwcIHnF1+u+ZUUedRV6gvq4Utk993CA1In8z+geNL65Cc
en4gELsOnU4ru/uocsm2b1eSEP+fa5Ozt7kaq9kHKnWY5h+PCQ/wxkcpn1MsfE749HVZmKfYsLP9
kPbq4F0KDlRVwNOhh9tYUMjL5LynVQLnxqGDhNtZb3z2F39+E5ho56OlcGHhsbGtxtONmLqev9Rb
G99y0qlAewsYpt60+rg+dK2y1jWHpAb32tYvuXDOVkwbl028NFq2glKtL//JpadwcFffM6+ICq8L
fYOpBs4ncs9WdpcP2PE1g5qZ1XhL1AjLdf02rqOvQMlYScFVnYwUdv0Lahx87o+ZWperWR088/sH
ZYku95zBSa5DgTPYPDyJVQr+VWx63fvUavtVE39VsuhFxlU0CJtS2zIAMJB7vbrFj3QvnoHIc80R
jEL63u0fJVe2PJTkZSu0vIkMoSC/fccXWoVkY3o52LcCdOsLzLJr6NjeHJeMc/lqYoufGpuih/Ah
fPI059k+tFZpjwedNxdqZjmGgPRs2/VmvGO2BEoVh+N84J6YIlLPBI6YVVHGQ4r45R8khuTRMf4j
UEP7H3p1zycQOWtW0wQ9/rRKK/j4XkGccJkTDNK/FOMq3jz2pUSz45ek3ua6p8reWzUiM2SgSjhk
6rr5v0EajspNsWKi8TJyzkJvfR+DX4u+yu+uOKFaSyIMl7/hrSVI+xgDW32vjDcMNErY8K86ic8j
XV71LVM3G4jma7Gubm+8lFn14vGgXdNSsnv2R1GGVDlqeLsbT/dnAVgUZwTsAjX7N6g/zhaOS4gg
wXKOGBcGMtjyfnm8sajJ8cvRk/9e1OWU5i090QkhlLgCXMBXCRiOmyE2sbGZ1onChBudnJ/ALcrN
PDUJYCWYzioPrHes7XR9NXl1pUyMFqZSJqBsn7INo12rPSnYAAh2aEIGdpPJ79Kx27WIuYbnh68i
3vH+RTnaLU4iXSJof8zKO9zFCgkRpA47tNfjMzRao016nnm7Q/2R3PyYFBTGT5seKve2FMjGHc+8
09vhbelg6vGigqy2MEz14wAbNiBktsH8494VAjhYXFgn2HLNZ2Y07IeJ/Lz+P3QRuVwamNkgkKI0
JXYPpYER1WG3HwYPxku9c4sM/dmhwL90VcYh2Gw7sLvQMm5t4Oq3b4FJExX67IXmTH/fPLTek+Qx
AYMTfQvK5TUYqUazFzuu/sioxk3Elh99fJFEn4a6taazvybuI02lCgOwKoS4COLtdY1zXNvF67Cv
9Uvj7JGXCbQWCRb2mvzc+tMduTg4+cifduTpDDgIMphQwsH74DmBiy7hGGpdFZgLHf7OWIbw1lCe
Oj/pgiq57nLuISbQPZ57qhcY96AduqaAyKNEIhLly2rvM4AUrE6QaBXzzDp+0gF0PdMXrZUouv7/
1yghd1GrDJgV7BFkhrGZIxgdjdmUthGucvDyGlBGm0B5ZqSUwgW4lOZYOgqxB/bQf3t06QiT6Fnc
sgv6XveLT10skUPKmP3eSHaQJUhH3I8wMZB05ODAZJEUGT1QMYr8lxrrSkm3lMnoS15Fxw1cxODA
/fI0/p9t9Us8NivpeVy6xOb9JYRBfH5qERyX7YT/bgG6VHLNBc32CTIOSFC4UuKDzNLd2cetW//d
goIRXOJ/Va0c9m9uSQ15GoQzIjAKAmEk4ZtUmGYvwSecu44sMK1VFjYS0QlZ2HLshkmO1mJssx1d
ZzwTDmrFt8EtyJIsaioDTQpV39ypyTUJqvv7POhyp7c9abosuMWf61gRPl2pKdOKna3cgRpHKtW7
hJSjmFVIxSfO2L9tuNoK1lxcEh8APZcUbpdiCFMfF1WqFKjB9n6JqgrNcDF/k1Zt0Bkgw+ivo131
Tq+lf4EhkT0AcXv0CIGpbmgYiqXyTLXJ8n/fpQ9pQEuEvbSq+e2pcGOo3ZOSDZ8bPpNTz8n69Hbo
hGTBiwck8L6DfB6nKDS56z5PAg+LckPrzZujokFlFAD+kd0Ek66PneuVlRkRphMg0V/x+yhlmkgW
4i5IOOMkqlCWZXJ9fTxhhimnM4sbwxkvczbGWdBqfmVBPbgEgbuNshsEdPaKiAYJwSqleYPvRofH
iDNRVTqmr40u9/bYs3qNlwc/liqD04mj/OJjNmMxCnl9Pt8S9jMO2F8y+r16TDdyqW4fhdKBAY1N
HPKY28Lkq316zNt8LIau2DNJZMq82z5KbsJAvHSWkIq5mdnfbnNhQ8PQGsTBXVJT21+lWJmlcRTh
/QNDW0mj8Qw9WEbz62pEuUbCkJ94BNr0uKQ2Im4RCSBAn+vHV+7NA7lNzFixKTe5dzxE/Hig7fLq
OedcEZPKy9Hp/buRqec38wFPAo1Qw98rMas1cyGa5iYn4XwJD6x48oWo2TU51uxLRGQ9Jxrtdi1x
BBoiYuf0fZ+gWIq1IkPWITa+JxPLC2VzI6xQrQ3MRF02t+ETMrkhGOeiwSTLuv6Fqz/nqPiK5VEU
uzipJrSVwdvQUwMNtdAi2KIFiSruF3bgzIea3NIOQIq6t7YLxbhPHD3FD1LfLjpLKuoxmlu/hVvt
YJYrkjyXoN9/1RqzMrHRJkJzpAPnN2agTUMSLhNutgI3FsNFUltcVMAONjNhGLj9S5h/9Lq0Wwbv
CyJAHhC1E7UVX5gV97KSYwdHHPfY37Ddr9zxgamtoOI0qYvjg07IMuxjCBV8i3WhaOi3T9fHO9C0
e6/AcyzukUD8uwFM3RvT4KZ7Jhfjex33iwJwGWXK2UPYEGeT9p+6eBT3GsAMZsZq4Xefj0uJwSz6
x+K4qjst31q80nRsXzyPGtwxOtI+HOyV+R1SlEOFxU+6I89FHh5HN3c34/MEtIjOXVVe6+0qtOi9
yuUIQmDnEHPeL11270O5msr4VyXG/FdR3+WzwKYLvn+eooUoSaFPVhbFIVwx9YrMFYHCWuMLX/LC
wxDF9YzWarfee4J7YlJYhFvPPnQlPD7vPI3XE40KO41+80vTg1CxgitMh7Cez9LULc4OgGFD3D/N
engaeWXdzMZmRz7KETKDZQzZ6pplA6/80RANi9t4Pp9IvWo7sFkno/KYl93YBW5MZDVclmThVTGA
Re7AvlCAVNHPyg03mu9gMT9jR3MJZ48F8Vgj41C0b4W2cab8Xm9vWRBAuI4vQRohOryXBiNyIf/9
A1KvoiKRWbwaUawRjUxifmnzKCu3PXfDkl1swVC7QOoq7RIYcfyEu0ZlWl5Ygbwu3LbIEYVY9Xfd
tME7jA5mnXXw26+CkgwgRuKXSU5CGWmz75mY+fomLwsz5u48xkHRQs0DOhuRSBWv/E6sxbK779hY
E5D92gYADztbf93eqkQFpyg57y6Q5cm5jU7nxYmOB3Qqj42uehc2gGOgd0GhjhXeXGdqMtyG6Gcf
uTuMRqsH8NazmBfDi9DIXMEQIj8JgIYfvy37d8gZ8VRRLA0y3f96V1P+6dcaDG9BBpxM+UzOUagC
HxO4TKmbreuKDvmQ531c9cg/m37XC7xZEluVILmA1RK7egE+dgEOFKFh8V08Ofw5u/K6kZkmdtEd
cNquFPctNvwkayWVP6x2YP66KTnHI1XDGe/3YAZjEuKGMbbHS1XG4nHnCRc7XDGBrwSSgPxZtJEz
2K19tr6fZqSZA9e7ZO2fZE9WS122yoMTigGMXguHhviJlYFVGQjvhATDbN9MWeD7OOkPzpvOqYnX
W8yewpI3BLPFASTuhMbj8mJrlg75P7tbayRnVnCfdUyT9CPo7w7PzGSD7KJXlicOv9we4F9NYfjI
d9NPird64CHluecu6sORftLMNvLH/n0I3n8zhn7cX+bpbfNm/qhXHrCW7Xs8r+QLBSEMekfmiN5L
D99ImVer1Hl7OPXr9WuPpXtyNx6GSmi85EDrUemPyTunXHvRroV/zScTIPInEsco8ZTa3BqIdsHi
Sue/ZJ8IidS0wa1RvEzDCrJzWwHzYeRIdNWWdgOehpvAgVENONj9KuNpnMDc8EE5eVxNH4v6MuTk
uNnGOGMmLTaXrkhDiTPgEVpTFDxfopR32UH8PH7jB8ZoBK+ahVay9rGWT4H7QHiE2cfQqqq0UMtT
e4OwxlFHwlA6rKOqUGVj8WIScLrLR4UoHSwZMH3XgG7J0hmwv3c+Pmx5FYKywuE5WotZB4tYTzoa
R4S8+RAJys5AvQiRiMGj4cczvfh2jEE9+i6+ZlXhVJxGwVY1pXKNmv0+YdklRjup2BzMl5iG64k7
8hiwrIUChusGT4CQdDR083icAYvVBrly7YXNp5F/DWhiPXSl0VtcFzOAeGUl52cYeAOOBHlKB+LB
VjDmPBFESNIkx2j6d5Va4rg0+Xfx9xXzFJAJml8mk9v83zFTPELxOJzqdDAV5m5++BPONeYser5Y
OAQbK1YnSAmB2pQI4wPXM4ctMIyXwknb+DZfy1/WIkdodC4dceJutyJtwLZfsjZAfKlCMlb+pGU5
z8zW5YowpU2ySBr4/yHOtGmhrnb3GDT0ydD2zhEXZsMvUHE5wsPI7EPHXInTr9fhTxerpWtW4nbW
si94YspwAyDThNExGipU88UyEzH57PZJwC0bq6r8Gzun7ScZbPrePy1RZvy2swZtFEm4LHvSzB2O
Q/VWy7eJJgMitnPl40BQ23uB2bV07iGEvn3vS8VbgyYsRhWgNbEdugYCsKdmZ4M0go+qMyxrKnei
blSxv1mCl2e8M2o7K1eLeXS5JITutIB+CkaU5SWN57i0yCfynNViXw9L9fi9Yk9RGHLk0l0E9LyE
qfClupU+BoXquwlz/xp4NpgZ8MEjWON8SXfu/03m8mDHkSGfDWvWgJK/S9a4nllzSsRw18FnXz/9
cNamyweBrg3yceBlwVNa6cNdQtR8dTUscBWUeL+FaONk3C6HnELD+d3ztuIZKObiPt3xn9abNdUj
SN8H+ZHqSOSu8tp25fi6APENae/d8hJe5P61TC19jBTLvjK1A+QXZZwtsKmyyMKxyU96VWKkH3i5
1yExtG9hbMuLMTxRitFr/FNHHe0JjRTEQWLVoBjuJO/PZxtxALC5phfw9cj9lZzONI1xjSzHkQF4
fbGDO0DdH0ukwBzg7GpZRUAdHOE4gVNjrBIBQ+vKj/rbfQPUmGHD60Cxmeo/vgzfFZHz/I+E/mY5
nCwLxFwF/4q1by6QS99+dQRfwjb5L7gVpsS7PEDEY1/dXcRBJd7DkO94tUGPf5m2tJTmSPW4/6RI
GHtNibEA2j4mOgyezi68bxNrI8y7S4MjyHlAVxXQ5TrQNYxKWGtQnX26dgQvatxPfXNSB1D3E7OX
rwj+6HMZDtJw9U9LQavp29AeyvidjDwETC/1bhcUPayM23HRmfenH9150D60gaUHCB40bwBB4Bjd
3OL+JEWaGzxoLZT7oti1uft/bwfdqKMECjVc4WBIhva1cOot2q498LpG57qNLHNmDHzuMPnukkx2
A+0RF2FIjnIXy5gIKrXFT8m82qSNNXl44yf7AAjHf9bKqCAFmPkJjyKQns5hrkJJ+B8kOvnBPzme
rbLBCMG+xZ52H4FmgP8LsT3gtjIQCgV1t34XbGGuxjBBhktIGZlS1R27X7Oh/pSGQCUjQkU63b5E
JjaIeqYvHOD9om4Vik9nASLGk5FukmSBOP3DEv0a0GFxf+felT0MsdifaPM1jsl/fgn4navSfkuW
y6NW2+dKVbo7p6QmfKLfim4FM5TY6i6/WuPimTN/78AN7CTOaIXPbuwFT1627o7B8EJWl5D84iZQ
gMK/dZxc8RIIssCDICfPYZ8Olc704X8LqFnKeySC30yaKXtkbiCYKcn/qB09bvWuQBhSfoBsgFED
8IJTr5eYhgS9SOpizCVB8SnlQBp4/E/KyK8ps3TOcIEWxV0v2+2D1BZXEySmslE58/HGEG9292EM
FuN7/Khe3kJWu8+HpeMROXe7sUIfiigSDac15n5AbJ58/30VIgbn3CkAsfCxkwBH6kCG6JIISULJ
BQ9IRdCCH8NP2gj4xaIBz6T90Bzi+C0o03aCIRoDENtxwAHE7BI0aJqz2aup/KbKrf0LO3CE0/Pf
1eQ+wDqAHRmKJXhWosJ1ZXnDpes1F4pxK6SYRJOSqbW1ccDor07KX7pVnZ/fzqi78s24WxyFY8+J
gjRi6+tMGcUqERTwQ88Mky2dott0VcQokqmgcFNKOnpTJX91yC29XXrp7v5NkvDHwz/R8FAX3B0P
QwJos3MDTDjkL9getXKs104ZTD//SiLD1vVZwcUQ4vuUJsrsuml7jw79gRX0IQLGBmTiTfiel30R
jcUFhqnJReQCabfOQHLk8vGGzerPZZsMmmjVAynlSK2aki6Iua952tKhMQTbEaOBOI9yRhC0/6hS
6SdpOTdn/d1//m8VQmuhNKgSMvomgrc279fHjWg8RdymTuGfrsZgGzPtZ6no5achbuUri2cvJJro
WRaxZjud//8g1kqWDMjL4RCx1Nj8tZd+cjm9uZXzZpCLSfnlf3PFlL/T180vw/RrsGcqz49/7TAv
277d/QRgAp3JPFC3G8iaDL1/6Sc7uGsQrXuinT0NcHYLOZzJtvbToEvbPggFRDqLKzEvIIq1bzLt
uebfCZqUHPHDMsanVE57sWPRhzC5MhgGHnJqLrlJHA5LEaa5V8kCaf2axEYnEIk5ADsRhNkQHMpR
foH7hH+Mi64KzOkfHZxPc3AiSU4AOMbVd1uHvp+NL8CNlZt/l61/jkdAa5BnG/ZJ9ZLIX0DgmXJC
Im7OSOFK4mSx4YihBcN9pdn5hkbgXPQaGVy71cROj5DFopmQojxiwTKWDwDj5Pldr4AZUvOoDGsk
pA9ByP43kHBYW4Jm2OtIBPS2s61I0kxTRQ1C+ven7iS2weyrSiy+19iH2QZOjzd4R9wHnFvhVDmw
VG1J+DVrmCuFFhzZqEYEWKcxdUezE3VWv15EmigEuc8IFVowmiYFV5JISs0C9AB+RQhiOLPlYf4D
Nzu/QvtBN7fc8hUngbwFfyP31/eeORjJlNRc9FW3Qo7QSNLyTh2oAdCld4pOilH+oj2ZpQltm8zQ
NwXldHFJiimCHwVOKzfJzc4SBCzyW7GpMvTbNe++HEu1mnOgGMRzqauteX3y911QkedMlgfPfOCc
xQefZbBbwJRCShtd9OPYLmU8j/CIwhF+4Yh35Ktb5nWE+Av1z8w+yxM6Pdcl5kn2x7LemcEt0thD
v62rZ020ACZW2EFuucl+oFDG+B6/BdAcp05FeRVCRPnjXZ+TwxArjKIuhYY00wZXrrxbdii/G7WS
DrwlzwGvoLlSMyHsiE2n9y5zeOQQkB0KlVIjLe6E+KcJvBGF4U68HpvS913uM6xeq9lpneXsSmE2
8jzFsqcjmEYKlLMIV3UVatlj488xkjohd2fMcrhXu/YxQ2AtIc5SZYFvdnll9puOWcQaPEOWWFrL
bOhMfaWhhu4tBtvQeKTe4CfpvufXh5GaoVvM3WJD5icmeuhOnViS0e+pSZkJpH6AzkEHo8YE9mog
TWV/zyrGbz9uAS8PE43sff4y+vFm1OUm28vKMoQyE/PoqPuVQ3waA0fB7YhTD4Ykq94TxamvcEOg
zPQQzVnKbmXJRFyANCTQG490bsnwzi3Dd3Hhg3THQalZ0ctT+Nz2BgdiBuMl8C8/SFjSojEC56az
7uPqdzLC7Zr7OaQfZpvcXQ3+0+KjIBOqAfX5n8UUNsKxwJwtkLJ2lZIQiuHZiPuPJW3NhSN6evAW
FRkH60ZI+hynijHrKOAOttArh//o0yBzsl5rVkXRO64Jh8j4ORluU5Ede45qkkG4mTEV6BRKIN5z
JNHecHHzTk7IbJG9iTgHntBzdR2Ja6x307UMvt0Zrx1vrSaHfkXjvQMJacjMIHWddveH+Dtk8SoV
XZN6xkejbgaeJXl6ZopP+Yx4cgWD5qPjph+UMkUbeI2BFJW49cttvRj/RXLKp0730N33OyAOopXd
amklP/VBqQuRvzqtHtw23FCnt6o89gwjgDihvVWNqf6t+FpqX3XNCC0m0E05LU/ZKI+JT4D3oY89
D8zqenLHRScLrE23SUVgW5DdtiQFuFecoQYwcHrmMbvbhOWSHyafJ6eCJpH9S8I8OvH+K0QBTh8J
byxAF4yS+j/FeyibNIQxidyAWI4szwBhB238ZeLr5vxGznsWiqpSAbFDKwT6W+nKKH3LM+qL9Uvc
sDjLSIo+gcHq+sdxuVyBQUFsuRS8MKEFoL9YgRWLqZRV+bxDil9urKRd+0brLZ267aWMnVuLe83K
3V1KIX0GfJWmum9tc0QinKcG8afJ0JKMvec4aflxYobu+ZcMeythK9ac+3dOydqWSKaQATQOlak3
+tZQdF555srOynP0O9bpmTaaazfpslSEZDjaQo5hj1dB2MingS3VsTQ2vURs0cqOY2RI9JmfOY18
cgUH/8sybGqZ2S0YXQ37dvC/NRpBFW1ZaDdIOnUuqDp4hadAHMcidW74VxVcKNx0axHhiYZFWkko
xlOeiB/8/cTzZXbYzTrp6mfX2xMc3z2gV3zJGXFAnmKlye//ThTfefI0W6/Pffu21LDfxXou+Kfw
2JmDeO3L6fC2SYrbJ09GjVp8EfCn3MQt7pSGaQZnAdmM34Xoo5k/fTFqE+IH56V+2Uvcm0PIrYnt
m+ARZXjY8hBWJVfzfQStMu4iV7UZwCc37IpOceJrf5S3ttZyJBbIC/sdBVMpLYMcLeQKV95Qsn74
c5RjjFtIMGEn48HLvKYsH1SIV0xj+mlcM0xTfgT3EjTFVa/XT9hcJQ/JwWPHu/WXEkdfXcxwJsF3
oPoMQkTWDd/r495ZNbyapwAezvuTL7kVUjL6coYDxO9L3kOrAeguf8ihdWW5WshFG6JY3UbMkv8z
VrBz1dAkggIURANkme18FgrTQqjC9wxi4XXo6AdsWg7rA/Id7pyGi2UKe7+m2FFmF1oqfTl/lUgp
fIcsKZ7Wbhqypyk2X6Yk0GKXqcljbLkGVlymNYxH29RTy52Gn6Sel4CmqqRMXdTpBuPFPKf2yDnV
3XWED8RlxFP8bZ1GuEQn4FAtrG969+morExmQzActagjlWwkpUAclzSXpsBGkbFnzYcAVeBlSxT5
7XPqKvicN1rOPIQqDl9cx+i3Oxkb4ZLKDZKAzaFhkyrESH79thJVvrPLl05dseKQ3N620tDyB2lq
P/bV7r5lsewwWb38rXoWGdpYfjgIM3q73Q2O+wqfsZA5kogu75wdfOUIVZjuEnBdrh3pyAp+t1U7
4olcbvzkalpxS6xk7pAgFRoX/z2rGWFXUIrYJN0WMbmg9zv1ii+Wl6LlX6DU5Ib1Jp1CEfjoYToe
gAyHpmA7rXhD2g2o1cdk3mtvdkwTUfiGPtDA6/TB9Xpxw4khD81n2w6sZrdJdaC37ifrC2sqQ7DX
LSAQ/LoqQi4Iy3pZRrm3PDyZJCG1fgFT4F0wQYgcVQ12Qv3qY/aBXWfSEfe3HfqCJ2mkh4utrSwf
bDSnduDWO2vUenvfN42qK52n2XF2hghv9Zqkdwjkat2H1x/RvR0HVO6CawG7Alh/xBxmFeJ8OHGt
e3pczT2P7Vmcmesgi4kGIN2fOmSPktI1Jol3/J+Bo5a/caKiVwBHUBZ/S/R902QsS7t5a13LIkuc
650EShRCi5Vimu77mqZexNE7AzPwioHEyNpAL0vHTSV6JQ3DTYltZBZa6qgtsiFQzhg9tFBxvqTX
JjQBBXoAc2LLJ1fgxOvxhJ018HyDEY/R8vkdJf7ynbjlLdd51IqOjVCbE1KYC2M84pzoN5xHQMwq
T31vCdHamxJ2RIkVH5rIvlzCvwjUaTthvBUgOmWdd2LElBDM4FctEHPcUprZnT2dHN4qrG9FzpJ/
RsJBohDcjgcs7v+McThDbyMl7PECqHKQ1ndROKqiMy+YuUhPKuFdWymEldqELt9OdGEZ0pT1pOvk
Ouz/iXz9HR9wRlZqCrEcnLN29wdYJ503OJzL4xwdxOwMidD9s0NQV7ImYvvBwQxnAQ6UjkgkhUbi
0SUvWxz8hlevFCAVd2XwH7c2M4VeWQrv59WAhocqDm9epNQN4n+d8ZQ1r7uS6lQxLKwk1QhVq2tw
gYyVhWz3W8HeFfISA0DUUrsVSXm5FgUHGznKGu7MiImiZ6Xw1MHd5oaxsECEsFT14C92EZRtOOFm
rzVx/gpHBC4lxBYKP7hyLVwNis4Ulp7Ut9+AcHJcn+anUtlWGykcjAcXBMIs21UFVPIfHqGShUHD
bOzgN+fqx0TsRTyMlJOruGUTms0aqEi+3hsUA+PYknIJi0I7B9WKzFKqjXGfalvlbAHOO1acAG0b
VpboNag098dQPFYYbRRapzLhNeHVOSCLcfCK+R9ilpm8/FWMKvb6j8ko5P0dCnBulBRJRi33Q0Ga
P2IQaLIzrom3qoK/GwuuDP6pmUrmOLfyVR+GagvxqXcFtJRTjaR5s8zHWfGPDEtDUlPb7LXuLYQg
jvgGAAy1saR9v5fOAlnWdC0ZAW+dWEmBhkKjMjpaU8n1RnFAxrf9OeUWWDChSZfIzeouzXOx9mIa
NRoslhJr2TbrqRS4KgCpgofnUz6V9EaJe3LeIhhABJxat4f1kaTf/1oSYCVKSspTMilq6e9PJoV/
X4eUsJYqzql8SrS79JJQt8HMlCF1wpiYVftjJeRUxhI1SUouceI2jGWQb/7II97KPpBTV8gOikHD
V4zK8zhm6/oCCLetOcYaTbRpSDGqjvCioxoIvsyHxS8LDE9PON3c8UphYLSCc4sVDjgve1/NnCIA
RamQvHjX0QMoPhbh6YSrp6Lj/7sHhz772t/ltuq4X8C6lzltJgnQ8Xn+AgPyOP0TRGEl6jTRDh+c
r084OYETPXvSqRW82lY0DlFzJkm1USvJ5uXIh0p1+T+sboaT8Kd0wso759dK6vNESzZRr4Hh/ciG
tIoXH2iZi5nZbYjLkL/40scUbWiLMk+4y8KInPYd2T2Lm22rIXIRPdAKw4p5J07yTAcHkrct6pZn
4MZseWBBmOstfFtthaHfdsW4XtQTDNw+G3YX8EMvQ8LvCQK63AVX1G6myTa7FqTIotK0144pSDre
HMT/ULuKPdulzU9pDO/QLOjysg+dXdEi9VWWwOv6yB5IyQmot/DIyEZFpmfdCKV1fS8AKhZObPQa
/lVi+14uNtFG2Ca8YUw5IhWDgeQLqXHtkB0DfU2P/pIaqqxIT+GBWInaxdBO1ElAmRjavcHeHaAH
a5BPKAGco/wWK6rYLsnyafLkJ5JZBnaVdLNKdpoxNE8FtwZzgE7+fnbqXakbsOFbQeGulZ53UA8A
iTVGmDKr3/HScBT68wKIn3oxtxJspguqtnO7GYg3UQIGYr0fuTfr1Ov3VwSNunpty+qOdgV66bNi
49KEMxfkY2Tms5Pb5SdVO6e7BoO3QI4VuG/R5PU90iKqVa8nJWXDs890ozlN5zicMYblBpbQoEXC
Vmd8SIRFVFEDPf2qAM0jF8KNlpMohDOg5fTSt6Fk18NDI3K7HqZ0uswoSrIU90ESoHX1rJMjkbfP
mUyKCuDjqkW8XqkUncK6WrA+4YeDfxZ00t7bPSAWWRk7gD8DEnFBZK+gI9z6QMd/KdOPyuzuRTpx
AWuT8E4kHd8w7/IyjZTbJDoelEvs2jXTE5SYb5PfBL+D8msSqnD4nn3L+lW3K0/RnqoEsAQeHHZe
44GX9IB5/2arvN/8KDjyseMAwukZlTEGD6o1Tzrn248AB9MMyDRScJmTRo9BNo63ETFBMjKeLdZm
CNJccdBB9RZz6pWWegJz33RdkxXK2Ws1sI5AibBxEUOrfKwNabkXYporM4ZKqlj9WIwUI6bDe7Q/
hCUSBj+CG7biOB8f2st6PWWTfAbej8eeU7onEkN9SZCHIc1gUnmJ7aht/TOjkoxqcMqsG3c3TzE8
NNNIaIaEWNpxTLxCstp1CVhKQq5vVjTU5FvNXFCcKXC1me4X+XAJZASCgScRae14UBCAxHzNf4k0
Ia/Qdq6ZkS+kpkxI33RnWwvi0QyKI7xRg8ybUqxIa4oL9ZM6Mhee16MA9je65Nqjc+2GE82KKRk3
S9dbkHv5MUqWrEiqt2q8iPAoGuUjQAC+1dzjfsUUVE+oKCwcSuKyfUCG3jGs7OTRpyvgYn0zdIoH
GpuMYTictd1hiOnucqWgilcWqIY2dvOsz9ICdwzUfJ/2ZJhl4+Db70tCe+LvE3s7kpbg/ZTWA0Gp
0xivv9KU1aWM465XoYllb5szQIlzOFPotTHIkXAZ6tCs07MVBU6UbnxmAn2G0rbAzAxQCeN3yJc7
TVq97YHY6R2TGp5xl7yRrij0JF3ENoqigC1ofqAicPA+wOdRegoNsYDKVF/IHJl7dTrZY/01gBzp
iUsLQ8/FzG/Fnj4QClzwXOciznmvh2UAeR0uqnTliwW47EvcHDnsDYhiawlnPhIweG4S/zgmHNrX
vo9edLLMmkUbcggtKjFBuuXCqnBfJhjfD//SqRiVLLy7J6MLpN2ewC6JoRwhqdrZuBRUhPFaoW8a
B7WTYHWjio4sd0LysaVYSybrrgMcyrYaA1GM7DQdHLp87lVi1gOD81Urk/+cNHH5Akul9MwWNfXb
c5Xx0SNsai2zuPEnDd9kPvFFJvM1x6Q6+yakWq4q3H8KDAj+jaRhH4+aqFmnp621Xl788hKnBTFc
yFtTd+hHk9AobRWcN95VgtOT9qRd63LDl9FiT4sMT1peMBvRrBinFZvafbtROCYf2VAERMqoYjL9
XOL6R+stYRBfx07f6emjpwE1sFICvDo7IJIu15m0hvQLwctXnAP6Ef7+SS7NAAOf/h2z0PMfNl9f
rZUHsYlrfETHmI0Er6eAhF8wZzzvyM3d+ix4vJv6Pfasw8WuOFq1JeWX9GyvMeqv7q+FDqyhvZja
1O4zEKz75aWWatOV4YA5jkeEWXNXuZu/TDokEjiXI2cFMNIKoD0yP2L5ZGHRnagkJJYJj8XkRADI
HeqK3GxrQkiFbGnIVonooAT/tKLbbGUVbUEhLMsKE9OJAnZrqKJOkt9IUB/fItbZjL9RDvJnVZac
G/K122OMoDssT/saGYNLoaP5Un6u2S3LasRbDZYpY13TS62NTVw5bAuLAhu1KAIVO0h8iB8X+piZ
mPIrO7yDbLZrACkmDGdrSJjgM6C/6uVEBRpGB7nJfl/8jvuiebAMOP0bwH/75tTdOgSvnzFo+AWr
myjo00XUQDD9Uy22cvDVPHLGVTkMfs67elGFzpQuDnqylnZU+EQB27gF/MyVbCImE4ui6eLibhVW
OkNEbEDna7Y/j3Jx4+GgCGXo7GMCBeflBTRaRpIGqKnhC511OZR3batXDNNpL/uFaBBSFIK1mvKT
DN9ncJPil30NrK3lpAmRLc77ff/tNirZRCwgR9ckAaG4HG1Cio+I0FngWChXEq9gBkEPDlVuVdqv
RD88X29GgUvAFaf5Jf+wiUXLMobsA9VJZE94ZsjJStI9qT9Pl7TjmIS2wCwrTlJwfHIKyvqWkldL
7AU4qbNQpYHqYf+Ly4tb34sgZxfGPZPY+lPHQEiDq/POa6DCyACpAVlzMiPAz4mBdbXWHFJCfXtD
0NMS3r4HOT+dy9XDmRcrHgSCEmwCha3RhLo7aKTD/KlIyW1NBJjgiNdS86Ms08+lu7Ph5fXA8yBj
W1cXxW8XQHKws+ViH1UtaQceDMZp1Ii5SmjQoU/pqyy0hQsN2wMOTYiIZiyfyQWxa6uMr1h7CKw1
iSxqEmwH+sAnqkKqNNnr6Zt/XRjnj0hiRNhEN0oEPpRL5Y8uNit2N1HmwVsPGaUO5JHhWqlxXsIR
NOE2oZKLAQhNtDONyXeQJQ7WohkL4c8aSf0V/ctXxjZWG8IwJToGgfklpo+Q8/qrKc2C3qs9wlYz
C3baQi1fgmpEmd/nm0022KyslRgKrtZlEq2H2KVt4E81FKgqyBV828RvG2uERiMTNCnfVVDhFNgx
n6rw5FGIPSI6a7hpnLLerU412iDNHC8TYDuP5HEDUMz+bsfrmZVqAt6E3rOJt9oKn85KHuJyoT0M
aHbZ1z3icMioJee8YQJ2y3EoB5Zdnh8Bfmvoq0legyKkSWa8tMiP3VeDX2/1x3zTMbjqt1pn8wPv
W/A84aSGdlgIYbx0TlrDCUmJdTmsi+KsEx/R70TsQiXXOn3aF0j/sjsZk0p4xTVqEsF+Jyvgghf3
AoCm1/Gm7dEl76YR9VsT9ek8jUMAP7F3uBJxOh6LFFD3lR/gpEDKX3i+yidCr/PZcAJw74KqPtlE
9SnJlmupFp+3IY8LWZ/Kh+2ft1b5z+hdgbIhgKuwTPRxxWKMKX99UKukIe8Cr3+1wwh1zKNICOoa
TVXG8QCONs12Z66Umnzw/HAMWrmiKHvWaEWCjV1+iwyBnJR8Ta1zDFW2pYRP2cKBdmWeqePwf/An
6cFgciMTRH9mfXUBrU+ttyQmS+PtUMwnUogZFDgYJUU5VgXigBelU372tIw+LYlrTtsHC5riqKdo
6TOaxFeSFLr0z9BkxmvchDv1Slr6ruy+MsCsiqZEtMU5CfymIK8uHF2CNVOeiuGz1FAuCdEUPhGa
yROriEMqqVRjU8ElpQ50iOL0P0+gcuCeAp+IrF7pHlPfF4mldJT4vc0A0UIgvLeLdmsjfFtQLXoI
0WBqCviD4K+Emv+7PZcHywqAvu27H/qz27U+SrCQd0cQSaV23Nizc2AgTbstgCKa5r1J+vaFjXLt
mgkixKdoUzv/9zr1HH/Nhq4dJbJ/R11/3RC+sa9EhZuto+rTsLjMW7SlvKIQp9ImGWXrCyE3meDJ
T2MIAsCpC826MNk7lhdirh2UxtIPlekkAecQWqA8p6SBTntHrP2cu5mBSAiBKDj6zWC8eTPHuVxO
cxfGrTKjsoj9zi+AeF/FmON1d4LHVai/by1yMAOhtlN5LBLC3hEkzmdqUSsI9DWPcuHDhcQM/Vng
cDTrIIOBhwsRKEf+vU0l0j1iuiREt9PguwhVWf534C4ymtkYqcGLRCTSZbGN1mJ5dWgNyF4x12uC
Y8xyMKuSZvwy+1r0bqMLWzeAtsOpderllExyWSAMWm4ZhWSgrEDkXbXsHN+r713qDfQS5BokOERV
xlcTPrkJYMmZwqKJPDjoNBT4Fx1lfqK0r+UmBlJJfphMu65kRPYsxPpfBMpfayin4th56c/Ko+9a
6lDPQiliN8T2g/B+sxWbHyebL20j0uHYr8H9wzU+BqqgHiKi6tpJkpXKBITA31d8RIZSLagcHxdf
/pA3dv0Jhts3zxaDXc82pTD4ILbU/9ESdncfVzEbLsKtRb2dBl912V8zYY9XYkG+DlD2ecGyh0Yr
kKFWAEeX+Es+TUO6KVrJP/zDEYGiO9mLvxiHMHnULv4vB2YmByMZbbL+Ojw+WIwwzb5C+ZXYct9c
3H7hIYrpuSmQUNpRK5fn2dkW2Cj56RyfSeTtzcWYyxXcnxcFGXwwyIgTIY6gI6W84K//2VNqVVLU
HyujfTLXIk9j6fu21LzEv0+Eozwokbra/OLo1WhpMtDeA9e/BY97ol1OoZSid97hkBLkmmBQo3Wp
qkSC3SZNQPdBEMYsd6TsgiKGP0ttnTExev4mQETDTxbVNR25+YCiU47B7muvYM3PSaiAjNnvS18+
ga9j2LFOBSFgLuIN/AoN8T4Rdc9i15se46cT/p2GKxx4Nv/XLrYDtooDNiKToIjmE01GK7pj2Q3W
J/Zj27khHUy4aVGv2XdIZ7FXPGpNjAXMJ5gaB67YTr8g/DqDrhGo2EltZzHVuB5B1yNaUuWbL6w6
ewc2hVVoOf3PtTtJvrVMyfWUckQ4BQ1PvU+i5G4H219aF9+/rCMsjfWghfuhMDkiR/Mkvkx/ZzHs
kDbzqKmFROFubq+RzhdI9gMq0Lk5/ieASZKRS/E8TwwdGcVEClZXLVFoqSwACsFg/Ld+Kaa5auuN
D9Qw/Vc0iqG6JSS8RDRZLZ+m+00AeavVIUc7fmm/b2ei1Y6IMCEuPsHwbNLJfXc3aTmuYVhN05GQ
lmnhfvmuY9MOZpAiquRO/LoQNwTkqS0wqdUn5C2qw7l2NxCYPhsvuZvRMYUArQor9IapLZlVEKEn
JVKbqVnhGF5n0Ox5bySVc0l+PvTTwFES21tL2CZtaRoaXWCpdQNKaQeFX6UbnTZQ3Fwdv6hH/wg9
qs1X7b/hXAvaV7NG3T5HNK3e3cT0X0w5Wqz6/rVc5Oh38/OiX057Ev5e0WrfKa5jxO1GMLzoypNg
hUsqJsW+ZqhbpaUUmaVlBic3i5xW+mshtG6ad5VoY1gYB7Urov9r6BwCQIMTOsRcAfRsaikx446p
vy1xR3kwKoRv6g7BiOMc4p7TlHPjAx+egPj/JNmDMORFeufZQXre4kQn6tfYyrCWF//vwclkRsB6
XBg83PVoxApihDTHUw7yUIAFSI9DoqUmh7lNOrnxjGCWAzK/bpOgFHWUIfXbPR7aElv7IZy1i6Uo
JIafzng4E8ilhiMB5pSEKmcXTCNxChhhy65DV5KiJMfVIlgXNxYNkcHM5P1mi/eHlP/4UVyAw8FA
RfJgu5d7Z2n36DGgndo/8OCDhhL9Fg4Xwbkk1+TDlxAIHLz6CiFnqqqlb2UVZoJjw+ss+PZPPiJV
h7mqb0KOwZzVBJ9Ao6Nnjqgtzlt4glAfe+ZVkVv6dMmnjKJ7r65lktiaNxPh8E9Z888QXovEc4iz
p4e1e/GbQsYetwjNfvcZGfvjF1kGkxk30jfR3/7F0Sn+CV2dJv6K/0dd3fB4n17qfkUG5hx5BHza
ZZ6WaRDotUjOblR+thVhcgY6+ex+UqfYzyUA3Ka6fkpmiQpRDGyAydlmRDBacD+86Lqil5hND8Hx
Vl9wKB4qQCXu3RXIkfjAOngWQbJ4omx8fxvaXmFevYVsEqEpPp9bE4JbGffH6kRUDSUAJ+h/yUa6
UF8e1GbnaHj4KqkwL9bQaRfrt4Mv7E0fhzq9dBoFnihl6Baktrpp9FLqOmCHL9aHYvy1CvPXfYRa
IQoltm8QeUZDyN3ZOSlHdP6hCnQ6fkBQrS7xyhRJ/zGF7Gfv9bJ0z21zLGZidZM824jTmA/v96eC
Xdb+gs0Yd2K9gQoHChONrjXc79vPsJExdRmf37dWbCpbaBaCebMYilojSWl1gEp86Ro4I4PbMr28
uurm+zOASKpRhymWrLQ+rRNIrgv8TcVAHswMQISj2fpEL86ICKJItwdV4kmFcVwqN4+QC0/rZCxh
8Hnn08VRaLOnPhBRlzcW2DtQjX1tQ2XWCBKKYZtqUWJzRe8y17pgFlyiqg+XX2YyUnOnld8494Xl
Q8EE6hQ6Ox/JhN8NdUScPkM7reyshOhGCYoJyTLaTQ+BF2245wmUmkNDzhHS31Jdj0jQKeGYChxS
NK/s0yqK1QHsyHnVvaXThbOykdHVgDUzl3T2mUpHX66TcBX/ZTwcSSn4qiF7GzU0l2LvA10e490B
Wc7Bj2XMUUV+sT5yJkBa03gaGmTgCK2JfgDKyz2mApWKF0cBEHMRBEAtMXVhNmmTicIJ2cgE4YhL
jzY+kN4UfEL31LqFc6MewUmAzKyYsiaFG9NaiqCqNH7eOU3ODGKTpC+88EER0ed05NON+mjDOOna
jyOQnafQ5m0sSv8KGlBSejrMMb9joWK5PgxexfUeaVK9NEl9MAJ+c3DHQ5//VtcQKGsHkwr8NAGB
VVeBl5myFze3+HnZDvMvTIQCdpZcf/CWABQauPD7Fn81xpRBs43Ne2Z5yEE5uHWGaikyEcnMEUYk
Z68PNsfR9XN8epNxIxUOU+vRr+GEo9gicTq0U6qRb5vYh6xJwAEs30/6J74jsJof02hKkO8XpZoS
4+jmLdXyEG9N2Sr3IdvhLaksh/YZkDv4Pgkh4rAuBigZ7qrdTOpAc2zqHqZa/H3G6O8lETGQJH3+
TdXid6EAoB6cEAnrtFLCxHKICGsu8JqvbWFsRCX3uxnJC3Wjmyi2ikSy3zCKctXUaMlMUGSVf6jg
gUP756dI7QGvhQb326+glgfxUGvEJz7T6z78Jx9YiKnSxNSmkIPZxulhqcYW3wusiM/rZ1KvBiIU
bTg84GWL3SaJkKG374cF7onCG/YkyLSbRecb3QIL+9r7OM8VnTXZwKKzWKm/Y3TuQmtqNWZ99KdP
0nAKo4Rd3OK3I5mJmsmYzMN9fkg5511QCD07FerHlqLYBZIJBPI6Dt102lFaGLIw2LhQfZkCE3b/
mEZqVzjryPLhh06PjS6mbk30mOJIHe/JXHEfWM10IeoWvtPaQPhCJYstpm/EqO88pTY7gxUq6vRe
aGrFDP9xwcQj3tajUrOxz1JbWADxXlbF0iGjRBzccnTyAHSyDLsKjS+hU8vLcVJKbhvUxdfakbtJ
iS0QK09odphNV9j3Az3Hv8Zl7U5iWLkndmBpM7CwMhX1P1eyqRD3hZXtNxwVmq4Y7dSUduqcPXuu
RhuRJXT2S0/zlzBdnsoVM6ImM3Vd6E5otCTBITgLGYU6XoJlnMT4IL5HTi+JsykImOAsI8kjfJ+o
hy00IXSpQ5DD7UuVdmpVN3zslu49Wg95UNoAwaUTQNlwciJqOu093ZYCJ1Gr5sp13y2EyXo2U9us
WKMOmWlwl7WkYTlkYPrlcOjUs941XPen0CigDlYQ0Oaba1ETtXTxYsffGPCMYn18T4Bv5b8xNfJy
4IkafQy7DsSXfhbGtk5XAIJ+PkMvwqG+sheZhvEHukoPeSzNupovRM+0Zse76/EFSHZaFYAwTG+L
afys6nRBkFAb6qhgbUniF3/1yl2dTYbpHp8GyE15xxW6q4wN19bjFvj1di/RXbxaRQGUOFhsM4MG
Z3Liqs8SOA3cV3FY0q+5duzL88rJUFcBdwG1O8IvcZ0sV+w+ju5P4/PvYEEx4qi9w7jRrzyWVY+K
1LHSnQE3A/e6ChDgAL/wBuPvuqWvykkc89XhSwdtyaM3h+UYbOc6ujLeey//tu3E1/sKN+5LbdvA
9tobgbq+xeT/JlW5Zxj/HU2mFnit7NY300VkwQ3bXwrOjjRoogUKiOd7AjWdxAQ1Hsvc2xUWmmBq
ggDHerAMIw/OlIBOJjkhyD4DoYm45J7sHKoihD4VeeNeH3UbjmqM0JWXgtI54UG50sVGsM3U8yGn
6xLnu/OWZM/kB+Suj7SHxBZV4I1LYZB0LLNtFblmczQAVuYNcQtN1E8hEx2EqxwECgbSdj+fRXP0
T1DltVlXEjODT2ER6CoU3hHzhp1un8dQCObegP6EjhGoIh55QGl0HQLe1bNXs95NDgTECJRpUHep
CbUJLoXpCAef+yQC2BnWkS6iD/BMqRZ5O/6+IhJ7a+nAzWXnO9i8WhtaqbGUyM2N/hcdf6sPNGdc
v76R62WnfRXdnZxKb06j4+nfLJ1ywi6+tMR0ws24WxNzEOsc1JfBMzFni7Vai+kwDNJgGRQfk9Fb
yXZoUleQTsDAb10+KuOsLPn/DwRZ8mTj9Hz8qGW4esBOw8y1YoIPEHJkRQjilsjqffg6yUxUgiox
L505NZTUBBuHkQv0OTEXXL8brI5X+vIQfz4iYWLQhlJ7IzOyPiiuEpdU5mJ8h5vsMElrpM2G4fW0
ADdRpyBaYsHUNHWYZODJUk8sbO1E3pKpGSreWDCstnX/ZhzV0MKC2AzRaw8Hr1cTQvk6HS8jx4iI
4MtzaakJx7q2NfGM51a8WdbxMdZKNDs7EfAKs+jOiiy5iEqyPsN29NkbSbivWfhFU4cHv665bFaa
fkXKVwmdjCOHusONxWi7TZzCzAX+iaTBIgTelHj1HgnF3ZR+nglqZABawzZKuv+uBNM9NldV/CIo
p1W6oUQYiGWEhmhflbCYsLLXiM3wH7poEq3G6laCrkhHZXSsfi+LbsNMRCxpYAVVGL5Gep1AXS0q
p8uj3C4myNq5tG5BQXdmvQ5/2M1LmSqSqheOm5E9xe5dl9onoJhLCbb1gUJpWIla62F1WFo/ZsB6
y3P94zEMoWK58Ru6KDAkKnCnejPpdbsJce2DmuZQ9rjDUp1Ji1Okh/F46Y/bXts2Xvd5h6uJ0eka
NvWI1Nn3fuhWNerjuPGhGCuaj/kgiBkehUtBZwmy+XYg8Hrn1Ud8Dr1mdIsIk3McFTtVk+5WoRaA
gYywc1YPKuSneO7Dyn6oNnpa4Rei0KE+P+zWQjBqIQYc7vLIE2qeKIzot780TAWUymEzHY4Lotgr
Ut8IiAEpg3ViPLEZd9OfJtghWgpsW3Y1Ns47vmzrgtR6o4iPKmgWMec0/IfIf3F+SwGH5KjYs274
7/rIZ3ThiRW9XSQ0n0D3oVk3ONC00f8kwyvu8h9yhBJ0s75SqfJ6R5rtjtS1sLIyIOHw1tCx7+rH
oVqFE+Qar5UDD9Ktl3oAGUpc52xsV8N+cJ6MKJhc+gfcsdf9C9yMTcYPY8itK3qAHTT28z5Q6tdF
uDhao4N7c41judfRl3dD89v/Zcvrl0883gfOXTR7XYJT2Chvf1V2bQUvTSqlfkl2dwXU61eLaoP/
7E7X4uAB4H5fCdDpsZQKx2GNzjcTmKgR7qX60f53mKBrV/kYfHaECpXB+xXksBevFBII/n+q4Zfa
ei+PfCCvpWP82cU2ipE7yc8T76pVdRs5UnRSIWVjFasxkDs990MgWKoVWYICsfn6kdbmfG/n0q6a
Blb1ZPB4IRORLBg4AD9ueYZj89a3IbhHnxruDYtmFkKzeYaTKbsLZevHrjXg9J97co3R/mSLRIkF
I/iBQ5wrLJvSSTpFY53wnOQ+gwBBoDhN3lTBOSujVb10ZH6n+B5yMwsiMQWT24mDa1lZcxKn/5hq
fH1CBb0yqkTS4w5D/FrmBtIaeJln1H9z9xwQaIjd/f5g6oFLxuef5wiAkrcxexwmnE/Ren3kQdJi
YPASXHHL4Dj1Wy+4XogfPLpajnBlt6YNypdpeR7bJAWa/51pqQKZKa70HtSMKEs6tkPUyaZqAuW3
ImnBCCVhCXYEwQME3ebIXWaq4yZv5wg4z19U4qlv09gBsqwu3Hyx7zWzr4tIlMAErIYIvEGaqluU
R01JLrMl7SylIuddln8t6EwaGZyavANUIcFl1s7mUTgMYDCYBtj0uI62HEW+TVJcC64g3CKF/Ycm
Le/NOfSnb7+/jwvWtV8KUG9KhrZMg6YZuK805aBydPEcIoX3+JLsCbV9tMcS4C87Sh9trSWU51iI
YcZE4PD3jXiE5hRfzRkvubYXiw/P1L+nZG86m/zegtQ1BeO6B9G31iidM2PeRBOkuq/4kg9+FTjJ
KSU6mTdBvMZse6Paa1drwsGdHo6p2QKP5QYTCs7YpBABCkf7pkxGLtlZszwXhfWEiDGDNZ1OLDMu
vGXzcsPtFfBNouxVkxGqiFTvZUlm1PTbhgcZ00VTsSAi9aGlSh2r6R8Fq3W99rEyYjk/x0Fd0bA0
5Nua0aXiIgOPXr8HZhzLcoi30ZF9XzNySeMMGAcaM0zS7n6K5Rs3FEqglM4ok4tTIoDyytFvwVVp
2GvIRIfa1h4zE0E2XVzt3x0XjeTcpUM01XyiGDmErnpbSd9VoX9m+TBtH8Fkb/vzBkaLIHaIPPMi
Uq4fVU0qxIFxaDUbYKpphACTKo2hwdvDWlFGIlQFG8NxRFejgBMmhS0JA1XRH1YqTUZyOpTj7xAK
YgCmdFY1Ub/TvdJfi+A+rz0rL54fi7a3pk2xTJ7gnmiM1l7Fz6wjFjdwNjEvf2OvPEPGtN2RAFiN
r9QgC96H4Y4S/+enDnAaHj/O0luShkQ4Lkfbx20QMZ42K4RuZE3o6G6+6bCk6gIOTXLboLSYojHo
GjUUT9WgwENgekepr3ZqFid8MnXMzZT13dbEuU/YCDXk9ajHDU3DvoaEw3ap3doj5Z1Bi+FAIUl5
NPqA5cII9CiJUFRf0AnELftSJczLWUtbL7yg3o8XXItoIVcdsVgZ1FNuv924zyvSXSp+wwqLbEwn
Gv18PC+44t10zOQt5woK/nogkDSmCpu0sDyJV8jtnOPF+WzP5ySIFldHyEf72C2C5Xo5s69qZPh+
nDiMYPhmf9zTgNWXrlG8ikc3btaVfL40DNaP/ULA7H8xPergjOQNJiOB1FC0jQ57eH3UQgJQk1Vx
bZzrGdnEcctawXnHXd7vm8BwPHF9jonO62lqhBO/a1xcGMt/1+QBSqARWWaaVMRJxoLryfUvgwFj
JQAVUua7mizqFe3aBML53+m953sjbaGef6zwWXzejOGChiDpcqHN48NHGHZpPuDwYxA1kM6FeVgc
yaSIoUYeAUuMzcvbmUbN7AGQ2AF5d3x8pZkS24Rzy58+JPeXDel3IzQr5M4R6x5gI9brqveOvdOJ
POntRih8QEqZqEN2f7N+DD8DrKmVonZWNCONrV9Y1g+KMD+kXO2qUYuiuDcmgQasGb+5v53XeXzZ
llH2VPe0aRHdyQF55PBqxvpbj8UxVoQ1+jv5jbZ92yIEi7FTY7PbwWcy4RgWzekPaB9YTvJ54R0T
dg2+Vcy/H33jDnKMifjltwGnQNQtlrrqNLVQlgmdtaFFDUGin3nllbT+9UhlTRtx8X0euAI1WF4u
g2SmvgbPN7qe/N81E/pDgV26U5fswqqLhyVcVT+jjseYn0OTGOyq7WNtnVDCE7h0NTtcUjPYSklL
93mUFU8JQfvHea1Qs6y9orUEj9o+eiT12vYmotGh2CHZXMq+mwS/PIFYoZQOfFiBqNywTJ51QmI1
WX6MfvjY7VnNJHvoAyqVbwRejz6KllvTH8RvGjMBzL1rbT60WAoKgT0rdLSMyCmEfmaZ8PcFGOVg
UXpT40tQwBvEGqOfRoxTGxiVe78zjqG0ALjSPA85XnDoFfA4uw6qxhOFIJZzdP7z/583Y2fDaLHz
0RqW/Gy3RbYtWaIkIrN5Zu4kj4SHfRvYtCjxAZ5jhzw6YeeUgBd2hmaE4gxbdlwFejXk5caHabQg
X346JkgAdWl+xLOZQyHV56HYsUYa6hsxumxdFw35OwphbfpvtpcZ9fujXvMlP4tGzwaHT2EFaL3l
c2aFdiXPg1iIsf+7QOIVUhhF99Cy1erHF2LoxbaEzO76tifIKwNoQzKxeRpdeMJF5eUYleyyX0QT
DxmOeEJesD5e4lhUmaxzcRpnWVeQlXy6VkrAP/tzpNfEJDH+uTwhHRklkN+bOU3Ir7HEQgmHYQKN
Z0aV5fkWjW9KNkeqx4Z82gFQSieTkv5itN7IGaJvKVjO+0ZOCq/rpnYHhpC3WoidXEHe56xi17D0
NnwXCBe1xHeydFtIyX2PYgBGQR1POw4BG2eXzpYELfJ3FuVGFvvHGcUY+jAJf6UT9Xpuqs/ssw9B
n8+JtBjl0MD0NzoxQasfh5qu/+NTUMp0W28vXDZAvbbjIws8mkikBsoLhPf1mdWbwP8qWEKG3HYM
Roke45n4pi6HbHsz2cQ2lkwzReSvqnIDYuXsKqkfuYOFv5EscSDj4ebhkuKWE5lTK9lLQNPMBd4x
7zVo3SW+zrhSY/5G7qWAerLtxMDw1tC4y2RUPU3QBNF6bNZr7FZwGe6bwwwrj75wIRE1KzHAySR1
0P1GWMO0nRQa5JOEteElS3PUZtQNwBx3t9UU1JL9439KEWeX9E3i29rSGuIToa6Na2ek7buQpSdT
i2Q7uVOvNvTY04SZMRVfep6/R9J5YmrkgEBB0wVUo9d0EsW5JzLMZUdlCiPHdIpoj36Ak+U6ZopP
MjVX+8gz8gtZIOKZyyw5ZfgVLhOXsC4IaJEn6uGk3Yl40T2K9hTyS0FNEcocLjXXsZKj8LIOphR8
b6OliGENMh08O3Y4FT5DSwSAZ21gDBzXlxRpP3VuaNhtP1melGnnG6dYRGHkm8rynqnlfO0izfra
ao3ISpzl/q3+Hq9gL+qtzgMX8QhZczfI2XKHSdSzbwHb5BgPOCIHMw2V8+JVS3ox4hTMmuptq8iC
LLGaGSokJgjhLRbTgMAqaO8dVPqFs94h98363CXcl3of0lk9uFCAO7C791t6PAAkRgJ9YFIipHO7
wdfX0ULU2gLaEhveLOqdgnyS0D1coPQGiD4pcY08RjZbn2O9k7voLOncg17OkDCsZd11TQJJV5UD
1UZ3sOv0f12G9+Cv4YRiY8ypAv6b2WiZ59q6wP6kKLu31FDRmzbYmImlfWxZo1/A1y2eFwuzwUfr
bR1o8JgD39J6p3Xsd0GTZ6FBM2mY/w2t5JY/iJOIcaWs4oXT8isezmjf20WvR0WE6yOnU4N+zKxp
JgJp2Of0J6WdXfXi3/CldO7sibuu0yH69LM+Izs5JXJK3025aTgjAeZAvvV41vKYCsHnsNE261oG
WcRzVRBwrDvzY1fqv8Pfw6jJvmpK1KWuvPF77Wj3jt4ezegQ1IoqfUBnlq+g0L3MuVmOZlCPnYaT
LaHpWNZLmQ8EL5tWiDqtNt6rdzFNgn8sJDQbcMONdtBkdaMxWFQEEBZTUjhmh1WZiDXpXwdLqdoQ
3NENlvorQJAdd3hsqvj7VNTlgOPQfEgmsEi+9kEcWI00NJIOC4+ymXt2NaXeynIZit6Z4VqEInMg
xFUUIe8U+nXlO+dlq8aQhSpW4gu6jDZ1s10fK4UsuBNE3YycZJTTpMYzdV8X/gm7doVsSPcsbpXm
+T7KjN0F0au2e0L3hWLo0ULiKh3b+B27yBjmefT73puytLPQMYjYutvUd9nxkb48Aa1SYjWj5lPV
NR1AEjFzlIsICuzwWbiR2JsHqDp4IFHwoVT946KutwIZCTqZGPzfXEZZOpdPE7NtC4CSwhumSblr
z91rH0Xd8mCx6RKPoOFAeH4yEX/HGziy+PhIoZdHavwJT1QWSwTlRGehOGebxk/WU8AgCS/CieEe
z28NokjlFAlh5zZ4K6mVVuPWfVJUm2L2qDXa+ZLtN3whrCHv04jLlSSHF4yMtl3s4WNJD5Vux4Yw
bcUrIe8IApoLpX0bJzwQ1Q+KcF61GH9cfJ9nUhZ4dNkVbDO6IukIgQbq7Q6MuSQNwUKeLBIp81AW
ChAEW0/9ZS3KpdCvx+rD3LpjYhxDvYiBjpvqcrIsMjqQMhEDzaKOt+HuXCy82g16dJFBaKVTl29w
neJbnWY5pLwEhzLjRcY3WFA7asLf9EYUWL5/akgKhmhCLCmm8JhspLD6rj4SvyLcaxzHK38KSl9X
SFZ8x2qclfRR0bY6B6exyah7/r0rR4jK1o9rI5Jw/VqHpL3W4zFSiX5B9yZS8yHd9YF2obabvrLC
/zPAcmz/9hhS9vFj1suwR7pAhKkmQ7wuOTJm4DZpwMSFIz8Ym4zzqnxhKtV99R/XZgyxNGNy0H+B
mL+1+yo43NoJqq6kyx0ILx3rpTCSW5ajHR2iEuxLSXqavllKonlxAXU+cdkKIUs7q5N9R3/x3nLp
MgmEL2+VVnzQz6FR3lBDlpRGb618ozs/RtMjMTuPsLu919OwaWYBCeY2N5KiYzD0PdOKYlmdnO/f
0m3DrwaOuC3IQXETYIlSiy+Fk0L+LOVcDv+MxP/rSRDSudtkhfdKM8hHbQCghXpe2DpvuAHS6ngp
SK9QlV5/AG20HYpQ1SxOWJttVTFXe4nXdGcx481+Z7LfNrFO63nf70+Kvy72eqxv5uWLx8Y+Lnmh
6QABGhho0zStvG1f83fg/AOSdeNHQeMvLq/ZuI0VVHE+QXTlA4Syqiy0P7fsg57F4d4QYoYvRNMl
2dJmy2KjO14K7MxTkYwzuxif05Trn6D5PtrFsKw/AE4t8XR4L5iojSD/tymXAEsniJFNXEIrUL3H
NBkewQYc7Xd1gC+dGfcWpLQmXMqKtmcrCnG8pTlz3IKci+upF9ToR/BtiaRaB8c2gmFrU4K77+/2
iSgOofKhT6dGMVzTICK67UpFnNOhxHZ1uyd2wNThW64BCnEiUIGlpHOyCXkf/9ustRKqYItJ5Xen
WpBRgpmEUuyH/3D3758Che8YOMS4FjQMBr4LfNnbVxZ8quWa4ZuvAMPusEWiX2m3MNGtZieeNx4k
VU8lSCwZlDRWYkzAPhJ+Nsrnyvw1i84lubBBXjY5zjDNvchPQEOI+faBXYoncfSIsh1q2rp+F3Sp
/moGFicqnELBK+COGHkgvohPCdTNTY/912dkj6/FmEzL4bKbJamUDfLhQ0vjhWL20H7M4QU+0xtF
S/IFlhH97wrXnJzgXcMIvLSuJPfSeJe1J9O8G3LlbgJEjDr1P9sf5Chj/anJCqJDJe32O3lfCUHe
1gsze5fWV2LDA/Drw7lMzUuU8UoMuMfdd2Rkf7P23qyvFDtAnRv4McK2g17k86Xh/D53RP30xTUD
uHfLT0aB+ayV9ig4VsNcE9rdy4D5LaKgwFKtuKeF5baqrNVUKnwCv/+po5alRzxvDrI3H/nOM3Y6
5oSM67KAwyfYBJXNp7HU3WyDYYCRw9Pz7vcmBu87F7DVnxJQe3ZymoXPZ6esqsWpk0dE0MQWQn5h
DMpY2jdeZznofBUxj3SrR8KuZivIubzY86Rmsl761z/AWgcBEKA+GwZJCa5LXG1JNdR31NpzsOfl
n6kCEGVX/W0mzXDyOdkbxFy/NrsRVa8kSnlsjvFKQEMcXxv/ERO7toH9WcVvzV3s1AU/0hVt1oap
TT00lVRSuk8t3LVpwAf9CO6N8/5yehOg6exqyyM+9X1nXo1io6E1YV0lmNAU/8FU071tvwVC1IRh
xuQthwJQlxzqu8gbWWVua4mDxQdmU8BwRViG71qBXXtl0oIvWDBeyg8GtpRBeh6ge16z7SGEt3+M
hf3Fk0Pm3BUYguomWYJxSN9SwzQB4g8DzZ2UuQ0nFB18AMLN2JxVFH+ip0BT3oFh9HfXc5EXw5xj
hAoN9lreURZseLX0assJGX+dzkO71gmJeLHEnEhY6MFSordst2zlYc0L+9pS6buOvMwmLHxOI4qr
33cfMNWOfNCb5hG6m7o7+oY8v7r8diFJoDHAdEVe82TWH3KBtIIJnAzA4/Lp+poAQSMcQRw/+tnA
pRLR7PLHz90Dxwr9tmj3WvWjC2CYndTdtdNnGSYNTBmImGn2BdhVOlSKuZW58UiK24fUrm6JQ5Ja
HVRCRwE8RyeOoLZipSWluZntzLgxlHaTpDpjG9RNuCe1n9EMH+NI/dNcLfCDK7KOsScs6zQr/Smk
4tvXzAxcLZKvbV7dXQpUq8Fu/QBrymBf3XIuhgCDpleSpmrZV7lQmf0r1qaSzrPXP/VNEr72oGj9
QDcN/Mt6rxjwvn3F/MY19vDZGuoEKZ3DvCVoHpu5/fDYbFRKm8wqTv5IEXl2tAK6jg0C9AC+Opz0
yyCnmHgnmCxVaYnYEbOzIeG5r55p78GIceZeC37jjR1xAm4JP/g+S/mR0EcNnknyC0MpWKZjdTnB
AsQkRoNS1n/3fF8EaWJtlpKlRc1bOHOmIbudgyU9op55PM7jD1Ki5zslzFt35rj9C9yIKYzL4bhD
B8S84NQUPK5SuSguuNuvh2xP8QVwfsefDG6d66L6vsDVUE8ho+y0eAsqtqDcUD2/H1Pq/1cxjvJa
+MmOL4HfVYHT9RqQGvvzqYr545j/Hq6cLvYqOy7sypQO7Wc+pAIpLdb5sB4x5RQNgxtPxHqxqKpA
SQm7Lly8OR8WH63QadMOEJkwb/EHxAigT20vAIyBxqArNNyMXm/TSetQrOMwPIGvVFVZYq7j7Jnj
7gSIN1BVEA36F5YcZ9UPJ76CN7Z6nGB6jxzzz6kSTZNRpOls4qOIoyoUmY+7tzp96LnesJDGhiy/
vSl7gC/jJ55E4qg4G2TZzVKJeVwuzIAqiLgrfqYkXQblwfeVvOhgXhy9vkV+Y2vgJNr0jtY+/Ot5
UZ7l63biqHNFYnq/Vaz6WMVrM/T0yWbwbIVga8i/65H5Gcdpfs5pDkOVu0NQItJABIBxYLhxtR8O
H/7rddvtoVRSeNa5BpyhlB9OvGVFWsL0Rv2XLhQuJMGxYWjLdrqBZ9/caagRJ357ogdeoqEXD8gK
rkYbuRRCea3lRXX3TT0eqCGp2EUDuwkLEYh3cdZSBuHeKYwAkd6G8Lqpl+yrbeX8Rxn9PdanzwpX
lCS3g7r8OPAacd/FLKb3v1lI3C5y2InADXvetoBkYutNC9ZK/4I65Uh2XBCDugOOgvGEFary6Pyu
QtsMo2nUQLtIDfSMTDF+7DEOlGjALaW4VKbpgx1lnGr61eNhpOe4UmHiR7c/IkeiO2nEStQtSrKW
kMsRPgPAtxTQlMH9sXhJ4xOj+ymfirlHf1cljzCPvQcpVGsg0dtkpyjqRYmPP8M/2ceC13yvqpRS
iLs8iNADD0hLLvELZVPTnnQXoOay4U3XMnBanINg39VJIl9NrGxd6cLhHNdXxZ/dvyox2wXl9ckr
zcSuySQrPO2QqxEWyQqrWrnsiEB07WkbYBkPtugyYaL6wMzo24nLTtN1T2UgFQjOeRj7xSCwpRcV
wMity4dhOlk2Fbi75VQTXrE6R0ZVp8XqBjt87SfUjeIVo8kXSSL2CKaMSvEdTc3lwjZctNt8pv3+
xeK0Iu2FtsgadRAl0KkV09E8zWV+k6Ng4WkCT2j9iyMJ3Ww1OzzLDxF8YVsFnIM/RWkBksYVyg9s
kIJeXsyqqxEA5EcpZmStRaEhHVMl+L+S2lwru7pCUy9zN9DTq0OBgs2rbSK6rfQx9/brpOPXVb8+
SXd/1QXkVJQnPxp9NXwmYmAaokurCVkliWNsmVwJoT/1WLUVHAGLq3yxGIe5Ruf9Wb+SCOTQIL3r
tkO7b+b79HrD40327VgUSvY7r/k7TWbRmkKxuWudbYylYiXye40BLSqH7xarKnIyZro46KKaHAbj
1lTVJq167sDgblpKtBuuCB3kPFnYtbEB/K65oeZYSY92h6udVl2LQ3czRtmwHCq41Fk9OGt2FRJG
Na9FE9jAz2KvfJZuRBY6Y5sJ/+mrce23FMd4/EZ00abHPt5zsE0XZeReyi3LPh4QjbWNf8seMcrO
1jr/66ospadYTxCt4Kb5XQ76WakDh7NxYsyOxevEGrxBalaJPBJZ5S+Aflde3DuIlSvYJ27UUoWd
Ec1sYQq+l/AXpzdiEV+HBrQi3QvQGoQAGkIdnfCORCSuAlepgM+J2D4hODNSESJ9cPf8tYNrWvGK
e7hSSOkOJ152pSJOZltetOGOR42Ocih4IBfkb2kwcenI5fkAGdXJ7ZCO5TU/mA7tN0jND04S0xew
jTYs2JXfV+EGdGpNO85AOYuc/0vxBOFeOLBpoMgcCmtk7ilqu8lFOVtUNX1eIIbacFzdOLPcj+En
0FZhA4hiyNXi3zFuuVyQx/67XdZA08GGA2DUrAzfK73FWQSjNad+5eehEsycKZ7STW283zQmOate
2Vas/l+gPsS5KR4tP1DuP5ltT7Dp92dKDv0KCGZXAIGQKpPcjvWW8fPEahszPQc2Elnb7lRdrBKB
OapqCIwK/ONAkSULzXD5BCmHRMueDeIWEq/3k2VqK3dIUqA1YkuuWVK8NZFw/9BM9OXTNmQcgrZJ
uFwRG7x4ScWF4j2OH2YatKgXpBNxawvuJJfGsiWGlhjwv4nnhM9sdky/uySwtgwsRfOC9rmCYivA
iO7O4IYJAKv7SivvIaLHUINZfv4Epswf9Utj5TLyYAHi7gTzpgoWnAl95IGYkkZigcAYxhhI441M
LKUplhtbtby/ia0Vqvavxdw8bAorh1BVzBYfJNCwa7/OOc15ICWqWOR3IBdHBfDcLs5TQwLrdvgm
Y6sPvAhI5Falqm8lo+0iIa5lmuUHDtfmGWlCSB/F2jB5cC8I8jdS85KKp7oJvoC5j0fvsTDK9Ohh
c1i95Nj10ai1mP19rKP/o96tRI258jNSVPvlnRsC+yqumi8mVzF77mjTx6SEFucc6YXHo5hl6Cvi
5aOPBXcQJUm5ceIsHf4K7O0bdMCpyqBC8F2TI2MOkpNgDjifWuMdCJHWuXkrBW+NrfbdI70Uzdkl
1DsybHY4cpo/0ggUbeAgz/dDJx0aV2o/YM1kSu8g9MiIn76NfWarKq9+HBCn1IXOur83Wrs8Z8aC
GL8H7U0tKcalo9QjLPdkR0EDD3nipk4OKv4992y3CUFq2E71fFla2zEUVlJMu3b9dBwTM7nqh4B4
AvWKuaoVwDbldiDRkvHorSZjtDwCTUrU8ZWYDALnGHjZOhBFkSjCmQ5R/9K+g6rHyc0apsNyPIfj
DxcwxkmkPgLzzYTw6DWzrL/aS4WYT0rhro+uwIFnFftMMxXVeNSFggaZ4gS6ipzOcQYC7hNbnrJf
0X8R15pecQczCsArOGB1UHou59I0ASyjiYfyLGVbexkpsmWxwb7ViCCpezlGTVL6m/9dQUfpbMLW
A3jN2MOLHY+AbjeoM1JfSVJF4ngsRECvcj2X+xpJfT5a50XUEKffZYzDGLH2VM6AysxjGY+rUFCR
bZ5Gt5oaxU6XiwGfvJJ7k9BNDLuiOfxAWrc85F21/DZHBsRheFlFk8mIQqey8jURt95h8/q4JPaR
pJC7rPpnqZbJDoCIPowZ+DSR8HTL+211A1+DBGfhM9ZbmuuSvLPsSI33nG55W7N1n4dULs8vUAVS
t4YSGotFk5jHXXkP+E1THa6rFpLd2ug7D8suNMRBlRy9skRvX4LyqhCYTpUPO4E4+xFy5nys5icU
npeNhxbNXHX9C8QAy6rSZzlPPV9BuzBr2q2HgW0YN6aSiwbhnHZPXCxN+umC8YfsXCvS6hxF60TB
Z9DzE+PDGKiqnBOiEy0TwUniMIi91mIkbZK0/qKhFv1oXxmh01BuppoN6xpLlIHo1esMjOWt7KD9
hN3WMZhToOIfN9A+Z/bzqpZBm5mwZDww1DrTTEZEijg0AsMVTKiczzSxyTrxDeDVZeRLeFy8Ynxc
F/OQFNLxTmsFTxuChRm8ZGkoigZa8v9hkVjKW1J79La6C7jAdCyOfuIynv5BGb+L7XuHM7ePItA/
7ZMYO1IEgupKRvuM8xpElm9oAZv6y17rGDIp6AV49tlyOMGIpbegUU9Wf5Q7m9KW0zvCbtg0zLby
3Oi9jQSO7u27EHk+AGd1dXq9WRKFe+YPDB8b+7t4M5a4TRDNafTNnoJEZEZ7sbQDJQz3fJVn1Xqt
tS+qW1E+PEltA5hVavvORiiJBPmyZF1u+E0elqI+zNQpue/KA4o5XurfpRHwmZARU3Ef4MdpCG4c
O8zSZ1cr8me6MRJXV1jqi2nvocP4p9vlNhFgN10iwH9c7ifHFN+nCI1pwtrMtMAHm2KfuNs/IHow
Zb3KFm7OKe0EqKDX5kbIokxk95UFBWzY+SknEdT92/HM1BOnVsSge8kEk+vQh05zAT970dCKim21
Ju7jw2xnMU/ctWtGHbJ/v3OU6GDgv//qz/EfmsenZ0ja21/Wg8jgz2nkFA/+6m1Fcjg1GUytOwgX
tqBKbKEI8oalZVzVlWG+cbluRRsZfs6giWwzrWcPCB2+LUBTqbAGJfKh90e+6lgn6l43rctfEeHr
miEFlCozTjFy7CdPLByyeqnvtCwNRrtRI9j933B9FXvdT34OuyWkW+crgngRmY4RdgC/jaqxb6nF
VLe13LeMijR+fgVGEjUEonYEQ1tlPY0qzEfKvXw9Qj1qRuQC9FsWZTb9+tEte2ZxXmen0PzyIl1T
oCW0YjYrHou4nu/qwK2bYN+gzDCpMkBoUK4dZE+ARNLfvEKcOlQDQXZkAv8CKT6VPfFwUNyDpVVk
my5loziYRGnkVQGgKIdPVUzjO1Y1yvmr0XMWIqqWkQOLaRptaeFH6m6/WU0eMf2EinptArTMKRvk
NQZkci983nB+yQnzi/O8ZrF9+uVCxaLdjCKcuBfkg4UIeQLuvm0LM2a3WbYRoObIFeAy7qewPKwN
ysSjKyQ9T69eCMdXe2HVW50Dpa4O3/3dKg7vlTrbNG6wM7RLOMP8d1y8bHWVfdlb3SkQbV3SSq1J
aiQi8Nlya8LSnP8rj4SNd3e+EGEukP737psqiRaXyx/3xELVCocuedA756SwUPNe/naHmE5Qe3i4
Nq+2Gr1LhJ972AWij5pBklc5rzVgPHxB8+S7adVvZyWZfQK5x1nSAnz3rxbJ5Cw9TMWO/UU6Wn/Q
qSZXGyn4r1BRQvdUptZndmg4ELV2IwG+OZs9gZNdE8jvxpujtREBtPpxHJyzqyqNjXeps8xPuZFe
5X7pZyA25W4VEtObs7SQvcAdcUmKI3fkexQjsLtTbbtWpZZgMw6C1UhucPAmYKHOMxlADfeBK9qK
5l+mbOgrV3s6g9U8rHl3m8CmXTPoCEwDAEwxAgzwElQJX63RmYA0Xaf7xUljlrTgszozPX8AysSL
vcEFrrCZ1CBEiTpKY3i1y8zeduSZJ4PLWdfW2X0wX2t3UL1pac1vdTbWg1kJzDy/IEGiTowaRwPi
spZIZzRXzp0WaMsjpnuCbZOoUZJueZ8tgsCHhiS99eA7ODpV9TGy6WHJEjKXIzubfw75YOD4UCJE
QnDp6zfY/1zmZslAvcwoLL1wlZYlhNpf/wznyYXyv9J9sxH7hyNsDnm6PyU8a/gRtJCDFW5DCIlP
P/BPgequRlhSKcxXdId8zFwjIraKk2GW5Fne92fStwo8XYt7S+09yxts1/krleluSQsMZNYaN8k1
9Q8btR50Oc5FyPXx/cOJIJh+mUvcjeorbTAd/0vsFVcI4XJf98EkzVAVAlI82ToIwog9A9Lfryx9
5xR87tieAuLICIhRsagAUksedlqCOM61Rj+AMeWSqDc2Ppwfu5IYjMHLzUHbbYAnxvPXBu0OPm69
HTHhmNJcH2WMT0QEwyvtUnlfcBuM7jWExLnDxzNGzpOgBPgYO21bhYmEYk0+E2FoJa+F+C/bwqnP
vrcSGIy9NkNZivlCfsD5ESQZRnmuuZxxQECkQBP3F9O/EVcqlt7sFieN68PgrT6n5iLeoorVQeLg
EP0+/mZPJdSEGdgrfD7Wy6JAkpyyC0UgNcHZkhElFCvMLEPJ69KFJ6MqtGvaHHpnhz+aYSuERxBD
gOYFb9hIYoVbBFNro+M/dSYAS7yruzuyBXlJq847i8IK5jmi/SHHDSVydGxUQqUgLA1uBiWy/W6t
aBJVmJYQyu7MkCzd3Iu/tguszipPdOcjV9Ru72GQ25a+2hmoDXP7ETHRtU7STvMUhgfkqHr6UDve
dMQGPbUDqhY0Vpkxpsfzg8ixaUuGJiMZ6QrmC4rBSObUwI+pZ23CEU2JzFeD7Ok4WXtjtEUdAfhy
4do3H8Fr1EmoD5c8/N2lK0ROOj/iaXaUas6pza7okvw6h3xAfZ95QM23aQOEc/mX/NIJvxJfVBL1
b0L5Vbdz6Ss15VGwTCsu0tyjCObxnBmdS49kTD9zjaJP2jQX+DW7elKEQl3/gCkXIMyRq55x7ozu
byDbxizOPvpLHyHdIy6Tv9qM84KGNz9yx+2pOqNDZTdHzt0dAJU8b7TeGFHmPn++LfzX1ErEjlUT
ifRiQAK2a/GxBx3BHbFpQcso4pkM6tmwhjeO895cYIZvsQdkibHLRc4mdeeGmDPoMdIJ6v7+8Ldc
Oeffwn+okDnCwSPKjD6mYUib6cEo+eDYUHcWdxBLF+hU2QA6idgao2QN6srlrk5rBekCRMm+/XeS
UO1IrMT8wVHf2f8bKqy/Q+Ia0DgsRgGpM9fGrJQekw6b+5I9pzpa/+LI9NoeCUDfSd5/b7crTzlA
vlo5xWHlmGviSXEIbUjP7BAiL3Px53q8DFv4Vw37Qa4SASlmSxHg+UZy0NRg3hchLvbM3UekZn+a
EKjG3NfxIMEG43YCh66i/qIyeRKAdoOckswt+2AtFpweZKCCO3BITKsU0o67PHW+sFcAouClDxD6
Re3ZqYO5rWi5AZFvPs+1jVRwoRF1sTAVleitCqyP+s4pc5CVOfsvrVNTm+W9BE9sNwNHR9HPOSrv
E9ycsdcWzoCoZSwTzpRo0qg9nST7Twa16dWcUhGUI0F6ardTt2Z4yuzCBVI5hnaocEz8eGetLIs0
zEEi8cZTkn5UHICzTgC36dD60hvBp5YTyzDyBYYjftX0HlxjKXYBuoHWJ5Em72lZjCt0dM2GcmNh
elcxjP/a3XbApJhkHXEvv+xuEMK13RSaB10SxcbPonyal+FKXfwLX876M+MJSdTgR9AcFhRAhe57
gd0CVFCsGHaW+nZgGYX2KgfwMkUgtcH1khUu3YUL16P+sAgf/rGwtd1U2L8NFPL46GvgSypsgDhM
zV8jykncQqHPdmOqSi9ofv77vpxzSjkBuNSKUkZrgPJmrq3aZy+ge5HxLZg33vIZb6Rtcn4wKNkA
SuEFBZoDTxkVhZ1FAAy3+mSyCqOB6ByVDE85VbE5Y3jWCh5ojlCccS/i/uXvOnuRrMXB71y6Xzj3
vrwOy/X1e0b1IwGZWLWasgAlbywKffP6QFEmfM8pMDeojYLsPmSSCQ46s9pDHnztz30PANI9oa5a
JH17JxvXLYBrRYfy/M2CHc33U9u0O8ex9nXWfso2hnObr/49HZ6MPtZ+tH66lhNVktx+Ak+HjSCo
9xy86bU0gwBdTUUQ8Ejeux3/AqASkd7M/IjlRE8MwHCINBAUdwoQfDujJDs3nb1RTRzgqZFY03A/
6Zpc8RhErnHlbcDNPZwBMCIsCCXzIT7fN3aB22ZI9ufXV3jeS+CBXhgnEkNDHYxPQIqmwE+XRw3D
HBWw5qjzmgQp3GrYH3Fb+MKCNEztI4jEkRhJzQTaHh9TyE0ReQa+T4syU+i+d2PyZjLKGfkWg0Sj
tF1GQYMv46EO4b8h6eAu/LxXMHIZXNjT3aNgB/IrTmP1i2rm3KEHSyunxTv3S9nykdp7tsk5jrqH
CxzEf3w9mWm7o7C/xJ/dACRts8VRqlL9dPpGOGHqYbInIwEQxKG/GoQmce1Dr++fMnU0Yy3ESagC
P0z9PPXZTk86ahGTgebww6A2vQkiS2oIRCKO9QeQdrhKMyCLquKnkMrwAxLiFN1wL9ot1lF9/g8/
Pd7eh6O8bLRlRE64wAjdKxJ7/L0fQOiK0SZtTr+o/KMmg72gI0Mhe5lSl6FopJ9vaBUhUAWHuiq9
yjybbxUuAyiDNh8UWRgYyO2UrB3fE1GcVw1hAHFLMpD1aoZt7NUHHC4jxnI2prUOm7P31f3XubS0
BR85CqwPUIX7pxjdnjg3zoaH5ryn6sXUkHNeLYQMMAar893/DHffyWnLYYCRLCHU8wM8N7/GPQy9
zu509IAmANiQEVRzLs18VxIUKm9Dw/YBov5K1e2bmFBMiYIIOoBB7uLSc5ZqyKp1vuC5NojG5bZx
MNQpUUKqT9xSivCJTOdjlRSpmKJShrr//4lCl6rABUKbHZ/H1IV/01fhP7LIHDRYDb3CJQ8byPT8
kL9ekDVQh0W00BHOI3pRBCnyI4gebxuLRyvNCfZ/ayDAe+YB557Uf81rcvWMKstRCLDnS/piVsRr
hGTb+bb+Nbm/PET4i9yPnS/kNd+ojAg2ZHuHTWuby4H00b4Tv4VmZUQaVbwwHz1Hn+/R/viyrOzY
9dvc9RgukmqRvys92oE+VQE4ltO0wNlA1Wgw/S3ZrgLnU1Lsyu6MscNO9g1miZ8UeqK20hlQL3IT
yWLX3+noVYovbSzm2vperrE7AOKo3Z5kFYpBVP1i3iL9lRFlidnHraGtT82P7g3iS6xkXq70fVL8
2uI8MVEINpslIAZ07ivy1Exw6xv6rodawHPnzKTciXu9cXYjhPuUQT2lkPRMR3KUXMDGeTGAfFyB
Fe5dmbFtAlB+VmkqAmTNHzzqV5Obbvhao+buuDd0uPOUyKDgosygMUNAFNSopVuNcBM08GSjqfWS
5oiFblY19uT0GXDraCUtTYzaYzprMSiF4L50kJQEUplGKpryxN2CPjCv82sfgc/NCquFnzK9DgE/
BM1RKTsLq66tTZdn6EwuMYJQyuyiAvgggw4bER3kfNrWeB0vMz9xRlXNgy6PXFZRqwJ1ba32B1zV
wEOH+XWEKksUZGyb/ymBXdkdnzL9e4GxuXjv3cGtUUwx9ftIh5UZ0+mHkYqnVMgHFaeN9a9WN5HO
jj5FjfNzh7qf+U4d0HNIg8fWz6yThWpRuDatz9XVHqHPplmavY9iYLjoOmElSCwzlvFhPGs2ha6H
7EeO6JY8B3tdOHDIHad5UDcYa63EVU2bTbe8dNxPxruU4HN2sMNv0CWPw9n2siR91NiEUzTGgvXN
LHC0LUU2Q8vjI66/P3cqfj/lyoIRp28SCpmJs3Of/NtxkKXBBlfyixx1SY0NrYmtnXcfPiz0a4k9
lAhX6/FX3u2PBjIxY2h+okAXAnLH7wI8LCVI6l3h9tSVaIGl17KnO0ID5kLWRawi8zqmlM0p3vgQ
uAjX7QqmRPuq1wRYVq8eV4FYp+A3LvGmbqDOzrTKmuYSuexYRv/j1t3/Ha/mqv3iIQjcUqTxnPXH
Wcn3U/5HrxOzHPwxOo3zJpK7hHrWqu4barof6VsPXeDfZkjYlcqSDvnZABlkGCv5vnTKioaROv5g
ocRjU/sTHVHDmd8FqQd+5XznuS78CBtdeR1wCoiRUYWCoISewu7a4ph9cnP+IYfDjfYs52Y97v3e
wanNQoYTm//ibK54WlFTqakKgDVgYtz0mDOTbi3KhAK/MlExwKpajG/jSUo+PJyNH/RiZoRWtJa9
iXhZT64JJWEL7HcGZrMKR3xD4oxacGQsDtCHf+nbAzDWfEjH/7qD6392eiz7gmS6Tk8gqXFEimHR
4HONaQ/agBSdQfRKSk2W38L3KUQSXXwY6w146LPtKEELCoMGr2NEG3xVi1gRPd5nyR5xhFyxDumF
ur4KCxwuulo2HUOZVNkyq+3K7C2Ccd16Lnp5Gl6NKpyz0QR08abrzQbvPioLmdKivG7Mnkoxmc0x
deZJEJG1dR9xtaeAGuzBo99LkJCjMeZgZvAKFLpEdrDIdk1pqC7prpYgcBKSJF3TxgYb2sfaTKfx
oyrG8gP+Hawucy5a50cUP0UsjZ/6S9MCbUVEXmcZzsbg42kOHuVC8oFybzSzv/V95x/7S83utk85
BrcjOVkQDWo+JQmoZ2l6kjo+x8+AO1c+3D1+7xIhbsMoNMypBnYKY19j/t7LblH0cMxQ46UCJBXB
dadsycBO80GNL8gku+rakCEID4gD1e6syWJpCGC094A7t/ogoYE1bBSt9lS1KhYcfIS/lYjOIEsU
sxqEbLWW0I4r4f5/R412OpkqTqrqttksrneHKMswJFHs+c2bboj6/bkiwmpMaOf1HYwDj/qsvC2Q
XPBlRmIksY5MulXX+wNDEg6IuUV26k3+6uFrUcbs/pa/uh0KrRHywafedD0AyK3TuVFGo9TTmUMm
Uq8+FMmF5SzlUoaiRaBvcsmkunCxRoC4EmPoREXiX80Q4gbsSTxxrRoAb3ryvdzwFu6h9gqieq0c
Hmzjp+mxwJFvakMoB6W9QUQMtgd6/4lRN1nzNQwN0wny1mfc60jNJyf0Exr0ZFOWRstukH7dGKqP
ybZJ4RK/Nn7I5MiElZ2/kCEWaa3P9KCHE9nfs+I42/M15jJkrhc7lVSIBLEQE8I1lNEe039g2QH0
wvlLQfeLsAr6WJDj2PIMM6gMWcWzaugrIgCI73ACKTaHa8RSnF36fUmKq3ZjY9+DVNMteqtET67i
g0PlxEaW1ZjYy3/K68Gv5/VWXw5fJa+nFt2i++UdLER6gtf0bApZ5kodB0kC3pJXWWbm08qB7kCW
7dVdgE/gKNwOsRQdvmXbiu9sr32GBKJgoarfANYRebcqJ1r2wy03nCfOmcmqF1+ntQUfl1qb7d2R
mMQ4Gedovxb/BbkKI4u+KosKVK6QVGKyJ4Bn0uZ88/MWK8htI+Gu34UFX8kl9B+GTLhhyvAmHe9f
djHr59wF/JuMU9JsDx/j7X8pxSWtvftX1RffJ7CjRYeC3dl/A+4sDTBVizCl63KfnmgZiQrdHo1Q
SMXQOePrOxDLT898Nqi8NMvchKXruLIK6FA7YbmVkOvjMFqjJcq8DrC/SHKc2XvXw9uD4oxjq58R
uYbMnzN4eGaBO2HIABN8gjk9UBaShijEE1O7/MVhgVd2zB67/8ZaAS+JQRsy1WKB/C41pV1MBgYo
XNEU4bsjYdcmv38upt8ixLxLGDuAVmFigA/vkozX6fdHdFa88tgLJKA5VPp+TzccZ8+sBByjD4ls
mARyIQuqoBoOg/mtJO7fJimwHbh02CqZth8trX/SaDpA9K/KcmSIp1BTw/N2IRtbobbhfruLQMs0
yXnAfdmkxnou0wT8x4x9oIsZAnRgD3Zybrwp4Xh1FMYdrblXxSDm/+xocYF1ySQ9lBTULKkUn8xP
TPDiT/QPLsoEGgZz6+y9tlMeTti8wKESYs2vIh2ONvLpHRraoyjSZ9G9hOtxOUOOLoebh6UW1is8
D5o/N404VlaYLKeQYRNYU7jqbadEe7hrMgwWUVIn7jW2KK1ynx5vJ3xLNy+DPvMgzLkg4KCOjZc1
0cjJQpHUCpg4v+DdL4rMhvo78Wy58XkwQ4LFNC4tMhnnnAcF863fzdsepe/qvXDcykFUW1Vr2v0i
6jegdvlgB5KtBWAMCY/mll956rHSK0Wu/IbeeFXP4JA4Cs7d0PnOTykSSR/U6kjZM1cofm9wvEp2
+X8DW0Sj2YG4E0jgJ4Kxrpy8wwOiEgO38F26nl1Ffk99D5E7jdCigH1Z8dMm8KvctdGr3SKwRhFt
t/NekMtOEg+IP/BoDLwzYvdeGl7Wei6x3lfAKuotq/tcnjQsckcAZJDE5ZSGa530R3noPWnxJW9e
Xv2llgoeISDlyLqFgOvzU48Grozg+kqb2p8zJQq+GkEf5j96yMVxlDNKBLQaR+KcUzbQsMm4q7DX
94AtorJfkABnmxX+NcWrjLcPhVJpcIkjTJbXpwcvUWxO5WTpI7FIASkUu725An8Hjav0DC1EHZge
9+dZx3OXgc8I832Tm/WZ2kNVqv6Cxkc0MhrEpeFIwyH9IqvzXxSGTRccPgjgcnqMsXHxqj5t19Df
1ZBcPXFNxu86087hAujTFJxkyO42S0tUqWPntr8ZsWXwypTzHgkzchmB5OD7w9qh86fxnWpNvS2z
OfRFY4KWL0Vm8XOcya004APSvX+WHGwFVBJmkaA8LlO+2c8RlatECuBkWA+7tlyoAhnIJaHRYNyp
+K2s3u2zIxKoTpiHt8MWeB0gI3ok8dNe4Y44XWekymhEE5f3hvCyrcQfhV0xrLEnrUjvw2ttcLq7
HegyvCO0OjcRkKPiKYhJI5bcG+3cgzSvOqhsBg2UOWGMfNwJSmFrQZN5CCgvL0QSzPgNYZT1VH+s
JxfSw+IXIcuHzNdeTHxbK2sXpq9gn7OBkNYPby7AVyNO80BYggFrztultVS0iL9OHsxuAA8QhlS7
BkrGoVk3M/xcotkUc0P/OqUT3DiznVBY6/MVVtkJs60JiqJHgZWkQ0BRQO5cPo2p5bj0OVBI8v/r
3N4uVN5WZa0jOI3Ql+9sWQTs4VDC2slyC5zULsbGpGGDWAy6zFrFupu7O03AK8WaGbsA5UTZQQol
kpK2RH0oCyNTs2xi5LnPulsAOOmFv8aFPQlpsQLKr6G8YUeVBOChy4Opnrc6fJTEQ7K+rVEtbgsd
1JbGSE0rIT+kQMe5I/C+qrZy7hzTm2xVewifOKZTj43Td1VxszgQ4TNrcl0iAscBf8LNuGRsDmj5
pIopdtNiHNxK1tKuqB2pqCPQbjS/xtUCijYyNgQ2bsZeHlBUlZxlQnVNsP1YYpJW4RHm+xXvnn0M
IHRwQ319QZ+Y0EeGmiYZ0uszFp58aHFi4aIqJWYhd4yCykSBdEMA3jyJpsYfcpNc4jLo666S03Ex
4icA+uM/FG7ODo0UqWwnpwgwIayG438VXRaOPPAqA3hu9udjawjMQbUUdzVDGT4TB6YG0/D5O6+8
dEAeuJdJCZhGDihyF8Em6oMFlQeRlDx9ZjnCsKHgHGSPxv1/93je2T9yhYzObrW/Kg0PA8n07Npb
5dr6nkNLX4NuKlozOM96g7Uh1+2kD6L08qAlH7j6NaVJpdF5pYbXk8/7MBTLtHbYyeOS/+36e3s/
cZmFLAsqZWSeQAfRwm7dpL9iMWmWBRmwW37jWR05qY81VO6rcwmny1Cpk5oDM+EgO9S49akgOpLG
kw0kpHoP2dIqzDse/rGTRgZEDilmxkI8TNtVXF5lXGd8O0GioYRPNm09lbhxLfbi7C4u5Ejp/qvh
AxHRNVqexrULnaX2vQgOJ6PfJOb5cVqFpn/RV3bgsffBayNL9j2i10KojTWfH9UwXZeAHwlyTm8P
VZ+hG8O41aR5y2tG4miLZVIwfCzLQZizsoSfyXIA7SUgsG/3MZ1vqSanF07jrbSc9RFa8SRJx/Bu
EuQdTeBVLUTtIJNSPLRGuioj6RwBEoIvMxu41hr1fqIer7w2KSGLFhnvcl+55doA6lhAtUGP5Si6
LUfHXhd9cIgofJT2DSOovMpgmWcPFWKu5nJjCoNyb7dpo4BgJrj0bxIW+Lp3VPkidi0wbFyGBNRe
LBxKbygST9TAleT/Ev2CQSvoUgbWwvuuvRIKEDQDDD7q+mqdAgDKAY9JPSBoBmpBBHUf6Pq/uSO+
gjnAj3+RFq34l2MfaftSVHyCxOsekPxFFrOYMcKFP/CgbYwBMkhJbAO8elFUJbc+UNdWA/7eXUBd
lOO8ZZ/CfBHnGAKaoqciCrbeh5r4/FPcIGS9e4AstS5nvSsIYjaCBD3AjXTnI4x9tUhaBZOE3Efm
gGf3j1cvEy4qwvhYIdIdMhQF3WY6R7HLe+RIrSri2KJ87HXt6lJ9nEjII3/KWCWD6oAjWKIon0dU
BlwZNwXulJu8Ah+SyK7+7BxGCzAC3eXvld7J48dCXbGirMeK7HQ/OT+H0OVI3CZ92GP9DXckspVs
PpIdgUNbBeNm3RG3bqImpjv4bSUsaV1ngdKtJXudM4YDtoDnqR+gjD9AuS9GWWcsoni6N2uKFs/l
tBoxKrqImI1O6ibXPteDWwbttksuTCotCXz8eb2JNj3PUX852FgvtZmHfNlQQshLoOHqI46bCz4T
L8FSsQDml6H+4OLdG6Ap6rdXfFqRZZFGUNb/4tu8rwkanU+aPLxrSfueeocMJHdq4a4uBIbAOZuh
JsB2VLGRNOnJUekt/FVeJCPRRemCbAUw1iJzwA3DDrFb2HFar2GizMyBMCbOC1fsScZXwzV3Zh2x
B+NDiNHZZ3PSgekI/rUyxZ4GCcv4NT32R9GfPcOL3pQU0DyahRYUv/Dt/gS1RV7MZN2ug8pjMGW+
hAdfc2hWsB2YiKh1qYIQf+X5GecyhMRUVE9B/u1ggElabwVDU4MOft1LkK8qmhXtHLX/8RM7xWxX
rWvEhhpjM3X0yKww8EvPyuEBC7P9z9U7ea2VwVeWwtYYpmiWWhWDcJYxD1BteoOhgLzCtWPSkmcu
UTYcl49wJ8R3h8tyLrlaEJWFpK1kYMyDpISAyjjwEybYUyckANVRI3WigWo0RgmH3sA2gGB0c/yQ
C624Y308bfly/XdEFT+QfLO+Q7YevwosBLKk5JRwIL/hICT+UVPL9tHd7cEtL0isGFkeBS84sa5u
jBMe3kaIb7Sfx7Jge7jHA9/P6DL3m95ym2Rr5sY2XQhcNShwAsMdKxoC7bDpAhSn3F3zZnPNUZ6b
HZdi3/SOzQvn7pYokzifmwmF7NdcO2a/kMWJU3VaSoqqQV9HHqH82ISshms6/hXJ4hk95EbKd9Rs
dewDsSeNMILXp4D3ttivfvOWuXsLhSN85LC5o5VhUywIr8zKHLpWLvWRqJoB9ajZTMN7a8Vgx4fM
9+Jb5wPAWKuAO02QF9SJ/C5OrZ45Hrs1ThVBKleuzsQANEj8jsZgHG4nYFXzluxGsUdmubnIuxfJ
4dMgvbFTPTWuXrOvnyyKhx58i39MoJ61mHJ6vPaD0V97Fd6xGgEUxxG4wn7+OlAZveZcBo4JXNwI
jBC1iC9feSNHNd9aFUAzg4q/QF3Fs2W+YOqLTW8ZZsBZ2JWPeiIDr4wQl9vkHzkoEM84i1/CXrqS
Fur/QuRcrI+g1lWgsF4RS0xr3Xfb95FwdwPFcWJYkj/EsRtbAOD1LG/KVR5Wu/C6ZUg2/yomVd1Q
KJ2fqStPxK3Yf0WE5je9eyjn3NXIm73TmcLP1x1OOcRAfzklPz91s9janWFXMHxYYn3PCYjnOy5w
7VYLDj2e61733WGy4Xe0kc+dfgf0oW6QqnVgbHrZde43nkJ7Q1wwKNZVb2nOKRq+/fCqaQ/s0xHq
/0gFYPgkD/D5m2bKiSyGpPZzclxZewFgQSOK7AprKODwOT17A91sws1GZ57iStSCQ1/xutDgOhGZ
dH02e3uAl9aOuM33AmJTwMXt25oz30CjoQimpIcvLn46zuQqmf8tN7kbVFofDEqtB3MDw+ms1j+w
3aaNzAWDG0KJrrZZ+D2mLCvXpMd4aB5k2xWTBiInsgyI+yo2vczE1/9tmDQZxHaDm/VuAFkl16DL
OAl/TCt4h/vFUgOlayqyraHvlap5Dvc7T4RwPqipy3NHzaPd0sgyQg2NWmcK4qmfNYMmyYLBY01c
fuxMk34KnM0aWUO0fdyqknxYeXeYQKS2rfZ1PdmAH9kNgeQsBpOmjeOsnt4bsmqyztUSKSKZkwLc
VaXT0G9pcpD16oELgkXSt2qDmbFps/bz3aansKNMex8a9/HVegSSnzuYaxoSpaTKKo5oicdIfHal
0waxDQhRtIRcmxLp898z4oP58ENyfM2yeEZ6YAW3FG5Y2ZtSIGhPWTXiXOdK5Jv5L4D5scFPsqQK
0LTH2lTciGdZjXcLeTWtBSS+kBePdl8uNJpU6FL6IxhRhSmY6pPV9fbUtGYwM6jquYY/Hxw8JJdZ
WttRraaEowoJQkMHHGFaKqtuYmjHNvKVPNeUjRjfrLEm15QvPJYzSm5EF0zXyCiffA7bwW+pM/ZC
8PkF+tLSDzxeyxkE0WAqcqUfAfqLMH6x95Smv1qbqEc1hBiiOIo72QfCQTMtl/H7dFe9SRof08pK
OzZWVELOKxS6lHNUwWA1tbb/ts8oNlgFEQ2Ulkfy/AQeZqUc4Pq3LukB/QY5JTc5ov7k0Wq0JJsl
a37oj2A6BRle8QB8Yta/TR912fAoR/NMlo/QZNVm7h7TTGa0nPEvxlTvRbTYfePfhfp/Le7lbrdm
/ViDHm0G/0mdIEREcidvlI8MewnNWE7emt1tUQ0ndZWysde31ZGKSUQOU4maN13id74+4EmlEXIO
hyfoaUAaeAEbPaoanj1iIzaiHfbJVm+GL0SYEak791XGwDYGteVnxIbjS9htFxZn49Ik4+o9NuFp
wtmsq2fLK3bA4DqzfxO2N/00QmHyBdyncRNR78YzyqDkN+u/FKtz7Afck7vZFuYEEqXBffo+uVHB
B2HehfTK4J6S6YZ/yEYfAvDdXzUpHpinKcug2ijrTJyuruzWfXkptkmx8KQ7vdrXDY6xqpfhoWcN
FUNpYZEz2uxpSrN+AY3HbdgvSp9LOEAqcluGPE3/hfs3iR0M1fvMK7HiT0SPEwaUY1hYPrC6B+tH
zV/N5Bv27FEKoeieN+ndyFlO0fSI3JR2NG5JKxJw/N5C7vXiSgfI0YJrWzTOY3g2sQbM7DWiUWso
GH7K//fqS/u1/ijNXQRX6cjXjQMiLQ5Aj4cLmkWCYUB7NcdNPBqtCf3z5afFqYmFFWBymOfxUCbT
qO3J7x400PT6Jh1ZepujQMDlsrLYQtl222kg6qSqPl1irxY6Mv9P3eO33TycA4UUCm4sajlQpfK8
usLNZOf4Lxm7ogGcTjnBxBr27lQDF5X/1BdUVkvnkE/v/RvqBSLRya18MJeThvbrUre/V5Y4WVou
R5xUnJIBP1oKi0J8u47aQ1VZ8etBYGx/kP79sYUunZstK5IpJ5pTgl8DebkmcNu35elXK/KkVvt5
+YhazuTK2rO4dKWlX176zWWEBKVr9yf5IordbBv8NqCm4Jj0YmwmsLzyJv+gkhWOATEU4hCQItgp
KDT7tjjzyu2/u4JaTHPhjBQS9NxfctDz6xGMyvJDV+ELZKH1/Vgd5c/c4CwwmKeu1OU3tBA5ido5
zBYUKvDH4Cdl73uqPpyVFWoi8FHkgn9tmPZoU8TrrzDqP5Mg4fAgSQCar1gKuQVFE3vlZNbhfqqg
VMDkS2rZg6cfytzVr+qy1VAeCiJTV9GXWyhQjZ+xfz/D8HEpozYiNLadVyGFJSJoyfr5m+qgg7zH
LE6W33blpCxYocNGXeMX5trrY25jNELA8yW3hJy2o/dXDH4allTB7ykgKbopIGt+bCXS89oMPa5d
dXA+VgWcZj7NyON/MkFaUKfIknJrQAbdG4/DHRELUDaXfPhLhnzrx79EsBSOGaonYgtmzPN4WQ+K
76NsZcbvrx6/GqrUcxySGJf+Wc0b+1cTB71v7kyIqex5y9Ms7jfPDxF+gdXfGguONg+DUCHR80vy
VsLlpZnadW3lj/baBIpoQx8cuIbK0hFlDJ8t+2etZQ4JbWLL++WNBeB2Ri/nuBz9kQrIzSYV3Lla
mvol7N0msoqw1uVK3FIpXPWFdZiZLlH0OiUGypoTzMKC1k776HlmyUSC8KFXzEVhcSE8oHDeKILB
Z5SK2LpW/skOs3wGVL/w+m14eP+qbEyfc1HPBc8q7s86YDbvYjR8UwH3ovWL8rnxG+KdVeveyHas
HMyAWcNzSAn8KKg7c7viFL450Qv6jlbxNzZ/kl9Pi4Fpo3gqRAY0/dg9muoR2ftyabvr9EHAl1T5
Sdq8DOUsF8UkxJt/h/dWnjslUWhNy0ne9vx+4yOn6QetKrqlnhR9+2wZ09t4+vcoPo4YuY5gfKSj
qESSofrOZ7K7pPx7JV9BwRuB8gC6oqqI4bT8N6g0sFzlpOUQkTjki2G6bh5BrlFrnAkgSmMJAhv8
wSK9R5kCpuoWckAnePMT5t4AQyFt2rAVpIvE/EBlLOb3jTyKoctzkBuNHHwMQUQfHJlKJl/5KAGb
MUMjl5LA8UNBetl3y+VB1DMcZ6HVt36cQjp7xyOTd0gmaeN7TZ+pzD+4ilYaX97Tbqxr+wVtNreg
JykrcEDR19McqaQyEXT/MoS+0kMbU6qvyoaFP0rY9YsN+pGMOkPvHHUskFxfqkCmJopugn8V8cVT
4AI3DHfLUe98EP33Zz6vh/vDcTJ9yakPQ4MrSBcFAKgarQl0f0zzBxnhtzZTHTmXY+XiKO+4NT3Q
l52waUDMrxh9vtZ34m2gVVfU1hUQp7x8v9GcuFrJ1qEtjhFcC2R12x/e1DawgDrh7qHkTgremQdC
KncgBndADXbkN6gp5m/BS2tV0m4rxEtDSTcZ/DBq8p8yacn2QV6R8HiysrEgav4CpZEVFKrpf5DJ
9eZ9d7jxNj1SHr63PG7zW/Pcgp0axKwdZ0q/5uixscrGdAAOYaMvd6B8Srhkc1E/MZE/8He6mmwR
8lm3yKJgV6dVp9KbqNYxHbV5eC59byywo+MTIFJDIvimkN6XfVc5WA65tA1WK3HDu9MWd/mvrDHY
a0y8l2+ifx3KIbiH21WHxktE9f4J2iLAJTfcHmGvoW18ttbSSm9DVcH2uN2keA6rfEKTsEvMU8k1
l25c4pCGIvG+fAoMajuHUhgaxwsbd8fiXVJluIEk+w7uradaSujJqL/rfLQbRWDhbvcIqPjoaM6y
3c5tjmcl4hHAulh2W18Lxswf4K8yFA6JPIKLKQ72+hUC8dE2P9Inf0GAbe8wD0xTCzMSfx+JoIH3
bk+m7AP8gnsXyuoFz0qj0TTzcv2aU9mOwCu0r0F1C7PhONN4bO1oKVSTWr0mq+l4zP5Iljt81rwp
TfVH2pxsa4aEsC2sFK6szg+uB1LOecdoW5g9COoICDsjltmQj4ftRH/Y1XeguylgaKLesmwI5Pfp
8TZDTbMoJtmRJGW2Ypi3hnuV25E00j072Weib0l0FvYualpqlR4bmuAnXw9vCMUHcNx1UiVHFYiA
01ggpYGHmNyO5cKOLn/meSUt53p3XaaulCvpxMa0tRO/5EEm3MJSuFuwipobu+QBmUX/6dQxS54n
26mmCFSY0htIxP5XzHcC306loMvEyg6LHjUUR3SpAqhEME6llzWyHWt7pvsrLVsCPtOqXhoFgRxs
fwr5Yt58/lRLAh5NX7qcHrtay5Y9FGTzktpWoDaqSM+46pkUmWnXmbBebbUFoQpnlP8PeGakGK7D
C3OJuB4Drpf5PJUt3chpRqmxvk1qL32UZY6QzeS9wL0yiTEmzEPv3T5InYehYp2+ELK2SlNORw69
IbWIeD5D3pQopwDDB/H3jCdxyUMbm5xrslHbPiVcC7unWO7s/e28+AL1nq42JGAR2ezdL2gPaBmh
xSj2lQUZE+6I1P/0jHpXm5x5rEgC5E5sl3sPQxGnf6O0aioPDLKcd40Xtu1Rtm4Nfq/aLYSUtvtl
+WGYMyPmGfhFv3LQSNrmVLW1S9dknpoWVOZq1X4i9isciZoiKKkrQcRgHcoA46iiH4wD5LJBkMVA
Z3c5zahFtG/mbR/D/7LlXxxKMBH+KseJ9dY4lb5PzYr9UhWF2k4lPb1jN1+XDg4PjXY14rJxJ5Iv
rITnvwVW2cTasOKkyiASpL5Pbpy3qWWB2q0fZAZ0va0u8DWdrRIh80917ANU/OSMkV8Y5YUYAEGQ
IfAgcVvq6RL1qAIpX6RUuutdly7E+x2KnDDM9KUI8m1l5QCvacrfh/93SBbNtF5GOz4CXe/jOUKa
2eu6ucPS+NsyMAbzps6FzIVejf9IBZMGsfqAH04h66YqDDHGuWYsyGI1kxmdNcHVaJegzlsBCJJv
IW3jdmjyC+nEC0QtGlWE5Z9t+1qNaSpx1OJUDyweqHTgLh9S7NTXpgGn62wzA/8NJfuYKalzrFt0
RrFxuCIHtUq+3lau6ZSsaV7IB0UsTkxjZgna+3RXv27d8aLN4w13yVXi6mblY9uv1z7Hd4ZR0Qg4
x/sTAPsSXtIYwfD9sVr5iGAU1Fu3szlzXyYJz0lSf2txFzGTNGP1vtxMDXxiOl5h/5IZgHG2kTde
JOgSmIOVb2uwYXr8SpIPT8RJlSXCJonglBAYs5uu3Dxmz8roNoW0WW2x1e3Ec+gU0L/IemVhIVe3
QGgcaqlOLwTZosc6F9JAuXNW0SajO19sp2dmbugSai4n3o3L4GGn/IIR+O95AMDP/5R9mvnjI/9E
C/WLsUgvd09Ur/VBiL5NyuSPrg8FdgieWjk9cKaQ/OTHVoaoyaZ6bM3K82QPjnAgeF21BdW+JyvI
vDOUluwIEvpbU9oAgXJHtLut5eoKKfPTckh5IQJ6PaWR5hPOzckfRV8KfDgLZrK0TqGJZpinDl5L
Ve+jaJFyWCFAVH4+FLl0ycgI9Ys2gkhStu3tLoFp9IvjnLyEe4bAHptlkk984wsUko2pB1cMrRan
sAHSwsVFbF9LVexY0iD8TamrBqoFj50oeDDn1d7BE724NEdXStEb8vmePfdXYGvTqIG1ZAyE6seI
0UwY6+uP7PC38PPIZlpO1OqFOBDfEEO76gLBdiVuZ4BZt24LKuVEK9ACxBZkAaZqul+Jh3ogbVXs
FYVyC7RINfV2oiYPXGqov4nfknA+geyujHGlBTvBrfP7mGmht9Pg+Hcp+GWDe2/dBoc+QIcUhjTy
qgLNbvD3B3hZgWNAoefoGfKwIiR9NmrOXQusWL6kYOASge67CwmXNagxaSAsFgtg0eTLEiDu+fTB
Fu9V6Ps5nKX6sxfr2569+HEfGhbBWx2rEVt8QIDDAU2j7iOL90tYge+dRFXrsGGASqDolJokVmsk
VsUjpp4gS94OXDR+kN050rban24jDkOfpN/vPB8DFhokL9js/mKs3Pb4luATZYxpbHG59TMQ1fSj
dNPXIEbwyD5qTWsUPgtVwMo1c6wAIVCUAv2Am8XqQs1rPMSlVLuXbUZu1IBadoNB3ggdsMI4m1Zw
53tr0oiWGjXdHbq8koUR6q1X202bJjp7Iw3Cr/mUk9y5qfwa1xLu3RkK0RN3p0NvEDnS0irP4M0B
dngZ0r6G2Te60I4MpBfttHdjvjVMXtwhw29aXEIBnsI7mE98/Nz2GM/zM7QOdPteGJh+0V15o0Ue
wEZe26xEKqBKJREc3IgLGO9ON8a0o0Mtc24bDPVqxjeSjH1SgM8LDZFtYdj2XJx8+6if/0XFkgdm
R2yDBSmmnropm22SwJMFVlmRPwQY6xazorOtRhBorXrJ2sgrQHDX+6wHbo5n2aKq+u6GGzdQd3HM
lO2KhmoQWIrIlhZxPuk6cJ4KbsYQoTESBkNnMIrIBYDMMKXZs7i7DY2P5CF3W2c9UYTB00gbMWIg
anXc55lvw17ypg7MaEJ2pjiUPACzoS2eYA1NbfbA74w5eEoogoOUgE6fvnNIgkzkNYNjg1AFz/BX
3eTVBwvzQqvGLc04HO9hC32aO/v9GB0hUqbMtA5Wtru+uvphP4eXvdN6oamKo/7gizQl2OitPMFI
sBshSI8ADHMCvMe2kb1LswWZld04+MPFvO1Xhz6wiSxo3a8NEvjHUZaKZj5wPqJhiqIBa+aAwEJS
edUSkxDPQec80r8fwmAPxXOvne3r9O6RLgWr7chuulzXc2B2glTMnOxeKNHQVpObZbRgm1NUYalZ
5KowZJLLw+oQT+kZdDPXnaHeQZ2QVorUZGP4xG0ZcupoNT/m3tWLH2yuogdKkWZJswoakQyPbbDn
DSTkvd7u37VWt4brRzorBErkQ/IuHspWdcAmTv8n9tvjmsy1HXAAhRisqegZDmKN1OtTzXqJFpOs
P07AeeBAdHokBQuv/RuFnfv4z+7kYG/vjE+YWIXCyTJSg2UfInZ+TElZpmgQi6VaY2T69jyyWCZy
K/OevrK83/nhxkH9/VwyfkX5AG14Z38dHty0IY2cLnCGnjRVLzyJx8ao1BKnYx77f1wlod3OyPQH
XqA7e6IcenZ37NCjV7OtBBABk7X5A/WfWhwhRz6IqzDnezps+IUWcDuUkSuJr/EvQPZwHWxerzhw
dOp32TsSmq3ZLgaLqE3ITPIlKBqM8QBCDV0Y8xxmPpvpTwbhUYJy6ItI9jcXRdBYvbJFd9iOGaAa
OeZ6V+duNRIKrm4BxVrESf/6shQ2H6e4uK+UFg05XOtMXBf70ahpW9qcjlSbwwE9HCvMUwLvkfmF
Z8UxL9TAq9BfpBJmbHtavA/+NcRX4L+C4B6w/ANe8BnwpIJ4UNvI1T/gvTLECTXQ3PoovWceCJeY
4j7o6ILSPfUc7Kb4mfiB5+ckR2NS5fyTS6b3lO0wx8zhzhaw9CFHG/J+9KSZCHOH6+9tvNZA1SIM
RdNQZNQPa7i8ARCqA1W6Z68UL1azM/DrEv70P1znJ5He5LhEy6yNnKSUnWphdaS3uFxfcAjzWL4N
RdFPm79PEaASpTVmPEGrl6076zt0IVFXCc2qy5jPkXC8B7vKxZ2hIEykPtt1W4oBQfPPC4M8iu89
AOrD8sgtjTh686JB+tZR76iyHY7If1g1eFc4ZV8Gqt8SpO+VQGrhRLBbVAuSEMREq3OT35Frq3J5
49hxTb915YPfW7nuZ4+rW8UsFvUlMBQsZQFwymPw2/dtqKldeKxVNVRT7k+QBD1Z79hRdCFhND+Y
TpAfC03w+mQnEsImT4ZfxLj1yssIow/OoYpNJS3oigUmqV4OFfRgXSotikYGjeekjwnd4+7h4qx8
TT35gNC9OoFgCMRAQgW+uHBlRecCL0H4bV4t8XLr0seStfuw4cqpC0jA8aaoPft7t4O9r8hdAN3U
6wYsDQ63snBMEUSmv09By+c08c+VAZLLRhrRZD2GPUCRgGfPGaHC7xIlMQG6zEZIPoCjowqF0DWC
gl9nklULkVatiP1RK2YKgvCM5DOVdHCQnz0ZDE0LxxCBdo/sfy73gmXzyIx4k41SCrPIrb1Yvinu
t0KjVi43C54SUz/NNDxkf8EBeRl3n4d3qszKripBFM6fSVegtOnlogu+rWvyTYM2sL2ThXbNIJ62
f15HQMl1s5I+TwA1P82HFnOStqSJfpNMH6Vabynh3QYPr9fBvWgY2zWR4tSGnC+RWTxAtSR0Q05x
DletwmVmp88fstPxmV052qmWG/FjRJqEPngzPnthe2fa/+NWqsFPkA7MEeXSs49bJCrNxAMuOaf3
vphRjNvoqm9fGOgMiMgoIixwPrC8G/2gLsnpdt8Y+sZ5Du3lzvCgznMJu3TX0lq9JmUeYqGr9t4I
UxgPUsOU9Aze05rgCqugsLNWqtjDZyn0bSjYI95co6PENsCdkTrd/pLreaTKDcJSpMPlt328xQSZ
u6U1sPRhEURHioKnAGrDISzERHJMk176XijIex7eOeJWVTEX7J+KGRajo6CqxRT8h725TiHElCtI
Yu8jLgX2rc68ElIcFbWPU/ehn/qthyDS8bAsaQ40HpsCOi9YnRiRG7JNgOSXhi4xKTNkltKSRSb6
mviqGch8HRunseCbtR6BgQnpD+DIyWk63QU6F2QMqo1RLu+vFmN5Hm1XxrcdClTxFvD0N6PsTzRt
sppeHnwsMTKRe8Z74VqvBRrikL8ZUChIPukI+dy7T2UcQw6+aZx8DNpMtEq3nU/jTpUq1buQjxT0
f8i+aLpSK3fFoWgHzntWvl38JnQ23EpDDQTKs7WZyqQbEJyLIkbrczmyobXysJxVS8nYrrS0Xfuk
A2liJbDctMES8a7RPhu5YAABFwwdKB5yF75AlLg3R7/59L6BoSl7Wnhvba4KR2MQ7tUXkMXk1TNU
hIhMTfDa1hLzKgYzkU9HE4EVD/9FObyLwy1GmbeFa01Dg+8x+k1MWJ86xtkn0BqwglZJBkNWzTgZ
Y8l73KWjVJMszhNHB2b1ObCnfUutwYNvh25vjHtupYfRropExUUq0kMadbbYzUJGzPXNJPhiWycZ
azMiUg++OJHhlIFyESy7k2mXqoz4xNoHtE3zJSUQ2mLc37o26WV/uh9rOO5EhwdFMi6MA5tXgvPg
zfqbLkArJ6uBeQ0+zvdMJQnQ1m6t5iHYIvWh4QullVhhLX1bvcRxFmgrCUNW7vsodEMVQjBu5ZXT
+D1cDLTydBz7lqwZWai/IgKJoj/k6ty2uypQDQngpdgrXapdorSOINF91ve2I6fMzBrT1AsOh46Q
Z6jiJiWwaH9QZChBM/aJ8jpwajmO4ILKFvY+b4Kl4y5P0Hq7dpVKkZJu2+dfgjDoNfb1pAL9hTCP
BVcsZf69nD4xcl75dJZnewm5f8yDUltX/XgY8S+S3d88KLkNbVhgDDb33WP7ra3d1X5HtDstX8V9
juP0rfzK+cu1LAgs+m20ZtybyGRfiZ3LThXgQxuE/uuxyuLRZwD10s+pZiOlknVYbkHowdPSw+c8
DVSpYj9EpZnB/QPLpAaC+GHMPd15j+SysG5x2wOomF3gOALomkir4Ehp57Tzb0b/6Y21+DNbnVMe
H/uVuaeWlqAMJ5rp2h/fAgDmBVbXCE9O/5QE3FL5Pwa816XS7OiSiUxQUF1k2Spnx++J8Ezmh0J3
Zbtw1LgpZ/rv9GkYs7JaF1QnhdKwgk+iy6XjpqFmLNpUPb1Sbb51mSjmrVxSRXjBg4eszwQgSxnc
57ejBD/03PqJTpxfuFOQ1ZBlTVGMKwGQXnZ4dyLIfTlFV1n2ecxXzD4PDWD2TUs/n+9c4d8Tcvk/
ksAnwLg0fM1TSoQIe5sNoreeiVvV9TZwuVmbFJt/6jHLER4iwyCg1uHHqgv5bM9aPQZSUjagbYTB
a5Z5EUjBVJ1UHWivmPP1RAYH925L+xEfnaaKS7OVCD3fMYviAP+FkrWxthi2NK3TF5Iz2HRR9YG8
u8ExPAimhvzvFkLYUwgf8pHkNPh5Dk2YEoSqjbSvjpuf0wyMWR7fjQq92Qu5xruA15+pLKzzrcAS
tDPqz60Bi2pRAoVoMKkJeN3uUfsxB90NpCpourVqGrC7CtaqGU33VWHWL3E0LlqG87ym0Fx91GJz
W+yRH8yMxNBVXmk581E4nqVlivRDHdCwo9EbEG82uIpF+p6iZebPSxck/ewNlpbc0WMLjz5pEepT
9DiH3C+rbrSCx8HhSjvhVy+Hm1Snk1dF+YutTbuQLRp00eFgdH+dYWc9QyNJxyxPjtc2iHvZ0uQo
YxPFocR+kK9PKWiiL7HmK1f4XKt9MSOxP7eH+0O6o8w71Z1XaT245iqU8SHi2WQY1fvNeunifS5N
aAtkEXHhV0ueL1fpeKBBWDSfw9H5IbcqBC4bKeev89K3DMIDDduC+zP6xaQhPe6c/9mUrJBZfThy
mKMsxykPtvwFe17lG4ywtEW8urrsLOQ2KkXlr/5Vr60/gGoFEbvWQpyINAE8VOqFbKQA++JwHm3M
Uru6nxTL2UnEjaY3OzoUiLRagBsevZyolGBRmXjFjdSZt5LwAIwYds9mHk+BoAuMIVciup13hVYm
SttOHbGKjQMjcpVogZwZmfbT9C0dakghAuQ5tJsR7QbEUixB7oQJrR6dsk0ymOkFJmjmg3aQpA1p
rlkqdFfyTsB9UmH5WuctSK31HcpJdIY9jLD9XVGaAniEcxaF7q3auDfAu3oHbUNySwooa3VBjQ+S
2nJ/jVg8Tbkt2UKFZLooJ0ug1w/1GxJ2CTD7/zQo+rM2hQG7Db3p+yASrQ7gnUeoQ6F/7v+J1sgR
nFjOY0hGh9JVYRqVZ/XpJSmaBlk8ayemdRvYXcAlT6+rnrWl8D3u7W+ydXzJr0pr0zyBAb31G3uU
mFxZ0KmybPodVltNHXGfSyZQizacQBuF18NK2T8HaIDHH4S3qP3I/y7v5dycAhnV2V0APySDPSDd
ROutGIyG+Qyv0qifu4xXvawLkBPG1eN4RkiNa/OMfAH1UYWcoYn+i9uhJ3L6kfxnVI4/4jUVltAr
Eq38rp5BMpuQw4eF/qXnBs61EO8x21kYpJWxv5KhKj5Zdi3ANHhRdmtKoGZFA5UPgh3Ez72Q2OKa
chaVYv2KnnFOHF41i1e1Xstw3+j3qvKFZgxhkN05cod27LFaZ8seLofwO1eie7rzyO9EVc8oIjDx
7IOcqS84Woeh0x1vxy0vjn9eM7GQ5JD8wfRBWqIvSaRv8iOznZeLssHm5BX5r/X6lNfOnow+Smta
ZZQRc2blOTATJXH3JSPru286q9HPiCDMfyzy6y/uGl/rJ2qXBxhk+U0k3lsHFGr+Lz+//5gk6w+F
kCZysqrmb3G4F2Ln4ra4rGQZuh9PMzDJztCsIFPNx8E8wKgPBrnHLOfvJVHMMMVKemOo3p+5rnvv
9n7k8gQ1gOM/fOdmS7lXn3Ec09vbrMtUPfWCP8AAAT8LTXpAFypj0ypxb0XCfCv9d4HOSUiA6bed
xNKuIEuWkLHID4/vwSaXWO/bM51Q0e1CalRBaZzszgETZ35pIhr7KC5y7k6/2wOhvRbPIaDnp3h+
uVZ3X835A4jkc65EGBvULO13L6fBSlBab0vfwnauj078LtF2FVZiQNkzJb1BvPYBxfD/x5cjoMVX
2Qy08lrdCDDy7It2a5EBWWEKCW2xFxZ8VqTgdOcwe4yjv7Y/2y/PAw39711S3nSDhioDA46z4lx2
/t+uG0lTZPPxzUoXapT6tZCS7HYu+WZwEJzDigFc/OeprHMj/UgSejibqkGxHJIDei4x2CajsjMz
oUpN3fhG6pSlqMqDUgn3unNsVgoOyiEx8ZVqsiuznu5jopk0FkUqCIw/tdUChm10s9xel1L6wcpT
w5StWyGydlF7svGNClxQIA9VllTA2JugQhg7HKzAX67VkCsq691yQoxP3p3L1o3DWSpblfN+v6UD
FwLrztHDZH2swI72E/klPeH0/cPJ97M+UpN69nJUU7vZfHDSM/K8WHUH5DUM8hoUl19sDRe4SFmQ
lVO7FCR8JQ0Y/xmtnzoROBAkEZPDEHPW8Egc7MeRgVmFzuHVu3w1Y45yOF9JG9epptNObOv30Ywr
kVWE/u20DI5HFxM4X9W9m3wBOgNTw/iC+OcPsD02ut5hN/KyZKGWQxFlqYPAgPxYOacbgDIJiqiN
yId9ItUHOY9d+84WWyIETc51RJVTFM85mTBD/uCy1xAi0Trdc9DGwv6KmaPSJgUWZLwYgg+uV5t7
yFcHZ1TW7JqZGZIyhV8GU26BV/kmOFTTsDyFd6fmDBBxyV5D4XBThOcWFwwabi8X2uoUP9eq6kV6
LcPi5/Ka02j+befr1LRb6N0yW5xjMghICyNioTst6EzTjSGPFHjdTVBsg3uNSsnAGvHrE4IO4jy9
y5VLLwWNpha+DeLxiUNMJ3tl6KZkdMC2iyZukBjR7I5C7V3K4YnmCWMZFsyiVdVR4oGmv9lnIwJJ
/z0eQLyPivf2quA9+kdK+DEfbd9HC3Ko9VmpWT9035rga8BhKxSG5DkanVm1n/j8s6DH4ogI0BR7
qOhfRJ+Bx7CTrZlvjqhYBBovmCaeJfeo70NHV+gPPzsh2kfjFm/ffPaQb7qNleV9AY11De358yUL
BmgvX6EDyD1HTk2t7cOI9SFj2Y+/qXluBoXeNlOBfkXGl/wfuqmYVGH5fjjrt5a2Kqon6ZpuSAzN
C3UsPYnXRJ1xWiR5QJseW663wFjc0QAWWbJ+uzT/HPOlD/+2LMS+b474DXZeOdg9Tk/qUGIcy63f
SSn+mNCtXxvOUoIjrVGyfG23uBpXtWjzDxr2RaqgMi1woeWY2gbvYWn6bqHUZ80jI1gMWV6Gaxh/
zgccyr99mFqpxJRcvsiz0hz6KOZo7BJlcaqQ3DXNHwU1LdWVv8tLCmqoC6cDniQrcLcaCD60QhxB
jB3VwYwf2ZPAfJ86apGHEZRytsy9KSHjicWmQtdi6PMN/R3XVTkJp3SukUhe2kvK3h53TxRVIT5b
CJiNeagzzXOVevv6MI66bh5HddYBz4Qm30UCeAIAj5RP8cNc9Qy/moR7pckpOqTQY65/80rt+pAt
Jdxjz1LY3N3zRItSiueW15lzPoqhrnQ6wM4d8x3OmyqkQ9JUdwyjcrxzFmYLRVIrE2z3zdjsjO79
SX7GJPIWNV6yLptuz+RBgUDFmLJt/CPtiQMCCwrsJAnZTx9b9F1Tf804xBmIrtz1gTnKLGJ0b/yi
GB++BHAfr2SD6eeqxWLe1Ie3Z9KeA6MKvapNB0ygZ4VsWmZG5kaYQKNmw3v64h32WuhmlqBO2xGh
74CBU2nxY914E1EWPb1jquNfDaW4f9VHoKZx6zbkcr15+ZyHxIRuGLYTZM9d5fNFBqHaYALXDpkA
L3nxRgu+U8/PgUccSm4vwcO8ZvoDcb1YTQyS2I9VRm74/SnqHnZtOoFNAC+sxKOaEYGVbf6KO6z1
hPuhLfTVVzRApl9rO264JHelHMmzTaMs9RDKP7st6KTDFO5Rv9kSZ8OEKsTr94t9D1I6hpfB91Km
bafO6POCCVvspk2wqwOMVy1sUe5t5LrFiLIibv2DsMQ2MiGZf/PfR8UaXffNpL55t6a1zxFzL1K6
/q68xhlzI3bLL+Z5MWQZ2Yi0aUag7+38PArb7zLCIz9jHuBSzwRKW4Mka+XpCDSFnHOFHc/cuzu+
+drBD1IFs6XGDTTv5AuDdZkwoI7edinlcq/YpXZWQLoDdiSChBV7tJ9gRjEuKYAKhLCtAdJDGchh
AQ2YHs1QNyxaCfA+v6q9DlPalX/I67V3N2J02F4oBbXdXiplOCgRt8kzP6E8nrsk3KsmnWZjZzQi
Y7plSInPhgRj/wkKTOY1TGiQOAhtAwEXMksr+1q70QvOIusgtkNxpJbHbeeLTnTxNf8Njl6Znpov
pqy6rbt9GWtiDoy8RqJmqve+qTxUUnVkcTWPRbiYcApl2eqEnbn4ac8CHGUbIHMBN711Mzap3jqq
YuhmtFByqTqI9SPjdHuWawGIjjNv1dzJhmBOlISN8BqFx+W7Wt8WHhxDUUxz+p0TxApuHwxRZhM0
551OhO9GXMk4z1IWm/vAhEtGcSNBJF/BLABb4CeM14kYnF2UGB9haovmuCLyySDV4xX2oAcMm7OH
ZIuBsfhRymGxQOEtMlEfIv7nrvE/kHbIu5x7f+C1NGFejaCePWNfc+D4rFVbn9VGfZW3qPswXtAq
P+AtpoPDYRLocZAmeFpc5odXo9kBsVZG8jkHa7aEF8Het2RBYemu4XBuErna180xWVpWedlE6nv7
1O3lAcguPbfQeMcQ//3h9ai4rQa5sPDtSM68tKGzdsKaLMlXTGLt1cPqFMoQCM1ljv7LHjP5kYt/
gxq+81K+bjHwVka0+tUYSUOFnTbxcolA6dlYfM9TquMQfPVkzAsxKsMConEDLfXIM07rvvsBe2Ar
UCIyWgV+OcomMip/AIr21BY1Z5FXLQrIvbf9iLVhyK0Enr//oyRvDENpbJtiQizVm7gHCmVeOjtS
kit3E0o2uJkaUqnrVjyszv0wDaM3KPLlWMZLmza9zfTNH6hAT7PgM63F/wylyW27+47v/f2rsECh
AnDqLl16w6QKqDdrmuuwyjrIHe5WgCegb6ncVlvrd7Gi4Ht82hMLAqmTjnevR+jJ3xQfC5PWfbhC
nm5L3wrJWhqH+CE65i1ZX7a9YgWj+Y3zTSkfYECoMabugFci0ZVHejYHO1uwI8aLv5x7GVmiTAip
/c/mF/4YoSR2su1uNSJEKBc9Gss5KdHW8Oa2CjFiY7VAkSKdU+AUn/i7NTLPU9ZVdPsOm8yJ2/jk
x627Y/OtlWcyDkbu2bEwx08FU4FznTYwOnOedZ6WH8QWlSBkj8ymuVHpsFXuWGpWxkK25ACaIIGs
lgD+4qBzZjMyzeK+96cGeMbt6YhmUEmIr7hkElG/v50+2rv/HmuYAUsjH5ppGd+BqPWUIoN5HTo3
BvT8Aos0JG6z11lbpdv52vidAIWh73kvPUpExIz7qJdg3D/O0I9JzmT3H6gmwKY/04TQY12W0tan
PBRfTrTa4CIJZuv3QRAV4P3tPecII7nuFwRA9E6te6GJAmu99SlJbC5yzV3GX0wwtw8q4RmdbOzM
Kcadw1MmI4X3k/Lxd1R1lg6nKsR0KOZDA/Jepowpd+wCFec0agMULsPUrMNc/1zlzca7BD8al/FK
FP+1c0dCsMhMBNuV5a3IJxSIGF5GHSiNLFEMFTC45Ufz6oZRT83zj9Jlo9xnMFXI3Tbxw1oD2ZUM
J6qO7WSj5skZpUh6EVdhDhtL1YN1kMoHzyDIrDpVf0SbX9PCTQc9m0SurN2DSaQWHDJPnmpY+TS5
vG1D2WpQmuIkqIYZa2ccXmhl2zhqoLD4X2//miaysHmgzkYLJMTyxX+75vI3hGgRkKloabb64W8X
cYcVdg1Khna1Y725JyRxYovru47R+Sxmr8worzcaav9fggY1ssRSeZK/udREBjOqJu6EfppfovXF
sdqL+y2+GrX9Ol/3wpQRkBdXgGEaWcgODZx6ipTXC3SvHiMVwbX5olzsKd+A6FOIwUZB3rGlPkiT
7H59BdfCKN5fkn59+TstWSJ0cXkZfNKLViq2UfTgc/e/hKUghcxc78ppvEidLJuq27ESKkrTFNc+
kvpZVgug5GHdTTSmdHG+Kxpnw6L5bYP6VFc/teY1CfQd4szwscNKWFt3KqR6fXbHv2jryutQtzWJ
ZaPq9kbBOGFWpgMC8dwA1y22LTajExlTLqrrqDYkxXqxUxSVxseMKRCdPH+duPhLDorepeFh1unJ
FlMhxQRllK1OKC0f4opnF6bu5ZkbRD7nqjx4s6kZFeVst/sF/ry8jukzHfpNAsQuTfYqTJ/+on/u
oYdhWcTddKZwiIfv7noshE+pooi+VnxLR1M2Oo7/NFztptEA2FBKrZudnkCOUUmOF6QH8M76UPwZ
BG5QJUiogENNIXPrCEGpca99EZ6M9BVpDmQ9C7WGHCUQ8qls49DyBnrkng0aBv2F74tBbHlw7IOR
M2sEtYOphf5M+WQgJvI9oMyUc8MbAG/sSotHiOTAfkMVP1j/cK5XWJ+PXAEYMKInYD4VWUMTfGvm
bFFjn6/GY+yE5B7KbWRyr837x76VskGQitwkZ7KRTB/aOslQDE1/2VKhHYvPKoc2CFMaIEZclEqX
6hJe+lqYykjSbO/NsGMNciahMWsj5kTkSCwXCqhct/rSFerqMGa9dcOVIqswioHF9ssRLgKiurZk
u15BI3qN89dQfBrtXlb66l1cdCff6f8Uq8Xs8AwEtOCgvGGsk3zXaBOKyzTgCw65G6VXb1KJY+VE
j/7dW2TMBDTR1Qardu4Ow84J5iVszrRRhm1z+QzEsdKoVb3f1mlOI8LOdUHq0COQBVm9MqONWpKd
j+LpjS05FlZqNhccl+gs5pNEDEyOr6L2FMkFWOEej/3hiiSARCOxtnQ6s+uTVi825744g0viylot
W2oe7jGIbsqLd/BWzEtmIyAa1e8gUca+7kYZIyytYrxvKcfG6oJNZItITYXviWHlKTFsHaeNGI4s
fP1xJSVhXSdKzuZvezjOQ26KoKkXvQ4UBF4zrD+Qhh9SL9XNbhrIL1qDrPJ167IekPky3l1j9JtQ
bQ+8RK7Rwev09s5J3vYf2GOmYzL5YhEq9YsjuQkViVjQCih84NF9GmrlfIBa+fA+cpHz9HjEenLQ
+G+NCkMR23xKPUAgLlGQjiWi8gUkfksfFZpW3l3H1tUkiIX94zvOt1SEroDSt0DhTvwuPHdAfrKn
h8C6EHB5ZzIxj/+znNonV62FMGq2eCKktRWco8iINuTwPa/KnAAUypInXN1qjuQ6HQ/Mo7tBoTY7
BEcUnyNltHe+Y6kPvg4CAyXPlW+NBTpEpkY/+IwdcaM744Ap0ixk2wEYDIo6NJ4GsK0eAHJ+C1En
RBW9w45yO2Vwc3hGolOpUXUMoZ0CK8amVuc8uW+xe0Xy3+qz8fRsO1mFKL/LtObXW55fBdq2pESm
zkaztiRIg36Ys2pVEcnXFGOcT6ukrLghG9P0T7vA3NQG8wlqFbKt0VW2XKXrZ416+SYIEpj/NJDs
g5p7nxqNz6nv55oYaX62JPRVp8ptJnw3ghMJESIj0GYtNMC3vlziZ34icKAzL0xCjlZ7HUj3fPb1
SJYvxDwU3QRiIIkWNQJuZg/+OXqjARYrQco/7sFhOC34wIQnYdL1nmTByYoc44B4C/VNEPh3mBGo
YkG/r3h+1bCm7FtzwUAMh00s4dM9hBRQ8IcCOhaZHVddhQSUrURSCKyqnwgRAutHfVwxDfBGHAyD
zB6ycJtzD/AYyjcNMMn061c5Z7uDKV4GANuEfKm7CF0FVcHSwyuZ26xNSNkn0jREWdd/+l6qwdvk
f+MHAWz3Dph6jOgHZtj0aO36HXk/XcsDpHzOkXJF16AuAv61nmSgP8BVKhwddefq3aVO9TrE7dOm
brcYIEmhu+8KdNTp4WLjG2BtbcZ7RK7QeirlN+G19zhSSbDCxRc3hU3wlrhWkI/dUVPgYRhRo3GZ
tSs+72yKHk7LrQy6mh/CO3pZ/xnLA3t66SWjC2mjPwxFecGXsKRYYFubzDvU4cs0TCYIjI9CZiJW
88px3l76rUcpNhxSkipCYje4F7jvoGriRFEEfS6hKXw6zZVGNeKcN715CR0NWcOEIen08CqYOcP9
bolk57oaJU5qVauz/5AT7LKIx7Kbi0YTjYoYrskgzVR60E8uoah8SjvQgeYM4/3Gx+0QSVYyMJnS
DA18i23BBMUj/0oSFRcQ0D05/5FQ45dN/MQ3jmioQnuPfNWIV/yAUtnfE25kt/kyNxxmzs6byMMl
K/7JLrS+z/JSFRj6vSp148YC9GGDiEa/mpi5h6c8yCeNohKM9NWgKarsAZLMhWBEdzFMZfM3vtEW
7l+Q8V8zamu02HiT9QvWM8E9/KgRA+p2qI3aB1t0DE+Z/1MUh6IauNhxQYu/EAY/B8DnkDfHP5Kz
uhX8cpLkpYJ8M+6IgmehndGS9BnbrnBnBqbZ71kEzK7EqIIHJIyHu/vhCo9rU4ax3D6OPb9oEhtT
AcRxFb1fJJT6H7c+LY+zbfaaC56DWaldb7NqYOS1YhhWTg2OYmM7LtwE0pGzCocPMTgo7EmRCE70
Qeu1T2NNgeeLo2n6YoirzXV+IoHWLJDtSwABl8xDp4bjWOR+Y3LRU3GeFl8B+otaCSdyvihEt+ww
o+1jpNnvdGPRuoJqPVfUDPgo/WtvWN5e20IjoqRPMWDkKyDlNdV7eNfqiYUUGjUbWmHqzsUb2ivD
5m4cnOiY+8HvWHGcUK1t6fkMhOqaeCdhAAjXszOlA0OZqPGMtCFxj/k2mRhsNdqMZDndp8RLzO/q
f5x8zvui26m/D/j6Jwlw1eNrJGwn2yjB3PgTCDi7E/Bp0SxLuoP+fSHyRWu1qrZecfLNWX+hEgoU
o0dqxtasDqfbxtsr6HB8ljHdi+4TTNFlePQEX0QJphRhYcaaJvHjofS8hZ7PPnuLrrFbeUpXElRJ
esEEr5bhjBujjhoCRfRpwl/BF4P/iMGe9LbUDCgaraXNC2AJoSO/5DEz0uNRdTg6+vMyYtEAm15f
HRbG3YVHiw33PSE2RPEP9Zqm6qYUUvsoUKlTTyN818difYGyEL1eUVDclUKiQUl1pcQD/RSsb6oC
j4R1wnFyO2fYTeTeLEP3MwxuzY9hjTUtR/szHrS+xXTjpjJndZxipNc16iVIwqr/0jYPYrpqpZOg
gYZ+Pnf5yc/+oOuMupjOrFXvLlkBzDzMuVgpZj2DcRcNad4y2brjH22Mg/iSF+nfsHtb8k41M8/M
WOXpH01nrQ7dXt6dExLNi1Tx9fglIP7yCNPsejICinhqwC2Sr/KtF4mH4NXL3pC7WKW8Bz/S7UNg
Y4pVIO45uOnxQhTGQu250+Y8syL8TrtVYUJ5ZcZb25TajkXv+9guwInTihqaAzojiQ99KSWnxiyo
Im2DBabkx79fLujbDRKVCxfB8UeZc21t25PEl/uEEC2X3E3Yge1YDUDd/ok5hb1MWRP0+0a2RgmU
CI7wXRzMyt9A14rudNKaQGTO3rM6h7dBWG1Pmymd6A8i1OfhfHYpAtQzfp4/SpVme4L39a9PL/HT
g1po5pc8JEh3mQilLOi4fl2bPInjJP1T76Kx3Hvx4UwVBXStG8wYybsuZldJdOl7JWes2EyPKAby
M2sy9TCXZjdy8nlfBrjgqrQFP0iyoYvOl1sFfuyES6Ize+KKlzkwf7Tx9x7NgGu6SuuWvTp/MIPP
R3opefRmQ+8FfLB9ntvYWZcpG0/687p8nQpJGTkqjl0GgW0z/wL9PWJvVnKcCi5EBCnLAcnnI44a
ofSJI9799I49ARRHpGhhnMI4c4xs05cB58vOJnIJ24xtXPD6OBChPlDgpN6nQVHiaMETbFbKvFLe
JLw5C9J+wc+bNRTFyRuQ90u/N3AZky14tRuHreCNH8poh+nEGchL1hcHD+0u6xxLGOrrzPnNvwWa
7Vlnar/TqrOhRveOd0XyC13cn/3+dkgB5cmpdFnQr4e3nLnMon2vz88cUpd0YbyBRrMYWkpdpphQ
2s2dQG/ZN5WwUQgPB9ZY7J9oRwrRIfdGreSgu8LCuSQ1bDw42ng7DCNtgkOSoha18g72FaTxvW+B
Z5p2n+B9wOlbtRNQY76XIA0vBsf/Tr/PeJfOLOc1gXeZ7hu15+6rPVCnP4cxGGF38Tfw0Jr0XxwH
is+G0B9u5s7SUYAWbIA0gY2aic0IjbMRMvjvPQCE++92owbjoTfmPkAETDG7bauzZmk7v+AXMuz2
FO6gYpMtDiXHwb5GI2pC9YgYUQ1/gj30Q81orLOp/U1JEsO7ZgRwxIJxg7/sMKnTO1Uzbl0v+Pf4
DoIPd5p4MEZQZbgyx7Drl2uX04vHWCvwr5WSzCUuK7kM/EXxvlizJVgottB24apAQpEGCx4rO3Ty
EEIGZujCyTJsBVXX6kLWtsH1+3I1y+wJoZxklQqPMIYL3sq7+g79bke0B1k4ybIp1DURkpgDSq4M
hdkdRbNV9Sk3DcoE2kGqMjEMChg/uHHBOsya2jzDJQbkck6dCGn4gGED0vPbqfG4AVE0nXwTLW1X
SpIH6hQjxs+A5RdCMZ2l8MasojY515rYNZdTgtPQu7rzrAKXpe1jaL+DAnI6oUz/0bJULN73kH+k
pzabjDAoVvJpGAWJOApG3lXbHIA2qjo2tkJB8JByRA64Y9FnVFpdvT6E+iTPpOxsXWvtcQ2cHmIv
LLVZYxGV+uW199+Dh6wugat5oFj/N5TOGXtOJEyDzouuHUt3XObePerSbFED2pz5K+y2Z7oYjEBl
K3Rmf48yV2PnGhUSbfmMXbbbRCvYpy/UB0AfbkoQQqUeAzHjFMD3JTBFPtffqXaF+DpHN8VbtjxZ
w5XXoBw+PV4Gd+TipyykZQv3LNDpJnXP+k7hs9XhDdeJaIphE7IljEnwySedWnosEHXUkAKkgyBt
sgvU3OPTUOpwz/C31cgTN6MaO+C9ftO1EyK+3dRI9fkcT8b6H+ZD3YENrlsxsU45iIuDsM4eRzsl
3PBgPyePp66F6o1oYC5pWvdOZrDeBY13TFw14QQ1+yLG0DslYLZyM3tpRI0ePQZEKTN7iN/aXwV7
UkaM50bI89w6Vy7BsLd5k98qd6iSeD57dTD33xBYLCW6gwcjPJfwNCSDVywisWi7R2dAsUwu+3k0
2ixIH/5RQBePc0S7/AjWI2cetyg+Oh9EgsG3yr4Nq54r40kqbbyttQkhyDZZKJoHTsetiLXSVSOo
IbLYVXwnwDeqYapoODneYuGaQeyxLUDJD3kW9YjmKx96SJzKEdgKmx0ofLdFBepfTKt6BlyNKC0Q
2UsMcMSKHLXgzufYj2wdHZHFmomoFjvUQcHa2RtIpQZ6E7CjHQssnzeCZaxBBcvaeohBPsVh6WaG
61l49hZ/9g97A2mmH9CmcAPLIdf5gl/OdyP7rHjfgqFMvhMIcLIMeIiQlNQP+ZD96sKljo7SlJJ0
lSc1cbu5W7CL/q9c24mMrxp5FMcaQ/XNiZZLV4LbjRijQb+Q2CdwB/Vq8a+br0RySbeqg09NiR4w
9xJKBLKJ6tJHwVbZAYOfDbSeNTatWaDHweLDU99ubfxNX2aeqNv/gnD0XoHNloTKs3Rk2gjU3yQ7
df7udi1xQBKU3YdC8qkZxTtcBT/4dyOx30S4nbu9mFRhnp0UbftIKPvb2mvnONvDgL5rPp+RNCUh
jMzrdFj/obl2oldmroZ16ofAUKUD+0CcvapIzzANPdj0JA5UXFLX+qvyCKqrzz40p6VAVnEfa7M/
m+TdLKcJY7vuzthOdxLPQNQ2R9E8sIs4QJBdjb6EineUamKfTG7jJ8cVZ3HkgfdhIuFLDg/UBM/3
objjCDu20yUVeW/D3p9xLpMbEgZBxlUB84TeAywIxKH71uO6YzmzbtGlpyubdwuMZNxQPrAsZYl1
mLxkTDCWRJjnmOlhH/CT9rGf9nKnnsQacdUr7Brd9tmyiTQxCycua7azQ3HCWxz7CHdIsU+DcL0M
1fTEq63t7u1C0QQv+4HlrDovgCzXFYgpQjZnR+HJOccYvzOThEpX58ZVtm0AQrk1fycJoSBWVAVg
VY2OoaZMrmKyuH1tFmzxVj+om620CAkezw71+82V1Xgl3pmotY3BS9JcNA01x/eMelHs47ZGYQpd
sXB3NT/CHQpNIYjUn6fQCYLk53QZOav9upVb3kPPi8I7z8AommGecwkKfuPzrk/RgEeE4bgzYy9S
JdRZYYR706l+qij6w6/BQoxDVXzKRIpR60RmHvaPKIZ3IMWtk5+Rxdm9mENAEnMWAXgOOLa9uVf9
hYHdON0e/YI0veYaRLx5f397nLVQ2umvLjMXFO9CUTdQhHZW+sVGZsuRqSwZakWtRWOjEQyzRy2R
2PB+hxm9N/ZI1nJqcHLsxHVHv+NBfKzlUtbkgx263bXHhycqKqP14dq7qQmi1uRYSy2Sgkx2LHHj
URr6D+/l4tgfKERT/Jx18cD/xFAdVIVfXaZXmSHCXApoGVfnjyXPtGR2r3LR51/w2VO6It2+JBtu
CRyme6o6w1Tm9Gu5ENq5Z/mT7fWk4wIAoFapbQFUgkx1FxQVci5FtgQpeqF9IZG8bqcOxWM40vGw
JB+iHhHxxWzpEY+m6npnzxQdsLzhIPEIB6ojh/OpI+HdZLoXFMJ7Pc43mpmyqbX99uhjmjxUSj9C
6yMSFzolGFJT/e5QINnalYsY/xp7+i1AvsUCxC2iTtnCCFnfOt9visNbhNDiC5Wb8Nl5Hj6ZX1Ce
9MusSO2i/Wqagqs/oxGRpbFcorDK4fxUPsHumQknQVBGFLZ+IIQMDaOJGsS3OJf3rYUbaZReLQ1P
Sngtp7ndtSo3AnTK21Yj7qDUzDoXC8zIEnqv8FgRspwh26ViWRbSwqSdKv4sKzyM9kzPKBQ/MT4U
5kx50UZ3O1Vu2/pQ9zPuCMABVU9qMDZ1/mg9G6i6RbZuP+kGktguI69OUrsstsMtNpEkhbyaNjiS
HhKKn/Z2LRSKhJhQJYsCxOhe6LDjuBF/8L8JtrQjAmCxd1hgh9ZwrhLpaQewpbZd+cwxKmuYX/lL
UIsbecN80lOKIIWNxLhgZq+mXgnOQbp7vlKZE63nsE7Kz+jy23cxH6OTbnco2jP1iyqQYc9d9WcE
58/C8up5kRrMSuFvK9f8AO7agLRWoWL0G1BRzyHMInB6l8EPdWIszDwcTUfWqYXnLw3n6RPPybIF
EHPV+fyQFB8xcv5hyDyiBaz4/4H3qjjY5qroA0fCSYhl477H0LZkCGRAhnsHeJCDQ1BwLt4aTTj7
y4XQBHDYJLeX6RMivYZKgy4jmZNUS791URBqngFhrPD4YaGGb7B7HVSCoWtQKrSE3fzus17tJ3dQ
9KtARA5gZNBjxbzxlIdOJDekxvDv4z063z5vbU3/GSmW1IwFCruCH26wwS8uLVD06FYg9AKE4N3O
CsE0f+KQYHz99i/9Sor1aMceCHZ5hpG+Qka8hPqerF/jI2Hh9UDIhhyIIINfGCpUeAZ4BwNuzX52
DiL1T6MLO8eoEfuVfvwbb3wlHex4R00z+OqEP8ci2X/3EFjeDjG85o4KZEadhL0VQZDs73KPbZVH
HkMvzt+9G0OUpLOLsgOnZ44l9eESsXeNQlJMCrJCFrN1dIENE5ewdXwObefWaYtcUdia5sJbcutf
K1C7my6KWdfb2HZPz5Pen6onZi3ZmjDV76tJgsZ1eKe5TmkRxhK77KeZ4Y3s3XFE1xA+mZnN+uER
II38xtaIu4EUI/aRUg2Is0QF3njQRQhPSZd9bq5wNv7dMnZ3cyb0b8qYT6GysfNqbz6ZQiqtfSXx
hsaT/0J/tyZZ8tmwPmHsLA+HYPlpldOMlB8lSZ37NxJs6uv2OlSWIqmhC43iKzf5St7NbkfIbQph
GUOBxxU3dUybZYIRjT6J/nM7S1Qr21woPnBwiC+dZHVzhqna8by65YRZQq3s/lsz326zKZpYNmAy
exdKKDOODays5o0Zbbo0MqDPlUJFmKqw91VUywl4oNV56QgK5JH/g/JCrYKfnBe4lXrP/U3Qe7PO
by/hC5qo+A3WfY4a66p270kaPG9KVM7ok09j5rMHQfDvKA0oBi9+iNS2kzoMBIA7F228feWyfYFr
LLVeg0zUh0F3D8q1gwZGQ0OMfQqOV5gTluwY9Jmt4p/PVxR5Xkn+YsNVyDOVkseTFh5FxzkSUTCN
qzbWJvWHuk1CDhPWl895h66hQJUWjOX3w36/K/j6096plXJRsTdjhPnWtxbZK28jQQmlMpwAZntK
DtrruHUwhsc9+IVaHiaf9q7X+IZjqqL88dVWqgemg1hI1PNR/KAegb5j8GLZJXd7IycfnLjfZh6b
KfOebeOrZECNmFDPFPXhm26qOacLb8vYRImjWf1X3mKgsqJxEAk/tWuVT7KHUBfpsoxh+t+Jy6z1
+X9RzJEaMw2h/BS5Gz6m/il7Dw1QXJMdyF34DeOV6sAFzuTaDh3/4mKYmQ744Y24P4OaXDfmuKsG
4t3qyOqxY+Uzsles4dCOdTJ0mi2Q5tP791iHvxrFjvBfuaEAUWmkO3EPmp+zJ0ciiegW0cfUnxui
5Bb0ynZgzVlnpuJU9HmNydUEm0/3KFzl4J7iSVThrqMP4PpY0W6j7H8GlHXVzA2C6vd4dOogwjBh
u9GQbX39JP84q24wJdLoKsNQB2qqqr2nJrTmYHYz5KDCo6RhgGqrvlRcm8k8q6CWV9Fm5pxKYoQo
cB/BSaepF1bcZKR+CCtaZ2KzBaZhH/o9iT507W4mQXns0Y3tRwOIIvV+wcJ7hO/OZ5PU7vfV1PzV
BZhZ9exfZ3paxCEh+4S7CGqmkZzAl3ciZhGOBsOh5pLqgBQREWM2OhMhjphnmxAMN8wtu+ey8lz/
aZi30553KcDHp4WD0Hz8qKBd88byMrmv72Kmt+3xF9ShskO4NqoihaKann2DF/mXfTrkl5tLAjln
pmagZjbdI71d75k/OWX/duR+qmZJ7ENvmzI/F8uubr4RTQxi+1LVeCtpX5ZG0yt/59Mha869eaxL
8t/dFIYlJlGxiONFYG+N353YrpDNIuOEBx3OadCSw4/JNCJETkRixW3lAgw5g0jcsLDrh33Ztzq3
/HdPGbpTV/MPh+sUaaNTlh74RWe9o9fAGpQdJFG+8M2nHZv9prkL2fwdaP5rfFZo9yTSuFmxVdBw
LELBw4OtLZiD1T02AvOWnA/i1NRdIiIerf5KE77SPAi6MEYzJdZMUhlWxplKO6jqUaBJO8V8O/Zi
YfqmbQSxcawpZtCgrMvs+8rUf47Zj1vH777AEeZ1SOIn+xeSan31b6l7dTAY8xoKbGHLT1k5r2ov
y8fprDtxFu2AwcnjGl7hWUdJ9kEVkFqo9/9y/E4nFZLWQWN+e12N/MKe/VoAZLXyxgwOZAvKRGG7
313JqIobDimOSVs6DB7Ju1R/QKmqc+FPd5QyMFmOEP0K/mMsqrziDQwiD1nI7QmH9C6ylsA11/dI
RuuyeDyToggeiITIUHgIQvPsP/oNqX0eT4zUeHPt5T643Gm1bpZIdzQ4W0OoHz93YvebspykRs6o
l1YZwPJQ2a0OQ5gPKwswkqD+HVADVoJrMOLuSpq/7p1JEY+VBodwkIXAjK4eQYr03MiozQYrmMo3
IXsrtGiuW1zGmKANOnuj+rLy5vHg0kot4BQdKI4tCys/X7S0hm3R1Zec8BMZ49WLhz4tPhBlpooI
RF9JgnXuZilMDk6Ae/6jrrhvTydys/m/YYyKWsP8wTO9wF9B3I878V1e6ycAgJ1lhIsyMFNv7Y+D
/WXawkLfXl2P46b7v2HxLAkIjQQi2PcobUVdEdQEcPI14sBHzCA3YzE4r/hrL8IJZ/YqL8fPJSYA
bohVx2jd1WOgI5kdFBlqQLUb0lZx0jRSo/PlUetVqSdrE+4+/ajLMiDtaJ8jcQN/wNVPixamgVqu
0vWBGDqFmi3CzyJ+DOXrqH+2/FS5E2fAq64e0uyBF5Cic8oGDE6H5YY5WVUMC8p18MS4a843IwpW
xQzLkL0yAK+VrywI88Io3GAag1+WV9mTjhLKFh+W2HDiGIJlGrfsLyYQAheRqIkQPfBaJBW3hZ6+
RfhXlRQ5M3LnP7fN94Z0BixoXhMNM0+DULR+A0sFVHAb8nUGAxTHb1tLu1/dx83+eB2IocmvV+Gl
cku9pizpO3NJmYC74FF8cOgFh1+b0f1KvooPPvdUY+fsu6LnY0xrOCHg5m/SHQGTg16jvLd56ASl
lacZZT7Dk+3wxuifYresAaCsYIliJ+p/5/JTztliI2HBx6LV2ulLxqrAUY+LkuJPoveD5CTd0M9h
aYOBP3YmHWnAr8IiQ5161YhnWb5oba9qOyNMUmgYYz92wnrx7qxyNwYAN51pP7Or/d01+2u4/hIw
RdfLcmBqPUD0VOKRRsE/iDdi/miZhrx1qYaWtA3+7Obg6Xknw5PxlUGksWfG+wc83IWFvY8i7Kmh
0Lh4dWx6d21FhNSXtHfz50LSS7112/fuonRwsa8cwn/Hr+w1auMIIikCnnmQsVD3y836k+LlyZXi
yUtl7GbC18pH85RbnXIuqQcbptcIV9Jc9cV5S+xOG8ee9fV+b8ESvJSB6ccOtxQE90vXQSGBfxV+
Nh5nKl1EQsGPQh8KGWlpL5ovTQJGJsBaziiUw8yx7i9Rc3M6w6qGChT6iZHRhlM+zqbm22C9+3bZ
WSLpG10c5Cy8XC3dnT+xJYBWpUy/HgrFOvCcGovMp+WODe2c1KcRrDlGkjhNlEXUAdOGdcUpxeDo
w/Cv3PBn9owZt4lBJ+3lLoA1FK2ySsnpHr9xAIwAb2GlPw809Jddq52PNf1AIFXW24EiVDl1EUBe
Oqknf87D5Ot7cuJKzWaY8t/o7QqqqNPuAP+lZzuSWbkND1KOEsZCC7etFM73vsYF5OO65A6XeY97
W5/1upevWVsJZo0Of5iHZIwMoz+G2FPZ7XuklN0uQOQZAPqDKJl1kWRj5EGsdICKqR1O3npnF4sR
L9SuKjPumbPMq2AklwjV2bIRtZFhqFZqshQHynfgevAAZZzTgJaDzaK6Z3FTsG27UB0qKfyDA+Qm
e2zQuiKVFjV8h9PnFNXQleCE6R4nQAaGtvJBn8KVL2rXVVQVAAekPfeUY4d5VaXVT3M5t/6TqbW6
IQHHHlQfhlxrqvjIgjVrjhtDc8CJnrzQIYsZChta6r0Gm9X/8Qa9NZMfdTrVjcW5gIoCAsfl1h1H
qy8sCvPvuKtEDke4YRCJJjqTOQTq6VsNc8rhFHs/t7kBMQ5vQGle5J4CVzM+BTa24nvKNRBUSJ6t
qqmQCuYtbHwdV7N8F4cG20QVp3xsUM/eH7wdjPN8ucx92THjQF2TTq1PZ4thaKikyEd9jjndi4of
WSy1yVJ1oEKAyi0cvYW+FAPjZH3/Y5Jw2AYBE280tgBB7uzsh7h/1du9Jap/C+4VnimduiOidFfi
qop13Li2ACE7Eygxg0hvorh+SVKgEsmx/gjbZI2Wh1aNLjv5SB73xVFEiiACPTRR9aaUXnlV78Od
62T7C0ikXTLWH+WkWhrGa/URXIczOlKUwOxHZ+20xjvOacPwizWDmCwxklyui+WmzhQoG89GV8y5
buaxJMsmX2d53VCHS7fXn6CTKBTb+RWSu8YHMunDdZl++rYhE1u1LeBz8iuA8YkdkpGziVhmglCw
Tu7fPjO1K33mWX2y7VaLIPOXWRjLvFHdS3mmbKFST4WTsXl8B26J2eQ5aOfPvSNYzNMgtpvd2R5p
1xe189ZKyzY/ikN3bw86tJfwj6J6htrIDRD/RTuCLyuwmyMTJxO92XGy7Q4+eOqCxfidN+3krWBX
HI1UN2hhMu9iomvGl8agTMVkOZT4v6R8NblXL8D98Cz+ajZTIAGvf7GdmYw8Buq5CG3QHFjl2c7l
HRp501qUP9lqzgkmvCKjCGOazALxiBhRc9nO2fknvkEXR1zcJyPjeSnDJuXsY2FMc49NI5pmbvyy
0+q1mUvZ9GliZhHcmrDd3zV8GtRuLivktQGSZqKxSsJS246+SvEzlQvojmv0+N8Z2UubkddGQCYh
lU2LDpYoaqPW/3KmikX7KGyQvjP7Csxqumu5v2yB8iOd0MyvDkJJXWNfEoJU3/LvyFajMMj5H7Tm
Ps0+wgztCIJfQvq+uMNk9Y65NEonjOC7O1EccDzRbOURwuJiR8GHsoX7WkLpaueAd0e8IUKYktqY
7FBo2ZupmAB2ftZ0qI33FHT8YquE//Fhb88QY2aRXglQQwMn8zA+T1A0QR7nUwo5hbhsYLJQYtdL
iNlSJPdSiaClBUxuDlqqGXYHkOTpQ/qdY7AMOqirE8U32i92V8W+F8kzzLKunfxThnOmNxcgTcHC
Ne4o45qaMAmVPGoCl6eaIZNhtAn2ValpCfSj5M5dbAagB32WrQRlPp1xRTGy95c3X/UJrVgb8AjO
c0BlPXNHSVeYam2ajNpgvt4+0HTvtUCHMdRaDqgiEnu6zi40Nh2Al75733yWY55iCym7iSkaPboG
KxteTpBEkebV8tpFMcsoC0vDOJ74poqGGaqzCC8mfQsM/35oi+EQIl0Eea5aG0rFTGC4N4CxiG9D
wZoftYfTUDBsO1s8W4QpP2IutnGSgl1qRgZyNn95kVnbSliTi3LGvj5nwkUYlKgOvP/r13waiQsd
3juI2YzVTDFtwDcny2W+DEtxiW+Oq3F7i+gT5zcq8ec3g8/37yCNFZrOjlq7APbtSVICKnEAHQn0
CZCPm3RLHEIs8mdRmRHWZKUrs1fuCKf/uNva0CxgoCoNEnhsrevlbLki6U45EcSrSd8uVyGAVGs7
363gy6Vv/42QOSjlkTlp1Y3T1Zqtbhv8o54/hDw3Jt8PXKmzV5xuOkznwTVSY+yRjVY/QwaRayrx
XGE4deT6YiqezI4NtlIOkMJn0fV9SsNl2O77fdPdLkZyBzktPRnfz/C90EWUlZc7RU6CcB3mOEbZ
uPx0RDBGsAb0RHk7uuClC53bhXWV0SNGQ4j4rCvi15iJlfx5W3+a46Iu7FJhIgK3z3ddPzVg/H73
JD/Uwkl1tGD738f4Z1ez3NLXYd9+0rMOLlpxykVYmXQCoXMBSMVfqt3J1d1V5M0r8CV932/tPSFJ
NQ/u74ezht8dtKadeY4vNjudWldzDne4FgNi90YO5+875yHtaYHZdoOKCEU6aaira70FHrn4dnah
VJNFmBQTL57g58YTvOLCd//mmGn5L7KOdtGBNbDuQgp2eJQh1VuRBwRxuRbrbV+tDXB2ViAS57bY
edafPzOkVDxNPymrXCju+yihrcJF0APGSCFuKr0Uyl5ldRRA4YIdwa0R9bylYRwum/kk1Bq7v2GZ
sv8uu2TE5AWl82IwNJGYFQkNrRGe7XrR6U4dF+XfuQrubwWOt5kUxIElHb6v3SZIP0qJkNcz4oFj
bTHptdCO0gs/f/RdC22FTqftglnD92RBKwXSZQShifpprxj4E8YwoyXNlDA4th5BcpK1TwmZVVbB
upyc47rBTzIjOndx9gcvr37MVmIBUiG72wIcUI/wYNcmgYmxgaF0Or3BNH8ydPHB/m28CW+SjwFp
wSHV8e+MsPhC751z2vtgdSPBH2enS10AqRRZDgjlVDyf9elYfbq8IVs2JBNjpgBCJBHtQsMYmC1C
iFrMAa22aDIX//f13x2osLl4S8EFFN3mTH9/kekcOR39V6r7aNgPw7DnDafnDro1lHp3ELCN+4oC
TG8w15YnB8HU4WxfORAqkCqssmBJHANhoAgpe26ogj4EK/UPKGqn/GNr8Gff3C1+DFzALxwktghH
FJMbETTUfCj5aW5DCCyD33gXcN4FnqM5FJRgiklSYvi82hY7gL0AtMc3dUSjYS2n+mtY39GRCJ5G
OO3Hm2AMSAIMw7nWdpsrsfcRb0baYPrViSIJkqLYJNF826rWrTUp1AUIJ1OEHMDIy0okP5UIRcSD
wcyjMoRutBW5WiRX6khSB1DsnhX8Jd7Er7PFgENu6iE/PFFgWkDmPisEYVybEUYqNsBzojgnxl/W
r1NOaXar5ihfGRWohwRLXPMh9v15J6eaXfeeUU4GNnygqHQJQqD4KKVrNpre7ztJVToxn4Xhnl3r
mTE/ksfomAYbKAAjfzmhKQ+0YA08IRxG9WhXXblTBgRlckVweNxhG+/8RlJCg7ob9dTExtsGIUsp
bjbWFUMvFeSIIfB/u/ieRQMw3ZoK04RVkkqNwRMVOZaV83M14MfJ5Dwc9dRWxrWICKcdnJ/8x9g1
Pz66WIkAdJSUdJD66aqJUx0OUsguHbi8Z05eg+EAg6fkPvwVs273MvHVoGpf/ck46YKQr1cyc/mO
ZS38yiw46FeWJK4A6FWKmN+DRcdGLVyCKYgOJCDUVJ6UEmi92MVKhjYhHLKn6xjNZE1dlejdl7FF
bLfSNTGj/dC7QzYtswYgfh1XcpvMgOKu/RXh2lQah/Dp40Qs8TBVm2oLESk1CKg5u3Lmwmqa6Zor
uihpSBallX5uBzm+LWbCqOx5U+36pN720lPA1Czqm88uvC/DDTnZ/H5KJEMBIGdI8NZy428ImXcR
108gFzfTkT2HitHn70sv09pzowRqgnDz/E84nQatKN2KBWA83yBUXJbkoYBPF20837z6e0gW0H5l
UF1fiEYVoUU3bkN/lMpMm066S7KZlmHkfP1x0s4k37ukUGUXz1C8vmk1wBidjdKsuyTcfRekQy8T
nI+CP83371K20zXFJsySNob/XJKW1qn4ZDKFNRBPMbvhHT39Dsxoq2okueRK6j22Jkn7+Gb6D9HA
7l5kESdnZmkZ9QO5oLB5Lk9qm6iMh6l5Yj/0PUpE5EK7huidDM3kFh3GpwpSq3NhfRoftGSR86Qi
w4ZNBO1b/hzxC6LJQvr+nsrUfNCwCSuYaI7niqLKwoq4opSgKX+WZl6718oN4gTKGrg/eZ3dKj67
dLLQryB6CRjCjO0fJzupkI6nVOZPUSTn9zgrccj5T0TpuO7P8UH7DN7kjY4tblEjIEoRPFjptB1h
o/ZaGYpo4FIMuZboD5V+xxaO4wwQolWwk/i3razhsHYfTDVRbSgnuSNSed26kh8EAh+rb9Pxm2bf
2O0ZPa28KHCOHeqMJnOQ307lrQesrM0vnbV9oW1nzIOpR6t05YjRWuGxWUQLw52+ezqNgh1fR3+E
yhFVZb8meTwyulrhfFqgY4T1x4h6mbVsqCLBoFDyakq44derGrbqY8/T/OZcSwsG3atF6k5zsS0w
PkhMWNLt1fR+qZMlRXaOI2TnEvDpifPZb7CwB5JlA2AzM1gfdVrxAuigKFmF+4Qbt9N+s5K30elA
8rL61UgQNeg5s6S/hliBiQpqQDHkyhXjyn6UcxMtt50wtsKP6K3/62+geEuLrmyMD4P5G1Iu2Hv+
hG0+gBxCuI6EnT1kYpk2XeWGh/niW9eMGPuHIBxEnuPqpIj8Vc/kCwTDeIdVO/qcCXIFFGrtZcGo
CjUfNsoM+/NOidP8baaQTCHzfvVR+S33F9VGuRykB5f/v9aXIegI87725cA9Vf2b/OAYwxAFSKTR
cXJ1cG0CDSoXL95H3BYdcxIUwB7cUDzb5LbRxtiTey3AhFFlBfo9Fs9iX8zpd0p8uijohkBlyT88
m1eTibCMzmMcgygXIYglAB1dDZ5m/Dq2wncCfvEn80OaVR+bay3hQ00ZQgAlOy6/+tFdHZWsti0n
efwgdhkjxy16AYsusVrnUHDZ9tbrXlUgCAa3d12D9zUoXMlIk2agMmFh7ww/mmt7uCu4PpHrVPRS
yR6hbTuZ5OrBLFAYqVLAufXUbuM22CvagpjiOfFQ6O89eu4Y1kk/Qs5nOsvJ4f334PXnFcK7GOxm
Ssb0m80/UA/mjd0uYpu6RPrGWOge3hINSlcsASJU01+XJ0rjNHReRw+FZtElQORz6zrzENDAORW2
pRVsvUHG1cs00RTF2C/zSdL54UKvFJ+bhqsn6BxFU1PL1gdkuS9H9m9JUQJCosHcLaMjic9GNttO
FD7QzvjtJQKwmLv2rhLaNZn6V2/MK6Ogy/FenX5ztj7eEaDgKg5DCuEXjvb8kn8h2xel8aKgVBYP
BB2ieSSnTwPbeSJ3mmveXY7GZteSC7IzwacPSs1KORrp5ZkII+jhdy6ojcTA23DLkPS9kTAi0fZt
JR4rwpp/hidW+17zIYjhntfbQd36lQM+ExM9/H0hHAzimjoGhzRzqC4ZFYbYiykvPV4d0d+O+zt9
IrgsyACjtKu1sT4+7vUirjxZZq90jfGNVgeZzny4GJ0TkwO5hkHAQxo2UZOqQd0KK4rKMdo4iOxm
f8EoKkYo6ZyB/cbSVFlfiSBMK7OlDMQ2Puw+q2XvYeMIJPllg+XJI8W0fka09hIrZ2YvMpPUOEEB
O2Msnxb5wSYjsdtLp2T0viCXWvyNy+XCxT+OX8ArXfIB9165YwrsSj1ZerBXxxFa2/W4qKUn6I5C
6T0LA9hQq6bBYVLaMc9+FDKJEJWtPYqJXq9MnhBkIAl+dkdO2o++tpQJiGCyZ95jQMHbv8EBlDTH
XVjLLVq8bwbcvIaegZdLdF2y0fQpaEt6b91uj1w6vhk69Oaakb6PEu3oPov+otFykh8HILVNfPk/
qi1VUxuyq0zZT/wX4+t0XrrIiva+rUGx+TfrlKpJeZ6GyKDKCa3Gujol4oWzgNamwEaRRZaXO7pf
ZHvxNxowtXwdIbfc2JhvkQm7/sTHY+IOzMaIb9EpsLr95RDBvGdJZ7YV/mK+WtpJ62+1l+HvQhq7
+phKy6GY0nzkqaSvb2MW9r9+fWMLxPJdA3nDFUzyBZpnPpfDVaqXmuv00R7CfUZhZoOvWkFZoMVF
s2vw9vcjQEiijMrOrCwebV5/hBxjnjAs+rX8LBqZq6+Y4PGZmycp6G/qeiJfo0c/n9UNnl9vyx1s
KN0GzuHs2kAieCZ6YIMulZr6eJ178wsa3+olMdBPX26qjPVDqUmd67zimb2rA0TMGt0zWxEWR5Zz
XQugdYm8/nGsakCmEbNLzYpyo2wBDZvBTGlJCNsZADJfbJbHreY0BcTpHyYuUKXL5UNu9BywTQWc
KxDwdBTqtKvVKUk+euqEJImep/uOXK79HSUt4wsVnerwG+37ZdI0vNY8u2E4vFDUmpY1QVSVRazo
VvnGAsWu3NA8y2bk4vaBIfitbmzHzh5KNn8p0az0ARqqz49aF3DyM9NBMv/644bSToDdMFVlU2dg
creEmICAVO/4zbQ7slUawgIlS1ScuwNyzINlC7kLo24WTpiIPYRFM01FA2sDAPSOTh3Fv/GaxbXe
Z0SaNi7j05ee9Sbu/1zJAjnNBb/Qtw8TpDMaxx0g3fK4HDSwBIXtqLHxbczEnpz0JNUw7FEUoScn
Nx5doAFF/Vw1F7rWLW8gbGuiHYr8GG4gLcoIU+nVjzah8644gV8NwEihfOpewCopTUXg5OAnnojT
Qjtv20xzIiFCvBkiz0Kh5Dmw6kOPJ147fq3sBmvQtlMRBs2bjCrdU9QuxhXU+u2ojd4PMKGmQvqj
4YuGX/kLFXvbDSJpxepdj8vORxvtyeeG5SE9M6XLMLVR6dsBmU25Z3ZxLRoWSuZEv+VfiiTuJtah
vNCY2/uCGxDdWZ2AabpVj2qd1lFo09+jE3HTPk5M7+ZBlyrRIT+wsmQsGktLFpQT7TZgxlgdZ/q6
YcA8WeFXMNK+RdQAc3nzyNIjJVUJw3urzgETjC3vubhdrQFTzLMOjQII6Oa3WsOMSQW/6DpieJ5x
mf6v0u6r3qMS9YuH7cPA0G/fJ76YTaPg5js//VATFfAzd4xCxgGsvvqfvTeLfvMeiEfFIZTSrWpw
TQ84O+Z+09cr1OYLa2xHnprjFe65yD/mhW4fS68S9FMDTWlriMJOkPmWhd4EZbA320nuSmhN3zsP
UnEswJgkeWLhDbSKtPPX9PZlf/EAxvRbbjjDdlwEUi1qlsnH/N+rFqt9epJbamZ0qLDQKa1j6cYV
KjI7RWe8Icvjse1bRBSy/FojhxpupdU6ZfYbjQEYDX79oQdeN6waesQurEiHw9eXWKNcQ9zIo3Cz
rpnXjsuU0YI2wVfidcO/wfgfmvkrUgx5HsXSXCfgS4R20l7XpJeTN7Owjsext5I2JvtXbdPHbCYE
eJfFMSqnR+nGD3vUvkV9skD5QXeQvZ16Ut4Qzi0gBrcyXA4gHZxXAshSAO0qVgNJN56qlwDaOODe
gzgwK0I+zsVGaKlMCSpF9MC7CvJIbRSOP9v5KWsgx79ZZbXaWccynKrA8s78Uc2pIUT4cEv9MPqV
rgAKewYyALnhn49dijufLzKZi5cloCJDcUWi5EElek6tNY2grMs/984QT9/iCFIV3wfMtAhz4Ktj
jtIlF805Wfe6ET3KRiYX+cdwtM50QfADKzib3tgapX6WHRXuEeUof5jf355QrQkD+ILAe7qhgjTF
fF0BnFPPKbwAlegwTyRDWqbDBkBMn1ulCPOuyPAO84VW4xqRF8NXceZx3H+vryZ5jn1xvErZTyzD
VTi9pq3uk+i3Yl07CVQldPWtfU/GoVPNJqA+KwWXLVhXL75ji2lyCCA5Rz9Ka2YiqK1KYEFTgAkS
CI9fDmQWisyjXTT3DTDKRSlBSYd1Bm3frQl60R2R3ceStaRmhiLIqce67ua1g+mVZ39OPV+jdnvr
ReR2Fk63akjHzPk3p5S85UnFJMRWN5jN7CBPvk8r1jbJTAt3DB5t102UqhXTo2l2BubWukfCRVLW
TlJhQAgW+dZ+xYQG/pQ3XOS1JkFWqlhkORNhLb9ZINsa2+9w/vj+dDqof14j/M7qsqiA5RaBJxiP
xp3sQrBR5CP3ugmcTF+N/6pfmi23WlRLitSRkGxj6c8e0QrjSvu1MuJROZvGIKTRwJuX5c+2xhZs
3HbGG50jTKXvr902raKvMelHwWSwTeL9u6roz/J1Lfb/dvbRKFU0PU4SiXz2A2AGw03QC/x/I/wM
hKMs51s4sUamNlc/E2/rxLbTq4rZ3UQdUp7eIiwBWv4Bx5sD2pCIdDKc5tk4FTSdNv7q1tILyKkB
iF8+3cKq+/hDKyqGaLbH7p8UFxcibjX8N/Q7X2SeT2tO0EUIexM65gJZYu5wutOODD11cuRc7ppM
E2KGHhCy8MMxrc+AFdg6UJaPy+C0ldfvMsLM7G3MRszVKk9vHsKmMecyeg7gchhJNQfJfCSWwx7N
NIEHuJfcjblLRRFBULR/NE8XG59DhNsURDGqFCovJ76P7MR68lVzYKZyxpgoZFqUWSr0HHA1fzfk
9TDms6P9n+BQImgLTPD57ibqoU/f3zz4loqt7VI4PhGZ5ltSisLeNnqd7omKDMSWcilVXHzBYr1C
QhqJdNM9AUGvxOESrY7OwZodVoOFpZxMrW32QWvpL/pbAYLbaySBSVvhV3TK2FYD5c4JAsEl5umP
qjUbLcgRVroYq+7HqvCoOvYdLpYGRpItx9SHa1p34rQoBJBY56ptLokMfw1fS9Lv7V3l739YKNK7
2Rq5VVr9JRZWNi/tBlfjjJYmoXwjECOH47t5b1sm5x9e26xoed+i2mW5sP56l46jXhetXVxVt9D8
b+ssUzZRP0eoluDQlpxiqQ+0luMe4CpRPeP30I4E+VHGqN1Bbd7x4C7zPTx6qFkjS/AaADBJlqUF
6pl+Ic9Aqz6c9qfdOMB5sm1IwGAxKrQ3KeouAAAaIxJk7V+PYUDyy3mGlpbtaxybSY3AgS1FXYZU
9ew23hDwPSwyJLf4l7/ZVBnoyMr3BbKhahEUnpWYTK9OX9MVJmAH/YHc6fR9JKwTWNojeLXvXYtj
Nn6teyC1Dwi4kBQh2AHnAj5L6bJ3S7O2gljZ0aZnOReFP492rJwY4UGl+wqJces+IQZqafuC/L2V
mlLwm7Zj7MNg458ZaXJtaMBXJRVdjdvPKyK3uDkyKLfhhvE3m8h+xykeCLehbizoCl0wX67UNH20
14XIX8TsyYiPa9n3/3gKjxcBcFUqfgIp4WSTE+RevA1WqgNOVVyni5EFQDN775LlPNjPMMk8qrJM
LSkcdHiL7IOZsX9IEvoiiEz3lpZbpXIH00lKsP4OG2oY9Tp6kC2lHnKMxSfpH18VH5Gol/64fBOh
slbAjq9dUp1FIQvsFNvQ3Y8kB4vI+L5b/khUFyFXZpvcncaUQF0wpUj6U9uiM+KCigCHqd7pmzID
/U1l35m51vtUEdoiUIx1RPx+R/jBNPBb0HumkKRfncwcKpcAP2vjSImg/AScvEJDl82sbttfe2sK
y8q6FEa/yInofVznJnbpe5KQYtPSrxIoBsfVGSKtVNz860vSuLml8R4i0Sp/vPYmavCA91IXzG05
NpV0V4tdym2bMTZKMqplrS4+fOsvrNGTIKBnAiPqi5dqBvwGmDAiAvubSdpeTkIBxhIu2AF4NyY9
x3XpVFec+4l6ts2nLRNSWtPBWbeJbYqWljTryqFv6EwGAheHEZHiHRqfVS2turoBawjk90WrJD7a
aZmFPIeQUvddzTSxAnbVrUkmtpGmhGTjgngupxPy+k8Qlh2n3Xdd0Zh+Zry0tpP6C1sQPBk3jNvT
dtJwsfBH1ZmCa7LolNs0YtcarApUhhPEmNVUu3vwhZMGmVpAuK/9f024N1oMC53GfZbCzaoMBbBS
wowh5Vw4fkURMT6nPg4RSR5wJmGsBCGV7J6i2LCSy1eJnKI6j2M5tCH2uXZg9TVBZeBdP+OnZWia
iDN6DOX/xFGDtcHxI1Qc0viiUbo6UZ1GUn4fJh8LdScI4loUmL7ck/ARgScuV9N2Asi/Fcmk0CGs
bNWkV0T1t0jOAQtZn/5Pr6H5poaLTWk/A9OY81qIpDPfwlp2WqFG1pOU2WL1nsbJrxqgojlo/d+C
GYB8cNL40LMMJzufOdKJ2st70sBYICmycasFTfXtrNzcoNUINoTfeq316oHy+7dJVAuQvabrv6Qm
WquctIpfCMWvgA1ABt0d8LmuzY7t13dFEoUVdEVULGIbdTFn4o94D2VOQYbLGa2dwM/zjCokv6J0
+PGvGY2qMxbmAwSFoeMeWLRgfE1c2zucboSC57evaYEpTd+5Kf0fMlnozJdI0Ga7BXg8ouoVm2dr
56QhAgY1I3vqslViP5LguVFPcXc7O1MT4GLwTR7jokoDZu5pBsRFrc2DsxksBcYsTBugXWyQFqQu
Udtmg8RI4bwIVgoElFwR8soJZkVOgUoYmCcWloAdsqGsD6p+pcfCxRm9/hEtohKItDhe6PDRrQRl
aFvyK2AZGg8EKMqDoewXBkY479oIiYXYZ1FPJ/ojdhRAcEVMmpkUt6TmOcakjpWq0XJ1ODdglQjn
icOo+EdXpNV1iw+fNSIZVT7VrYHzaPTNWJfWD7PcssADnTzzU2lIT6SJ2xGUqs5oFHemxdP9Lscv
QYPduAFlnoHB74W19sK/52+Fie4mCeW3EANI2gtrAQHVV2083mLSK/6R13WeUabnYE/U8XBVqRt+
tmG6ubWc6k6Ps13gKKRlQTuvZWc7EJMA3XvJG9cHx41eeDkSVo1Y+z6aI4mikKq8Y+xoOW1vYHFo
umwjM5p2kT9sSiNfO/PdJFQTF7uPsGl0XAPrCtAWHasRiV/6Mt0Rd2an51iT9LgwcuLcBa63P0UH
RjF1kr6SIf6hBZgNBgf1cEOpqHzdn3StWk0Puu913z1i2SD74vP6I9K6TyEzKXMGDetWwZ717RUL
ibSDiq/BY8zQc1xkyu3frLhdvfvUzN1/+Sq37iQqYzbWTQ+PT/UzZD2avaerHArdH9IA9409PY4T
5y6zlScnXs64tOkb9LLWQS3QXFCC75nNBZifAVdZbFLyMVzUJIRhaoKE2EVRZXuZRpjOUjEsQIBM
kdhmLoz1ztahQ2O3EgE2IdhCscFIyo5QwCJwHKOyTYb1eLBeqgGKerV+5+zBSg3s/MW50Hvtz/79
HbJDgp2OQblditGxfQroJdf4YZDY1Vru7H/4/y+W461rky87fNb3DXYBrinEC8IofexoRoGwuVkf
L5CGsP94U3suNjs0yNL6hKgvuWmJALa92+SIdpuFV7HBjQMuLPwDUKZuXFVseU6hCtI3yy2LiqWF
quxu5D57ISXP+DW2fIcm9O7d5frRb7zqkEgdEU68rJ5Io+GfmoYBRqXtD/yVBAHokwEQL+YMyFJY
meWm8jTpg5/3P2ZGx1So9fUxMere1aP5AUEp1O8SQ2+Sy6d5m/rP2htvDYpr0cRNjPB6W86wyUBp
hjCk4H+bI5XWYBXg1y3u5sm5NAVmXfKm+1WOfzUrPAIKrK9GUQx03vtTdDFh5Ag4kcxsXkbI1dqC
QjONOKJSvH8RnExrLHQb0tIhDYBQJidvjOHQZBAaUW5yZQzKIkTYQr4WZIbRvkG7NIZiQ0MmuBwb
zr01nj6Qh0mOtSprn8raKLS6o1hTrmu8DRPveJNJ0xulZy5EtyD+Fmu56iqmY2B9ZskskxN1tmAz
AZFsEYIxtQlqKSLLqwnUoPI2p30vunaPDEF2wjICuRFj1wXN+KWcEWi1NLT2an9gnc2IfwZajS4X
pVbR7BsEBgIeETmHxfIbAGmc/02Zd+pyWBlYmb3+T/zrdp3LBa8maRDimLIhAp/r4E0PpvuhrC0b
P3AWPtwg701aCW4gBSXgtLdhh9JDzxbyx+RiEzKcNaJH4o9hhDte+sXFSD4tmH8quCdDiFb5tIwK
ibUID+qRIAOm+5zADCxqEPxWQdWOPh0lTaRbongLMaFB4fF4molC1QXE1XhP8ABmvwRZyVT6yJUF
vxDgRTl0SfXq6CuAeUhjP+EjcGLB0+am4ah/Rk9c0Quiy8U3MQjKh/ZQ51Bh13H8/JWVIVVwwIGA
lPWW+dVDNV/cXWMBZucrCDkAKHBNxeS59x8MM1/tTnkEBZcQexeZn7Sz3mCTV/UFIIRLyylcmI2M
jwXZXQr5/lCzi0Pbb7ODvfxXJhBkkbimp3qvYm+9hOE46g1OtBn5rBl4/DR7u12kXDD+QW/3vvqE
6v0UlHnE9EmE5vjpLktaD0US+hP2SOh+ClbL39bE/nb7881XRGAgcol1xuXS382VoT9AvUUgWJuu
UAXHJE8AuNpdhsEtGB5W13J6g8Qo8qS23i7HxfN5uVze5CcrnhQ3QB0J8oG1wIhb4nepU+pclcO2
wZ72UtvW7EAFBhqFs0UHbwfCtqfsyuzwWYsitKAILtNmoWMNzM7MQ6gVHoWTnbM5w0FNrBtymUiJ
zsuaLinOVu3siDcG0XEHhCxhTYzCgjT05WuicrCZC6WwwRBTuRkVdnEnIwma7szcanJp9PqW0bgK
XYNU+bbuT4O7oXi1JSB1JjWIUk74r26kqaVLNuNdUUazQcNGSqc/JS4S5aIQAuRN1iDq7kaozztf
2+JOrPILQGIylMuiiTjqoAiDTfiStUi6g5z+T1/UMdEYvQSsQ7A98hsN9i+RNxVZTJAaL3GuqHlj
GTEH55/eFcNvUez4i0pdAh40l/7sJhTyXWtzOmRzkDEjthcqxkcla5QAtjMlC8OxbhCqODyZ13Xq
u62Fltt7SssHXGm4PvXRUgnN69GvDu+aGNUT04+BFNdsGk7Mfll4PL98ngGSUe+iG4SZhls8PGh3
hi6H7A+GJxfSCEUoaSq/Acxti4maIOtnpkP1fhsq0qnEgv4fKbJAEL5+m4GE6vqa3ZbZPCpcDUKb
PBWJg31ymej6h+o+YvXDGe+yO3KZsxG+ibFTlWNDxa4tMdrWalAV/nW3QzAXrM8l5NgytXWJw0j2
gDXgOCrxyouT44MYKUOOvnbRclZbf8L+uFtr8uctSfHU1Y80vbhfLJozRrSjwcjaB37/ggHDsypP
Y4vVXnk+8Xbb/8yWUwhc3OQ9JjkNqCCCcxIeQsmVd8g3TnjqFKcUqxV7Nm6TjX7cNB3/4tky/HMS
lDTz5OisIsy+ZXEzVn9tsQkBNhrVXAXvlkoNyRFwWiA/x99ZbP1GotM69SeTDbqHp/7joaF32gnV
jxPTWrjGc33iIgoE+hJx2+KCy7bMm4ooEQK+I7Y0VuCLYa6I2SFKi2DHXVD31sc0ArY88t3WM4XD
LEC1eI5Fs5Ev33fsHkGL2s/ZVS2OUTT0I2ghbSD3x+C0+Ewl5UT+t2uyR0UiMCvLMrqljcZQRaYJ
KX3SFXH1y7GuXXoK5aByUi7LXAfG7X/f7+fadmG6dtSIKpSaFYBI9uQlYJtywbwpKmMeITaqMY8B
6G1modFop+CVs9tnrkK2kumfozrWDJUWs7sZC69CY/mpwenC0yb6YduHlXch8CrsuV+0bS1ah1s9
qgHenIEgKpn1sWm8tQjvGxb2FIVbKrbwlBI3SAuVbHz34GBYwgShig1GJyPkNfH+1AWxo6PgaslD
PN09bZ++C09WsxLJ54JY00kiM6NkPStI3x7gqi5fsvH1YTKMYoSHc+oUOHsq71DaMIPQgCiSQwGH
j3zwKX1oNO6lqxMOSMoZmbFpo5/nQhF1CJnhUEd4xT1t7E9Ss4CgoFXs+0onaLq0SGHlevjBXUJn
tDPLc5DWkV6qC3wtH7V1qKR1iC68hRB3VrJwTWrUELNKXBxzF47x6eCbkRIGg3LNzYNomoTDEuWf
UE5tsd0/ii0VjiRargcksmvnXmQglMzli2gChGconJIRajoFa+Jxam5zyqj3bQYPX/2U0xmNEYQx
ru+XKFS8K2oWpfmfUOdFGkokE24awP9SBlJKckD8Pc/sexY1NvhbEvjqLsKN+rk4vcvtr+BM0Aua
FmzjKe2Rrf7SDN8vSgIYwEw1j7a3odZYL6o4RjUdZSTmvgVmjKYCURsphroJStWl9U951E4MMe1p
VgxyPoUXYr7ql1Ot43vgTkq+SKSeRx+OvPLIfLmamM+BSIBkDXLB7BBJVeuy2VoVNLjICEsWiK8z
g+LteQPrgRS/V4C7ficSpZnMrIwPXGIRx1UlKZk7ZsWtzWpiXg3JGTUE1+aZDMk2A0VFCKKBR0N3
eP0IZBIoi8mWv095fNzOHU09GN1doh10q4j7mBvqqRBmMacG8Lz+61OzRIBcmqM3F/j28NK/qqYX
ww0OdK2x/S5hmKP3FomBrtOvprVvHbCdKUyj0wZZh+W16pIW+1f0rLDxo1+x1/wvrIMmfUdq4x2k
ir6y/0Dq95EXnnDWoSMvTwvUwY/eBQ2ktulAharNph7LxYlZs0I13KSWxlmpnFPX48hkR+gqWdo9
wlFAUawerjA7fVv8WiJUpCou4gTLTVxvoyly7diFpx686wTPyODq87wJIQY0YOz3MEJswvg7rlKE
Rf69/ngpCIc+srlUu/k67UgX0yEUMfm+1gtUABR2Fo6grL+FugWO9njmHyrm6SVpG85s9aqg2Vp9
q6ShnYFd3Rv8/56Hq8aqhzGHDyaHtxJs55MUf9ir8n9hjVtHtLTZL7aQaFrY5gFSQIlWpohPVaAm
zkOBUOUphRdYvSUX1k+3hlJSoJOgLC/O8Sm8dbwhEE3t7cwL78Z8SNbpNTFo6GNTh9ER5R4MXy16
umUyxBeOAvCHk9E5ftzCbCShYeHb7mcJtiIIn3UpaBiyjUuqGh/MWIQXfpxhoQuhJai/JVEMI/bG
7a2XH69RL5X8/wQ8ppbY51Qx9XzmZt4dDYKwwMNnLNd2qm2Ie3XQaeYjqJ4B2hQMt9c90dFw1Wg9
eJ3YGgy68h/lsJel9fcYkkl+avK11KnJF/P15F+sxwnqY7tiOBoq6Hhrqdu5S1GIlBV2tafUJD9v
CvW/6YNGWKMzzYyeAPBG1YbEji1nSjMucbZ0IVqXfSSSniCu+R+0O7OBfr3US6EasvQi1N31pJkp
gFBjEcQaR5NKAI9uXR0ZqGRC1sZTn97u8a1HtXGLBUm4VYPQsG2miroe+EsygSXF4dguun/4knTd
E6wH1rn1OgbXSeEA2yQ7YRqoxRKtFGKADvy3uhMEertLQfXZ9L0cP7X7WHINQUa3v9EBkioM5Os5
kWk8lLPyKEMOzC5lkW+44ozVja/CzRw7ZVWCgf88UVpwOn6AaQS10az63xZaCarx8HT5KTcMXjDE
uWDq/3OYeY4qtgpLpFu5BixpN61+zW/ge+fDrIpL8iHx/MyrsuHV8C8RbDiIa9AxarY2YI/FqBsO
wvty4/G9s0o999gy6cC6oLsLr58HT5qv9J/65dJ5Vk9AaQI76OTYhq3cp3rtlg+O3tRf++1i4a7a
Ko829qS7zq8bKg2wYrraYM6ak551ueeNey03/CoMktqAiPSgUekNBtGOnmRITi+k22LZF1ViRguK
KgHBpPTqCui72ccxa2sg2aVMilKs2CvbIEKmrgl/MvVTSpD7LRwQ1nGjxJbJLO4JT3FOqPZRnZic
3Mtt7ZEYLiwF54af8klC+3CZT2m4iJ6ulIHrSzDfMgT+6Upa5rMq0JG3zUnmmkq4xu08rzteayCX
TooVpfKvluTqHbw6RovWorX3z4GAFPUehPhsTcBYU2F87Uoknazn0hagJ5TxSDOeTlYNt+CHWiWG
481ZicEB5KuLpYByBcVUTeqJNKYYU5uPi7TtvEUrxGrA7PV796Ywr4Kk94pDWz4QgyB1fCICjU0B
s19mAPBNs4IMeNtTe9+iBLFtd1ptELQ1H3Kp/CVVm79ME03MPIAcWQsE6uC1/sChi3/4iei5lyJM
prI/q95u7mzDoPWyJAuRIW0AWkhgL+I9TW78wthNXHiT3SyB/BiEwCdYpcM6rIpjre5FrLjZRKti
R11AEEDn/cdTCM8oJCG4GJZIh2tADZENEk/xZ17jkUYikXemDgxWHqRLZv8/7zhDUbTkFqtrKaDW
mEehnNlOAyiikc1gpzYaHrSvkqj5v9xRWLflY1E2V+e2LaV/R2IUAT7HwkhTPlbf3JIjAWkvzFkT
Wh8UVJb2zgMelECCT3HpLPyv0CZl8SN2LG6N9LgGVrZmHE7YGlGaaGFoXASmLUkOZU/mYSgZDQKS
faCARlWLKNql2BBzU1X3dIsE5bYJadB0PG1iTTIK4ifvEUv9McmIB4jXZwZkdOHEQ3/jMeH8xHCV
nwPjdR3QAKgPOCo1T2WXDIAZdT9OvJ+X3JPyaXEskzb7kKPRJHG8zbfLXQ1IWwTSG6QmRQelkaI8
ZLbtyEgrHri2BwzlGFNLCEop5j47LL7CBvLKbeuIWOUQ0rj8Sp6jterTGNCwK+w2l8LvHGMBc3Qd
TARLKVxrSjtHDO05KBUIYin9bWaupkdGLwrENtcqyZ3vbs4MG7JaDwOZ0Y8iHXU7fWdojhcmlb82
jnVvJ31qcEFWCzXoAFZri1+2Na2lhJ1pCEY/lDTV9j9n3zGlXW8tU58vHG95F3nMT6igsfAwh1uC
Hz+v6C0e7RE78cmxGzdJKTcR0Ug3QpJUXl60W3debCkpssQlENWBrplRdmcK8csmhk1jhr1cH/Y8
vci5pwyfuQ/fE3bnxnHrosznQROyiztZPg8B2CDU47m/Dn7KoE9Z4wXeAymhQtZ5ygY7+1IGs309
Bn7F1D5OYIkce4UQ6ctlex9s/6LpUGQ5x5tcOEUjNrHIcVkKWbkVazYAxF6x78AwNfDyce9UaGNg
ufcs3W1diikkkYauS3JBaPF13a5dmVVn8uuWeBj+g1LROm9X/Um/Jo2UWPotvqj2HqYGyXvGMwLR
b3QcNve54KBwqZx1OtGJoTnsCelZqEo3g6hC5Bvybpf7gEAfc0UHzS3hARkFl7UlZ0eUHGGr32fg
YNml3UHdZVzbIAmoEo7wIPBAaqoMu7SNX52DwMlwA5HTOHvrTGUVblIG3yIymTT5kTkhN0kqWLOX
Y5z4JPTGjJLsVp1VtfAzmiyD+LScwzWxhTsPoCw+cRN3UUZFzsS+qCYT4S3V4dJeun3EMRnrnUD/
xGvANrKUN3lbwSlpM0Cs/9WQHayt2J4UOt9e2zIYzyNK+xUT9Qlz9OH7OpSGiqNLRjf+xZRE7sxT
DEL/bKCNJWZG2/r0gCvYiZ6bbHXJakVfA1Dgak8BuHQACfKtm39/M6hXFZRn/LznrRIKjd3M0BDm
P/p8nXrWNxwqvpbdzSIztPuspbEVUsp54GcP5LYPeN5IvoVvwqXzXKAxadIMNsV8qDBdTS6hgn3e
L1x0M3TCanxdnfNBAQpIpWsTp0qCQCPxNjCMMuUlQLr/C3cjgXyPLBbUF+Jcn/QDLWvRquIN7f/j
fIdEAwF/wnOwBDf4CWZcePayJrlyWnEKOeL6CQ++fk1EWRkF44RjeLLsvyb4TdbbKIUqlboPuoGm
uhwjiStQU14KrCM8IBmSKArqGnu7s+qWy+0PFt6DuE4vhW+oEbFgrtQiFNRzQvTU4lfd2LAkuMdy
UgZc3XZe7S/n7nH8T5OTQMyuzo2Ra/M9EXtpBUI7829mnCf1f0rTFmdzWIyvZW1HOlt6QWT6aa/Q
8wVGe0kvawiigBUSsjfzgOnZL/k2k5XhbPT16nLqjGF/bLYQZDvyErROEhVc0Q/BZVaC3PgGOUYP
ViBaC/RUxnSAJA5r8x4j7EMCM7qjLJpQlGUcjfByV2WUa0GGmYMDOvXlItPrG2/CiA4rrCdoPbPv
cYXww1oPRSOnPF59kAulBJX4FWKxZFKOjb8oI1Bk1Setj36DZFQCBGdnuHJgDZYo5SbTkbQwRJVm
sFHnIoNQ60L57yf3wYKBmsxx0edfKSfcIkRX9AN+mRG6VdA2YrS9bBuhOf1GK+sq7pLDP412wkbh
OsSy+m0XigJKs0+Vht33m6a2vcji1ioW+Zl0ZDEm/Tv7WiJrPs2vagqXp6BSoFfrjDsx6BQg/lVk
QIEOOiY1RJu/mDrGbLSUdbmVZPJdiHCfIhe4DcS9ExKnRk1JVLlJUObdeQ4jAdU8xaO0qWwSEThT
4/T7fm/0xuaBGcdVafd/iHcO/FduCFV7OVVKGrPcS9sXiSH7ySjJ8w58m+yRNAb9plQou7hbUgCw
hkx9KY86mDD9nZwoKmdhwm8mib+3cnHJDVPz+i/A9bMBS4LcCdc6ProqPIxd/1d/dKnxTnqicGXl
/K23pj8B+GTfHnwmRN0mJxhymf/qKy8akAOxWuqofyGGjktrOguA2s/QQBmtce0WemY0lZw3kMKd
XOqvYknbLPesdKIZkArFxkxkpeoIjjlV0UnxhumIv2Jmtv6T2twoPtacso4KoOfOPF+HnmEkXAkh
ZMj6GUq/bEKDJpdsLLInXrNQtpnY46iEP/Jtaz7H3VwWvPuNpXm5G3XTWyao8J1H4td0WIu7eh4I
xzEUJggMvJLndwG1bYcREl3JSNN0woOqxrZsIM0XKfOeCs98Cakt0YKsslMBkD2FpnKH1vuR9dXX
U3/JfWeXJ9YsAgpoAWhm9ODxnqUGBdtbzdkjLUyxTr1eAyb0oJ2mlXajX6URT2Jy1zMnjTkWLLjS
8n+iDfM0E05kARiO9Lu9W6RForDwHSGyLp8cAgFjZtJ09Lsl+lpju/WBb2PDawOttwbOAxtkznT2
DAzDeE3VAjkju+z3Wbxy1cO8MszRHSZmyGk03hpla4p+H2oWEvyEhivLeTna75gwGs/qthsIR1K7
e8UEw+9xrVMeP8XHc5prurHWRY0Fnj2J3fr+8HWQweoaYQu2Y4sPqiKvd0IuLoq24/2ArTQxPYlI
Xp7dbwNAIg4nqW8TZzYasFp7BTQw68Y5s7q162SuNR1dC5/Gq5Izi3C9hvTCx389lQ/loCNOZTxt
LLLJEkvDPPt+Z9+LMZKyuQ47WFXp4rJ//D2HmNlxwqdTulbVow7wF2CcZlAnkW2xhQNH4Vct4Ttj
JSqn/sjer4aiyeYbgeOA7hyT3N9PhFNAC9cTHdUbMdN0ufvkl+epJH64VQTWqBGi2GNDuFrhRFbm
S9CGySt2JzSdTzeh8hDL9q+WB8aNcITORxo+cZ600neaG429bjB0sfOeU6NKrUiwoTUX8P/0nZOq
FSWw4A8R9jPqXoQwBaKg18xJWrDEiDD8YSqWxUdGzjGo3mVun2Mv9391LuqOFZ8jMa72nYCOpKGe
t7yRSd5QHg78ijjYK0IQsbwAbObz83dV0CVCMIax093dfJdo2FrY1yR9e9X9Fn9b+4g3jtEoz3i8
35wTJS6V+cRuYidRMxtXL9XkjTLZUeLIsa9lfSYTJs6UImuORHY7xb6thurzm8a8i3eviKfV+4iX
MOB/fFhV6rt5XEOU7ZQo5wmFFAtfNNpSa4WEyS9wlEIrpEOKfQYQummioPqsEmT3g4Rw2WpxBDOS
Ly5vjM42VVJA58OErxm4umzXMFHFIVFP6/SrG7TRYBcY6y5UnUMIZLqW0fJxhV1oJzVaPoAomN8Y
SdNUMFuVxS3SBuC91xEwYGDmx7kXyVC3ovp4TJ9BaGT7tQFH22U54ibuckxXBDdyMaqqWy15HGXl
pdpWUW3xyQ5HvtA/lxsDyMC7dE7pVWbKdMY0xbNqBkNEt/sICRYhLzNvLC8a/99vSsPBqmqXPppr
3tLSu0tBU6RLOCUz3uFwMe8uqBLVPl8myLafIMCg2stoRUNpNYwofmW1UsfcbukCZpKc2Z+si8C/
GIE8jEz9pT9nYvJcG6Acof5l3Ww6fFJMEIw8Vg0vH60EXvO7/KTqQLduMhkM5g0mo38IldKmxJdP
6yJ544wQrTg5dYZXejxKIGrL7e3Dae00siNSaczBzd3mzbr+DSCbxLUbj4ioLOsILfghnUnx6DW+
IUmvYg8FyPlCzx4iGOWJ+UvmxDxpjPIrInv0ZFV5XII98iKKnspW3VkpYlO5Q0C2yjgWLeIAT5BD
yCaR153t9O7YlJ1jIqNidqLKcDghWF5IKLWz93FAC8ArLZnBRxzv1k5YV1QIqrvM/50aaeiyvL1/
Ws1KCQHUd88EbFC2uGccbJFwEtMLOl41DwR4+66+tqZ7ZUf0b9qo+/LqJIHJ9LQdw+TVIT6SkBzV
HvKd0LtUklbq/EqIzQVrfz04fKooDZeYq+Au5WUipjLGBQkaOgVOzr6NfZ4NepO0LSPfck5dN7W0
eApwfzXso9HrETMpG3QY8+BIRWjXFn2n2l3CnThq4a2gW/t/nBd79QDNO/CYsLBWqmX2WyqdJWmw
oZGpWKU1722mMqTypBOLX5DnOazOqD8jb0rZkFSfavGMkpWLrWJ7GncHe6hG+wmdbmkto3zpMWct
ABCEa90vx6L4x4vQURAwYgAt9UBII6onxiQnyILiTiv1AF+vr2DKP9Q3ME4AWiddjUsHtfcj76ll
gSbsY1ZuCTRHHzcCYbI88ez5D+COxLLczpIh8lk658sdQpOTj6D3KhDfSHARL3WkcQX8ak9R/Gb1
NhMGjVMkdPglJamz5SFu5iES0z6rvHk0L9GuDDvr5NpMWvQnwGkfPigh7zDjIldVVs+U2vsiGywL
oVDk/lOc4FnveFaAxE7kI/1FOIvqCN2mW2Htzjg1QpFXFM+Yk9m0+HpavY1NDNLvwO7IVSbf/6jp
ItKFh5A4BSkmF0ZOLcNhKqf6nYvjXmJaG5zZWIZ21Agl7bV7MuqBuz3ZHi5BYk814SN9FfdwGt9f
sdjFOvB/2S9Tbgbnb7pIvyfzPBATZjHux0m8WR9I4VIMTU08fg8oVNiWfHnrFWuPb/zLjPmmfj5L
KC6Lb7ppICs6G4igL3Jww0ilx8hCnxaZibuCmkKbD+RtrbnCaJxqjiM4QwWnTTUK65PnOKhhHQ4/
JQHx8hIBfQxgUCsCGsFTc+bgzhYR6H9HvfkwN9hOufcZ9jlMEVlK1nkACGxC1TTe7gqJLBi2A33m
TKGx9JFb2Y3PSbavUix78THIJEZPHlQmGkjqOA0dCY22+Lu810S8ionRy7mJSjW5Ei7vw4L/e7Ti
mTRon/ZFQJXK6ZpVdKtq0vAQLocbHuvJC0rYR0aOnPJSsH3TObJaqpwSyzqPoHCmMJTLvj5gw4o1
GL+szH+Oneie3gCjVUU8GmsFgWEkUndeRA+W3rdvo06J7TxN1XgczmqRgorn4DFl/ufbqllsxLES
9qQZSxJz9484569elKvJb/X4d4ebRN1VgMUel+RWWnOqCDM9Iq+O4bP2gGy7/Q61k+vf2mWauRgv
vlxxPBdlraBDuMc7dwSNsFs9v7pU+8IH7TDxxIEUN91gIAHOU5HmzcPWgzjYNk38BGhhR/z3tUaA
lltUeemCmmIli/lZQWT859a78u6OaVgTnWCRKsSX23cK1v+sr7C7RjzaGtl/NDTy0lqGEUT79PIX
xumftVL/XZgu7iPOsXqgRsbPkNVQxlsPR9RCdjVpHTpqD//Jq4joyMoZ0OsxuJpdDSHYe3nZpMFE
/S2W1kBPdSNM5Ic/fNbSy17bx1gt0xmda+gHomVqaaEelgnVPJbZyQRmZaMhd2svHxwwtODRspyC
4IwM0tE15QzQr1SZFHmiEQQbDVX4U3+2DBCSBdUlOdf+veJShT1gvTDHZCNvR5Y/bb4AvJD0QmNb
bSqmwvzbBkqe7eijl1MnKg2DiFOd/YOVfl7fH5rOzV6B3uuyAQ31I2yc0GxgGLaAjkpkwOtbwv/W
O3Ds5wHj2+h1mq9XKO/DW06lPRtiKoF08uNJsNSKstIrG00So0PdXO05w9O9L5Y0xk7lcvP/2B+y
j3AQt1XjmkKLytEsSpXCm0KItFuWDAzacrtlogavgEinJLdYmAKmPtk6a5PRkUJtKzwNQJHNnBZ+
H2qkhUqVoXxS9KsHO4rcmr14rOZ+bnJC57gQUvoGhH+cRT/U+LO7EANRTR/Zwcmv4DTvz0ypIICm
IukZdhGZyNaLtI5/vzaT/CANDC4c4nup4bPyNVJuj0AOgAjqzkN/TK/UyliCqbFw0fap15H1/ZWw
3i/CDoprLff/zg1rNUpJooeKK7RgdvZH9EJVik9iRoOAz5I+Hz7puI5aIoqWPMMHw/Ksu5oMrvaQ
UKCUO6LlKv81lWpAoGg90AWyqOpSecUqA0LBSmLC9z++ilh9plBZRYAU6y6MYuyqBdBviBkYfyFi
Nyvz2ZMb/hp86nHbWBRGYHPAl5acRdAGX9oxBj8E4H8n3QKOVn6e1zStwy1f57KDJGPUjMfXXou0
B7TVF3F2bv6d821Z7c7ZJ5TfZyRmXlHfTH7ARU26IRFNsXyBghjkDqNUrJzKeqq4u1aZQwHwTiRQ
OxfEPqN15puJUr57/DM3Hh+uP+xAQwossZ0OZ8E9sHW5DWWsIsA1tzv/2X3VrElePdVughVWbADe
6s4VAsK5PXerimNCeYWrAJtie2uTQyFhBYsyKtDLCp+017UM8wWSZh2qekBAOX0ndoNjvOOagygv
nAtkdmX+mtQNRyD9zAd3IB8WFe/YbJQAhGeBbXltcH1a2iihNsAbNn5pq0l2nwyegyh2fFvL9cep
UrvxwCyxQxcN7SBKZkYTz2BKNHrVtPfscWD/Pwq8SsL6mqpbFsABAAflKbz23U/IBUe+xuA2+QWP
MpzsVaxknEfv8FIHG8xliQFLXXbYCZ20P7C5LVB1GO7ESqLlEIkuBhdutMu1F6WUfY8YOG4/VOKh
YDdq2PZTJQ7OeObyXcSbAa/1P+q4tN0AazziSA/Ss0oXzyzWz7xlpNpihq5tGD24m2Bp+HAQJNyX
OOviHYbpdUQT/HCMYkBXoB7Orcb4+PiY3pBdPGwVDrBIkbcTimOlJ6oDGw+KfkxPFZGiXQe0eC7E
k2v9nWpICeHC0hxgwgVCFWa4kMfhFlUXowfRyk2qzBqBqN1VY9M5VPToqqs44AGLiB5RFhj8GVIc
6A3OFDlAYPOl0wFdF1nvYopjUWbN+OzClSVZ/TfzizKH+7f3jA2EZRl+QTHF5tuLgGZ6g2ME8Xh/
MWUveOo6axs+CErMWjUtSyIkiGAlit93Q6DFVA/RsGzdqLjHiNmL6Lv1FljyO9uizjSg11J5/VbA
1su82+svCtweGyVcCwedd5RaVUuIIfRN93ABluUUIUK9Mtjaniqsc4YZbJNx8cQ6lRRQ4UFIkDqm
4JQf0WSel/fMxRu+uxfYMBVctP+Us/eCPdyqUKfuwktqrLSufy0LpJ+zlf0+0qDDu8eHkOUowp/9
V/3ck7r3oWi5cKkSNA4zYih1IiSmT6U8hqy7a7dFLnbZa/5eqTfIMf2DZqPHSOw7DmRsfQJgOHUY
2YYNnO9fiuetg48NmuKa+m3YaKevF0QohyZRo4Bawa4rGOXlWncqpP03ILYQ0Vu+p6pCPrqaiIEx
rZYdOyOObj38eN0bI+BqTPW0JmktqKqzTbXtRUxJT6MWdwOidtB/xMF3b8qNPs5CI81xEwd1OAfn
RKqbNc1g2xUiKNWJW/y2xvcQZI+jttwW8gz9ZCgPPrZV43Ohz1Pr6R4U7GAiwcaPGrk9FxOdTKB0
1Vde2LLJmWukWXKXZjFE2R/2lTCM2+U7yrkayee/K8t3pDac3RbpHJz7TBTaANN9UXZFymqPnXRm
cPM2DQfFZi4eXJdpKMAyf7LPSozYC0rQGmRSPuipa8hVA6P1QCi8YKk3VfvdJbOzJW1aw0Z/Yf/+
R/QNZqqZQhOAV2eUKeYhCjvPBVk5G8iLq8hhgjXFPNWGBhY2vNpfLbShDBFInUAI3Tazs/JafgRJ
PVe0Nvwc80mDGBnE1ff1MTifNNwKvTkavcl09xSi1+OI4aSNUIvGNvKzb756DJbCmBJ0oy2CKC25
YYdf/IGY87WxY2WQLrkkgI5+dqSriWqsDq5jjb7iitpSH5c1RyowvDe/mb2mBlGGjWCS6b2VD/ms
CAJUUuf/8zCJC6OwEGK7oLr1zbOlRss7AbcS2L3vDdICltsMWFZsu57DbuzXIjIwV/1jNy6e9Qrj
rmjTNQTOlXi+KfnFgyeW5Wjic+dyIsWFyYvTriywRDC6WaQEGQAdRjXrHW1lv/8MoHEELwkb68Zf
05O1URvOFO2GHL0doqOJkfGYFWPNJzqC5bDWP7K1C2g+smRmHf9WtzFcEz5CnodBqoNNYSY/mCuV
78joG3Yck27oc1hQHfEO5jhMpB8wGaeNrwMMPjjJ1Ki8VFZSjdhlA2nYTtv3FEZtnYvdLxO1gr6p
R4omH9wrY/uAFHU31kRhzP8G7vKL/nQPdFowKQh38yziliTDE1h//OLSWYU7xjPc8zFWBeBxtnK4
iEl0uippmn+UKnKY9VnorFDQWjGkiQ4r421c2N4z9YUgnFKm8ZV/SVpE/Yj64kPSVzmCYjaBs4YN
kCdJam+bc4BODJtskvSYWwniPjUxv0kEr6yDHB1GZTYc2I9Yph9dePfPCmr+qZwQ1UF4JHpzIXcN
ikFyKBMNzvT+Xv8NVy8crXiNlou3o4Y2e517lthgo8kJi4AWXUx+Luzlk+Iio2qznfHx5ZC0se2L
cr1QXid6aEycDh18F76zpDrb4l2h24T+PKMrGbdFHCeOmjV3mnA3z3adAklxmVEPkijnOXRKgzWU
zf//4oj9UI2l7QVb14nUICKy7CBXmdAl8jBEVVM00Tw5RL9ILZX/EL42Dl+FiwU/UWYWeArw5l0L
CgOoRVUg0xFCSG4SH8enuMGOfAqbfoFBsX0AbCu6iSNsxoClZB0H8WoDDJWjHtrnEyMLiA77gVNL
Ziri0PRvcBUV7Gy/tKDaXdrI2YiPREMNQuIrnp/roLO+WQtEC/tw1N9CJzjLtzn40tM9iqrPDqo8
PNRfQOBQN8j5ocVQEG9dzo7PMSSZzzmN8IIFcG18xOByg3yQao25BZ9ALRNWqKhh/Ba+v8/sx+U8
OPw9RAgpLz6WfJ8mbzv3msELQ8AmW32Cm3HNOl1EuNnf63GjSmqXgJpC3PN89iVbGA8MT1uWHxx4
Ut1BV8zOi/WWThZZTd0j/6UVnYyS1mupZ+vL9HavrCZ2VLystAmWBNhydyJTR2xAxCm3SgasaQr8
FRNoUw3y4BIxGVSVaZeeoECl2IMRUB0dtru28mFlQc38sbE2Ch4ojvhOXb4clpedhwcfhk9fjNXQ
3ar1hWqzkMaqcQIRmW6QfF3aGI1rAEv99svdryIwLNTMwQglaUGJFybtsmzUM7SM7Na3dFlT4V51
QqHdYZpjdJib5rJPwirN97J7C9USz36WWAqKYJZQC2X89Jh2FSHRAJ1qoDmvzwhUJV8XKTUQTSTU
qmta3cTdVTbDPhJiLAdc9hPaWquzfV4qoEIV4vlu+2qxtpImpRhJTsqOnggo2E/JsKFM5V6ZGlYc
f+RojKeqmj7xwGMjFNNnT1dmQfeHC0KXh7UWXyLNVMmRwRo0Fd0L1ebcQDx9FGDLH3pCoRZtlb+G
Ui6/xTXbCVD2vMu1U8ogjewLzFgQcaPerEhLISP4o9cLvi3l5sbT3je2GoNNhR4r4sw7HsOtwX9+
3SkY5OWHXP1Q8UCypkQWVL4bDEDYu06Sbl0r5e/RatJQR2AI3fW1PcWRIwW5UBzLz6CBDPcXlFhO
lx8qLYiomiZSQoR4YFoZoF0xHRgHGDdgyWu9bCCdkq0wE5B4XYchvIJ2Lkba9HixSPm8y+UKNBDk
TbnJ+05RuOmVeUISuaKIaIt3mmUKDu9mZLM7g59czPL5x0zaJtYI05pvu2tCeUsOTnOBjQPqcl4v
2vRWhWIWTK2hIcCHOHzyfUlpVKoRR6KpDhSUh0ZeSKfdfito2gUxHu4NlKUx5ZEL+IQ2adwB/D0s
pdMway1oXBVmISwJ+Q6gYF0LFecw71DLIKwigribzJM/Q7/p/Iy16OpobNsKcQBWrLFCMSG8IArk
eoBP07HFAo+o6ZNY9eTKkqahosh4wIFhJtCRzFM9h9DljKxe59OwiuxAXe3D6/Yk7OKkmE6JtnSG
IW5GVaGOxU5e6+GPExl6FJf8kPgxIG4JrXHlDB5XWAx3sHR7T95locD+l/obbxJjjVmstbudg6zu
LWopW0QthPfpk+kjgrYUfw4P+NBbw8IE2hFjD3UXZAZ1iEzJ59ohixT3ZXpxt33uDA4esYkrjM1c
XW1FfzOvXz+7K5kVcEAH3ZsKgjyne2YpYmH4nFSszyGT1DfJK7Q6NIVUhMgHwASSLC8MafQgmmrQ
39uO/G3KKFp0kyXvko5m1lb+V35vbmWcNrFC047CfMq9Zfi7FW297CM8x/OK5aGr76yPAX06CtuN
kKU8+8tzxUjdQjKWIjO0XruKNJ72fyx9PmQbuE15sRrSAGJ4sB9gD0tGc1wt2mrIF8P8GfNUTRX/
CPLatuUG+OCLb4DYz+gcGPaJIvDTcFF+4vW45q3zy25Q567l1dMfgdH6+Qv8ybCQAT7GT2C41jnF
wm7Qj30cNP7lqOJRONd4lflqbDoFIJnaEYeLkHSgB2NpIopCuRg8U58+zeNk1SIB7NiyqYGbZRqC
8Zs0+idtN5kF5/nWcVleMzErgIGpb3bT7UpVlTHtUPjJfoGoqljj+Sn4p/otWY0SGfqCvDvTwo0u
8Y9AT8S9OG6ul27yE2GUqEKdGyQFZmknTzmpnWWOogC4sWA5jGHv5kf7TkaodNb9Mx/XpCiipoON
mD0TOE0H7s3DykOMtu7og/3vzmckqCNstGABRig5S13e+MPHPjxXqk7/r3x8F6EOzy/W6cnW3c/X
un5cExD1IML+r4uk6XHlAuO7rKO+7+N4nGvSUGRTBvIAWZ/iLuXqFcZmLypAENcxoGFJ638wQuPP
3aqL5p8uMO3OaUQTQ/suvZkRvD9+kTWde89EBeMQGpIsBqxG8OWkJzLOhH8DXCnlfXsbxeVD+vOc
ahppHa5nyB2UP9RevY4QFBu/nyRZpfhkJMde1l/874izoopzqXoeY2e388e9a+66jHHdpPa9A+hR
9WjWQDlCJDEkXCym/GqyzPtVO618pWb+hW8wKZ9glIHOP+AKzRppDZ6L3M1skp6LoAxp1BTRjSqz
RVcPZlFqELjA/SeOkpX49uhLevTrrwFXe9bngfC6NS1/N070B4t4c7NaGGoIjY5HJiGy1EOtFsjx
9ySIELiwu5jsplKxuSQgLitzrIlxqQvGx8VkbnBQ+W6Y563YHxtYs8Qov4II33vkOtutaFvtvcMx
O35HysQ254B+Nuf0YMrXl1iwJCXQs4VRRi1GFWby1H7NO7jgRRdejxh9JGfBhHA+M1tPLOaig/q6
npVeE8/FRdoT2IvhsflzyvYTOoazI7SkihgsaPt89aGiaJBHWlte/GNGQPsuqc5D7z9rv3MUDAoQ
XkZxucY25mNyTPXu2pfQCq27Orx5SWNlKAmX+As6yz7MIDRgJI4Y+HMROXMCLOOtPB65u8tOubjj
zXPF5Jlzmsw+FxrPM8SeB44T3ZyD9qGG/6fUoFRQbMexZQuzvSDZWZMjFt+LJA9zijxE/MSkqo/E
ACXDtS0Y07UzecBnY6sCY3ONBMaBXKXM0mKtYnc7eONq2Uv6Re2tsFPBia0H2TxBOKzf7S9LFcty
ba0lQMu6JTTqZUebo7GwX8baI7n63X71yf2WOB0fUsxMyp1QGiYY3nYZ6eHtVcPyr//vKAzopwov
OqMkO/0f/vibLQySQHDSnsSdslUQySk2EK1k3Aq1aT9DmiDLHlbdtx7Q5ijva7DIo6VJFdK8oYBV
YQ8fNnetWa6s+8gszn4T5WOl0IQ6qv6mnA9Bjj+k3UjHtDy09xZcF/lWIekTXtYaOUFMbOP80gud
lNHwLcJ0n3A58+chRv2xI2axQtK+HWoqyrhesbwEdavQ9iwVv/3svudY/aP4nnCVTqEE6Qd274Xc
b5wQqW/cEDD0GQ9tBwfsqB4POcDt+MUM8xEyUpfLIE4i76iDpm1QpNHloKNCG+DnTK3Y1lDs/Ro6
sP6LO0SSRM+9DLjHmx3GlGcJuVhwLzNQd0lCbpSJoVCOOJfbMRZpFISY2FqqiUZuEhK4WApadt0R
O9ras4soFQ6efU46snmaTlARQleKZuFrJUA1NsjodTGKiN2LVn3URfN8WUh+2qtrK4Y0yEanGdGA
Q/is1PmMX4uvXjGhyAE4QCgQZO6oMuIhH03d8qWDF58EbI5Cqgkp4ZDoHR3RNtF5W+1FxG54WOKe
8nrJQnFyWKagel5RqDLec2rjLh+npsOXho7vtMsMKEbAAwzbTknOylZILYI6w9+skD+q8IdV2F35
zolfqKFMheB60qtPlV/1L6SOQXnk2AhkhhGHXzfC47BIUVwv3GBx+L4JHfKuwyc2X8N/uiUXP+Fc
2I6qjsOKABzS3m0zleRP/RAoD1xqJUnaVfcI76F8Kaco5tnEXN7YWevgzYER/k3Oi6BVDGUboLgX
0g0ztaOz3ilvwGLh3ruD08VmObCf/0UKowuSz4fVtA992O5p1UaIT6/C6YhZKEgI2V3JFhfZCLCW
QoYprQ0NPSn89JG61tW4d+837r8R7lbsN/CdAfJEhxW9hN69Hpz9p8KHSsA1FSbyEHY6CWjFJeUp
6BxggfkxVVJKaI+Od0PVotB22JsiWKkKfKhkrPkndocJfSG6+oZbBrCS/PQ8TgEUoRHr76LLsn6Q
sJYzKUPdJZMZXVlOYiJ3DSiaJZLHKTEspsscqX7nP/1im5UFk8ToKSmNRn0c4Sm1fN69GmTgLaj4
scLIKqK0KzNqMTDxGAtO8A3FPEPtUH0RTG6fmMPEwHouO++H1/aJLWYD8YJAU4GJ9P1jnpBrfQzL
IGIUCBI2XyAgGO9Zo3aOnPi16njRmvrTFAjLNXXs6wOPTqVnHsF7qT91q2kamYDqUBPRiOsk00hA
oA3/hCDinMUgyXDiQn6jRN/w3cPxzeeaxeiL0TNtaJXgik7z+Z1IyxOe4YXr0LALwNytk19g0Hyd
wC3y1uCHrfVRwfXBInvUnUAe+OIPUtEgW+3M99tveP0lIrxGos5FTCkshtH5YIkLQ8X06MgJuFiI
DIKuZ0U/mgHCEPriV22HCuvRK6HK0euTGLD8HNe8WaPKTadPm0WY6X5PjlbRsDtbGfFIR3IOj+aO
QlQCB0+WMMpAhR8AtcA9R3SciCIvPASC1XHFq0bSVDVjRMeLZeZ2pLarF+DTxGwasITgCZtGqxFI
O9KhT8L8VsHbRFdu/hn7SACOhSdkqXWawalry/ZTRMwZiYzhJ1ZiMXUgAP21iHqmMhiqyA+L+YxJ
7CwpOY8pKzyMyrzlXDiH/HJ53vhkZ+qyMW9G98NDodk9fmuEfQKmIxXpl+PlK6lMw5o9O2cdLxVx
aoiRNVFetBe5D8wbWe0XSq0vBTl4sCXyVd1Kx16VWSzIAMsq+fcUdK2mORhCM673qLFhBWefk7ZP
PQT4mryo5a42Vs+knUqs6DciPs2e3/7XqpBw5r6WTm8gjI5SW2QO+ZRLotd8KdQNG285ORdPIaKk
b7a0QXd//TBIwMb2Eysd74jL9h3TMEHoCV9JzFDEt1FMB+KygpB42d8UsAOR/byb5DZ1zcaT3+Hi
9yqfIynk1QsPuzWy1UTHsN4uLhdFb1XvYVQuCYh1XqZmtN9XLTzyda29qkaPJJEiexhkDfMOfTjH
1QQAhy+HNMaU12FY/bfpj1B0ORsO7plaMPqrfsIYC5LlnZOzSAFO7fqA3UUMwLAt0s8MPo/Vxs86
Qm9oDkwfUzhvaKXqY1D+xSXIOViPnrhGFi3h5vMKseEo2NByhe10i7ubIJyweExYQI/VN+BFjg5b
XXhqroH85zcnqGrdFQFetOSyAd0Lu1VcCW7jKzS0lLdFjijqxruVr4n1K9eJK0YYDnFTpnhXttY3
rOlZb42RQoP1tKW52+jFGNreje1e4djBQy3GnOlFdkUVoQd+MBvL7c6SDW/EOKgVqxkNrmYJgBlh
Mqyvtyy1AhJ8Z5HFMagqhzLG2m+IOHlWqI15ERCJs6YBVff2NzPmEF8mxjTJOJ7qxVISI/n9OwJz
jfq62VUh0bLI/+xs3S/IkPdN8f4zY1lWWjggy4XbLg92SZ3Woka4nesSUE0D9LJk+rjMEHo0H1Mj
+XJagvrVfGBGGorUkwinmTCgkfZK92eF4qccoYQ2isg6qy9+XdpYiitt08UbDHcu04VIH7T7TfxR
PH3JavJfSQaay6u4oBMxofCTGWwBxPv0UHKTDQ0ydWmgL/nyPhTVRyQP2x8JgtuvTjQFJVzJLZ/Y
sUpoXxo8R0ot37dgU3Swd2URdb4HiNwenvpB3Idfoi1jOVyqQWV9aH7RbwQtExoFJv6FsDdDfGkn
pYS2I2A9CHfPz3JpcUkSDcUyq3BZbl/W++TW0NNWNI9IDzs+dV/VHecyonxm34hyOLg/QUuO+HJI
1vPEG3JjuLYW5OJiu/GuOuuNx3nkqSbOCvOm/sWJ+Ea2Oa00ppw/RG3UPiHWJnH2ZRlmhB/rUJYH
c7YxkudsDOFVvKJf6NETpgkZEL5x2EwEaAce0QnqSqe6BuEB1SEOqaqdo1VGL3Z8ZbFX9+9aa3+n
SiJQ4gwMLSKaknIGrkPVJudOSxuery512b/AI7fAq2n9HsRqXSe3mL4xuuRxF+FjojyOKyH8YZ9R
UZBXT3djja0cpf/IGGGjrI3QoSRw5pm0hMcGHTlbyEZlYCSEZ0laS2mf4tl3U0c2I7gTyUHtzvhe
Ii1CJJiYsyK6D2T22OvxGGdlyMwwaLSue+Yt2OBUflOaizZp3Dwre9NlnJNTnc/KC4eQkfwv5Ili
MXg97DuKex541a8thtCl9bpSZ0zwAmRJzvjTPhKAyF/zZiVF/3YLkNlS2c6+abbW4WiWA0PFnqjJ
bP82Cc+RmofN75e9G2chxEz5THnGFVlRjfmzg87Jr2QHR+etavpBhhjKLnrjjksvGSFpOI2b8hAm
ilacHUnoG0OIAwBSMB8yTXgZUVhx6yzeDsMa5SU3o3qKKCxjkhz4e5lU5LHeqUf2MhogTMRD7Mal
an3LAkHngrGPlOrR7G9DffGF8au+cm0CX+o6yDp7Gmq8t6QOouqbDLpq32C7bNrz9lmWYRuZo8Rr
WcZK00G0wBUpLejTo+a1WuO4uznOlWB4+f54H0y/GS1IUjODsufL5ryMF7r9Mxxbe618zoWQDIjg
VZr4YUjhuxP0FTPWAg47lVPdDlpU3i0zHARy5QFrqziw6VBZ6Km2hNpmJXH0A2jZAm7umCBxqvb0
oWSQPAuBrN3P3nu8vBNpFcF+4k8vsGo/ZEda6HR2QSkTwtjKBk56Us9RRIspyVbBqn97VtMFnqr5
Uz86+/o5GGeOOct+NrtLkGykFNIVu3UBc7CYUO3XHp7xlSYTwYsRot3TCnT6NzAE+sIrt1DcolrN
ttAxmPU0LZyir14u6cn6w0nOenCcJVXQEIUq26qYLDAYnXFTSviTRiXIK0Tj3cDUNxC5XXhSoVHG
p1zADZPMRuW9IhQ/KfqZ4uxn17ZU4BixbMe3bz4LViENXHLLFaSPuBisG2VI+z5iOKPrlLiNcnVD
Rr2lD54p+uEvDUvzF3jqvMNxnpAzUPbihomRIUfaPTqG1//aIYwiAHyHaGeBV0f9r84idMD/OaAM
/82lZUPO81fJK+++HcK3+GRfAGw2eLqHvUandl+B0hA33xaXWYRLpESZpjzN/KSk6ioMPdyCLHnI
6NxxXh/9uYU6C4LrpVdcHx21wlVubIltdqy/FUbTNJjCNTrBZHExCkspOeozCWIeLvPIBMtOuwE+
2zVYCVEsUiCcrA2IW5+WjWsFmIk+IKkVapFnjizuCh70AsEWDCKcvkQv7AMxKEsomK6wxOUOE8mQ
gIaO+6x2E/dRJrnP3HdapB2cLh763aDA/FJ1CnR+sD0F7ZAgtScLQrojfh0FLDrukINEKfY61IRP
5o7VViVcxXrzR0nqmtmWDabIDlHgvL33VOo9GnrQ1d3tja6fCrFv5d+SiNY8L+HO5RZX1jPIooIi
YBZvgXVdlro0ieAl6MtNW1esYqWydKjThpcxUQqDP2nffLNjtQFZDn6iMxE8+lWp4KfsQ23nwQRx
XurE9GwYE/cIuu0WJQ0LU3k+alsuob7F6b/GGE3xcxeMdA+c8ik/+Ne7ugXlL51PmYRwtDBqD5rm
PNJCm9tS4TritMg3S4GEiWdUFB7HtjqX5vqkiAt/8t2+bnXKLX5H7zRqkstkBwv6Ib3JrKmGORPg
kedaTdu61ztjPJWW8C7WJGLY/4x+tralpBaIqlZQuDSG7CamznxugwU6mq4Jt8jca+U4ibQws4jQ
IaHCdRywnz1Kjw4+5dejKQ8FgazQMgVC249XXD0jlXPl9J63eAlPB/beIFBXrfw+KOyFcQ8/VanZ
/ZvchmpFAvOfQv/mbqT905yX6sV0bTuypIq3nRjx0S/wqj8YpLwlhneSZxc3pf8ih91+kCBAqBQ2
wo/axpZXF8q4xwVmFtdS8Kss60N0JwJ9fhomgH5ggC7lNbjq6KQe4wqlzGP3rVbKlJkynAFC55Bj
+VoltqzhRBZ5VEMu/SPO4AGfmTsVhA15xLhqAufwyZsCkuDYSQuNA8ri2HJ2rPm9N1qdm6aOOMBm
q5klH3BxyO6tn1IROoIA3RjKQUCRj7YlXgxn5PPqWVBqA4FhFwRWwTzkOC2x+eAsg1mKTSmNCAZx
yxLqia3Zs7yD+ZdNFmU3i7K0t2vnTdKjRBl85AfP9yGlvQ7x9E5+16uOkAVSzaUK+u6c/u8e5DMY
74r3S6OuY+Q6Ydr+d8xgRFwjZh+raupfTdJaYWS1Qpnh2SwJ/5qiOgB0ZDt4YdjNZshhhCrCYyBM
9IeIdKC8Be4llS4PoiBqc5RSWe4YD4qW4dex/6jhbc3xLWnjecqdNuL7CHCGP+GTzqJXfv1l27FX
ddnu1mzp7lFDDvFpiXta+xGXeQ+DHXlvGb5aq2Aluw975hRc7oFa35x6uAiIYAspbCV7rLBbISJ2
tyPD+8fz0RFj7toET1TVxbjUQqU0VOaNdUcSOkLId2/Yk7O2m5OJPq0qfZ29foUr5rWK/HPZv44F
XCkEx49HOA6I2a/Wgt4f+sHe/AhvS78XD4C0Vf4MB0WiJgYPMCjA2LnSZ0hQPY8ls+KK7qU0EAUG
8M/3BzQnIQUuwBbMxAMK2oFsrUWLzZE/vLh6JHtkLRCUZ19zvZAoyrBRCMov7Lgt7Y2PlKd2Si0F
SkDxc0eAtmuUsWraQN0b+D6X7E2IKUWhUDbDRMVYNrfqIgxh5H0qWotDzZl3rUG8O2kvGNSE01bw
U9YuG0Yqdthn3JIcEVWAU5r/VgoFLUA56jPJIFzmlSHODk+LNvBwKYBxIxo+0cWqJIubioGicnle
Dh+eXAvFRjvrWp2kM/yBzbzMoXeRP86/TkHyVJNbtY3uSZBH9GKWVpf01EZJ8a2s20tAZ2QVNHk3
JIpT/4epKEH2nJ+rWdQ0Sy+fqL9AkN/ds37aDWEsm978pk0Jziav4Q7Y9eV/NZ1gv4l5jdvg2iKf
taJgVGfl8Irm3ZuKXyn1tFNd/VEosehkH8DgaB/AHDQcdnE76Kf4OgIwrAqLt6i88A44bpod59jC
WzgjdKyX2lH0Aut//y+x+eeZQhnkLRQJBUoV6kW95j7pTF+OK1lSxFmxkoqJXYcrW9IPlLgDx2+p
9cHikw2xaSttEzRdEr8T7y7GYBzpuB7cfABUs0WZ2xVtkUtgIteRIIjXW9jG30fxsj2YdyCfeR4A
GMP7THFPKU3TSLWG2XOTZUZteiAd2rymNVYQxFNIn15ky0dfs+P7oEe6Aw5iOCXgpPWxfgA6aDy/
GZ+/pYTY9LaD15Hc0/88G4vakpHhA9VbvuciBN3cTvAoacI9ci064vxg/PTk9700pxN/hBW3I8I9
fLPr+Mts0r3UG+n543/MAIIZdFSB9QdTx2Uqe6n1M+Uj9s+1DrpNGmgwG3vChuxvRcApzmZGMV7X
e5ou/3BfASTohJaHVb5a6CEK+hZly73dc8cc3jUKZ9xo+qJCBVhM1YMqEj0VpS1aa7DpJSdOLg5D
qVfat9uAPE+cP0lG3L6x4AxWfc7QrhMmHmER7W4UEeXr9mxH9FWMoUTRNpq9Q4i0DcRBt1qWBBHY
jJ36jUFf5Mo7L92O8EiTq8V1VMM1pR1UROk+m08XYjhEP6P1vlZkaFglY30cCUOvX8THrLNNIF0R
aCiiAibxMm7fV4IxOEmQDO23lrddE9yDFWHi3+fqtw1hNrX8Up1FO+bCRCGT489k6tVhhtc+U8pY
2f18PxZRpw7ptUuOg+jZd5u+ppPDJJ9Kq9SYaiIcGjXh8qdOWNFvHJLt4bN1sRjX4L/FbHYn+dvD
EGnON1vhpb+wbDu0NtGxraTG/q7xyITUeTk31DkKi6fbmWZYb2kELEceapzRRCX1uAA1TPfeUlMk
sv4ABx7TmdFo+/jDDIV/JVimoMunZ8s2nIY1msJo7ikF1U8kZVI7iff47+p7ARduLlMnOca3JTcj
mbIGtwetOQjrk+is7ISd9333SZnjAjPYNOc2IyqS3xvt/mmzYtGS3aybEXtANAFJ1yqEJwuisrpS
UG6P2iFI+holV3KHwMLejOIAfOCv5a5dfD79Tow1o8Gwj1onDb0IW7NjT1BKdWMXLmf2lqK4yc/w
mo3XNpHqx+THq1kZ3pqYw1+nrTFauER5mDJwitzUhyUp+4jKLNLdIoOzdyya/0n3HtWNnksMEen/
IRJhokuAgNK/kSio2PfXQOLsO/CVVxSicz8R+EhsMS+Wg8o69KRlwz/lbm4iI15tol6JsMx8B03X
fjTZ3kjds4bE7SRLlceiwAo8mvb7wseLPlp5wH7FK7axd3Zm4i4CUwbFUefKYbYKIE7nPMDa45sG
3rhC0r6QtKxO874Fj6r3jprsKmSrTGUMOAlp7INlmolWQhAIUbRw+A0NFh2raOWOAzuMtzzZSOGO
L1QZUumrnrKZxatLxjq4YZvn0KBdFMQKc+l7URkQHvxAtJn0aUDGzwKTGL4hKnFDd+NugrUoILnV
vY0iga8awqtXtPlk0XrLodnGFc6m5zayDEfIn/Zr30Gwn2cMR6EVkRytXCKdB0e37WA/rECcVWiK
s2A/l26M8u/aBq8TNX/kBRzxenh7mXQjMJYrQgyh+QqeKlgCAUQJa9OLemCp8RFQiYcVmJO0CXLc
GDXPAJhWVK+CV6dh1NGp5uvyE9Wy3aTgx0cCo71pJYr/nQKwoDEJ9FQ7TGwf7O1Br3p3hW/xFC+c
V+JBcicdaevhYVfCxlehIl5cZzwxA+x1UtUecKcN2NyiTo0igccrhAwECSTX2ILHm2+7piyaMQRv
lfDnTXEscZ5fYLNPnQWiRxpfXmwNwyfGeFU1Wqzm+AeyqIDowTTQuvBFSzfKGtPOhE++/8hedo3j
Nyd/bCLBBFXZMzqiRlWImCI+c8nY5M6mAfs8J+1mW5ASA5NgfCeb3c5umIY2P1NBKBM9HgDc6B2D
VLD3B/LQDyM1la3kMYs9GnAKvDxoFfh0yAhFx7y93SlcuK5jNMA0SfAjxGvk/MFiFZ2EepqV5kEA
kxcaeXt/NEaAxOUzJNGeQr9uwmdywbWT4daL4jlC16YX7GjVM/n4DX25AVBwEdTGD4csyCJ6Z/ca
sM7ngwJQpCm2ZcL73oIh8bfD2+Np35mmxiSpLIkt10In8ZAeoe8LfOoc7PsCqZL4TvsMQbTVDD1c
kEfD5hvy+5SLefmOtXFTkSX/byQBGG+/W+xXQcXHAFwND5wKIvnn89jtCO7nKYA7XX9LXgRiXe/s
XDRckvu1QW80gK8jCMwzUMPKovR6hckkSZruuuqEFYntLH66yAd+K6UXXDX8QhTFCVK7FwVZFM1S
k1SYK4ZeGnbjhnzAA5QMFGTDnYLPg0XmtEBrGVVMTqQaGYAzkJsCqkgr7QHElSIVMmDKUt/FkIuq
2AeS3kSVc6j4MN/AJclOcvQboYcBRLXLzLg6dizdBOEpKb+a2QEN1/fmSvgtETIlzG/CkhDv7HTT
SfrzSsXIyYrPzCtpDLyQ/uR335nvXrR6fbu0b49UvtISAXSs+hnFZFe7kONa5fhvbDZjNKNdDJQ8
ISQ7nd7uAqiRVJs0HjToL6hSaippFXMkArx1BHp4bFZdCLVUl8Q5pA5c4B4BocYvKUakySziSiyN
tAOwfwzS0gw408o29qcs6u0uGgBRj3CwO8a55Px00TC6PMUZipKWd39qtWk8JI9oweNMiHysh5A8
d1waTjoxZcybal3yHMeojan7ok7wTnIeLVFCu2iKT1GWYNMCy2WACKSYOn0f4s44CYjsbElhIq5U
ZUbCaIBAKK2Fmdmceq15ztiWvSdBdZC9RC+3cQkfGZAjUANeeWDrHAt9bwQnr7X4D2+rYtiXinPt
uIuOdAUaIOW8V8xc8N0DUk+redpmfcKdpkxpJlJwviwAgh7uyJJGjrEdgRPSwyUfwNgJesQMu1K+
QqXuVYXRKIPhmUbvCsmhon/5PsLGBVMgRfg+OoRJCjNH6sjM6PSV9HCJT58S2RnKh8/OrHZbE4lj
1Dzseh7HPunRlIyAa5BowEGCEgjbSuYwDCt5c1GK8y9HspfFBGCu7lwhmXKf7c9clWJKd9kucWIL
HXb6owUYfNopmlgQaw95v3+krmMwmTQuG9GZ7Z6g8fYpy6fmQ1FIQZgRk1Y6kzPpgAZ5x6BXMZ/b
BO1a/0nGcgKBAJ6/kttDKpT7pjYwxqPkY+H/EPkER5cjkiX3sVlIXnwz6YxUYGzHxxFYhocXzXXb
+xtnifwaK+c9B6+05uMESEZEK6wqFVgVCUt6Oka1hdSy775cgzzGRx1cVlbN7WywcR5Wvk01i+cv
Rb9JU9YxRzfTEEvKLeZq/ifZX/mN8vdA30DsK1yRUxs2tBX9rwL/J8FaUyyz32ovH7yaO4hAXqBN
3qVLkdPvC5imdTqYe7FdSBhfqFzgBBxtse7SLnt0ZnLDK+QCN7mJQLiTlx0CFViZJS/ecDb8nQx7
0Ddl+bCW5N51n/zTN6Inv+hqvoD7nqCAJsEsmXWdJBANmAiHdraF86qA76PPeHIVylNfAnsCX8Q0
Dpi7Nd39U52/GKm6ig0P8P0HAxLpHANdiRZgUPAA6cv73T3W8BjcEhF3DIR4j3Imi37sZSUne1mN
BpOJ56Aj9l4/IKF+z44mTNQ7joBDsRkQXUnxSXUId6L4xd2qDrxI5MHtnz3QliDF0UvGg8m7DbVi
WSmXlIjyUq0pdjMcIHSxiIHk7yEFPMK0+hYXgu8XEgZ7IJROtKE5zefZpDEqkPm/mBoHuxcXa+N4
umDVKzI2uNCaukQheIX63IWWDxpwdPAk4xVDJG5NhRfSaZQEIo8flEwTzIO5bIpKPt8rJ5VLvfjm
OpEvyUA37ZVoT4rb+5ypJMpoURevtEil1q3eTOdyWYKDOGi685gX4vqrjSGXzll9rWU/jcrRX0QJ
GvAVTM/vD/AhjtE2JdJz0O6whI1X/MIYZTZoex6dKMg24/9qJQzZuQl1NP+DbekzJJfRZyJVXkgL
A2Uz7EXHxOdSgQTBFC4cyQqjG4oOIL3aWarmkj1N7Ps2+fNLDo1+FwUOeYy+w/MDFleQhjWB64Yo
FFg1jaVD2Dkyh3mnJCkJfw1z9ZE4Vh3E/tfM7V32GsBU5dij1zpInBRqRfJY76rvDLwX4LUokhbi
NFQsR5/hXuryhgFlsDYb9V9P+oqRbRwGil4wkPse4hDXEshbETqTeCjjHe+biBj2AlJtslwUFAV8
/sOHxjAxoamfVz37T/qzY+swUgrDbmWMFx/VCxho5RRNzzwo0AxXUobpoH2xMoMHunoLRvZmswU2
YCK2wTBgMom4w10lnwYvOlhrGtZTynwum4A85le5iWpw6oGkDfakv4bHRx7onLh6NWxKVEU8/BWF
PGYN+vBVhQlXMSZ5rVUjFYP3KB6GOtTByQ1S8ZCmt3jk4PSqxK0wN7To1CaI9WGv0iR69VWkHYEf
itJAexNjiPoFf+HRvqvOCpJwkBhMtMMf5E8quuu2C81Sd1mUOpghF/Xiw1QjLyj+xMhW0czeW31Z
kn0FVQgG4zd+yZBH9Pn41Jbb38aFOoGX7ZXGmOgtdPPi2mAZ88KCzsGg8Ix583Wg6lEfkxROywut
6HH7nwyfR18KfrlqLHm9MvEIuCOr1ads/5V0RYdRHEOTrMeyPwyasGyhYBAYgMEfeCnTup092py8
/gWBDryBPgZOVEqnbx50mBcpTL3E+X8NIx4+onCwDpnPis2X7fhK2wP3saqsoHzuRJAlN6wVKThm
t8PgxJOeyQ26zQ0ofH/5TEhrkB4cu1UiDhqBMR9RqaBn69DD1nz116BGjfzblm20zDkyPodSUVji
cBDcPjew0WjgniBHLyCQIjGNxCiXZCHdOKKXoAmmzw3ZaQ0D6NZXNbCOfhgROlLmQ4ui2mNdPTa8
HLzBFUZy6gEqoGTyq8VM2B0BIlcdiiO7a+MxEBQzR2Ur4tbJhnVGwyBedtlJCCBeF0MfsiJXaoUS
61zd+GYcWxsMt5je/N0PkLd6M1t4ECDzmllyfC1PWWVfYFPOEkhhx16fC6rY3U56UtYAbe8CRcIZ
k3kMP24ovZSxXUjf5PmTnJkfyID/gE+3gy0Tbv3z0LUzF7gfNqdf4Tr1cBvRFL03grjuGpvm+BwM
Y8ww/cDWKmeO4jgTAObnKR8ciUwKylADpl3aSknd+qiZVfVHUxCtAW/ArjNC7haVBAg328a32+ec
FY0YBBDhDMbtPyavd37tJmkomj7LwUY6cfMeHQxovWEhB1InSzM98Vcy7ZPTLQxj/JNHRfXxTWGh
rT8d2I3DZ8Ld/XMiUynEgc92A/Ra6nKId/KdJRFhdfbSz1VcUZxwbZsTMzgsbbueoSrEQcFs3OLb
THLyIew8G9IJAdUcQs/AtoTwXnyBaI9NDudjAs/XlVyt5xrPL0ETGe2+1xozyJw7M3JjXr2F8mGn
UgAh5baiu1MAxuyetzoTRDxwBYRGAiDnfzGfYKGQYkbU+oGg+xWUxz6XYHhgCruDFbdNFKdGqTBh
Qobfj/9XBqRh/Z8YHK+vR4VfQTEC17mLyclYX4PG3WGxTYwJNLQS8duEPmsuUyr+mf1lhoWdvA4T
xYgzM9XbRy5HTfHWFgeITk+UOu7xNXWcWRcFaFufWxvp7M7B9BQUg16HFQ41ScefQBSDrEmUapcd
n8ovj8Q+MaLaDtz41YyCshdr/IxYQxJnaIzMLcpfhcBsvPbEYUEv8qdTQeMtMO5CGZQ9DIaz32Lu
eQe7yPBs8eE2/+7ZuCpdSywD5v79JpVVh79o1bol+B2vAFTUAZT7n7ykUbY3F1BK3/uhUidf4LO3
EC1yDtGtnnwVr7MtB1ZMZq6X6flA2CWsPl5Hh28lk69agF/CZs+q1ehzikA7apuilP24yWIYakb0
7mZHwdxIS4SLl7mV1PYYxxY/1XlV7aylOcsyymPFnCPBR7KgvuWcNhWZ5pkeJSXYgI8tZ6onLgix
DdxLT/FS60BJ4vTkXm/3YDQHoPQ+QK7a5QkSZOBoOjPH5N/3U3GTLTTy3x4mTD5l6Q9+nCzhaPO8
BEQ2z9gVfuzgnOgZikE7Lo+txnPTNFgwtlssn2ey6k5HfRX0cASHl7aROn3eaZHtMgWWGOzh0N/O
a6MboTori/HHHi3HP6ppCY0fbwMy/xljTgPRnQO1VJGzhEI1V2zUY4GC57RN8Ja+hH5KRebUFYn0
0/WbXbS8S7H4Uv2CZbOqC4a75c+32KSzxCd2csagCMQbWdW8dti5pSa1SVs7pUifzvrTHcUQXQuv
9gfjLOYlb6iDoaQ4+KqOH5cMAgtB63IwLdYhpMxBx3XqScMwvg8ECo+j7z0XntL+cgUvFCOZVZlX
x3iAy0TnNWN4ygzX2TOCHblu6hRxcK5Ys3wrkyPXIN+57HQ2xQmhDFFJ6DDOtwEEQAyTSgY5cuDt
fcJa0b4v8SW6lucIC3u5XpXpcb2zxLgMgifM41gbNZe99MLAoJH7sHM90gmYA4LHRqi1aw8d31ag
G8QNBzywBtv9hdDR2rwA4t7S1nb6UKLYyXklDblm3vmFj13/gK0szRwh+P9LzspudQg7vD6IrKOQ
BhgBDR2r46sPOLOKj37Dnv04A9xYZPHF5x7dOLZVs2Hq59mWJtjSZH48+EO4h2o4pyeUbcdhZxY2
ta23AUGoTJee6gWf0EONniHLxDEYJPmWs3qXl7+WpmKWqip54B/04aqriOdpk1mntk9524El90nw
chdHewdq5ok2kuwubx1I2+weCV+0ChUJayVyad3Q5pakKm0/1f3mjlqsyIAoUGlf/wOD9ZzpRMEx
WqH7wlWvbik7QrN6xPHMJQ9UAvp2/LAJqu81tiNBEO5GVoIPc1QGtrrK/DPOibTBSz1hG4Sn1u4c
/rgJV868/Aygoo7W6eqf/+nuVedHJEpcUg/7gRcD9fHXbSq4yDuuH6X/BrgeMvmIadKyZ0GzwnHo
uZHAVXYBop6HQsw2wBPK/wbGQiD5Rjrlv93xB0fV0/fkFZMMnUlcDeVG77CQDun/3yoz3VWUJ5Fs
Bog/enkNVjXoD3fTL7oEmFUeg+7aoHJGdaBYUfMdkkn/2KrdxcyLp5WZGUXpMPPs83wwmWCfm4Co
NcSRZAp5awaL0hvM/VLva3cNLStWgbWSMBJoTgmne/kqh4ciHuG+tllOhkz6F1XKS41BYVU+W9Cn
CfsrCeAcJEKWlSjEMDkIjftIEJtpe5OXcLG+SrRqMxZZ7BoaKwXZsOPc7wKb1ZhHu/IPCEQuoLeq
k0Xx4ciU8qj0wp9paYkwhcNJuoWkGTFSxpVC81MbCOdpIzbLClas4Hg0wKNvEc/IMqlP9cJdYxXG
9FFaJElsJjNkLoBbaJGOVENK1mQUZL2sR1a82/r9mWidowwZpGbfN9KCWCTYdS5hGxN/1ODdeRoM
TNoIUPJLZOAAFbKHc3PxDzlab72pNe04eyeT6cOQthW+O44z/BNjXMs7yxfW6hSlOG3wxX+k3ugx
ZxgO6WF+GHeiCFi8wcgIKv8ptQv/FC5RfbDnjA6Dkr9HBp3gzAitl5V1Dclu3Q1TGGu8tkPzZL7T
bQSXpi6VDFIuQUuJcyEPH+/w7XGXSiIQ0E0YYziR92RXOd00hpsc0NTmBWXxrrGDCR5+n4GmNHmy
xGIt4cLr6+dLScYWmq4IU0m0THE8OiTnf4KSIud8FGWvSjI4Djd0xj/rThJbFM6OalLuM3bY12v0
mtjhU6XXpkmvcpB104F8BgrkmFnFsR8HPvI+u5wJntTJ9YmNnfQYCA4rWIRJ5btABq0nrRTKdycp
d3KLbXBR/nk4bZHbtCCyzSPkBq5Qglp2uwMabN5djU2a1fKGXJMWKBKW6pxYhmaD+m9x/3MlmZRF
QYKkOm0xodkdPJ+fZ8b7cZFmV+1kxdQvLI6I/mG7ZOOp7jroJzgF+ANb50E50Bqoh4lrLYLgACyf
Qg+OTr5FHoMwCgeyrCVorpmZa0GFQiAN5eKALwslkkmq7CgdWoUKfDaUSNmnJF67omBaSmUKGK04
qnSGu4PDnY5BIcfFqwzCfRv4YKox9+jNj7SHrzytuvR+7j4bN1xKkEfiJ6U21JYbE0vmbmQ0Nnpi
eryji1oexnoBJ73pqEOcH/JeP0Jvy8+6KcHIvvOHJkiKLy7XVC94SATV7kBei7CgbBpYP4dZpXni
Y/odg6nWYv+vuWUVtkyN/PWYI8IGAj3ftErA+C0uavD2edBx1fM+V7Itt3vywmpkTzkjQTSQloLB
fhJUSSYpoU57Gmqs+kuJ9yZz4XY+QK+CzlypuePjddNyJWqtxEQ1iT1TOCRSrpLj3QR0Z9tJbJgv
Vx21u9gvb+zQ7oD+AwFTbm2fjJRh8+eZUEo2w5wCROJz1KiI5AR11wTISDR8NPM+vbOPNIzNCGP9
44gD86GGSlseTzd6XhvIyH70jmWyUgzpoDqH4QoHJMTeFNeWUvR9P4WoKK22ztU1CU0ULcMC05Kp
sowFrRDPWdMx2TBkXBQ9++0K38g9H9qdnX1m6KE/PGscPStFDEH8it1NqDl2GH4gkf3K8Tnp+BAk
LqZTB2rOLGWKlKxP/FnwB8dTo8k1TzbvYdync8f4F8Y3m4q4fEMRLwbK256AGRrX6XjrsdkbscJq
thd2cUvipie9xBSJdNUweeF2HOzq3NFGGxqpfD8RRMcjURXGToanwPlHzdxAm8NQs6A6Hb3jouIl
73WEkaiMxTpyETISRZTxo4khiuKyH/TuZL+lPRmysCjBHGPebCqg1/2BLjTmSCGI/DbY1fu3mcIW
DgIcr6kNGk5FJJ1Go2OcPKy0dD9omgoF8KrpOC56gHiJPX+FrtytqYPP5YrXKBscEaTkYmRErEhT
p7nKpNIFOwHuyYHq9xX/Z9YH0s+XlRsggnG2MUz/Vnz8KHvagwFZnZ+33sEjPAgi+vVIhY4b0HLv
/mKXmpDyeWowQ5Wi3defDK5acs4tESVfuNlZy8ntve33YeckKKpuI+hoeJAqvVYPbuwh4aFdEt+n
3+Gxsm7SlxBhBz0OrOwAi3TZ0YWtJa1AAIVtFNwNXZUmB2k+N5pnB+4153H1LtZPVbpghK3M+LUH
RhLSr+/U+vHDxjcnppV6KntlW80TzHIso/nwHvAb45Xf4wu/8LqhywcAJhHH3+9rB1dMbUzSlSkP
JYT6I2Ce6d99WCWa8i4Y3R/RMY5IV15bPwKB68T+QblcsyIUYBP2yzitt9r295xWxIcXTNv9RHZS
MDhfrI85g9LyvZ5I+DWQb143Y9pMBhdJ88sLdCkz+VMqb4iJlXGNo/N343y/saBEti+kfJa+sdUB
GCkkbNLgsANuTgnj9oQrfz/H5Dh8PAhsZXOYKBNvtOmNAMB2mtYBmg71JvtWgsZgtSglDCRWpwa7
uV3/Pe/Uao3YTgbR7sm1mX+wGrGUupY+kmrQbbkBuaBjUlKwL0pD8SIIeOQFQAVljOZTkejmFSfO
EXrlFLM/6Ec+CzWMnvwnksdhWV6aRyEkbG/21+GaoNG0tPN1rXCC7OCWvInR4l374EsmhcqHpzea
7qiUQSrmPqwivtd2fyAlvPhHtHLNyy//Y9DLLLfRgtqLgc7Ql+GXlQ9Ct7fXYmJRQewdenNaWt9z
urfQrTHoYBjQmnFeHcxOCPTUWb9ghzjrS/VnS0m4bkfOmm6s7KLgQeLr7CvEHVQwlBa8AKPxTR5v
j67zcJvpJGEdvJD3Ofh+IEqJ0G96b8pA4tFzmquJE7+MBNoAIYsPqwyOMMrtoOtGTPszPKkQcR8n
r0iBgwIQNqG7rePEfS8KtMNOP7I1Nbh0ASPdnp+MrcWVQ6Mkz1kaKrq6oOEf+bf3xNGr6mBpcST6
aoY1mol8KnvrWoagf/r6kOyEqAr3NC2DuuqRJk0aF2Kh8erDXs3cY84mn4Qg9xEvlK8VWIKiMISh
jdVwBJGEgixwWZtKoG9We7XgdjuQyNZN05k+s8lEBgSRo499bKBtvMjSj2+FEj7ev/hAYfBOGWIx
bhC4HdlHIBwPXxOR3a//BzLXQqXYvHCKiPZJlNckXlXacvRt0mOl0sjNJPDk4K13LaRYUJVtMEHE
QLVDi5xgQBrUuEpyf5VNoSZ0b8wlMPiWHYGgHnEwdwMBPFFU9nJ+uIkr3PMoay1+c8z7BIP+zu5R
YhKA/4Oj2N+ToW72Y2IRG0cWrhH/IFTch39T+VWcnly0LJEutCTA6uR9lrq/uolSw1PzDHZo4gXu
6uNGafR3XOwYJ9W4UNJolVPSZ9WD7rtUqreSIUm9pE6iGST8VD11DXXRkHx9cKyYF9liMCfd0JNZ
C2wtic7XgZGI7y++YUNEeAaBAnLJLxacNkp7SAWyp64Fz/35e0vjkl9b36tgBzwRuMISkKh/Eip2
gUPAD6bGpqxTUko6QYXaXfQEF3Wc70xUb+cXP7RDQleByu0BFiAROjU5ylhBjH/u7oztZoyejRZm
ZL3AG2uCzxDE3vq70iOTd6Qky09ZW3SqF+MbmYtbJIoTWB8ysk7wIxnI5niK8qmod7Uy77xgqkFA
NOJ0wlb7cE/l66Ptd3zMvpwlk3zYHYhPqWqMAqkBsxbkcabtU6azWWw86MM+iOfiPP9e87gCwavc
w9cFzAxX3AiN3jhkLtQZgQmL5nYXni9PpSVQgad2L+aLH+chWWC54PhU0NYSDmI1ZLyDcsVLjqnH
8/sjNU/47Hg/Pq0go+WOx/UeqrMegc882/bu8py05WIZ/mHJsEwG0k4hfqLpOpk7E1VjxyQ5HBUz
IfVZvwmqV6ko9Hii0+3JwBo4yPJW75kZ1cpnOG/JmSUDTjpmQ1DWqLGW55QF7U27JE5mwqaNPr7I
LLNrUgFcn3yhjHG2dJjaLIWb9g9Z/t2mfO7xycwkejcDQpCxI3kvcLympy9goN64vtzFvUGtv8Y2
jrud0pWkzsIGA7qLFFCX+Oe4jpKKK8ZYjLRaL5iNErPtokYRxdOJROvP5w7thirvU/gMNs3AMsUy
xUj9+NV4z5i2w1NXKcbtT/lg+Pn3NL38sa1d/ffLRxmKUKuo1ZngautcsaZ7rXSXXvWsF/JX2BB5
skg9TCI/17s4wM+LjzQP1dirrmXguQi4hPfpZQZMrDryCoovn93C82U/cyUhtVpYmrdZtJKwolhz
hG6B5klidI48/p76Dx+35UgIVsxz5N50y9UHUNWmCZh4uBiqoEfefdvduMmzqhUIQkkeDi/gPCqM
lVVtAtlYfNAkASStkeLXY6O/AsyyqyfJ5fl3sMzeBV2hnCaswmqQyj/izEdpUAeqPk25iYPsI8sV
usgBjH3HfLG0shRvTKwcju2+9zsf9sbOypDNRhllNHdareiNfYimkn45mJMxvXaR2C3aIyXpQotd
1a3hpfEeEg2cct51hpMctjh2KbOsltNGKxTCm4lYc+qJR+J1BSJzcMJoZkfD+g/jR2oAqTZyiTKS
uHOMq5fb4L3N0j1JaWRfDlNuBu9mrQCjvnMdaRCHPsIjnjaOSntM3E4cnUpbLgvR8T+Ncqj7dh/S
KszSpl/WLg96ebQFQOhZCJj+njYEBwZgQDdOk4Q2WRhl5T9RVOi3yA0CD5uAYHm7SmX6fpRCBM0M
1nbbdhYF/W8bt0WnvzPUunYYBEhWG8kKrMGzE21RpKqT2MXyTHXoINABs0l8wQg5sg65+SmJB9R8
bMMTYkt9VAa/1Of1vq/zxIu/jxYCrMyxUZSeD0GvNbzLuMtZL7W4u3WBl2kPf4/zs27FujNkNvXM
OXuYTyux7vIy7Hs+6d+qIG9csWQO+aJ/yIV3ws2YX/RhGZZdVB29O0XtkLd7q2AUIBbVO2REG/96
MzNYnWu/Q+DjNzCYDfVrXkaWPo/RQK9srC1svP/utmPW8z6/l0e++spuO03K6CjGS36Xp4la+v+7
ubVsHNER/uohdtdBIuPtQs3twHf/4Sm3Zi89hIp6n9fvGqC8liXmaWC+ym/7xb9Abeghhdbx4uj4
xuJakBBy7UqQsYU9XyWng05bzGydCBOJV7/Msb0sBoctYHqpEpXGR8JeZZLj2WNfF2RRlHqxl3Wm
W8RFTUYKlo/q3vUa0odyMpRLI16vxNghfKi+Tmr9jEOXApSMpcQYfM5b3ysEY1sZOeY0F8YKaJHW
R505xVC9c6n/Ljjj4tOBBjBj7OYqoUWOGthM+mJO8ymHG4jhFCLjr2qwTOsYsaFN7pxTJwofDu//
JkrPD/CSc8oMpcMhkjnhfTAk+X7uXawJ/TiCaTMaIjvxXjrIvnlyZIfqb6GztQb+vGA5WArDF5zV
rd6A9CvyRJ6uur+dUBSmDwlM7uri+XibIcj3Ze/yeDDzs2qARaO8TBiLTImykin36zourcZLtCHc
KA5/ISJB6c0BSzMjVithACBfVfK3CwCfpHiQoBBtm15lH9iQrwX0QHSfohIEaH5I4aGlt5D44bgY
Mt2My5ap4sd4KE/j1LGSlqxQ0ZWAc4ZH+OjTSz1sPgW9mrSyesITaDg3Fjd8/D+0mT76a7OF339R
EJgXo1nqGXWs0fjm1DW7V1UFAiRTkga2X98kUlAQaANiez51gUlPhc5UztG31//Apl+dK8FedqhI
WIDz0bpmsH0NhQQWpHQc/tzaBg6TbiynQ4mXLKCeBIX+e7cZRIhC+z9a8YIt7rWk7X3JvMztI2ct
uKvBCQdrNbN4Uc50k6ymqM4WhY9eI7WkhT8o6aJQ4npQ2XYBaHq2q29yXE891OcGEHlSJOz6EN8d
hVy2n/gxtwGuJfwmkJGw1ghCp8UJDXCYRImO6VPXHcl2Hv80dbynn1RnRMkliU4xUH3V8iO4v5lA
CjF5FtXKDnDMfRjGd1KR3kPTrOoDfERcmoBM0xUkmw3at7z4T8dcPLAXpxlvCsmmP89Gx6tNukjN
CUGEB+XoFrAedvLsiEnyU2u8Q55m2DzsPi/AnCyWrto3svitRMtVkDMdLlishtIngCB3e6iIz6eU
LJ/nt6oFtZqMkScZSX5UBEJWc5OY1JPHZMMaIKnpF3j5M/pjp8TWw4chEDYeAH1V03C0aeB+kzJy
2drV+hnKLAJkuiIQJEa8nF5N31AsEURxoZ7ZbA9hTTaOP4KESdu+5KYPJYZinDypJHL8eJO1w60Q
sfy9XBIRvwaeNWphDnJaWH2hRdfG9ezbbsdk9BHl+CrbFI9lq2VpUtoGmfdhwz8FY6C4TUy0pgJA
UsJOWRgKvQpdiKz/1bnG5dgWqZCG3HKwEf6Jr2IiAxp+JcHBmAcBccnmqBcFe2Ax7rcPxp0fCr8s
8cOWwNNqlF0W45eqF/XF4QcwiVD8zKi05ZIg7myFdsGi14h1wd2iXWGAoNU3H219JBxmvl8daDJt
KcFAgbb6LJwiybSaLUp/RMY/7Xeh7HdYpWGxezdABQzIu+T09BR3qWOWw5yo+CQvVAC03TfqJn+y
234jx+JpSsis8wwF7tgTNCv/u1qhDkR2RAhdlCzb5oYjOGLtg7asFMp5HrrLHQbis1C49JN4rLIC
o5/1Ti7NE7rKXmgGeDJm8xv8lyoYZWumpoKgjNGcfah9Fpgfgx4+rDq53bN5Ku9+gZQSH2OgK148
IM3jvI3rQAar04Xk4BdvWhnwUdSa+tKq4pLPAuT1yMDQFsWruNSSsTuZZr5X6NmRlZKa8UvUlU84
aZW71r5RpuF+s2lx7j1tgeDY7Xx+YGU4jRp/MSu5n7soTur+EI811nW2Oa3Hy4scvdwLg4J6UAV6
Dh0Etbvvph/56YHjti6RitRPyc+6bxH+trNZ+zd0z5nN1NogC+5Ph70QgAjhbPM4U1L3jWSQET4n
z/71GkFDwzFM3vpPQ3wxK872KkBd+vD05CUI2sEqjqZEzYA94/vxVX3Wg45R01AMXKgNeG0ME20M
TFbgbWL9ODuHnOn0P6SMy8Jw4R5XevYvjBmm7oNOa5IrNrUWPeZy77HwaFa8ly8Lvhi/QSnb95ZR
3rSx/30uvGXdwozjxcI8dV8N9Y1zTSD2M8ZjKQOKSqV+SbKNIz/EzVU5Qet1BQqmEGjUuTkI+MR6
xIzBlz0HMw1C8rg+b9+BEWKgJq60ksZAhJc225/Pw86GTBjQzCvsjQl2v3WjDU6IeonLrbk6mUTS
VUWTHvNCRRrm55ejzzu5GX0JFaBYy7FqWxfJov6pOxuNHMv4RwL/8YSCS3LJ185Thz0dBNpudHhw
pWznunab+rGyHjTwOsBaXK5I2jh7qmE6JOhffZg34Zdy1e3P5Zn4pWEcT0BIaTvnHhY0/wt2RvoG
REFNnslK5IxKs5yenMJoQo8tsxX6lbB5uwBXquUEmnjHrmjoJRi0QABmw85o2vOQcjk72wHVPDTf
HDjhHxGA0uJl13MWPuM5oITKMei6kFAq6h01rti93q2DUiWXlluL7tnp49cnFf4oe2gAgfeyxT0n
n3kaL6AqWzJIRtyswzuQXlMTT0bmQAz1mIsPckpPKV9PYdSmkDm8+K6q1dGXy02aN9guGkIl4yZd
pyTYCfWYMI4y8tOhJ+obOfXBns3mRu/RQZAZskoYr/38dEs+Ews3UGPIGCsfTe93i9YVKy3DvW2v
w6Z6U2G9OdJwe2VJktk6T+KjRTxclhWSY44DWIj/147dMiUDONqvGC/b5GG1s6VR5t4vy5xyKaum
m0Jwmk2xpktoCZmSZlLdvE1B8ZA0fSEccpVSSPAMto4al/rbGOD6b5Cm08C+le4V0w8V5SlorZB/
K1KbGBIR6HujexkqsO/buHZ230bk+NfI3IuHdHB0Qmuo2GYTKTz+jaUNagbKwJvZkFO+CSB5hhr+
f4GHUqZ8Kil84tSB/NRGCxjPhwB0PjbuhbosqvcMoG7eLCuzKFsjsn0F4pmrrrbkM1zZxaOqYm1U
nqJ0COXee+KMDKgw4qkW8i9vhPVxzme8DRHH0Ft62LqknmgmdRIkEz58TsXu2K0oaJRVemkYZtLl
ZYxDgQ1ueQCPrw9vfUhkysv4pykStvffxwbpJjfZ8GpQmmB2uDP6HJqEKyytxHG5ojSCL6zKpUnL
ZhFuBpqDOWk8wv7GHdcXZNpCSFn0eCMNrdOGOEe9gDyESZEmOK7gMwGil/e9+/WY1jZp+kAaV1FW
ckBy+Df//o3wCLTg9APBWQ8X0aUCAjtp5wWe/+LDTYkG/qwCwFp/9C1N6Xgg2WsQ3sRlOlrgpR92
mNbwU5CaP0JzSzkpn/X1dBIRjp8/+aOUZHKLN73VZIgF9r2Q5C6a0L1aUsqa0+ufclp8yHm+f2Rt
a/wT9uKE0Zb0cchedJej7WLGvfNuF/t/jRa5bLph6d2znYqt0KqokmV7HT+7+x2pXT6uapQBMgIe
A4+UtcPmr73RqEw/lxFc8zBkpCCFh0yleCno7qJyDdwgSx0zOXzSko6AxOV8HGZXczzTxzzy74s4
NHQztSgO0BbvGwhF0EFKe57noLAwH/TYrb1gyW2L24P1cibeK8/ZbsnJaPpi8UDSLE0EoFn/ByrA
Msw3m8Ln5J3dkccBePKBEWQ4BzMcDk8+Ck8DiJ22t86ZPCweHgyi5ZlglM2HT584ci1nj6Us9w2t
1wbSF/lWjcuIzN6lSOAczhgUOf5r/q4iSd4N5pljkwQsRE+T0VJgsemoKYxT6rjWNlzXVvOtgq+I
JF7o/2YMY2pWbEal+JEQG0c2rPdQWQnIQ+Ptzk1+Vq5+VhSARR1FiL8jWXSDto4XOHVttviNjP8z
EdzoMMl47qI0HiYQtS/sKRwIyQZKDDl3EIdkU7z6FisxlsX/BzSHoIZ8MI/rFt2glPO2RCFqGl51
O9d1bKswOHeLCKOEWFV3TIqC6fvDQWVdM01Ao96lxtib5795JhFqka5RVEjYnoeogLGeEaF5iQit
buHGrgZgYBb2KHEDMSmk30bqJSfC9ZjJqQX4H3bOrCmJc7xBbKALBIOESBN6ywjPigRm1KcPExNj
D4GIzvvlGQeK1zI9qlmmvBsQJErujuynsMWJI8c7BOMW2JjSbCmZ1TTdBOpj1CWTy8u0D0xxa6JD
xT9k0Ynn0KhtuRrfpQKzvIPDF8q67glCfJKpV5oTXB733ihZxJCsMnTls2/lc9Rn+IDDJHDABMa7
Tpt7FBNNo0Kem7/TGpiSP9rMEUjqnBAugQrlWHNS1cLOUnyloqqzzCbgfnMIzMBw6EFOvmiOqtti
DuY+Q9aBHirtthUPjUv0mehj+l4d++jibHj+OjO5uOYsxIJasI837BfvULJEVvbmK+zRDI9M/N3t
7CAMNqZUXfayP0IjCn1kSC7BmY+rX75zcHca38OG4VrFqyQQ2Y0fkOods8RFWQ2FFaoPA0lCvOqb
/7YT6FQnJ4kevQbr6U50nH1E5wA2gYm2jtetEipszL8SNBY2RUZScusQ4JMwzMvrnLhlH5udLQNq
Et6T+jXXUjU4VmzySWidriaYAIWV8FXuOLodb5KDNFYAcSX/kLxAgaXQ/DM8WaV+bHm3fxdIH1Pa
py0n5qQ9nIUbB8ZOQ52IuIw82leOZ8EDN5bmOsa+xPUuhLYb2iDOFeFxj3gHUCZTbW/fAd6PyaFC
liBpYwe4rZPOQcDCdZZa3OFnKBCfOdpZN1Up47W2Dgeol/Fh9RrqtP3w0Ad/YBnwCJ6OUlGePPAQ
pIenOPXJd+7q5YU89a4LRoi9wkOx6QP1+OzGCBz/AeEJYmhC50pi1RGQbXmruC5yIwciD3sWjzxG
RSIDL5KgRnEJmczVOIBtY+UlyAVNNsMUO8A1udvHc4YnTKaqcfvEkFHC/Mv3Ehk+hQbiPgv0968d
r2Xr5Vbi5C+Dto/L7f66o6CZOA+Q274qvptukWJSW/JHNqFd9OX1SKNM1/uSC1Td0UeCiE4etn1z
cyCN3uLvG9B0jh8EOpe+gW9YIR6P9yhC92MlaX8htoog7IaN2K0poYumnTZK9ugovnVaR7eaCYP1
+d911kfaSiYImbs95vHIhSXCWuhQaTJEXbaSUdS0kxCubzW0tjj5ebQJdN/2CvyZsWj/q2hYF2oB
sLLaONvmFRbDhFrO2Xh1lT35f/qgclL1QsRHNBShJRzjo8y1lWY5pXxc0BclGaD5+vycCaJBJDml
bheLLvYLQgcDegHVLdbu11284CMb8c8PL+CvnJ7eP2Uf/4remVeBYsvO4Se4IcdU3aeMSGhTfD5+
PxZZsZmrKujxQqVXeJWFwwpXGk1HrkEI+KgrYagkSOZ/gGzMUgnxLTXC6Pfb8st8bPzEPbNbOEHe
FJLKjLFPD/3v6ZNPMD3pdfnxga8yjcoKe8GIy9HBB+Z0+EfiNZHHgIK9rq1tQG3CxuJQQOnLhldg
kL+J6FzcMl73Ex/A04+NuQv9qIpUmU15/tCILuBHOhikxlLf9n8rQ4356NkkWFTrTzppk6QXLvUe
cM8geneBMiCuqnsUh5+XLEQpAJCJHxuVrF6cm5n+8aUNwpv9XWbvQmxHPFHHrzeU5gF1Z8xEAiT2
f3gkHlYBCEpBUWU+UrmGHZLgSEbTUjdWmhROlCM+xqsgB2ZhToWPYqi/2bQDqztzZjxviobU83iw
zzIGJbm7gLJmveTGjnVaRfddEGb6NnWsz9aWGV8tT0upTHN4KZkB5GworekfE1ymFRP4LhbWIrS1
JerA7/Cs8fpjdojPClrTb/vYk0gfIhdFWt8iXznZX7mHJSi/xbBQIsS45LVzGzuGkSScUqy0rMCf
VbZNbd0vwqwMxntotk+aqdtcn3VtmuOlvNd4Z6ZK8BECTzVTHr8kke+Kpb+B46ibfBZudLpNvvwD
nIDMMmZGUqOQSa+le4THbzO/9hMG/bOQ6XgCKS9fP1TzN+IdmdGMrTWM6D+U9og/C7NnQGgiDT3Q
Wn4yMKZpMKZR/eDtGasSmwFVM9rDPrqbD/PmGnkC6GniHwGRM1sv8GA4HPmWwL21Pm0uf4g0+u4Y
3iP7sHQvfG340lfLUoDHu07ABlYAFH+kZJCi5WLHnfzJTglvPWGBeXd3pVX+PMWc5KwluijtSIBq
IYzIssoGNUg7iyI3QwyVgwtgGk1JSY75tPUGdUnF4STn3tvEF2VCTc/WSTIPLlIRWJqUzbGKEUte
4mql3Ir9yLeHByGNpRMsAjzgxzMCEu4aJcxEgBrGBI9/RmYkvJNbtQ+ZNGMSRVyOxgaGeBXXOC58
JgunHE0QJowxHrOGoFD+M4L+LMdavzH8f1a5zvj2kr9XSud/BXWeJk8KThgCh6MPz2/3mK4nF1lK
9G/oKQJdG1uVuOvcKVDuY5x3ffqa2HUJRvJ0cmbi2ugtWO/SF/1d96K4Qb6ct8eDhniFMOxzsYty
hlEp6MGiVDpWlheRcAfQh2XMKGCI8dg1PBAChn68VgGHkPiMVsAP6PYy4A1lHwdqcK8OgSprBcD1
9Wtw48mjPvUC/4mqS5lLQmmtdOZXdbX/X5AlsQwhT88UfcaSTZbdanuuDM6I3OBC1q0SVJ76zKAW
sadbgXKuEMvtNx2sLP+LQ3k2gDRB8/XLbHDLEwrqOrPyP1nbRQsyQmE5X1Rzyr3Lls5/OW1gJDnD
OLqqf62kTbtScfYV3ybH1Hn/6W1jkV8e3Aj5u10dvE6F3SVEjQJFrNS6LJhyoLKvWVfS+Pm3QXzt
El+PIOjDcp48kp1ZOELfHyX3PWTvZB0WyxWMAwLgmPeQSML593phdiCK+0Grx53FXaUH+GHN5TwX
DypvOTPKMyILNsReHvwI5JNrlMqkpDTRS4kD1iyM8lDDysu1WBgwXQbTkUq7OaUDlw5REMtfLude
jXXddw7UmaIvSEPFdKMLG9FXnK0wO6FIuwrVcvMfsfrIhscWXfo7f0HBpgRjR+Hyi4eit/moTqav
nQ5uHGQ6YiK7ZuYChJ1iZ2PZLJnCCWUqGoJ+lYLDgzSxQ8P5XgywYj7l8RT4GDDo8LlpVCcvXU6s
EDnx0MSoq4hY7AMWCQyFWMugq6c2+xvEAAGSB/68P0vGDL/2Lb3edrYG5H8zrRDwwvymPUND2ffv
uA+Kzv4nKl4vlY8o79HmTGGYR3wlNkpPoTn441GM2QPBMHHO3a0gjO59OamGMzzKvMfeeCO77a60
IEAZKpsikdAUn7JSHN8jNJoHkBlTsnclcsUwsCAFwM14W6+mnZYGUv5G1xeBHnFvmAlYCE8Y0Asr
ht9GHDZ83Gb4a3xE1mu4pLpqX+lCzxJwadQWHjps7QHEhFsd8J5sjyg3kf8OX/euHFx6k0Svr4kb
QP/Mul2G4TOhLWoxdkTrNHXv6YR5TjZrzaeHE6699w0h9QCkB4/Y9qttCMZxF59439Qyj61+c2o2
boMW8FWocksF6Pzn/wMkTVM4quT95uiFz+dch2jFsYo7jB8nGHA9LIlXov9uxeOBHiIijd23S06L
x+pOi0rJ44mzTClf4isfnULtrTDqme+CxEzaHcnv0sXTbgl8OeYrmntOCo1Kg6V1+t/Gdl6wc3Gh
tC14UOXKAQTk4vGvwwTIqWHf1SryygXeQDwkYDZRQEW/peXHOY/9dqJpkUzwV7C5jKZVuGmM+nAN
X3qr2A7TRBuXV8ifZKoZYnYqZmVVeeMmjp+tSerAIsrlV5lG93jbz+dSlVGTUaMwIZ9r4eeq/Tut
sJAPWHW6MwfKKapXf1ytcE9iFkeCz0FU0LEX1+4uA9EwhtFbkF9Sk5H3VKkvmuwq8w0hDKlKyokk
qNAkQJPlV8d6cnlDxLw+4JzihG89AZR6eOuyVrydnGVBPOq04hGew9CoH97Gq7RS/g1PVejuglD9
LIgXj5AktzsGDUudJrS/8WY/NCrlwORknEKtFl7cAWlw9LqQWN/iY9kIj0OLTXEmRfaH2vB6CaN/
bZZVR3CZyReW/3Gob0aDsKGhXLU3t+T6MIEkSKacj1xyFsn5TcCd7uTBYUfhTaXdqNaWMn0dIuri
5Ial8VVMfUX3RkNXRkiTawkJkjx0QqYRnrtp4ZdL0nQDgri9WtWEi9BOKgeAnwVdyWQXCbzcnadV
zhex6MGNZ48QLAP+scf0uPiZIMhcnEuhadYCGKSW0FI1TtBmJ2VfevnI8m/PaaO5kVoG7coeRqDp
LSpRfzpEvmvy8EAJGTvkDU+LcRRPCputS3yu86Jpyc+nNVAwHcx7l5tpJ1vBGTwNODgg9S9pNe8D
71tzhaPhyLEnspAstSwq8rNDj+cSWQ1YH010GjLg6oTpreGgwh0csPlg7W5Sk+j1H2wqndOmtURS
nLvC0uPcLT696Gqn/auIBXN3pXSgG9ywO2x+ZvSXItIgSe5AupaPDrXH7YRJtChEBsJhjLP8k595
iJCF2qyh/xobp3lC/3e+02NYVQpyayLexsfiCOHeC0cihAaqNQYLwZqKAnC/yCdUWmn13UaqdbLM
1Y5NptvBTdF8javvSmlpgdjsc2IYaTSQcvfs+tjvguyFsPUjyYKwjiR6FAn53AkGQ0+CpWB2JrfE
CcX0b0Lz7dpBXyRjgWo+bqZKqvs++1WoYMUKonUL2IaJvEXazvXwggK1f2eAOyTG5bojqSDCHrus
5QaguNpHd00Nol3U4pcgVAvS4Abp60j1rqZWBTuY5ZRp7e8tvwCRsqJk5Nl2MILbHDoQuVDgNl4h
gmtNHSI/+VtxiFSrxleWUf2bGiWFfOM5yzyxCGmvuZNFbGy6yFLsPd0Dnvoqd7k39cxibmxIbMWI
ahoarjxejVBqi2mvD/gIlh9RV2flvtdC4AdraJqloBfry7d6BGiYJVyijW23DzXa3juzxt+87Ocj
xhB12zJJrbCVjcN5TRrtnKnas+cFSSn6jTVn6YZQeUWyozZBRQwpt/IZ2QjKOr82XB2krZ+VeK/U
C8i0yhSDoH6NL22ZhEOCCKVHeb+2+A/ZSi9jEHtDsGo77cTvtwGu17E84CPI2M230VwV1j+Qg1n7
iwebHkwTa0wtL2nlld/yfvL3GYuM/2HTEdFAQdt6YumsKKrmxj291HZrDKQQYTTDQ/KkY0tvMz0v
5tF8fN9gHkqEU4310pZABo5EPeAahGs5wVu7ixCyAAMZ3dt5oP89UauAlq9lpSTh4x42+DHejZD7
z17suGQEXhVc2Hjn6eptbl/gal5bRNhq+Zg+Hb6eau8tE8CJP76OBxqRuKCSm5s8KB7ba+ZXnAkv
7L21TV4BnenxDC7FnbzMQq3SJZStgre0D2ILtA+WDnT2Z3fpWJQD4oHV57sFHU5JEktXsBwmfFzt
f3T3DpaFNbgGXWX86Rlcj/2xGaAmTdwHUUl0ve7TtYXckA3aK0atXBUvpGHXsHcXlpxsLAuUji/d
TQh/EFSlyOJH2tdNEM1D+jsGRbpxW63m86owby4eRHWbU3DYxj3erWd/W9gIgG+/mUxrCKCFL8Dq
d1qy2sNDVRlki+Rhhs9LwSzTwLFzEJ8Ajn3KA/05mrtK8rrCEloq4uKN4MT7RQVOvMhLIpo00dPz
p+Pofo5adLtLlAi9JGZjqb6LRP5ot78FMH7H/622EdSCEgpI3TrKOQEfon9b9pZnl8c7lDF0t3Mv
l2GSO7crZvkY/CeeAmU98/3cEd+pQ1D3Gylw6+5Ayc0mAYYMxIiIeDH8rIquupRnljBWBbOe+ggk
z9Ac7nQ5yWk2j17oNUBwVcR2MnYbcgVlB1/27VBgvj1FSaXmmdrSzKF97rzgDi4lLYxYV7c6iX9g
i3qLK7cIGGvd8uLC3R/rNjTHu1Z31ciZe2QAUIEUOCzAMYbwf/GdGOOsncZPHO335q+enqdi4wVX
ugPHG7Ti09hTHVUX6yFXuA5jHufiYSz41lqhWqJbGTZoM7PMGOcUeEkhLcVfWkl21xL1AwATESjC
x4NVDzevyjErj4hRuvYQRnC4a0HJyew/HXwtsYe8eaxHRUpfCb9hNJRPk3H1Z1crmrOj0xPW+Ig/
axy3ZCpxdY63zpZ+ex10qkgYrxHuTNoxfwe+JpLTT1u7cSAkQ61ykl286yTsSscN9gk7d3zknFE+
Yi2WDq7muv1LMrn8UNjH7OdVHx+0lRBHzbhyRO8rDYusWZyRPuhNgFKWdEqzyYVzjDZFnlbDwBZZ
JLlbukPN72izckNjqbfLoyxUvkZKnSMpC+fP9VtVL08lccVCOW5ctsqB1LIxOwKhTRoenQF9s1fL
FZFeVNSMQvcWhzxGHqh9TRA+5PYXCEL84cxQLQpGJKZuKqG3b378Fw3DXImVn7K+5kDwStvPRh8F
JmXzfCxv3KzDWMN2GLD7c3S/n3p7r4TNbboiZsTTHr1B4DG5XUZmrXEPngeGUv8jNrZX9KK73dAx
LmUAoZ0sRu2dKTTI7F/oevm2qPXixZp8Q6aqoFKrHPizv8i2OE/0JAd5RD4IYa8ePS1798NW20xi
bBIt9Ro/5irNGCSq7/Zs47kbi5j9BGtmhAlxQtx27xvHvsGC0wrbg9G1FHv9F473WmlzP2ZAUjjj
VAuLcQ8mIGcnfb3In+Ea27V5EzB0I8UKa957HIJhx+4tvE0OJB8Q3XowtkX9Y4lwHg2BtuXEsC0z
27nCSKEHS/lxWkBihbOnpl5h+Uyvp6IFLWEJteWJDKQ+Vk31SIyfge+kjImC5vJYr6CrOUreRMpa
RHFfk+HDz/qsR8gKrm82CRde/ahR+A7R/CgroQXJtWIJ7v08D3uQfhE2YI+XvmJI0qaxAZGfD032
WIzxJuNVKnRAxd83bzZG6cpxc7HV337iRg2CarcCl7c6JGxeoB8S8wu4I3ZE9RhF5DRMdghz+Nau
8n+pJiWdym2jVtY19A9RJs18rGdEtMNnCmKPR0OWbiTmbCc/iEwPeCDdc3Rx/mixkLGzKLmb04/R
YeQQXWgUaIFAHQ3YU7a6DcWCiLXQw2AsuQ11atIU0zav2KmIgVP95Dap0PowlXnjXUogfqXdvLyK
Ky9v1VbpoAMQoVJvD44/jPBtVmWELvuR9nM1jQGQFFykrTO02TkMj2SaNTZtUY4PzWm+yKqbye0Q
Qa2uTSGg+lW/XOgHzdKche79IAjmTXjM290UA7cRiHJrRgRjXnuCQNyyLDo8eH8mIzFo1b8BjTn/
SphrJD2+0901SXL8cTfdcfNEkQzAq0CC4qWLaJ0zEt5wfiaJAJfYxjAk15SL5DNIOV2Q27u2Vs1i
0Z+QU6OC48h9+2cxhcIMin2RkcUECKXdkl6YoxBUgZIquBlr7ndhgQbobV6SeaQPz5ObmTT/oC76
STOlVRAK0OBIYHoQ+TcjPP72Das2GiIZjNBYmliTDvreY5omHxCHt2ImYM7WslOJ6TILgnSiPS1C
rFoL3WHmnC7wS9gMe6EvgsNtD8VoK95xK1ljMv76WxxnwEjRFwNgz9bmE5eRL9pNxLIz+GEUFA6G
LPRENDvJpURuydIKQ9B9AkD7t2ryN0ji8nCfbrxjFZj2vH5iKQRTVvcEvQofpSVVyJbyQoRAQYjM
FHpx6DMhlV7eCg92nNZv+0CSYgCfsT3HMkwXG1cibyROyjiuDFyy1eGRZkFyPRuu36r5lh+NE4Qw
rSnlpRiKNYApTYoafqdsvpDjM7ePcJNvo7vhO9POCJhnDknsKu+x6oHvnhbl1JiWI2FfW8Q4QT+h
LsUwY4ly3egD9sP/EU6TeMgbgDbKtVYyOR/Dx006Zef+vA/qddCtO6vuqbqBxbqtgMVKne046ANl
mvjKNqxt4NTiGo3hEqeUKWhR2fprjyI+nWay8y8c5NI6AdTe4KDA0H/OARXB6qfN4Oo12NGjJ8wt
Uc5AvttJrOyVQOE3+J7/T+D2BC46QvB7CDO2WrAnkMb8gl/tG5iEzsolW2LfShyJAlQNfFLuMIak
QXhMyAwbKAKRphdtSWBS/UwMMcpUz2j+6Dl3xe0ba6yzIBqlA1p4qjKUejeGKs6OuG7cRBdW5MTU
Y+aqGCMRPxAQHrb6WPF+Ylkr+9d4qFb0RazH/OVnjqwEgrWjsnmWEJu65KTrsDmcjDzA7ho+C6II
zwU3ouUJAAer+s/YL927pIp29xxhr+/oJu64TnvANFNdthlTTFIXkqT2blAHVLsEWNO9jVAhneCu
buMCPAMTu1F/mv0lrM5ZzB0BLLp2DzFY+kezCRUAVcaEdYFCdSlPSji+lj2D5M1QNJbEBBQwKBY2
x2xrSAV+lmr9UhYJp/WLeygxXA6lfYgiXdQxvHOkEWDG89pr5BvsYcgk+dP7MQnGqGBZ2RojoD55
8TRSATnP4DNONlLAnvhaUWwiivmWVsjv3DbbxjsdZhN9qiYoyNOirwNPCAiFKsXnh4052XXJWSs6
H5QKlBhzwbZszz58wBpCwVasCQic63OjHgHm/PmeGt5Lq5fYS77E98vrUmhpkTFIawZ1WCHdmy9W
UfMcdPuX7TyppxeVgmjDM8yoU6BUA+/xM/wS5oPt6LDDgE5OvHI7fJ/CeIywPdpIfc9rJsa52al4
wFNO4GBYbcKWh7zNg6LdvtgWMjLsugzJTjecH96ACIHK+En7VP69z0CynSvWIPKkChGt9H6oIu6N
7J/NOe0QJE8Wd2ct/87QVKWfB78ZlZasuDYCELXwVUnb18nfRATVvJr6dyrc0tJbWnM11hqwervm
7XrR5WjAZanw4iKdthjU6QR6CGMSA13Q1Ajbex1qX6VnzeVc5Z9hfNSijWcA74MHEmj3OBe06+L7
jUOq9fB9RDTa4uvW/8bg8jiJ80iqIZ7sxsPsRdBnL4OGIjujENPRu7PHDUnT1rfQ1osPNw4Kws34
Pi+f/tf5P54l9qRU5cbspg75BMPpNGzrSeM2EwZfksFe+volqhwu1bItTI5aC9qF7Vz+GsRJVn+Z
UsEa10XqHa9/pK08qumf5qOcHKmfuF62JmPXqm2Nsy6hbAno3gkbSLyXf3YDeM+O3fnwzaozf84V
05VOyygtfBrgFSg8mEptgI6PMjX6hQNnYRM4Owm7Ar195UXyezBgdOT6MIZTE6RpdrF66iOP6wm2
sa40NruZziinVQgOiRq74mBwVPQTnTgrpGnD8zp/3UDoQgxwMY5XptGmmpjYzcBWyYYFh9mGzgzP
olzwuA4GTYZYdR/KRfsClPsCradf7200nPprh45JGyY/x55t+EQ+10duPOkyTQ+MR457Girdpjm7
93/j6mhH47ifzr+XXb0/iv6lvoxmtB6nagemSlxkT2Ao2QTFKXrIUiFSJvR1Q0e9JY3U2AUMFbAW
o36kMogENzsdW4VpXUlDwd0MoGmAFD/J+Rgqp8AHIUV/Fg14CQHIW7BLqhUNriiDzhVnW2mn0Abo
mHwTzR72xzWww12UMHnrp4OrCKRklBDrMoB1tHtBRnCoFFDlVX3FaKLcBPtgBol+2QfIdsBJOf6z
A4ofDoMWuNO3X8MPkV26po7UTTrcMMKh8y4dzdL6dnBc3FdbVCPtXsmaM+R/BPBCUMFh8alGTS0h
hGMPU2/PRcRqrui3uo5QrTBogfgBZYhJfQlDe86f5BHLEMJGI2kNNkplthYfSK9Iz4f1AioMj0hJ
5b045hbpukRBO/uRgfmqpcoU7noL4gRf09cbSbcvRYKMSePlSbO1P1S46JSaSb1yyip/5V6q8oNe
jr2dVjIjL7yCUiTln7q606G5QnzziOKhI4G18kUYfXGwcbAVthafQ6/DRE79q6Vh0uECccUGaYSe
VnR+vZGJmcLe2P+26aX8vXVc1Oi6CH6z3Nh4OSk7JWfibhaxXmRMsiq3j7PZByUpxbfHQjcrcdPl
CUn/VjjrGq7B1vfsYhe1i+Id2sY7lnqUEPP1GvL41S+jaE+5uiRM3Vr0yjtkpQSz6KZRpaJnwYvP
rqx9eMHCBtZ0lKGjKFPBiR3X5AyY3547F6g/V0metl5URlZhFRAy3OCIFi3w1KIjzS4SN7qevEPa
Ye9gHFInB/uD2VqiSFXAeusvG7huqLB7+UUSeRp1wFUm8E0se0L5PHm4dGMCL1JMmufeOUuxo6q9
6v+b1R/QlG8PEDVAuy9Xr2b4PJqSErHI82xEr7EhFhbuhOZnxRpwum+4ukJdZ8gcoLMJu9i86wAo
4KkVi1XVFS1Qcfy5+Mk+uxROdhpL9MgZmuAZ4xJ/Mz9p0REoXTmepUPK9FE8G+wVzGEnS/Y70o/2
pTAGzeTTiuX88ZEiDmc5WZp3Wh6WNuKCBOIZzXEKwBwXvxW9e6cyyKitnaf+DgubsDY4wWWHkRUT
z53aWXOj0Z1afFuJGNKyTadtF8N9e7HxKSRXKiZptHLy+geINPg/sAHaPHKWm4/wSQkgn1oIDdhY
S/W1+WBk7q7dMBGl4uq+kPAkfUEnVzGlKrNo+lqRqGoMt8817E0/cCnox4O1u3MzT3ja6kjbdZha
GPqZmv8365VmWLbZRJHLE39cRgUEaAqlDErUC2y4/Xm7t1PpwrxVBLQPYzzQpoEazAt0lkGtz4k4
Kat0xIbihxY+UQINls7rRDhqzfN03THyTYqDtekByzM5BkSSrxwvl3HkmG1mDks36AuEA+VRVHNk
NYcWWfo9HNjp32r1tAWtw4hPkCUdlaknKzGKn/v8Bvz/8aTFv1Dal9T7GIpmHeV2ja/cP6Gibntd
aKsaJGqeKgy0f9aIyR4svP9RhfaVPHWYNNrFFTHQYv6O1Ugu8maTtQ3s6/60qiGymeKJgcurKWLH
GLUgDyQJ3RvSN57KMBjMd1Ck2V3GK05YfLbdcJVJ6LQIZBaCJGlw6YZ24Hj1JklMxjSNhF/IQK7v
ZzQkOU9YWM4+kdQDZXnnE1FMgwqv+utt2vzI4COPvra4S+xpbaniPgCjDeRFlyAAr5dWZfR2eJHf
g1+7pPgM9SFnJiqEc3aVbl8ogKWtAKgiMV43KzhJenW/cq1xCaquUM4JnpE8vJys6ix/4PdRqRq7
fftmQb1zGtdz2U3xMGoZJZ/Shx0SU8y+vg7OEFLXTC2MA10ZeHtjzLVXcQM3XOxGN0ABPF5F1zhx
+4yeBAzot12gkcT4KFc912H/fxH2ijbyrflNUT15Ff/gQR/ixDb0GLD7H9gg44RjUICY2uMzoNnj
PA4mh4kO2x5Q9p82oLpjDYfjjv1HhluX3nt3O4TkxdisuZAXAl6wFY8W8QEOwklSsoVto8+eAZVO
nouH7TJVA3YbuHB8eTSAMTI/PFOkxtDkjx0lXpHJm36Y7MOqJ4tID66UoMOUJ8jZZje+mg2MZIGR
gB9B/k0YCZIKvtL22nrRTOA10SFJ1VeyQ3e1z08MvEcQQTD83UDYuZ+AteOZtuTEJFrFaBiv6PCf
TCxY7vMS2i4W1yuL/+FF+4Rg+pF52aCsadFO5tH33ZwvJzRb1Y5fUj1HwiRH7PjFBzM/PPH36LF+
wLMaAC9WG83GI7TceKbXbQiuy5KUdJziasdadqoErGbHrEUZd8LxKkourDt+jyqnRIBwHsYJnjcQ
5vHixtRrv+UIEwh+MKhKRZyc7jzW0/5EBScCbT59gGa6y6ydQkjXVh9FefsNRk1nRek8RLypOxO8
QNRcw0g3c+R+X96mQ4glxK9idq+ONnPfF0Y9aLq5+VPWaI3Sho4W0O1NnRG7O5dp9VNYQs2YqyM1
WpGefgrOWLuEETqMVjFT48MnaFZL9CMrqjPyWaw9moQgqTnGHOnrx2r+/nLG+sNGjWiSObQJbsmR
KmblS2K42fLwuZyn24xQ21QzXTdA3BvML3ccs86hngatSBfSXGnHQc+OrJ2PUR/k1vRZ3hqVU7sC
wjt3KYTJBuIy3NQmhfP1BXCiFw5Gy/CZxPSUZU0ptPWMeO7X4dmrm1THZDZRlAG/KU/CL7+4Ms7H
VdTfbgucWYx8Ghrlm9YgrY2p6M0dnT4i4wryQmKC03hLv4DEaXwolPm9OmRKxWxHvfMBtw398DZT
humrC3QfLgfbeCETkFOFyZLKrMb3h+XVZXI5ug6PFLqDZfWyVNoEhEe2iHgvgNCZosdFBcEJRrLP
RRCVmpTDQW2Tfpwku0IydxE5VnBB9uLWdic8L4udSVgpCYbmLj183L3cSZY1l7A59ZduuV6WYF+G
ElbZ20TGvTn/Yt9LBqTVKFJ/U0Ag3Dzs7t22K8CzfMs9AJimOvf7fvTCPozpT40gDmsduavsE7NQ
DVFuUO0U3ioJ0fUkAyhI2O5wvYaK6Upp6HlJ0yT5dRbU3aL/QY1f9kwpS6vtRBzr9Yu0hb7o9y52
DICFvbp94theUD4BU3093VCaKhe9L0fxvgKoTpfDAJVklNccDcni2xcO6oLMP6G2UrVH7tIdiFmE
OoGEBLs7NAWEru497aKCxfLORovr9QishukGpEfvX248Q4lhAF1+ywkR04RCfsjMJZTQ8TFWitgL
7lZ82GO9Nk64GK5FzqYfUXmGHVO5D0GG2FYC22taUqaYPP0mim5dPrIYLcbsdvQ+/1MjoEBLbB+f
9daSr5JvWQcqXExpA4VGqY2vX/dHQVT04xepkqCvBHBiSg7FU+mYbk0nDwKY9RORJr8mbX/fINvL
MTDAvjVG3ShZ26iFWRPc5b3dM4tr2/+tgkzkcrOJPZHpr5E/BIZZbM+PeMb4IDOhPapacr1Qja7u
aunCs0W97enRUIrYOVjBN7tb4qeqQKdepGw5U2SzGAKmOKFr6h5TFA8PbgIgvwMRpVXX5NaAxSyW
8DIo0AnX/euqDq/GK9ZKPgji9GI2lYOjwBsd96hYdwBjWQafcuquCIMTMAgmcQRObmfN+BLawpPf
pL3X8oDbbUYkjKf73jhDNXEaCBL4MnCCAkLpRwDVZ3B4a3kEDGiYAFEn3pYb1KuSA2mQaqc+ZvR6
1wRi50mkaOFncnnlxb9lBWvOuuxx+4MFbUrT+0LoRn/qiO7MczLrCeRvcT3Wlq57jYdpNeK9LxCS
bOsmxdXrIuzGf9GA6ucxp9jEtwAAezWNhX9j9x0mpNuOinAM+ZzY/8mfjA+JoEScA7GvFEHH0VUr
Pxo/piqU+Eao2iw+xFa0Be+RYIZ6dMQXYgpvfQh62NHnUA34bdA1PuPG2x949QNG3MtLBjwoA3fY
p9+GSdS18t1jp3zdAc4Q+NTDGNfKIZYH8R6zNxsyi1rcHd3NaT/nwbbvjLMqCkIfnekYSk+9AJmO
+nl+eMycvdUjFZcktGFXoQF7MF3DGY1bLulkiofIyk5csLxT3Fp0KAIejmWAK8XBVrFBej7EV4hQ
vK15w+E9sYJONv7TlMA8aAYPuixRGv5mHChcG0ssl4Hah379TP4UZhdDJikfnqEoLdSPKx1ZHrWk
ef1ymbR2NcxF4TQA6bh2p+HAYfCPbn/75d3/XV4lJBNu014m08nQ2S8iw5Ir9qklRVczZDsBbyIT
T44vJz1RGZk+KFLWMRsf4uZH1PPbdOhXaPqguF0QqKbMYGcPO0Gc53QVJ9euPRrlj4ZKzNyVhMxD
8e83TFe1GZsLwhkyg2bS0GIiUHWE2sSJWtFUTnBhowINQZitgVzIrEPXSFvLV+PpbaptgsTnsZOv
ex5zAwfzAKxUU+gYSJJGXo2c7GhL6LJ4ImzFxMxkWzDWT/VaGmvd0CZsQWjkFk4lSxl7t3z29fxv
Su5qFCfhSiXGFiZ+JOTS4rXKzRkHqIO8ABLtECmiDNBgKwJ4labQ8lEJQ/lF0wKlCa8EcdbjxtuL
sL2OWE3oSvhwJaxA2DS6rAhXTFpgtX7mAl5UYiknWNRpTBRXwzoVYf+/qVWKen7z2m1LkPB8Wg8Z
9/IPcRZf2we+KAGh0l4vsmlguWZYWQyT7rMAxvK3jHxGHzYAkjrYhspPu8IHqYKpviTLs5ERkXwI
KRkk+c5Pv51BoUFYnHUdpzfD2euGY9fQjib/vrNCspnx1XE0KlEHW+oY/5V3A0DlnttgsyQlScuy
sEzsCccBMvlanRtDCVwpKonzGpTHpzuKt4VDVCZwOEc19XX4AZqWINRHOQWzbOl6FcffSMeJCUDF
guN5wbAo0TZ0ZOE80ULtsE5Ic05WPxES2j0fIudcyITWaCi/nj4LmY6w9srlWvCV64494XSneAkB
rv7WjcBs7H1BuQhkZZ1TuBCApecxIGguQ5p/VzrMQ0sppPnbeb2Ft2krLPCSYILQIFKQnrQK1IP0
rsjijUKrazziaPt3EEx+3TICpKyHbwI4vWhZNGKYNa9n+dR6ldPtS6HyQfJkvUWzV8tKrXo8CgIl
83din/myfsEKQCedTe4ejGs9S+OE5wpIff6B3+SP4RHz3IscIMssrnNN2RJ0VQbtOYyPQmuQmAN2
pw+DntxxgiRzj8QnlS+4xCXWMxbBMHzImhFXHh5E6ozC6x7qjfdcPwsYxyMqlN9g1IyH+AJory5h
Qlmrd2Ow/eNbSZ7PQ2wE94oSmBmCZmUiHuo0KE0bp5tsEN5j3ErFWoDowf7Rn615KOE8dAlkzBpm
d6M7m6uxelgFpJLkZCIcP8hfw6ScVgCEo7FxhGNQIPQKsc8fouwajfLkgTtVwS3rJ283FGXKKuEn
sxR45V3Y0lPb5mdIw2LtbzALH3Xzq3jD2ArtOzf+NiXa76G7lk/6UyXykEpRyw7TYkeGEezLF/6Q
lV2QAFImglUAI45fxJGXtmj86PRDennXOmYdnBk8+ORvc8OKQDZeZRajhD3eJw0+kd7CUfxvJsPB
15mRR6yq9g6qgj5CAjBqUpQS/4Bu/hGihE1WGcScZ0a0WLmUX669fP0ggtvWmRmDfB8oYw6QpMjD
5ST8dFwqq8A54GQLnJgTK5N90wxTWxM/Mo4DvTZsDUs38XOtJuspKLml/AWcvX3gbwoU5b6Of+HU
e4ofD4avGqKbGJHxi33m/D5e2TeL3rImHfuwPW8WdcabrCgwzhp00OU3HqoZN2G/WlGV4mFovmXP
X1Uk3MUBekEFecLXL5v+FqV+62025lu/KgQ8TiOKB7+wWVnJnjYAgXOh1agv/5yC8oxg4XM0hzEH
0czDvDT0klaa3z9PYSB80GfXKNboVL1Z78UyAQukcuQL6Ch6uGP/tTcRlxfCtW+s2n52iGvAS+Tk
IT7iXHTEHddvtWWJczsEKAiA0iR48FDhGlSpa4IJeLdffxmz+CxOYpqIw+4EB5Bx7YvD8vWU7VwH
zFc8GaJdUKvhxeI4Hu6sFtW8Gbe/NhEF1nFO8NQsK+DF6m8qNe4Fa790BBxcEx6rFYAtXxtmXRCd
JlSWrlhMtil6+wWlrDes+S7h/SMTQP6SEteXouf9cE+KrUWR6afRVBigez185Cx9KkzzU9ti9zMI
LhBo4/7sglhmHAKUZVLGyiF+ly32MwIrI1p+vLjHvLx0lyDTAzltOw7EZjCT4wXv1KzwxftYjSWR
O1IRYx6GewpvxhKZTQGjjlMA7uEs64krwJ2Nk4WdxaFGC+7Vt7kuJP9ds+aprBJFGvBNPax+5rrd
aRVVN1PujQUrHghKUdTxRkUlsCULb+ob3BLnUNi5TDwG28BsbYg9LbQQzE/C9rxoL1OAeofdzsK4
l/Jn77/JAQqRvKcnWRzgK6INrLvolUGdfmkN8V5EEHWEm+B7zzw0qHSbcSHMiruHRxlbvcOXoTEa
wOfJinW/e1q6I+sqkQGwF1u7Pb39MoW5s1cAUiVH/Nv8NsbLFosNEs88JAk2LV2NWztc9qgORkvr
xAfUpYHnoHrH6zyyekBMq4L7fYxRtaUy6j5/F++WjOp/prjqBXv5McorNjBq6hVd/VkiDHTFMz1p
uah+gozVsgH6Bd0tb9YbdPoU6s27IUo36syHQ0XjisNdidRA4Oy6xPFAovLF7ymGICxO/RIoiuqR
ed4Ro21hCI5A6RkEZwMw3+6kbcnxKGsBqtMvHM3RvBDPgJVDfeHWC2fb7O2Ou/rLLH5X+rsfboKy
X/r4CAAsvX+RIpJWBl7XRXgTAO8QRaW2SKfwATPmKkX5R3RDywxFHGiF9yPtIdEcUYlZ/h/uA3no
KoNTpO4KwTFi9XiNFgZwG8Tfxs30h4heHSJOyjBNohIBM4+dOFv3bhQDx1yu6BMrPAU7NwFHDIyG
g5OxINx/Da1D5g986+SN1JgRO4/OyDIlfIaUhMCMpnhhrJkxNxln25ShsvLiEFe/t/EOcZSVJGrp
xr9U/GIO1Pwj1btXjSm1oP3KN9Vk8UbPXDoFrUtzbbRgP8/XjG3F9tXwDhlQTr+r1mxNCOCFFDUd
LwUrlZvEVIRP3r5NGNdFbrw52YA4g+b1hIljjXj0MnOsO4InkNC9zxKECXz9pVzu/6qzBGGklgzG
XAgcA7Q3H82exeEufVj+gksZnPEAUIjDM5V54rsBRMnVcyL4JEi99MuBN4KRtsrbDNOIt9DvClOq
mDk8jGnI5GinyM7LoTIAoRH/Tn5b41NTjCtsSbbMGozuPDlSdbofjLHcPOv/2oEIRWym0Jx/zfx3
44qF0Tk1E274zDtIQGlW9uvRH1wU4xvo3G8NI1K4QmL7teakfDAECTko/OTnbVd/2hyEhthZd9JG
8Uux1OS5eDQTDRzrjKnAsxIWVcFFBuKpqEnpa1g+wd1U59dDoXg1JDh4A3Rhp9yaC+REy/GL/QtX
AHdwFWd7mpetUCRejDmp6Mfg8LlZ8DsF+6GSac8BjUU+8gCAS0VEtHK7SCAYxqf5vRm54H4TvtOa
8VoKUG+DcjtR0JoeL2kAAr/Icqjigb/65W/v5tMmxunmP6LhxH1M4MjeOM8pDyYvG8wl6Z8L/hRV
sXWiXpM17J/SjsgzDbaSlx+kbjlR4Zs5CJm2PS9uxu7eXpnlFoly7sLZltlPA0Kao4h8SxbWX4li
ImfEkGTdVxUqsOMP4yPuV4eBChcnAsPonaF94KVC0TOKTOXbQJ9FJd6LgAeFHerMf846m82l9OEN
a6fV8ctX2Gws2wWpK38cBt6S7sBlVelopbHVO/5MXsxeUtSq6KQ0ry19owJ4jO70Uw9JQ2RjyyUz
VJxz+LaGyB5DC/CuX1XErsgkxQ9Qiw8dMD9x0gHyIhmXCnO4Jp2HUr9EuxEyvbn172b9GIf9lW5z
sjUUmqH4piv82ShPC8sRUbNTF9CkZDaJdZ2cpZJDTB0p/zEf2vdRf6ACY80Uw9Whh0MbQf4MYE1M
87wHhlhT8E5ddqcWoXjJ5aC/jMQ5Z+xpiHSEuV6qFtcpt7K1qs3yELDTV4oQWeN0ngPbchEsxvH0
xY4hpfEPjeLU1xDsrJoOhydmTucgLSsMl7uDJ6AchobBuD0FRd6gK2Pq/Is/uEwKsZ7Cc/LPoauK
Pq6U6RJFFOyiXvSgewWZtPzKvubobISJsWlAQNBbtwJTv283GtD5+nRjUy0LtVxMOYVnRkOG2i2A
ESaj09TAKhn4aPbqZZkJ3fxwQFy2kgoKH/LDzy4noG5u1lGtSSU9GmXkdIYnwIjPnjjVG43Daft6
O0y0Vz2WtBMX6lKG2+S9S44s7H7J3xQDl5PLpJSpn5IA9ttD1veBDcIGh4SIka3af5uJGVCmadyw
c8YycEl2fienq37+1yDfpCFNyqGSp/i4LpOhbfAKRLTKuRoW6zhnNMtJYbjIav7vsQwjDOvgY1Mr
QVuvcF629+7w2mpR+VZgl8RUn83Xx4jbVGoBNrVeC2C5KLgip9v9T0+aZjk5gqL/QNy1HzcSAtWF
1VdsnoZ6+EKLAPkco2tc5SlpsbiP6sMUnV9dU52oDEDEPJJOyMJ/Cp/a3Gzl0MMwb9WjpDxNTsqv
FY6irvvR5deuDh/Y4iop4EqNcJRCVJzCQedSqIEfcKS5kjpsmmZ0uP4pEOh6eH0iU5z2dfTX+FVa
c22BvEP9nnXiLaW6AMU8rq37bg1b8fo8pNCQVMzCqHllMx2lF9e2JfofNmJAgzahmtxsRPGyPFcG
baGQ3pFZDCPXOsKosqRH+EXoQ9Y0vnc7J/F2qGQ8J45uIMKri//pWkj8u5VWAlxZIfNcPEC/Ko4f
GguHONzW/vYWTi9LyOtX/m+eAxCgzXTCknp47gMBTLiavUgIMKQtD76NvR0XaN6U84k4lgtrhxIy
PzkLKOeaIlFRodmsIK81Xy+Tvd1VRmnd4wkERfjmMvn2aLvW+ygN36g2BpGBs3cwPtok/7NM//6b
ebv0QzYQq+WwE7rWKSzJP/zRn1YeD8pSW58/IEMd0jpn45M8yEoCLF/R8hv4Q5G1QpY1NcHnwh/h
wWQ0r8vIWA68F7FXJUwWRB/QwBfnv44akIzfkJcZr36E6LKJbIb16y+uL7dLWiaA6HtdGbWnC//l
ruFSEq9Yve85LLeTCgq6Cax1JPERHyXmn2V270Xsip3VuczbUk5WYkzBXqWbTvB09jKblb84MmAv
B3hUuKO4Gxb+LPmw8LUELmTeUSH2EbsHCzA3PxsnOGcpZzh8lxBh/eTwB7UZsKNzEtOa6TNQRzop
d65zWidKz9QR+rsKCg1gfCNRT6H/3bNEBQR/wtwskIVyhA3IaTSEelVo/egZy5OYke2+lq47RVJR
Qmw3zd5BaiT+eUotJZxzj72d5c4hn2rBaTdHGKK6eAJZoLBHO9zHHZA0Cy1TmF2BHBQuxto1rQbg
o6MwQpz11TxhLmuwKo6tmFrXddFGrpqOlw6741LWTw0Sene/f0oy7kgc/cNwugSY5GCc5RmePYyG
w+Zz/pwFBv4EQGZgkPk9uHCWbhBV3kRms45qzlZ6807rUvaSLl0B2b9gHfB9MhTb2yKCXTUf3h/E
I7qmQ1yC6GwpLGPUdneqIGiY4UhbYc24MbGx9rkcksJf/Bl+3xSksDiTgTakz1Phk6AGHd8GnDVv
4Sv1XMMGbbBTQNZeENbOWfQb9EVY936kvZg9gWQNKY197EIdOJPtaXxwqxCaiX/AdD5Plk/owswS
CFGLntzBjMr6vZ6DGJc+yirbvRiUbnEIqAlSV7rZsA+8lS2q9+wowwIhqAa1UNFlOJQGOOIhm+a7
/ioVqwDBB1O+3R9ZR2srGB7bwK0jLD81NJOuzRB2fuFG2AwN5Rc0B1teFSnLTd31WFhBfX69MDPT
jlbNK+zj2xqfV6rTc3Zrkuj6/YNVZRtibEtvcfl71S29wOlfBshQ6urHHwBrV0QjQR9B1RLtd6ee
jOw6/MtHqgnanhexN5KzmX5tm0DhdruIcp/ujLEULHjQoocYaXlASSlE+/2U+8fWxoKgnYZSlj0b
sT0HXsMFmSeicCiR1egL7IrttqqBKxrRtY8bj8WrpgFSBk823Oks8ZCulxtqlcwYBx6Y+RMr2F72
p6Y8MMa55u0knQhJwLecRWVdjbUgfnXf1BGkggdRP0DIRU3Ar/X45170o0YKuFAtlvmZgJsdkFUc
6lHimAhlikPY68KlDEfj6LVoKlvKwHpTPSyEDkGgD5YecSsgSpcOsZDifniRkMfNvmPnsn8/bY0o
DrGUlINsfXWEL9qNms7GlAKy3eMH+hcnueCfqokYMFHTIzZPsPed3aFd9Mb+iqU7i1XeyW3QHx+h
iHwyEjMhTf4E4xo55YtyZ5hji83NlUWrgeQIxWQlOSMyG0UXsup8ukeuPCICHbZkz+zW7omdMSB4
1eKOIGVl/qBuRHpO4+pmJ5cNtI1GUAKxWcKTlQz14VbPaXMOpcpr6IQVcURF16fyPSIHetgBkWl7
bb9i4gHBidS99At6IameDJZByx864Z6fIuXmywVZG3og3YHfjRVJuZNyiuVlm9JF8evk6ZNXDtkA
Cnr2daZh31qqrEe0o4+PuyFF25La6doO4qi2PRZwQn9dL47z73/O+Gtw8URyCv9IMEVHOV8lFrtw
fqUNfWsaGITJK1YoR407545eFZukmQzB94KBPMMtVOlM6cFJRFnb+s3yp4UhpQ4vLfHMN7CRY2Nm
YTJRKBkz9QggEQojKuyTC7So0FaBCgcGWUPqjV/pUIlrhs+B8IivCxtwLdAPS0HbQOa8sKdn4amW
qlRdX/nqp7wVP3hchJpdbpaSJafknJhwa8pDW1jjwEtWzNttlneF1yFtYs//4wWg66WR45iO1sbc
f6SCAfNeOtnd7kHXLKRI8eVyiX5pqd6Vnc1xsGt2vOVTLeBiFneprRN5H2QyxiztMHnhrxwrtz0W
MyitlI2waK8uT163CwyiFxVrMbzTvoOGFkD1uFOP1f8gv8fI/xRVEu5E6vPBAwmm3qWm1NWH5GR/
ZtHSNvuXwrQT7e73qpRylFsckWI7jWbybEd4hIAhSEBoawpPB69XTXLm9s0rBuvpVeVuUvYIw2I2
Tk9ysZxC3kIgLh39TQ+2GxO+SouDCvksC1bi3woAu/+w/8w3MNiw60jlytJjMcp9INWiQ75Dk6sv
X/2chTEZo7Juu/34o5JOND376nwx58cd6dB8wY3UtUFT0AHMu2EGoCSPMubjk2kvwg+dfPy+0D1V
wpgPMsCxNEYaXXIyvQcZBmkz1eoh/YW2UeKin/VTaMPXwpxX9cY6dlpeEzHJxRNjVAKKGm4B36li
/vNHxC5ZafTcyrN26eoOB2rTRaUU800Q2gQUiVBsh4/d5Es7JyDfg6pdwHocw9f+4Z3RYsKgJFTV
rZdQiFEcHfz4vFfj3fsuzcPn2gesr1ovZaT7bBqdsdfytXEuMC5Mjid0gOESAtGKfoQgP5pXPTz9
9IQi+aS0jzHYTGL1EpXxIQoxY+PAof92LmbUIo6GIKBr8qLUuIUOjNpuu6sHCinJ9hEsKEFWTa3h
3NyLReT+J8VK3DhwrwuzNjNddyt2cbQMhVJE3s3a3ohNpS/6OV6OWF/bbqLZebKJm4+V39tj+tXi
eICSFmF7t+2FZb8cp6dO/pcoN0NElV/jlXAjIZgJbCZ/iNNYoYhnRdArPgVbz2/Q253uusv8Rjl2
5mstR42pPmTX5nQRgJDRuDDZKRqDZwHOHZu2pXPi65pV6c0zXYZzvNhWF/uGkR4LYv6PGWClbFqb
qqQOqWLzI8DcCfLk7RsShPAZUEE/svXneUrZP/Dz0N+daje/5fSOfLvFsNrs06fZzSTZIpcy8zGv
nQuHZu6sZi3Hj5tPeu3MniAEJpFk5l/D8E+fyw64Vj9ok3QINideI0NLC2Mg2lxU8eN9Ol2dr4cF
auUugohEySudoWY4mYSpodwNIK5sqS/+jSmVLLJEDoX/7FraGlZCqH3UwA8DhU0+1J4TuvTb6fY6
Rjhct9zv7Xadt9AEjib1TSa3TgCZM1purtpqB4VGeRe7cJo3lvkic4F87wEffbHtocyWBPw0vwID
fsUim5RjQFeD5krJ+yGeirlGDrgcXjeiNY/nRB6YYqAdGX7qJvbZWVyTFkfuXPrPXlg6pT6r3xp5
X/zagFr55JB6cuWsg9GpiFpH/MCi/gcNcXc8sS40T9G4sM9FCrukDxuZeekzs1JnsGPAcx28dBRh
ZDlDmMDlFxoBBZD1Xxqoki8a9MhHgVnq3MQpbfEY7pMNVEgu3Q4zHpGSnBeppqUJzzovUyDjtrYg
mJzKf0pvqL8gu2FX5OM6449h8qFfP4XkL5+LxvAyDJikR5Gpc/jXHVieyV+8BB7Pozz1emw9owYC
xFj/cInPseWdmN+1n/EFDskyQz80w9FR7q2XXcSk2dRHlEoBV6dlMvsoVttWJiHnlwVQcDoYqqWx
cpcjnCQcTjw6xlkYkSaP82TSBW4pQC/v1E+YOwaLtF7jZafEci5pJmiNdBTqMLB6hXUPnQsB3RFr
QgxTI1j92aicsyjBUgrsdOn5JQe60hHhJ2DxL4I5is2xght4to1brh6bzFoF4rLguhF1zN4krPC1
ZVoHSUj3YUhXXBOLS0c5cUpJEYgkfhFgtKTPCWKNJaNARoAbVFR8ng8tevptPb/lj7SWdmscGX8e
HJRfgHUrGZWGOMObaLgeSi4CyWJKbXMPeCYPzmgwwchPVV4mIGhnVY9AjoIhfVJZLPLHdJ76Vw/Q
Ipi0xBMnKGsVsA9NrdNMhGIecQYnACnTsbuu60s6Ta3Kko568wTufROkeYzxUeyQVow590CYlJGi
R/7zZx9xHXECfinteOjXmFyYQamJX5XNcggL5WFLCtxsciIqfWc+yr6PZMhF+KtBKa3jQnPjUw7e
k/uh8pnFgoPKnB1KETNzqO4lJeePZ+jVLS+39dfNzODnQI2LS/jCIKP1sRJk5KrM7MTl67t/kAUP
C6NYTqH7owJc/aIdwoVvXxBsDx/VgrIBH2zJZDesk2LTS29QzYIE01x2SOLCJ7yiixRzFT4K3Ypr
0p1+pgfKd4uKNSmenFaKk6bqTRKZlnThwrY7gt911V0GlqKr2MiMdOBqzYuZWMTUEavGqpaxAibZ
BNcQNTLKEOf5hDVV19bzmmDZTqnWnpyXQAy5aHk4P9lLy0+1UUrz9a/YcVnlB9StbTbps7V5PdDU
KYBewv/coC1f/IVnGEwTbiSMAO19pCyvEvNg4tRb+SUmdfNDK1Bw3Ll6b3g5XL2RbxGBoHncAFdI
KizX4OLwSrTARo7KIRRd1zw/ue2eswfybyI4kg3qKbsOvLt9sPNLl2OfH/coZl9V7CSVp+fIe1kN
RwwJdoR3Us7up8R5iUiI9qPVVrGAbhjUTEVpruH0TxasoW2mSbVpXMXpU57WF/BTsJuVVM5jJIfF
nD0Ei+rQ1l76gwJvr2E/VcCNpPz2LBZDaa5wfFG4cbo/K4+a8ZIXN22kE3cETqhHhJD17OMmEecy
LlDw4Z9wu9Mq8f8H8zIcGfee6H58PttjrvbWxenaphXDwocNE4B/Cuyxgb+PVmRTOtzzmrShh4my
a6hSPJlhK4xttQF9mjTQ1QSZJU9GdeAWlVr4xuTOipXNvrhB09NbB8+kFEZ3oLf8+Kl9oRVh06wL
5yP0UZLBBo1FTU3iabHy0293g5/NCusYAqpadzD3vxr16nOEBo09ptRO2wQ2WjgKZ/GjqzaKb/5c
ub0MMoLLrnRr67/cxUvgT28MP2CKAy6r7RUsl5dUCyWa9G1ks4cUD3AYs0LhzxikYr6uCYrITjqf
etColZ5r3GWab0CgnScWaLVDsZtT7JQmbNJ7BtEd/JDpbNkQ56yElHR2OyRRrxRd9T5CPe2HZUR+
arKRMLIWXtKzyMzQq/Ei81ctD8uwhoCZpCOzlv7YENZV/hmmO0qB8ryDoKZsiubhOJHG4h2T8/Qv
Mi2bSLQ4y8pcLjRkdOG6emjUojzAv0tCDheLa3tdjaV/O1IMAfKlKBN6+owWKnv+XQGIBwYNU13a
WHiUq4A1hDAFLcF+7Er3dn+MWNg/RK1/kkQQ2g1CXEPCprbio7Ch6q1kZBnFjVHVMdUbLC28hnKn
jRBet3j8/TjAYT3jKGRaQ1IcQA/DqIiAdKSNwMGvOCfpCbRsl0hS8pAGfPi0hTmY9gVorkkP028L
RIU9jcuOM2767CPUULf3gGXyTLSJSp7JcI+8hz0u5N3usj7c+6a3xHGNy6KngorSACnyk4gcdbkV
+xmEO2sJpcF9VD+t54t8qTedoqoAVkIUvBLRu5KEps0Bn6Ga1NexJL880VMWzVHU3Qc/rVXtU9kf
eoqvJzWTuO59X1PPgblY3sHWOGa3wItISoA/aSiBCCzVlYuLnfrTtEHHRsRSKdtQ3XoRkBWXRKbJ
r2z/untB2B1TthnQzUmOLUdRAc6c8RxTEocwgzqUawj9aYX+KRekT4AME6Hm11Hmq8t9MpyKzyHt
l9svIu+9sQfSuBtwnvp1WVtU4J4khbk4KMokvcEytubQhVMbgHxDO/6jPf/+rvdaVfV8OVsVh4Hl
u1skxwRDz4l/8ZGJ2seN5seAdeB9HVQh9F+kO00kboVeBM5BxNhTrqQC9uE0NOkL7xLy+wrUEsgR
5yAnPgXJv9RYH+EVLkInkIgnSf+FhZVjsOkIycZ7xEI9ChDtKz36iNjLa/cvyfDWirvc8+jOWOFp
f2L9vFW6DveQTAzypYAt7UrTwbuJQBBQdMfhPQZx2XODubV+aBnqFRU9w0J+xoectyGRUwe3vETr
ey8fRW0QSmWwTtEQRE+ihVpBMRTeKV2felbD9xAA0VSF/pCHL+xFU0bk5dmg4LfMqEQwFCr7Js3+
7nihQ7sBaaM/UffP08hUJ5nsXoPWIf9tBaxvG+KimjG3GyToQMoJwsrceN5B3eFKUDoqsJ7NV4bu
n0xjULPDgeh2fKYNWZKokT8CaHsca8QfYXbAgEpNpFFeQU+tEbRWb3kaNOPKaV/0Iy+3gEjj+07h
N0kpOuBMCduBDI2ENrsNKgus12sjDwyhir1oG+lpEYieiePUDDq8DBwCvCgUQT9nQyonCnAJNqhF
fvpPlneWwPqiyS/wMrb4Q23Zup4Elmdx7MtzAswFV3NvJC3oJCr7Uj0Bf+15bjBx3kXQjrMySdGc
bgNZZyOmQ/7xcSZOvkZpEd+7hfR8fvb7RcN4R7VtN1tOegE5r3XRwniCmjPAmvIUnjE+jP2QSOht
KqKfI3X2qPgUG9gFIywndWay1R7A7O45iU+1e9aG6JZ+k5DaPMvE9wdzSV63kcaQ699chzNpKwD6
kjjPI0mtOs5Wu7q2jhctKgGNtlq0fu87vIqKURFIvyZP5CixKPBprSj4fzOOLSE7IZ/sghCOrkFA
R3XgsWBNG17vj2YFsNEL+mPQqev8hyNuyrS1n4t8PV4ep1ttQG+Uq1IEuYU5NbsY8tlwmzbfsF/e
XYTBVix9EGJ5XBJCnkVRzU7vOgwbl8qL/zvGFMCAFClLNJuJdKIPKuYPMtxGNsIFYzt1nBu2pKhU
YUYL0bHkERnODMG8EglTchyl0Lxm5BnlUrVRXnkl/RDz5JWbzzu7iN8IOredCIH6hb2Lchk2u45O
cKLuniTEERicDOVZfgYY7+HgKWMxD1ZTb+1nKA6D3u248qyKFFfJA1af0vqwkM9JfkwyNHYr8Dah
wU3xYblWaNJC9zCvBPt1SaJ2GMxzaP01JxWFHtZlvBrzQKTqudfFL3WQmX0jOK3UjBANYGEsWz40
8aj49JvT56kj36DOLyGAlcAyJ++8h1g+KD/9XXrIFhZKdPKJszqkB3rLIZ9UfQUz4y6FsvevA/cP
3yLOe4NHr/d6dCIZ5qV900n6g/9uh5OUs20HFZZC4KrD/9cCUua/Qfx2D5zUyDoOQxL6zHqkthGJ
BtZLHeabQIBWBTM3bJIN+tBUcMRAVOXG1jpq1+kgFG/UAHZjSy3ZJ3HBIej6e38gjXecjG+LTlre
ZREoAXXsq2M8Emr1eDTbR+0sE4y3tkHUEHPp6rosSmx/Z+Cqg/5osuXe32q/WQAyYTQPQkMO1qlf
vrTpyyU3uK5MVixh4BXYYYBYcVrNky23+SqTOpYlWDaBODAu9FXAd+vUDEO/NbNeyyVA8PylawvH
3Cn2rGZFqTvzmqssjNGH8CrjoEqwVpDcNqmjvVN/0tm4ELJ6e9pBMuWsGiyI39rO/RuPlzXqQGXc
Qq5PZeNukUbBFJEQiCElqLcpzwhYglPA/FVTeIvUR4CC0lvXhnAkSnZYXon22iyJjg8HeihUpDzD
jCr8SmNoWbAr7Z9cMguE1aLbQYWsJo2UYK6UE6GnQMfRb76rLdgjA9C/bewfZzJ0JKHZOty6WrVP
CYF42tGL02TlCldzgtX7d8gGlNQCnV6gAAhiJmMrGQbrlVdk03FlI8zLqyL234r/r+2xKgqxL0u6
uM+JgwlhthyPhZ9K0d78INfvc3q0ghtP3zqpqOYaYZ+VLBpcg+H2E/9z9is9IMwcpQxrSeeKxtFb
iwKsItM0OfcIBnVoqi44nRgUNNOxsQsr9+CZpliGyjpfsfzcUHwlileVXZXQCkvu1ESx1wU//ZPZ
rSrwjnoBHoYPemWgyTBFMppFtTOCytdkdAZYtySHKWoZk4+0+6AXCEFJawbk9bB46yoVVApqon6s
pDaScSi+v8Jsb2qJ7K4xDcF0w2ZP0HGVesaCjR1Hgxa57AeWZXbget/KJe9luUzeMvTbdX4jha12
f8kL3kCQobm2rKmolPpKT3DwzEzZhb9ChyONxwd5LMhB4BM34Xzxea2aEC+LBREq1ockXoz6O5b5
hDCwfBUGGvw6LtZ/ItjM4bsBFwt9vp8nz6hpGVdzHSXe3T1/U5SlRKj42u1uxToVPPK4daRsXlX2
hQY8qRJOc3GLBUDRNJNFzMZdLe0hvwCLa4U5xcD8LvXybFQPhzGz0ceDFUsPvXGQmnYHRyhgrB5X
7DW627t65czuf8HcSJo1j7FztPRPXZXoiP6i4lZJNAOe9J9BaMXlN1W3yj1hSlWuaMOL5ttLcGxK
Efy0BSNTb9d5nVe+qqvb5vfwX+si/aEqRtuEtYuvUH3DATgwFCYXztinvZEb1xBPaIqckxwQ0YUG
StmvFBSWmTBQ8nFoSdlMAy1hxVbFGeks6QXpH7g4E9f13Oq4JZEEX5p00XoVvgy8N8S9BXPZgida
EwQ7RH7k2HqHODgynGT9xJQYDasDrPpPvD40cbk+28o8pl8kguOEl6K5f/RwuOmQ9H6Uz4Vtwd53
oscGTrp3hmQS/9hKX6OUgsiTPrTguj3cNF54jVZqyTbPMuqWQZDuvjO5hMvPUT9ijCz8fQqUbh1g
oXaML5qlNZf3YeK67AQM0N6aSihXL3x4hbgvE8ZLc238PUOW7PPK3EMqbxJeXE0CrK74m15dMOTl
5qEdjjCjDy3ZnjzmZihhOdGfys2oYEoyyE+sbQb8/O7hVtVCDI0KbDJMzg4nAnrC82cud3oUQz4w
lxBorh8fMBfmZXmm+7qE91l/GbDk9QKkj6z/AZJWwxESBv9eaDbGgwO8Mxig7lsskQyv/qmCtcrZ
FPIA+5RDtDBnqk/n9mdLO7yJ84xzOYqNNBaR+ioIuWXPd9q9Gc1dQzWA7FTleHswIvEamWGbMY7h
0lDn2R4J1UIY5OodJeuA8Fcj/X2rxpzOnxZLw6SNtfBsx8SRHEErXPKmVaxycKG0zP9FOd/6KlfU
RMyrmwInpeeaENY4KKn8mBkK7rqypXzyXJaiGwFT8g44My6XXAa4dEEzqh56G1LfsyPEWDZghnsF
rJQJolweGa6FU4BOijBUm4Jv1RVLL5It7pgYbpSIEGSHb1iQMUs6msip/ofIaWf7bEt5ysbnT/2n
t0hBScVKebfOOTr9xh3nC7QDFv1GXgYf6wuAuZcHFeoATuP01PqdaTpCKyr6v2n244RszVGgIuvn
M/T1qm3XgYmfzd6UDVMagl5Gq9+aHjAUdonefvrAAZP/nnQQLfZ2TnEiLsTuDKTt8ravZTaCPRJq
+A0PrXbWA1nyvbwywXGvCRz2Pcj02ulQYbH/golyoRqK1H5s69KsZ5v2pCH3f8MeLOOBI255cO8a
FkqbbPCy9CEhWAR6TEV+qO0OGtlFJI2qJroAfHSVbf22CmtE7CFERal4pSgDhyvCxMpV93L2yfdG
8WZWBuZI+C+eA2P1EdIcliP0yWGk9fQ3UB1EyJZc0/0Fs2PNGBDNZR0veuRibt+2UDbRtiTyF6bq
1gMW+eINAbBXyQ/WxOsH6/uOIBzvJOa6eH8UHqvUL0umUnChw7gsIvw4bpVHecPfyYVQs0dJQwlv
xRVSBTJItk8cgdOvMe7QtwvaioFpu9F2se0C59yqjQz82P+gKmA5FcRKQL9zhygrR0O+YwI3C2lF
gMC97ciKVLzrINHPtIfvJukmu/zWO3Icvg/CdeZqSYn95DYE5rW7XHZ1+VawlJE+2tIrdXVx8htO
uOHsm27ESSn4i6Ock+KTmOvOrZL+F13v7qB8A1WNm9a0aZrmbRB7YlSZMTQiZbrdjx6abR2Dmk51
Sm5IfJaYFgC/ieoONJojqcoN3PrGS0f8zCemJF10znZe+MNRswuCIBq4jQxvhQgOGMsLDQHyjt2j
25g2CXYLcWGxevgc6OJ9lH281us2c9S4lHFZiIHxdYzQLRa2sRBeGAwahys96bQFTFPYOMiUZswh
QYs/pjbhRLNPmxAFnFgG7ueM+YmHf4eeHJHYZSeSJaaGTm1/uE5mI21F2Eid9NkAfEzmD/nxbNGd
92O4kF2ExE1X1KuFSlRye+MUTPHVy/36V81JrK7VuFp60rimyenjZiqCKbNLX29AAJp/LWkxbhkh
w4ed5knXgmVH8fbGL8QS+GMLQZvTCL/1K+HaPuAwgkiELsAkvEJt3GzAT4P/rPmOhvRQrYZEcTOv
NX611GkDWN8CDdvP3ptQlbfeRtd5ZfMrSK0svHc/QvVOe4LJIpFWUpP/ewFP7haKSInzwiVk/69f
OospTUyoHYcOMFHTvTmy45BPynmJe+urZrox1a6Ii7Ho6f6pfzNDfFcb931f//YPV7E3id6GoxUW
ig3US/4M/G4IbvPolkMjw5n0HBEeTqw5jpkkMUejtUNRzxUbr81r5LQsEaVUDQ3eE7DS7TJdS6mC
axa3ZrNFLNkeL92fvtB6JZOU/3jOf9Zrlh4vZOr2W/OEEZ0981a/u6VAgOfL4OOH6J0ixmkDjtyt
64wQmV9W4enHit6sJ4QJ9WZJsjo8GuAZBZ0EhUwGq1Tuvt8istDuiQ/7VXPp5bbeXicZ2FfYyLEd
VoxHhfSpnDSlWqzntqmExzUBmJwIr23bdeMLx1qWTMg6p3plQYfskf1AFiWMPEcsv9y5aDyWYRiD
zr/dUHbEY7eMvv5GdjltGSgDMgPftLPPjMtPvEVo9fpaSVapRHMvCMm0xbYUed/0yEw35pi7fwmn
0MI4gLIqsBJu8yQL3yN4N9+wn/GS3mKwb6FyA/cqA/Q3nHv9q3o4AAUF7IaulLvLOnPQmNOyikKK
FT+xlkoBCwxjuRF8x0BTRa3oXChJitAXFfZfeoMMPQEJoVwtDhmQe3iQP5UHilD05Y6HlxQUnUP8
4qbWX+WH5Qky4Q5NogxOAIpVQgusecZXrGsfmYBm+Z/+3yyUfwVuJ6i+hbrwnBxN41vkpP6Y/t5H
LybmKe2ZxmJ3vYKhvDA4X9QqljFSGSlTjwZqcsDpdOSxKJUaL70AwEVgyrr2e7L2yOTa3X4hp+Um
n/pSrJBcyEzYB7g6CyIN4/DRed2wNUtYWC335Wp7VTGayHZtvXuMdsvR2U5QNcgNZ0qU2BvmVAUe
aQnDHcfSknJ3qwYhb1wiDldVYzEC5gOpnnsKBpvK2iCBXlVFcGL+cab+yR6m1b0RGpypmEu57IvY
fqvkWrnGYdFj/8muCixpiYqBQKGWChZbEvMkuotRd68CqQcPDh/UAkqlZ9oxZQTs4OYO0zHKdmJl
nS+SeiTTdxMOf27uGHI5f3cqyHytP9V6G0gSiMjSquhPPWrAxKuhIiruoIJfshJLvH3J5olbod8f
muGt+KOU09bEsFFHgFjfCPDi1GBGfb/W3tQZUY/ar/R4yO20goIkGZfjtUshReJzvk6ngE9HwQfd
qq6C+sqzOkbbuFi5+RQrqblKuMCkZ0qWduuD4STslXaR9y9qDGDl5ukKQpjkMFfHdqNJQ75IRf6h
9u0UtJ5KpNpt6n30uRj31W5AzTIrRT1PDcPvBwQt62/S3fm3CIzPJvlmsGnmw5uLdLv+X+HyBpil
O8cATnqlZdrIfIMQwaaM3mkZSuskmB7Vq5YWmpCNl20We7rDfYFYALEASa4pyiPmuRDmf27BNW8W
wWCgFdM7ymN9yMd/X0cLMIYY8O0NkOLTTrdKvxv478pyo2BLnb8aFUcZELnXy7T/racaR0ofDIBU
X1j68t5TN69Y2tcvjr8hYOTh3/c7AdvMGIGXFnvgdu84K6DsrvQRZ1gYDwV/3wV8Q9fzBN3q0+a8
7V4yPfC0F6Py1qc4ZYgH51k/rS9ytF8Pfq737+NXZ9CQ3BEx9HGq0akSCTRineXtU4XjjyayLnus
+Zf4oPSdUPyjeVUFpIiz2zpAbFuyKiO3AllvHnfons6pKw7vu1yy5i3yzNs9L/vR1/75xXGEnJxM
STr1EAaGmFKH82aFaqhADeD7JXu9+vRRqE6oZfLLxV5T20drBi1Mv//df4kTaFhz2mzr/jGJQ0RR
YMFbQTPrJ5keZfInvsHzm73oiKsWfjo8GLTPc2DE3iGDWnsACEVm2VA3FI51+4GVu9pEHHEq5byM
UqXdiSsQWuk4YPw5gxElN1I+VeeNckd+/hEUQWBRpq6PTp/VRZlxeouMvT/z5ksyEsGdnM3serq1
BbMMJN3WehQex4ag2QVDIrKtEeb+QQZdF5geSKi6ZfOOguANkVVZhjAcRRA2FFKFYrugn9QIkJ8D
BuEyLTTgqsJ82VTx5UxkDbPElNaHtO9LbinuRuAaozImjs2/or76iCmtYjNnpp6N0gjO35BaI/hw
EcJDlMyETsC8uwELC9h4WY4DnUwNkDpVnXemolPXc6uOWjW1Jo8WBGPVVv/RN36uFrglNtxICiUd
rK+N25Cx463HFtf4mqUSsv/JykQZVPZ8wyINwptLEAFIAU6fRBEqc24rsqBDpLWhzsFBv02zNyhS
1V8WRaGgOcB9R9CytXDAU8rSMNlB0WEkuCtIR0UNQE7GjdrpuGwqy3HFhqQUntbdo4f71PCdsSBv
/fGglELYSP7Fyng1UQUj0DjBpKVb8MLEVgSnL4qe3SiFayFTh1SBTcG8RWUnAI0cDlahEs+ZTmaI
wH0Nji8gDQQb8NpPF+L8aSV+h2wisINH2y/O3DgXr5OsSLmnQ3umgRY70VXl1G/uIxvYqSO1B/1P
aYqudGmz7FBlfzRIAx1S2RqjR0kQ175gNfUGpDV+56ESpvDU4FdZj1WZGZ6iTqyNM0youSe0a/y3
d8P9nF7boBky1jGeFHQxpuzLO1rgGU2EfOV59W90OZbopXDQGT7Fnmbq/FAklxF+DmsNFV9L4PJZ
tZ9xigyeiIbgyo483g8bHJRc9YmPyXMNDBaP5WppHokEq0PeAzDjduJ8zHknxqDCbpMTYJtHQAS7
SMAn4M6/fBFHRlxATfB8tPkBu+9pwRwwB1GDXqpdl1KNkAwHz6vAXlKmckXD6uc/BH0aIhepopWk
PSpCGpDtUcKXut4Ltfl73eWgc7qm3grenJ9rlEFG52olwx46M0z62qHYwGsDfrJDlIb3hRf1juOv
kMBLjKm43OTIPuAmUzQGWTTFqh+BxjuRk2MCETtztE2/5ViJr9hCWds2ho15dDw0BdvwXKT8oPzR
F9KjQoChEEfOrOG3uPCkSz3Q0edPzrhu0YZBOLPcZ1LXUBw4YdivTqkp5SCPPnjT/MtG0yqFPqP3
f7W3EcY/cu2lds6wN/HR9so/OpuPglQRhMMouvokCkU+UJguVj2By3eeHnWGN7sPynMxmdvpQaAR
Y3y5FFgH5Xqp1NpsXL6O71MbEt18MN8dhVH1yFwO9PQ9BKV0Aqmn5kXqy7UW28mSRQ7H/cZPfek7
kYRTZJrXpjxSenZgoRCuC4MRyXoLbSDHKb2u9rxJ+EPwIhv+uUwPqeYxh4SwJk3ixCdxJH2e0R8l
QlpNrfs8QhoAwVpWDQ5/Ft8CoyIEFqKvXKndW93frfAtWVkdHRVlnQb1kBYfRNDs9Y6Mih2Ku+ES
APKR7Uaj0uuczQIbR9uA/BFVPkB3TcpIu4P8Ynm1psC4RKj1zWdP2RNCtk6u0ZyHpeFJduJzJb8P
85olqIZgmz8EZ/9isXaLT9qUuqDXdhmWQt2sCdSBzMf6Dt2QD4CwgVVpH+NNSLmE17E/+QUGElPi
yixS82tByqDuZUzn/XUREBWEzY2B+OktAI8O3WFAzzUJYZyy6OxvGytuGwjJghpbWjMvF6p1Hrfq
wDp9ZesCyohIQdRMNgU5zFVoFUl/oaKUjj5gGoXqBUMwZro7OkFmBCENKdh20s9TaZtHHZga91lK
bHxsEaq5zDTxwVQqYqdTb/Qxs0Cr8b4C7N9y9Nl/4BiARs8tfynWK1jADCtoT/f8p5wpTtkwYpQH
dj8wh7xEqRxCk5H5ygFKMF6B+5LpKNeZsyjE5xdEvITOKn4fLioUZDneIX+23LrTjeu1t6RqeJBY
2rlgODV+keLjE3D1CkDN1vl/BKCX6R6enD/ehYHzJ9sxMqZCzGDhmzu+5mUqsf7sSnPTWU+sXruN
3wh/X3HTVFF8IH1Iyzo8winI/6Zvkk/XhxDPEkNf2P8QSmYIBPnK1IUydCSGSLAeYeEe0/d5viQ9
/FyPdWtVGyueblLrokeBAcUHebWRMNydcoOl49v9wuZ92F8Irm2kFDFTTju6/OtaLujb8bH8muz1
Z3Lo/zbFp59VL0S+aI+XANLF02aWU6VCdWTxbk/blbSkBE6P/M4lb8rVYiZ+OVgfOvF2rbUc09vM
27Fmr5xPTj4HGJeOU64GZ5tEfKv/vtY+hGQ75DBKzqvgr6/UAgZsN4Wq8z0yz4/qko4ZB4iKnhUC
1NaCMsMq5zUq3y4hPP8Ci9qZ/tr1xK0vZFzRruQACi4TwV8qvyclQaYc5snDaP3+G1XDSllq5/cg
VXPyS71nkeBx0osfwC3rM6HqL/i3sHbCbS8Jz6B/32IVnOlkT/vCn9ar1K9ud/4UJ/ZLkh3xT7qR
WuOyZ6D3uKGYdW1f8qSLtY3zzydWqonjMmHbuUGkdOO08oOjHF1hmC3Unn/BF2qqwFwNXk2sbrhv
hs68OSvpRni2VkpbEPJHqKp+S7A7lGfGVoRZcCpzwmdFqoqpdT7EI39ADXPqiQYgST0hlurrQugA
yevALDGuB6Hf6W1Pi1WVoWMfuFLoXC7LGeib9N4pmZw7DueM3NlkTtVCKEv4f1fsmV9QxsssSRqX
XC7ptxs+NnRuDquBZgS/TnSfZrb/DDx9Sdvp9LNZ3Wuep7H+CdIfhu+oyHLIs+ngkVuUK3hIlvgm
amtLOfMdHTa8BogkD2PD6aorWs8lj38uBYQWyD4RPWfFvY9xhM7XSSCkTNT6hqmqyuWGFCpc2Tz7
iiwgML2BbX4Yyv1vjx+slYn7q5uk7PKoSJ5zTX+wYt3CUJVdPvRFIo2owMfIcVqPd2SJIDV7RZ4H
JG9bmvoX7Kq/k1z4hSEI2QEndd5c3vLij1NyxPpAEyC8BxwesIqoWpcRAhYRePTx2ANZMceb7mmA
N56SLir+fwXh3Zbdx41+qDs4txK4vZw/mkK7n3Kz2ncBkuCYHmTYhNfkWPAddbSZXEK9E8Z+AVij
eNAF4OIoDZgNdOfa06B2dsz1ihGC3mQ5DXB7K2xQcRb9kzVMbhoOwIdQfW8buRHinHeQT9vt3GCb
HBRl+CwiuXr015Yqs8+tmg/CLErjmRd/iXLyH502k4eiNxBdzCZ2+i2laTcAfGxiUzuKRrpZWpHF
piCgMfZ2nQUOoMbGQYQ8KEjN+VChE5ziokgvQoXEY7RLKR9sYGJ4yWKxCmBPdfYa5SDpkhmTFAX/
qnf+DRLKaYOeO3fcGMXlSzuiX4/wPG592HYX3KzLW50HzardrO4uNsPSRy0iRM5D1vLYi3qFMagg
Fj5GWcYOX7qrN1HBxEVdSbwrDmS70+xagkHCdWWjwVxvorRPrA5D9dYjQVUwrg56/lfBDE/TI35Y
rD2CYCEzq7z5Yk0aPUCHB/MfWwrqWClgwZ0GBU2KhCniTo6wkmhqwXc1saDho1L7rWBOPh3WmQ/0
/lRzk40ntM1sJtewv8Vm3AoenGygIaVTPbqR5DSzSzjZPDFxDcxyiTZaV9C6BaVOnrE7T6n1FuCS
yL1voWISdEZ0oy6mnxNjPaD7Pzk4lyaKL8hb5shJO1evENWOy2iTzuwoCcEapvtUpXz7pq9yKYsc
PK974zWRwilNRP+pHw6b9l3YdBA45DSNb0VHNeRygxVtlOcY2gHZRlYgZPv3Xr3CugI5b1cTiUzx
OA62R9xVLx2LRCLba6K/TPFQDYmmJUNeUhETgzWrD7YRNK4uXTH4C7yb8SNKmQJF8R2ipPW4quxo
Hw5zNWLNq3T4NydU65d0IkEScblV5wVtYINNCi5t5DEXz8oa+EWy9EfeSYOmv3nc5dfWN9oCuHys
73szGlIqpxCrmQhNCuOm9MvQ7W2uIQm8v5ODzaxeVy+jdvy5mM976rgmXFm7Kd41P3iHzAkd+OX3
jIH1vNKrCoUHoAQE1DQAjdhpoFTsCyXparuwsZFgk1k5pXJS7KMabd52OG47TVrEVDLuKN9DKYgB
3LD29EHvk07565bdRNNwXTVraoAl8DExTFKI6T9P91VXDMKeWAkUMkROF1w34gZr0276e1mInPQQ
JGygCRHWgU6ubiZkWyOZZ1Ie2liARn3QyD0g8PC2XuXFxvum+9Dh1pKS6Ad5C7f8arKzUrHW2rxF
qGi148nXIic9W7SHeE7yFjW6v91rSA8dSXYI3Pk9tHmqASuFcBZjCzBab+dpGO7ES+J6qUNEH7Ec
L/g3itEaCPZNM/vrekhZoDSXoTW1Vbhn+YcEHhuIAIwPuUrCIQShZaqhkR3L42pZeYqwXWeF1lDy
HSpBJHjy/P5MkgnNDlNCOvQS7+c3cPH27EEk+p15tZnE492kw0MtHxGtOlqI6WKjDjKI8ppUwiJd
HFm/FGJvMYB3wz4KkJ/OEf1OB3ZZlJKjxmt3Dc1F+h89dQRK0tAWIrpZwFGF/hXFAGvLaKQq1yTM
H/wAUF/O6msEswbS5Jo82NARR/IGMpID5bqWRBRnZfBohx4D+NjT6VG+9GAWuZNSKJGJ4DDJFvsd
Ax34se3nlzZdoJ1olLrsfXrZ5seuVQMOLKvHuP+sJCRZONCTfRTGLnm7fSAg+rJrld/IISpTJ/4F
6dZlG357u+3zgulehZGqj758P3gDoYABr3piwf44iXOg87pDNhxNeh8nUktblV4D3zuKnVgzmYEC
M4tP8NcAZYzAHzyvfBh8YOZrpWPpHwgfFiKxY58M4Hai8C8eD8ItTAwlmnJkiI5oTKT1JyxRqvrw
6EUyxF+A789NVjxua0EEUahShnahLvTu/Lp7TC9SQHGWb1rlYS4OAA9P+qcl0HCfFJ3AcbrODvxJ
sTdshw0kZ8ly2zphH1RbglwQD886FI1FWoa/GI83USP6t/tQ/VaWkTR04xbgwPkUzURSGAs//POo
lV/FdqDfx4YrNI6WGoMFNWGWwsC9xmzMiQEt7k+uwzKLKoVj1R6d0aB4BKc+Qv5/Vunsf8fitKfX
CgrCvfM9BEr7+I2ExO/FsvSWVFhHSs+pgZJiv4Kd7W0aP10zcAOpaFIU4VOuO9Ml9H0YUXeHR0E8
RJdL5pH2G80LknZfvhx9/CmOtyG9SuVcgUAnMQUxcdA73Q0l1Ibf4DFEsstswqxRcA6dvZ/9XfSY
5yx7aGmRgdum2LEFJnBTaCYV+Dh07yQmqzbwDgGQMBURWoitY8CFXsUBIEvoANs3aO2tt+IxevXO
T522jxsDK7kujpTAahs5Xg8ESeAxJ5amSRv8L19IQEvkPk1jgd+9eBVPPBDko4AjFdMbO2J5P6GE
3F57XdIznCj7mdgZHeHPCkUJvLmM6a/Ig4tey/D/cV95QQ1QpSFEi+cFtPr3MuPYmT6em7VoAn6T
0/RJNEhl5vzoGeT090St+w0GFL4jxENUBKHnWO5xjhLl/MUN41qBRZ9BuzfbqdlU2ImDhw6k/pE9
vKsTIUtv9URJJ/cC2yuKXsE/KUGpyhADDDuy8bSF/ljiG/I4T44oSz5c2S057ue/MXCPYzMTmDnm
dLTIbBu3GVkgURBdNo7glk0JTwyGVlZ6Rxq0D+L9roVnogc3O5Y+ZMSYOTaBmR5xqodyWT/2bmcT
rpBc0dYuGY9n/HPjB0FfjA14dn8GkdL9pKDHK4a3e6JEYsYdBNouU2RvjMk8A2PNGqI2IwNLnMJH
OHkB4V9HX6oxalyZ5XTbx1D51Zaw6s3SQzLKfX+FzQPXnn0BZqyWHHJ9C2cRN1+SX87wb/Qz4tbc
iBvNFaXRGVObs8RCaP1iR32azfvY0LVX7JB7uS34gU2uLjwQgYH0cNGllguW3yXJaJTsjFDumezc
SfG7QTLlMFiJBDEuaGwqVFb+zADpx0DGnsx3/b2UhXaRJi7kBBSdJpUwwW3Mj9kRCRv+qQw28g+1
BwFqed4f/BL9oKegTKgc6kof6Q9cAhZjnMCcPMqEDkilTC+eiIz3z9tXr06GGLMsAzkjnZzK9ysg
N5tAfCiWB6NWfERdB4EIBW502CkQkuMzL8jFvxWx2IPh3zdwD7oLesxvqYJjR1bP9ww5rnafOQSO
Cb16A2xm8Mq7x9rbpj8rX94+XCr4a6PrBQrV0CRKnojUBfWZdxHnpQt4b7J84LYbywQBJ2mFgo45
sCbexpWpQ1o6A8CHkfZH4xs5r76u7m42vShN0r6qdHNz9idv8tUiHYg/6bj5XstHlF8Gp67lj8Ln
OBb/ewtu6nzly3BarwAK3TXabgyYG7w1zLa01lmCXsYwwZCjaS5NghiYHBH1fO1LXA/W+D2GG4bT
QnqaMCNwwBYHS6YiCZh8XTQeK6k8UAYzOyiW9HlsskCvFKiRtW8v17swEYUFP2l8CQOpdLXz5g05
tkRaOdrYzads3FJvMJYLtmK5O+LsrcFuph1ot32G9XcOz9gaRgSdPb6ww834nDZyy+x6PVcPscqs
kikq2x2wVUIARm+OqbDrN2phKID49B3wLCYtYAh1NmRHjXp20dJgMwPu1GLl2B8z5IS78JVlHg6c
0oBnJ3H1Uq6Xr2XyUcVFq57SHz6TOSzi1DhATWQpt+TrCaUznGjR2usElxrGDMKdQFQ0demtYdb9
dAl3bLnlPGhAOS0edxND0JrGbKdSb1A9YrfF10IUWEM0O11D33g5iIPxuo5TdGZFJC0Pygu7usNd
mlMw6FyrTtjsGIpdKCAzcS5ZmPVsupMK6vUWIxpxlm7QwRadYQ2jICZ9OrQczPkg89WGFB3dxYPz
SdwBZbMFfxOvgnf0HcRRiQ9XJifhlB0Y5xpN+pDXtcrFMSHFkW6e86gSDJ9jzLsoREdwi1VjiTwu
t7L2/LfuniXiTXDnZxt9swHYAoBLNehPw9y9XpOPXP8F4CU22KPmIDKsHXbfOAatOf6ru7E82QR/
dKoWrVcKEZS5SqB6p5IrnY34cWP1ARi+DdwKW1xMHIzvsMxPnMllo4WrWIAcdMyTp/q0l4iKxB19
sJqdA3R5JEVioUQkVEKVObo31D9PFTVVU+LHfGa3SG1Uc7zLmxCACnxK0F+FNQIeUFnZ4x+bxDtd
L+zdPHau88fsPOQDkWqJ5mnwltrgNcNmM9/TeC/bF3Kpparr0wB2yfMHsKEvI6J/Ce+UPSpS7VQN
EdmZhBDKrE+g4ApLHeocqm5CJeAqB+9wmWRrkcX9ukwhBWmvJ5WwX41ag8e4VkxQkV0QYLs2CexY
WwysIrVLLYofJ/ebtx6Ltm4HcmnIM7BkZL+pv/OJIBJ+vAtoPfxHEUWBLr51jTP00nBxg1NxBqNy
rN7K77fLJK6bFj01IcC4w7JqTeImVwt291+pxYaVK3fbn1jO82fbtd1+MdLG+tAlAjNSBJGiZl/U
BLqt7u1xBB9xQl8Xzinil69vlaluk0wPBHxwpXCiTkDPX/BtDGZbNrK0VW/RDEpWlB3+WT15Si7a
mf9YuIOYTOWKjfJ38P7Nd0YIF5iJf+VqPqf7xmwuqIYqAzLC5M7H74qheHSEXmXBGOMPreYDoCbr
bsn9O8ducSxRO8WszAn2fQxdqBRJk3UASxuGxQzsKkHeTepzENNUZYDWAokAB7mihGIKxqMkwGR0
HPBrJdheqBmXIi6NfGzW6/V+q4bz0I+aQQK7KJT3TPvF8EJCimTYea6p3bICjoaBuJTFN/2HjIXO
LbVL5DxCZ6Y08dAtlyrwifp91YeIokXNl/duzjFHBmn42Obahw3P9ClX5DJNUvBg9w8uApFKh7Yz
Y69Zi9Rhe1Tqf/OlF5i8xY18t3qjm6uK2H6KVrKTfFtprPSvtp73Edk5NMeFe6mMwJ4Blj8pIKAg
U9O8OudhcXn1bO1QHIXaFmculwudZ+zr1IOA0N28dVst1H9waSAyNwrimKdoBYXRKMpHBPvbGP73
BXmai1/PfhX/CEWC7H6zMHq16LOG4Tz3SwvlpesFnjSK/QQlmxc7SdAHG4tnDbUOIs14pw1syi0o
OGbaxnRCDCwXMy/had1aN8DmFXmeDh8AW3GVYYO/k9Tp9HBKmyOulaiYh7DFF2Qw+ee3ZxY8LLUT
9BnXdunjgH/9aPvkWktLeJwbuKNsv7et2vJ5ezjrQz4XywnJw9TgjYYEohGLvsTOZn861SJ0mF4m
Bn+IQL2KpMr1W4efYB7z3fv5MGrieKNw3XFMh8seRsLJ5K738PEvuMLDKQ/8bSJuGqsw20yMegPC
2lcgbQnMefS2qN8vr6zrixEofb314vsoX98SQFBIWiMOObjySG/eiuHR+en5CdrbsoRYqluB8mH2
RvCZTrbUK6a69nLH3DtQLuc1stqmprx2W5pXKRR20eisDzt5iCZW0DGuIgqT/qjFJV/lOrvH4pdn
j5VNfREsIfl4ExTIX9+GQBclrCdhNh67Q9zi+AkH+AoK4IO126GF4Ik59LiflCVHhWaxwe2Er6kb
hhDT/ogkj1EFgpEsaoDXwZKzv122lDKckxmHdj/U0lvc+4W0nr4KLpBsUw9fY4JnnFVjqbn4gWbg
cpSmxeSJtuWf+jKGqCK7oeDV1ysu8HnObRBvLvH384HJPaGq45/ZEHP574bVODAPj6NADlh2yhDC
B8U0fH5z6T0S8soF5rMffjsja35jYKNaTEXlMJVhrCNr3F5OaQv4N7yXJDzFuJlmv6lpzEV9H+rA
ahPiiglDnBKaaQEnWgOTyXzr21QpfBYqxZpeGx3ohQkWqDnY6hVogt0aJ+UHoweBF6AkzAuNarAI
OSIqPwhXrAFFiyzWDgN6sf9b82mLLEkq1UpDrlDXSfJwHF99CHjNrKtBTiAe1PIHlK/vnSFrZcA7
DobBjpmUzgg9BmIs5N0GSXZg4oF8Swei4aqIBRIxYPAK1e3evavjQp4Kn+JqpQ42SpbtaO8X/BBy
MNGW7BVlVZq/XPqmvPZ3ZRN3LVqMlYE8YwIJn19pbPKOptxXGLedeew5SDXZ4dflMgZFdrsRkuV2
gTtYoLocmzhUPtfDCmGQ50yYvqXic9RAvmUPVkFiqnTOTW1bNYkeOYIFUtirJNyYUs0Qf6eEMrDv
ChdNR21Xpw539tfQaORMwCJhh+XHlZODEhMnAr16EGKGtpjUoTkXvmI7Gtn24FRiS9GKSLMmyVA5
clEX6E061vdhtyj9sWPCyZxwbt1VEfqMjzEb+JOjM/hKqE99Uj7Bq9rvs1RF4OIuJdSTj0J31oMa
ZTrMJ+ldLfWvoQR5D9uQDdEGnBoZgitncVneUt3c+V4uXrHgOICdOqhhl0PkCWadjR97rpI3mx4b
NvePtH6RJzkpOx5dMY3VuAIo4+Z8zUPZUKlZkhYtQN9pzQfSSq/ZLjGRF+O25bPtjyt4iqS+npC9
SUW6miTqjW0FcMWLmi6c1JWP3c7RHnYp9ru+mUCi8yDvk4ubGb51aTs6IiXiw0HKafilRxmV6/ZL
mze6XhLkudXy9vLStEWinLUpreYmt/T+P0XRuwTvwNdekr3rjqJxo5B2Nywd7jEsA4A0WWZYh9xh
85gygMZ2aZh36Inc6Y2dZfH68JvCDrFHDriPbfGyGPqrkzdwGqQaeSLd29CBtfO/VRRnQnmk44tx
r8Vc7rKZB6jGiBz1VrNbVJUl9sFtes51tjCq4Aue7m3hZR45W5blin6PSiUapsuSt6acOXgB+6QD
3qa8gpdzvB9DAItJcFD6gsIXjkuv0vIclJp+YJr66J9gGgtOmdtjMIxO6pCtiM/Y67zkzxc6HOY0
VuPZZDR7jLsVqMl6+ID9dybJTgNq0G8Jdi1XTkTQfFTFu8hbIO7PX/Nzs/aehMnL8y3Rm1fa6Dsn
o7dR28q+3jzqUIJtgZJLYQA7AJWQfgKthgmJX/Z+p23xUdM3FM8ftFPauLaqkNDT/a4PAF6wlR1A
QiiHfGCjIi7TXvOftPrbE0fqulU6nGv+kriFzrNrQ0Y7KJCejOAvaRiDyAt5ZYJ4U6/YEPZ1juRt
o989AIEJK8suZvf8CslapwPVEdu7OKMDVnH8xu74wDkXwxrb5b1tQrLMHw4xWuhLGt7pbJDHcQEq
qrH0hWOEgqhLDm7Q7g5pggWwLHkhdjmqnxNuyw37kvTSA+EO/PcsXbUDflPiLn5k1myMXFC+0TC1
nme3anHueP6MHFZC27UuXf1C0a2d0DkdzKL4KsisigGDF4orSKb1OQbkO029GvnqHTvnBQghqOVG
pm5/fSw+Y3hpnOD/rgu8Q1LnntZlfZJRhrn5vIdF/Webvdw+i7SyIg6tderR5yr8EmIs/5uYh5r5
49PMYVcPb2ItalUFvOghHiaG6nP/91d3ttWMLoOLSMO7toTsxviyxOxDByNuIpQfzADVP19WYzpw
n4/6oyn91gtrNl6Pnbh7OdfsX3yaD9tsF/iPGnUX6YHNvE72GnGHQ1/uZk6FoXstEohCPFLO83OJ
LZN86BYyUq+T4JLB3Xy0VnuibiTz1G20jM5xfJ3P4uCQKKvinmQWmYyg3uKkHY/4A2CouxDCAVVn
jUUmoV/uYY6+CEpdrkk7395e5ogBExtqNADCa3KIdX1wpPEAp7FxJ4MU3sO7HZBRIEFsiiu0C+Ue
7F9BOS0D5oofmyAwKOQfxY4weI+WmwNaLpPbx91i09JV4GRJim5R7KIP49u19pGkTUzxTJw7Q1cG
DdZRxt1fHLdhB11H9RLhXhODp8IjfbwhSjmEUMpEfsmm09PPRbHYwbzfKdooVckgirWtQVLV/boT
5zt75wPaQ60C6JzMeocWXz80BWQ1c1/fKr/gmcQEtvpId17J+q+HIZPOnncwnoG/rNORauve18fF
9Vkb01yS1Rk9s/+O2Lgnyu4biSH+MFMDG2SQ636SJUmUWXkMLl3fePl/EFnq30FUDkWuhvFcCzSf
KQxV+PWnnwWyDLnNtVcV2xmnLx2h/IzgXoiHfWdTHVUXzZmpoBpmqf9r6HrtpjCTy9IyFKTnKXq+
gm+rPuWe+eim1D1q69TxsyGJsVYNpZ3PI56B3xSoNsGH3lHRjrD/RobDnNhVMnuPoa5GgzSbVeN7
puUeANUTjgbEpEBIkQzOdc6Ms133T5QhChcXjxBDnCoR+Q/VAYYJ20P3xoBIhtSQ7GdJbBYRl7DW
P2/KXR5VIggSudOqukQ4wp4iYmVx+22sMuqLTJUtSwcajV3i4tqHADtqIYMnTCEtg5xh2IzuVFUR
U5wKABC6rIL9nklorJYFiw15tLrzSb6a6+0q8MXzeaQ0zFKnfdDIVKCOY/mNwoCcI5VHOIl2wpzY
VrqnS/RWm5lk+ksKIOcqPL6hBQr5DDU83biriEw0t2h5izY4x5VzSAcFkfaYp7zpS3RUe5Yahb03
r+qAcP7nmUAya42XB6jrz93OWGPpQTPTql/zP6WTxT4esZ8HPw3Yt5WGGhKLYn4JgIA28H78WneM
2LwIgUnICFCFbHVt2oWh3on9USuSy1HUqNOKqt5A4u4fN0CY3O0NIa9BWf2Jd9IhXg6+ppMqiaJh
eWlxxFXa5JvRxFiivyip1jHwcy3jEAcEXUmTuRyf5P46NNeKh7HrojtiK1MQhEhqq6fcGTzm5V8Y
nSDivrq4/Rh0HHSKoDSNU6jbnKumOHrxNu8Dfu8Upfv4n+RNjPEirXruvWL3sGIzxw0i46qpW7Ab
iYqsGPoe+t0dfirQEnMgSmMIesP5kWwrL/wNYiXN0VY4qlLlyOIXMlqFJC7SeYp8GJtA+2M0pI6f
B8+Gn7QNWTJyV2beznC9RbGgKJ1UYHFjcJV5sD4b5nNZFJyq+zbCBykA5fgkyrSyCHjyY8LIPCU3
brjGtU4iX3fStW8PTqvKCWySY2ca/HOFY7P36mtL5luqupKUesxSzjoVBH1GtinR1uktg3C0wPvv
pimMiagepvQYvbOpYs7T8zSDtheoWB1UMi6taFT9/utPHNvsjjFU+shSTH/GueZgTuzYPmhoC62x
IAstcKaTzKmhIRXpo+PgKoghouuXpVlAiF2F53XuE/M5RflIrIDH2c+2cKWCW+5pth6MXAuUsAnl
snvauU7UTAnu+raN9RbPwdR/FAEhuGlnnMb0jePw1JIBoG2V4u5OH545Tl7BSTN+Syxy0dLE9NZP
MDdl1BKBrv9aJ4oY/PkxENA/d1tZ+wj5Z6dJbL3mgQVm/cCL5RL4KF02HcQMmsasU/AZy53mM4Rq
dipMQUDO5f4KNhlxedcoO1iWjq8ITHrag0HEGE8EjDyB8hWMzwsOrScchtrfzJYdZYOvt6MkpFLL
VA0CMMuY/3oiu4XQw7kZ9wO85EL9qs6XfJseGsbDL3p6OhLZuXdVWnKTNOjzEPhwbtDWiJsVgQtm
TXTn14Q5+a1ohoLkgct6yah8gkQQXIuk97MQrKTDpittB6oj7FI2FwXF7Oy/ifCd9a5zcOAOuWwb
Nk8mSCUAdu9wnTPPcfLXh0kdHoQMUWdWD7mK2WytNDa6NJvQXzyHTCAfbYf3xaEVIh8i1Bpvk9Aq
JcippXZEMLYLBlj/Pnwn1O7NjPyvY6iljXbjcwIR9zm9m6GqxV1oe3vNvuRRgVyXFd9gHiBLQRg/
UQenxZaJAtyrxZkvZ4mT4WQ5wv0QTmdFC+mDGJZr+oPvzQTMY50Uf6ojhnLMBhzG+THr/HrEn5Pu
KvCY/5OQsb29zpPMItswhvmPsXwT+JJRFMuPXjQznB1FY6qMipO1abLQsKu8tfaHQ6mMJVWINr8E
Z+Zazvp1zZNOulc04fRJJ3U7JA5Wt5Q33IgueBRJjj18U+d+sWQejuJrnHx/X3htmAsLM1YdJeqF
+rRB7Aqp5EtwYgTbfdDjGMWqZszpnMUeQUsj/03USKIpXIsELnrv0A3tY+a/8nrUdftZ3POMKG7W
lEfUNAgNLhjFVn+iChq1st2Ak6dWOnRUkXgKVmqiIg2PX03s1mX0+pOq0MRGhG65ii8m0qO4Vg5v
j3rWhM8XQfgd1d9SSgaas231+U/96ggDUVbEATL0qX50Qgw7xLDNz1RdQnsbLjVQpvX47dFJDqJv
l3ogjacs3QYc5l3RKatB0qEBWIHCDthMqNIgpmbxaO6aBiTzNOxVE61aWFIR1zfTyxbTqq/r8xFK
Dh4KplXCEDkhj/ziy3sL7VWRdMNCK5WVXu47lbCalsPUlRXCB0HwCJgUpLFYQVd7cMU4k4wUK2ro
h+O1Ux7uIV6hc0RjcPXehp5LVoWssxl0vXINTDVivcWosO33R2ymrE8k0sNn6Enxc3qJWhzvtyv5
FWvpoShEqX5jYqkpucpUIq1+yBzaFZjfbT/zKQGi5Bt/4rAe630gf4frEu3haeFi389WiOE3sfPY
TmSmROr3ZHhFx9GlG4O2adJ7tJF5OieohRHyaKaPjLJBo7S799ndmMufwucnjdvd7JUm6ySnylUA
DK7NBl1koYQo1+tOfbhBPCQTFYithSFptEg1E3WloqGR756aSpCVGN13Xr03VDMAr46zgHBWN1Nb
D1t6KZUHTSVlJjSGfkDCMlrQuovFvDOr1tFi1x6Ic9y4HunqGUEyhw8lqqKN4ErD0n2ySTrdWIJ2
7IfInfzSCkQ2+x941JXxWv2WOUyXytoVlsSBMXri6hVJSsWT92h8r10KIXfS1w3WdIPbaeOEhgB+
58pBb5VUW/0cDjj5nPZANXddAXg7Wi7r61r7YrwNKp5nkyt9rqXksqTgkPy4L7sgMjSqUBSr9oUP
IMfOWWX0D+NeDosFylHub3B/Y3C4IsYR3n5pyoEw2OUX5YlYhC6Wbc0J4vebsRys/DFY8UdwcuD9
L6EgmPQGOkJh9VQZw5zxYPFPNUaenAU/++z+Oc5KzRxUKmoy7R9ewxfhtER8d6cxailW9G65Wm05
kJ3ZM3Xbw6UZ7LlkO/gqieAhEY1QdAiKQZ3GG21RbJi2NOCF2KWTIe/vTL5i+nAEWX0va/sPGdD8
DDMyKjN2mySi1msPGSR9lbnZ3cKK4izZ3prGjtMBZYkWROF5615pqTOM5ypeVCsz4zPGei1XG4P1
YDZKXm8v9gSQ2ATDQwG7ehSNKm9266AfBqG2TAViuVEjs869xAG6PQ3GtEwU6/Wg9LR2EhqoG721
5Eaein57xLYR0eShhUQBPWMqKnB1QdjXNEjjU0xF9B+zwcsW65YLiyDezR0n2u+LE16jF5g6U0nL
yFJOCTs3mnggzausRXbAfnMKECBDUMAcHsqwbiz6Htsuyp5HoHQKSMw0uHve5spkYoOcs8DD6xb3
prGgDQRKMeZbJbl6zhzegC5ewkrCzvPvXDIcsKd4Wdk7itgzTYJQ4laGzr/IjvIZ99qXiZ+tCOKI
DzMhRxNLtsFdRZoFNhwVpTl9KAIZiZJX7+HyOhr4E0aIv6zu44xP23+cl4AgHKtG9yOHoKmG0yAN
vX+7F4wdfkTrC4pCJivodM48MVzHwqIdSo/q9NkMteokTM1GPlRSPtVRIuhQ1GGPUkygHnDdfVcP
tldGAgX0LMBxTo1395PVP39gFKEU+kyj6o7oggkrTE/7IjxeyxlvmuUQPq0QwKqeX5bda+cc80Zd
/3w7w0CZSmImc0o1bzaufyeQKWTDkr8DG2ffjI8wlkAcklUq5TFQ8xxvFS+UAZfz8sy3JvlKM6Iq
hJ4D00wPRkfy049CtTuiDIwIG69VZlxAg6cz6ovRbl5c4rliQLkpEym3f8UUGfkiCKsEZi2LQZnQ
7Sq5ZsnpQSBrRlasaCmoQfc7AwdgP0HGFVJcbqh63BtjMvG9Melzy1tis1hkHrZcY85jDCi2NUnm
tfYxvawchjso5dgITTr46zq17djEnIYsug/99c3rSaTsnj5D9kyWY6aIFcIVdUvpF/cO6C5NsoUY
56+7+v5nyb9zwwxRlZJNPi7PLMAHE0fEQG89ikmJ0hvkhuHydY46pnyifv1NyAocCn32w+1ALp2g
CerHP5IkEW0R2mB9gHAZ8zZVCHefgWdAQu7EnbQUG81yfTWBUVj/63DHeFh3X+uWNtKJgsGxDBPI
8PXIQ5ct7b5aeC5sslCVtADLEzSCWPrPDNdl10ROBppF/7VcDx8hmuXsajw/9q95XUiBVSRAWAaQ
pSw5PLMmNH5VM+uaPDlWeC9xOuCXTpT7CIT60U8yBp25XJxF7g0m+7Nsa3ME9C2gwWvRRrBcDdmz
qwMKzeemyyxDvEMPAliLv36d019j9I6udcnb/C2OFygHYagXXpGwH27NHV2uEExghduf9aMGdNLM
4rggfH5C9xe+Ge4QaXV/sozm3eCcLLlee0bNwQXv2So5nasjjHXtGOhbP8f+5nzY6ITe7ngjp4Te
rmh1lvYHCYsJAGw6IGcgdq1TqbAbNveGK1cyRWC1M5ybzEHUaNnLnmuiH7EJDDIByEW0M8xNcLXl
pQ3incMCQDwL/l/amMVy+0/nDewLyCYyoxIFMrdeXzXj7uNPifDC8uuDhuRqVLf7BfkfcUIzGiNx
RcsT/FHm3FmqSqT8tXt1IOv1EBPDVleihzZjPkv/aCL888qy1lNmP7Vd83ciLBZTvLN/obX1cFHA
oFVndX7cSMPedDjAr+NP8sGgNwHkjf5cVw9NfpW0Ne+ZPRmoqPLPFz+aC0D3es+fLDLUS37/G8cK
LDz+sL7B/WdNuAz/1/AVubMGXSKtBkZoozRc8hzAXFWUw7RK9YNK06zlwCHX9/NE2Od7OCn1TY8v
tTa9rAU1urGKGfeOlHWU/28ypq1gyv4CftcvgpKEw0+bAmIbiscM0xmMBURgIxBJI9hy0HQwHaND
QoQKAVbE2/YPXxFG6ywEasBKbnVvjpcogfk8MwKw/dhumJsz/cwksrO6dV+5WFiMhOyff96uQxnL
9CG3Ke7L91R2H90tEcxiMhyWH7+qfe2zUfd54W8Tr3xvOxuIn1fSspCbWMwyiKyZvJfk8sr4H2QK
Kq8GXJpE9KHyhmIVNLssdg4q2EY90aiylRi0qWVi651jsIrJ8qrpw4CCt3Pufi6O7HdNF58JRdSy
fAFZvE8Kthv0a+RFRqB7Jjm9q77T2mkLiT10u5NWEOI4LXSIomsBoQeK1OLlu1EGWmGt89m1qbTy
BN5V17nFZeP/EI7c4yharx0+k2wRpVtGY/k5adX4ofnng9ZdiuzBJJO4jgyzxjNNdjaO1FBkWQMe
SzMw4WSdy6pQaMv8oqfjYBJPMYdPhR2U++gsovcUZBwwCxlSiBmL6Xuw/1pfuegXvr538cTAbLZG
QY2kx81arUTeHCTGJM2VAoKfepXWbjUAFU2XY3ET5VS2kwxCY2JYyFa2eHt8wuMm/tI2nSKdL4I2
1Epun4ts++rsWzsVnJBNspQZuYKY+LbmLWxNwh+KXHLAhJ8ovKpQJ5HHTWMlzJw7ktliCFC8E7ai
iwLyAdnRGkYz3Qrw3FYpa42bQUvWaXi8Gm2GVp29CPJ+pHiwH1qrlr1aVEGKeh6fJiMHZfP3rp/n
hKuRSPgilNKjzCrDo3VOTFLYW4el2A4QOan7upCuYX/kQYFU+Ro3vlIrde06QJVihW2FCuy88xX2
VFrS7iQdKxTHBRUQ/luAfc2t0vFEECizyV6OfXMJyQgOaoLuadpd4C5NdnQZpYnGYLF35pwd9BpS
1riQU2YboG3zQfWlK4pJLFFur2axTtXiPrFlKRpF6m9kNrAsQrpAmEc5ZPPmaPRCN7mjFhppTixn
WQWds/x7AU+5MZWuUlFVyMn1CCHE5LpbhwQiCJj5YWgd4KCOeWs9CLMsKl/bZ/e6RnNqainlg34w
Rtv33QASDyPhGOYlVGY0/vfPd0mYjg6Q26t5mm64r3tgP5Vx2TyROFB9Z3NPf7AT1WWhiWa+Gykn
Q4JV6QWYRZO5QiChbYf7LzKHrraWgKaXVcrMVzqVr44AN2xchy5Sq/vltP62bcF3bU7Bt08MvPyD
icmKrzeyVQrHfdPbljtrxr//w4Rvb0e1UD/PxIqDzjGBsWCAzaIjxWUP76NCKJVnpotUNREEcinc
FBtYfT1vc7MHHUEYUT3CtjmT7hLYRNIL4vXZbxyJEcC8KsrlOli8Uf83l2PEJu7grotL2ajYxhHt
4Cx1DVuxYHOBx68p7pWBGSuopku/U0KEi0MdTX8I/Nro57pRvYgIsyHYf8OJf40yx1EKTb4FQBVF
lQgweW6ctnLtIlZK9iMW+/KA7Gu4YhrA++h/VnBsou/ytTWITuz5O8FQaRWHz03md0mT0jPF78kP
MLIlO4v1fVb+Ik1gse5njxRAPINHiAzHalkKSDSqTjI+V0AvoctPSR0LvFm2KUYhmF00k9o3vcjh
uZKvt0l6ScR0JI56V0JMsWE66EbDF2ltbCfdr/eSd9ctO27gU16kSsGspSi+imrn9/K7JeH6gIEh
7frvdwX9jhd3upZmt/w2OFxbkisn9MvleOi8TmivKX9xhd+g59s+OyYOqe87MZoAa41pJGMqxg7t
2BkNwVwdSs1/Wh/zz2M/5p1gPiLRWWSy8NqbNrZ99OPtUNG6J+Bf28Yr1gVlk/M0Fo7XfnE6sk5+
eXpeVoN7rwlcCcCgLGFhUUkEpHfy4d/nMgL/LjLh3G6G9Xhp6BfBtTHHi/bXrcg0hTIgk/5LuIKM
fB7wIDeEy/LRI+xjlj/bQYAsFJWAvw/tL1DB4cNi8iwxhVbs5CH1rRL8BRFbHiAG5nJHT0b9OKuN
xAXcAvoMixy39GLpaztAMiAlTcaX50YzG6YSadmocL6j/4YCXdfz7xhblmLhPGVGLdA6hY3BfvDE
8CaWW3HJCx7yXApHho3YzHNQAa0GG1iq7CidSumsrKeCDkGRtW182oEr36wV354dDZOKg60cQg9X
5hOsMx/jEJWcgA9ngxHpRb+G1KdRXgCn0wXOZa+5OBgzx123r7tPeFqeNBzO4c2l6WY1OwQCxQsN
Y9Re+5p5gnx6teS6yaoJ9oBZMVLc0JRekD6IWEF4O4VrwSbGfQ9Dfzc13dMCyJbKWJzK3i/HHw9p
oYSwoz3dkLIdzZRWwSIxTQ0Am5gMMhYOKTbzANlE4eRyUpklX4Hc6bRsBnwHOZwFDAAn1goyIJIz
al3Y6EKi4Wzvf3KMJU0zArfvBCdX92PLOgjt35SLdCYvKXJKVM2KBRFlz8T9hmHbRceqfzUPgqkN
DcNvRQfGLulWP/ge5Vr8XLEet2BW5303BuNlXUpSkdJE7Hb/nREAIEdHRkHYu6lvDT1+2XORXRs4
/SA4+Gar4tQqUyAHN3lPQuVM0YC0TadoOrEd6luehXM08h1+NrbwUrVd1gkii1sW0cbhSSi+jfM4
kp5XxS3KB45prEJDvO4oGyyf7VeuGiJl9MOvOu3woYPutriF4aJRi084Rw1Ict5Pl7Ul21OPKtI5
7qV+A2s70zryFOdDqj/87WrZbKuObfh9ObmNfQUJ32mTkjfSKhoPP2jNuXQF3Kynxsgb6qg8AGtK
roArpElOmM6D54ieggs8zWvpXram3aNFlUTvQ4gG1FKBqp4xuAlSZOAqwEDMZInWBbTnoACRbObr
bxmxiBPQEOStLtEbgRTzvaZ2e3Xg+npXCjKboHyjrGTuxFQmR51DwAzM830lYL4Ad75WV/XHJERa
Ffi06imAqRULPlk/Mc8A1aDXRS715K2R/Tch6K2U8mwwHN6jyreytfhXpvHDY93inNJvFxIeWfme
bjwn7o+j2l4HCrxDkO0Ey4TANh+6/GooabTa/nJKQmD8x+ICXsgYtz2u9egKo+lrhts0JfWCoXNQ
5xi24jPc2iYMmwo7/KTraCuqBsoqNUHF0wwkGIV10EfSYihdNukjePqiZ8PA12dM6C4J3PJ3yHrP
mIuWpu3ol17qwCgOaKtsHg/dgSTdEAY6G2w3WonrVLKWz96AdPiRZJ94mqc/td8AZcoTLFEnydai
jjvP3I9PUIR4XzNZUE2Iri2bsGncE3cFd2vbFzzNw67j9vGrP7/To+BbUOf3rZqFqrrY2DFU3uik
do1o6T72uemJIHe6ap+KSF1pFw6BsdnRpS0tqSit3E6cL5NXc674Zfk64RytXWrRQv4WsbNBlFBG
2OjLextParWtyMFeJP14t6G7WDPcWpsb+mcQ2UEMsSABDV/xupWcam/2MWq+4Ovw747BjRUBtlTz
q+DHVnVIlZeQOPf1zwd79ZKMIOZXjkDUG39bCMA+Dmmk3/c3H/8w78815FdDalvqC8fXNfEfU3vy
Dwndzf0wBuHJz9qSx4M5MLQlhZyvPFrA6QD+EAe0Yg62MRHrhRzn2wMZrWykybNAQK3NQqrKLcrc
JVSf1XIwtuxrgZrIZUy4SrlMbfkKPWHADdKxbCV8JuCdggXafPdQzxgpdQE9W5gV1pDpzhoPIIc9
qqhB1R/0Zg6hiJY2reRNTYikX9R7eRUUBuBmI/rkRx0ep9Ha5kVT83VyCjSjz4q0ju+XQlhCiD6c
fwA8HDlhxnAI+tCTAnbmyVzhPkMtPOI4s7alFjjpYcpYXJeLd/EnFAfIYIrS0f8Cf24XbuJhWPF7
V267jT1f2X3fHy18Lye+wUcNF/ilxGKIC6Hl2/3o+4R7+hVK+EHVMjrKt/q+PkLkyHzG6vcTKCsr
mMb6e9RwPFvom5Fw9CUjxKA8pNpTYVijhgdT6xHfYLIJKxlcWhi6xpWiOv3m957iGyg57M56vIIo
yvKNXiExmtkvRgxebdPgOApmoXrrX2e2zfb9ffqW2UPSYITZAEBL88RBT8K8Q+64jxK2n5wHt1B3
nM5ITBSOnBX8qjejdcgWVvf+7V41ZPmusuMGsRyURpiYHfEImhKSQGrRVWngW4/H5PT7g3xJy1bY
UOYKOw1Vhhec4PVVVQS9hBBdGmGTu3pMXSeotRlV9B0gZlj/eP8G7jOskfGnhgybeIppOTuZnBCk
g8/IBWIQ1+1uhqYv8TfDew7q6BQVeF0jDHx9MDjAKw97s9y75IkPZqRbgEt+Y/t1sWiVn1dW/Qyj
IxeBKDjGwAkg7cDrq58W6iva5Z4K3vpeQax6o3DxMq3N7vyM20wq8gWn8uNWKCv/zWpWMwKgRhtO
Zwyjs6rkuaEfSj4wbXFvbHYMHugofiC7a7hARKZ52DdhtQvE6OJZXFejPqLs9rviGWKCNiDGJV6u
unH49zqAY5vSsywwk/v1Zjglz6pTVWxgbQnNgCbmxMTp/G/aaboj2Eep5A+od+19mwq8tzyOQE06
bn1koEmIKRz6DkM21odmvTTqg6ejV6xZpTRLZ6GyTrHUEkzuhoOJoe764LlIu+hauawGB6MKhoy1
SnmZkUwYotyeHJToSqB3VtKk4nzMu/syFlUAcQxAWGjY4KmIj6ZkYUa/yBvsiksfbLkyG3Q4uoJ2
b2bIJsOiH/bqyupnVcEi54CPKwzycpYGJRBH7dxIZt1c2sDvUG1QvCO+d9v0rk0QIHIaYVL+wL6x
8bBP6VY/13odZL7fkvPmuQ8EIaUPmspSTdrY+DuWCLsYJDJ5KKlAKLcX8Q5Y/1lwbjPeqh9Zmtvl
DUTx7ogmrWPGme+EsfwPc+IHN0ge74xHqUzXHjuzlF2R3cxosPs2OrBRZVLfn2z9LpHwHRm+wNPe
C+hTqUHEqdhalsd05TLD3OhbtuR/jHwoOmCwoTLbjIggtNsF0bGLXdfnR3RPFq4zwlBqZ7jfQ0KD
XKOzkd7TgJ1W3gET9J4eYdtLsBzuPybOavKNays914rd180IQtEIe4T4zPSYMMX/8U+nBKtUDP6t
CCPcpihCk/Bnqnzty945jjrUWRBi578MCNRi5M83ZTRzLDD35W90j0+JjRgVd6Yjr2PSc392AGkY
+TAKW13FMpWu4D8ZVlnSITyXOX5KGk3QoFf0kCfzOZ+XVuvEOlyZmUQTNglK+/I3tFXYFw8gehcP
m36SDzYSbDYPq6Q4OQekcKHBfIKADgrVcU9CNMQpCFFV321zYmkiUXSFPA5e529GfBO2jtq7MLo/
lWFTdNHbJmYSLgbo7/jbtqIBiNdu5VSmFiFi1x8MocYNDEJlQVI+tw6KJ3vZsgu3KaaBOaK/3jmA
GqSIA/3nKi0+qrbVNKISIR3tDwYOeNvUEua/Xln0vVw8Ks7DBUIPgMhhtEmuBuiMAZ96EC+VQmTw
KLJR4UBJwnu9D9INKeqvO1LtKwo6KlS9p/tnSbxfE2NoedQwyc13ur3yT3GjijB2DWF1LxyNyVdT
M7R0FswlAxd5f6+i2bHpJIrB9AWEVhR+cdn5A/pyMJ4m/WTjQsUj13CSj97OUS395OG3YTZlKsqr
O0D7hfijLLV6Rahwtw1ccxek2nYG/Vy6+I53RtXUfEI5FHF6XRNMd8b1kr+irJBtnJiSGkVa8wUu
XHAYBpUCftc9CgHOdf/Ozuq+g7erXSJ8wkeMlK42tziAY+Z0nL7WImKx+z3RGammBBcwHpzyd/Sj
F7bqyuvcmM6l9eKuen8+CP07xUp7XCyp3GshImAqNT0z5WcWeRz9zQ4rduqoVGiuP8xfoEACm2r4
ZUOblXBOr1/10E9HV1n38+VNjGGHdv4zWJEjM10tCkxCCLvuC6MHaSBWGwWidInuFeRSyjT+XYvL
vPqRlWU5uCKNApxDs2uRRvAym6mOVqGyxBbSUS+PawDzeS91hHsLQDqy67lquWiO0ibE4JwlpJUC
jCmjrsK1xMzOETpdAAFSCIF0OL6Cz3X2KhQKtG8V8Yen/ywggp77D7BjFW4iPLv8x+KTLl8xZJun
pmKhNgahHO0I+d/Mt9EzgWANnyKJuHISOV9o8ATs3MBKYx0kscRUBZg1oMQQom9bx/A+1ag9UpZC
zue64n8KbNiKTtxqahsFH3T3DTExc6oxc4ckna5nI5VOI8xOtlUy6jBSoxjzYP6Nc7j9EG/yMqR4
jVv7DeK8oCyCkCVAie4X2bXm+b2SLQcrPTOVy7y4sBOABk9qnZTehKA3pAvTBPa+PZagVHZtBYhw
PtmK9UFkTO0roLwBnhTAxHUgt74LnLJg37GdMT37aqkVxhs8PfaoBLsOsu8hQk1cIAo5hAb2EZqp
JdHZ1Niey7yaQzRoFzBWfDrv9HFvb0AkKxt59PoRKpo+syfSjt2QszlpLCD10XED4l/saNqQddlv
WBnNKzzPx9nJMOA+V/NpVl2OmDhH0rsQIyQgazECpIV/DGSHDeqlf5x1dGyucc4ACxxmTlD8JqVb
e0e+1v/S+1XzcxbrqIKIceW0WbV5+iiAfrWlXAiBnhAnIlVklPFKzi8jXmGjb2IWHFLBlgOUX0Ns
4GxAvcW3/331mFmo5T0CfZTC1/Yr99Z3Ke6dqXbsZRxNwtnYtczYUJ/upzjiJhLG4PAWEJ5LY3fP
eCcxkCxBpHLWQm3TMDKQikBppH8KxXWMAh9nNEM/8P7xTPbuEJLVYVG6sN4An6ED0DLgBPSdhSvx
UnolKxBJ4x6ClCRJeFiQXlDl5R/5cnsUkMBdwvvOhklUiO9MCOB0IDcsrwhyWTbHf43Knd92DpBq
+JXDd43uLeaC3HR9aBYMtv3iwuPYsOHxgqTD8wYTB6ToAVQf2BDNxfV99+X/Dj43F+cOXgkQFnZH
BNb48tUJ9jUq/P8DQsg6L85ycMAjcB5fsMGRiJ5mwWEJCXmn8KS9Aqc5pAA9TPJ8UsArZZ+9BbmO
jrOTay28dwHEt6uEWywvkXQSD3U6fJrzoiFuIa5OTeQfbR7tEV8InkzVYD6tdH6JYdFc/W6OC9q9
UMNvzwZuw9t1mE0XPnEqOjFFXJ/TUM3/I6tcL6XyS3bTx8fgnbcGEOfgBMUpN93yGGsQ1xrPc3HH
ghKcOvgf5Of1dgo0jQRXCcGGV+O4lZU8E40p0pLgpW3Zq3Ds9Tgw0suvic/MnnEURnUk0zsbFT0V
a/UnX8yMX8nQyGISlpHMJTXcTHeJ9zsANsalRu3XhGqv+NmwFLXSUfRYuRZaM/7FSlW1BgFbAYwx
wdjqM4hU8kPEKlDbA6zHlgSzwPRPPsPiDZBRnoif2txlOcX+rOVQlhHyaghOBd+qy+RKcEgWbb40
G9WJ8P7MpFhF9Es1NNqp9+AuXi+5CqVeoMjXxT31PsBoTLXcOQcZdCaY/oEM3VeEGqk3X4EwFv/j
UnYupVKf9k2gppsaONbBkac+OwdGyx2Mo1QmLwjrPv9uCToURMiscSSQRjLXJ3sF4SRtUdGqVUNC
io32R/njSVeTWBTGyeC8mue+IQaM0dY2jT7BI1w/RS0dItDad6nU7Y6Itcy3D8+KBtu34OrW7Q/W
e0ByV6XtpoGC9nnfhrHf7VWEnI8Xgr9YRnTZXNuPBfFILVO2YLW58ITENwL5vnWj1CkPZVtBlARC
OXYtS+s8HSKlOPjUi4pShaZZwBpqJBxJuD7HO7dPR11N+zT9/A5GcwqEWCK4jzwlz55HD8W0i+aS
Ee3Xw8Y5vJUkJqRZqSDX9hRzXWRxicWD0UDDvDg/q00jHGA1S2AXRahj6F/ngPxeSf0SlNWUAroO
A5M0CdvyGjv+K6lkIdPnymXWG6YcPWdbHcml0U8FPNVgH7QMiC7teQM4jS8NS6cNsZW76GPkPOJt
PdevLs8XkouYxbh2G1Lnc+G225crn/fRgOhL9wS+Brsiw4Eo7yFNNrmsB+z1c0iPaP65f9aqt/zF
Jl3eXqj9+HUYxECslpxVSjk+aM8sXrvFg3Op43uzv6qH96UtYyFQ41kLd/jFi+3UToL4JTMMo9bT
re5da5kzau9Q0kNPqH3l6RJjo8Euf3fLjWXxq03AGVW5HQ1DPgt/8aWHEaRh9cLackgHoeUh0jzT
no2pEamL+SPkxsTzvPvUnSYUdyyZV3XC5u5ju2yfYGiSbd5AC6IHciY5iKgDrihB9KwYWeEJluSb
BmC32XG02T0QT2QdmARuR5U/1HA0hJzB7pejYuVRbI0p0EldF2i2XXZwUdRjsBOmPqmdfNbDgD3j
TzwqSTmmCuMBNquy3QbFykiQyTmFREN0hN0wfxvBdojUz3svGNjFqQ8uL+DeD3FQELoWWHSburLc
KCfIiN9pfGuhFpKNd7UX2A9kpewk7dXiAEUosvloBP/D/A7lcmtO4gA9sfjnlnbp+45baOjpebxE
ULBJyDOhg6yaXA44XmS9LecgnxeORew4mFVSrXAFEUxLff+q/r8s1r23y+FLfaQsVkHZPUst/USw
LyN1t+IN9OMKPIu59Zeir9yEe6Qk63Dx4UbxP/5vnpY35IQVWpbTOKnd6LyHJ22b3ns3FhHOFTNZ
pwZbiw4VYUVuywQOzdU1KljPEg/76jAdcqFyvzsSbQYf2dqyLn31jDlY/UdGf/NGtoDt4srZM3f3
WKF8nRb91FTUfiMh/2RRSgS0/lTHQydH4bPhj7/Z4VFJQnnHiYcCDXqh4lzmWrprBsEw/L74in9L
VJCKyQ7lGoAmJgxvHnKqUIPRuhIAgSzf0113xgU6CbUOqDwfgoNTtW9O9+NG47Y9rY6nzN67q/jr
W1HgTCLZG5+r61C9BNtWU1DVEl0F3B0Rgkj20sWVxvn3hs7K//ohXpik03Hw6xBxG5A5q4ZMm0tz
V6cp2gCbrh/fnuw6Jq3VhrVSvlInpA5qMccJBeIdZ6SmFZtWzr9itaTYWY5UwAlCSpXEU6AjuDkY
QDILoEobJ4QuBE4/xPsM20LIXyrnWym0ShWRf7RoHPwvhU75prrTM8VfiYf3ai+L4G8uQ9bV7tJV
HyOSiz2AOuMTew5X1CxBuLWVBMj5crr30FUFQFegbEJUjZUvB0yBJIzAmDG39EmM6PuPB6i3X9wX
gjRseZ6UY658J7opTRxdkBjoEhES7ov59OL7A/rrXg4A80+c1X72zvvs2YqtsU5vF7Jv8qFjV5gt
athO51/P1EmyBl4PpIUUGSrDwhYzWPxINXDYeQbYloorboYSwe32/G0LdrImolHdYPJjKBTbu+aR
+mbBLFZxK8hX0U727l0CBdHJC6EljUGENSEn+f0IUCobAnPB7wkDZ0U59xhracocPwhqwvnISHbJ
LU1K2dO4/QOY9tswOzpAIfaXN+mRmRHR6HNiYZti+pgqfRzYGHLCHCYCGcNiqV2I4916CBSH2NXU
002VLfTEtCffF0i+Nyau6Dha4SS01U/gcVI1PMGaFtXMdX7dRfrUbRHo+1nm14q8m/CKiDkeS9AP
+VJiww13luB2CSGsJnMs6ORZFrUekgODTloCZGdOCMCcn9uJ2hGIue5Cifd3HFN0ZzPR+0egHp/3
+hWJ/yncJ9D+2W1ntny3iG5MKbMJ+BCwLM6H73nu9jEqgxwu3yAr5T/NI1CCGOs//A7yUXaNDgaZ
fhHkcPFU4RV/r1JLryY+i0lmtg0pjHTmBqIfwgpImzVF3NGK/zuEviUJ2MCO7dViU74uGb2A0la5
lXwInjXAmqhXRENQ8ocBBRU1aD476q84wSNllRfhj1MiQ/uQcb2dOx5mp3jKO/pI0WrJgq11egKR
Efdefj+exd45kpLtJ4VzlgLPPrBmNltjKnuv8U6ZTjKTZ/G6/BZjMmm5uvgPZMTS9IXdxhzdTVgu
fZtGxaJV0xVKK7w7LPERXBZ2ilw14M8qeE3iaQLSw0NOxbUAtu6cvYQlQJ7DMxb+mrQIteMMeGkS
rI9nxFxPRinACKAfTEezVWcKNiCs7E6TV36UwtsqDK6Kxr3kv7daIJAV40otOlhj6RN8cbh0uUu2
/1zYHQohCAELCpZ4qVrsHASSrgecbu0lE68EBI6K5wdQbrhhuFw2nChMZE5OtVCTDdYqcddqCS7I
wwBqANEnmKU2otiWs0qyscCC5CROE43GHx2gNb0D6+pFcpr4Hq0Ih9yQlL4zz/4uFLWQv84kJhKe
hB4GF0yANfN+e7Yaxy92TqVu7WyTU3T4mAJFlJyFNT6WshSKAaL+ltiXUVG2wWuQYEuFUDXSFsKz
ao3S5wlkfdPAJlFWhuI8prTrTzBCO/BFvy2Rj4GKWcSBxyaL6K6bpQL6/PnjwhleAGOR93z98vtd
WNqB5KhHz3Fv0KUZO4F+v9vlIoeaCIzXvGvsTsSUO8fv0yO1kBMxhJVd1pk8KApGghJ04lJVnohm
t139QPNNewveeNPWgWUIGZFuxnK8XSpTlxSwyLI/nq7opwM2t81/9QWs9gHEg6vCbMCDqCKAjPGq
37gh4Bf0FiGBAK8DOEq/9LHHugIuPwM+ueNa4D2F/t2SekiEejlH4lfA9arVzrm3DOQZBdmGaTx/
7CMEOckMVsEhOIU5HNJKB8aP8ezr2JNakcN7AEi9ZF4GgIpmLrpWQoJTh2dLkmhXOr0Ox9Yd+wS8
ra6vqZpBowWFoe0mDnuJ0ooKR1Y+/cKNOsQOE7zyDgUHcQ2uLXTg6rTG20kIuA1V4/+tsBxdFNC9
JwGn8fGN/EwOl4ykgXvKimlE5cC/XZcaaoznuaP4PGilLNyQiesloZyoQVNsjZzy2XaWHyNWMIjb
N1ziLUmPwtC+wu0ZMInuUXGC/H7VUOBSdnXsTsosuWUpfeUCH244aHYIEexmj3sA50d/q7TIdwvB
YEAhR+2JieG8EXEwh6Gur1pHMs8kGupWCwtyH1xIlSzJJR+Oftdco1tw/EQ1VUuxF1ka7vX1tkpK
O3uckS8J2j1b5kN2REJzlKxAOUbXNBgnZP1J3jK4X9KOjTT/pLZ6LZbb9oyLvHCzUCHxoSR92uLl
HfHq0gS/RoFLA1zYM1BqK6VKPdoJ/DQfPiT2O1JA8X20KjfDunTNTTx4qKz0N76/QxtG1URWiN8F
p4ZKFNQh6l87oRCJF9xKMEakZpLvO7xGIxGKt4Q9n6OtAjuWJvl70MDGyaB9pGzv90EnHfVwawBU
4C758yEYnEa0hFg5ykk2JxKWuEJfFqA92DbjbD294oJBYANS/JGxnGd0GhAehIHIe3nXshZ9Jfja
lAUinALFyIqB5t14mh7ypKtID/urFfNaZ98kJJIOZGamdWzYOTN28iozzvsv1BFfcIRq24vnnbES
ve0v8+pNM1mFvOYcm1dIa0HUvlymYLnenxapisoT3cEl66J6pgUvpOBoJsRVahWI5JVr+X4Rqsv/
pbDZfEIiEiTV4ofCYAG4xRl0wxohNauPv8AtliXL1w96+KgzFsQO9SOjxhGX/fCgWW3qeFCRiNNy
JpGOBwFSc1+LNJhwGeMMhu3Qw5IDxiqHO5PITuMaJ3NEnLQC//Lh+JTiVWNbgILjSq99W1IlIY9g
RfjivFojMUxKQWzdCIKMH676TRZxakbyrwVmg86Lu7peXOFSPyjyRoGGuUDy2DZazQ1fZjKcjVCI
N0ZhinNTYailKAK+J+jUpF0/8jaZI5AovQ0Yi7CCByZ1lNJH1zz8P/5ypObbbK2HQcUh1f161P30
2IJxxLCM1O+IdoYbTKF1c3ohTAXkilRP8fnbe5hOm8zmJhxbuTu5WbWy1c4u5qz2Uj7JwXkVXwwU
6eqPODXZD5Tf++MPAS2xiriioaE2iw2wsrI7WZcZE7cJRTJfClzAA0zry79EmxnGEgqCb5iLdImO
exeJlRvf968PEEcnDzGZ0qDY+ebTueYykaKKYAo0ft1vLFu19Lp5ND+2QIm+ijAiDhoeV8qLN5+c
kVoiG9q+W/W7ar38c+6SJznujl1sVhFxFC5MVB4Kx/4OpttJq0PTY30mMoQMAABhuyPEqU4rMzOg
NVWhA3sTlPRpjUC/hH/VNMwByw8PV4u3rC/l4LnLpb7dRy5UjsDF/bSLQvcQG/MQwUfVfcvvGnvS
WdvaWBTqOifKIxXH8eTTTT+45mxqRDAoRd0LwAeWxIfksDlrz7ufrf9sJFM2V+nt1xgpcZ+IOjL1
EP18JSHETydcY4KnOfe3xc5+wo/BtMWE1G33DHWZ9nvkNC3ZiFousFnB2b6ONCjWnGp5GtFg0dVJ
dxrvm3YG/XA7QeOzAApDdgfaTRiWahMq8pg6JlqFsSr+aO5sin0NJMU6anA7F1cbJ0pkWKuQjdMx
mMyDQ04QPMh2jtIWS4UWXzsNoyd0SuRXwX22n+SWmNAbX8VDKpSu5RgYaBI/4L6VwnhVqlMiURz5
AdL9aGbTe3wSwn0XvXlt4V1GTEAhqSAmWk7aiiM5A9L3Pa2bVjNrl0uaCP8SmhTK4LbxPfkXJob/
Xt4hf+e4GDE7Ka9baqcxmZVYcL5HDi3CTE4jyrf5c+wT8w7+cyOC3WpsQpoX8bFfWgq7NDyuB8yA
QfUUnO0gcjVIf3/1mJwDxV26V7B2J3ppYJ5uEmSYveP1VUbfF1sdTI/7zqB4GRV4lF4a6uTztyaB
2raxvPCOwqG+8vrGKn1KWfOUj/K4hA3wrft1LFJBsRwHBstOGcR4T3Bxt38DZV34dF4JaWdJjMTY
CHfH+ub0jqpFZo7agLZ5kFrjjRJNECLIP9TNvZf39bNDZSyJgRJp+WE+FKWE/O+uo65THxrdEX6p
t93bsrjQmOrc1zSMOHQgwRXUmw2/IaxhS+rd0K6FYvQHPWira0yuA9HRggkxm9vw4Kp6FuAPXD0A
Nq2LuLtnUN6zATMO1bOe3LvOHttfAGArYwchzayLFRQYeQfzVxyJh61QZNcU0ChdHQeBQfBNjAx0
UWBG6sR/hr5IFL5rmC4846g77PuqJW7Y30D7TIxkBhQTIR+l5ouo9nythvaQ8dETTcTj4yPde4fh
Ih6E3cS8EM2z59jGbk+T3uL7BP/F3S/OLOm97e8gHklvrV8gLOJoZ2TzxJ++m+WAMWJbpBogRR7U
t4lazkWbYL4q+zNnZCAhZw6GtjtqwZi2w2YWPZFIPvco77DEppL+nkFWEFSGNy6A6NWd/Ipj8tjp
i5g80oV4fpDMJfZymOj/yPAmEKrf3hKbsjxFbxrMnLnYEuL0DxEHG1IYoOwO8r5wwHcoQG+TpFoO
Qb3kq7+rozVPD7CB7VEFOnql5GHVer5FQ6m5+4NjseG3ee3e0/JdhfdljK46/2uGErmXRNn2WC9/
NnTVBkL5hwYyzdO7daTQOx+eaF/KtMBnnyQCVZ4+lGVAGT7BByigx+GULkMGw9ixnCTy8PXbRHxV
0LUSpsVfYTilSPzCN/SccOvjnJt5X/bwI6XzabuWX29azEdnyOQ95YWJiI5mKLZ9WtEK1uZlr9vs
hOULT2WJK7YH/D7LO6ik4hWc9RNEbBBpBNjMhxwYDKJTcaaU1F3DVqMoZTikRZE/QbKch/rAtVsf
Wrt82Tv8esRwCph8rg4Hm2GLL6q4D4d8RBM7RyEMiSQbR9Go5e//9X/aTCG8766O62dshYNbMo77
jcohggieMKc74QhmxPxMEPBxFjCdf9R42N6mzuN7TTrrXEn0soQZj67Kq6/qkPldvBqP/2yj/TPn
8wwl6mbyWkp0fULD6BUgzvNOjhDyzeBh6AyaktOftCRtaNw2PqSEpCz4z5a9zK9NkAwV5yFZ5A+y
RnDENoGWVp0eSDpQO/SQmZzGWjdME8maooFglMoOzMJpaRXTXXXgoA9HgArdDTEijNsrwnKuDLhT
42RVbpJjZ+hzvkBxSM75qzDlXtxW4l6IGxUXqhPnOJrpsiMicUylBX4M/hDTG/fhUQXWBo9LEGSH
IRQPFvc54480Nhuf5OriA3T+dGtruUjOM6m94oHXg8ZOXcS7q7ADFckLj7ZkIj1VoXhsuTnf26H3
cLKP9XQi5rH1/PoGh/q8U+SJfjE9K6lchABfJEDtzWwYAqJsBgjz3zFkRHZ/o+2cy8E1Q0y3qS0t
u3c1+N5riiAl0lWBN9bj38Fy5+OfOlkTC2V2qUSMbGs82KAE2pb760FKe57I6YBtwnhRT1gRrEJP
kefQBaGZ1sV9Z+TiOlFn4daqOrTo3voVSBe1mshbSHbA6ViYKUctC0CuEKpp+hYSK2Jmm5R62+mw
8jdSzLX5MEyTd5PHs1x/QUjj0uHelORE3McNIsep1qC+iTeJ1Uz46pa3IrTv5YjKZzuQQOwqGVaj
sPJjEWTOY9vFuEcXDqvwdDn28ibeRaAtbyedarUsAaBa5AdWSuG4plpticCN9vYo6FOduhVBxn73
YmPpWaRv2hSGeH4dDjlHagg3p3ALoSrHuYNcrTK+xD7Dgrzi2DCTHj7i+z1fZaV4PI8qI3je8m5I
tIeMbHTGyE26Aj6XJf8KBAcM1iYhoXWcXW+xEehyS0VO4zc/r+OM5WbJLVti9MH5h1g0cPLZ9vyq
hXslfX2/7gp4WtB20HtcPv2PntsBoNXfr12lv7QV1T9PgeevQ/wpvFSa07qdFBPhHv44VYmvsisU
1RGXGqWIEWKRA34iex3NkWx8zphryq+zTIkRtjCPe5PSXlmkHCKFBoF5D6UVz+siKKzpnO2NesIg
OLBw+hiONz0BPKDlVIa6fHvU1xwXiFonio5N+1qz2PRhnIJJJpq/+wTSXJ2QH5PLpmw8GkKN9KxB
6Wpe4znsCiPpQgvidxFEWgc3lw+KNivZtJm0w/v61+S2u631IVU7j3TWnNnWnHOr78X0fsZpIvfe
QM8IAX+9bjC/BHeFbN7h6nD7Mkb7hM3VWALYeWrVYGwTe8jW1U79QwxHuZhtDurjT5bjdQWMTH3+
/YyY4Zvj0JR+92gyPfcQsCNJ9NyQ0CYOaKv/EVSx/zyDnkdtLbjnxFDv2TpJqOSfpLIz+GdJ8B6h
saTRIWGjyqu1fNzLQNchn1ecyk7Nf/cjDYD0yMXhf3tHsaBkM+DEHWdScWpYLJxjiMCZysQVmOYi
pGuL8LVDL2QLrKr77NWqzP37mv83MKX4EaoQAAB0X7GE+nI4lkwTD36HkFX8TTaLlSCw7CV/6+AU
XT4bF7sTGDI3+RE7qy4fXlve0VQM9uIp29jg1Qab8wbg5GmYQs05B66DizKNMxAgUJZrZU01z1Ug
D8w75aJPTc6RuToToc1jkAk2RqnGYNmsmX7pJseCE8R50eWsDjku0tLRwSsfocPQEq3FDxjGlnQl
c9BvwwTXO02AEDy+Szy84/37aiJT4WM3nmEnryW5zqSGvFV2tNZ1zvNB4W1adRykRXNzgdmn1+/c
FlTkUk+dNTm7Dug5D4n/bfHjnBbimiuultOPFgCTE4m4kZ24PDg0ry9QRqgKCJrylue0yWFaOhXl
MwD3CmfVCdHj/hoYoMFh42JHvkPHO3QCRWAQ3n8Gen6FCyv1ywwqJmI9dNKk2EnC+G5uq5fAGxTo
c09iOP0JDI5TZRgD/XImsFCrHKXNFjgb8CrW3kjiDjfoVB/eLfU/LeII4VLa5/eSRfvaawFoyViP
cbO4Q6fJq8gtFmtukL/CiCORnVWd3kIu96MvhLjYtIFR7F7uUK/Td2l6ujkwClUv7abxrAbhj7Am
p8t1b5dlTSNhSv+v3BBZT58rYaVtAryugM3JLPTgIaQeoZeY6VPC6foc9o2L9y09+ficEWsutFdq
qEJ/L0GnfhXwSZkNNoTevp4aAA5F3937SaqIrngQo6JWj+lgqPdQFGYitfSMQVwvCvvqgupeDExW
5+zCrmGI2/IyvvTEmLxOuSn12Kxfetqr5Te8qRBYNfRlhQvLK+T1OplqgmnvYQTZN076F6muk0EV
pftRHpTPG2yvLup1T8PlRUKXcCrCyQCNkSM7W2Cx+h3KxnQnWRuyhpwI3SzJdtHKOoHZof0+cN0w
ylXEXHIlEUJWfNj+kR10PujzH6h3i9wqVLPrTJ+e/t+M2/AOexH73VtsaPoIlCUS0cOrhaG24AGq
UgRL0/n5HjFuo6lbNqszk5S4xedKJqNbHfXUuQiu2d2cPJyr4j66W1hSCeXJh4tr80dYnh/a7OHB
3JUZ8K7XCEzj0kHp4Iw0pQfmBPFLERNk7lpoFWwSicMJKgwb0o1OUa5TtWLBUWt58zLhvsNgix4s
U/usFB2Xo7eswy7Q8CRNqqQqa8ij3C5pgbB0C5yv8MCeX83Y44gcu7xSZx/FB6ye0WSXC1Dq5FA5
rBqfAfs2Qjf6739VeDP4dcDVghsMfIh7+Qhy0933w00bRdO0oQhG80Z2xYQBjdzdI5Ys3OXtLx82
39B8XncfHWG6NwvxUc5pTfS5VuT0mBHneyoPyJ99HkfDnzI84Fkp1Po/abw05hU7feqDheD9Lv1q
MZ9w7/0R3zwtMKEqUZ98Q2FPVu9bpfKVBDdfUGOEU9DXbX2Ay19traeG+ChOH3EG5n9j2Y3H790T
eKW3B1Fyxtom1Orh5T4Ex2W4gkcuAxwsaS2LNlAvJQus/722JqfYhhEAKZuRzKSTbjmN1C3t73G8
nMut7wGAZz0NQB3FncBjNIAM4v4921Dmx4GZG60wSoP1fcbQ+6Fqp9UTK56+Irtf8MkrBkkKTKvN
PSLLBdQGuxEGxQWtdhjTmJ5Z7OP8SU2ghXyZQgYbyzBwWMGoauhMOfaoxRxptEbZ5NLqhBfGpEVC
+cAVXJJxjp+XHltdWKP99V/ECULVG9BKRXxy3MqNhLqAjA9JjfU5yD9oLCMiegGZsY2KT9jTNwUw
5XqxasaMiMVm2nCWI//qKKELtv85tUdPt1pRN55Of6OXDumncGUfAg1Yq0zzOT7iT4fixn7MOjzI
OaFmLnxs8qtCUHl78oOMy7bZMMFOPdyRliB6hzdgzLrw2UvZspYHolNrKULoHsutEQV2PY2bhoWu
njI8CaCFiu6orfJXlKVydzZYYxYX4EUKzqYNGE/Wb0a5RG71Kiy373feLeXZaKhxoGVxY4IZLpAj
EzMI+SEZurKATSUXfXdNpZylP9O4UAHaoVJ5hTX+6gR/sLvoPU1f2sjuj5AJtgG+TvM/1gJ8VPvM
bWHYoqrhw0v4cjquYJET1WJjzmbS/jlpWQI0sqS9ykOly9CrdiienK2LSMZJ1ginsCBQSpLygBnC
fNJ6HCztlbipC43T61B3HjPsF0Iwk3m0LqEURc5ED7WdYHaUqpOJtdvd1lXymmiHOhElEJ6mS+3D
GX+6jJ7qYiwhWm9Wp2b80K0DTFlrQmRxEZKBeeTgKpHMRV//M4ktgvCEGXIlOamw1pSqnBamQHmQ
IGShDsMk2XUus4UioYUUtzwpNQzKnCjeDA1Pcx4V5Ogq1SOOeIwLaJK6z6IUYBScDxAwsRDblYBa
aE+73G4C/7hfDGDMrhcTkVi6+BhwZR/ZK2B/zqZqcoOmsRtKYYPoG4y4IiYq/JaNIDrxqM3TZNBu
u+rmq4vcySBi/SNnGL3wTwCeh2sJSg+/cATMvW/ZRT0yJfz6f/IOAyi3sjyFb3aYwOMAovIVqF5m
yBbCmUSvssqARQNmspQwWARDdAzoXy27MPrYyHslXdfgyCFJPCjon3o3qDrWfzKR44S4kc+qoSGu
wvkB2WmEQ/FVtkAjfU/O7QiQx9Isrh7PuA2zw8t/E75CN6XFghBapWd/bWPuO86AmmGU23J3bOok
iKnNMCxDuA7arzbIOeH95SkZpzLNv/0JYI9FIzeyA6PMnUNARaDLl0cU8E9nITr76msbM1i0jSAq
dg/JWaz1phsmca87G+wT+GfumSoWvoBoaAncsf0cvHrEhBPz2g6tVLyjJw4vPaRDdrkQXJGfFs6O
dZj9tTVRKrG685Sudra9YRJpEMkKguBvJiqE8/LWUMQGSg9cPt0JitiyCEuxwliLilPXB0tykOLe
pnCuo4pwa3R9hw0rVt2g9eOwQ+HiUgf5D8pJZg1dWrRbLu99Iimq6ZxFUpuaNyQK7SlJ9ZSY0Ez2
9OCzqUdU6AdGodUHwnch0eCctqRIP84cGYYrluuA98uHN8eTnSw+k6c4eHTdkwwbtjfNAOs7mW29
iYrTuIpXOSjoTvedy5FrUgJcRo60TxzKNxrVxKajuNIskggdN2RXrkTMeucVfG5xKTCqzEAn90At
j2QXPjQGFGXG2Uafadr0ZgJCyJ0QhhkaNkIVxPmmAcw7pPeVziiIe6mASCf4EFd/P3BejRpu1LhX
r0eHt8Mri17rgehu4V1JWJfSmrCm+Ilz63Wh+tTUTFLZQ/+AFq3X9Mh58CtgB3vIIQQbwR+wgO9a
HHhTtmLngXM4nFsWreeCKvH8fyL2Qj/rIs5eVnTq3euvtMzVyld5/qGHHRfiHsROkt+dDKvuWGus
btv2ybBPe/UpaACIWTYhIPDbGfs2aS04SKwKYSBjQrhjPiniGXIJhZ+xx271PvICI5b/gqwW1Uri
EMCwSG626pjhbF8+FNWe3B/D67j+2ogF06buxXt5Ktv47yxPeYM6tN0C5oI4TxI1Rkfm5gqiZEuD
NFcVy7QotTc68fMDqQ0HVzh9sz4ZqYKChbb9MRg9XWqZWGJ5OxElNspb6Asvu4sGLIRej46FeIwL
Dn24z//+1pNirRB8z6tN1zJfla5t6JgjWnCJ6Sv9QgZY9Ak4IfN7y5if5RuQCrz5uT5l3XzeqaEx
nNm3If0y6v8bMR8YNDsQZKupClgAgdZVEvXWYQWOvKvRRM58RSThYVczwsiQIiYQrj93FWab/BN3
MFAbgtMvtXgHVhDmq4SGOW+h2IKux4701MDifa+lcFxLXzJXFXJEox1DKGPOYJIbLx21AkLDhnDa
5GEjhyAOUHKtPNumg52aVYJoIx8TBZUdxcxEoVPqBsaU8iue7K2qRmJ01JW3VF+PTJBnR4WHNbir
MwMhjjKARruztOIDrDlYV750bG/Rfwtnj3w+1sS8jDTHcHyvZ5GJ6/cJy7i6Xb62NA6UR738gbz+
o1ln2W0T19ZCgkuEtkIDEGGdffNUsRG07cwjYvdCm4AInPG/20AXn2KxJ5XswWuGvDH6bMROnr3h
XggJsYpBWINy7EclbKNHoprFIVgd5EdSIUAvQQWulgaRuJ/f6x2bkKgWYC7JmmnOnlgMX5ti2NI6
KFDQctxUx7CTEIfQsuSStSwSb3iL7VoHZ3CMpqjj2vHrhzFJXCngGCD+n1/YGdAYCQLmy5l6P90s
oaDbNP+bIEhaTbvPCU758+6ApAvEnYPs3yumvMCC/uPT0HfPzKelOY3urZGZPMhgeUQ2lRgmau14
La6PojjIRRCM50urNP4AehNyzQu96iaakNMAydjB8xWnrMlF5dKFEA3B+N2H2bKmPThar8y1PJ+v
uDIha4snWP2CncNTxQLFaURmbOMJAQk9Ppoc0gn8jBSoA2E5Z1kLxEA45lOLCShKR6CmDaF0/rW3
fnGKsMc7s4DeNM13s4Tj8kZVtAPGwO8AutmuC3Lw7d4ajPkdHfX1ojKa6p8b1AEG5gDG1h5iX5ou
78VDaUkdomjbUQVkmR/KcQ7I7avhPKvsd9XbTlhph/LQ+Kz8hPdkBsv7E9FHOYmnNvedhJ+n37+L
axfyRpLDGQYGRUb8BFQHegVa2oSjw5q5igpCLYaH4z3DeZ8qNen/nB3ceK7R5IFU4NFy8sTgkojd
o72+m2MhesuScf7KhaqrHpwaT/iFuedjwL9JdHz9wcOzP3i8jWE78r6+C8hXF/Y/ECad753nMJzW
KHGqz7UdaOq4IsTehC6wfME17PAm0ti8XTmkuoCbOJrvMw33HyHrYtIuEyk3Xf7w0BxGM04bTemF
hzhE/QqfeYj86IfPQoAi8Ctuxye5HSbaFUXVtswoUgJWyGf8iL89AazXcU5GWgnOH8TDCsJNrvJb
WWUdxZIQbIc/GiSIU2l/AgwYgF9sHeFVDOeRakj+SggH38yiTw/aq/SoK4Zc2jHz6/me2fb4rPim
f2ADSVm7VMMfbmEu8fTPzRx7DLHEa0YcRgRqSG+tol74gW4f/k0EfMyhwblRCqsAekBl886L/gg0
wfm6HT9pJbwfuXqkL13FusGDpiLbw/0+EywA2Nq+BPckfgviXq8lLGgxnThkmiTT/fyOmK+P/7WK
SRJ/hGulAE5ET7cHVhH2Yjin/8F6P18nQg5fu7J2OX2M1UN6l0ekS0HDh5ORnVhwDtpPcX1qXX6b
FZP+3H/msKCI/Bk0XsBsWjyHxcCaBvuKawLh2DMygqi01KVX6uKT2Kgzjk8jBZRyGsUfbIiPiMdh
j/SYqdFNfguM34gExuclbpe5erUiVKq6OEa4efaqrV+oRYldaCpCvYd+jrF81IiHJ6GaIHtt5/lk
Bd2Rca6Nwh+4Z9Pk+HkuJf9y3a/kNcESVB9javEkknIob85lA+fVTufZTWSbXdTJ6DoMuTroyWXf
mCC1Llwe/GoOxLEEwEG7Dxj7Q+iMq/zwE5gXjSFc1uKe3FUd1iJSohx0iKDFa3RYQP5Tn7fl1l1u
O7cNVBBFriza/563DgMFw8Zc6B84Sf2ULvfsDdC7MSAIcHsnARXgVk2N+zaMlzNBE1WztHSC3wJ2
HwA05dToP9EwNe7cqyfMI+qFd9ilJFB2Ot/HlFWOPCRUYGgQte1B1/RaivFO1ZXDgFghBkQNhQs9
KT832M5oSqtKn0ZVwtyDHAiD2l9+cGVN4xLjv+eyluyncKIz/JMajCffHkBEpoPErW4BlKOVeKlh
iDWHVwL0se3daoxOi+fbREVtN8asD9KgE7LR/voPIaGoRDIf7aPPf7SUessye465tCoWyRjBk/9K
t7cDHWQnG2caU+Zmh8khyoDq6Vn2ScyUhIpD7NReWxHNX49oyctX6iFUo4HQiTy7+WuCVOohVB1K
PkoqG2dyVsC7/p1KkIOKk8BEdItCVxd3/nkgle/mWEd8hZn7mh6WeWJS/pXHKWZiV25L7xL0/waB
bBnKf6eQ0GIHE5zIgnvU1O6lLPvI7OAt+6FMlbKnssPNAQAdZT3we4J8hGaefLfNGg7YJNtLVizM
aQJvJCQA+EUt66TdWUydUBmyp8qkro2QLMNT7c937sVyO8cVkVYE7qGOE05cF4S4D8HcUtaiaH1b
wiPae4J11PY/FC4UqABZaqndiyzezLIx8HkwokURnQS2PcenpF+UgsDpoE5dMHKiNJEWSN826W+S
vbW2zV8uxEfOPXqszBTlgx1FNOAEYTf3HQyPi77IWukx6y2U+txMCAamzgw4cMNvFtBVQCNzvjzr
4ovMy2hCUFkQ5ElaOzBWS4R+5uKOSIjnY3IfUx83lclTrPjW40JN+kwNZPzojjAgIP5VhOtdtHRU
W1E2TehPhKh03vVWXVACG+hLF2sPsOriATMs2WU0Mj0XLi+DKFXwK7MFXxOWj9DmvliWEpDJCuuu
jwEjjgsfauosY+REmkZhPHt57Ofe2x2aufHjabXz9gpf2jfnuPP9f/Hhkv21/G4EaZPWaehf44pH
937Q1t3ij6ypzBde5BYgCpCyxwqhkMf3lzUILSvZgXzPVHqo4lSQjJrFonvGUdK09yqDyelWNMxP
vc/99uDOpmj9kLdqIaSSyhu+06m5gXt7PE95yHrYqGHGIUaSqtgr8U+KguhIRO8Z3jKeScfhz3qR
BO8SW1EnDmDmWoJoMlghbDrWro0FJzcrekKUp7s+FRxjNJlNfp+/98wxHA+m93saE5GVt8qiIJNR
T3IbBkaGhN0pag066IRqaeHgTDwOVkVVsIuNoxyoiUZuhbfTyodekLvGddPye4XYaf2qheDcD8uj
sOvLP33aV8b8TRYhEHPBD88ly3vKxHs43VrvrhBwGqf5FDPnRsW0vjegvFH06NJ+swJEGvj0OWMW
hckuBDteVEtbWUBg6mMAx4b/1AX0M0rkm29g/zcJzhFAgmAqF9jgbIUAgqMrn+Q57K4Yr8hkk+jh
cOWFi9f1KbIV1PzSqkCOKTxa/IX5tz2VJwLXmUlexjj3aJ78ILVO2625YntYwjlbfP7nmXwA2qu2
hyFNa+Bb/fe0AOJRLgdndfRK/fJCTM8DQ5hXOYp1T88t182gDJn1Slxy5KGko9tzooi3uIm0/CsW
Jt+wHaDuFtACH1KXKd6cZ3ApguR9fGiAsN9wLAjLTd2vYeagGtXGZw0NhE4VJdqmWYUP9qA8APfV
k5FiOPWktEmREPYdiLugQYGRzPW5RVKJ5xXeJPxC+k2575pgyaqdjfgw4AMnOUtJ6DK7DZha7Ba9
qpGesfBefnWdKCWWBvuUaXNbVkeyOH73ZMakE2VL7LgJ8rgs2IOKB74BihRbUXiIZ/Prt+wYWQ/P
k4u0AQBUx7qQI7FyPDAIsd3Ni8cUUBEU3SJNwqzsPHp9zs4YHGdFIkINf6eH6GwEDh4XDSHFrEwZ
yXR0Oj2SRpAWDaZtd2Jq+y/xY6McyZeBXgHihnP+upeMc9Romi4Ira8uqPWsOjdsLRYqUUtyNznU
uAXXjiINUvIBD3k0qA3qD1EqnWWR8jBlOEPFz2AGlnYQBcyZFonb/K7suOp+aWhlgzNGS/v/st6Q
gm3CGf4njae8dIKRbwnoSEtQOib5CcXo1c+l/LnE/sNfIk9KJaIBgZ1t829tzR7o4+4j+b8pjR42
LHvhzSJB1/Skhey3r3wwcFXGnbYTnTkM36T8KWkOoWIhRE9dhkZuAFlTcd3ik1ZBk5yxjd/xH3ZJ
Vs0/Vc7Ai5nTnfuCh7wPlBLUfitUyu2ATqcUywWkqRsgRqr7kxARiZw7ZfXT3G207B2btjX2l2rY
WO8AERdxii9K3f/BlJVaksVBgUq20gLOAHMJfkIgLDpIS+9MnmC1B6pAqsFfQMsxSaVsxz6vJsTS
IwMC2rGgQ1nCm2kg+AGFAt2T8CH9x2s1zMBi/29WRyMRiZJeB2PlXGpLkswRjbucwjQFHOzwXkok
KJuTpOyOSx4omN7ZeKbLSmDfHvfXqaPpfFEjaIZLx9i2x9kzS6xDo3ciUN9OYc/gG104zqdQkWbX
42C1wth7mf2ubecNw5tK70XSr85VAL3mfosG3FxetXH7gxE+brOhsPG8+fprmB7gWTzOEPmR05tp
+jSEgdNt0RBOc2yIZAkSYOaHsb7E714VADXDv1DlOtvVmyC/LEM+kAt34nP6sZI/APlNXvqC5wG1
XqsVUR9b4+LMJ9WA0GUZt7Zk72hGEXf/BQctlLdEcj/nq88bWhxk+FDh50dHyFEsFNjtu2YO8Q3m
vxZEO6hg6lYJtjXcAEKf4b9bKGJhUsGtpHzDszI2x53MoXgm62kn7xY74Z0CpjvxCCRveXSW/TN5
+7qm9GLy90aIbZYMr9hOk4LVRBkHvJe/2MSRzMiKpM/0XF/4xJ5cDeYL+eyWvbZh5/dnzhuAqfgM
gcpwsPJeBFGIePrkpLoiF46A+297VZbrvJ4NCpNRjHOgKY+UVb/6reF7vLkzkq3A7vMugGDDW25+
Wyk+5jwd40daHd5g7peoQLOAnUyem3uN9c3qC83SLXckjwaCLDlWoOQE/z//BMqjQi6CWyduTTFT
4pk3p+/kd1KUAjcV1ypQAO697upCG+fDY79wBH9MVKyGvC+UlGoKrFD+pVJLEn1+BQhVENEq6E6I
vGjWxzuKFSU6PIvialNuqJUU9ofXkR9j9fB0W0W7J9WfcPq6fq7grlu6I0CWVdI7v+qc8QVNph2v
UIReIDQw1mkbpgaGabvDLZyF5vvJU81AwITR0fDB/W8Oru8y22/+Dmgr9j5CPU9UZdxsvNqH9sDa
3N00KmLohcKhICfAMLeCCJQhACM0VOlfpbh74DKnN6hbvfF0sHJv5PU0JTd2PAx26Z4QqmWahaNM
MhQG6ZnQHaN133rAAGfto6/+2s4JuOKfYaEMBUxM0ad94P3YGMyzKll8m02CpoXrk4Cy7u8+WJvx
CUbDIZj1g4Z8+qRrZnW9hKlrxZNvaGOB7gEMWCSt2W2dIacmv9tUJovnCsHdVqpJy7OmDxqwfY7n
+ZDoUTc3K6q4ANXlcQbURNYW+XtF5mKFUqUy3q8cXF+z2+uCd3W3Cr+KLeiG3w7i/8XTYxHg0gKv
0qJHSoOY2nPif7fgeQ33uXw1GrUH2v6XIof+xXVfiKBSGoqiiDYUpSxksBLP9ALLZygiHbxZiax6
7sAQ1nTTeYcslgk/ApU040eP7DpfFMVP4dQTaXjFFWpJWEzbWQy2UQGHclsGpjmYgT1JgABcMhzq
cfX3QQQIQGn2VkIatCy8AYjQ5T1236uta7DvQDJ7tbhPL2DZkFzLG1EGXmOTiPgtpxW/JM3tsHvd
IJiDWURoso/y47expC3PyttWiu0tgptWfAeO+l+5nRPv/NgeGoln2+90u7Rj66ONvUKaVIeLnaFA
j5PLnhjaucRLmYUrNFrEDoVoxbaQGUEqaGjDhg3DjehcHdYu4DOPInnJhTfXrnMWsZp1ocom4vAQ
/5+3TKqX6Sj/HDEdJeZxl0S1sPRHkskzjJJ0fdBwUeC2y7OB/G6LhA72FF5M8+HpgrX46UrAs+eR
r2Cl5Cn2kDgl7Mgon0EYcEq0u7rRjtsx/cfQ8tGTz3pPhLsjFs7P0oqF7mZbXIte22E8cmZnXnC1
Yw80c5Ep7yNeZirEuTEm2yq4B8VuMU+hwrEoiOOURlX1CLs47z3W/eg3Oe1n+lFO3DDsAJr4YkmQ
LoelOqAieB1CbX4hpek4l/brNjf+XWvzKjKrgGqGnTDPCnBe9Rvmuo+FhIifnFq9uBy4aUZbhcOE
Al+Kv1w9o1x4uXPw85cq4A0SWQHXp2utVLA9g+oXwh5JEJkYL44Tpbe/ECgO5Cpl/s6B9cm0Yd6D
h36Tb/iKXdb3muKKVOO933QCWyAV5pBv0wre88ldZIEIUF7HPAgvXkPiEI5WUccm2FGxxNRuOh//
UvDdDtp4dZQbdBMunRbKLd2v2D4rtUhrScE3GRmgOBYITN7X6KAr3uRWqcl1jlDrECtT7LqAxGkM
n66WX8so96+m0Jq7h+ffZ+xFSUyn+DiK0zO04k3gXpEAy1RCcuvONtfYdzkvvtpmkHLsV9TFlRqw
AGBuFkWkvUShNmi4DtSdQi6bEvIYZjVqGgS+tFhGrfdvwgg/MkqlKj8qTHImW7fkp8QlXbkn0KHA
H+A9E9OA1bjeCV9GShT0URDrvqNfe4HQ5OyfShZpX1ZX8o5oRBesKnvUIjOlNN0w8LCSWQLlV+qR
IdzcFg+6oemTU7DZcaojU6cEJHapfKPSeMlOR6PwfIrIH1laNwdd15rZwzzQR/Vysba5WWAWr83M
PY8EjztTRXrgkCe9L9fpCbLcF/W463G74BVhfKkU89R5L7BUVaigb4ix2cwJLlRmI8Bdw4L4h2ha
pLao2zDD8JNFAHyB0aAsbr8cmWoGGO5iffc5YCvP/AraPAYAm6EpaLleXFaHadG6pYx6mnNCYu1J
IrjkXoQS+V/y6PfOX02ms5xcgqWzQCmp5Nbgujo4c75+yv1HE1jerSlAkmIRwyk5sqD0sVoeiz15
BYh+Nol4DU2+ldY/hmciJ/Co81w8f24MJKfG2vTfmIHxVg42yL/8y2VXSsnutmpnY4aDKlNs7bxn
dIIX3Ak99UT1gaRLfT0Ajj4nJzulvKK4/nYH2MtLzjFu7xzxoRGf9tzPTUvGlIhvAf+C4yVk35kN
RR27uzzlBDiefn/MciAJBjkS0MFfX8YVH0AIO0v/m+5/Po3VtDIfltas3RF+1ICkGvmFZqVNEI86
b49uKJdgFfv/aM51fMvxYOKldW/Mp2qBU6omFwozFqEUdaYOXnTPNjps5WUvLyDFjcxjdo/2RGUg
6atp7MetZSB/5wxFbd4ZU80Wu3SzHvQ2ib275oO3vjbX3Nur/KAVb2rD0YU8r7uzjsmwaQHx1gFN
Qnd1MRoYaYLLxhiEFgHXhurhPvaK68Go4kPyOU18lw4ea3YzhTE7et+2xUwmdgUeOJtEXiJGIfj/
QklBfdUnSNgKpOHAKYsdUyyYa/dgJCnsMGXgVNc5tXHXjnglKqTqJvCVi/6ZaPzEzdH4Bw64x/IG
PnOZMHc+aK/fo5Xc3LP54cYNoAulczJNfuaAQp+0S4cHxHEMwkEq48XmyafqWnEHxmNbVkkbPXhE
k0orqGm2TdTDxtt2uVArS1tDsbwEU3eKgvEybi0JVa/wKeZdrDOQgvnabYjRhr9aCeFK93R9u3k7
EiGlvAQHhaNelyWwChfRqGnibC0kTFlUosWIBtZhwOoEJoQdwkl+gam5kefzMK/4E9FXLi5plijc
rmwMbE3OBAgfzACDGtzA8TqOpH7v36zhpQeKTeqTA+z2fuhbGgFvJN8fuuvfU27+EVMmJUOoUhQU
8/n86H4BlaIIpPA2iDFhQfNjmQmNMZlSA/64aRr2PEziRX0rI50K52VUv+OIZlvXIl9xMcYrUU2E
VX62exKRKLccK7aEiKkjgwxHoqBFHwLwIY/W52Qngosb6Ev6BVJC87y2UFlgHWC6oAYTo+BzG4at
ua6x47jPWNfO0SZ8aUQRjtLmEF320RTc0oKvQjrS/BEdBPA8cRVlrIMsMvptugbuRqxWnmK/Yf89
NGMSwTzXyQs3dhkNPXv0uW4inD454xBB14LpOte5L8M8Fc509oMa0amRGjGj0hnn5fGjFhgQwDZX
61lVNPRJHUgUyEDADFXHLOF2jxX2wOiAIftyLrFfk3Tq0vE+sNzt2QiUM2QEvlc0rpHSs9KkEe/2
gPEATk9Qgh5QT7HThMSlMwAY1br8TlW5RUtahaf270ReYsRbpEE376qHchtY8k0RDYlokheLbxJX
fSb3K2z6HIq6cSPrb3NIEszFz1uCK6iXJhq4O90S5CiCk86sh0b2EesZ/ebbPL7iBkBw5pOn5IlB
vcLsaQx1bNdYI65NNMTP1cQL5DXwijkpNaCNXmS5Jyd2Twr5YjZcVTJ1wbwPXoJE/GdUEMEEL5hI
rGIIeU/aPqNMFqCY3LpmkO2nflpzCuun8GE0s5Z8gzUUDeIzbvoKt1TEEG1AL1T4AJisgWdCu82G
M8uuMZPwFbltxSG3HmC19OxJjvxN0L5hwexRkOeEyyL9PxQwwUbtxVGGpNZ7pzMWRgMMzWiVjpDu
zDHpq9epu83jn8FzkJzRCeSeqsn10VGIZusXI+j8bHb4JxcSbdQeyAhEHy+BPAeXlf7RWTIDwla+
MZLaU0tk8QpyfOvIbxkgtsC8oaVbpYbeR4BuN7i/OEPjj63s5lbkuhciCmav0wjtgf+qdAjsCDfj
lWyty4uR/wybbEnQzn3vrEGYS3CDSu71R1EvLaLYqM850jyt/5/VgdojJolovHzL71wOKLhAboVO
lLn7S+jbR4HBjacTyHy7+EdHllB0WmEnp2QgElhxI7fxcJ4VVyskfVFuu5qCylDdvNb2dwUAjoAu
OKePsXPAqJ4hgRR69ta8ina6tBifrE5l5w4hPjM9Kbj42cKUkKqiW90R3iP0I7vXNr0biTfIBZzf
oN9tOhBFl3O5Jk2tLVOyg8Ps74CR0P/IVYzaDNJeyQ6TBO1rYr3Dy++IjGzCWXs5t81mr2LOY5c9
lpQRqypjjY0VoCTEy6t2HEMH0b+PUz8opADK2cLrHh7SOXOrWkREg13WaVMIzAn9ECDYI5MrfDar
SsUiO5RDhHMVxYhv6hfVZeSwGQLlgMUv8K6KUvEKwidgxIBD5hcLk+K/UNXghSk5LemPLI5H7yj9
LlXeu2KPhDk8SnXpsmXZQIfpjoMhpXGM7dr5akYrllVL6+CKXde5VRgI9tKaXxbNYdue9LPlt+op
icCvR2O7E8ieEamf9IoO/RHH5dNQQMaBAx9cN9pikL65vg5z6R3xTbIj0dAj5XTp37PCUzg8Izid
ZLKVgIvBryD99w7RrT31gUajrzCtuOWF6rTC5pmyiFwDTd213yEYU+bW+vbu7KhxWCDiX41Zyqpb
pkzdZ3bvRCOxn2gMFjfOIz43leeIppVKJQ10P6MXL4i4eU6V6cWjk9PeWl0ogMa6zlQU8GlAmYdE
lEfwdOq8aaZFGcQHEcULL21b3yXqhKbGMSeXxqWzBXnG7F8ohmAX3ECTMkXMsj6+sYMbCB4HV2GG
C2fcq/EmLZgsAVI0gJ2m702WBuGaSk2asBQl3LV1bgRAbdvOm0NtCWsKnqQagA898N7Od/6Rv4Sa
CAjUaW5j99td7AA3ITx57qRhC9fc017aBHpWRF4XftFXWj3TcKp1hRSPXGMqdutPT8MESFYekwH0
YQJPPd7piNG7kTQwpW39k2YBi/+gEe3Bg8Urpti7BqeH7hrXGAVndWG+hubIYNjQ6B47gvzSaOBB
3eR5huV9eCKGWAX9nMyJBqyW5f4RGPPnVHOZKN4gHwmWZVtExpbkUZMV5AEg+/UCti+nakkqmfnB
m+9FRYH4Eb3Y0qiY26lrZSSm3Rd4Iv4436jMW90ymasJnhMoY3mxuGTY1GCpnI3qVyVq55IqUcqn
uRDNM1lf1paZGB5GYjfghRBLi+4dwgIUEFXIW+9jjNpy+Y1t4fGf9F7rcijRIY97hbZFXyC+dgYI
vVYg9CxY9YaQIenqxDbeAYYHCP2C4s2zWPkl6TRO/X2Kg28gOxfKK+FmOOCk63gMY0kvYbFihEmY
LtLvZ3BuEBmMtpaDeURIQ0RWLLfdUt6LYqDypCNqdGeFmcDCub7jauugtC2EJ/QuHRbCrXRWWD28
UC75plBSiNV3cqYBoU6Yof1H0nN8HkaeQouqgXE8H3vYV1vjGQDBWWQ/NJ770xi+vHWSO/9ElUry
whkH4i/a15ZpV/Nhz7CCkGesQ2e0jeS5VtQF1/ZO9GpsB46JLtFYJE5v4qk3x0GXrKDDjrMAO+fl
UNfwalkgqhjRBVTG3P6ocvR2xpkbFzD4H8/MYLEh9i+rqGr5L63svz52ksE86oJeTJmDiCb/vqFx
1LWNk8CeL2GFJWqWJpKYvA6wLQ0W1i5XM0hlh4clweWSx9yW6hmX+wGcN0iC62Y6y/UGH0tonuFm
DfqynLAaL9LWx3fkgDwCSOPfYZKmukOjXR70uNMDE4unTUG2+CBBvHlgwiA1ZDtk0Uw6tU0bDvh1
+WFDP/6H+yL+C6LlPY3hJdKyqcxH8ZZK1wYAaXb9LcDhWB4ta/1tYte7At+8Apu9wvqXzM/tCBdq
hspLGQgB4BtFtz4ZIN1dGV9ihtU0GpDD2YlPNg/KObxiOrdxAvXxQbOufosV2FEmF2Qt593UkUBm
dH06cJELt8zRuhne4LtPi7C8Imh/do9sMGSJ0DzW0PIKZSqatx7dUWFTKYfLSnsOxKm6KZbEw79U
yTq83+NF0rGeSO0aYDZQMzkYlPCfmhyE5twGt+/zoJZRAhELN9/NZ4IJykHUSPK182m8Q0STJkay
lkR5MYpyMxcsBJXcJRv5ixhJf/ttKa0B3jE0WI0KFoqNutEUkVZTKEpDP3ele2jhdJxRRKkBpJah
Y9CNSd6vXKUHlK5zR+dtkzLahpceOiG7gq83NPoLBeb/XS0nm3YBCBvim4o1bBeNolvkDRrDDHKe
zhvk7uC1BzjlxwsNlrrIjIVragCaDbuVT3AwO93My1veXGUR/og5fGBCnBR870KnoVGu0rkL5ChB
sAiSg4OOUnzEFSqN3lurxFCZWvXndDBDD+ilJWIHmbpSuYSPccQTZ+l2cFqqvVw/2ZZMuJ4VWgv/
gX//Q4gOtxZTsZGp9Lorq0cFaPV2uKCbD58xYRBxYYLnONhRW+BxX09BIGkFISQ4+d5+6uD1CeSM
Owu/G6ssaqaJWo8gTKjxh0cPTJHlC+7v8dxo8J9xLzmQScPMM187yeMu2u53ek078WagdEJ0G375
q/fEAxjw4z1eb248d/NTa7bFsWwqA8qRJHLxYAdM6ZH9lhgob2wCzX0Idx5DdHGf8KyNSGrYZE8a
OB5KEVl5EaznTTrC2Nf+fF2bkNi+M2f9bMH4KpQaPisUQnLavRRvLCGpsWPlg68Rpm6wtidi9b6S
07OY3FHjZdJG6YFa+WxErOtDtAXiC4UlKqvVH403S+F2U8wXw/eSFhhRXDDzkhh/fmOdd3amzrtW
rjJ+xduL0onHc1Z+qmQqitAeScFv63PLElmGuPn70VwarDw2tofr3rmP937orLArtHlpTFrXWG2W
hpub4x1eRAjFrmH3O6yM0lAOpkCbFkzCRkxjM4DJ4jTiEC8On8w/ul1HH0Ih/NzLObMRFiK8g79E
SisOBOKwX9IM6euMfa7ShKymEIdG+ttqGFouzRuU7IG+lQEJp0u2F8+HYAo7BCIXJUtnNntifnRe
YSsGVqdpjbrtqyROEfpMKk/wx9NCXxidcOmsvzVkeLkMKHym4t5GFgQ4BXk19/GUzBsMSRWtoWY1
ZJvLfADDC/GmlAhh3wnYeFOLd+kRe3yn8Zt9RshT4n+D6CBolJkwkuw5r+rpQdbOb+3oswIKmZwh
RXkkKiuyeX2Vk48Fmiuu8PahKjFvZp1tll4B88pNnf44+TRhwy5KPrdPkp2HbnS6IXMSuDNx88xe
n1x/ouQAXddmbEyZYrAry1qPad3od/ocAXVvF4uj2EpUUP/YOqtLntyosqfFBYW6Tls7ML8id2l6
8QbDbHsWf9mH2bYDdBruZ1+iNF3qjxLwOVS0kBw7vfQFPbEi+J9csy/9y/V5KrHyr9dMQ2LJ3G4K
Bswmea6GPI428yChnbzcYRDfJWmVoKToOdzOsTjAzkLSrz8SNiHSP+obhXCfDvxmx5j5AileV1B2
SmHCOg3RoqVwz2FYIvDWiila+dM5S5S+B5tZ0cicUucQu/EB4q9a8IBfAQm/jxXcAEbphoRjIA6n
xyEqc6iBuYnD2i8xjT3+TuV95bFvmtQCsEfsYsg2q798+FLuMZBoDhozjfdUSFZleo9A/QOCCIuf
gkxCacv/2hWIibJfUXD7e86r2qbC9WheK/Jy5OkCSyp1QgAaZO5NOS7nU67x9YrWYchzsfiBYiti
tjjheit4aB3Se60ddJVdxpPyh0DHXXyjMo4HYevQxrozozbS2pW7opRiWf/nMelsSn6g3qNUWMwj
PPVOopD7Guyo3YnXZDUNfRDZ0DlpEh8ZsaxfiRzF3Nav26L8h+OYtYROyHn4sdeQBgOaYnFgyHF+
dMYi+KE3SZXSWYQxn7FJMjs14rCqJ+A9SumiB58uohjZk5rPFOpsQwiNhpyLclcM9FZxVp1sdjo1
e69Cv2nZYtNqVMEE6ZHDBTyNKSWetquRaImvIvK+lgbv1cav9Xeu4fn/m4et/NmAQToZsC0hscW8
SlWd6Z3ocO1TyeCGCiiIx9XzZxc/sKvR5gK6tm43JHRp6ITEU3NS6tp1PBb6zJrvY8JzZbolO+0X
gdLW1ykovZMxOfuLNdwhwpGkYzoLuWgXCC4D8KTHU44knb0myu3KhMLUIU+0fKvUR8/gvs1YNOUX
J5/9QMIKV7ze3XsCV9kJHHqbWwAlCGQ/oWaJnzcg4et25P1wnP5DlMAdaANthex1rVmerx2poc/S
7ndGCLpPb2ZFiC0T+8BU8Wv+2MVK77lX/3Ab6e6SpoBNbvShe/c6Jdy7zcdUSL3OS8UvkcMYPwCz
lA6US0WpYQqtEzcKEozZo+brqipmsLx7BRVrPE8cDeMWPU2STIa//Xon7KXSTBYKSEFi2MN8cToq
VL1neoX3/zh/y1BEQLAv/u8HDS+Lgf8Hb9b4FhJc/4DiGurh49z4iDE0WsHzgAn1N00Lx6HsTQSn
ucPmtSF3Vn/I5sHtiBkSiXtmzF0GjiOJ9/MjJZV85smpThPbMXmf3RfgthioMsdRfcFoYvZWqURh
9/fFJVUvXuKaudLAoK7sAff+/O2RV4OIuyJFV35ahS9nlHGXI0lMapBL9XyU6ZCsk+mTTBKQnf0e
o4AdHwx2wzjVcObItH3x5qWmwAUpNUE0Xa2YZhacSqVJSrgZ6hAu5soRrJYBouFoXw6ixsQb95pS
Arkb4hgkfoyyZBQjeapcttMVi17Re1GrKAPwLOdUMQ+zH/bLmphznvpv2Y/AdxwLhdBe3ILovy/B
F7puGZN2iAO17T8eDa8xxjQYAOxGqfPBGLdOuG64gSsZxLHY+7R8V6movL+QNCgnnyJfCVoCNwZX
0mqIDIJpZBHgkVfFf6jNEfmjDQbAqSq/tZRz9/fEiwdY33/8fmMtK8vAKWLNjmGrOwZjQKF7fliB
G7sazJp9CS85LRCCnpM55FJSBgODA4m/3QE2a/mMhqGhcitZOXeCVwmYpiAMSpkBgkd0jt5YQqNM
+C1rJM0lwqZUgSh9fOpqe3oi7s6GFH7a0CJByQTQNvdir31aVVw5Q+/I55XEWOLLww/H/ZoKdplV
MFXvWIL63VgACdsjUxNTarmKyrjdtlKXoju/oBXb6UH4ykmljTJCfZ9dDnzkDjjuxo/m5U2qhVQ4
SbovFJezyw7i23q1C9mysf6v3gR3aS40kmI2g4zS4yoVnZWOreXeDfbAc5tiOjqc+BbToXTeJbCg
kE1O+c48X8/eDK2m4CyAmhslhTt80DZrbIZBFQ8nIqrpxXOxTcj65m33tOXKIEDihP3PuPOfC+Bw
b4brSwpz6NBwTVCF/c/LwKtysNLiXZDAmC/G7y9S5kGIam6fTqraOFUX1qQFsD8p3iZjA69mcijY
xI4UlU9pB6Os7NdTJQXjRccXiUgsO9URchpTtWJsCpYNAskCZYaokPYzkf/AHY3egJ7OXnlnVpaz
FukKX3eKviNEIKJfSsFmt2WaNXaJGPAEwUIx9Xt+Nwr4I9Mm0a3GoAvK7jXNAfTM5lOqgamQ9Xsw
mMks3xsNGHQdR0N3TBFwRT3O7sXBGZNptr26BVWV+eUqQxNv4nvPFre11Tb967ye+ird3e14xH4N
0iemmG7hM6UQ52B2EOf5mxR4oL6lcbSUIhvGRrZDwq9QVyq1YaIpZZLzlxV/FPGTPnX8oqWnPzA9
XLOVNw4BkWU2OxEyWOmq0/rm+/PYt8/vlvzNO+dsgD+W1ullLrPZkT9M02vPVYiXgW5w702vI/Bi
aZ1IViKS3JOKEF8AfiJSS7VqpDm0LoFY2dt/RE7/LzlqvUdS0J6IzFE07iHm7BE5SZNjwX4+PfQc
WxSoEK7d2IyEvSGzW+qUgp9EIS1rNUyPkNwvMlSY1peDapi48li5mw8qYBqkzy9yu7OTDjy+3fZ0
fIYrNLqy1HAXmQy3WoXphwUGGZU+CM9EfqyPQiTePU3giJcZ54+PRFoNv+iImVSUSpV0BCcXdOnr
xCdv9513iZEfokSsyEavjG8bct52mmcpyospipRAVlgnq4FO/OxzHh0p1YFhlZbfo7sPw8u5kKvZ
GNFd3BZ/G02IHErO40MeZGomZw+NGVXvZ9pXV0hUyzykuq/4xXRyREvnGRhCFw3uKobahJwHFOJj
Gh8U70hW/bn7nDV048ChSHeHsTfJCMUm7GV/1/DaIVWgowdiwj96G1cjOviaSGyX/hL/Oyn5hfud
0d7a5G8lzjv+avIsnDEdQKqRw5yEESENkljXpJaSPPqkaYbLnzjBsNHyNa25LN2e99o8Vwv2pn6r
UQdGnjbRRXUfwZc7wltibhkIcnD5kN8hCz1HdX2WD30od8s2vqTmnWWsbhkK/XRuT30WacF7/5U2
Oh45WPSpBwV6nQUf01jKLCoMppVVof4ZPJbKlwOSQrYvIBDhYF2DnFi23G7QHG8nKFlCxNEhon4J
9jeIU3unCk4E5h3Le7Jp4c4w284HUQAQWICAjpDPsi8lM0punJGOL7lSDkGnvGxg54lkPG4h95hu
4q0mP/VH258xvvI8DOzvlzOZEQeKy7inB8YadpqrkUnHRSvrldnIAe7uBSSVboWFF7sqnuzMcjz1
DbJJWs/KxaH019XHpnCFMjSbmx4NLpb2Pq+XVXD1Mzd1BdaOA53NJxkT0iOPViOT5Z6Ca2M/KXqg
8Hh2le7QX35gX1ZgFxdhG+2UHs3lGNrMuh12JjffSHqGeBZbniEzAqe9BPTtJ8DonKZMWMp6JN7y
U+gfFo+u8g6sOr3Pfyu47WdaM9luCYEP/pf4h/RMDpk2VOe31/ywWr6J7rQiT1rp1ccJaYC0SAo2
z+5c9leKWqXwohzpQROWu5ewe63BsmcZDN1rrbysJFmBt7GF6Z11wHo/Xf0iR+yAjx18s5Oz8WVz
t4yb3OY+LIUXZLt7DNI1qs2ipgIFu7BE/UgJGX6WmAxHbBoPd0JjrcD82KhwF78dkhNGdkPPhxgr
7wxFfo5y4iIjC6unpR2LdFNS1c37Ckw/bw4P6UOcmOCofVMEaKtUtkm4rRobcOKS8MVTYYqKMS6u
5UnADtrfdWGyuDRXCciObfcfLeNyQgfhM7HXjml8GNW5+i3Cfak2gBACW+tVqJqIb6Lkq81OwhCW
ymWXtg7JYWtlUiI5549n0P9kBkuUbjl3OnKVKwjGIgMMh8IJjQYvTn4UZDCdpjov8NE6IPfdBcfw
SpCLDvUapUYa23SZkX01CCLn4JFsbc1FYPO0LXF8d1QKaPmO/yvgGvdaOXq4aY+8TAZddYmBu2Zs
6IN85b1vNMrwg/QO6hj55fUBzC6gHNxo9Krd99C9SgsRm7HYhBjEUNfvvh1Nof1GGpmUczQBaFFF
qdA6yme28PUwlNyYbnK93jYkcjZ0wfRgUEn+/3tm90XFdZoYiFckL25EarrLoB1/2ayT0eT5zqFs
DqOssJSniHm+vpDCRGzdF/EUrapnFZJsaX6qiFiXbccq6tRLfnKUSYpeu95+nQW3zzLGMC4bQunb
IBX56GwxoHHBV6GyQsbNQpWg18T/wMKzNzWCIkeu2HZ9pxfD4A/k0q9HK/dSoqOHVk/PmgPtdRQ1
A4nS87W+dEtRbfAmhPwWA3Ha0XMzBP5Pd2mSPblIzgCzfoE1XKaANS2xdkH5Ra24LxFpPiUtrJ/j
KpK8iuZYZA+1DupOhdKwGrXn/AzlMoNCkyA8XCnAuPp/iqev4VnRN481MllmjYdQ/uIkc5GQrqcn
L2QrrZT95ea2bbo4sdxH6GnFmG1wneLpZOvuJ/q1i7uio9iDMaInUN22MrKdV1yBmmrJyklHMABV
BWhruGq+MuFLbP3BzGqabJrR1rFj/CFexfVWrdgfU239rVlAD96MbjoIL5aN+GIG50+srx2ghyRV
waA/yuqPmp9i7RZvyzH7h51WHyZhKojB9JcceyK8gDiD4w9xVLBxHZg+tWiRCvo+dzrzcobX94pI
YYtb3EgSDjKFvBoDwOOGG3UIfPcXkLXVDyyhrgWgvCo08V3ylxi2GrtxR216Kq9ZhO0omZf/FL4C
O/ruT1X+Nj8RqOq8mT0SCygxS1zZ/b+XPgPxgXMnIAOUmrvr1XyG9ohbwmoEuf03g9DCZLh4w7a9
BpUFFOx4dQV8VdXcibbbVsZAplz3wieOTXsr2Kf6oa01yDoENCnyNDVA/5yslEeiQ3bDEHa6lS33
z0H5X7x5R4uVCxO7beTud1En3EF4iJSCh0BzmhPG/8dmUU9RGjw+m5/HtQ/uzLPeFtBjVNntYF44
k5tRjnaG3HO48dBk3XpkBxvlcGz4yAxZYw9dYDaRuTqrIq22zjJ5Y+w2Hv+f/UNz0JGThnzLm3kS
QlKwQpdUtv5j1AeEhoD4gOsuqxFFi9K4BlFJYbWv/hlPsQug90b15VC86YhM4tkxIROSFMwfIRst
B5zNWjZ2u4nUsEJ2nYinC2AttPP7Cw8MMy4lvG06Z7mhMSpVDXcZdC+3OXoxvUxlSf5qdOH/7tKq
152jUMxkQUB0QvcZaFSRuxzx2Mc7QMkTU/Io0YHqO7K9AeaeUlbj6TULnEOkhm50oYjplBA3IK+g
2wQhHevSMu+kTywOldd0Z1cVTJSKGcUEsHZoUb1k0PRw75AJzq+zavtk/0zkDG/xHrIgx7iMctRw
SFvbL8LvFQXozMciDL+AadVFz5OmHU6+AzViD7nBnRk2a8cpBVuCOCYSFkfOzIvFw2EfRS49rggb
jYzemlFrwpUNG8MQuTtfqX78aHi8/vYYuniyj4Uin/uPDHPbFlFjKVlu7BvFFkZe1a+OkyJa6lls
Ql/SEezXqsh39zbLzy9iwUDT9xw5e58M+jllfZVveICg/2cQZP7FiISbjDnTiOVKJWXMcGyD7AAt
/cuwMB2jlcxHiln/EnmwU/MlytCULxDMluwgQFyzqanjdecWP/nT95SWlJnmvB35nqGELcSobLOo
sCsbxwLF2EUkkQSAPnMMafXMcQtodTg49xjc89qIdjoDHLXwfRgG2FH/312/vk1T5xbCj8QrSGsi
Aa5IsYukwiL/VwjoaN3L0o+XOqCr7JroEkxUq7fw3JVygOg/470T7Eu0aBEdozVaWi49XLhOEWDH
XEGgWD81CM90/0i+3XSWxDKgAB94rzesXzvtiozGKeWdGCVRcKc9ZTXd8t9d5dkSP03vOob7xwCQ
AbtRxF4u1PbldkQElnmMwoV4NKkgy4zbwztHRgq9zGZmscu5lRjZBXHI8HBpWR8YOH7JOHU2vHis
IDbci/oR1jvIRspym9Upppy5geejQf4yzc9Je5EnJHLP4gT+xJLasMwzNdy1OKJYqTpXhO/5mw9I
ddPQEMowhcivu1FkCOAuTH2Hkqcmpa0Q8bb3F8dq7afx27tws51RIMn4UGDe2hTt2mJ6tqzzfGj9
X3xxtQG5TvlCWxRGR2veqqwYM2xcpPSHMjFcW17UgiwNCpRxJ0Z0UzSBV28+oF6/3PRLF2DZ92j1
vbcql8cUD7col4TQgo3HAobE+a8LBfnWQB3O8UQqSTADBH1kUN71LZm2HSZi7Mc3+fA6ILGKmXoS
ulOmgmPo8/1nQBsBRZS2Ul68nUKBeLpO7VzxG22Ivf8plDYn+jCJGR/OG5GHJR2NO6jigwzqorXh
0fFTdaYGfsPXn2YHRntnoohrf1tyNOSlN55D/2XIV8GePANxqwlLoTURzwv8/kphymZtQK3D8Ir+
SFO2r7FbnFGfw8orAJcT6IUcGhZ1+rRjKiJiMSeV19eFldEI0pngVi/G1y3Q6fzWBNH/Xttsz306
pQdME6CCYee/IvzcF6LVl/zkUxpz84ONAq0Ujb4Vec63zwLkHz24XSDubZubJqZoJD52qRM8Py7U
4yONd7VdxeysSzGG9zOTz0yzvVOCZMS/AkA8w6Zs95z1A1nJyLvtCKD840YXI1h3SJMx8Vu6j72b
BfWMgvgPDqKgW5YPB8mAWqgMUZ1PlA6T2ZmVuwlS7UW3JxOUhe02dWkVbZxZ46zzCInfctAKm86+
H4bNCgkcT+VTwtBjmPQN3B3dsRPyPGhZ7x9M4qzMz8eNktmtzz1RTekU/Yye0hQaVGKBxe9NkMrr
ucrqDjNM/IZ8ldFTB4HndnQVxRiA5cdeUEvy8JCeFjAlPGGax4G60MXxcTTXClBEK4vHU8oyd8kC
M1dI2hi0KYwrMivfP0YWlLvO+4/jNwfyTxV9+wBSUo2qtVasvj85n2v9vCq2qKvgP5novw3nx483
SeGmrtyOmPdE107A9p+jbyEgJICnEMbXRbKQR+YtGNg3OHMSwBGv9Rcau15oUDjzObFItzY31XXY
+a8Pb5KUSTVfHuleKK+bkjlOdTAUMV4MF8RvjaZ8rODN64nF0C4YkZBh/mS7sco0LBAIKpbzAgu3
5Hr0z9TJUyMV/H6/4JcQoODJvG0jOyiPil5W3b3e6tHV30vfD276LuTTzLFtFYblO0dIWj4gO9fr
Mio1KiyaLTgv1mD26QeIvNpTDadZzW1yTbUoEZszMrSif0G8uBEs5TB/HHOCJBf8+73pfnYCPE4w
GmUFdlqe84Ds8tFCQnVEb03FQXwseuuqbmuPxdmeynT52wfghnYH7ybpafTXOpJvOuFWKElCrJj1
L/wXOUPBPb6q4+GSsL2H1rwcCwC2/FDwhAh0UQc3b8VtzWs7R8Jq3N3zurQLoISAddwS6QDFvz54
BFlNt640aNkiJRIuZ9NCd6Z8kxp/lI8Ufgb+R5+JXORv283izOzEqmWOoFlprUV0AIY2QEaRUrDB
gn/g5R9+s0Qwcko3L7GAeFwW0blVkXidzBhQYnSZjH7vbALfBU7l+snwp3HMC6djEgBnjOvGzrXp
h7ulNWcf5Wm5OxtLmn6EYqOL1xVSofESfc0XFTk0lTrz31bJTfx0irUMee9eXhI+EcVOQNK0Mm4m
4iN/AzG1aoexn9wo51OrC+SXqQQPWopWLKRiGGXWNhL0hZwfUrkpRrRJFo5ch3g9ZTiaB28PNjCi
PhmLOzTrz0TxqFMJH1iUC4wB0gVQlnbRqHENWBzjamL7QetFg+1ltL2dXMKgNGRdbn0SWEHagCds
hAL9Qab2nVZbyklDjrjiVPlvSnXw6vwzQ5sFEZagSCDoLlIclC5UL5ifIYSKemqoXM5wDgX17X0e
KjbAMKDnn8U3HILXVudRFHBDa/DpS7nbcKkLvb4fTX6zixKr3r0w2YFmdkg38OsN6STPYOnfLBna
td2znN5/z5z9I3cNiZOenUiNVgCbMdxJ3w96reagKyOhEuypXXv3f1pWWIcY96F13MK4ebmQqgKS
0KVcxE0kNtF+1iYXeWrndcuagc4h+eQihBzzM1Gr67+P4bd6/bPA5W8AspXhccanS6bhbdSxscOg
g6ZQgD5MbO7zU84fe6CV/pHGx3iDvZnJPGNleZ9opC608Kyqi9aW9aHZ1mJ/8+4qadfssL7bIuAP
9Bv79x2q7QYbl9x2Iyj7m8xDZ/QXEpGxbX5jUTOoJgSao6+YMWmK0Zp524G8tK6yVbOHEHp616xs
x/aLQv+fIhY+PxhePFwvbwrG1gKCwL3KeW78G5IGCSn+sivhVUzGRd8AFwJeJm6YeK5y0ra7z+RN
rH2orl5gLiXrUgwK3pLOFwcJ5bbqdKfMKnd+sfeSfrhlao5QAxDmdcBXsoi/zWdABlFsPmMlE4J5
HWS9+9LITlPDSNsP8diZ7CWUZpKeY7m206gAMbyo1PSCgd2QfsHuvrZiOySELLfPDwUiS0DKIr1q
7bZ+yEAo1sEFlkRGvKSUyS7MoHIyZCN963a4jPWrlNF3xrDQegFmNtAzz8cW3VG4Yh5dduMTIbK7
1rWC/OMUHG1HBzrwLwwlW0Swk5PR7VbPdGmNOFu+bO+bb3e4doMHWGA9QOE6RGp8zfPLQSWk17Wg
9AyyGCW8n2dsrwmhevCOw1dVsEgn1uW21MCeSMLrtvfK/6ZVb1h7bZErBVqlgiKbQfTU7yhikb7g
s66vDTx/vOMBGMc7Tj7OUoWcIXAv1YVL6J9v2OYABT3Ae/DP3U+/UDs2V2/d1sE2qgN4p21iGBJd
DxnkGl1miT3r3qzfKIrjP+LeqXkslLpY6QOZa9pLYUjEApR1cYyeVgwHh5i8R5OeCJ5dSYjZxD/e
nmwgALLvffHMNzEU0rkkiNocvins78Gk/GRYrQTZBE7Zo1aXeb2sjgk7Kr3cOXqRINjCdbOdrwbO
NExhYVP1H+OOlDG5iASml86F9U2sUSZXVR3S5j+DXrzThlH9MNI0yOht3+cRxdEBKvx7iyELflvB
eqRCvQ8jjvu69qtiifYTQw15JWlHKHeESTPfPftOk0SGUoBLoCxyXEvGBk9/JU34urI0aBxNFYaH
6rKi+0ez7Ok4nBx8YSqe8hN/xhEA5RUDvlJH+w6BLlurlFMU7dcuZ5bsKqRKiA8yTRFiA7S7DNAa
qWBPJjezbkAA0g0dpzbFKQ7FdcyWFZfaJabGvhKybP7aiJCm8z2oIGqhO0PL5pVPuHMkqg74CzUq
OWIgBcB1Qz2QSnPhH8ZM93f5gG/geld2xbmItrO/ZXxomqkEGiTxjOOqdRx6BglMmQZQletubWW7
ilmifSj/tpMokFElrDSOHVnA87gxqEHBGTN15gBrwGhTNsEI7K4xViFktIChND8Y2Vo5rEZv5c37
dL7oxOsxi8NlF7qnOBv3yq4YsMmlQAPw6XSiUvZjyrMN9h+6RUO90gLQRP1Oz3KbjjOHaABBh4fS
/B7y12oQ86XPd0nhQfZv6b/RSBOVThspYQxm6RUn7Kn9kV2wWyleT3pzVnMO7YmS7UQXuv03hKsf
xyQbaPw7Jexkd8RpUeiETkpbxWbwz52+mhkwKuADD0sWV7IS95KVgrmz7LIxK/ecJ3+lZYxdXKKN
jj3nRBkf9Oz3xLcYnkOuTLv3HDx7e+1fdJz8+1ZhWbLvLtG1+GGg67lixQBrvLvZaLY0GZUjCVyO
NivnansPtq5d7G2btZQRzjesvI+/bI1v5i999JjMcOZrsn/ss32istlLEn9okNJO58nGp7ATy96Z
GsuCOGJb81uJmD4kh9bM5+Pwdn3noINzZQiMne6WL9nKgpLN6BAZp4ImtOl9LTDGoX2QZM5nlt7y
0AEP+SnW90RmHSXaGhLL5vDB6zVJ4yhhWx+LSdGzuQ95XCML0gnO2QSFV9jiIl5IgA7hgZFh1pkl
I54yHy9pfj1jJVyreFpJfZKnqfrfSQcehOBBKz59/56cOneDW3CMnH+nJttVpK8Gunause+Je8AC
YHxSfUgXTIRJgh8GHLOHFLyedxd7yn4Nlt/qq+YF9+xcxo/uFlr5SHCU9TrnGzZW0B4IPyi7Kay7
5h+bePRiS19pTpSnQ2H+zmlhQ72olLoyshBqJfYbH9DarL3zNDS+f02xliMMUvJb95xqcs8D93Vx
6zkx8l2uLvBpLa02OxxMSVUBpAjy5z5yLZbxE1+yTNMra131paRRbKfRNoQerTf/bJeIys7QbyjV
48UmBr+7exyvJmAW0J/d+lKSTagmBCLAM5k5LWPoWro5uBA4dpcwWoJiUcRXYu3ayreg68/ZvBZ6
VnLd37RdD/cFMc/kTJItgsf00j5RgKDnQ8YhxheuWqLHrvwWcpr4YsLdBbtpkXG94WDuvbYB1QXJ
eSPlaLfvxS6emuR5QuNmEZOILukJ9tq+gbPN1Bx5hzBWiyst8FgPXzwLcmUbde0zK61nRSOhrcxB
Q8U/BjRT1c0LFPqpF3QgCA513YHUK68GEi9SfmhAvXiRtBEhJBzg3b1xqFevvUbLW40BliU4mXlh
vOHcBRUBL36WAOgS+XaOIxZjWia8KjiH5fAiZ1SuPpJN5osX05OcwN+3s+tcNALfzCsNVdMjnQMt
JcjY8i5J7Ec9ojE5AoOIy/hx8Yqn47sq7iXuwhAcKKvHlJNkFYu7uxqJKTaEzntJlTewZrtT+RQY
aTpjY9iirqXTNfXDRZanggJ52VwwTEPn/FfVrUvuQJ9HWon5ChY0xbxZU/mxCUxoBQERkS6UwCMm
bX86TjmXD47DMK0PIP49yjiSkza8pTGJfKFaM3HpINvf9p+ueEIIzkuJyR1TpGJE+tVSo1AOIqpF
1CX6sNnG9AmoWpLy+Rf5ZFSQzFh2BLmR3uPyxl7gcOyCqPBLNGSBHeTce/YCUyAFOMxO+Rlg218f
LRzLkiwWkcPcr45c2JaqvE30OQvmG6d1z5aS03H5ifUPg9rlASYKuU5ZQeSr3lc9HFDNBY3EN7jO
w/YOFXMfZX6Q8pg/nidMNAShKNVbEZTwIYXekK25AfbzYmrQ3kArePHUz320K/7TitsKJwYUU/Qp
+S0WmkwGac5wdgab4EpskubSEffwGJUxpA8Q/qPyH/RHVUIfX+rGf6bYhJrwIIfxa2Lqr5ass6fP
Bg4oI8Dmkn2eXr/G618QukzCddVeLAUEqzKiI14/9918NlpePSL8G7LXnXi64n+5nJlV1lKnsmIx
yX0WK9MQRicn5zEv5BAaqjJkEx2QgF9WtLgztG6IDfjUWfha8l9j0i8ITtVnICkSQwog2AIrXESW
deMZJFXNUwcyQpWldYnC5wIHQn4f6d/nBlqg2QnCWcLWX0IHGjcQHR4NBYn5EBFKnELAn0vEx6eD
rrHvHJ3QGvts0WMeVKRSG5fBdHr+iqL+XKNe/q/PQ3nYCZ69Ej0VEG1te6QIuDCpOFZzyvQnYjsa
t9cavhjplzZb/DKXvhILYNkty5SrC/XKDitQxtSgu93AXXbvA9l/tm/EnbtK0pQZ8wy3oVGh2LTV
jPPZYI5u+OW5U79gXrHot3ACh4a3/krTCSfGllRZ2UNZhtDhRsev9WAuYV/rGXn1/TvRKvovlokF
cvOBxvNEAV5Sx2Ii6Vl6H+wVi7t7mahyB5YRxubcfHm/Ypibaa4eloLQ7r4hZBOEHnNS7jYnQBl6
Vx6liDevy70NX1meyD3EiFYPV0w0Vinqr70DBpFwNVUpd20VUJKH3mVVcWQXlpr2+acIgIeQY04D
i/WWJ9cqINai6NlIBSLmKbHnB8giP0weu7dtJRIRdwYslmJ9DhReI1Gk343pthyr6XNgQNtGguwh
BpovqsdFu8LaUzJM9PZsRbztv3koghNv9xt1KTNdht1qcG9ZtN7WAhuHGzliWB04Lu8GlDfF3GXD
DDtkv/YYpygDPV+y4dEW2qB9m9rxK77IdxugvN5k67yt6j+4bLfR27uf+ABy5wQDj3Tz6LX0u6jU
PXc0TO/bWE6//HK/J3I3du+pMvf92XAc1XeLeecPRjIGvgb9B/u/eluOBWRRrXjpr4P1xmpzYh9s
P2T43DD8C0rbgrlffYTL+6DIP9PkD/BA4ew8Y/J6qz3kJGiHvGXAscYxHo6byH+hC9hfYPpkLr4H
jeTAspNo8T/rmYK3cvpsjxUoKoEjMa2skBiNI55ewsaAUBwIWIIeAID994sRMhm2VpRVD3xmSteA
EPaOhqMkfH8k6MtslmYaT9Ul6othF8OkvjZMWkRqbm8faalB2PdjfuVeNJFDQZ/lBV31yjoHqTtQ
AJGAl0b39McsRk2CjsmGFau64CFsax/A3afX+zphFSPTSQpEtK1oKQiwUKcEgGMmlZn6eMQtcW0W
BZLhA0CPwsjFwdUYALdDnfc2EVM6oYClpOZKCiHP8xm9hcSPeFs8FhvQkLg0PEJJrb+dE1rykMk1
KQSVpvcGiInSzx1pHQj85944nbwK3FI9aTg2pRiAKgZntOaFnV3IL/qS9GUPTbwaVBfvWmvY9/vC
g6xfgbGnVsKRRpBr0tntn0yuiRiu/hKXlSiVHHeZHEpEWPMRAmkeFvnEotiIPL8XjMYtTXRot6Kv
vH4KIoCOpOTjS45eB8n00SReYeBrv4YhK1bZg8g6QCifh3Sod55qDu4fgXGC4EFQYbAqQAxzv1Nx
8U0re+WNEVJQVTFcb6yo+H9yqCxhAktsbY3XXFaSPK8niwWX3WZJx9PuR3kmn3R9Je8Uy1tLq6sk
u4/h4tz4MPjVVN1u5b0C80PEulYmHSCf5EYvpcsbErj+CVeFTcZCcS+Vb638MRlZuY8RaVYZQQN6
bI1NoZgptqfSQiDqfvbY26M3o7WVmqiRBZ9oe9jY9ev/Est6eODVJwUvbjvckZAQNJICLCgtoTIe
HDHy4aPlFBAmhMN+BiU0BOlx5pRcn8Vs1sxFmF1lUgvLwcItZs8vaHB6LHgMV8xI2n9DZCndawJk
ixQ1Tt1L35ty3jAG9LLj9okMh+2UHgZVNpj79zEPrGJaNpHbRvBbEjtG0pngTjGRp3cjdBOj8Gek
nojnMLpHNCn32r2urVg9C82z+oMThU95KkFYmqyScxSqyRWpf2qPFYKgXt1XmYA9W95aOUi7+53B
sOQ8Uj3oRVvXbF/03ysqDk2ApdUanjIq+2rfWObbbVnAgFQCbR/FcVqjB+RfpSYmD2KGVkE+6dqd
kKu24fX6hbe5qKayp3UopzHvaxgLShUo/EHL9y56oU5RU5lzED0K/g5ybGdYLIsxsI3MZYi8pz7g
3f8tsAF86d2703iQmR4+R/l9I5FCKXsrJBf2Sa8MU4LXWVuKWQPSYdIaX0VhioQj2TgE3aRvWXXT
slQYnKMsqmfppqUF4b/n+55PuqkDrTHoorOOTpv1LkJtgYvpUWwoNJEttjnrbnmwMUuP8iGYztGH
Q5Y4JO/2vkjfBskYHdoTZXt+yISqc+8WaYfBOXZXYaZxC3HoPWyTf/zgc0e9wo3dWbKsre9zZDQH
BDhgchPTAbTwb+c06Ykaank6GsrRGYHvh4I/mi5j18XKXxHC3HJUhKwWeNzsYjTG0/36D0nhjtpo
Fl+yu+C9+IlxglKBGHGESFQC8LAW06XlBvqrgAR/ZOaCKJG5cFCZ96se1Zpes9af58+2HfvxlFhq
/UEl5E8ZKqYUtvPhyqFm6m65VED88QemkExoE7u42i6R5L6BA057AOUiim8A1Xdt6E0AWb4sU0z2
vYGlYwMOwpmb236KnAMLdzLE9/roOCAvK6rd/OwoQMPcJWwbfzusFpin8TI2fyBq11hRDFUj4wsY
lhxA5F76jjHyp5pmmdoKr+ITxYl3xGqw/4rz6Cb2tX1YfO86gMcsU+L18gfZcjM2m9WHwkYrF51n
5+ah99K24YNuwhstr6NvzWwdmdjVon7zCgx+7uEc7okQDSmj0vIPDrdnaTWyLMRYgNxzMwqURYGy
LZgPXycWxdlxUFiX7o67GPDAcIANdIquCvw3l7HQNnsRQq/8rErKeIOwxrFYhIUFBSZwsIKWoNFO
5wWUm0j3z9Uv0ej026bYpzCw/ANcPE2KUlhSoQIQ/0FondwiCIb+p1IHkjc66HmQVQfhDQeqNzns
lIJo3ce4wQWAIzWw10TlgcVgnGHyV9laPwflpHwQ/Erc7Pol6GS7ZPKs73bJs/uKEpSqTvKMBfFr
h0nyKgAlIJbvzzAw5VwbCUm/My8E4x0xgAQ54pf5vX4HBhQfbIGRnxMLu450MjEYdT8kCzCQcOmk
eZGsxBk48nz5eO3fGIuSJRbzWh+60ZFzIHIbBzJIXNIlqdt0NFE8Fwj2K3WWqZZRh5jzeTeEskhO
iQKu5AaJAIYDk8YUIn4FUKGk1yy+kGtTZ46x8LcBwmh6nQlqLxrboQOV4FVoJj34C3PphtEZghcw
+zIqO6Ld84yHRZK3TEOXJTuT6QqxXbb2ZXkLLVl0wbs2/oPYnkdP/3QO+HHPgQjIHNIZ0wmGA5T2
BfLJqJm1/TNpJYzJGlwH5zdtOPp58xTr9PWD65J6sm35diiguF4ZYTykyg0tv2nYBblAWskbHaOw
dIjldNHfx+IjrcoP/sE5dL7zJKB42JL73LOSA/n/UFCcSqb1EIFwTNxDrqamgoyqQZFfFyYTFna7
Wz49dFE8woM8qbQHJebnA5uQu1OoQECzEWf/PuEen8dKPDOx8vexI7aGuJ52juHo+nsfiQuhnO9c
hn5kI4hhyLefB4qHHJEZLqGX7TGgx3wPlPeQkYSrW+6rTAvxjRbyuaLCup/O9gyFzg6YPIAmchfL
IWzEbn3XWxOR4kWVxf3Rw/DcBO3ilCAZdjsic6hXHHR4DcKYxgLb9wLweO1iExlxKSb/n/Mk5Aos
NxmJySEwto0v2SVBa+p6o6YLYJWuzqm1E/xd1nZGyea34Bx2Fk9O/PZbLKrYPHdmElzYAkXaZvqY
Nkm609dsjM5MJlfWR6AXtxsPL8WH7rG6OjuDtKruFWVFRA5kINeZCVgj5h7PJdhMJRxrk81OUDNd
njU200B+EAK42eNfUQpXCnNgMvKitPJWuXOWc9pm7nREL0WLhi+btDsowgoYwEmIUqK+e3vyh1kH
HBn+mvKMVESUEjmWqYkwQQNDQkB/tIJ+WeA0qnNfKqI7ggRxHjS3A7oIZbG8gSVHywDvrjUIj1L2
1pSC5+r84gFTeQx8U8/MI4YBgBwXTPyftSOjvpNqglIu41NplodMmLQGWNIsERcB2G77paxrZ5Rc
5bIAguaxhb/5IByK8zTB1FgrEC0XUu1SPNEOelYxa3XelSlZRhOMOoH/8Ft6Ndrz/dbAKQlDvs3B
cnF58eVnxthTC39y2wrzcuOXvwYO1hNWxblaHAsUX+kF8A9Z7r2dIgWoNMWpV8C45YCqLgPk4CFK
AXc1KsOM4iz6slWU2vb1gPRpUqy9MGGL/cBxYqDW1e3BgLefTmYhtkBwHZeQJdle0nlSKxRmoT7I
eEIM/MFh9UCYClZk/5Ehqjnsj0VoWYjStumoXCwHOvHXmu8s85n2QgsJS7syYmiLP9u5Q8p7+vTk
WEPe2tsgqZ6UURQYM80J/gcSVkyhXbNRvs5eAQjspjYaQJBo8SnopgOj3OSiuXImTzr/Coe7mVH3
fRoUpttQfF5LvGxQfChe0su8521A5H+RxVjzVtxeR1KWDCea20+Ds6NWsgWikWN0tdLXX+aFWiAe
CiY/H8lGBIgWzb2Idzy2vWeI6WuYArEuWnLMQi4DyI7DAncv+phsiTCi97fv5l0zBnqt31+v6x5P
AChot64DvamyFS2zSz2ccjcr38l73ENDNaM1wa/HXs6IsEawPEX2J6SGUzM9A2gT6khamhWfso7t
Wz7ILR0GT1/s+oyy0cDIAMBp1iRienrinTibYHtCMWfl8USx5/FvC+2G8DWlP6TNxPZnzqfnZNmk
MXtdF4Zn7b0MwqI+qCxisRWjfmYwFY5mzBcQ3vPzNITowcGwW+t5Ax2MblaiCt/RBna+sxLCj/Vg
RTmm68YF7U/hwVeGZeP3jR9t9qmtgmuhvIhiX4PPgyJWVu3BevW7mOPyM9jJChJ2vhhlolgdtsRp
mhbznrIS608PKVJJ2ZXIbwWvHeZ+ALvro9ZQCKOPj0OtIa/1UZ9PpSxi86V+Dy/Y7t8QDblpDilR
gRzRaKUf2IYxmW3igM6avv+BjwEMv4D1j+DA3ezSyHSU+DY6W2LjfienmdwtKsj13MMtKnip+2cm
YXfWJm9ediQ68PWS1YYHkmp7NCGJhQxK9RmOYeuI0KvrKBIRWsKpkNc6ChKSGSRSiobedpqtnXQ9
dRkE5cLWXZk0Jyb+PyANr5pPnu8XjHIpOtYpBaioUPdSCS1kmT5y87B+S2zR7AvydFwsVlUevWil
tg9kA02ggEebyCMWq6LQe7mORqPa3islbw1qWZckzv5mm1Nzj9gggsYJXfEA+Oe8td/rLUaJIx1h
U32/GH4yNyfiuGlswxLZGt1UMj5+WaNyL0KPoK72rosmsMAm2ZgPTX4eDj29Am7Cw93kaYEQmkbU
ymPMenoTqpWEBAM6mIOZ+lYnXchd7ZtR8vavm7P6G+7HI4s+TEhznBMpu7M8UQz4vPhbAdo5pqpo
a8cuKIknDtlDcm1c+jB6KdqAx+p0Vnc1XfGP795DBS5q7czg7GUvCNYQmdNcTSLeNBlSAvORaRRE
cni+aXRWmNaj9QKaqI88XTuhnaHIjKrzgXdlgOnppTl0EFS0tE5oNl4yWmM1/sYW6f5AWYCPONrT
19ZIqk6XylRJ+ZC13/pgrwduJO0NyCOWBmR5YbjZne9DFzm+7NMM4ymfbHhPpI3rkz+KJtz0nRjA
TnOhtmVC30mR+t3JSOm1WcBM64olbXaRrcA9NoZcHdjSnkMvf5PubRpU5HJbzK3Q0pRhUIzfUiKv
KZ9A2MIIjz4EZjLag5bUjLTTiW7o3uFGTTXEr43qXIXkJQ4HDLZxX5A1Wycnz8Cc8wXQKfPrTHKG
X2xjZX7RD4ty6NPmOHykyT/fb7MKeSdMmOZK2luoo5QYBe5RYsNNbexKiTOOkaJstfJDukCP3tmW
X53E4ALQrp70b64diEllPkfG84563ds05XYk2pQbg0ic27JUAZ/jAPrG2lt6dOSLi+jrLcXGRM3H
LDUjWqaCS7zUs8RcQ1iRBx1kyw3EdM1ThEJurFM37vqWnvzh/bYCxHr3X4QFoPYcQ9eo1/kwT1I9
oxAtvgo2Za4V+E9XB4FUXBZWxkygI6YGhlDh84coBr1rb6E07yHBKs7nTC9ssusD1/uvxZr6p4TX
K6EbANvzl67Q+QA0z/tdRAHZY2xbI4GuGNdh8nTIN5wA5+rYADd+QNe52DH4WD6Cr/sM3sD4LBLY
NoWW5CkzGO24xblpsN+ZDdM80PbNz8dDZ+4yDMnVmgBBKm+/tfGmJcbEqF4U9xv94EGJqltCwcQf
+eaH+EzV7r/YG2wxMf7jEUKVU0SBxB5+KUrzMRyminXkko2N4pgsZIuojm68qFtI1CijhZ6DHfNX
fx4nRSmC/UJ1csgE5Q0p2T0WsaEdz4fjHBusUcES09DGE5gpuL5LebwdRVh69hTLBZKv0+6BHv5n
QTrRhLn+wDrnTJKwqMabIdsqjUKKlvwYdwakv7If1IKK5fCPLyarWPQS1D7hwG8N8BOW9MRcsApx
oxT10d09KkA8LHdK3jYaQO9qMZaorHw97mGuYvPn9mZMkb5frIsr6GUI1VYEhi6EEodB/cHykiUv
joevmumDAQb8+ZqgbYsodDFf/hpa9OIwnfVuuSTnBRnY6z9/OJPy0t84fAbryVFsrksVYfBiL/ky
u39QpYX3oZc4mi+TOzjz9lzRKzLnVAafQ+2ZhTLD2PyEuskXzl/nckU1yohCZiXtBp32wuoV0XMi
fJnNr+opbD6J1Trw6X+q6pGkJkRWQV2nBwivy9ckoI+dFCp9ToDjday+hDwnMLx50ODFw/Hbg2LS
ZLRdGkAaahY3wLimAW3EfC3RqDo29i3Ge2+z1yi3/WcxAqaRx+jpE5xWDBuPGiteBdgfb1N2QRlT
3qyaviW4v0Oi4xSKA9UlQr748wIUrKAeMEany17DSNSSjcEwBzvieZhlolAdeEOvy3h9RWgZ+2df
KLGE6xuWVlK03aIoShYbRU49gCbEDfKDNtYtgP/DjFPp0ibMC4umYQzR7F1oYJSsOOd9F8hPx4Gq
YKnhXgF/Ppbs/CVj0DdA8VLCGrkBmNXBg8dWtPv4l+6YEgjJiuvv8ylgGpdd0YgUqa4wf7K9Ih15
5hQIvkLsBCWKe/W3mEgk2DW/r+5RveZwuaDABbUTCazMejeNqSLdvqfQY8qWTKR9aBGzxRKJj0qK
rF7TipZP5lKuT2RaIoxtoSqSmsm+fgDF4N3s2WvjuRdJy+E13/OQjDtb89O/P+TTXIyZxMNcHuqm
l9gUwYKulXwKn73Cpo/p7L+7HYDvrlVT385tBB/FZpv3QF9XOcPTl0RwueYYC4rOhxwPA7AoH94b
/+kM3JXsrBfUvVMagsbuv/DQMlXUnQe8f1g8eweuNAFgoDs7ZBoTdf0RIygs+br9Z/1WV8nuSCqJ
MARfeHSHarJB56rBmrx2xwObUkQTqb4pYGTVrNV3Zdba2ZEWg8hSawlMuWOj/BzReeU4YvCLgAxX
y+XD0NvaRhnosKW0TxlpZVj0/9b2l4o7fTbceb1RcxpTQZoN9oBcyUeoesfQzEVRitmG5swlJHJL
r/l4vdQw+Y2yfgqs3av+z34yQEVAXb/s4J75oel4kaAcwVEVYmYnMNe29lDTs+ahElX1smqIcF1I
d6Kd9bRjxGm5GNmdWf8HIMxF3hnvI4kuhhvIaZvv8/QWuh1R03OMBNFHw+7JXAeRIg2SrmAC2apa
VIa6tfSAI4GxqVszFktaYwC2xI5Yj4huArGAh1wLLr8Szzo+Rk9Ka5/AsVOyVQqgel+/qgYQE3jN
1YDUeyUdcRfsEac0PHwce0U1Io5qs+xhlx7E+vfbu1v/f/6tPPUAtiRKLd4KSCzmwPpAUXz8BxLi
Ykpn3hFVuXEHlOPW7nMN2AhM/ZKPJ/ahaMFYD6YXcY8uHiDPOokTeUbmOHFZ2D4D/XLN6q3atd2Q
hbNxv0S4okLwErQ8U21FolCsQ+7FJYw3XsWpe8X3ODiZKEdZa4XkXWm5R0eLLel6Cp5z17m8NMI/
W2GvFw72opv3bNcJSlgn454N526J6BEpPHLnrOLtsxWpxEFozR1oInyCzSGj7sDy3001doyRFFC8
fyYwmFM4ntTdsYOqPKLyvGIux9kTCmhX5cljIP55f6Of5Tr+x4P9zN6TQ3j6Z5mMNdf5s6snu0J3
m38n/6CGAQ+oDoM9yvwyu31+nW9U/GSi4t2Ur6tE2tbPpOODD2pwxFOyEWu83vzVLMSYo0q4Nv1m
W0d0VrhivpXs9TJNAgAaqO9oVlf767VikCRl2XEJlY3uoWBYLcxdFxtvOzm4dsRUzy1/m+bAubz/
YMl1J+AbebV8VsKxGsS3Je1p+Gz0XXIoSIR9X8CjCt0imxwIdgusvZws6tN3s0XaRLdiW9WYwcD6
WRYpRgkizYBmpMd86hXjD8giNSFwRQoh9n66+dG/G1k/2mg084qXDAudXvZkhVoBTaVCpl6Km4Zi
cYOGLn3TTE5EQL7UuhMFKCxhQDLkvX5lRJVsjNV/G93nku81OXLXON5+1pZBxOYC/4kPz1aUZ3DJ
jsjcwP46/4jWw8UZBkPw1BLCF9Il/tPQMGWhRU6rZMMPSTdamwP8wbHtGPIjUAyBoVAGZBtuvPz9
TD+nZYstwGz+hT2N7U8n/gLrcv5Oxcksrs7RB6WPtvIZ/gwwVtgxoZovsBLPr0WaY4jTYLE6TSD4
b7rPgizQaJ+jDzT8LjUMcdb6OtW4uRVYHu2fCPlEefFwsgvz78ypk50dsMqRiyC4cyWRdf7l0Z9f
Kz9E2e6v2GZFN8xJ/O5EZla3UlH1ARv0yf23w6KfCgKg7O2RNQVsRkylcnRpmbdJ82If7oyEIrkC
SNblKDMQhva1mPCqD8eDN0b0idu4Mj4Rds2sKQsUH4UQZvMdrp9n3J3LaFN74fxpfsCugjdBaFUB
z3REJU1Ar0zgtzaHt23h7oQbbgchKdsvLXiXG1Lub3GknrEoaY0pWSw0OyEniLY8IClJWRQUhM7I
ub9r9TEPfSC8tn38Ah45p1NbAD2T5eMf2GiIJvxHHZnntHyqN+YGQEMF7V0Sd4mc/DRPod+yywze
+nnLFmDOr7gTtnj7ialPdyFNecj8cuEM2dzwjBTx1WToDXmKOCwP1vng+gwjrZK5GuuPX2y1ZFlH
HXaTeZCymAaIExPh5EjogpUsqL2eB2SCbOy/vogXcc3bv1NPjq+2dJWWXbguRO3WpR7kIcIl0nsc
n/H1u/FRTgYKfjpYc4W6Yk87T+BP/fTiSs7KJzCio/wpE+mF9xrqZTXC0HfZnKtQ11jlw85ERpzv
6v7gyT7lXRPgf/hAuNdBtR7THIzISpcilz7fbYjDP10B21gD9wkQgRJhepxbTf3KBr+oT5qHxWNl
zx5XxDyeLAbHD9NdmiSPIGpjWq+BbPSE3pRLzfh0YpZ9qOvDbZIpuKuERShEZL+LVR8RjYBNlOfk
trV99qqA1Iqpke+qHsbQhRSlxg1+07cSpVhCBd3qzQTTXglaNTUCBg70MMd8JPZQBVSWvL1xy8k9
sA5YtTZtMM9ayMADyXwkuTJLOnbsVESfnNIih5M+dhnJzg+2CXFmnYFsCz8Nkj2KF9DxJCFM2NuD
CBESs7XfSfsp5LpBkvbvKROPdpgP9FABmzmhNvxaQqPqxNy0/PxMZfjY4AI/hWF7lkd6+YIN1gjX
U56+xaOh2EUHvaGEwn79Lw8OczdLv3Y3QEgSCZXCmszu+ra7bQSuD+GS/uM3R/zpWKuGnFtXJYTj
n4yTJAxBJzivyJBEEt18S/v4RaD1/ozIyTp3+EQCDmdBllhq9HIqplDd6wkoK45Awi9O/VQuv9Ny
h0vB+jsxzF0bBhG/2rtsB0t/gU6RjbBg3fdB99LrHVJvSkA9xKUha2Lng3/NTmtFnN6WW+CWbseN
Xo0WRuZu66c7xhVSqg2xRYVZX4sjU8Q1YoTpExv/aqhzMCxs4/k/9a8TjVnyqajesDAFSKow4cEz
W8j3cjHafWOmQYAPnM/ZE6k++dI5dz9rJ5Mz/j+tMxsj8fQRcv3G0fJjyHJY1cusbPhKxcQWEPdL
NQ+IVvGzQXlLMtywZFkz4RuElPnFXC3GSkTVwWqWiLyWrXSB3yhBeU7N7cjEjVChwn5wki4pibRV
Y8wr687wxVJDfgGzSBezB9tZmMumFLZRQ/rMDU0CrGHVBjE20GdTBewZnjMJHCy2VTiD3R5SSAPD
7sfDUxWah9NstgUo7Qa7xvculI+MfZhVijG6cqptkJikE3jZv2rnocmxWHSDXXNrf6FqAQjwcuUo
nb4Fmi/RJMkA6443SJQuoz7IgmulAPfzTmvo/ceWMR3OV271ffUIACcwiYb3QhGpI/s4Y4dvPTu7
e4jWwX+Fvc2zpkmscC5e5TgClrfpyN2JfXIa9fWlIQ/3hB0qYb28/+R3hKqxaMRpy+V8uh9y3rjn
4IiGNJMFVFqE579wdcpm/gqUVuvJQ1LPHymS5F6yhIy7bOPUqSFz257LbMZGSrr3SEIcs7N4f+Je
v+rOjuoBXYpErxhKF3zIeh36oazTj7OptT1HpAUgH2Ft8XYoqGMdIBMiJ9sgS+bC9UbN1nfxdDWZ
IY/BTeJaXEtmPZAW4eK5rg3j9WHO52KWH0EB6AYlg7+D1zUg4hlHL5C7icixYoEBgcd5c2n+yDXS
Cec0xXAE39rjxkIjrfbj+w0cOL8Snr4N8J6Bh02J5QMT7zt044TnvPene5bhxRFxkzw2TckZLXSf
TpGqgMrZVYlYzjevSTxsyJSxQayBOP9L5bIBsRcYnsEGDBTR+0d7bDBuAqoNTNUwLnoulUmSyiib
1nye+23VdCO4Cmuejl/EIunJqrGdpvOeAQHIfxx3D2cdUcW05Is41EMXDz2LTchPAHgFyj47PKv6
09vajEWIU2YL+TB/3a+77mDO1IaEb5qCIz2JMXUJdkNeLeueeIxvnqpIlsc263CUjAvInxhF+v7q
6ZKZupBE6srpuMcFOHbQ/Q9ZePat2j5peBlxzkNeldlRW0ErxBZC7kpQkyGhzNRLaGbboQil6taZ
HWPfjTkr/dFwOpP9KtBJ6Z1zaeVHavFLql4FtOKnY5Aa4vny2RsykD2yWHwlBsb9r1It32gjIYUL
kYggBw1c45uMRB7C/hj994A25ND5z6ZpGnN2HAy7ATGBXiVgFRkg27sJfW33Hsy4eRnHtwb8xCgX
nx6psYkBZ19wMbg6Y3iWWlmhxb+gm5tBDPqn90u1Eu4CQ7/TJTWqwdsYC17RYBfzrlDvQ5zCobqT
57ZvTNn4Cjj6UVVXDGleKQutk6Lk/xzMW+hiquQjdr1yrswalj8dCWSIfECYPxVnRRDSjl6ltC8I
jXuYEjh9pPvjyxOx7CjaUiK7cJDvWKdQ708mdwB8+JV9XOzxPj3wamAfClnuriqkzW48q9L7TFG5
bD+D22+zFKHAk8aktZpVXzrJsKu6pSoHrcpdbnjD/SdyUN10G5rGEx4+bklbDsuyvG64O5YOfU8a
rFf2RUB2iXm2T0w2fbWXfc8RNgfwzifGlww+BbsEzj5IQ8F81FU2av7JcSxWEWl+jo9TDEM5ORlK
9E6RlfD+4J18zVGSDT8Vx+1SAlveZ7sN/L3eYzLyoEkWYxn033O/tG61tSbnZ3MSIJEXsn51aPhC
H9oCEieU0lT6aPCQ7rL06RmCkZjAaP1Q2BkFu8ww4wbUC8J6sGDyVeYLFEynu1DEI6ZF+4svLhTC
670ieCte3VPWzydn0lMRowzYsPh12hWGBDeR0qB947RYTuJnBqorBK/GQSh1pcLW+b/cJNQPp+h+
alFiNyVq9YGeUwN0AAGDGbaMBvDbYo6jPWWznATMrJCzZeeY4F/sEiI9n1GR+fLTmlz4c2xa6Ffg
eXp6eeyzTy+JBmAAbF1XVuJ295I9KloKJYPKFk8AXiSOEKZeWHqK9pfe84dW693oRGmpOb5mdWlb
9RN1ZQ3ad2XRnKBkanW3wpVdRmAAxFgHTuequ5JKK4eGd4MCHmB4U3SEez2NdsrPlsukbP+i98qn
WYXpznb/AJ+tGo5vrIxNCKD80rmzg6+c3CdnPJf9XZIvYDpFVAWn0DrdStoxKdRjxen+eRMmx2ia
ZglsGIjnJdj6JmJrVATp053z/j82VVspcr812Xaofs++zVVO5k9dKWsTVBdaRxbo0CpbfbPEQoge
1of8sRsPK8PvmTitMiPICn25v0MitnZy9sitMlKdc1n9g56KZD9t9pa/IVfPs7Q+iFVwvUBT5CSJ
5D0in3BUw80/lUk350/Ay2647scsQlGv5dgasdajIoPcRoEIWRZcpIkR5Krtw+o/VG4TtLFkYbMw
3S2g/1jRH17ruzRDa0Knn20llunoN3lcWK7OlL0UD2CMeXReI5ZzEtOmFq6RyRLY5VRwXEISvD/l
ZFqq0jxASLw6676jXQ6jM2OAUNwhQZZOUefMYTkUC5i0f3VyG/o3Mn64NQCXLgmXR7hv7YD/6Lgv
YOGo6855JF8sr2FnHMWJ2Y/zeoVmYXBe5DJjhrC6FoIqdt22PmT7zNtEsngukHBZYSuFaS7jNM91
ZFG/YKYzgLAJDonwROK1jLZhZVYtBaDSIW3MEWSDaNifFqWF962F8peCPtSwzjf+lX2s8L2eRi4l
IW4yt98xdBgNkKY162ghDRGAEXlhEOXuTYciCvONfraEiCl83EniPzpSamyhGRoerPm0aL7kThxD
61UcoBCvhb2gsFak9wraFJqfiDpfGHuD1sdBGvaNShtI6j0tjhQfhLAv834YXim1eD5QiCZxBlU9
OJFzVra6hHkfYcplB7My/egjx2OGJ5KIIfr1edNQ7HDYFIhphqJu+419dVmoBXfKPXCOhblre7/H
JTixAutxUWxjaFfMTNIL8Q8+fElM9NB+GHbLR8QXwon4I/WBX3midPowZ+QfEE7Nln5WQFe0QSK8
QLNbqd20tLMA4rwU7ZBTmm5olFiimz0cKp+XoR6bTd3LaXgocoT0oxvUYrwguinOdbjC8SD55yTm
PDaNR+0Eqz/KTw/kagB1juVS64ua9vEsFwIi0H6FyRrPC86UJCBGbAJNHIJFqcojLOcREa5DcfEc
Old19pkrCA4BJWXiUe2dypM9V1dLF11EyYJw2FVOj8rO6bAGwSZKq/Fqn72rBsHaZGGWSiADf3Jq
i0FnOE0tttCEh7O7dxWYafHEfiPzazR+20rBm3hi+AsTBMcm/rLt5N6QUt9LwvgO90uKQEPxJMaB
dQAuVsTiajyPL4/AezMtHdWF9asCXfbQn9jO7tWAjGT6xWO7ZgPo90VjkMizr/R69RpXTy7NvZGA
CxGC6c3U4V3zU9HqHKGVhGP20sQOxQslI0w97+genAkv3lYbHTTJTWGNFd1FhIzNOJhuLGoZfFah
MoWok4TYbjrDuVS9JDs/PW3SFcMAzCDxSebciqn5huo0yJDEtZYX8KzTVht6w8984yD98p68F5b2
4Tb5bvYqXyx7Ta1iZ6fHrBl093rrqfIOe5nD3Xq9ItYp8zclmUz7gXhaqZ80t2o/+kTzGltA6s/T
F7oVlcTPS6AKyW2yZaN6mAtKgKNyXabnjltRSNlVvJvR0x+9zPKxJ3oIT66Vh16tbOt8HYa2RMQ3
5A6lKs0O5OdwAfB6X+rGgXhFNM3wRBy+IEuDOUm0eCtzzFWrrc/fmY5a9g0Cip7BsG2azYCDYaXQ
0RVlgJbOVwpiGf+vC1X6q/4TdxXwBaiAhDKYXMr1McYtX4cdJiUagWvrbwajGOT/mKVoiSm2SkIY
gdWycfyzUdgDb+WWTiCAfsHNpbnpKGxFzCVxNgbDapopCRYUZKQyWBojUXq/pbeWOkWVDhrVA4b8
eQ7bJTwEqEVs1MYanX5L8mpy6RavxGOt4/NtT2pxX0lPIr+3ZyaV90QXRsc8g8EutmOWJNP+83Oi
vfP0vFN/CSJlGETqE5Wdi9aIM4nsH9VGd/GtfYyiV8qtNbfQI99eP1SPbWs3XmwGNkfx2reNHBys
We9MAwIEG4hIeKGya10LyvKVxJa4gvTp6jzPWjS4dLGjsEwDk6Re11FTFEqVX9jSN0wQ5wX0/rVb
q9kwzQ1J3lXHx0p0GRe9OzubB/9d3uCXU2kPvL+bBEAzAjVoQJNj8eUN9g3TbKSuZ4osjyZfl1Fz
TbEKkWtvrtGzW0LufM21ExVwU2MWzaoxb6wnCTOuPBKxYl78LGpJbwP9MMbfoKMiW3Jdw3VYccmB
NTHLy9VBlWmFu6po6a6Keit2UkHpdjgZNzt54lxBw3bH6OPUXJ/cD6m5CBAfCqYq/xwW2EoM5L6i
zz32MZezkPUVhBh2Ve5CwqxLQ2e7XLU2CkcSqWoGx2o7uotqKo8BlYm5mykYygFQ4XqlhPDsDyvv
1yfxILpz+Fx7Bctc/XQdpU5LzkJRM+twFJKEfgMHT5+XEDpJu/XW8Y6W4Ntnrnz8Ak88ikyDavSW
izHs/g1/935f4XZbUlzW6c3KAO1AfXr5jaX+kNFYjFEBOUFIzBAGWUSxCVTYwZ+yBgqI4kmj0XhM
JuiLZh2Jyh4oAvHEEb90jmy4vF0WGfLDaSMSGXZpnIBV50iM4Ax1cFHqCd45De9iqIf5YyHh8q47
TzY5/kA/0axf6+84PxQFs7t5DA58UrhKTO/PdrJEnUisIumeuBlkAi16leRl0P459hehcfXOj+pp
i9QsiLbGsIeGonGrJjfl+ggZ+k+skNdnyYe6EEXOJVDz9hTVM87mdSbDYn/ozFgMzKokSEnZ56zD
Z1BHsoVQGSbD74QD3ZGHSJTub0G48l5uT85IKW6ab2+mCu+uUYgtGMB5nypf8B6hFFlCsk8yEpi/
sjktte291OfreWMmCXgJJBy3TfdF2/xB5poq1hYHVQ4M9EOOtyWzQaUhmrO31o8pOJUIrM3TT4oN
POrlYgsBcH6bmCx27ep12ZIkDo4JpEqrR/Syb2mykAl5D3i9Cwv5m+84qwCADHA9mP1OmvA4a60w
nAIOL4arNEBsXv+cOGDZd2veDOEc6tTbtm79mzhRp/Ds9tNU0dfTuH6jOkRJsVHmEDZcZF280c1T
uQR2Uxrdnbi8dV45G74IslIV3HF6gyyoN/oEL1+2WMI7W0lAP4CWL5LGcaWYpJPb1QsZCO8fYdEI
CgwY8+hVr4yma3ejPSWVXEbSS0UT2gFqoQnP0bnKpM0pbNcWdW7ORmm7fWYPW0ehhZxO/dADkflr
82hB5ud+nsyc2Wr+WgxjJ75zAFBg6trbRzP+3PREnViPnHZGar6pfBnAmdk95ZzChyK4pqViePkq
zh2RnLQmOZ+Q8kWigssvdBdQrcqOrhMyQ9lEzWV1mf1t0QLNUTYNQG+occHJoraZCk7zfXxmZgTo
OObZBJAQLz9kmk4Iuulb7je5vNjkF672ZZIhwmPZ3I9tFPMT2G0atY5bMnozS4vrGNVUTeCdM4i5
tjwC/SAoyJDaxPcBEM2uPhU7XQ+yiJQovd5rLIdIbAjMyrpyXejACKO3qarBFFJbuw5GV3bMIko6
j2k26mBL6Pp9d4HRei3XzF+w2iuEQ1/8EheGc/eCsnqOp7dNvK6NfVNs8MPCi5i+qWe5upSGQdxI
9Mhr6c+Seq5Nk2c9/U90BiaXKPK7hom84ONO/2IoBYl2UrIePHmiSmnS4uOAQpLLg3TvoE+Ht4eX
uDF3NkD6QQC56MUCbmMCNYx18dRrdCmVlL1zsLOnw5f/fAmNaSjRYGvfIARzuT16T5xjf4iFmD+H
cyFBPKa2rCtHlsj+r4NmiexWmFPsXUDKgYGmR8OvRqksgd8TnTD+DPiU+Q0ggBkbw5GR8XvkjxEW
56Izaa2mB6JDkeYMaDIWoftUCGVueLRAaIPVlknbDFvt+KInP2I8J7gORjdiW0EO3t3EX/7Syb0k
8iJLnV14zMYcEnik4cfNM2P75hcYNr5n6AhDnNdWhymmfBovjUQfuUgMrKpfRKszaM+ooSbvDx/i
N0rEY1aTA2H63EGlCkBZVuALRQjgte+3r1QQuhsjQGUbANQDeihknFqq/2OK/IM7wY2kVRL8QNP7
yJkrZ2PBoVHpD1J+f0A0W4jQKa5wVFwsMkw909m5w+LJxcMOjyiAZ58p5oXeLg7VeV0nmwlAgb5w
8aD2fi+VXa7h3BC8naz5CTfyghOPqt9/KMDv8f89w/NY4nZ/Iw46E3nacIyFLV7FeoU5p1dGPbTS
0KZzs4LjSo9pDnD/ujzL1bLbhsmAe2pwst/Ipzjsd0bBx7LJBr7sLKoOKHRQWCHhqxj7cDc2rNsG
6xSCTCurW16XgD7lZY+Kl0g/y+VDdeSLrM2I4iI8igCrmNsBt1a++PVr1A31z3GbsNj1f3I193Mv
JBtGClMzM7hqdTzPupKjlUx6qOrdV07NjNjMMaZGsNz+dfRw4lKT9aKwXcXFwGZ+jowlVb+X8UfY
iBUnp/aDsBK0tzB7LtQWfyrmE0BWE7CklRgvsvDnjHFm9WqXMnt0zBpoR55qLvhof81YKiusjzfj
CqX1tw4EZGO51AtDcRAny/LMgJTCgaptgPXit4SsKm+uvnJjLCaxD1bP9sF0VXaVG4iahaWtLMN+
n+BJnLbs/H+ozyQYx7MKavoWb30SFZ1swZXhS1npAnhZ9OO1vyvIXq4lL2d3HwoCIvNkOTlmI70d
I1S6Xa8Ot0IGwruqajeqwV1yub7X+Q6+ZhMoQTw3Czt00ciURWUCGBXxHRHXc9LByCiPIge6tRqd
PKL6IvCU0cVXILKnZmmdbwHdFCp95A3poABhazJAha7Q0HVdT/0PqFOMZISneRytXH4pIgIpAfaU
xIXfgWhGYMgyfdITkw9UGt3be1kcQsDzHC2iBUyxrx+xlP3wVs4IrQAdjfKuyeRvbsuWUKnYhqVH
Omrf3+bJPGUisvlrCDZO1ElzJRinVElkmpkKZr0AGX8+phGSy4oRH5Apt3DUa5X2KM2sf3k0QLhd
KAUq6zfmcD+ln+7xohcKFCHPee4hMXxKWgLvi6B34qXgxwFb/M02BXcldfEDYmFzJYUujwlpqPED
sS58Mxb1emymqpWoXYwQ5SRIA9i5wCt/TzOkGe9vz2+cJc7hCSnTvR7/7KR46G8Jt0/qIxdwEp29
buu8pFIDBVtaEmXb0CqCsnLNveSZ9r65m2jQfO6DnCew8O/Z8F2yrLqaM8NIK4Eoou50sqCOKfpp
r9ei4Y4MxUm5V9c0iIYsLUbo6ubEzpE/6Hqmju+FprTf/HK+NZjHTC2pRg7BgUiiMWbczkzCE/ID
y94Ts1TF6jQzJKfemT/444gD18DkrPEkWLvZu372PQPfTt8tlh917KS9Bb45pPjzNjeoV9z/7e5q
+ffN0AnFWn1u+a0oLdnFZ6lESha0ADreLZufpWWFlee2P6PgzC7Vp6s2HdVfIgU7ycrYXTgmkpBc
LC8emyUJn5nquPQbuUr6GeeJkaDV9P3W0ExOkgHTAkExCwoYoy7o5L6nQRU1i54srEkNLTQ68rlY
c841bLyyNYDW/KgFgRGD1dTxGeFUjMsiFLhMRYIAuSTGE3FjnyMpKMDOj8SQza8xwmgLtNXh9HGj
bsTeLZC367Doe/HAF0bhyMJp30lGNvv1y1V8XFWyp8X93sVD6NIkt7DJfv9zdTz4ZZtHn3Fq1FC6
YTKjab+UpvrJv2mzRWZSA02rsX1Sxp8zUJbo2Q6Cw1UofUKEg6O7Q4LtfKGjYlGl5naCQWL0w/oL
7xI1YyBxh+jkDzhNweAQn7zpwZB7o+I6jrxfoGXz8Lj30XNDMZEZEa3WAepFiFAsE1upMt2YqBwr
2H1M0U+SqT6QuupzrwYgyh0vv4KoPFHdCHDkZje+8rGQIsz5M4GZ9wMCjKPr3h2I4YEOwGP53hGv
PEmwHVHum1vV2c5jWXIIojX8zRptb7TqnSPpP9LGdWtMm9BtDTLQZRpUMOtDv/2iBuAfQCDD/7rH
OjfLwNZhwSNekpECQ6WCl7NQf1QufqaDVwkfDVyDQsFq3gH2GIWAz+e/ssQAp2FywwBkKOGDjhOd
+IfFi3cASHYIXRH/KXpoLId5eZHWIGd38XzAy24HBVsgFtcavrfxDdILq9ajTkLUsqhu6bNOgTUl
UGXPqx2qFEyv4uabMFnie4WFWXwgvViXOa8AwZtoyqMlNwgbxPzGJW8pL/tjxE2jLPIfwnznnaiQ
C54XA84LPE2u/VNxVXw6IhWmNRH5TO+TsMBBbmDl5CCdzAr8WKRE3ZeCr6jk5rrozVA7KkXNB/n6
9IgZOYA89TL6H56qmKQK1ZeGcrzLw+Gf/03FhHezefvT7KIK6+USA9ybNntvBW6C8bg4y/rKPEEL
QtyoyxaRrPwNjjzTtA6JLVdpqcjtyIj7KznbaeXIJnYqLLG5rgDGCyEO994XA0bAel6fO9VyB7C1
n5NCPp6uCiRD8PN9E+p9gkYb/wcNF/s6GO/md5bDG1liNrwXC7lQ5IQt2sEavqb88ZBU8Ws3emes
ryNIl0cGchSZashuBiX6YKwT4/KsIfvsOddfgRPXRpiQ5fKpk017otYNy5T9cnFg8fsvJQvgUT64
awi/wZZ316G2lzX/1MKclWJm+YKotfFa5H+zSbm0BgGG3EI8osCW6uqxGb4avn713Xdfo46xjXtX
cTJkukkaqBs4avyWVtaJsS3KyYA8fJDXbn4HHV/01QzVZv7miN4l28j3oNLPrAgHZ1pYn8EaJoD5
+urNAuBf17d5jFr4kQSsFPhR4/PhJAPIZe73ENLaCKN0SQ0mmR3xCvrRQRGms4Qt3JKX7d7ahjOG
MBgxHftod4RGyQvGePBtxfoTkPnBaM7tSLdmOIkJKVsb76vVZq5mkk7a2eTGnX91BMr6YiIqh/ct
N65coeC55RPfWAXu4Jnqd1WgpvwvjvUYztCY9qliy3NJmjKBbYZsNy0VqxX+1gpYrVOT1ADYyzVj
MQAF2yS5aJgvZsns7KdDb5BsVbJ8D4h9GgeeFNMUQW/79iQ5g7s/etx3XQFppL+iVYM0cJyeUN+P
fTJFKWmFvXrSpVykVV5FG9SFS4k4RfHGvhvFHXaQMEDPJbuFebbwLiy82Swm9PAhbjqeT/K44bqE
S/TzNUWGztaw9JQ7tyLLbhCnSPtdnQ5RPhMsFgXUtOgV7ozvhjyzhk5gugXHaFxoHl/EizjuEXdn
VR+2bBGcZMBpei2ljgTxdDsuRZ8kAmzIAotJ58/+AuetErIh9zFpK846qEIANVwN5UprVQqpQFkC
64vvtzcufCOzBohXCEEcbX+7y5C4YDwdrWb8Zaiy6tm9Hr93AXnkK5ss50UBJ2959ZfYdZj97rcQ
wLEE4CWk5oef41nQNTcXFaE1dA2wnv7+/851iUTCDbJMlJkb5pgjh5tunnTq0ehSpZSuo9Ph5TEn
VM6e7NUxUc9oKj8LPmJvLH7ClK7w0lIpN4yPltzOZ+aQZf2NrOaaAG24TYhB3m5RIdLoadWg9s90
Ni4DaVaguDbT0FFY89NwfkVcD67Ov1g9Gv8f5XsWprywEZ16l8r/+YGxUpe2WivFm3ZfalWk0SnD
dqJCDfnqkC4gOoq1zFW7zm1ySFi1t2PvJhVZ1L0HDqNw8BEG07XOJBUHDfxI6GTpdiRf5jfqhGyH
Qt1YfzP6KsIIE2X7FmrXNVu2eKbrYKAYFXKqmSBjGykHdlaXGBwhHjCTSghZuh3Zlr3tHQTQ17Mr
jtGYaF9nnrV4W8p+6pyfA9du3vdLSE1fYgW8rDg1HuWJWuM1o8MqN2P7IDz5qibkYTEP4jGBxaMb
uaYn4nM1gzVjNKT93CKACL3wsCwdDoxEZKFxeoRLGlNW5EDoPBcqeEDoVM4rRGBLLGU4pgJi+2jD
JmmPIojyDRY/gHZIBjxMM0Ojh61u5AeDNJYngtyq5zSgE388jj2CDuvjVIJ6qe+AX7pLXPqFLrlI
qZkJKxSFVZ0OeIixB/0Vn1DDnmRRQb5alEX/Ah7CfMCLQJHE/7b6rJgTN6pQR8TivfApoLRqUK30
x/RTcEN0pZPW+tVX8XGRBH+qwsw2Cqp2ZIyxlEF/bnfF/y+gaHokhtWRfTVYl4bHsDCp9n6oWzny
VqMGldA/D2KLvtWApY6loAlQoMdS/jJQULGjcSHjQFd49Q525QQem0nrWWmAGI12znb/KS5WfNkk
5hGMQb8VFGWE0Yx2h3ZSYxTEl4/BbJLn5r1ykfjnbeylAW9uSuD8XIqCD/RcCY6cmk8wojeG9n3z
apQrd4H06XuR+EpEdD8on0suf6O6uoq0vibdxBXsPUA4fXVHpiKCY/IWtgSiOKsYqVY8YS4p+O9B
VGCYvgXyWNHbmWMgtxjSf9mnbH3uAGE7PanW9fvqdhlfWd9TtmZWvCRRFtx508jiSjsz2cG40EAM
QO6XzffG0C65GVDPp0JnM8gLby1aCuOvjUo8O1IETBhoUUTyzjZuzECE/8q0OA82/VrWHQ0caFL5
6bf/4XpYwHe1iZxZwgTthN+B5EeRNMMHjtdMHKk8ksoj5/sPJFPQeCstMmNYH1npd4qahKoM4Et7
29vIS26Yh/C5Zkogcxk6GsjEdL8rXLlEtM+h5aMCpxf0lqGXJAt5wQ1rGZb+vQaHYldclF7nDIfh
0aNBYEth4s/vuWpXK5YdnosNZSefz3f0+emcZNA7vnR1o1P0Nfyj6sm0tsmxeP63nDoeraW5Di7N
Wo6kjZpPfrxWOcUMvz74mCQcy8TmVSZPbOshmft7ltEKDS5SbCNas94nuYkScJXMJ0QovDLvs+gg
ZqKtxuNAzl5WMhdlOMMlvFTCNPK5IS0UQARWs1KPEihJrs5wgbLnWs59///PxS55HRIlkEq+XW1y
/RwjzzS36YrngsLBTvFUl/AWq0LRpSuyOOn9xPa2VTki1Y1GcugtJ4AbuXaVGBJZACZ3kTaghnyv
rwe6iQrUTX4EYsKoL8o/I4nBZyq1pBZ56VzGeME9/kUeIR9z3+TXkf6wQ1s6/qkuH4jy3jtdwW3h
0HMgHmGqTUfyIVuarxA8i3McMcQUSvpv+BrjhS8/2Q//Sv1kJUkpoa734Uq5ChM/NQr18r67XRGr
CkdIPhNeszx9x+16DJuMkmDToo2noE67EhMjGGEUXI7IvtHsnr0Nc2zU0MNlluWVSRps+sjrKr/v
MTqFro6j6IcLOEd19EVir+oyTEaOTAZAHW/LkT4Cxm/fRyQgjPWfQoNpEvR+rH4E3c9Z139sLLp0
awtUme2BHwvzht06TMhOK9XKS9FkGXJYNQ9SDHdkThIi7yFhO4wMJzR0w9VV+rIY9u4Z6gS3R1h7
tFJRyGC8z8WGctVoavvRS+U8tJBes6E/ot9F+m3n05THM4s0POSmEkd0XBzV8r11zJPU53Wt8r4D
7wXy8zpfPGs7XS8Pi1+/7Lts8TZbGsnCpqJgzdZHPXSIAGI2tDrvdtzh2+ddHQNW8ZGiDGO9OPM8
A1RTU8OdxPZwLCCnZnPb9iXwllcVUBfg1O/Z2ezWyndj+V69cMycpG7PF652NGc97fC2H3UyY4pF
As1guITEnh90iHMGrRWi1K1ccpCET3CW2dhypiCR8srN/Yln9iM9vJIhury4cJy5fZCQ/7T/OPhX
wMW4UC7DJQA0ZFgbRF3jtVCFTW6bp7yk4z5eUcVgWgvjpsxSkEFigTJLf+TVvSEJl0d2Ox1UVsTD
7soopgDMWkQyPeVRCc2ajBACw5ClnrMLCruqOBGyOY/U9P0v4wp3wzvVrR51bUCPgdzeAP2nV7D6
OrQ5FjrcAPvIFwOQFvrdvwEyOnx+L+n6X7ytWgpVVvyYsr+gzUVoqRcAhKROhoTslwC03q3T00vP
9J39P8lyvX6buB8SKespjVpqvrHiSS34D0x8piVfsAiNBeNPnaM2dbGdNkwbicwpOERxZIlcNbxw
mJwWzr3MYWpU8QW4wDc6aX7sP/WFCzw7G0tjBNK1+8GBE7Z2EAfXWRIDPTWDyR5S7Pu6ge4Kji3+
xnovRctNAOQe95Y+hVQaFVQXDeMC5tNdwuljhdfnsIPr0NtmOErmRgs1L+LTM/uDLdmt7dPORoPJ
am5Lug/xzlpTFXz0ArBan2BMC+74SogY0XzBtdEkdU1JuKq/AkQOI4r/Aj5BkQyVQgBZHib2Lgax
hV212eETdfkeR0Dxjs6Q9Z+JwDMkQ3VPmPJ2KCL2w0mrjnz8hCQOIbB85eMJJYxWUjI5E8HVeh/9
IQlFVhDRnuw8IClm+PG70eJcx4RrvfZZ4BhPVeqjHmzoH7e5AyR9Szu8uvaOpDIk9uLtXBAIyuUY
Nr6Ad14aRenNwv2yew0COkKGAdAVDNOjftTcLe/fnfrD6Rn3DBt/k7PJcRvmw6hRI613Pw5bIKzW
KJb68mnOsEDX94gPJU/amZF2ISFI+1/AvdruId9C+m28OrW1zbtGWV0IYCTSdw/tFuHiEpOwYn9m
O8QYoX+NwwL0VWb93FVJUaO2+NsNv+ybH1MT/690shRLXU4U0UrSiD9DgyvNbrnQpmrSQeBSO3Eb
Q7wXGCHJIFGXL8TUpFNxZnv/yY6q8X4r6/f9tCf2jMQ+A++XJgk0wxhefBAwXk4ORF9F2T89NvXM
Wf7N0u6HhemEJNtOzxyoHu1WnWVmmH1QCAIWqep8kLMneBT4UO/3gf6+AfakZ2XtetfENRN18SvX
8f8/xCdcO/04BoAT+Nf3Zbq0WOTunKWLIVM8vsq8d6nhKhjZghOLvlIj0sMDUxD22KGFB8dFUgwm
EcsIno6LKzMwmM+avIVg/jsr8Y2xeR/oFSTrFSzWdtm6hKEbK16c+Ck3KX3H0yRp/v3s4h5xETlO
doVh31Cd5xC7faDxmScQgPdYUAKQMuz5yKZAdtF8T8n2BRFVhmXgaWMugr1wcfwcRGEYLirlHcXY
ftjg0elCUPO92cW844qfq3nAA6iUSTSeWJZX0PN2IMu9MjMHc+PY4IsBCfY/EMCeYDvRFZl2YBe5
nhV3/MtzRw+K5Ic3lZPcCSDxcwtXRUtmEf7v/jJe/Mo85Navne0XQitx9yEnIWyBOcBUw0K2Oz9p
FFEYxRYkOF9V463bv+qK8bW5fdNGVYGhbWo8rQb/U0IFDS6KnTPt3ppIe1YTQgxAikpJ5iSH1O2m
VVonR83pIcHoroOjBOTa7nI36n5KrEU6FG3SsdeF0u9X3dl15QPM8Mx6sUpkBXiy7o4rGfZH4ntp
PMrcOHL3vJLNgOOnT36sByib0oFa95xx9aUc5CikNs0KydQo5jwW1MCc3JHmEi04SumfMlpnkrjd
5hVx+XOt2uuGniAAX6vq/XRXoVbqtouuD1LRP32DR4KQYiWe5TS1Qy57TnJd3uirGpUNyFgECKaO
KGOvKEpvL9o3hJrucX/UMFTxcvFHN2J8RCcl065wSWVQbTYUPvz9QEnr7QrDDoHnLsN/HvvErJRO
edA7P95Z8zwR+cnhMTiJywYe6WfQqXIJiHrCpPDVUBwZsQ+YXjLazEYbCVhAUbJSQqT455doSQvZ
QVvf4E97xXjzhnU6qu6Rf/ZRFOZa+l9lAaO0LylS6JwRJ3+VcouTmbFHy4w0Zy8108MOKHUdD8ex
94TGwJjaYyd1eZMgc+hmaqbVtGkNn8IKWnTFy3mlxdKrAGIKKyJiahi2MG9USjFtLHK8eElBQPPs
GLxHbDeKM2WSWPge3Vn96cAKOaON+KA78n7B+QrxSSMj7ZkXYrWE1kXyy51pIna3zUtqUOO1MgJn
f5jBsSytMTl24OBc65FL47c46JhfggbWPezN7VDkDxku1zQVKRRp01tRRQcZAt2VQOI0Cw+Ma42B
BN9dz6HbAMFp3ByQBjJMAGlJiyitloTYx4P8Fc6HGnXcUktS4fRy9iIFLw6d17BUOiXUuSiPCmVe
YKTMSOR5uvGlo/fYNs6Nywmj6fwUe9YZ4ezumNpzLlRyXPddwaiAXktqIOxGKlQbQ3ROaEsWjwAd
lzH+43XJjwjQGmCZifqBZBdPv+IUehRNZZpIHDRV0BuCYDrNaStTv6FwTOouTF5JSRzibVFMalVD
u5u6ZGxKCOplHXqQN4p6VDKt2AfgTvz0uBEqQvEZSIZbfZ7CTEroqH2QaMilxm0yLQosaRo0BsLf
r9ldvSmBT/6mWYL80zd+EXCNvgOVY9IpwT4zvzIKTd1IKbu70IKVRmtAm3ixd/gtXssI532kwFyu
QmorRbSc2FGInFNiBUJ1O1UI0BYbnndD+gCO4k5bOP2NeoBoyE0uhMyZgwwAH1ZRLWzE9cYtN5Na
b82t6/82I19hTiS58vmO1Okc5B8g/tli0DCyH2OWNS406VgVN2cBxRFGIm2rwec44Lh6tsTnq51q
Y7NFQMhiT+hCNj/vzbcBd4xwxiV266LNxkVd5MGkfAnjWhoezdfwIuuD3Jo8rFTKi9qMMudYQU0n
abvkLFRB1bSBMdQcDHRfit0mEK2R/6qChZrlEN8ssHv5/rfaCJ99jtieNpMB5NyrxNeGCggCzLYv
D7lpldDANMobidiXY20VODhs68DxkLPBtwtCd3fnRAPd46dGL8qpGUpSjcdO4lSulUQciky81xNK
lJR27vhwQi3ikYv8Saxk+N+uhzRFddaL+wz4ni4FnR7FlpcSqvO6v6sUSBx6ohmVMY+de8HUIBKm
HjTDuHY0FMfSuGSRk4XmkVi8Ktas9eh4R1UX4F8IAXC92j4VAx9ngbojrjGBAbva6RVYYPXoyFE/
z4BmmH/u3ShDvqVJN+E4Yz00qhpW5S84+OV34bEKEod9nkxNqcy1qmppDYblpmLWEeZwfOAeLPt9
wnhpegUsiNugpNeWC28gJ61923/nA4+P5PKRo7BIskqH3Q2AB/BTyYkMa/Zg03/4/wYPNQkJBeAL
ceGJ+3CRtTo1UbfqPo7Ym6ZsMQl184BNlITZkjo1dLZ1JGByuBkmOtuzRLsEYpJC53iB6OJO57fo
DtynAvssG0FG1EVTDnnA2K5iQGzLuxeebFtg8bm5wjIRhMiLUKQF3cOR1V+PUg6BcaFH5hGGWie0
ffccnlLH/eMHzzyANBrlyodaN279IhAda18V4Y+uvMTrtAJn8mEa3Vd3eyasHPx/3n7YVnssF3aE
LwSb6ofQ6V1t9WsmeqAwy/f8MWW56cUXBXbhtuiMumhE2mM54gahcAJ58/581IA5+c2fGal1YHv+
fXvkNfkk9TxIO2FkRL+MNIPH9DBPzSNB0vuBNjX21ING/G06Ir9mzM2N/sEopIHFkUwnNCDzLlkt
evQ4DGKQyphCGNuj6r05WHX4Y7HwiunKgNYonehT6Q6Q8uAlTT8dBuKyuhYUxMN0V7fac6HNaz7x
SM1y0Lslak7PPxfRz17klCVftM0v4o4oyec1KHkPBlYvg95ja+n95FOWHCj31X+Cyd5MGCNbhvZH
ysVTQEcxlYDo9z0MSZUHJBZsCDbclE+Z+E+IYuIWDseq2P/SJRqcKQl50km2ku9DSZ2P4Uf4OJC8
UcDXUIfgCbfGMh0owLd5Iu5mGkhn3AmjEHl9byMU5u2yjF1OerakMO11kBm31/MelbXAyXmKx0I6
FWq5SlxdBhOue69lCStRrCJpDLfeTabxJVgUI8o5fru+EYcq6Im8jewiFPQ2Foijdx2yM6IKi9pH
0X0e2vrBkgsXQZNccURvw7TgnQgqMct4odYPO32iatCJyFuf6Qa+f4nsAshEtvrBY454wpbJoAjf
LegxpzIg9sOzJcHva0IVHWB7PcSamVnDg4VAozvGZnchsyhZEJ6iAtoWUgJfTlQBSEKa/GBjGXtk
4I524N5z2Qtg4pX8NWWKb6c+XeibLXkQzPGIhW03/dMm2lGbH8n5qYU4hi3e5Q5GWUqCdaR/I9BC
Xv1VA3waZq3f+QG+B9hc46uVVEAxArfUF6m+INDHwyOFSwZmyitkYo2wJoSPXhj2zL6IcNo8yU4a
Yw3EU4W+JFLYiPIsv+Pongo8ZT1NyEkkCUQISHuIyw1fW7BwTbuYjY9sY1EeCj6uaBMUx03noIhj
fVkrHC5+BvtiSTttqOOEbUkp/VO8oRRhiHHpcGMFOa4a39SB6KAc8qLUOF6ZHZvgIQnAbtF2xUdk
RFnbNaR0yvyTGwBddokQ71I1e/BFFv2orixBimdidjZTv0nSBzGp0jwZc3T4agyvuoYoeA9S+i0N
cS6l8auXNIbyQCQilyDm+6NNe0JIhWTY2gJN7/Wwl3t9emBhIbKq0jF2E1aWyL1q6w4Segvt/Mdn
YbxQngUMd26R/XCbkZoGLvL44M6AqnscfQmlsJac5t65w2Kc8nnALjNrVCAJlWk9feDcOfy2CDHe
WAHahlLNBnYvPlb/1rLZ2nm3Wa6tKyrT5NqFZCVW/mNSr4K9iIwpofRcsqgVg6vJpbxFw3pFzvob
uM9EO7WvO7IYOTTK3EI32cwKinPu89SVwXYLudZCZwID9qymczE+doMWXSTYxcafgYiu0lADZgtL
H0LyJXaiic0mgSWf5Izbr9JEXbIVv6srrGZWPg3NFgsC5FWGiM08UdMjPJQRkT5hcEqRpmXJ0sqf
XZNzdZRhz6gFEtQXtc6tf0Sl2pGDyEBRIdAttZgJPi/EU1zAn+sfSy5iZJjhvZXkGA9XVEpgYHjq
uY7LTE/rJtT28wjQsI43evmiHXtX6v3nf3mkJd9dv5R/xIAOYbAuysJb14vRi0zeSPDj3DNzvwVh
uey39DT8EOf6TrteYkNSmlE7lGPghMGPlul+ohgT0pOdDRqz9JhqqJMIhI4Psl/2Z/WvslKBojEe
WQaFQ5yCw1mdpzrDdk7VbtpILCLcIGAfhCNuSppxsvqYWLiCu90W7Rz1tO2DXyynih/yrdKACVrm
N7v+iE2ZNLqw+LASfABC0uLKjlCzPhtWHgO8VdnXBvh+QQapGWOZsbxE9HHrkg159L6eRRGbFgrF
vGrEW1I8KT6xwpovtxxwPWsxd5ZsNi6WDteHcGY9mexOD7R2oM5pjvf7zSo1Uu0siYI2GP3eEeQO
23DD+roJNCM2fmhx5suj8waVMQ7eTcDnxwYvFEGvDSSgBfALLJziopj8Rgci/vSoVSinHnBpx2Nb
5cT2GwP/2Vx1WfVtKcIUdo5XWP84tjTCl0PPSpTDq/C7rO9onAPl9l5hBv+W2mqCuHxEADkq5JxD
uSdSdBWwi9QMdYnGcvMeMTcj2+ZEuzZ7bMzy95kxXt16bM21YzSuAKFg7v1+EpuiOCOGJyBNmOUG
Q8H/rcPoBQiXoyLaHh/Ieyc5P+kljG8DKWhlZs8/h5/Mck0QoH1jyCFPtZWWMkuTxwqyXKuwXvxM
8r7iGqbkfjcocusJywMd6ybwFqQrShuQL4SOeHoRHuWczkJeaRn+jrGPqzig/znA21G7xhzDqYrg
JV/qWKKVt5hCnqOjJv/xG5U9uD2LbKMDLFu7j1Q5AOLjx0UVxFNNMasVnDXbH6RsbFOG/Kt1wApB
4v0Y7ShUAUJjXZCNPCzKn4/N42gXYCHHiCux3J9cfhMuFYWjcYzixl3kQZK/B4D79vWonlGi4QD5
1ztZmZdTv+73D3+oC2YnCtgD7ZMO+2pmX+m86WEh+eZGaK/Aaj6OhsNfpJIitnkaE+rKPAvWjXHN
luueF9KI5V1RN16J7X9/A+9dauo8kfuZ3EtsTjlZ2ngH7JitGqn4v6lt1pcOLwPm4kTX8SnqpT7H
Xr2rnQSNaWsh7nmVSI/DPav1DYX3XPp4R7Hp7a/IECYN4iTEONFvlwSXbdnAKoTj/PPUJfsXohPO
/TpKrHNFCMAXVVRtePhuejYEHYn7B9NXbSlizWDvYnBg/BhC5CohCUtN7S2WrelzWSkw416f4fdM
nXVJ6rfYtmQcpuvSGfbGKTOp4V9pvOdoxaGVhJODGM9FOKo+Dx7ek0ItAn9GhZnewjkjMW1jQeAy
QiUtOOqChXL5Yk8736+AYRRQ5wiRKJJUt3oYNOGxgbZJ0KFHMNfh/N76cd4JPXh7znzkg5RTTCnQ
upO3IsNFXYPtrN08mkoQaMYPS1djFsZ42ifldvqW8/OZv3x/HiW/zvuTDF43bWNE8+gXTonBHyQO
ZFaSq2PwSnVyJzJTbqCRs9FyEDelNS3EpyT+6p+Z22lDolH53pKtOM/8Muc39cibOkafpnwojX7e
3v8tQH3+LpeRAQFcnItl99I51H8le57aNN/L/ZgzREUfqKMkZ1KYoqNg/7W417FMZ6Nlturg7q9q
x9ypdF52Gf/CEZsdwv36HpZ1Om+JELrBMwkQCp08igd8CkrwAFweXy3OMPRzKfCsGX152PTfXYWX
M/A46rn+LWrMGl4sllfLUZoT6IDcAmr2hyNHp8/Im96B+jkRvrxSqsobyjF6+AmbUo5ZqCR5lS1i
CJjOkYFVmWaUK4oFPzX3JZL+zi9I5K5iuBHakKT4UAn1s/weXMIVXHwYhb50+JdwIFEvhxcz+BNq
g9ttj0pwXhCBsqjSdWCR3cUx5N1o/1hX1B6UylWgdnQOgFSFVqr2pZOwUMMY2DCeEUlMNNYhoU6C
KRjRrKpZQCRpHh2gohLVrCrLmtiGmqzfGZOi/Uc/d0PABPa1Bcc9H9P8bKAlpB4ZLdBqdp5gsgP+
3U8kwrtg4FDA2qR1uQz5U6f5cdWG59wcOaiCJ2FPCI9WU5r9j4zdvWNIfLOlX06lBx76HLhwtbDA
A5Kkh/eGjPFen8A8TlFcfnHa1tpAuB3mNvVdfxscbyQYzkegxPBMf30pLEA4/mQzW35qv7ytHe/0
5HltnkiOvo2B94XS2ZLXGc5OWPPBuStkhiceOcFkt6PQfUQ5wpf563Yy5WpD2tkOx9Q389OO4Gfd
p1qjGdp9n29G+d9Drq6/LmOZKOA5S0PGsC42mME0BPrJev2ap2tb14kJxnenLTRd2HogQ4UD+qbM
AHgzsrkMQ0jpQGuDbA6RaOz07rdFeZRaitWrP3LflZ9B/BL89b3xguaBtDoPtYirGGpz2nZPbxpC
kyLdlvxGSiAGh0+3DiFjZCrbWsJhsJ8Ov247ddr/Bonb+vIu8eOJk4780QysBrtqTX1MbTIxnR8q
3b/oD3SmrA7dLEI9NGjD5YGoNJGdDxk+QBXnMc5O/MvdWx5z3lBfSo8VC4ejt/qY9xAswERjwXVk
6DN+zr9WSXvpnr2G+mhlcJZ5SOYnkflsvoutnMhvCzZHjqTSGhwuZPDIcwg6Dh178UEZTi+//+T/
dKtyi0sutSRzVsz99YxSxUQPV6DN0MwrRNctQNb7MACPLGlTde/v0dduvrE0pz+J/VtXtE+H9v3D
zPhT54aL/WFAY8PcfD8fJB6h6NTzb1UsSBJ7sBobd+Q2k+yKVHlyS3p0RAeWfXK8s+iOWtGfmV6F
E+kIqdkEUeTgeU9xy6MWf0q7DewR0x7wKO88R2Q+QTeEOHbz9c4uboT52KDMkUK3nhgdMRZ5hUrY
jDmAemLCa2BacYb3+pgIklzOtZXoNPNw8zIVddnvBcKfvnYPc0ru7w4IjLmi/feeeWaeLYVd1w7o
Lj79WxF0Z4WSIslyidbXr0/lJzdJVB5v3Rqu6N2fjHbjEVDCm6427QX6Soc/mIwz6Yrqu2LYoPKK
6/mSC2K5hxahZta7DC7ud81xbp1WDcWbu+i5GwWD5ifWmd18CBBg9OVQCbL+C3WION+rRAb7Re7H
JNDlZMWqi38kc7BKHgcnadT+YmSJr7NSRBfanrkLEqwjJVUJi9VEWYLWgiGSp9vcspKdUpugFnrc
1KeM+dMWfg636hNs3/YKWR30npI3LHJbTPaKFeJ4LhglzYt0JvsB0okzgahxPwOJWTfNCHU6qsEj
ROEPXdsCexn1alhpqG7by6KSd9CsqcAZi9fQg+orvIliWusdCv16pvZHvNMjDHFqVLsx/6HpZBZK
DkuWWJhVkbhLCnIDujYuUd44M9plOG7RLS6sZn8CGUobN7wBVxPpATEHj2caUrvuJQwdWqRAzfwZ
aHcl1wLDEoLI4b7se94uN98vZVukHK3+M/AathbhKOuZ/AMUjEMH0gCkXMcJFHR6bCgoriyE18xI
0vlC24pdSMFBKLTaxORfp2/bGfnzxxekCgNZmv/PsK77ETLrKMgFwmdrHSMMw9fYmbcefn9BYRKN
YN1gn0cj5+eRPC8g6k7/7bCoIt2TmVgHA0W6rQ0s7bq57aM8mqi1rq19bdskLkZs1t43clLBkfNN
nsfLXV0KA0YvvtewWI8qKwY3s6DD0GEjc8/UDB2mLxzLFOJAQTAxWhmwttrsmtEY4g48c/OlbeKa
HeeE4xm/NnqBbN/luJ9LMkXBELnISXFzIbmv9nf1d2fG2dT+3DdWNX3IrgGYMSHAUQzrrO6M9rr0
ke4rPqQKdInAh51RwzjY7tCO4Bl6zemRQ4R8/+fT+1FI6NH22rIdSAa0vdmRXryL3RMZUFxdSJJC
+bpChsPIN5B0LWxvWrJdY3+1LsNBWzPRu1UBZcOcUB2yj5/ATiFJc/dsjc18/Enelv238smtEGaG
ydVcdkgrGxz+gQQ/tBchXFOI/7oKYjyhQgrTT1XHKg08tIiiaaxFSl0xVwsnnm2YbCqcuDIdLn7m
q6nmshWJ9NYd9I2tubaPVs0o+VwVaBNiHWsQl0LJmyDKkCrmIpCwCL0xO+kkatRTEsu2pGDHB1Kp
NAFwg8trRNaI4XJH/r43oeyt6GeG3E6AG7gMseEMpYCvlYW21CMoL5hw8UbozTMvkM+1325Trx/q
IdKccqhEOvrBATsaZGAOZRc/EBirPEfv9ilOH/KpKZTMMwq+nVsWX7uwbCp6IFUbL9c9Tf/yclYD
Y5h6B6TK/a362+CWqyQ36dcXYhDpjwBz20Mk+i0BHPrXi3N0asyi1tIalI3gnBp6Plfsf+nl2WYZ
jCSlSgFFRox0lT/VIr943zGXnwIhyZMqdbqj8nbQf92llQzwByZPiQdAJMOTGNKqUHG+fODiQFo+
6uPFda3wYvN84Kzj8vyYzytcCeOqjzFGeWxCdTFBWLIlArVHTseI+lViV9O/fi2cINC85ItE9hii
wAFgtx+ehlee6whM1SXlT7uytm7VsM/fXYsiYLbbNmpgR8FM7U8I439xuDc5xeNcQE6MygkF84Yk
AQuvCQ4fBbLTKTJHIWaHuOkbhVygDZneCZw3RhzZnU7VLZTWOeio78lAqaLG29TByMbedxc9PFt3
mB3pzzG1Cz/X1+ELB0TkipHQsrAtNx4m1vINnbWuCV8fxZBD6CY4+YE7A/2tXfAqaUh6Y4UXoi24
1cuhJdu5Ioc/qo1FiC9KON2vpXBGo/KXiikrDttbgpIQPNQosiHKSNGq3Apa5SSIi7F8Abd4eUVa
TLnWRd8be8TthE2IXVGbfKN/ihCDrEqwUSqgP9ufFInhml3QLZbhcXoguMcSCq6rQ5AqLBgSzG62
QJz+ERFm45Pxyy24ngHFu0trb8coEzp3uEwVZRA2G1xVHbbexLkApipnZu6gKy5DxAjaGqNdVNt7
OnplHsVca5S6tR+RuE8S2TLOYvUV3yJPL5QX2g6wGVxfTwamOBKvaoIeySjjeGOBriMLovVw7O8j
YO1NyQ35RiIjrXngBsIBkoYq/KNgeegWBPr7+DdvPRB6ci6aXM18vpvCCB/15zugW5gEB98vSotL
Bm8Be2BB7S4M2UhqXM6qEzUJKUk7vjVuK1Wd1RoE4XbFq7TKIsrfFKx4S8OhIrhD8R7qlVLL7pI7
+xjITFbjTKJ7qAVjBzyT0rz+107W5pcjrlekH9ckPF/MyIZ0jNkIOurTThipuZfCPfoTaZUpP2ty
vwG7uToJxWrbVi4yCUUfm/uFe2aX21Lwwiiew7/CeYTpAs1h+h31to/ET6ZKEQ4PVCJWAY+OPp9/
8Xmn1qh4UfXHvDpS7DR8sqvLYTykprq1cw+uJGqAaQTcMvkbtyzoZ2bCUWVDOVqbJgjO1RFesJrC
PpaHvETRDiJqnkndZ42PgrCWY2SXikNsCKkVOTsl5f+JUy8vXAGWMKk9/dwg99vt2I5cdhGSVKMH
1lpiZy0j7WeVeYRhm5G1T9yf4LNRUDPfqJ09axMOiZVRlJ5OBPdA0r22Olt+Ai9ipIMuoUz+KF0r
ZdQv20zTONJl9oV7Yf0jEjBJXvLdolr5vlUOjqQaA6HFHwvqQn/Y0D5A24nut2MXGPeh6ly2R0CG
LXrfjyoA0K4aMplW89jWV/0YbZ6ByGVjOvNW+67Eil8E5MbB7japVpvSOiOXBq804lvBc5xWStct
PfLZVBCIFvB9Ns1Fk7D1/XZednMQkPUavGS4vkbdmaY1WaaF5XW04Fv6WQdO8ay1p6P4wWSMfCh8
JmkH8c0Wsyh2SfT2Fsns2F68v7sjmpMK+HHRA4F4vlohuXkbw6o2z+7GpQR4lsJvdh6FH7D3mPMy
ZmJnh93A1ehrDsp8cDDclYPXxsf0vLQ/GQ9XtV+HPxKG2u6y/ZKphnWx/kqIAAc0CSqVMKOmG0PG
jbTZEEJnHEw8w3N0THj75YcQGa29ZsTQdth9l9uAr6kQZsOKN2DkL05hBGJP0NGf7AquB4v5tHEL
wWk47KeknBgR2P0vQoxyuBpQYZuXVv430BCms+2PYDv6zn8z6sed2d7VRprr20iUGuzhEsQlJcr+
7lDOL49kFX70sETxu1Khs5+ohMBFx50r/egRKaawnkmJHxbvNgEdGV17Ups7ixV0jbMPM+W/UUVM
9l5wpQ5Up7nA4ye+sh6+XEbjepOCXak6Kzqn8e9ulPoE6M/40fSxBAunUQquM9jksn5AMHPSiZBX
85VXqhiqLMimmw/2DAZK9eC5LwrErC5gYvNlTYIxUTxjHMa7Uwe8ZxwABtZoRn/KKWWgC9wt9m4x
5IIHWkKV3MKJzyZp1aezsfhE0zF+jEJHzOAlT/y+v+MG19gCWqKvESibSsg9GYtwaFJ7i4I55uXk
+QVVCThLjdC9eifkg8lZJAOW+b+/8iXPVQCqurLf0zemfdRAcopaKArF2KFVQdiEwmrT5Jkko8mQ
j21ZWTLzcTRA9yHEddMH9DLdcryUQ6CY8nCF/NWSSMciFrERvgn9EsgtFj5EBZQzboOm1woecoMM
QZpvzocLCWh68atFs51frGOyA+6H5aor5zC2aQuYPxmldNWXGBnLDrFJS0HEE1SHvhgV8XbIre96
/5h+x0J4s6MbxecpijuOvv/NuBessZKdoBwjJ0AANZg3YRhzu+Ba1JQDtMjQ6gPwRa308RNzEkMV
kMJfDaf0mS804asSUTH/Anq+dAdmcpOVeX2QL8laJVSUMxs01uHYK24RtjFsT3pn5RQ1YFDEKHbV
yJk3UqicGWO0iWtX0WRbFQF5ao57R9X4tFvn9f1U1P5ImmcVxdtxJBgeTc53D1ExcaxXQi9/eT21
iO49BgrDNK4R6RsVRiZpWUQvI4iq1Zzh7HIMD40FjvZqK0FhYxGGmXG1usGMpOaixMvgi00Odh9c
8mSbffpNsfRorGe7G88OHjj6MlohS0z4GyiNkY3BrDr+bMWZn/K+9kxaXRc8vAwsMezblEJ9f9Be
xhHrCIK6huIqhzvzYyZkv5Dg6dFapvgpNkjAeiLH1GxysGtVkjnWAxFWu3uYwg/maaT9NnDpk2cU
B9f9AniNAiaYBIint+lPPxjVMuHfWIi4MY9Cfi729KxVhj1YK8MUzs97YsSORztvDgQbYzCa/eXk
xAhts/0Ucnv2irb4irAQLYLx5O5j56I/aV5liztVVu1V1pRZ7tP+W2ZWOAvTPOLUGYVTeA2A2pXa
faOhsG0m+qhWxL9ptGHbUy51GUXibQZpvnzbCeDDgQWOgQdm93HVoD9Q3HG0NG0CFPIGfMLAT24t
nuwtjQH9v1J13mOWdQQVi3iEgoxuOFkKMCqJ3JjmiIvkpKIPkbS+YMKhYbIJ2+nQaTxniAJ44zvB
ZS4Nl8N5f/DkOAUJwjXLMEglkOUwxsMt2cBtJIqrMX7gkJ6ANB/6vz5v5zLYgFagWTA9i9ff3xJb
volnOTBQ2/3ixMzvV3j70mKVc9RvOBwbdOMnE9RCiEulAx6D8+wSoahiGguq1IvSFAonoz6tnT/8
JAFLXNkE1FmRzifcl3qSMbke0eZnHTR74ZjLsi+5AAsAEpnK5UU/gDbx3NyXDVa5u8sQyP9XS6pf
vGheGnMt1CR8Su9PxcmSubqcMeuveuVC4Hz8QYc2NzodOOiww4StqdRJwFikAmlxe/mlq205XUwA
iXuvwvyB4k5X9kTCVr7gDmjjj5kp6WnRVdRmLYpg3EwfiwgAMz+wRTVca2FYky2HZ3SrNSaEYNac
go7bZdslt9Byxrpa9BYRH6zDhYCzSBKq+AGo2B8wF6ofG2c9CWCJ9NHdfC5ggDtNLh9nITtsJn2I
wBlPTPHCK3yUMqhSvLN6IbQMT3CQhlIEcK+Ywav8VRsyHRlQo8yO9f3YqAU5JBSqiWfDxMlkqIcJ
OoZKkeEUxXl8fX7qK95uNDN0vlVn6skjxcrh/Igv68rcDOkxn0JFXmMSb9pdlXPoQKdIbkuvQ9uG
IIUsEAFYqZyv5heo6uG/pWlsfrStP+KJqzc14peD33R5QPz/lODwDyzHUEOJhGfSZ4zM0HwpqXXb
hRjb8dRC6M1vSYOghOZsrAezwwqmIOTOdzEk/pRbQ45/uZ9jg4nO93ZuzXBLUqspY+7gKAVUrfoY
096+EvI4sWUZ1hFwuL5TcbfuJKnOB01BU4pPSOF3klP3ZQuz4qkkgWfncNEECjYt2/H2Y80db8YT
CeJgQ2fuw4YMxL6JcIeHu3Wbao+Pyp4VRSQC6kwgdVxWlmg8qtzQ5oMmsqRf9mkuRUWGOW1RnB+S
2qY3Zhf10Yi79Y+sWNAL+6ymr8Qapjr8w893LftdUe13k4kjqb7VXJSoA41ecxhd1tZpRN1C/ofy
TOdRhBZnDkjmz9SB7KgauxXU7ltbOJF6DrathdFPopvqjZSt3KuSe4T+CnRN3BJ7j/1LklASbNAp
HNkzVsJ/g+fi++2Duw6rBFYFputOw8qIUaaiFJmcGgv4QJE0LiMR+eHdmJjlL8YKejinFSIJWBA+
Jf+GwjW28EK8E+CPVAWMB6KznR8v1RQXTYJHjP9gEFuRUiwQ/1a8cTnZgl53WpAqAO5WrBQfzXn2
3bZr6MUsLvEnm7hZlv2b/1TQn9cKCve0JatTw07PG4BnedxcSSmQjmo23BXyWbcFaLxIXQdQ52kX
LRblFFL53WS49hEnL0UsI2wNdbmUH6CtHzd5YF9Wpc10+1T8N+voy/kpVV7KKHjjW4NUfEcpG4Y2
9TXrbXSpubWkrHH1mgdW9bke6YjE/M4KvphqoPt/3q2QOyWTjYbvZSkjd8fKw3vUNdkBHZRYtAno
JGlkx9ZyFMyzNH5gQXT1eSlvPB2OprE9iJhGF1e0XEugecYlFpGq2yoUiYGMUDrIom1E4ffCRpwk
0ietO5cPMriWwY6TyFq5AvhDohMh4ets56paCNW7UIODXJbXgz2wAuwnEfixSVyuH5am82gDGdtv
a6XCTDjSqFqWjBFGoMO6ZI1wxA4aaKpbsnDM6jrXVtb8l+paAxSVvomJ4lujzh082/MBKrUhO0kA
jvoF+5UMbZdM4YGePYo2/V13OrVAQSMvXFqZXhbyw1juG3rpAbT0kECGfO1fGCfQearaAekGnxg9
nHe2jJFVSJfQpFnYqORkZ5cDU4ighS6Qhb+QXYqRV3Me1Fq/noMNPBpb9owv7SSPrI7Xo1ubiSrW
0gGGox24tyAxxWj5s+AC2/cfuRA6wNReu072Fdx7M5pEsVKb9O3PGcT1G3PEvNsDdAk8J9sloikt
kBaDhUtMJGxZu3Oyjvo1RpmNSCTZG/rZLlG5+eZPehzly5dEG5z095J1kzgVvgmv2rF5G3cOInRu
QIAhh3r5YIprcnKFDOTvXx2K+FMbyotURcFUFxcJtdJGtbbRKdwDE/4YK6n+keW+rLJbcJH14gbs
NZsDCubkTDlXDtoYXhkK+ZQM3w74KmgtOmSORuEFZaFOpXswbb07ZlpCR+5MWVPnU8r+wosOmfx/
0a0MT6Tp+Zafq2HTDEDdMNv6mgbBlZKUOyh786JwQngoLxq9oeURbaAZARxnzMO5GBL4XEzz1Pun
kFW2wzOaC9bVeLcFtqvyLXN7MVxmfpSY9abcErhwfyzSqtRwK6asQlv8XBCbvKY3TpYYFBT37iDV
QGMS/avnQ/REDMlugPjsS9ZuIFPEcR7NnfuJJDnAmaMBFNVb8zHWiQ8b07OKPZmCVz5x7yXkFrsL
5yJSfD9MUCEplapkzvrwUu2xG1SyUQZwhssHcSXH5E0trRr4eLO6QhH+Z7zLm0egGlvz7JhwhFFq
ruBBNiqWqr/xcIdRTP4S6qm6BqTZ125fCusilGATXOV1auNotkxvGo+uO4hpuY0JHvB41Ut0Km4n
L7j2VDnyQDvsNEvKDFgBn5S7INMvuZUdTM8NdEfURcrhTIddFuiQXeNCfikf9q5kR1vO8pIlZVXp
o4WNRXGT1Y4TMwvJyZPD4dCVOuCpT4U9fIkIOjWEywTa44HD6n6LfiCU/uOq967GE2H4kZnls2o2
lyVH5Ohhdal/7ZiYQl50oFZiAPV78CdCxDgiV+JWUVctrTh6QJ40eBhDTW+5Hb9KkceNI4SYKyqG
UcLIch85L0KvfclUCrpRvnyS0OjVzU3RFz+s6b9rpELWNDTijG1ifcKKQm/90JgrxJ1xIVF0ZWgG
/Z5jHnincWZqWKUF39B7DZ8b/Vb/G5HUrOQPMoUg+5FZZFc+Gnc+1VSm/H6sr3av6cisovzqe1w+
iyd/x7tQcp43kwd8tfjKJsjvEx/H5Fm0mw5A1TsXzXbwX28hmcjy38yIouCDBXWZr4+YRk1gAzWu
QTW9Aez17t9tUo7UyDwy7/qWRzUlZUZHhL+wGxGeeBEMK0RN1hxDUc+ajPI3cHihCjmrZw1sflub
1i0nO3AegtGlpmmQkFQrhXqpSbarL6pC35Y6/lKEdeRrFEwSv2Yy1b/hCw/c0GLarZ/1o6qAA9sX
aGceoPlL+57LJZ9Ku097fW5j6Q/TB+vrq82iByucU3KQqjlIIqTYMFb/rFHjwahdlHkzy3uTMNQK
w8CbO8PXAXE3HdTUM4YnSwTlMrfzo4W75kVi8cCIpTMWtnUAk7u+cSdVCBnpW1mQqCybVVURefiz
JAETFYqtok1jH7hQ2WJMZ024AOTlfh1+U2R3+dA211oSmleT5q1GuF6BakHWrNcovYG0rrzbw2HS
WAiejLef0qY+Dx8ZHJX5rassIIQNgxh2eixdW/pNalhoq9eZ4RsZLCeej9M6cdPgMJgVcOEjKt1R
ZeCFdS9jgENwXy8qBdgRr+Su0pSBmfyMhEmQKe3VHB8jSStKeWzCwTqcg20VEZA4/qRa+PtuxxbQ
UAj2oUv9wMHzI32zf4F/C6qwq/OjmtxByGUu4WOIQ3SWxNmY/0uG9TQIUwKeYE7DJBn/aKC+gJ3E
wbLdH2GsXgkJSLnDzU6o/ojoV/0BN0EsggP85Yu3S06AwVrrB9zqa+CrabZBWrJBEaZvOljHJ5hN
BGKb6Bkk/FTlToTs4hKbtTbNL67oVYLjuEBzDVby5mISvODOT2Z2FHgZs7OZigSK6PON+xXmJ6WP
NAfvf+tqJRH+/szztS73rCFE7W7Aq60qckA6kBv6FvKT+iT3lUXDE1ouOS1O+IhwB9FY+1YD+R+d
xRgFSAnCnOqwjMs8T/kWbKFHdekw8Usnwahhwn1bAM27qVhYBnqtIhYcdQb0rZChbRG++cbDlAhg
USbDn4wggY4O/Qw5Aaf3+nFequQO7Jry3Ek+yHw/Coadgc95szMrYaO7c1F2IgNEhcVO8zYsL5vh
J9DhmS68QyUeFlK9lACJe32Uhp/BQlpxxfOET2oSDVfVlEdHyf0eHz8D8RmO6W6XwtdN8FPBj/MF
kI8ZZRYAEM1r3DVwZDP/DpTjapaYgV25P0vAR3hCqu0xlbIaeQIRuSAGh9YU6/SNtO4KZ7jcr6fC
3DFL0TeS3p9SLb7HgYpgr2n2H/0d23PFEqoMSwJgYbaQ1stYh4rNDgGf6wiLNVrltU2e6xBrGJ9w
YzHRx5htbl45e8lE/Rc6unCzWDLk0vUT+3p/9satMNjvtCqGXZ32o2Yt/LEVjBhzcYMYfIIsnmZF
WhRhJZ0uSsvOl8WttTWvdleB2YqEizLptVJDez2utacYNZAgigLQeaRC8KSdnv7nSe5PAkF7c9nn
2eJxAxG9OMBJiN7kmBIYfqiT6q5MZ48V6XnoYO4t44cbzrWHEzF5IDaMEGdSBF+HELOT4M/OEG9E
bJKybY2xjU3q0gRNjle+FJnjrePyftyvaxmTTCueSzjmhbLHizFS0+7533Mdjt0FwYm6quOn/J9U
8NN9eFv/g2BpUA0W29Gm+i4udlTCMfwevwzB3CDi4+K+wKhiecH0d7dBHw/4Nwc5rlncdyOHS8JD
buQGOh34oli0lbj+O9GZbbXqLJhNyOcytHpfvDThm+XokCg7VfHpJc2HufY0hJfzaSmLrecUI2KH
lFCdPTFeplRVrGWMBnvtl/l9bkca+tfgaBxFk1nfgoi3cwn9/Jwpev1jtMGoabeyyGRcUVL2p8eM
r3uZ5R0QnJIXaszDPCqq+vxvQCpSHtdH94iUNcwD4V3ut7+5thuvaMa4RfPAw8RnFL5D5mcnGvmL
rlCNErsm57pf9TIyCJvREXTAIVKlNVfWd8qrautYMnPPMgjDJynjpuJPbJd/T3FNXJrjh6BNSAUo
gwaNEMGODakDrc7zWtnVGpeN613k5EqpFw1nXDVJGtHAg0frlYnvGYOnXKM7iXqW7wTE5mYGIoVF
SQcvSexBjyNWrf/quP5SynNT50FvLYLlCwVbsjsprrrezLemF1Voz+MHLGagplsJXmOA0splwm/O
Ce3Kf0PhNO1xsCJw3ntq2ERPgr85HdUBUGacmJ+gFAI0JWixAskX2tRyLLhhA0L3wOgA7sthBdz9
v0Y48ZXI+bCz3FSbvJJPalmI1z+pKCPyHPeii1KS/Waqty0vH+wdBCFCKRYEOPqLCdL9PrW/o//R
Bkp7ia+yBNruE0EMLhOs8JP3ye8CixaML78SopMQDeoUWJTq5rnRErBpmq5bTtCCoHLYQ2C0g0ce
gb3Zvk6EneqabQb6NDT+hIizYoiqdCgfJMuA+fo2EOPR24BBINb2h9Wn9cItKVzR7/BiJlPpdLUl
iHc8vzLzQ4OLOBGO1urMkCb6DOPWsDrBP06ZkPIWjhwhIBnfaLnlYckL6UP+1TdNlLQhj1512OcG
nfyouZ/H7/3AGY3rWXqlUX1EtmMjHRhMVCRfx0/TjU4RTlIEHf1881IwQMmeoWKGae8BTfUhfNX5
Oe69xI6VQWWck1ab9i/6XfT319FGvfKvfVIojYF2QGuviIgk3lO32J28rA1nyut2cegzGkrEDH/0
by6CUkRsR8WcNTmKI5AeUiejXywOkDvYURF7NzVxfZzx93fxXlSrro3S8LOgaS6hkDnmZsnt849+
ssBJF+FxQHnXTXldK8d59mI5b7zunMJ10xjBgMRikuDqF89dhuxRGLQOC/4AjFD9+WdfV6AFRdZ9
vkToRR0NTGC/eoSz9ThDAgPgepPnkOkbAw3coqSWObfcVcg5K0YjxziZ3+sU4YqhIQOt0+Z/OOyy
lkOBKXLvW+7mCFJY+2BEZrjWhZx0z9mo7bPMipuz0lWXNUARcKHm3Fx/RMeu24Q6l1YCa1Yf5EMt
0Su+1DrN2ySAo7t9cDhr8ErN1TSdBCQEez+ov4N7hHfuHHx3b5YNYj0pDYgaUD6gEAqn/j+9BFrh
EbV5Yf+7DMEhGoCp6dM6eH9bmNHxpWaDCJ5aoRGjY/ogilT4envVuXPd+tOeqmH3cWxKLpXCAXZN
opKvK1Jt2KLBvLXGIdGTTnW2lx6g1W06E/eInYXuVrIlyEpY5us4adMlytra5niKWLGIQ7tllzG+
FDXJV+SJGdaXEamTGQYSb1jlf8NO2JF/q83BIzsw3vQC8Gj634m93FRcaz08CNOSnvYulpAC2LcR
UCjBxEX2DICCVo3DgBK4d/9CZPLBz+fBQd9O1C3+z8ykiU0N62XODXZSfwQ4Vg2SxUx27bLalimN
SU5zjPIRLtctq2ROwgCytWYOQF2e77iVj6/DHTzuZVOZ/j765moD+AhXw9fX/1KajnvzFkDJZUxu
s1JfE4wob3JYrSiq6VAn4nQbkvxqpcLZEj43v1S5ABmFyXmkTSpFYkMUa7aRsBsx9aZtthtyoWdX
GjKTQFezWL85EyCqiimkmot47wxgOCbCNHzwbV15ThLxZWUYSBBtKVgfRLgcYvoyHrWlUugoP7YI
Wcb5cNmF8/Kv6qiMQEbLS1iaatTl58AH/NCGu2fwDEapNhxuiE5HE0DmBC+UPCWIcvoWBs0ZEHwu
daS5unnlsQG9tNvORbkOOc9VwPhUGzYpGBVQ22/FyCfoD5UkvrNLCutD/hna8NTBhaLBoqXt2lxt
U0w7TIushpgB6kTh2WMjEpfzVw720qyldtgx/V8/f482jDhPvQaptiwHmsE3QIBTmY3NRJqDUVE+
fSDpnDB3wpx83NuO2n07Y19D6DSDw4muk/PaoxPgfx5RpWjxjFIPYxmTeplt6eATDLaim/Gv4ezB
i4JgaR/OU662LTwZ6oUBZ5gjDQrvxC43wQZvNzBAV2g5C6cyKN/kxVsLBkUgnG4S9R5jMJZF1sZc
oSeAGu8oMT7ctfoaMN3eTbUW4kAtC9495sp3mYQ7Y8vRGvkvXUpEOCozcdmuRC2uesTwKuTONJix
quEGRjyMSPFCPQWaMPLzpUOOqxl1jfH7VZTGai7BQYHl2T12eWAe23crFcSZddXYNNG5DubFJyXi
Q1dG2CCTHZgzUrHAJE2BZjgbJHQ6upc4FjfUUYvDw+mkex2rgE5WnGhGl2GqDU0KbygMpaK9+8JT
ZCm0/FB0JBZdy5+F2yPwB5/NTj3Q/JzpJr9h6sdRmvlS/NPSNx9J14DjsvcMCUBe5xSebslGv1C2
4xllEfofonGtgBSYF4D/elngQMtvW7NczM3FzWfc7lPw7LgxYt60VtIczUYVBJNsMSnEt6V8xZoU
V+waGuefj67zRIGBYv9u97rSE67kbrxyQ5XUKZFFp8c65GPGHhqxbuTmk/3SOgx/vl+LzrvuKTOc
DjJohpN4rf0mSKfSlzYR19B6GOgP23liV8IIpPlq1tA0toM7S8gGjRD5OiHG4pMnrZwQfP79R/sb
GWLr1XnIYES3OSSm0Y0aq7v0JfaG0uJ4NYbN05oPpIDAn+nWVQprOQtfnZM3BuHBluM5PcD/QnL2
D2k0HNCcbOMPTvjfFUORBzeZmz2O4IJJcNYWrwfGmqKIUhUeznuNHAD1bItCI7Iso8Cn+akP3OPu
XW6Lm7Odkj+rDciv9U5soUcZ4kvDtaBvScsZKmT7Cnb3IN8iG4nAFzhKmXqZqBA8Db9dIeHte/mV
ZNOSe6l+UK0E/HAAwzPUnVWIs7ak0ytl42CCyuR5P23BOCPl0iUVD/jCiyx/rXj4tWAGpecYiu0E
Bu99BHfxwl2ddvJhS+Ht0AAAt3E6D6P6a3ZuB1OsjlKXJGpSxyPhh3IkDu56Nl6FTXlsJwN4ua7U
DnVWXPWq2uVvB3udp/EBgV4ToeCIcF+qRVDRyMCpr/AH2wHnCZEVPMItbCytCY1hkucw5Dd8GQwy
KGh+L0HpS3aznopWvfip5sBOiJmfgehYia9IjOJjRXTfOZ4DMrsr4aOLI8KvFzyEcczyyryx+LSA
c7Fvms3ow05MKms23p8aQNcytIkJE1xmBwG1lgd5BKI9khstJLowekG9FS1VKJnqFVoQ8WtGr1SP
oDxRhZQEdOzYCUUN+l7Y3iPB5uAAcuUowboWh6OQraXgSZnHP8H06wArZ9v7f/LmOXOYN4aQgYml
R5aTGvKhh+VpONbTW5sTQGeNRC6XZh0FqmlQrF2JsI1nFC1BU/Zb7ewPSwYiUcOnH8jb/1ztBvD7
66nFXAwUAUzW1L49f7p8+YpCK0Ik2a0mWFDIN0ASLkqdONcQvMFoYVLtaKleVWz3tQ6/IvGEHDR3
epwrKMlgHn+/jk8YlolbstYXQuDt4amAY50JYXbkJSHzYufGEHEld3F7EyYN8neLH6lMGNGQAF9d
Y4YrXgNvB+5sM2g0ZxHpJJO/Uc9GGcd7CeOR7OWD0Btr3VcfGJ47ituGHOhfMGC5JZtNH1NW/UEe
6lt9B+wfpXVlvfEm/KLhHGF2R4s9pjpVFu8JXKbsyMkR+TBMyHwqAVkbrE4KJc/XiTH6ggE5CM6u
bK5wiBVW4IzdWDqj0AY4PjQFY5wuVlBBcgmky19I98jamVrjg4JvLWeJ5wmVHlzJJ9lT31W/QFBh
gZT4SRIxjHKoIy2qQD7TI/+2DSx9Rthck5bzdMY5EE0rYPPZglIAfi7fx77pDCq2p5cQSQ5rzRgX
VDq5hoGgFYBV+FjmKCao8Fph8p6EV1PF5BfMgspqhUZQTTKPfeOHlMSju/xvKF9Uy31WgDLhkgJ8
JGmcNIGsmZIUlLcM3YI8dPxiBSKtspEHjJyib5WtcK0D0eMCdJKDduKC64FJ7Zg+DsohE7WOKQRl
+yMH2P6eP68JMg3qEOprRPfavuCQdx2VOmZmbRC+uENkqV5ehrxQlmLgvJ3OHG0X7cEp5THWHX1C
f/d8l8NN9XQlMj7kz3nBL9cwY/bRCtrRXvUrnYJlXjT0NrZgjAhAfHr5xJYcpDSxFaOsoWLH4w+9
oEpnyg/8zz1vGYN4hg/47nBTXpSW8JcvZ0zvuerM90+Fnua0qxvL3iNkhkFz+GAvoUhVKjoB2Nzt
0fsU9x/MpeMVotSf86+4qRpD4N/Ady1OVFzuQ+7NdPzAPm7lxjbvSIhmvzeyNuu3g9jG5apc1+jQ
+tnBJ84Ep9oUSrq1cfRc4o2kwTIG/HFA8g3HOuGebWPnGiWAKVPwqy7C6G/HRnJV7a/zBtBPzbMX
ct9KTk3553llwJyOHZYLa6sN8ws/de/RmgPjCrFdtkJlcnd1mWfI6rOouUTiAt5CpqFHTsWNbv6T
bisKISnGPJN+gnpEk3xaktKSfUQ3fnZoBw6/z9B+92r7UxjJOqmdECqvfAZGa+4NMMOwHa0IkjtN
dmJOzmhwy8JaEoUJwoQNVgvGs0BkjEOQobZFbfn4i7Kc3764m1QMy4yENLZdzp5NdvnmeQQz3u6t
TyLwc6fe4dFzhEfoXp3NgkfoDBgLTjx1oQcQIaVIHmWzqwL/mr127On85PFBeLuiliVGjmmpQ8BH
ccxb1W2/APVU/YhnvRJkPsOALNoibkYno5PErx/IGCV0AD4hdfz54UA0yjnYVO4mMZ1dl3M2NJ0F
V604H7ye72XbpX5k9vrHuO7ri3SC+aDowlSAMIvbn8AJ6subHIv6VTxAmqqxW+EMbJk/65fg8fOv
vuXnrm1GiJNRX1Cl73wcFmWlG/5xcETfYewBFBV8NXnFEO/wpVjARrbsZ2o5LtcffoleN9/Hdm+Q
NLvZyzNT/guv7CrbJMc1NMjRGlX8+jeO4dyHfbePtxeJetgYuqPwt2UU15gbBrhDf8KBbKU4vcw/
UV3A77Sex/63GOGEZGvMcF5CXwXM9WdWHAaYEfmO0VtB7LhDQ7TK18pWW3VRoAySkjo5rhbry1/V
RKYG4Gw87wyIS5spMo9j9Oa/Amgy2O7ztpcs7kj5rpv09o7jDcKlXBZv5mKVQj4FRWaOYHOXpTib
UKP3hHFYQk9A1wPBWGiMI2AgWNHjbHR0208DUZN9nRjPrSDQKnYXOfR8Qc1URdH+F6urEbqMkUP2
tL9fjgx5QyPdZDWNrn3X+hDicZQ69E7ybVgaNEC06ulSiDJlaCCAFOZ8O7ZRZww4gt7+KjvBxeuE
7hyTpCquaAs6wkRIOCD6aab6FJqMZGgKHNPUcvDuwGAgtWiOn5oulsQU0ISRV9emRWX1doBV9JRr
EaVaFN8jbzx3FRAdquvWla/JLhI3aoPcguBOL92g7ZwEwEsMofIkTVUtOfPAYDirvlEzpoEQP4qp
pUvMTWNnpA4JNiHSb+/B+PMtyS8Uai3nMfHJNLTFUEm7s5rH1tyPowPD1S3kCjrx9wT02Yr31FyP
vhuTrEtfGDJPhNHTIDSVzjraEieAFKN77Vhw1xHWGP3AZ/dEhBDo66EfsdIG6QwpjlYKHgLTt/ST
41ThVbRYMA2l9YshIsqyt+bVzKyalmTYO3FHQwHM2zUs8WR2AzJENWoRXiAv5b74L2K2q5pmTC7N
J70Jwguz027RSy89b11k8q77s8RvhCej5oUte86NtP+Hurb7ymocGJ4V9ObiQAhsb/7VbnJ5+pVs
+oArXmaIPW2gs1hqLIGlMz0xikj9w3WY8d4n5N+ZDLsqdCb90pS18NKrC0o0+y3w9SpnDp1dxdeQ
wmtZq6PQiS2uX44+p+ZloqVgOZqYeR++uNatcKUDM/GDxyvMClnszNncBbfFqQuHrPbuiP4KWJ0v
Ht2QUrFwJ1k/lJLO9vWburPkAfFF9UUJaa0O2DxYrq5LSLGPgxrF4gIsiUChvqEQ8FP8EjUHceZt
hIgvCqVgMVITQCaNRQXzlhAlNXOF1baJgTXWxPbVxykx9DMieJhOFYthcmTiM7piNdB0KXQTE4g9
xBaBe+4K8T2ekgn50tzstSKEv26UjGWi1kSJXjKnkAt62/ZnL3211vErz8AXbPXAWYdDugCKylN8
6ZNuGLHx7HP60Z8Acf/GIyV400c9/pGvHEwtrp+0y2LO5Hr9aWBsqo0JhH5ljMbpyjWtW+HdR32/
2RWg2IBtiQqdtRxfNvhdWxCInapRgGDqUNO1lyvzV4Br7vrAzXShxE7XFfUZrOmNiuMAePJxUswl
j9osyQz48L5MMplLHuK/tMbQgEp84d3RdAxvefknbPV25HOnTRKDS7hFopOneLKzOiazL2TFN74r
7+NFXikTSHa9224pEteznk7C5sKvjve0bYTFt/k5wlnXC8u8+S2ENZ2AHJ9oyoZJr/a3kz21ZS1C
bb0mTCvWfeKALBi4q2O2jV7B2DmAII242B/Wsy+RrhMyBimijiH7GkwoG2s7LFIYYz4unRSNrgCP
vmHpJDYjFA6RrwvsURaYlgdgvb1xN/E/MvbgYBrTTXoet3G+uJ4MMKhC6rw06OudOI3w/e9B5phA
5rmA2kPDauwxClHNINBiMs+wIW18DDhAGoVLEdaf0p/BRwmkVsZtriRlrSTUNtzF7knDrgsG+cQh
aNVohPmQqnWNE361SUT5Esg5GrgCNXjB7Mz94bdcJtL3UxfXmjtrT5qVVFQpm/Zn1yleXatlhRte
afu+YrwJ35CAxWznWFWg8JvVWMM8xdnpn0cW8R71rJ+R8nDWwWiKzk5E3kz1CYODH6DcPoKrIa8B
3oS5RQPlotQe3DIYz15w2BpAuC53EJ0ehwShMdS5W7ub3C2iFJh1LMcQqvu9z4UAhCA0NvMPU/GW
kFq5+F0CSIyE55SupxO1R75cyifUDCeq6uBJpqsqenXNThT+2fH7yJIfIwsLb7cXj/w/tp2MgZto
42Lu+UGCYvLXNI0v36zq+z9BKX9oDUn984sL10FxdF8ABEVK5pi4MfwrcihKHGYisZahCjuIwgr6
GKJYn5fMmATRF6PH/h7HVmNLepuy0v3lzz7kn9h2PKpyhDTkwZ9pXRUjOJbPfWbuQbDKo2V/od2m
KDri1G2Z4YlaOJd+dCrg2VYv9ckRlkxweIkN1YX6txtiV5Gdp0p1dDqLJ6eX2+V2GxKzhb4kx6E9
Kki+fjO+X5mRmkkX6rJwkQedr2UkYQEnwLG+Jk/bq2R/AM3fvOCtapV202JE518J1syAkF64o8HS
nsYuII0su48WCRpjVfkeUUoSIc2z9KgtUhS30Eis0dWn92Qg3rkw0Z8gKBscLvpc5cOqXMbXjpRL
G38NEkqz8+ds9dl2iH9m+R68Z/99vJfWZUseP/gSMaMsTrqPY2aQCyV/+2F6+/EOVU0GFVcPvaQ8
F8lnjm71T6tyeGzDwezYINKU5+LddV3gSOT94v92rzDRwWYDZds+kdlPZ0RZ7BMylqCky3duxIcE
3khKV9CNu7IxHeu+L61/maYovnc1/oHODWrv1/JUDTMc76Hlwo2uyOo271ScNf8WQDbML7Zgq4iq
2uJyCI/Ef1s1CGjUajnS+hvNvxWEOY6bkCzFisJL1IG/stg78F6Yqd8yLbZmfcckFOeX5ujP0lwZ
vqbchlcWEvUhtQ/CNXTB8qM/HshQjvXHCx6u7Y0F/uEqm0WE2uPBeFlqzQt03627HmpgXXOIZEOa
yZ8YWV3vnztHIFlLXoeAstBSlYnruFJ1s2zbQzqcJ0F1pGzEBqEqYYWRJAInqB9KXSRt2T63dbiV
52YwgQxS517VRMBFk8gIzi8wX78LuE5Q1y7/ouM9NmqtK3lDSaki6iA4e4NCbF5I9TLoYQRrmQ0V
XnWMubkh23f+/InB4vEA2pgAl/sZ/T0JTWUR96L30J/2MZ9Mr969vZKI9lr5hCdnJUNmtzibFbYO
aGbNKX2OGFj/AN4+COnjoAoJpVXp67/NLt4F3om+dK0DnSBG4yBMBdTfD8Stbvih74X0btPXomf1
kQjTLWvLfhzS+pPJvfwK+SIIJHR//Xyx3PMrEBCb+ctfQ1pKW7BX8yj092Lny2vGmfyCRUhEtvAm
uyezq3vKOebBs876IFYjAdWLgs7ncwoG7PROm1tH72nOhfUixx5DLPB4hWS7I42pmrN4xOnSB2hY
XQFHU4qjtLNeC5F3xgNvh6Wdi804iC55zJx/lT8jZfjocIbBJacyO1EAcG21uEL1wRu/7UBVUDXW
F9TBUnZtBi2QYaM5f2JSM36fiIkb40cqFKj+V/nPl4mZxTpnv6f1H2PaSwB4xyrsxxRtTnjV0t4F
3h9QDAox/RdBU9Yir2QwspUuw6pekE6yxEXb6SSigoik3t713T1VRsg8781/TewAvFDsp5sHRBfB
a8iUpShsVD4NKKdQCl8uY/K6n9i7QDU5cdu5KmNSHpnrZw67tSacmZTOcNegR8tWY9o78jEqxBYA
L6zybxL6xCe8IKNsWFUSs1YVENVuZ0uJiYUGjXSmOaNgflfbabk5UBdEQQClmpxMelgs1JIa2Yha
Y0HAI4RGHaNqWUTsLfirim0Xp8dMZJeAlGE09BgR55/mmj/Jf5e1fpcyt/wYXsRVQwLbAZlS5hFT
GMrU8SQN6fB+eY+1PKn1YMnRQTwfw8Vu5fciVESsfU0hk+V7/fqJ7CzWh0Q0PUVAp49H7uniFVJF
Cpy5AoMN2FKprTDn1iZh2qViWvxTExrkemeoK6xVU60mvb2pY2QYZSGZDUu0b2ms14UH2ey9KKcV
OuezMJYtCwsZr9w19QjuSRMAzpTOl6+0A+UfmO/JOt5A6ytkQAlK2GpWGLSTJt04bIpgabRdqdLv
Ib4xk7z7QkrDHtOK1+z+wJe+oVfVRSNVpdz/grg6Ao75jlyaNaOFSO15ikLJNxK5tJmggvoJefiZ
bS8paKSciDje5GOgHBIhbQSl4U8OrQoCRVfi/I8VATxgFjPiZKZW8UtWCZlHIntEoTC0KIKNP3bP
XZzxEVKstssPOKA0kc3un6b8IbVAIf+jO8VFwzkgizuCSnA84t2G8o87CWPb+7UF7w4p+XZycyhD
jUj2/xl+owW5Dfitzjnyxh0T87qkhxmhWixrUAOS3NBFg1XxPVlLQhL3H/I3JGzO6P4QwisebHeM
LnCO7Im/QeSxEfriz7AyYadhcR0vAmXlh3HvTnnEoZD817e1jSS6zZcWUEkHLglOWWmfQZiB5QNs
CipNSsPWlIMolo593ubvj62pi5iigP9T2M5O8B1Jrv/99eVMCMe/LQDUuJw9Asccxz69N5bI5Ty6
Og2kopUu1Qm2gOMKDp7ZLJoBeJeOrPmtocZfLpQGO13IGzmKBeJlu+NfPUoZCOPKFa7Gk0u6U0Uq
lS+lIzsBHKbRgpcFTDKiYJTnXIw1sem8AJnjzQVR9F6j9ag4oOes5qnN1ZnioNMJIEbF1UUlQwov
gEe67XSgdI998hGzv1RwPrlNzj+JI8fGLqlDsLTLG9NzfW5/nvNpfFEOf3WDqmt6RiIspxYOSRcz
f/X7Tsz+KGlAM1ZO4Uu1T1VLYrtCGm84U18TUGUTRRTfHHaJ8hAzJ18azV8zbYlqPeu+vMBYSIgV
LyryGAkvlF/Kxb5BkWZ5QNWfVE+wdQaqzTKzquaK6nQcd4uxuL7YdesuZqGpxFmlz/ne6GFNS7Rf
CEwkgwru/MXnVDWghdmOi31UCb7OreqxpG7a22BHtxauo5ATIUfFYB5e85DKSAVp+aYkkpah3rh0
HRhPE7KC94kzXyPqp8afsdV3ZQ8Yams+3V/F7/NVnKgXRN7sfHFvtZYQXsRr8fNsCUa5AC33T4dF
/aq0leHpXyjSuQDvmIUL7PX3Wnr2Y7HRup4+xE1x5O1g4HpOa8e1cXJJkFxdIMQzG0zTIEKDqCZg
SxGaCUYrGCZaefZo2bHP9xMU1BxCOgmhXmfWWo8UsMBDklFJrq+mfS9YYJX+cejywKrEgecWO+25
zZ3YDpSwvA8YSC4u9Msswq92+n+w8jRanbZLYbcie+3h45rt/sFNVmsw0kW5b9uap3E01M+Gkn9x
uAb6mJ+Nfg9ahEo+MIrUf4kN16qWx8nPVyNUyKIko3U/huhrHjDJziGU/7Lo5EgbLgEkV4fOT0s8
wcUnhdYgUGg2BgSGOW1BnGNrqHcuvC0k55SjmlEdtsgpta3pxFPU/YTg/Itd7NqxBPuO8BfjM8GT
oG4CIl+vy54BOZsDB51pjZfuOBfaxs+A3FXWryBwgZp2uKIOungrL7SDYkCnTTbPmHk0Fk0BAWaN
gWB0+skZtJ/4TEn+OUFG1M26HbhXknB1xl0Zff4skgOkuUCoUlxZlYAWnEWBpOX1yUsppytAZhmQ
MOxaJZ9Yxgxa9f3JuaU/M1R0LcJ9rehVl0D5vfcBsrRg0TKo26DhJegLf6NpN1rbA5cqB6k3VmFF
WbhwhQrUO+olqGo34PiAYMbAuVpTRtakVg6KzObKlx3hZrKgHvD54iSmHUqwUJyvAWrkmnUhpcEz
z8tRgRMwCUodeOzVFOh6mvYxW9UJZ+1g3qnVCjOrpyuJHgxw0BjuZeLIVmO5kU3s8itPkGavD/7c
Kzt8oQ+rmp1rLANIO9dgfsro3NNY3gryMDJMQDv9NX1iMy6weue7xJMzPPpiy2tMT8/jWsQwMXZB
pQS9UnljxgJZyKJeM7iMrQCF2k0KIwQ6dDYRXFnz3V1TCtc2Xjmqo68MQwC8eusLV3mfGC991yXU
ZfBx6a911UsOEzaKRSEiMGOL82pZQmeW4mAvixP7EIu3K0CTuVeu5nqQzsn+1mcEoMZR9d72E1SB
VeXiFe/J/pO7ZRK/h9kr1ZoXVe7JCrJaHKGo8HDvsS2wbpzb657zQvz7haSp244jdNWDAli+AQ8w
0WQFg4CeuBP2j3UtCJsswtlXIrFWwEdEzIUAcDIivoHGzcj6smMTJ1Qe+UsEUEDn61iE1wVp3Bts
GAWgeeLdDoHBiSs0Fv5LyDLod3mKTKVusfaMDINjmdsVC2rBoYpCs/gwYK7sjQmktd447B2i3PxY
2zNHJ2q+vmLT6xfl+0Cdq1pj0q7RuR0OZ322h+y6POsvXIh2qAnCPbFyITBsrTt9CNkeS1YETHwc
s3UeTBaxWP9QigQJC2YqMXgr/zoxJbzCaNZvD2yF/VKofJ+//zu2VhexBoYaHS9oYft0M0WvkuBa
Spd5+tIKSzxzV866GD7iHnX+y9yzvcezrycAjAkv+r1TJQ3iKC35xhJYVYZjOWR6stRhyQuU9W3H
cuwuftJP1uHjEo1WwrWUoLKqTmDtOwOw13ogwRYbV/ecHTh6ejYo/oEDzAroyyOlV3Fhs2vvqXsJ
2PeZ5rNJhtkHuLgsyQRbEeIZkKLMc4uFq2Bn0Z+sGZ/Tegaug3PRYhx0LLJ52kbmhgL7d+rylaJ2
EKBei+Jw5I0pQ369JIthkJnfwZC2vf7emrUsJZCXOXNUvUQsD0YJGByDxwfmYEqoI4njNFsoPFWw
r+su4wpKmxBUqN8sw4mh3uOXwucVGB5SfpuuMe6TsKyMonjhlXRRMta9bphnWE2HUEx8/epbDyxS
cziy2P9sh9eunTIa7ijD0gB+vNONDA3/qHh7EoZYjgGjzIhEwKuNCQNHk3xLb14qvcrlww7slS2K
5EIsrr4oreMQD02yqZQfAELq8je9sCzLy6dfy4MK5qyEeDU8LKj7fIuyt8k42GS0mvax9UwUBg1D
9IYCqS3gVVm2Z/bp/e6Uilvc4vzeHPKI4vEdYoFCY2Keh9+4zmh/Us1DBenhanIVJqzHLU0xDRFV
U9hn+LVza4yf3WY7oOyoPMHpjOSzKgRSpC+YERKeXn8FLyoLn8tZenrtP25+P/d6rEOGXFhESxC+
xpJ6pi6PTJfkMLn6UdA8+mE8uFdVSfcRCsSdpoivylqyoSc+rV+HtP03rGUcyr2N2LHeDGxHKZUZ
hoRbeZXT4ACIRxzY8XHzB8whN0zhwvM/a0XQ5MNEBfpN9oBJ/7CG/cbPelwVXNYNfLQSV5gOjHl0
HQi6KdGHHpOYRM3x1gYc8jUEkmzoD3lxrgkqUR95PKGFOQR9mBxZx4PfMKd7CyfjFviSdStS8rQy
m2G44vN2aOYg38IGhmXGY6j23ljL99BUnDz0XwTcbPBThijZk3IJNWDxkXVibDkp9WqbEwHInpns
k26xymAdFadSWqmsWf/FhXs2qXgAcC6dZLgYe0lUijCrd7AYOIfmqtLDus2vO6CkMdZoajD9pfz6
EBlko2IM3FZ5DX17gH4cf4Vq4B70xW2IF2VvwjyMUbv9AEaXLRRoY4nYuUjxXF6Q9T18OZN7QO5r
4lRmTqrPLVqtTUmRCn+8VP9IbvBvrbYLJ+awrjSb8awVLpwcJ8GyoJXjSnRrLrXoyVKjWSY858VA
1f8Vg+NNf5DK1DBEO+OMlbcaKU8cB9YJnxUSNLMsX6eBREp8B0dO0LKFjQ5SEwIqNDUCaUc1N3HU
Grfrv7e/vD0iA84j5IaG906uuA9v//OZ9ERaLX4b2R6vVasG8IlcMjrIrbXq4MRag7MJQV7UsPTL
MK+ANWD8hlomG15fK5tD4I2lfr1tTscZ+pyE91RFHEbRcDlO2hN4rtKdaeTAp8QjVbaGo9f83ktP
vrF7oDKfVWhbwgUMfPtLimKnbi7AkPj89OhMqbi9xNtVt6fuX+hpWKwcFGF+aWSimhhrfy1X7m35
iMNf3dDJ506wpmMABp5vS5hr2XoWze+X1I9ZeVjYLTtn5p4O8CizE8zx4HrFy1fl+vqYdWUxz5dS
YW7jgpFccD+9IB2yrVPYTgq25qCYp6pK8Jn6eSCHu6C7sGTPwvzYFWX/j/x/MfKAzaBb7lL/rPpV
ccGw59AbwucwNZl5AR9uKqkAlWCXFoEd+k4VjmxYOox+4k4U4xIyHH6QNNE4EWP5POJeCWZSS30w
+FtjGoWx1q9YJYl211FRZ+tgOW3xYwcKo6L80kEk+VkBNIHlMz0VhJqfb0KhqoiOaSxkNbSkXYKg
IKynzQKR8ndVD/VEElv4yBjufSJ16f26pStDeStgEIc37HVr1usSj+2nDfOAV6uUNYbOXWAf+r6n
52Spy4+1M4gmUXwHKsihlFDXD9VvkftnFFAwYAk4W7Lo08sotGjbQoAbWid2ndV9U4fOtr+MbwgC
6cCvLHgz4I8ZgBHw8U/E2IsltR1fLHz6L3UP4P8a3weIjcZqpQAJ3HDjlmrYLEghyuim1QSK/E81
PcqoW95uzZMtPlX47KG1SqNlOneCJ+Qy92W//DTxR/41QKrvDhQN1vowysPV6g73lx6SRBpefOt2
yekp+tNvXcDU/ouuBDNPCe+JdMnmaw9E4IJn4d+h3XFy8zDnWQ9yPMj68n4AlfJw27CCpHrAoU28
BHX5bko/YB0moSq1Wzk+6d6HVdxvG4DmsVI4Pk3/qA3s0QEVu1pIFtVLwZcYs8DE1THD8nHnO+v3
T5BeQkgnCcsGTC6ohLZwf/c/5yIV74WwjmL/fRW7a4VU1OTpVfMuDMBxxmpIAYWVKkviDFZseVk2
FTepoKQuyGzNyBSkG/M2b8sPRj43lOPGpv92gNFUH1e0Ah79FTVSBzNg5eADiaEXEysbLAVxdjmX
a16Oeij9Iv2Ij7UqE+ZrLzlrfiVZfiKilslpqyy+uxCqyFzOZgwZExj49LUzu0CJjEoKsqapWCrS
NRn+RPqYiBqXnKmzr6Vm2HsH4DFH5XBjV3JE8TlXbu1y8ORmbsIMMPkbQ0KNpImC4OY/qJIrk2r6
aCkSWiXeYovgxV7uYyBUabLEMjflzF9hC+DqrjGUnWK5TvYthNJQlWaBIjB17eDnMvC3emve8i/X
AgTkSa/7R7+LWGaXpoXbdr/kvNjj8WsTSPaaED+j0k3oKgXcXbkvl2LWZI7B4C18RMcfPXEjonu0
y8Q6zfBffhP2WqAmBxhGIICIJrm2eQi6FdS/aKug2BbSdd9WSTD2jXvd083R44cAOvsc0z4zaweN
y3JLVPM3w2wXsA4xSqsalCpatm8Uysy2QTDzW/7O0cKiOybb0aXAC1Q12uP9NVOMzwxb+Nn393Us
1bOIkk4DJkkapgcUh5a+ss9j4hkI+84iujRtQVIgyPA2pYaSzTOqTHMsb0ehXwZ+AJ0ScDI86vOr
vZIOYDWh8eDWfNDO72tSj7Z9EVgPN0Y81m9NSqdYhWAeUp0X4r8tpsqfs6Xpjn64LPdKBY8eVJJs
0se+khC2rFG5KyluLtyqFeo8JwA3jHasNAKDy89ivxPZQ92xFS6xrJ0xNxbfVOx6TZnXfU37jrHQ
yQIAkgzHWPjHderLNVpenfeRVQsKkArOzwGIDhrS8c86kSNg3h1qOP56UZyoRn5nczE9fzTLLDKz
9atza7sste+e8et//Mya/k5Edb5cHSCGJNIfotmc1yXFQ43tyzQB6QndR5oNiMOow2I5HgpBpZbq
JIpIQxsP1a/wtNfRADqYjSBHk/Zxf42F4D033Mup798OocAhL4omQZN8qdXYTawrkkMh5GoQP9tb
AAQ5Wc7mcHu4KGCKpCRjxn/rfO9r1r2aJ29gQXu4/6fRbAwXZtXTWjmerFSXCq/UJ/hkJOJG/v6o
AE7fHEPAVAt7ZKliHwD+w+MlvC93MsC7OcxIbr3umJmmKEpydYznf7GAR6b2+8BoyUshU4He7O8G
0q9xJiiYozcaZESIEmUd3vCaAZs0nGNzkI+YPgoIVzGRJ7aHmU5rMzbpeA3BtUJ2B3GtFc2uvSTS
jPYliZOIah8DqT9YVQ68qPpQaZOBOUzf4XnL9pNpFDdzcWosXBYBenJnjMmtqg/8E85zsUBXmaYz
/gsqHRgdY8LSWHE0w124ZC46TWth0miwYcs+DNidJRF4CJ5Kd1vrQ15Wv+9Iw1XIXhxYqjn8tKou
PBPBnlnEoyg9XpVI5Arby0vN1XE6f973C4g/YVa01tssBI1czqoVTQBQPi8JAvkjG6mBu4W7D9ST
9TKLCEBGSqFXPvti54ctXtBbjjsoaIqsL4WIOKl2+egI8j8he2kNBODzr4Cyo6DuBZi/pCxPsNf3
r7/qh8i+7H/PuVnZwPcFONs5ujvAIt4/1+n+a1KgMFyOqwodyOt5nxM1b7ePpE4Qe1dYw3DGvOGI
S/jtzoq3S9tnFocpd13o4iW1VV3FPqStzhWXUFdoVXeRjUdsiBhka3f5maFoF+YTRHbY0fwRl2k8
4Fx1YM6dT8gMWUsfyLbIg29NIxvXQ9xz6qxOuHr8f0iu+KgoRL1lRrM0EpFOSoUmG1sZU2dNgyDe
g4nNPNKDMskTQSXspo7xJjtx4U+etRkj19ZFsSa+ipiR6y2MaNNkUQ4Te8NGnDzV4DOx0euz0kTu
RhyKeGBc7UDQUQKeePzaHgpqOojjQUSajOcj6qIHt79PUaJ/QvLNM9Qs+LD6zSCmQM+mUaAfq0bQ
tL/hQZND9Q9TxlbOmGzx3MIjXJDJV9PsQmS4bPvYcHjC6NtvkUU2z/BAG9rGXZDIXVe1RQ9E2wO2
gDwVxh9HR0K1OCw4NlJH83zsAKKqAoCTK9dKVpIGG/vAy3SNrRYEmmJs2B2qprsNkv1zSMB2EsUK
uCjtVrlgMFjlHHk7pxFTUgC/iT5g1dCtjeJNzkA+9y8Kg0R1i/iCag+ADRCVLTrCbFcnFgHxOsDS
xua0tyifJ/xzbzmNSblZk2xcxSXCEh6n7c5lNS4rP/7JDFfh0qXGX6LlLdNBHtKlevWOdYUeHehK
cUqCpczEMhX0TceSaRyRryFivQMzMRpAApU/3Oq60TcAH6fuX4gzPwR7JHo9pMWzHJR+lnvAe2/D
jbrdokHklc31L6G/wfBWISicBGo0XPdbnvAGNfabk/sdzFT/5RiZidYRh+XoJ17ImocpsQRoC+Dh
wHhKXYryjgDKFD5/Vgs2ZfV3IskJmjzgj1lIy7jIuh2KECozs+RCQJQ8OR+x+YS7D0Rt5MMGFyQf
dR8x5IZxYl6ZKcA/YreI1dAAvntXtAOl2KxY26COQ/51AO/7yx//6RLdLrnEvu2BiVbBaNMX3Gmu
gqV71SRBoIxICOfHS/g52JrWnofrGF+nh3VieFb8gJrugan7U0P41jen+cmzTW3zyFZ4Sk2pJu5e
Z8b4UMt9n9bSCJQzTGZdMriLiCTdsMpscEpGqNCiEQS6tVRu881HqlmCrzg25wZqeAhUCs2Od8np
tshFBWgUJ/rJBY6fuKsr2sBS+X5P5OwO5+kTeyIBmfLhQYUay6t3ymBLw6TxARxg8zskn4Yg6vJr
REApBGEl/QgxZLgsXTlaZE8vovh5P7vf2TnPBghyV57ecHjFd4PsVFlqlwTmYYoikWWpUxcCxROe
IHoF9Yo5cE8+HFUQnUWMUOqna1MqOKoyZD1VqEprWrXL0YjoJekHclU5fYrLNt54d/JSHCeZhzJK
XZ7fPUuShtjLruJVAXhd5+nfHzHRz/EKsmPXH4qcHDxPBPbBp8s0VkeVIpdj8VwFCxQInnPmk0Ge
b3SlADqeEyQscn6muF4/M/0QOSfCLikHoOyQaIrA6C8N9irLcoZU54hXg7Cb2FJeSiSrbmGxhPcM
skkw1CTz73SU0x78gk/HzGp+rNfL8c5h7idTJ+8lTmUebagprL6tqYBv6+pvIR/wKEo8edGCJHO2
MaVmCrcAPQkkNfUMOC/yi3iQqCwJisLsOoOdCu/CcKnkMDzKHnvOf2+bfy2ASxr/2YxLvPE9OxWT
34/qEHEDoTC4RvhvDJA5KZZ+3XPSYpBPKJcEKz6rk7MzcE96jDTZlPnjnMXSWKmac0vt2MBLdAA7
W0Z65s4FuEeTGre9ci1svXm7BFKjfp2J8WX9KdzJTTXZZtohY5OTcFCs/bhv6DmZL2U5NjZ2hHmQ
jOfYjKcDNvzD0hIMdCfeLa+RjyPK3kjOVC53GX55o6XRTxf6KT/sMdlC0XfdU8pUWwVl5T662DBA
GXghcnmGJEZO03bM9lMcIZ3/AZieeMIo2AEm8KTa2SCW7F5lLRFdXNw4q1Fjy9U/ClyLA6HK8vAw
N1PHCkldxB0RGQdzqUiFdjWjbzjy3kyqNZNSPHoOtX9wn+5BxiyczvZBKsAqrm17szzzXMgFIvEh
RnCfCkWl3S7nRpcOSKSnnZ0kneyMpF39ROIYnwHVDUd6BzCrHBrO9Evqkq5svCJGOtlDv18ma2AZ
8MTjhcJMrYUZJ3GpnQbLGudKD00r++23R43lFhWGymHtnjtzd9j3yP627wyW//Pi8TKrUVoFBoiN
xq08rH6M0c2pWBZLMh849kuhiKPo8Vks+RYUld0tC9PtV6YnpnuS5t+lGPEhCrDFlC83XvJjsiC4
Z+qf+d9dabQK4d1opgKNxPMFwSrbpZ9tg8eO8fHcv2yyNhOpZrC110abyfoAUJRPWrG84NX70ZO/
+4e4DFnb4Vc0S35SVoF4tWZubid1ph6Zaq4ogzYQHW0TlPIV7TJRAY87zxZPQjSAlvdKd8NLV46G
NDsMeACvhVKVEO4+MGmLjZwzN57O+eIjkglVmp1OcCosX2S+CxLLOyNYhsYu5bprAjH43lpM0vZZ
XPcKoHSQlqB43F0+PxdZkk1YYYfD7vsB731XK6Z9jvhDw1KF97+qWq4AEbJmIRd8kyVqd3cGRqqX
i+URelFij6NPVGUJJGwoCeyrKTJk52+DBrNLm60n4tVI87t8ZEMhU5l1GnZkYkgVT6NyKip4em3/
CyKHhjeuZO6UlzmAtJklc5BsVFLCjzDek/diEtwEsBhUr6tLgw38XbGra3EGxHWp8QsMFCJDzP9W
GS0hImHTzDSB0pk8EpBlOUunUzsAGtA1fClAS4mME0S6/dQGeQsEJN6p1z423zkXcPcmrBM05AVq
L3kvqSzze29re7SAoY7YGWr/hk2xyKjYdCcNvzuNlYo5ejI9XhogFNQ1fQjkh33GHS8CKsZ9UFEU
HSs9QDF6Fqh1Oj0gwSv5hMlIbpESWuNkzC0TgO82M0C7IJYZdiptNQEEmLJbkulFrxjo296wzwYB
HJhPmqpXdTxdOLa0sxB+VMlyRFshzqzOFBmI7CPThDyHUr8xGJp/+z5ChyKtQkX8WuFeA2ALbDWx
TmOD1dXudC2hXODuDLvfac91a9XLfI4aEdwVauUCM7VlXnvLLN+NgkcZyqPL3nGcAgqRIQ9r+kd1
xLDYf2cqFRPXkg9tqCk9EWec4YkvF0B9juXn1nXzm4VoQbYCrHTs1VYwqjfwaMjHBb191pkHFLxK
no9O2WYrD9UAnYzDEMhuxaf8YFOwmUavRSHNaepWtPdVQGAcNNLuXBt4VUpJpnFGgW7utF8j1Xp2
tQEAQnMgsIBf3sUXeMtXJbLIp3LU03jSHs7t6/vt38xa71Dl3Tf5b8M5yZ9S7E0R4KwmArLCjHJp
7EFB2WD4PKKEhKyNkWlOzhvoTLYXwWOgf2laEeNsmNzST52xJ8w2xuuorygSuQKX8ICIgALCpsqJ
/sCPDXm1evTupAtWTNYOlGuyZ8Wt1uo7Z7wOYbRV9Pv8njluc5n71E6bvIpO5MLrqp97h3HAczk5
bgCdCYpV/shYFCU6ekskXeXV7Qzcc76afNnvaS0cQiMe1JYOa3iuYP0ZwlF9C21pcGAbRcsKmlRR
MqifBqIC4AnApCVtuDOeE+4I9PWianuuKFQ8kzYCH8JCFeTknap0bw4+L5CVXbqKUyw5A+DpJCBs
oIuXWY+2JpLMSAib4WLT4pg5m/CEBtWbsxcKsKh6MMJ88u1L1uhukOR1RC0Ht/mzJf/ec3bGk6fF
adQjB3hnEx8E1NDCoe1RHstcMFTOUZMb4lqPXWnHq0baGK6kkbRI3PNECLWgm9O3Js7EiOid7DVM
/pEq+/zit2bVyHDxGWk6IP9XqTVpY0OMYVO3kz+k1yAcBzZPkl5TitkJnJF++CREkORFIdhMm1gh
ME+tdFpMRFUHzPdTiGEEbjKDUOvxIWd/1OOVK/8L+qchPf/DXfabPrLLF78yWtU8uO5uilIEpLHT
/d4zxUhMVt7qUE81rEguP5zursOB9EeHIFBwaKWOP0bRSfr1M7vln0q3nN5mJ2l9dFsVNr39TiYL
mAG5N+y9udS/OSwdSZlVMyjG1lUkHHCYz//2LeRVyZdMyoKThFTcTiJA45n9UVAaRSrsgfpJPqIV
FTPmKTnjEWwjajKj05W7qDtMmtLOmCr13Srnivd6JiSuOsvhF9/kSwhJGbQDtwIWjVJaOy6cKXh1
Hy5pNWVlelNTnDL43B+yGtMzZanRBMbm1UjxVihwRLh3yEr5F9YIi9mUqQ6+zBbPrz1ujmr5joTw
xZMmFqb7MFxiXfY/kyggHDgmHPeqlUEKuxQ8fAQoRw+YHnK1f0nO0MH98B224p0iOZO/koGaD5vH
pcmkGzdITtdzsItxST37eangmU8Yts2UV8BzOZPBuY2aGwmig30r9j/Bm7AAXWVHqs128iNVRT4u
CIL6ETB9xFAG7QLd2Aqmje3wKkI7jjwIErB+Sdtr/id4fzKmm1z6q9TEkY/Nhg15MvveUFiCOv0t
Ar9Ps+lu2oJ9kLBlE4gayMbTj+moA1WfFNO7i55xOwnr3LY36W8MTLzZdo4geDnz7h6RO6xhSdIS
iw6Umpbo0JBpyVtl+1ERZQ7nGYIJqIIijyVQUKlWZWdfN9C8yNQbO/DE8RkyvMntySWHcENNjjeI
GUEQr6n4ldPeOzua6cb+cvKcAADcbdMzBXUxid1r+JiqAnaUG0Q6qpPifRUataaLBLdrdwZUS+Ve
UDOo2Ef3hPUjPSsCUQ2kciPPWRQYGsyNEjba6BzSasZeK7GyLBygDHMduZ8iSbOj9lVoPle+nech
5bUo9nGp0y7awSiU1+5zYDu8VdHqfmDdnhP1CeYaM4xNVOKRlJOSK8JSQD61XwLIXYkS5G33OGfR
5VDBtb0FtJA9lE96p2nnEYkmJ3egiaE4MMXkDzsHy6hyUpNV6ux2qqdxpNY8ExRIG1p/XdsVddmw
Y5AgsdrxlfihKPFwOn43d3Nhh87F3gt4sAB783Xv7hk6KqsPEpvNG2iEkpdLwGKV9Gjf+8iK1DHG
XyEDJYSVj3kTWYXWHJ+TqpcQF+sAcC8gAxo6AC2tdDUd5ZXoYJ6/ehfxcu9bcsfDQoSL7RzBOlMt
OpNj2OCLT2xCZd/69Nfgpa2SnBuNh6KurN9vOXI2wwkmZ5cXpEt+vbDVcc97Md7sswnPkKsbHlNc
DERf1cTuYR6WWvVjgvy+GSQfO3g71kPXe0HcZ4KVd8RvW//WoMmKdQSflm0qTBfnN/40VR3jcIkV
wHaY2nOi770gwnncwQC5k+sxTTDzW767rpD73n7cVPT4z9TwciOHruzB7pEvopN1kJbIaLTzodDF
hPWEaVo4hFULuMGfvv0iFsz84fKnWYbwAJEIiEaF7xtn1mdTkdJ0EQPPTm5zevM/1PHL4Ucc6QOr
hR4vHn3fAAtTZ8QnrSGwlbVNL23gHDqkNzZ7qLPeztS/mO6rjbFinT8pkvN+NMT3FviKBc2zw86O
jeaHrleZ+fx8arZZtaRBR4O0GoTmiqSYws1wanGw6UKgudle6Z9GNmd0oVuJ+Y9yyXiGa2ZWd+ai
Y0Xfk6qLPkukqWB9FzHGnurMXyczAr/KjDu5mOSYpZMvQQ2HTQjZOaXoXqdDbK/ay9l+IRd87a92
4qZCYFZbm8MjTjDllea9OkMNhCR/0XjqdevbTJqpnx4VfVREXolUmq13WwenvuroxsHpIKfmoGG8
JUgJvjVw63qvXB3i1TthLr1fWkkfu4V7QiczF57q/ax+9SYn1wD6PNolcy6CLBwfkJzfF8kNwc8Q
/6BVZTLHyoMtM1h13ddNqU/vDu+1tRtZTkd+V3dPOYgH6V0o+VendoSkJvN19sMyIaTXmQ89Q0IO
AsKLLyAqR2VmxLm5elWy3/Q0FNb6EMDvS240euGUbmGB5937gW+6aMHapd12luYhGlrwBVAxCjrK
p9g1CyponJoSpupClCr8LCeJn5Go9DzzSV2vnXWJq4WvVT0g3jqgoK8NpaZBhTuOqEpw2m9blEmH
NZvu3ntYvzQxZ1AlS+OM1DaxpcP6ZElu54yvjz9iKXoVatiOwhp+N0y6Wo0X2klHCicK8zxy5o6z
q2YxbrPdHvBeFiSSR2Wqf67LTgwevinxd0hRhPR3wqJnz3+zTrMLIVelhxiKhJsJdnwvN3/eao07
FewGaXR1vSMxWzbQSZrrrtr6VWvOTfY3V40YKxvV7a8/z8SjAjqiVRZhE4YvDQD7TIa5YLBuox1P
F0SmZ7a0TMwyfT4YUhZ90CoqTTxJKG3PaU9ZTUi2kMriXGc33yIs6Q+3O2yaQNq2ggT7Oj6ruvIg
X0RtQdk0YFk0TRb8fIh15FWNCcLM/fna0ygOrOOQWmZtpWOZNoyb9YSWIPvy2rW8rB+zFbBreNV8
sxjEtRVab1JVHsHYvdniz7HrOiNzo4yDQnJKktzrWTPJF+Fu24hHRN2D8bbLaol1ud0h1ukDA548
LTEQsABz1HvTyR0Pl+EBc+UH54VRNDy2tqjGFKceaIysGFZXodQAvjOdeuahwbGoosDRWJcMwPXR
Sf4gI7F/6MChFb6BBI8Lj5q0clahd5N3ZLOlcZUeT3kIUpYkADDRvzDKfdwD2FMYDcu/fxyBgLv8
mWBs6hzBH8oJCPMPcBbt0EH3x2Z/W574mCPBBia1EcH25oXZ3ZNv5ffxpM4c5l1W1rtC9olwFWEH
hb6cuokeQUhlfNtldhdeH1KTu0GSp8DYiGR1Jvqv10a0d/rgAAs1ooIRz2xSix+vLgHO1kwRC8e+
tlJpphRs8o2iMKRpypX07ffdHp2Yc9Z3fe1ZbQoeuyB48AlhYZM3bxOG4hhpuaF89On1g7ky70jg
D7zf2pcPRcl9dsjwMZwvjT9D0bJeA4IU+IRSDlBMZ0nykhvzpDmf0o1LNcEqmxnupTAiBHN/DEVv
Whja39UCpOf96NowXDZJc3xIeVPchXCQq5LlFc8MMAuoEvJtr+Qm95jL1Li2R1uImM2PJcJ4Z8HI
c5CRa/2Dg+WZ38LLrGPoijUTmW65YQZm3zMrrNlRktbs/mGgCgR4PhyHl2wSxtM2xC09klnFqxYl
EL5Q8I/gaCs6Qj1Xw3Fx/japCIu+v+KyEgneD+001sizLCsifqHg7z3JEwW8b8oSFvMOk29Vx7HK
aasLg4BwnZ+iBDom30sbDg8sR28mDeRu2qUdTaL6L7JyZcDVE9jT9T9gl0VZtJ4gYG0lOgSAPRsE
a4gvfgd6zZ+cziMZE/0uH4W7c/JD/WMwlPD+8bIxxx8E+/iDlk6Mko1tk3IHeNxMDqJIauvZA44N
935HUW6oxvmV3zgs0KZ/MLTk8mrQekyPP3UJ4mr9zl03fyJlCz9upRp5LPBI68T8TTvW7uEKIQTQ
YYt91KkszsemkGl8nhM0IbGras1LF+VAW9M6P6tv6vSrEv9MCkOYbHqVmrWTpa8WRfL3eRsC/cjz
t8RxmC4aRRE4fHqsPDc8pfR0Y3m+/gYCdDCJp1MNFcDS5shAaqhxjbsb8fKgpB6QqbXpxKnmaZj/
mACooOYKlZFi4cBk9dF/nTYMQk8kbPcffibbYZMJHzA2nIirFhTFtV1jzEyX5HsKHtn+K/ApRSeK
IFkHEPtlLGZdoIW4kGh7in92kjgWZ1OhLJpaRi6Zd7U42mwo2kjnIAyLZtePPVOAMSpg7GJMjgJz
KpBTun2XbLgx0QuJ/lxB+8r5N6+y0w4BC0urh9LGqmtmmBSPW3E+yNiZKPeGZBoi0Io7zAMdx6zJ
StRm+n5hu3y60PoauBnBF8etaOuP3WnukhCVfOJqIhnuKMmRWtHw7ye/WWiwHhmBDp6pmgmb23mC
M8lNLOgyiVbTw71fcCzyHMpKL29nb7AgA4XPNAP3NmuOW+uEoMwnOVc0nh/JjaxJt0zSpKTftKYk
LAgbdynFRbMcMtUsvhzQJUwVas4tu5bTVuQZPuCDNEmLcYtULu6+exoC+tGrnBgWV6kCUo3AdjOR
lRoG3tkvCC864hKk3orK3tH8DWXslYuey2eu3/Q43lkNNzxdml+K/RdKKrFQIf7AJltkmsRVlcgO
J5c5iiuK6zhCO/bXbyC+h0ukAzuLCGgsifCKjzyBJcNDiUFge0YcZPp4RR7rQahqHMMqpHcV5DUK
dGTZXFknfa8yn8+N6x5Sy2tOWHObmg3a1hNXD+VPEj7AzM0I4qtfW4RtTSsDZAPrdYuCm2tTPvVn
GYw7pq9DCKwNXMo2sTZiZ2jbkO4rfwkRPW5/v6HAhSiyVuvqPLJUFImrbv1TOeA0P7ZAjhJkT1VF
mlaK2gVqeJg3Z4RfRbHuc55bmNk+EjXwR3C3Y7WTHbR4b9oFNPdVRKuVpSH37jAuHHn2DQTdEgi5
AFixtANnGM3Q1je+B1qm4Grmo9cQ9yyfdgyG2M+oSpxf0pwVKU+ylNsnFD6rJ9npfavbUHb3c4W4
dmLaMtk2oBHiNpMeUdjxQpc4FPTIHPNZB2gHb0krNN0tsHi+wyrfVNUvgeSRMpwyE+e1V9SsX7L3
L17Ho50ph9CwKMzgl6vM7abUL4leKquKgl7uLX7UbZQ+Kw+/FHkRjZ1cR16D10R9eh+9pvtd1qHT
X4gktSrjhzPrIJo06M+4DadtyyFYbDqtjt3HEba7UXIAd6BYd14m4X4zK7m9KJfVBlZOgvTWSBuS
62lPyt+K9oNY+wfTi1YsDlEVwUgB+2fJBXqBpxanfcVsjy3kyTHBwmEg+mNJhRrN+CQj+WPQCVAB
uCCG4qs/XnLDyRIu76y9tDLOEeH7HNNbDAxv6X4uINkOqRuPxMTHWbC0cln7AJPVSbXJyG5GvuSa
Dez3wyP2BfzNwnWk7C3m+nNTrCVHt0gHmYLZjyE37AL6DoiZgMf4s4zFJN/V1N4MMxKtPaeEIJaP
bVowyE4v2f2+QRPKwamK5VpilZslxgwzytR5UTAhfXhrwkUp6K/PZcMMOT5vlLSjzJMzUH06cdUW
+QvkFEnt1UcOADO+kCMxEemrki6A8x2U+ncgvbZP4kk19KP6nDpqnTWQlOqTQ7+4QfJyWtgsJ5ap
kJSqmEH/I2wnV55B4DlUlmbCW6HmxmlTz6p9LIJzeSIZRhGsUSYwuEHaPXWyrbEPCr5i9lnFeCjv
n4iZ5Rik/E305qdpAunUrCLg174XvWFjM6sr/H0vNGo17xomOZdgxDLjCJrrsWzTv3CH+l0x6T1b
G1L2jPqQ+R3mm/0cHc3JYWqrucj485vuIgIz0IrvJRtvSeQPSKNV38je44+/48wSuG6wFUNplClF
+GUr0rpLy/H2nYax+fxl+MQNGg/5o3vO/rw5tO0nwzVQMpdQct8jtKIGf5zFRVe4XugTl2b2SMo/
ZKUmjqubpuylvvMaKZl/AO27GwbeBkZvv0B2yw/v83z4uq+NtouTiJnAgIIdxlvdXnW6UeQRxqvO
EDchgMqgmMOfekKS8LE1bRGVOhuBV1H14t9QvY8r8QY4sk6q+tnYoW8eO111etJNOfYHs8RrVzTy
OLd6IsNk59ekylS05yNPgWLmCH1MSSPL1w8Sag4f6wwY5ywPx2Itd6aLqj3/DcelxeF5b2TRT50M
k5EfJd5IhMOPDMiakrJyhH1ewXly/Z5WIvg8VovAWRNySmDJ4vqqWyP04L3mS/5+IMbUP3+/sX2D
OuwGAKz9aL4n8OUqcgna1SN2Sx6s7vdporkOuK9nSkzk7UomYf46inCLButtabDAG1fKzkCObJek
q3XZDPedOPXQXb1L4GDRM5ePyxD6mhT41t63RwHcLgkt0y5cRaENloufVejtzvkvcZ3ucI95BMGt
IYdJMGQEzlbxUceGArx0gMRjE8gF90GXfaeJiAF+iSXUKKv793mzjWUuNZiLTCpr+2q3r7T01pCT
7xOgJ+wK+mxZLP2efwZC1Z68US0DEmVDkmnwUgx2o5zAq4/YvS79ZCz8cwBUJhnBQ2mdmbpIaZ1+
wT6ETwUXpNqDLhyrHXjtg5TO3PKHpXpOKfIrw7+n7FlCFr2XimiiqzRxu3pcepsOlTdjMxt0hZoH
lO1cNHaw77VpvLTklrL7P8wo0ZhjKO0EeUx52/ni8Oc9JHMq0UtrPpqIjf5LbR/sD/HQZDOTNcTk
gQgRyZobeDptVdqvxRxbORBi+Zn867fkxJSiZxMioB6BFjcjQVzSLdTz/bcLMY8vGcr5IcCnoN6Q
u7jRRtPRhPp0SHo1+xn57U3GnnUnv4qpruHlyqmxFIoE0Y1A2HAdvLkSr2jxEoD1fT/++HYgnLTU
aMhxN5DX9lavv4Q+/rHugrP9weQVG6x+1e1V1KW+KXdz517tagku56IR02f5NDYC8WyqCVKehSlR
4OayYH6HieXgVq7ckYQiKtXzHhB9YyXE+XjIbDIS6E4OcgEHZXupU9ihGdkKTxioBbKAxfd2Ur64
H07dUGHjdOkfPZ3TOx59ZbAhP+xx3Red9C1qLqenk/4qJsGw4YAOIhecNYxoyr6SJBYhmD0Qhee+
+7k5FiiieyEOg8jCtbR474SmXrv+/W6RIsbuWDDOyqf4PpKMi0wj12dhPTnXuYBEPsXQ8no9kQHx
7RhlHUCHWL89CbEUDgUMrfGR0GnxfgOL+aotxP9nFWVSzpqqvbqjlxct2x4CDpDtUlZe4zVX4W76
VDpDT/V3kKMGEI91Hed4y+NTXZfCLdu6gSb2buVzJfnOG3vEhZEACm9LKAC791PculZEgsjFWaDu
4CPZZgLMGyuzBS3OIhbkRUaPIzhOzrY+daBkKsZwusLLB9dbiIMnDQede7HQvx2AHUaQPjvMU7m0
yRX6Pyj+RzhabTFUCZyQs+3bPLnFiFT8/4CBOFLSwKMw+0efnoaZuUQrI5mCasyBKtz36h1VuOL2
Rg8vSp9sOF6pIo+x9ABNsdV70hrDQAflIBSs2uVfqMb0/WuhrUOWgQv6+QJCVpUAz8/Gz2NpwuOm
4aOKZP2AXkIKgZcE21Ds9WNUhjTO+Gu1f5FR8J6jxfbkn0XGuh/l8nz2B5PEQd7WN1V0gvtd7Har
OfWAaP7dlmMrjtkErpCD20YR+G7nouoS0Ommx1hHDE7kow1FvmbrcFVmHZ1Qitx0tkiALGZpHX/U
JwLjB6PDSyvoPJXHF5L0cJPgjd2HIBnjTkJQHDA8FraUDqhxs9XQq6q80yp3JQPM2oZvEN/FRmNt
1MW4YKq1VWkLVpyYV4DVaNoUw10PSJe3MljQJYbVL8LB1sWZq+h9rr7mkWpM2lKGi4XkYtNodDBM
yBb3dShblOfEOXBGmlXXMyc3v0ASYoKoGH9w2cxV8d53sDsOCvh9gxxijGjxKXDYmXWjShuPEjrf
vKj2Ey7lzenHn4NfKm8Yux9H+Fwv8iWtX8r7fqd8lEIqxXAH/Kqp3Xb5cpwC3bPTyCuXBV80o09q
k8GvUWWqro6rTYH5OerZEb7uJCBW+zzY6DVbDdLXer1pj+mt41yjppwQsdWtET987equewqgM3yo
V57WCakgyhvNphfMi+uQo2HZ6lZ5favuFer674J4vcMck0Du6rd0tTcpZHY2wCcpwW8T30VFl2SU
dA5mQA0yspq4L5tjbmSX37Js0AcUqtyLhVa7MBvM7evnshrFbXH+tNROvxH9DcFDGV/Lcf3sxg+D
aZ3QkhDyk+QtLYoxrhj6/bZ3lVv4U9l3Dmka/j86A0ql658e6PsesUV3tJLjgkOmJf+lpTNZEb6r
IZym3+wNqR7DHTwsw7D9QmBxgxqVCvsMFbcu7NxWVsn/LR5Rhtz5gX44lgQLxuZrqHI90BwGdYe9
y7O4Nbozj3CKJWm+cWCs63pKAPsDfI2J+y/9xnKtvzRbpIcPcrGbzThmJWy76Cd/d4YWbnfufoI6
zhp1PxiMHIqzLF+k6Hmd0Ht/nWVQIHF3Xxa9w9LTGWpxdD1HbMMZdzYPnwax2TfqjbHTtmMpnqW+
muGOthTwARARoBT/cJp+wgX/LPikUz0Vc5w+Lt6Yqcvdr3ZMZhbosyY5fWBUxK4CcO86obwJ2rTy
/koDwPe6VVObXoB/ro8/zzWGT2hWloRQzTWkleV5eUgJ4MlN3MGqrhi6haBQ0hcMHsNYPK0hjrtF
iYx8QVPW78yvwm63GsGeuRnuMX6Lk5pibRdkHR8e/NYkzUY3V6wTR/W771UMPM/8RH4L78YSN7gK
Ty97k0As2W+MH6dxfYK6FWfg4DL1RrtGZFjrpdLLrjMCFxle7HSSBzRX/bmySui1pikDA6/xmct/
2D2ThGBQdymDLAljAU+oSnRleB/DEdufbmkC0M6ef93OmPGEd8uyeNaxAvgoo8Rt4eyoTAcvp3Hz
c6164ZlWm+k3WHU6ZWitTW0FtFWq+9xBYWTD2pUn/ggT6E8hme/yhNBaHMnCyeeg7z8xcWfqFK0z
jseoInsrqBppEcDqJhDSewyDwlzZmY6YrKjeFCK9M9UEMLIz+KhNTBwl28zGT6DLiLsBupUCgvER
MTfz3bOQKWG2hq4VKs9Wb9OrbKaOMreDNyqHTOvz8UDXh+QDej+5XKq//TjXAb2s/PFDGfcuQ4yu
Xyr/D2XtUbEzUFzm/R8Q1lihdSY1OhZVI8uL0rZoewy8f6AsYiXz/yskQt192lkdl+C+4hCSxXlq
cfwHpu1y3U9fKyY+ushS00wAUHvLP59WEsjgg7xTIkBbsBinCepXOgmmkD+TX8jGIbtKEGDghc+J
PGf7v2ZWoTG9vZ+vPfuoD76jBcGz7MN58mrbSSVocb4eCQXcHsyEGO1RSgSPfiILqIuxwwhZz+dk
N9bn6lZoef1NgWOpbvOxhjRvx7t0VX5LG8RP2A2ooUsXLuWVIH2Se5KBm6lXH7zJbdUh0svOR6gK
Figg2VLwmuUAa/JPkPxaK61kvI0Htn5tSJ40BZ6VqNB3lulObdwAi7n/iV5Yaywml4zJMns5yBPE
VpCqhotPGlxsdrqv6L59APMyqICvowvFMrFhlueMVf79ayffhyhsMCrJQbWkc3J4O9+oTsNoQhU8
GBZSPvgko/7l01CNN7v7xeF7XcfwRmWGqY9jRtoIhJ/0HCqplKyoRu9j96VkzZSyHH55s/w/ueaG
Pnb833TxfoaQw9D9z9PisJcuxf+XpQIfnLlQoLOGHgNUK0//LZlzK51KMqvtEr7FnggYvo67w2DO
6wfiz659gIFiTxGvkGS+XPA+2Sa23IMm32/QI8OqoNAPnw2iWSd+Fu5vqMyXR1V0oKKH9c746lDs
IJFY4El5euI142MMm3Sx48J2p68IGWPuT8TEVEq8hdtIaf/mS6MEiau0mFECtw10UcSvsKpm6CwH
4RHJSwgP0M3URuGXjcDW5MdM0hsQsTHG/Tq9X/KPz+UMH7UjnfS8ti4BcRYKE0VxNa1f+xBH3HDE
MnPmOMTGTdeZjmYkd1j/JC9mISmE8V/WlOOK2lams03JaIZGGHgyPgfMzhSwQWHqcgT0KN7ltR5K
xShVslD5mDYEbemHAHH6FDgWFI/BQlEpM0Hd+hqdZSU21l4eLscAM/ow78lN4VYMF4UNq+p8sarW
uceTQ7lLGhQ+aO15RT7CSPjxO6/EbOuywCgaS/C40S4CuNFD+864RpCHp4sKbpDm0yEMogZGrX0O
dlfPcvH25VQBOq25fzHOeayZ+50OKjlAHejbwZjPBH2t7c30HQL01HY1yTafs47ZHzkaAedEeNw2
O0dzbeeS1AF1AF4Apih+wrLmrdO51jv8QefOmtTY3lo6Jkd2FGdvl9aFjm32Vzr+chfuMAY66Gr2
6PDbxwGIScHuiP9IU/TreZuvIwVA8y4TyCYhVDwJQSOe1FAcHpQ8BnuN4Fr9c5h9lachDyE/0ZjV
+vQPey97lBZcHu0PApNZh+ipD+eJpP/exjYqdcbNqlAouw2mqA4HdeWwUsdlDRwuplJvwiVi+oig
jRzIvyjavmSuX52xtT3m4G+8jNLbYbEcojggJR84LSRMvCjrnfdU0Ysz4vn93ISrApFPOF9Ibsbi
n1iGqX9tHbRIDuXjJNejbSkVatX505r9dnuHWu4l4vEylthRDEzQdLo/36kt3Wz10E+j+wdZ9oks
5m6LABAf9jOisL4VKSkqcgv3E30Y5ND3WFPHNUpQtOTLuF/3Pu1pJQpZuc0cCPsfkNG66cKZUaG6
e6Hc72Mgi+10LflhO1Q75OPkjzQvwI9Ep1WWR8Qpg+rt2XWTiZ/9pAEVRHqPz8JcLiBJLTuaX5wC
ip8QoajdoMjvnwIQxi2nNZ2bR4VUU+iQGVxvspUgatju9by9oSudFBQNJikN33X17uGRNI4/ykQL
g00m5rw2nLENrGlAFf+9CdnlVtgNxQ4E96xdH1lLuOldGoh7k7qncY1MVof0hiquIWKMbzJmiMXD
kbf/FhLA+DUQeZTb2MkybIWi4FoLRtH/eri+p08LavdXKXMbLmZodBoBvFgFlozNuMRT+DeZEv48
umfDrxyt2S5YOGA11eoGnLMMPiOWDA9DDm30O368ZnTypNVwqspWBSl4ZwLgeitY29k2ZuzqHXZw
BsRKzshmDZVxjfMoJmtHkRkEfQuLoSklkGCahKLDFSWUwz/fsagiq97e2bAN0OMbvj8EaRFb5MUW
6g3ymYiLuN7/UTDOxFJEYHbJ8idkDixfXJFy5/i2lipqOzg/kQDt3GMzAhD4RwO0lVc/kwQgJSK1
nxwK6mAokxHrxCGUFsBhfQM25GjDC46rpcm6DQnP/PKc917qbcpbSknDEh1dZO0nAwlL2Ih2/3bn
LI38neN6Ovc9/tjYJBvW6cAVABtqBFzMZao7xLVHtGrbaKkEfIBZvz7Hf7XOavhM8bgfm6tplSa9
VCC6VO0K84ilXkb2KD/IaVcyifeq3lqc/6msAjOXeTwkznA/qEpIZDhqw+9sf+4dEXkuWQOz9Qg5
I5IVCEsp5MFgT8zmPwxmo8U1F8Egl1lUfCn5h22vplXYWKddR2ZmKffOi3a58dS8ubbsKFuo7eSx
6/+nGb9OuzOz4D5tnO0ljq9AVCLnLDzyoGkdRAkM2gvxs3OcTGfs9/VVAdxy/COoW78R+N3A+DA1
nVQPSLYnlA29PvPUzbQVBQUhvA30435JmRqsUfn1jybeqJEjvASmlg5tkrH3wsfNXoUTQejFTj4N
kMujxsdmb13G842mTqp8hmtGw/XDlCiaPOevPkNcwqPZ+J+56sRk1Jrul8babUevWLc6K7MMav5W
5U5PP5gX9wKdevlN8ogNXs9I5Ha2PXMJY3pUeCIclkS8NqIyoHf+p+kJSbbtR0ooV24FKkiVzWQP
e3b13PArZsbGV5zkSPhv8C2ojf7lH6XR57hKU2EzokNSG7iE3UGeiRnCenXn18z1L+c8/QmMJznU
gFdCRUew0AGV5g27UTT1BeJC2pmLoqBxaXN2AoZJc5M96WRcqvoi+VsLTy2xHpbQA/iVt9AbiUFO
9m1DVbbZ9S8uU4CINWNLAE3lnXdCUUEy/b37w3n3CKnXvZOuQP6pe6rmfPDlKf0qgeQcSX7F6aQB
Kj1ahgqF4UmASynptR777hmbMlTKYenySz6Ns0Zxb03U3c9QpyhEMGRzkXPSrDeuZwRiLrNHu0W3
5TA9dCjazQO+OWWQnotzpF8JLDM+baRPmDIofpyt1T/fbz3VScQIfzh3uNymrSoFrn9VU4sCFtw6
bv0JvP78YrM3bBFdQtVasWuaVYG48529BFszhpOU0GYZeP9FpZu84pLn5Dr3EuoDELixTaxeCATS
9Xo5KQ3So3wWzf+UNV0d8q2jnuEHu8K7bQvzz2h7gl6HZv2TVpA41fMZoA4UkQlj17v70X6TjtTe
fu6EmCP3EUT/mTZl0nD79ILPMYuZQwxm2MPZyZxds/2zha2oKJaub2OEy56dyonzZgNOPqnzO40O
/hdJ8oNaGuu/RFI+rEcK6E7wTz8U7ASbfYC7dYQM6Ol4lNkNMthT8gOEv/ssqDBu7JBLvFYr/Bho
DxDFK9DdN/CK+VUrg+apFAJ3O3evB0WwstysEXmqudqrQtNCbMp1/PlDFb3/sdCUhx+fWvJ4iv21
TfJi+3hGXlsjw1r0/IlT74USxdsRdJmJ7YzS3pmdvy4csWVenqFnw3X0pVQ9z/vg63MGx6ekZAOg
Ch3hfzlG/vCGgnf0LXAcp1ZLRl8V+5UxERW8AZb/Iz+fAe7sOlM2rWqVP1kX0lbta+l8ewLwZIHr
AKU2krHzvfIxBAh7J1SzygVIe38plvz0MGtcvkzTFaQQq8u/USmSZI2myQh251MTmBxIsRVLcALI
DerrB8anlY22pq3XReLnXqFneMIimjGtbbAfYFelx4oe8p04iKCA1NPPkEFO+ku8keaeX3BDvjab
ru6Z4RC5CAGkwDGLRg3TdF7ZgtIeYQRWWR7uGJCvZRl7OJJF9UoAPKTHcY+YN/1RVqE+tFpm8mU0
QA+7MNfatnmA7htpncDSmjwbL9YoZodhxpwr8LqJGYoIAJpiIqRBEoGDu/eTGTYAQ5tMF8GxhuO8
+IIRchY37wmLJssICDvTnaml/hKktfziZOwjKgF6gOElYP/w1gRtfWcSsBRVWfoUTJf/lzPA10G2
tKA3fEQdX8ZOtDroAXjVulIrEvtk6W/8j+CY6bljGTnkI0xTDcuMqHdllgtMIiTFg4W1GPfRSdtx
nDQjEtYgOPsAgpIdra9DOni9UWYcR+LMpofKLFrVKlTEhw+wgFU6cIuCCPEIbgnC5rjTmSeoJns0
uBq2jLhc8nqcb78h5aUmeOcdH+B3i1xJA8ovEV/GgI9756SOJl4w0rXMIUfblIaJjP4FpBkYZoRX
IaJeE9fWLrcXad0XdnWNMjeG+dOJMZwI0xIDRjwT1MHzF2M7tKh396kt+mgCexdCjKfu65Fl7cNg
mwrvVUefTzjB5NuqfXNGGxtdlzf5Lkf4N1cdALo7WXg4G97gst+jENZMGuk5CDJZGlK9YAN/0nt6
rHp0FJ9r/yUwbcYXBMREozDp0/BoHOJ03UADo0vS69dIa9jiqrfPZUIw247Sqj1XbubVTplRDr0G
QkI5I1X7jssI2qlPxtMTEY82J+2/yE7GsKWWx38156BJDKE5ogb+51eTds40DffLT4wNYDhD9Acp
geJ25F4eaYyTsz7OB5mPAQe8zoWiayrrCHeJtn4CXBj47I4YdfGnoXBWzsoEOBpSTkk8ayQIq3go
9Ov2Qi+14i+fx8qiXQnT89wN19jaQA4Y0xvdeVuyaY7K3rOtNahMi632poJx/2cKFJRWNomu5wrY
UqL/7vfTQq8KdzSS4PS00arInkPV/bMAWdWD44fSCZhrwze58pXRygl1QM/AmQ9JUUSorgzSIYGq
zW1uDPbEZ59/wVdNXa2QMdTfQ7UO4Jhp/x3z1DzR9SxbOQdzmI4O9KVkKbiAauFXZVfE4F2GdDEF
Xlml9TC2N4H96qPy67n8k1zZaUBoGSsi1NEKCkb7YmhB2uHzxu7rFjIPKiOuN+cJcdli0dSIosFu
e6VnhFj2znh2H0KlVEjRanFAFZV2JAcspwc6yFf2oIjuvg3omVL18DXwcNMgyP1aSwiy3Ys9h24v
X6VXFzNKSKHD5jDxDvIZ490v5VTLvwM3fIksMVA8OIelbHYQFJopnYThuQfW4pKRP/eX4MR6XasK
hSLgEvIMXVP4FPSNSjGtoovS83vzmHPXSfLuYMprrUUb/cmroY5+W3WIJKey3s8QUx6on/+9pb+y
Cf80RZs+qpFWYJm0RQ86Jx2upQ1isqJ1G31Uyk0H90U6D8dSDcxO4uSWcIkGufKUsaKSjoWVkdZ9
s9jBYgELbM+XSFQ3OjoYAlit7pFX4zBROU+YJ1u2TKQ8Ml8GL+zNReewM9rYNtEnC1T/gWqGpYO9
NHhNldQ5s+E30TR4OIJzmfbMadj+Ndkug18WVqZ0sK36WRMC1TA9F2swUr49+qrdmR5ctfoQjd0N
AfYJr+ZOupRE//TphbSKAxodz+cjKQc7EjqD7k+xqPnOhiJRI4K5R7udJRBYv07q7O+n8NfRzemT
//Url8dYeWK677txWY3xNlf5u79UJjmSOmLO9R5fM9UmKRjoXYtrGgPPrtFJx4667TsqnE0LOGBq
wploSoHOnwC8xu6MXypEmHp3hxDNfP6xtEHILd4tpmyWn2w/iE2BCzIn2UqhhInqCAWurLIGdhdk
36rPqX4zSS4DqJxrVPJpJxFEiFVVLDSQSim04rbE1ILOzJgdHS9cDkxGNMJlS2JzWTNcJUh7zJ2h
jhnqjanVtZnVoAoQKAr9fTDKmbMeN/hDxZTeZu3BQXRZugpyzpRnfP4RQvlFJwnaYED+XpvNcEiv
wYYQx21mdFKnmjw3U9hzIpo+8GUVyObgUZ+YW8VO0eX7fcQaQc9ReFGLplgXA91fl8eCCTBWc1Nx
e288cQgaVzbAz+SFSPIjpWog5OJ0iD9ghnTiA7JD5V6uirNgOeVuyP4WNZ1oLtqssbyXxbwWB5+E
iD6/PyCM4Yr1Iu2Crv3Rew7ROOstrmNfCpCxz3DJcTnFmnjPvy5R+CrECnktLNWvf3s+Sxp9rUBf
YL/c+Nxzn7cH52lmjS2x4nHXZcR+CFpRnTbD3SvU/YIAr4/7c5hCV6ehzGNKnMMOfbkkd69ICrKm
iEaEzZnlfEDo9LlnsN9aYlQvDfgVEUsrJX8qbFlYmOFPgCJ2knjV3LrWlITTdGvKrvZRApUOJfYO
+RVgciMRXJmm7HW3lMzy+7k4PBzy8/oU3y47qhhM9UvX/2zlweE0Uoy7hNDECCQ+91gRVah7YVKK
l7MhVwVFBiT5nMAeXUHTTjVV5ZRrBrcu4mt3X7XXaz3aULaKD8/nOaDwfB4BpfKmzozEyq5+b/bY
4PCLmlskt2efUTe3z903AmhJGTyYJaS1KgQhwgsrOL8zZ8yQ6h/f5vpDQaULcIUn422QEs6xKtXq
UqftGvMmttyw5zUkeLA1E3JPnctUIGzaMmfMWkMPgdMyrvh41tuWLXnG8UosA0dpF6LXhbAQ+mEU
iymyPu1fYWMlc/PtvUsUd9V52I2tEJWu5YLDU1DQj6ZQW/a3FnuGETAhITfUI5707wVGnx0orHmN
3maMC+1nrS854e8poDm06uk7svn0dVpRAnN2WCnOnpqgxwW8B/xFGY1/62Z9xE2X3DItm1HRwNxr
ls/ZVVdsuqU9+1JcrqXHyeahSkV3+YzPHxqkiEa7gAklpIyl/fxHve5D7HdeufATTVG2VYSaJRjT
pZ5PLzIiU+vwZTKtApCy9e5NxW4cWjni8wM3jysXBoENicgRRkj68OXaxd8WJpOQArnf6ALhfjg/
vsW/2rV8FK4EAlSkMg2uDRTdzQFG0ljqX5fUrIfiVOMn2clFXdRgcaMsNbP5oEmWzuqyUOTMi0JU
Q5ZhUrGIqrVzYLh5acwKaRWu5wQXla/YmANwwD84lkn46flQ9wzbLI+psmI2S9aOvF/mLanBjZZ5
sx4iO0DbCNh8+OmIN482p8mwptkMDAzTLBGMl6SAbdsk36NPPbkYMgEelaKWQkVY00Oh086AjPLn
F2GbgUNN7Ddexq9Y+lI777mW3f/2C+ImGHrXWlavgfLWcP28q1Bis4pJkI0jVj11yXI0wTaY9WQR
aen+fih53/jK6xi2baAvhufnLcqGDb2gKJQhgjZt7325PPnTU7PD9B2paU8EbJQjr9fCtAbsCxi8
5VBp5XXYwsOK0hvBz2fW3h817Ppv7vLHrRkm8uSMBunq7lz2ClytIWKst9dQLQ6Vyav3bKG8Nel7
WRZavnQXQPIrJ2bhOixgRpZoJhlc/eIXlIKct1fLTJKol0KcXYqi6vecgIPxqiG6USURPQMkDLAV
HIO7JIJ9LAMV2nUOiqkihqT9zjl4V1SJTj8nbh5ouDo1lhgsbZbOHf+Rb1+9twbv4U5+hyeCyMDk
zOYgOo4PDHE+nKmIIhvHeN1Tzu7rWPh6e3sk/piYEh/AT2IadqVffhZTdJUQ55MOiVJxnkQCWe5O
vv7GATRc0IEvO+udehwgta3olYnOMoIW3nFo1fD6yhML5hTqVo5eZAXJ6q7Q7S1Ag1mEnyCiCLDW
Rk5GWNi2TVKb+HCsK5caQoJanAQxXInpnff+kAEIhHq00W2EUWhlzX+XIyV0aulsZICajhAMY8zI
ftsYj48+7LWwLQKtpN9AR4d2lfV74ukX8DF2xmnj7fS5euU50ezr4yUKXxn+4VZ4/YxLONLIV9oy
oVJwHPxTR74EJ5IESLz/wYg1DeZlBu5nIP+NTg0Ijm0BzcxeVCe9V2Ij1/TtNr+pmDC1J3ULd/X1
9NaSR+A5b4AcLBkbwn6k/Swruiy3K8Acp+kvdLl10yxpbUnJtaHH6qsO+lGNcewrzdCaBTL2Fz6c
0jL34ORUy4DGLJNpq+TeyNlRTUpEI/4biVGxY0s73iRNNdT1W2ve8+wTWo70mtqsJ7sThLK6qZ1c
EMg8fnCG19wk1OWynF5/AKE15K5bSHt3IZ1ztfi3/hxGdGoqH4ZxUKOUo4tWnShFs5jYdB8jld+r
/RqwnL9rs6icc8+L00+MNJwq8yOy6ekow4w6KGfWZJ6fBk8zaxb3atXGb4SmZqVOsizGLYFr5kPa
sY3uSkMhoCimJ1zmadWY+qGsj0/JjYeLpeaW3DbQWiAvEybTRG891BQ8vyZEkOrriOIJeJsZICLM
pW4NoNqNIbcnEhGBA7ju0y/jjKiYIJsc1fXbhpjEAhFP28GM4uD4IhMQatP7kPHIq8lEzm18pJHC
/M2aIpMiNLQ2TodDfLS4SjrC4w2kt3jGoxpgjLgcgpk15Dm6iu7+4KZV7uCpCEfmPIg9qa6IdYh1
UXI6GIXbWThV7w7kCrw8DpUwW82/8PxykRXqnQF6iO6M6IuFcXLz0+jNKI4WOsmdoM590tRSGL09
v8g22BnpkCAizDzpZ5VnppVCulMUPrlEVXiXQwx/y+A3HjVIrc3fROlZ0TIJB2au7hdD+k2fZRqc
M9HP3c/kx6z/g0MDVLqgOzPTBQTZotO2wrQjkJ8agIylM/FzZz8TsnJKZzyMbs4mF4mOdf1BnQBq
An8WQgn8sc7WgQpeEcA7697S0WbIpZP+l3EOYw4u8mPd+6eyXeC1N+Lqi2xqYhIPPgaskXRBvNdX
oMWZrmZ7DvMxmEIsG4Tj20GhOgAz0MVguPQWjZUOxoGozC1FMA6tPdblLDHhPwmk/xAhIIaABVUi
eM9VxS+IJsh+Oi81HzBXaANzzX726olu8im9bo7lq0c1OLEBNuvm893RL2pXbbH/D7xuBa1uaFqy
wvKhRPRobDewm3yGmWF7NG5otH2cNDwDQ8KI0gmh0P4ubaFINBYUh9/YUhfIQFRvETSWiXVBMMCh
2K2QDqJOpBHdTEtErSzE1XxMZmlvmN9yJcQi5WJ4ChqQAT7e+2PvwUnpfUuuZiLiybqMh8W36VYp
sxtIsD69Y3eSdDwBRfwwhSL5Up22Wxt8yiXZ5Utu+BXri9QONj6gtbFReERXbzmPllnmoySi8SZt
CNWAiaHayGGWtH5g0o4IIMgrZKABrS4o2nc/0ueG5d06sT7whjMuHuC5hIJIHrUS6gsCVSHQq6nL
kNE4a3Fg1sQmcF3lJuAZzn9uwGh0OYX5T6klLUHLc/2Qa6oZO/TcBGVC9u+4C0uF2E0Dm0TDjxwJ
/y5rk2ucij0Ai3wWTMeBXttT02bDH6z2dJ5q9W6s4Rff1SnLbL/OEFm3Ex2mDlcnLccSSa/wXSCQ
npf5fyaD0vLBI81u+OM8byjvTdQx3rZDBUmcIWDJ5sIvyKVy7zDPyD+x1M0TNzGuneyjYFj89nKG
/5Qs585t79TaL0nkKDlRv1pd9WSmzNv6bF7a300gb1bjPLM0AF8qKfyFVLNfsS9a5RkFwaT/wKwB
2l+oMvDgQNaZBIhS8mBuChmjjOqzqn32Ng5wtCH/faenKRBGPQwyKkh2sY4oM8VIr6btCsrTZJrg
oswlRC2SpYkxWq5D5Sy30GdFp0ZeQ8QlNM1EIRAhejMdgYaKjGihwRQIEING5bNtzfTxUz4S1aIt
YqSNjJgmfyDXne7ZitOpPY394cyJSN1Ct8KErH2ExFSMIKGDdYL5BCCB1uZ9I+ti+80TE5/IR3lW
1sMUgiisRNT5CLZf8BF6JezPYBCPAgOs9dHvJ0fah7aBwrIuf/pW4OMYPR0eEDGTU3isic4+HhhR
u0YDhztApOJd3K67Kjuy6wMJn2fPgnF6v1deGlaxXyp5kJM/65ZMSFbCT+UBrReLeusFotlajYoK
fW1jV+Wv0MK6AMUveHEeK/st6wuQv+fP/sA8kcQIux/OdG82JWZY03HZXY1AyMPLXJsaQcrGsfOL
cqGwcJd1OglDgjdhaXmEk0tYOr8biqSNN9uXP2acW7u7rAxsG3gn5oGi/wlhzMLjuSablluzsQAJ
IyePmUobciK7MuPws7eSNomzi9js+6qw6FjZgozVxD+Xdac5SIq/4s+7atRpqNOEGpevbbDAxKAC
B4v+EBLSVNqR9sDmxHlD1vab2HmplVe71SnhaJyJpwu9xi9zkfpCjFWQeM9gKLixonB6g7rCd627
urE2VwnEGHiDUr4kIDJPuCMKhhCF0324803HFBKXSs5kDB2sf7sFYER4M/lxnfVfOJqa7lcm+VfA
nzSho/pi7fvIgSgs00/IwBGqIZFZs4Symz65uXZr5iZ3HKx+QPB0DWqKtNyWth8SXXnhgU/Ufnai
EMiY+RnVIXqgvPdK+cYrTNa72T/+VTt85OzWJ7V2z8pQ8JwGV/l3WEKg4/G/Lc6gZlWnYM349s8U
v00YhmqRB5RAB5mjabZGNcwozGKXre2fkRU/iYMRrosEwjcNhkJ4/tPx8T0saaUjtzhKAgOpcKX4
NRYlGG3ysZ6vozoUijgXP1oytULyxzvThrOqrXhDYcj4bb/9NOY/1uFks0WdJGe6PSS9TeLAuiyJ
uBGa/ONLXpEIO7KBeaN+0urBbC3GRoWLHthxN4NQm5sWmsF5SbJk4JNNaSfMOhgKrlTjFJQfKvUc
RZNuDmoSQsMb5OMn8yD5iesJUrZlBAQDjWKsuF3YiRh0tF7X3VfVpX7j216CtE2EjA2FQHKp5Yxh
DaUveWJhG86/ptl4LHos4nWgLr/3aqiGsDIHKQkIlFhwuxhnO43sFs6bzGJsifjXBvHutNdSD79L
CE9OXxgxEgPItRQvkoPRSfsFHhdqAfpE3ON47OGe3FtG5REzyeyFmUh7k4fL7KF0z7oP9id55Voo
b4L6u7Dv6PSmmqxvBfoH6oI8yJEJ03FuXwe9NTmlzyBq4pkJvs1poK+FOBKous+V2gmibXk3OjnO
ytJ+MtFT7rY9wFt69a/Lohu+glwTzrVF7cIdhqVp26LPATVZoGXIiMK7zO+hf4SIEmmwwlnu2FJw
zMumZzuF9BeAJKath61LlKtPGmq947BQvJ8MoGVP+A33tgNkTqRFXxdORBMwJhANCEZZ/GIY2itk
OhZ7ib1BHGzoHMUfHd/9g1oMxP1/4KmC/irOJ5+FiAaStIgtJzQZktjrfHwLnE3NKQlIJ22tlTXs
ME1gY9kFAoC2WlhXw5wBtffSiKz5TjgVFRqNlJ/STXKh/zVzdIkeVb26YGAzbmbTtndC8MWJOcla
rczU0rUylnzos+h57icOju1iNmN1I+APAIgmwYDkn7+aB5lylpjCrGRJrwGCaakB4rlGWo5WVUaT
a2Py8Jwu1110NVOp5ztwMrzm3UR5egjTJ9eU8vcFYZfsDQsRymM3H6JLFZsqtSfOfXrRenypNc4J
zPfZ/aj/OQ86Wg4L3be9VK+WxQ5rv4YXjaz6Zl7+bjXPu4oEe4UYQqnmgBFa7tGO0x5toLCBV/Qe
27UbP5BJijlZMFzxm7F2APoYsN9glm5bgdmLarSCMZEZXlHy3t2yMxF7B6aA+6yJCTjxlkpL45hx
jX51TY1gx104KlgZ+/H2BljXuwiJAvImx9suQM1Z57qpweSiDKlwYSGrOWlULY/d2UHwiFt/UUun
ci/9VQaCBAjk8drS0jkU1NTQUTpyXSckcikRBuWjssvC1tckOKLfoZ3kwXldilx/Cnco9Y+RQz91
9gZFxv7falOWV6CID0yvh4r8JPtLoA313zGNHQa0a43genAFc9Fc887OgtvXVAmfvprdg2KQrDmw
q7dO+Ez8QdDUqCFrhg2U6NeXi7N5fbdCa/OYxxZmuxOK1/WglmTA8E2a6XE5/s+l8dZxubOmwu8o
Zw87Mo9FGUFsXMRx36On1MOh+UuIWbV/HEBFop/b9e9x3FlL6dpWOf5dbS5eSXZ8OWLtHpp1QgL/
cEjd/koaGukE8tH3p7WqmNIpoBQ40ES5lvbKjCX9Dl7dfZ4G0WmCqCmv6MkAI/OXJ0nMn8uBbiMU
lJWL8gPuvyztb/xdqL4LEvs3w/qTszjP17j0gNrn9JRF6mh9vhUgwt8TJlq4TDijYWIg0A2Q6KvW
bpYFX7IV1UFaVGqCR3xY9rXIJ7bhK6zxTxkV/R31ah8dcLYAv6ws+j+QJqMNEZb4fNU+F2EsM7HT
5sVu+3bNeZU9bNf/DFUV+EAocgnLtFF4bzb0GIfS1eQ4avFbMHZA+GS+N+4LXKYMSpJT3fy7HAyl
UG9UpApc0y3FBSKuGJ6PMLwc/MGwkecR9BZsicfC3ubf8a7ZBSvxOKgLc6Yetk4Sw5+YDFYQt8Co
aDlUGonrJtq/AUx5kr2JhBKNNKXWun0njr2G/um1yQw2TBOkArCamo8KzOKWsRaCFhit5uOW7uBL
aMf0L7CsJp7bhRTH7AkFmOMKca89zi+j23Kyz5ksgr+XIYt2pd0u4EaPLxTz1KPat0lJ/tJ7BxTZ
P4zKSq7v7YRvNM2fmFMuf74FsV2//wSJuDY69u+K/BzLQvG6tJVHuTes+SZUGHexxfVW8ExwaGtd
oMfmIGMmWeSd1pGiyvT5BE4VNX8aF8zqrhQjs7lOEl3zJy9G0IvDY6059SxfGuEPLvF3GfqwuE3a
YNBCldE9p101o1+jkj3M6ePIL12WoyTNis5L6Mb5VujVr0amEh/ZLZR0WNTwFLMN8lR1fiPZJw90
FgtFgcb6rd2GphewSWDgGnAFXxcVXD/75uYl7gHxzhQQfT/Y8Ldgb52wOPDR5eVx0wMXF4lWPQQ/
o4eInZ66oT88N2kmxw0+T7UMDLG/auNQTij2SQeKd+gXS+NaB1Ztmz1i3QP1irs4TbaSDX8ipOGP
p3E5yXFO9wxALq03/1mwWZiQVjo1gfV0hpjDd6djAwYcs4QVzkVwi7+qsOj9D1swv166Zecl0Mjy
++ooMM5xekxEjIJULFrFtDpo+PNbgERmVlHLJnB9y8W/HzY1a/Ukky5Z3747dNfO/lbsLrIXZlKI
iMpswYNTH9kd1y/daOQu2TXd/0yspXrbj26LoFBucfXp/26bRfh4yCjsWvNutt1Qg2D4beyeyn8e
6si2mdrMe+8zMmaOtHMCcPq/n6B+ApA6uexPdegwypIuXlcBj5l1KyLEGA/5yMaFEOHav9W4d70p
oyXkVs4oXL8olAWtBPQR1EJxuOhzmwDeVpXplyhUVVZTSh6zQQHwITId+DZDQ2c+fiVprsAkSDQI
Y3x3FhstHmND9sTWLLvX71Tiq4Fhaj+1ImNZTupu5QZKM43Mq/jexIPb7Q3Tq+qZIwizBA9zxFJi
xWKmxDYGXhZXouCRoVK5yWm0p0M5NyaZv96whHk+aGZQdXC+IptiwEcjQYVcTvEovKYMGGNiK4bb
Z5ygx77+E98jLYw82lOSCVDYPm1IqttztYwJr/FpNFoFjt8A5UPuqqZGxI6N4TPgBvMYdknTXVfE
7OOvd/xLoAQgbB6RQ2T9dZOekxWtVvZkdzIelmjlCmsH8ynx0+AuDIAsziAehxtIVTMi2Awn7Cf1
zE7FspavJqd4eDzWXmL2WFuXn+u0EHmOxWldXP0SDFSF/UTgH5uwkrlT7juKD0JSuC8D9ahNaK7f
062C1zYe6lwZHXj1oidQKwXg1id3HPW3uwMGc2Z9sPMNWGb1K5X01WmFrWY/A78+W3Uka46uAKLS
BPiLj4o8Ql67AoNnHPhTJM2AC0Wga/YvTj/PwXQOniv2GJpQP72pd1tMoHSRM1HMW+4EAd179XbF
ug9l1clvKE8UaSG/n+TICnIm3nbmOTOXWQIP+lxbp/qZCFRpw/EGIpY6QH4bBjfkUYafTJfK7Nsb
KLdRwg3aK/nka5X1MhYv0eiyoFn+vv+NFHbOO6/lUf8xZO7JzO3nFQGp8UijH4Y98bRfyj/CW5fO
onGVO7r/LdFt7BCNSdanrFtoU9p4gUSAsrbnsybZEaM8ESxlA7rtzw4y6nTvx/DIAgg0FBHLDnP4
XVX2qrOipYxqmHUIaQTbGmzDH3G8aHzjW1EoI4c2C8EPxThiyE83hqmfAIz23gQAjh26Dye9PmdJ
PNRYp1npdzW/sXFMuzer0tCqhkLoFjxfTBTFwTTmYw1HjS+wP3bAbJ5crzwq0hfLZFlWeEsDgxDP
vF5SmxKSOEwoUFt8+J120rdddhW7ZQjjNVkhkZ3eiDEZPhUkq9YNWRjLVY0bKl75N51NnW9VKPbo
3k3UnNnhHjAQMkWPiS25+cgzIT25ZhdX+Lbimj5zrDVnxRvPd/63L5Tclu7mgRsphZCMLE2tH6gB
9WZYlLM1+ltIabCHFiBxwlGz+kGtpvRiixKNJapd6PoSLf4gd0+nXWgS+SUvkgjwKhNNOZzLAqFu
N/XeVf3InGCq8nnRLjYaPcnk66IxfNU1vSunBDpKPzQ0omPP01KtvcgAghhISpl+XmhzA6hzLz4e
nohYNRY7t2exbbdr4kfMyu66wkmTf+vYpUQy+7szA8em/1PqjtJYnF+Yi8YMwPjYfTBKl7fMUmsX
xMgPLKIKzgvAP7VJtpiS+eTUihjBuA/Ie6ATYDYojA78pA/wFCEZeTcvUzZUz08CUT7QUUaZRp19
NibBOEVe0XRdPLzFgDzGpLOxJlMm41V+ecInk7kRiwYrZRbv42KUUxD/Fs7lKTCPMtJViCyTQIO3
gTv1vVHas7WuPVEDqBXobp4k3phHX8zqWzrJ8Mu8XmwUXgzVOUhVnA78Yb1spQEc9z9cdUFnCxK0
XJpxu0Dgzer1u4lb10zwAD6QU+eKM/IM99KEe7anTncBQ8PR1IAJD3e5v0vNr92zyS736Jo6t047
hRzO029Vj93dvB5H/z7w/zy0OJlH7RVzI6W3dsJo3eRx6/sN1cRYRgLsErRnjzRJndnvWCUEVjAI
oRBhUnB+UwuRYkvmKQtobCwGMrWfv/1sXDrnUkzCWbNrpAU7EtUyked6xnpuhWHBY8AGxSrHYp9G
lhdxIXTrMiE6zb+0wIFuP0aDSyzSeYpOdbBh6gnJu4/VIRlZ5du7sRmVE+Z7Ys9RSakuC/pAdl5o
S/D4ZU/exzpOIdEwt1ON4/r7jdEd3GtS0fdtjIbMj4VHOShqndYofEQTxADen+9fzu5c2NlijDq+
i2TaAO1PZFPhfWRGEyaNCH19wgQnjaOqtb9DmTXNwuYMzlXDdLvs5feHr19TqQ6EsfKyVBTgUSe5
kvvf7RZaRBPfe3AiiRzm9UZdewQOCZsEcoBgc8qhobtMojZvOZH8yei0gJs/T3oCYZqAWCEKtMS7
7ZhKhy3US3W8WbiIumNAIhtJDA9ldqdeDkDWiY0kxE/CX9S0MhgL9k8tvDrODpJvupZ19OLGB9RS
CvDBKPU0gfFEreT+LS/u5E7AzJEOAmHIrV6ddxXuG46GE4lNDRU2EzdRXMibu1kOYgfHknGJqpW6
liqbmgFY4f2KCOFHD/XclK2Sba7WgVWPcNaIHU9ue+hWX3JpKsVSE7FRRoZzzPgrOc2BeEwLueYn
IaVw+AFrC/fNHYC+NOesrqkwQZaaEUCUU7NfwuD2CDm0FTbqA7rZl3vaunxhxGe2lrsYQSk1SR7H
K10hAcVYILNh4+1/xYepniWz8xxiZbUSWIUMA2WY4ghP/QehbwsyjTxmIzc7XCddTwAI/UT6s4+p
cP/p+T2uUUcW7kNxt6XWz0Am0+YMkA1RcyK0ZgDYGjM1ToenYOD7n/DwFGLeYRBT0ysngW5Fjph8
AccXr/b5GASSehsKmABNzAhTJA/LAu2RyaFKl0zEv19g9/qL+aNG6KaUQCvW7kVy3CYE4YC2TO+v
S5v1KgUfwpdEk9OAhY16Vs8E1zjbUrNGaVPKwHCx0cvmWnGfP2T/bVuG2xSwaA/4CmFtt15GYwdL
rUf2698WcpePAKEnr+jzPITh3uqgihwCI8ILz1lSscDltQGIEvLhsvmMypc+utWWGR7elY6YBvFB
UME4yn4SmwRDSGUiA63ZXsxGzl2UNekat3BPnJr9QBXLMYU1bvNBpPKbwXzuwWHo+CLcRxobXUtR
3GpcCac4TBQn/VHOSHYBH0gYjYLN7kL5M81hpxuaIMj1/A+0Hu59gM5tjk7SIf5G5q80IsDILzXE
pb/U4qJi4jLh0HhF6RE/0dSn1Fx2CAeuZaRDFJEwHwRPVPT1yrNzgNNhO8DumEidmZJ7fNyuWYe9
2ilwh7FTQsRnaWzjVIjf638JmZfkkJXtl9stYbw2fRFYoyULHBVfRimSphHfqUwdZuqJk4yyRcE1
n5TYPqoJrGluEehlNXls7spgCvWzZwLz1FSYpXaohalj9P6guDHs9x/HRB2Pfu6RasmJaSdQKjwW
A7O3BdepGhX+rUoEnYFfRe/84g6al4NMTQqIxs73ICAtt3MsjHm1DhPnK7H1U3+/t85cT5HagAwO
A8T8k4vzVJpAuo5wdyP75ZzGjsdt0OKUUdZMwp34rL7Am2c1PeXnF7moqUiJE6Dzlj5DlixQk/Ec
o1tMw3/EVBW+uWcdMYOQh90sI5rYNVNJHsEd/+O2eLTAryDmx7AM3ktB5LRmFdq2APn4Hwjac+dv
r+9GAuLIfPjVULwGWpMjZWMJU0w5XE1L1H1HX7kQ3da4+0le6EKrHqH0d8eEx7a/CRKpXsaaJ9aj
a4oE7+ii60yU3UcUKRkicWL8MBPluLb9NHmthCNOkbEp7ogMipV2IhAC/3D+hOO53+1Agjs/dhZM
L0c1h0xT1Po3TycAAdeM0C309vKYOFYm1kM/hflgmO7anYbxp3LFMDtay+VvfVC70OjJa2JhAvP9
7WHlTpbT5NGrbdjEY3a4yqC8ZJHG/Md6It+q5C7QS0EsrG0plJLjI2432sk/6DC5zNs950xBTB71
titPnkmviKrLyCOLRsZmRvkc5uCpK8L2uXw7oM13HBtScXS6NTmwcCcbptaGWo9X1UjT3Mf0rUn8
bTy2PNVGdEGxDWPEnKgA43joyXDxWC/vG9ekIQ5FWvPUomFtF/czCBSBOJ0ztxwd7+8TFD9zzoZH
L5XP90q3zkqBlx2QKKZrlKObNV8/DDNSL9EXsxYn0v0RsoEsyDNe2endxSAFO5sEAQDvU50ybC6D
Hques2avWOe8qeCRaeqekiR+Xdj+WhUcbn63UyO9JAsClmPv8/RTXLBpcRN6ORW4J+Vmb/ZUDNHu
fCcnOX+fI800LxcdiqX8J04TEg9qcDwhf1mZLNFJldkPktVlvPCH6bT+qkikBvgAn7sVKxkEBMEa
6ShBIY/bv2TxsMpcFEMnC84m3eY4xtJIAXyvbE8p9+2GToBYAXMqJbXwuimfVSoAMRuJt5hwaqUy
XjOgPdCDgEdZcFQwB/G7O4hoaFp4D+mW6JPMocPUmuFN7xyUBKVTEhgrNItaZAruhwuKSCz+sdXg
0aVVwLEKaO6wzQ61nNEle6FHWZSPWAs1awQbctvm82HE//ktzL89cE44gxoHlSDT8qgCbqpIcarT
5HqtMl181S6yMIKOo4hOie9j0+Pmv0hsSvdVJI+Ec08ZxfWOqn608gwt+m6RV2Zo+OvCPbYUCuvr
RkvB2RWsRnCCErRlTsAY2Bm2cVTlYWqntNKI0DsSymhTlhqMDvzR2PJOqFeFIx+YMGSRN0hCtI13
brsKOHweszafiik/UHIbOulwV0GT8VpaNJjzExjfF3aEj0jIsB8NRI9lLcdn5Y/IS2/14227jofK
6lorOftO8lao4DLcNraLZhnB8xPJrcHbycUOcf2YQluAAKAHukqJnyP4oMmN2tAg9PWUH/IX+3GV
41uP1qxFClOGst453z1+RBPAaPo6KwPajBDUaYKhcw9n2tRs96gbwdVKvdhRan7o69kYyICwaaRQ
ktNoVUIC+iCidXtD/xIOp/nB0FOWWJ1ASpwJ0DDTQdJhv3RlEI/t0IxcLWiDMCSQntRonvBBJ6FX
OaGGDgE9BXh7ZDP3m/ihjiVVI5zWlkXHJa9zu530pD+1qOTZgx5YOwA+h7XMg5LJSSA3ak1tYGbr
gkxp6daAkVeQ/o9dFg2xtXmWZpXodvVzLSitV3Q2xX2lLF5HUr6fbSppezjafIB7g0nY+pC6PxrE
o1swhH6fJCQuO2dXyJKX72D45sOS6KUW9k855nVQ/cZE32EXH2UJGhtqea8m2laBn3MxZ1zoo7rc
GTfq7NXW3lcX/OrbDNPVXEp2fihycYs61/jwtEFlnzYsdMqzps3Nb4uVWJBkxf9MPn6rI8JLmxBO
SDE4MYLXvizyadRdIYvvnqLnDbiM7fqEPG6ikjaZP5aE/pvtjhiCVN6lkHfKl96I0v0z0JhhPkUq
OQeQ8ydWkpkbTlfo1HdnOsr43zQosz7h4jhBj7Qw69Bpr7Zj6lx+tYasE0CL6bfIy66DejmApJHl
m4qzX2REm/KcRvb5n20dPCigGTmXFu6hCybDWakR5hATgMhcccjQ7eew160VEju1F8N2e/NzSbLQ
BGvie3D2DMT4G0m46WtX+HuntkreWXgvs6LkhstAbk1oRCxo5cCYfQqNmPzoMoBzPWid1WD6ZQFv
sN1lU/hqOpaDj8WCzAWpTyUaxvp3U4ebdUg9jNSVqHJy+iQEOW/ix8yqQ/Xy+j3Ioajv8TgyBJMq
WvBJJIk1ZWD3yEuRkCqJVxzUBMYrrIfMFu4+osS6mpjABILYd5gyY0koaiCX6TfaqTWhhqMEYfL7
OsoKLQWW5yDh9GzOoNs1zdBBOevG1veyhjmyGpo5XQ6dyNOWktwUq0fwrorVmsipaSO1DIlqJykZ
M1ktQ7dksktKgIcIs0RMVE4gcQmSzDZUA2gzxZOXwXsUhMxtTR4t5+V76IpzneczP+HWltKZg5DX
jzo8leUcXYDU1lD40avrofdsl7e10Agwp1ygw0TSdLi46bepk15PFHTpLK6g4aSDeZ6XqEiIC9OE
Ldhy1PvpS9vWrjqKk8ShlmGkCI5Ezh7wlCaEF1bnB8X2w+DFsNMluJhzCapx5vpu4DQiCivN3WZe
5NaVE8Dwgzzqda2McC/SoQL9kx1x6aFKWnw7c5e3eeYMDHYkftYLbUEgOgF/Kz9EI4OhsWOMGsTQ
4GkaisyvZ6ypZ+cpYazYQIezkVOy2dNMGsWujJyK3VHR7ve6ZoyUYxF0dyktLnjKTjwZ41UHxLYn
THQLGzdmLSbgIf2InyUgPb46JGVmO1OcsnHs2rorsjmLoJ6TY4jvsLaM7GODnNXNtpH9Dy6I7nqD
wptGmeRQgj2QtTatjzEmAvoT1xR+4WEKCuu9jnl0SKes7yDP81R0fuiFNKzBWmzL/GTwRNW1HjtC
GbWXrV8ZCuBs+gSP/FL2RnGX6tLWEaDth6tF7Nl6Qxyn31Emo55EOY/Odj4FK8dDD9tHIstB3GG7
18usyASJB6uChpK0FCxD4tPZ63kER0q8w5ujtva9oztFVaJ2mVFvWh1gymsswP7okluqe7v37JN9
YNIZq3aC0XCpoDjbceQeRK1HXMK7sRi/iY0xWAGCajmxPHe24Z1bQRL/GP3XLZmGdXTvDsp06W6f
l4kFmFe+UvyJLZBfoj6xYb8wxTQ2cZ8nVWWqu21DNhqOMRYcKWqq2/zBPkLQWotrlofKEMzxsvR3
qLLTtjduFSteXh++fySR+CXJ7m9xhdSw+j5WPFeJ0ZeWvNmNSZPsiQfo5zzWz+8UGfYGuB6fmjdk
jN1/2MHeqmkqO7jacNhaZPO5OLOZSaYwgco4gKORzvSHT9WGsWAEENaozUJj9HtXdJtLBS+lOwF8
FiEHxCAqfGe0PI7cDzcjC6HkDhyQYoYRuWOUUm8NJSaukOp+zPGXpSvvIBx/ngKs+sF0MuXsXZIn
Ill5ssXjUd1JAGxI3ds733rZ5jMWWKaS75X9dSoEolrcmZZKXXDLAzv29ddRAr3iwCVboHMjzTTa
nKWS4mE9UnTMV//DVw2vev7e/LtHYCTMiga05sMgwZCVAt0sQ+oFQ8lHeMFAskSLwJgdT5h66/Cl
YzgCbKjtg1LCTXB5gTRfWqaGoZlS0SjlG3JN84sq5Htde8XXjV11b5LWS/C63hkz+tOQINhOuy0n
RwE8+vizOKQxNKWmk3u/aUlNGRGhSghqj80xpyEkNbJ2CIAXSq1lqDzF6cSZFA8exzpPDnITBojL
wnQ8atcpvfIHjZKYzZuhZVAAskRz+CwfVFUVcM8dQzzu9q1hNsBpyQ4qMWy3AERvv5zDobDJIONF
3J79ZsJ37dWZwKuaY4Yovv38hPfe1cYRZfkIRKV4DWGnCAUR37+BFvSyN8nNcZBKaUhCFfvx90Nk
0/Q1lybF4G8OCVX1zuOD30wA0OEkTrBUfzTmyt/+tblVTyk65OjmaskXgDVXe3SH+YELw5qqPNZl
TeMYLlNkgtyrCdeEyL0RoGmPyW6PR1aBCYJYOZm46ZPLtbMkWE0WQJfQlocRxiXTIQ/W60LURm39
9AEUOwmOR7hxvHkeSGGsiMnQMMKkqHvO27x6bVBkvZ1kTs/dTJQDomK37VbUNOi86k2RqYTQr4i/
o7mAAdjqqLYGk2FPswTBia2Hf1Ws7Q0to6NDVfjKCbt/jUb9U7ETRN2oXRJwTNma9raZc7y9EEm1
GwLcej7gbT/XP3or0Wfm//okBD+5wHMWR3BmxY5LA3gtUzqq7Y+cba0M7RojRfkbGzHiZ27TU381
+bu05mAOKF5TNvPy35A3RGH8qHPo9E04uf+Jz6xWbCdcjWQDDSKmLLFQzehCdTdtRe87tO1PVek/
i76c0g6TXLvMArnjfQJ1xWkpHqqqJp+zXQMSihX/JvcozYU3YLOGAPcDcEuGosaw/JLXgQo+q63N
MlM91bwgqN5/uX/YBFBkom6btmAu3rWkvHfo3/BgpfmW5lz/YZ3yF1V352BOUeEdJfNuUBJbeiYh
ENb2U7F1FJAFYvwo3BfIg30vpmKQmuhYTdIGW2krDS/6T8dQ69Sl+SrGnsyJJk4GfwCw7efE5HOE
Muw+yt04uEjSqYItUw3hJaB0kQLHpnk1Q7YEJObEzUOzvCnWazIhef8hG89uPoysLM/eu3HGd5ms
N7WAzxuS1dbGgK6H1YAGpT7fRbm9v8qKqxB5osq9j+yIh6rFi5eceTjxVcyfmwGPx0CCsxlJByPE
Q1/PsRuPa93yyzbapeZtGpqazU1UJuL0NUJZBT5cS5PtiEladFjD2o6tiL3o0Nb9ugm3YXE6YVLw
HyGq5Ypne4cXdoP7FUXABlrxWzZXdsVRgtpJHH8EaXK1YP5ooBv0nDQqVp+qNItOoJwUQj+GbdZ6
0DMziyLgo5+IZL3gd0vSzRBUHz+Yw+Mc6Kqq0Jhw1L0wi0h5i8bS6CCNQ5qGW5Vqqz/zCMOyWg5Q
5KO6MT6ssHpTSvV3FtyHramY2LcklPsDqeGc6ldkV0hT2CfdCJ3qo2hopCQ1VB5JSiprVd6Hb9ZS
r3dzysp9o1UsRMV8Rz+h/OhSyQMR6OxZ/pE+2AloMpeNoVxZQk0yj6DYvFpiHs9VxBIF0KPgxzFe
YPjbe+Zyd4HRnuLSc26+1frYDm/bCyb44YahUuZo2hSehKyqBkJI25MRjErJzCItWkvANhce9QR5
/n+PZSXSFYY9G1lYeVZPXrV88v1eW3Y9gH2H3AV7yrzrzV65XG3SkX7/muOPJXlTxBGbRaUiM7YD
TXqepXBfWhaR5IOpR7SMq4nEnSYwZnot0qVpiWOJcOVvXs/5y05ohPI8Vy28sx5Q4cZPZU9RMHbe
FX/7ncQyUVG97N5qHTrnzjCNXGC4bFLGZs4dmNuqm6oA8k8XwFiftZQJi3m3TmmLMKgYth7wbJPz
Rn7tYhRnOvBMpxaxvvpJn6hxoZu0wQX92qheogDyhpT50msnZKShV1JqIGRNvAU3gIxmvE1EACya
rrs5TMy+RHNRkPTMXxpfJ2yKTxpGmDev686OAcncxHy7keyyL3NpfcC+Al6UM5zpa8UdUmlmyIuP
/CFAjcs7su3bJcL6Dgd/iqfmGXjmAXSAgPIc1nT86OYoQeWLx7wmD+WETIX3CvRE2bpUCJntNkpD
JYCsukS30d+BYYpRLs+1buMwrjI7cbGzCpDX/V1c3wyo3bbCv0504UPCHB4D8pgV0IUg3i7iwut3
Md49vHY0YVMhEKkhtIH7a2+fh0ZcX14WuAuSonyIjXBrKQf//nZznnuNUXOEh8MbIQ+G6p4lJAiA
Qx21Q+3up8NLgHzya+SjHX4FA1FtvYlz0clSnWsVg/05dAI52HIgTPQQiaWB/o7u4+/dq+N+/6g3
EqQOCHGa474fsMkQjl+QLaz+sCvTkcHxa4rleC4pXvlzEDGpE4ZCFbDAEIlYcng/4fok85rX+frO
61AzUSkcM1o9qcWqOR3uFjDTD0xApSEFn4cWlYvi3f0Ddg7LG7ZXo9GrYeFkc0Dn3LQgwBb8Fpei
v0QHoEeb2AX/Q7w7YKUQrEVnb9u1Rv1hTz0RzHr2mZm3b6fL23MFr+rXTv1pfFFygCzmmW7yA1WA
op7RZdOMeiVlUsZvIiASvqntMRTqzCUvh4DvAYFdljRZRxYXqzFuSmaJaTz+ATk7ZqBa4Yp62+zk
4xfWAEMq78oKFtE3FtraL27hVZ/S2DPu5DnLqFuzxWuJjMG2uKOwnReFp/cRKsFYoq2wiivN1z3P
lSiWyGUBbMu8CBIdGDhqwz9Ca1/C1bwkc3BjGwCHeVx+w+HG3ph3jkt18T+TxWdx3QAKGjakFUbe
q3/vTFrcZiCwfVzLTPwnIxAdpz/IYKqHts3GWCp/U45W/N+qvmUuQZsTKZmzNwZ6Xq6W/5IJoAUA
bqkD3AJ828MbCqXLBLAhil09M/1J2+y1HAKgzhIDwd2aM1P4vAAASj340Kk7H+xGWzLZi8/4dh8B
ieYmtfSLI4JGC7a8bJG6LFqU6XmeLQUkK74wpbm+sgY7W4ZSHmD2s6Sl5+Pjr5V+Af011gxtyjD1
bznvbbC2KJD28CiQosIgNEjyTEFqYhcM4of8rOwcZjrEFXmVrJ3VsBtCVE0zTnaMHjiJtD0uIaqV
oiJI9DFE4SeI6agHj2mHPMoSehoAkmXaCsBN2C6az1/bin4yj2bOD9wtFDRWkgkocrPc92gSUG9Y
JZIUs+6iX1qSXCtYNOoYlxkf53efrWl5K5hRNqhhVJU+XKFcFvAheayJkMCvMh7jonF+IDocyYWg
Lr6l8jU1H0+vs48/N4x8pXrZTXYFbPk6LL5wQGldnKXyz80phSE13T7zKXrZ2LAwDn32wy2BXwAu
YYBL+wO/tnLVnB6St1HrYdzVV4jxhLcv03r2Mq/DCO9RqBQQs4p/IzgB31toKBilR4RTysmfhk/i
oeqafUQK9qQYe2eb/gUIkm5mdsmEd95kcdIkZkAtnvut2LwQtRoL55DT7fzo+oU8a6ueceIr0hzi
IhSoUGCTaLz6/5xOZSySODv/hpiCCv2Vu0+QXCSd2cn0EDwLl6cBt8g4u7Dq7OPM82yYMf7H3ZT2
eN71nImR80sJBBJR5uev2FCukrGD5Wf7YYyRvvw9puc5tg1EVk+twjUEvVNp5N7vSpWjdaPUuU/g
NrOZuo79x2XfZiGoQayqEfnAdCgI+G7nzS1G7HOw4mfMurSAr+E3zNEhW0k/3iSwMREcPduVVg8h
rRLYVpZDvTA9wO2fOiURMSnyRh5aDl68tedP3aN+o0RO3vHMQOHzf3DXHNZXnGTKwPUTD0dhkKih
R3bvrwDkLLMjeLKh9Ow5qFYulFcemscqafHgLdrdYSb5ibBpcz4BpD0PINKc4M6IArjQciPSYb5C
fRrEUh7rsAhND9QBcKc/poe+HiKhcZKK/6XPK07Sjm1Z+b0JbUduUHfmgvhow8SDclRJ12nJtFCq
T/j0uaq4yPz4OKKYmd2XUW6OlEyEJ0gKRgFrbvtLdh0TR9sF8a6J/H/9Fp13re4LPVpvzZTqwCcd
4ow7oDWJbx6yWMrSPjIPKD/EDZKkWVuv5QAyh0/PiRSLgNU3OVocfP1AI2KkEiYkjd3dCh+QHwk3
lyIcqWz//34L+nm2b019sSdRN6eBW2e1OQeG5tlIuMhx50I87LJ1t/rDgqMVul2JlDSJmorBEb9w
xLsIgHPEgTN62X6MupqDN/viYLObg6UnwOPkHHa+dQ5JRXAc9rkNCOhw1ne6kafqFp64CAi9fosX
0Uj+lBQesN4k0w5yVowfsqXGqM5WE78jC6FeB/ls6qOdAXWumNw6jKPb1zwmz/HXjbDMJ2H0J3ZM
yngYg59B+GpfkxI1CQ3XLCeM+9y1wuwB3dpjI0npN1Qyxa6Fjyp898NAUOpJAksrqbfHr+BgM30e
RVAViQYm21d9BLRMiv0CscISObSnM6Rq3Kb8JFFDBxV1tpaSEzEd813ll5CzhBKUqmzhlpBrlW1E
LPDUvpQHjUJuzrmw5InQAHQVIEIOnkYMewGTMG98GoSwNhJB3lYkWPCO2SPnV/2LTM9C1dGHGN8K
Se5hbYXiel1V5HbVzThO+FTNiO0vjs91r3/7u4d4V6CxoafOJxIV1UAULO58/d8GvO4uCnCXYOpr
UwrbaaZLzza2b8pB0VDUWNVPPuiBLVzOwjyOWLkXlyqjr3eMu368bZaVfOh5vgoJ7183VZS6RRyp
USgWxvd6xBBO2GcQBDTDcooh7YZy2LNIG/ON4CcX0NLyT6g/7iUfLmLOJE65wyvURG12+NqeS8ip
43h/rfxb/rzYerQle5LNkEqZ1U0d3DvTldoD/9mBngzPASrQVCwGNOOTsb2cRTY0g03FvpRBt2K+
BroCifelmg0ETnuecU71FFcvJW36FtKWJxXBZ9MQR0w6f7hMTTtuM0py7tNXZZAJJHBzMGMNBWfr
pwG7VaQQCZbRWtFcT+ZqSCaKzFK6ec288Y97jzDrDDz1+dZidYiGNKo99/5N9JIa0IXStPqY9rGT
udNHutKOw+DRG45YPrQaTjrUZH5EC4i+kDtdGkp7SSzibt1LzyGP38hc9sJOTm9TTP9aEubQUF1R
dnNCeMBn54UdZUn28Gk2vnTKE1t5RFsJMuS1xH9sP2McXMfFt0H4OrlcB9kBUJxue0EBEFQPUIic
5kj9z/vZp1gNbsbEGYQoiMBuX21bfRvQxGVsOmAaQ/PEMmQ3DbPnZrJuGko8myLx/p/Rg21iBcUu
00SdJ/SZ9vkrXau7Ms3ybjctT8v3dNhuFYaHqkDwwLPYk79iVuiwwOrM8XYJj6H3/uFtefA9EukX
7KLrGgkQ+eSKWSqccCS1V7cuRdzSCwjFgXa/wy6Ln2mzaa5HvWaUkhvR/nzOidfKBONPrugGznbg
Nnl4yMLLcjF9B7vKhVV4Xzv0IZuIhQM67s7DeFyHjJGs0BrXaMUTPQ/ulvZvkR0kc/WFD58MLG/Q
NSgvCuv3wWkqfkrjuR9ApE9yMzJn8JiGCaKjPblSJyL4b+MgppUqhUdamOywe7fq0u+qSGITr++H
+shX37swVSa1GYzZztRMyhe/R77izp1SwMUr3JF1BcMdBZD7PG9s5qV9GgQSEr43INfRz2G3XUw1
Mvh22aJEWn8q7jGMGuODVuy9VEbBCmVLPX9qvTXZlI++sSDQ4xYPUJRJAORrIh5ctBb1sRxB2H+a
XGKYOVl2+H68GFjFYh/hDRbbkYOf/oWKQ9b2E5tF48JopH7OeuA66Pg8HcFEF7LYEK8esHMWVImJ
1pl0uHQi2xSCREpXpKbLR+K0AseYxipfQapyo89G3v9VTRLl521KkMF4Bbd+LaofNrv41Rxa6CvZ
v717V85r/rq6CR0wxt4dU0hlXwO51Q088WAu6dWDaZ8D9opRf81jNy9/IVwrrV04Z5Sc1muz+8Eh
Hv8w/oMi/Bdd7l6eZAVpPD7l1OmDcf2+tD3nSpd4XjaONbn93yZHzk/goii72a+vp70boBsTdrzL
NDcA63g8n938dtPdED46HWGL1Tbkuenry1Kh+oSVSGxBtLbzZ40Uc5at6UBLzrVmcmNIhC0PBlb3
Ypl6KKtxy+BxUM3BFhGCiD6afCEexXzbZxr49ugKWshxsk+q40Wv4iwxDdfd21nuBnptKk5ARShw
SYzkc4kbDcRazC9Lg+ZzKeRLKa47e7g67daz27+ntQWsFbcn5MM5VK8ejnRfJTkRydF62FVFJfbV
NCXPqdz3rLNhkJWx2P4kPS3SNA+cSGMULjYvzY5KmzYclpm66VTrbC2bvYlvwTm/+dsWu+RLze1Y
D9M/haPkbC/YjUxQ9kDLMylOvqqodEh7bYphaM9E5L9zdaLtG+ctLUCj2MXBhtCG5Xu815uucWQQ
WZnXRXO8avrRS9Xc5V2EDNPKbECJg2un8Sz9pywqre4i6yGs8XEMhTs4sVSb54/T+8AGSLjxp4G4
+m4FkrWlabLt6+YJnMNwM49plSUaDONm7ruWwqH4f1WDr4knMvpiIhcqQKI5NKEXNMlNC5vJrze/
ZFcGRIx7KXqIc7KPoNX8my5rpUqGOiu5inA+atJWaV3rlbeCfqqT0z9rWOI+Sz6QmXghW9DrGPFz
k/CvAuLpzhF3FoLrvhl3Iol1V5jqQ//ddqbQM94qzRcc4VLl9mlvf47ThrC0ue2lEMgXRDUZAZMf
p1el2+GZcInxyAw03RZ+hZyuGjOHA/8CsJM6t/T+t7gJU55aJq/+MfugMgeo3TIZgZCf9BaNngnz
xb3qzjBnommVMek9DDIuC/eHRQveBsBTrOZh8xyLS6zlhlIK7Dv+qCBmA5Q0UVEanl43rv9FpBUB
NJZbFFeLJbHwEsoe5bhOjOkyXAcg8igldhEEZ9PGpOqnvzUGQbqrB8sWBPYzG1FYGamZT+Xnj/hq
V5vOHUimXSdEaGjEIqpCLva1kaEOAISKCWyIA3LD9klEcTGyFrrkx/AN9nCK8XbBoGlC3yPg+Mpq
C8WM1NkdT7gd4/iF6sRtDTKGRTfgbKVEVMs3Xf/+wF1pzkqBUKN3mJJ9Wc8mDwJkQ/2b3ABKXu5u
hobRo+/UiEzZ48LfgllNAlgMQBVa5IOT+m6I7n9cp4w9eW0a/+jr9glfEt3TORWI/LgtniB1UqlI
UDjhLCxrSMDQ9FDMP55Pti+hFzb8buxAOelsr6DxizOEXHYCeNSjpc9mVOamhdXke1ahTpboTfSQ
FJKN4Mh+Ga1+/kLdC6bLOw0Aa4eTmAU6e+AB6UJv3v0Uta3dn8AlxklORT8+C2V2dOnGPkYxroXC
knhKpKWRu/BS+pOdW3lyD5XC8aI5mjmeOHcSDzsyc8v+G27EnNWE/GfizeAvXFDDD917xze5jULp
mhFPg6c+k3I1S8wXfFxFyR2mgphb5XHXmtytR7s5oLiViWbO0SqAr2jYbmYyvJhYNtsOILwcEZzP
vQKrYRW02fUpXkmFUAY1WNGSCP3ukqEwGe+f1i7rJcR5ARn5EYCpfdMTTc+kHgOcOAAvH4O3Cj9r
VG257bjPvPNbZqTsky4SpkPDGYM5hp+ZckjhD66fu/5LRZAJrh2+vbDZBp0ldTrpCPQh08toXjVQ
6v99c8zTryVbFW8xsl6rPvCFSyzzQ7CJgRcVuu5RRZ+OpEkup/x4oOn+9fQsepBVQjwb9GwPtD8Y
25nnZwDeQ5yGY870aMrLdrmA5pvneWdzo/YWJjpWgoSQ70dyu7Is23qMJJ5NJNUIcHCmI82rihTN
Se4c/XMzNfAqnbU3SuoQ3APCGap098/j36Qoo9MNuBq8/aqV7VxQ2cmIKZP4/c2/tbblNfSvxkf/
SAHM017XBdOw8EhaRN4CN7rGAW5Kqa8Dl9Svej+Az3NdTTjZCn1s0PrUCcNmHPZoOHFG6fHhFNPf
3uzR1c6m1ui48cN4gpfsE7KNd7s1Dzj6BwHRozzpSroVdpNnsFNUxwTEbhiEV11pZQLcpKZGPeld
Iy0cbjqWNPpDdMe9+QMVt6SRMdPEX4Gbw1hp1BgghGnClOHrdzmWW8wpmHg/KWW56Oaa0AzeGmW+
/3NHNBtbpwmZbKf3rdwxv1mcRD1jJ3Y/EsKCsUWrwj2Jq8ysiCwOFMZFKLzbQqwMistQFgns/an7
kvlaPPUGznOyi20wioIxqDFZNX+DAxcAnJpQ4MJb3aao+pDCYPikm0MTX+kH2wd+V7MZzPdAa1gh
iz6XVrgYjRBwws87BGYQQPi/BAaI3vKL37Se7ScXEk0GrqM+GdGSPv/sjnsO1pOIGzY2pmQC1w0I
CVXmP0w95COwi5jeRipkT+w+UfSXWwgxjBYTDK5gd4oxBhZhlJvSIW7ndr8ctza+1CnO3d1xDwfl
ilee3Ciuu6qpmArg1au9mIZtRTrEXgBt9X8QNi3jqHOw++/frL6Dtcpq+B4SoPl1RHGG+l0ivNC/
qOJhUzian3cJ8EZGDvFahbkTKJJP2jR4Gev3jDc8kb25BsAubinVy6HZ5JEw7BfXjTxCgMYXticD
2BjfyQUyHiLFjx1Q1DvoJtLgUO2MvUI4YR84YunKV3ULroOWQMvlUt+WVu67ohIzq5ybzzXgJTEl
kuwb4wI1xVLOpOVfeX9QQBF4AYxKN7Z+glNdMC2Nrs6SPyVXMvwsf5jkB4yySD3rbDt9k1OZfcxO
ZVNN1Zgxy125OfgHeFWKiU/FWbjxUBMlNpnTIgEJX6wYH+uxhMOfO9rGaioxHNTQ+PJQLtJ6HxzE
mc4dE+9OIr+DIps+e61f8W2ecaZ/7tXtQH87C8Dy39h+6m5efnbqVLS5+u1B6zlkmYESXKwR3Noz
lMkfb6D5Mj5fZNh/GEoizDO8EkBYYrvqPfLkDBySVeW/ON6RPp/unH2Ybt97niJSzYjW3RdnFUCS
PBcuUn0dvZTWi+r+JS1aG1Y0ZwtPgZf8rrF+fs3a3J1Wy40yu2W2ik7zD3t36yqLe3fLRixHo8kL
So6/I02YzjZRTLFc7Fj2SRW393aagPwB6UxtDac2U6yjCcM7stEHnn1yyDq333MIj6c8eskuyEIy
u1LE57vXiQ1mmmzGHLXQDm3ThmTUdR7vHaIiU+fRH08GRsNY5qTED7a8pCVVj0z+pgXDfrRHlKwJ
CfQnMMtgE1WilI7VbvVlES/cQq/5T5yPyy4fGSdgFRaj+0x6ih6KtR29aJ6RYLlm2w6m3MeMSChN
xymj4rqlGaZyiHfmHhb5GrHJXG6uHus13viYSDMSPLl0iva+zFwgUzWVJ/oIp6/xvZrmqGAHMag0
xs4268T3ei8fZAt9ReOKZtIF8RwsZ++MArABOaIHgtmGnZiNzbtt+8twrd/NGHGYn7GsU4rvELS7
j1FVq4hQhnuL5Zoqoi7locBnkE2Bg05S7tkPphE7l+5WfW6rw1AMHZLWxi7uvV+V3NgdQfVv9a8E
J2876YILtN5xZUspE8EuJO+DyAK4q22nvyPM0IIr8l9gm45SdZh0aSd5ouUGh5/O94nmXbN+CeLT
TX/Vn8w5+w6irHVg+XiKo+2gnAH6vhIcvTRzDMztlr5oUFyVXC8EkUABawkXz2yEgGoEeAyMudhj
zhwCa6uXCgcTZY79F57GCyy76ePAiYwTzhQNNzn0DbgsKhMdaYVcwZZA4zdjoBQoceY2XCvaolDQ
gJUK+ySMiLGq20nTXM3DjvWenc49PknsB4k5j+u95Xp3c58vNkx/Kkw7GCz3IR5UkWBHEzqBcnZq
SApqCOO890z3hgsSToWKmUqTZjJExf31ZeF89D545NK9Cb1WAptf2GLw/Eh3j54f+3ORerEyUagX
yDske83THcjORU3CWIFFw/2zwAqZaUc6PpUgUteQ10wjEZLkLCfHHvK6YXNhi2po8cQeQuOei0cR
mrp3AgTncLgRNbFCOpABOIiOkRPPgjDZfEkUtVdwniiJKYbXB+3KcBLWW8wyKIgSodOD1z8Mm2BE
/E6iaaBMFrZEpNRSP2TTAxZ/ru/gD+JPfdV42lymi+zaXIy78YH47y4XJ8cnydPUsUoIRGoc/8+c
Au1wKLW2uWlUHcSE7wyAUFJOifcyXnFGA7XOel6bo1xzXkucaX73qlv3j0URjAcbtAI6REaltVAE
h57LYLo3cJzSJSZlmtP2XRPR2LVmsG5olp2dobRX8NUaA+cbXj2mwc2UaHie6V0oZ86Y7hGjrEOS
lvvc8ULEFB88xez9Ku8BF0LJ1So8WJ9XYPov9PnfMwXJaieW6bitSCDVO4p2gmKrtEltmpTDIQ4T
sae1hx/JSgrR8ulUE3/yEPiAlozoimKbtCAQBCr59axfmQ06ZF/B3ym/58jN/mgkjny81TFjBKqp
KGh8QkC0/lRbnWgHh8hmUVb5/wKsOmMlC6I1nuvoagFfugW5qeSCAl7RWD3OAe+emnW/Em7DN1lm
mtY6EOJwFGhe6gjFZQbM6J4o6SZE/hW6yPp2Akhg7Ka6BdmlLnrDcHkVrAZxs05TqfJCh+E8u8rn
mwQbYKH+gxbUCQW8C5AcLOtN0VxJW/8nRd7z/gFWqAPPLL2XOobr76KHNkm8L468sV/Uhm1+jC8U
+ezeDewMhmKK8vvJxTAp5ab14DequOjk1Kl6uSQyj3vDdx5NnhfpIbRsvRZEIs5xCmMlq/WVtuyF
ApEZ9NOMQrkS2bRPWxc9jdCCoENyh5YtYZP7aj1EJyAAXkr62SSr0zYHvWJOGUzJ9I3CpOCyA2PY
4QeqVfM2cZDRMeosGKSjcvW2HoUkbSkPAGxGGp07/3QUZwKQ2LMud3ho14hTSRY+Qr3K9OrX/V2w
nxknSfmgwsKT4G91C+50xSZFCfcCvqMO7HrKlSrDGovJ8H5mPHG+NVf14DM0n3BiQI4fh+GF/78s
0CruKq8nAmZE+9GsJxBBGIE/l9Y6Y7ShpIIf/gijahjxullgKDTFgOkxbR2x+etO54BbnNVdt5YB
FkoZvaeLTIfs7QvnIO7XwXomD48/r+XeO5D9rP7upvH9ueSh3Y97K7/1DFLAOJ/fGpj1h8bZFJPJ
zqIPIZPX7bQGTJtAKNp3rN8vrlF8qlL7se6s8jD4sCZsrKNGrFeiZU3LWh5X497y/DlMuDvSAjWC
J72D/bySvJW0QwgYjeg94bs28mti6O9fIjNcDLtQYtluGap7cIXn2Nr96FG0eSluOujpREz7i9AY
zgT02rfEculBkF7nMPgRSzeMQXyl1YQwpkBA8BoWEj81pp+a1xusC1WrYH+XvD+zw2G5E2qrPKAN
OUt2t5h/JcqWdWgXBXFEZGhV9yBYu5/PE9uEJhcc6tWKHwdkWGZPNvd2lr03KC7uKviFYc75QaU4
VkJsDdk2hREeyulmvUasokzB5yNkCbouxRGveQ7eRfJDwcHJ//7H/pTLWjrBhIKYAESBw+HnkRrX
ZenxLnXJ06Cx59qYp3jKYig1KmmKYKOEVp1q5V2xvUyq2l3MyORRiD8o14/8F+CLmBOF8xd8UU/Y
ZyctmXXub2kX9A2WmcaGS7AIYbsuBTq1ATcDf+KnCvkAJA9gg2myI4bDUJ6qL62nHtLe8iMfGE+O
0yJjJLM7aPoZJWNlmPKEXUCZM6hsjYUvqlbd9PkhaBTzPuuWM2mLt0zi24TzFSqQA+SIThK2KaYc
3KLZs11+Ul0JcCCAVi87HYODl/oCqbN4qoGjJHPYTHoiyhRQgs++y4+Q7YSITuGo3P2wcmfFsSF2
RqxlBY+mM1VdJ0t/8PFLiojrMaTk1TNfmTRxt9yQCv6crqRxpgVlVHQqeTbgfgaS7NZEQHMIeZyo
GSKsVb0Jhp05UJsemus9tnSXGMTo1AH9+oQp8b99vSu+qMc81dtZrV+ugs/mAjpWMpW6d0uKmxjf
x+iEa6SjqeJrZj/9ZpLXS6ZcYxqX0N9PXVk/OidGDTnB++5t3Pw6IGI48me3JALtMYHxo5x4Ej0H
iHap+Qw45Wp0xCq4oNQGsQt6tCs9wNheNXP5I1LjBO9t6w3TKIVAkaR9bXXJsn7AKEDEAPlgAXUG
xvEeXbaOlOxlwEd8yC+dD3mG7VVnoNvq3hnzn8mNhfhH1R3p9hW3j32apsitJy0BIlhVB7Ju3Tp3
p8HRxf22oACX1jvZWu/jJvN48ZhIdpFDs0i9pHqJ0/10GXqwGmVGrQIvMXrI5FhYYmAvamldsycr
tDfJd7lPWO/qL6KlxcZ3kJ/ZdztodWwKaUDmyMxccPLj6E/JMcr+Pi0KhHOO7hVuktai0mqdRYxN
RAUNPm6C6E5xv4n/b8KxMf6MU9rSBcx8EwBzc+VRD546vD4/dEd+f3X6bNmXvXdpacrAmdhvOZtf
tApRhrWAY9449Nye6rUyMUMzn3tshWxDXJqpwTGyTsPsRmzFFlIMqcea+SeLHXKl3xZDlwYZfRdE
saiSg0B3T73KH22v/2H/hq51ZOxozmXJa/ibins1SnN87ZSVM5fid3RlPKrapv+hTye4qV70BtKI
HfRnvbV7s1zNxs5kt9teJvtYJ9oA5bIPXncjYYitTtm5GJDKnm8JY6e/rGqCLBXuXL0uv0tohIls
eaelRgLCTzFtl/KLPmBT0mtBrC0ip8KnulWZ9CotiqphzGl4E1T7xYRX2CxIU3sbTh2M1ApibKbf
6IC+pugWg8skGvafOX+WpTlcdwx1kzuoX0RCS9YZFRWZjyfUWsWZMwtuE1mlqrolvCDWwHW3AirJ
e4kH1afpCZs1+rBCvjNkc899nVYxfz2a72fY2jagQmid9Mp7f3/uKL36fLkGYmn9zVovbS2T5pcP
IzoTzK8fLaWBQ3CoqpSl59AUYX+Uv3hoKfW4U3bmQ7LMVc2fXutREK0ZhmVU2tZMO+yzL7lKold9
f9Nm9GIUB+2x3gfAmmZMyBxcQcNTGXrPn8w40tZTYRZ/PPxQJ4v0bGKmPbo9F+P9TYDWVZ66mtOv
//k/A94H3rOFDm1abPv0G65r0wWjBAfn+CvvxCIwuhil/p16JJsCoGtvy1quPuOKFd3YKB1o43Jx
iaCz0RVO6HAR0DC3JwcnBd9ZQ9wCSPtlbMhWiYegTXKkUpY+alCoHecnQVgGoq837fc6mQnEERi2
S42o+WybSRfimFeyarjILZBuc44jiQtWsY/8j7e8Np76LGaebvPOiDHlycPN/qX/Y1VKeWAGhHl+
MI6Na28gJeSHa9eevL/V3MkVrztAKiPuajLVeYIrdEkfi1nTxOVV3DRBwEQIjdXetD0RWg8FejVv
GNsUIWWIym9QH4kzFs4GAY9p96zo1YN0F7v27nLawJN1JNS6juWLUNNBpmAa+j99kGCElFtztNOa
FcEuW6xTR/HNeQpMEe8lxEFohD4OAvLMEp5lw6Pn8Gw4LsvxNZse5UWH5BxqiN1gOsWm+92tQ3kv
f4Mip59hacTsAO4Xb4g8bdk3o7zNCVD9c0PPcgXAsky0vLMtdDaLH1ZfoaylP3D1VtFiXXcVQUlG
IFOJArLjGl0UQmWC1gjcyJQIxeGtbebb+8EVPkXVLoO6EfBCbRgXNaqBX3wbKk2Afr66ZET66mzy
2/kwQPZulrd8g5D+RZUqrrKFA0//jH7H1qvyAa+mBpIdV1eZ+d9kbtR7AdEfg4H9jViMKS9dziwf
Pmtp3g2DqB6sPX+EhG3z+HHMY3vE4THec+ojscA/inNFoZkou94jad0MKgrOFRSVUqPtAPqITwxd
LW14UxP1pnzOmhfyLvA10v67vaYDrhtp3gLfGV9qt6LGoEohpg1g+dzbmF3ABVNaVXt60eFivyG4
CAakXCU0YTmosunmDp+1lRErcQHeHBQ11fxpHvPBUs8amV9Nvn4sQppsEs0sZxMswFVXa0qjLJHk
K5WajyeeNt3aBM9ledlYGRn/gbCexbl7IsTHryOpL1QclTjZ9wGlaVAJlAsVyPBs5EKYMETRoZ4D
G/sigbFfjH4xKjAaB0ch8c1PSpIPhI6bz4IDi3tJiDXVflGXlyI+2yUplkkuXC0F9CIgUJXgL5b/
6OWS3NxG+rzbbu/0uG5T687r/EObdE/De9XlyFELoVbhjFSpwbIBHuLkQtUZGqcjfzUHNGU2OE2i
MsIGhshP/EW8+NDlVc5+ERg/aAF9rMEqmUy/PMOjaZ7YSg2XNMgAhm4ZcnIT6crkAExzLKOn8Sbs
va1ZaH94Y1TWLjBNTq7UHWjg+WVqiuLf1zgZfECG9JaEgaqLHaMYBdhh2n+qo0zDW+jSARAP8Kkl
QQ5ursEptXTSCw8pMYTwi6/x9umwtYpnsM8fPih/ilrrBE0TesxUgHHIXoNlV97XjfIYe/PUoxP/
cerhUliOccAemZTZl4u9FEZWMytqok6tOuEVPiZ2/urRPjcY1uZeeaKYz5Niuq8RQ6lVzUk3lZRT
C15bStfq80p7ieW4kGbq9YxjyeJZAjjmpinHpe+ITOm3Q7Zc+LfdvnpQzJIiCwvoQHHKtxVbQr4O
Rb8fs+ytfprLSwZv8aySuAZprI6kWQIaAZbvF3L9p7nphqUtDyCgHMToGxDh3Q0a1VDfq6StYHvE
FZgCXvMV3NnV9TCEcJDCuAhLNrPx9D5HRsr9aS9XV8CU10IffSbViy0kHEU6t2aUedecBr7lHFID
NHWmxDGk4KfNLdWmwcTI3i6YPfZV7X8Sc+8/EZKiXSeIXZfEni9wbbWZuPjCm/lnAaX19AL0tVoF
7/mgXZwKX/i09uo86tBfPs4Y++GU6uU68LQqbk4grBw9IWJH2lQsdlZCxFNyrTymDQTlr1M5DQgy
BAIIsb05n+tW6mxZ0Wbclm5i2R5FjTWkMSyW3EM9f8nAaogIftVX7rI0jlOR0AzBChLzt5Ri6S8L
33QPyJq2tKLzSXPpLQgD0YjYDv5VeQTlaUqCTiubma0n53tCzIweL8VGjFUtXUrw+an7g2mXlgNO
ebwTd776W2uam66DSeahFaGOBZZHVkSBD6zQiqV0NPFtl/foszwh9gHVJgDNtoJF59r0AjtWJNz8
9K5PTB3At+shHcPokto2KsSzXIEtuPT9BaA7P41LnoITn2MRzJ+StnR1gThKuG+b7rXOLIx2R+TG
ZUNvBoDAkSi/y3Y0kI3gK6xH2Z7NCcEaTEqrq2qmRDK39FCEp40RLNS4Virq+rsHUdcsYiIVGEwa
Z8HJMibu78G7+BHYX1l1I5VwT9ZNGxcPeSZaWv6mQ9HILPgGj+A5htRcodSWY2ieCL7j9HMzGo+5
DfCayl5/dgIzn0qhnxsxxBi8F11KwXhZYlOGcwew3sRLJB7+sCTcOwlwwiweBiKGElEtXKNmXN65
ymQmBG/Bp1uMyGLhp6EQSC72s2GbklL0+IFmaupbbWjR8g2ivtMNNesj/j7n++MiMnd6c4E251YI
izhUMj8RoEBVLp1+90qlSqPhtPqZKrZBU8uyUjlIqKGAtDdGQM0MoLENtiXro4IY5VC06vbBNk3E
fJMoMICo5EbVTjg92f2VvuIcck6MES1Xo3aSdCes/JG774n5bXPnsasV74kjSSW/xQ3lVBJjAUDL
ByvctxkEh1TNd+zDtH4kWVuVgw09Z8etNMu5rmRhalI6+AGpl/FmH3iNdDhckKePRxpRTzXPnXeS
aWN4dm9zH6qqCF7yxSrC8m+nxNA/LF9/lxlUlpjeFcKDnzFCyDRsZE0+2rXucHc9BKN606h23gGp
x/1qFL4Bd5IjKzZXwv6kTPkRs3pEQW0rzRqfS1R8XyYS1Xi5elViz17BLgLDXkHavqSRi8vB1gFA
FUsM7YE6omkahe3lJuZ9sd7jcj925syNRiJuo3p9Ujdk91nLfAgdR+Z/s3V2Z3lKC3HMbYXSC/ya
z7MT+mVlDMMd6Xc0IW/ZvJpBRE1IEzkhKUhbD7YqqU4g4MxlbQhQLQjhvSj0TW3AUK7sIwx3eDo7
m4NXWFsfkUCQkDen+bokvurd8yqK/7dLuprKcNkQsh87FCMDOabw2Vf+P4oSqn/QlMDyV1ij7xjz
nsooglk3ZVf2f35n15qdkMnnwDnaZgNUvqK1Nw5cgG3Q6Xiu/tVg6flyObCVsoOyZQmhp4fNDJrI
njUwp5XvtVjck3AYREFH06BA0cG4MfsaXp7naHoonlys4wO81/IL6hEI/0WTnc088fVkiYPLjH+/
UfSCSq035Qnvacr1rDkrT3nQdtkCDHnzFzwXVphlXtlppoLMAMP7bGsnzYcdByua1Ksogx69+x9+
a666eBwGsy1nzRRhcyV/tpEUY8JNlxVl09rfxqFpA+FctAVFRU+ByQbMb/YWXc2EwiNjJo48CP0R
OSIHZuMp9O/o3qyMLwzE5Cl4IrysRFQX7be4f5WriLGNHRTc2PALlDUDYTzTNKjVs53aldbHDVkW
rkIosnFtr9Qbrtw0zk5oB1jiUpIsQ50KKfBSLevn+sQnMirFnvxMZU2rEFpogHW9lM8K77lMUFHl
CuD+kFeEEhOepkhTZY5/zZdK7J+ki57+iofKzZsRVoI/k7iIMZ+/ruvLpknPP8ykezV7CwDX7h9U
bZR7fsDGT2Ttn0OkLuHWFsRwW1dpUSvTkp6avWFFimLxSfQBwsina7rIllUnSENEdkDrEdHJJhMX
79p+Enm3vT+QoeLBsy39dTUort+/xYnd4DAJbw6Okb5ClLO3TvsvkpJYRkRCDuTmMP7LKBFDWmMM
L8W4dRuSHRszSl9YjaxkFjFxFuhe60dQVBuDWgTBMi92vfihcWtcPadTODBqPVts85/FVUmtF3ko
OA6Wm+mWGgpYPK127WFgWxMx+es965zTYzTCWKkg2vEC1et4fiOdvkaenStm+It2NAY368YV2zWa
1GbSAYw49gCTU6Izsh7mdyLZYUWM2G4SvoQHR+QRnw3ZRZsxzzDXKLx7Tp4PaucdjLnfmbL+XG3K
rJ948qnxpSS0dGJtQ9GEjlTH49oO+oYzg4ZXuN4IoRjuX18UO1/i0ItZHBAKGoQO0xCE//gAD36u
r67tCbSTjdPmOldbHurmITpswCfjpYZN+ul/Qmpk/IjHhV6P2UQmsRgNnTBXS0YTj7O5x4PNjYfv
/YBdfc3DT98gj7OlZvLNrhWrSheP1KE2T+tyPLb0Jtk0ZAH0yApa0RvHbrrBNDQORZRudBr0Zfli
yku/R2b0lWzdE9eqmRLDIqGO3gp/8q2ArCAPjmxPjwAaZIGohtdP9PGowsdHDF2bELLJUvVkd5uU
v8M8xgZYs9/6faRhpSzDbYUp2KzjbDqjUmTQc8Nd/4dQHzI6s+b8jJW798YmUYdU5+EFoH9rjR53
PU3YZZSJ8Je52xZxHbAAsSk6WmVtyyd/nSVZdAU/33HbVAtYkbv5oBg9U6O3wBp/1FIOZxzAS7HB
x2J9JxQEyPZKCpDgR9i4Q7Ke/IDKBuxGXA3/bVA/UsDxUieT54nSAS02oxLveUa/Ie5d/v8/Gtiu
KEa42OdW/EKAEefJ2ogvmeCPVlFZrzTXNTdGT/mxJ/ieA9c9xc1qOceyAUmND5wRLAubG8uc2Rqh
BUfIbYW2hLRbJ5jp/QZCB7BAfvuGSVM3W/3htfBYpheXYULOlYhsdPsgvgGEBSjn1X8xd0nvto7P
zotRaadBWTa3UBjFCqSaspI29T+PwavrtCuDzZ3ZQI3h94SprN7pBJrLONaxWkWBHTn72Y3b720k
tE3u62ZV4/rMp5G7qyyjmg0cR7oX2/90xojtkA9QrFYm3W4pRAGFvcBn6i9WPtdrxySjKJI+cDYp
Wi6QmGsniapu1PYx6B46ALcEo6pPBk/EM1o2fVZXA12FhUd2l8r8GeQ4n/f8aa7XfyKLT11Uvz0w
X75F13faW4yMI3EHybjZSSgmT9qRTdTyGWVmq9EEAc1CReBCtjM69hWzj4JXxEgP94xg7e0uTeAD
llNXL2DNIJgBZtmrMcoHMzlSJLGBD03nJ7BXfVqgplJt/c0MOv6V3FjRbABchJdhHCCBI0XLOqk9
zmrzbh6gVWnxBuoIT9pqPmgBNDhAB1YId9LBroFa1Fs9qDeCuuMXs9+XktDS3kHzSgGM7IscCKRj
GvOotctFKvebdkZPSs7bxkwLHfC/g1i8TRNPab5Tjgv69SWXejRgCulePMhL1wKm+b+2+o7DV7os
U88Hh1T+j7zMAf/ddPH3liBxslRbgXW9KDeeyEetwjuysLaM7Cd6ANLSz+02Dv78aCjVfBQr6nPF
IX+j/TqbtiNpr3xxnGjR6o8tjLU+Ey3oY7FJqqiYegfixyKWHhkDvXs5o9Wu9+Jv3Rchh5bRtDjU
ikHH3r6CIrI1ioI1A03zSDCXEjkJKMlYu1n1GxiQfLKx9HREC8rcClHy2cJJjrfN7Nhdx2jf0pKz
zKDm0OA9eKTVoELjj3fmF4tfcpZMJzHR+fOwTFA39IzvSzXfsfLrwTAKyAUvlc+Gf9L4ibjU1IdP
F6NlFWIEbycvvfB4VsVJY2HlDSVPmJ7GzVxl80G2kEUuby6SF32CqoU45tHRUlC9kaWjn/X5xY+3
9YcIXNWTfMmpqxnI1KBApq8xLKEaUMmxA9nm6Z9aYTsPZrItYtjyLgYjgtJzBlaFYNCo7yjBoIbP
DadasIzJHHXD1vXB3AOXCkMlf2mZrMtDiLIpOOV8LMZnO/oQdk3aqLjRHUFH2x5s57nlYf3bZycb
t95d/l/JiuXjl+MUhi9xfefRJ3YtkxSCNgDihqF/3BOKihp8j0jXz1ggIcQlw0oaLEulhF9m+74q
CVaDd/ePS1fajo9rc0h7XAbHBw3uOAqmYxCd3hT8jHsLqHCxkMC8fhOWgEt2t6+sdt89FVcToEZo
CfYI5IxeJw+8/Rj/h8rOBMeRzr7rWwlPSgpTPOBFkfw1McSVKomUR/anXq5ld/kGrAkJzKM+I4BL
FTKQJa5XwXUMV0e13BjfMpdEVAptfyyw2+T4ko4fE37IWnwNTj4Vgp7arjzGL1oAXz+LK5ShnGzC
75sRhoU9fz9lcMNyAMr+yIogldgt51HNSLQ1txQneYhnJTt8YB3mNQWF5BYGvV/aRT6pZ5N2D6VL
bQNij0grBrMqfV5lzV4WfjFicszZLabXUtF72Zz7/eAS1GRbmc4e8a3VwaW6ET/hCOcVGOm/x9aJ
GYEVFhjDZ1jN/0ONQkvdq+qdirQok2RDghhxm7qA1yIttmRUXoncZsNOz7/nDSiS+XWPSTVMg6Qz
MRN8TQj6iQNQhsNi+72ezVReGPPF6acHioNjKknAfuxWDbcZeJeYtaYeXVRWx6FXxzDble+YukPp
PcSKk7Uaui//Cw1X4GfQ/9CsK+Ve4HGO96bPiOcBXCm+Ozz3OIpvSxUk0LRHISgMFySpKdA9Krqh
bhNdO2LYjVezV6zvB4hv1X7pr093y2nM0a93s7nnQI5yICYm0tEXXaKb7tvWr9raCpCoeKr3B/DQ
iAI2H03NYJp/l+tpD8qEbedZ+hRJ8gj1DSrwZ3G/aqUy2UUDyA8yDmMPrKX+TUgthWmEKhsfb1B/
KtWApDcN9qzQHz4YDr1yILfTo00chxgguzMx074RJ+DZ+KOUXyodYjMfemPszll1wRovVljr6xWG
BsxEhIUCzUmZ/YFSlWD6s7z4rgxNE4WEfRa8PqAdDdDAKdPpEYXoAA5MUKmD6jYFB3K94SHBHl6j
8YnVK/jqbGt9AF9LmYNR004wZ9a85S/ggcLN1dz8AqxnzFivPjcwBuDMLn8BdBBxv/kOtmmdK6AE
BOCSY6R49/19h3vv536D901QGs5YNRhupo8TH4Pv9Ne+ep2lN2cUDAdjd8zii5w7a/Sbib4ryiti
hWwSAvyDL4kcHy0ifi6AsASaXJd3xSoZaZc5/55Ifa4TxGWe4Xv10YGusbEcjSImo/yEKOPcJ9LD
4kd+wnhqSRVUgbDxeIQUhcMviVufz0LBKQw91bA8e03oTK8kMB3j286Hu8uzQ1oadnSD48ngzpOK
PjDpzcG4nmlJu0qUn7cxi5BKTILn500HeucNgaroZMk7ZqlKxEC7C6CAHWwa0a+GVUocmLYihMn9
imco76TbMyVZDFwUTyQ4CCjYDPnDxAr2kIIq1h0D/a4kVGGemqRBw0GP0G8/o6D/gOL7gPBzKa1F
pnXqHebLQFPLMae2Eg39ZjQGrxRD+miW28cRRfsHr1vfB6J5O2hdVoY2zTiomWxWD5lrkPe97krK
MQ2l0X3cmLKZoJVtMb5bdmJ19Qva2d8bgeU1FJuXQaAQWpTtwpAYelPDaZDZ7ajB9B0wcjeUlDZr
lhbx7fd/DUrsjtaafNngIqyzYoMB6xySRb5LCTQ4VR7KJwBrtMU2QhM2UFUARCf+85uIw1WfOjWy
LDbLq/bB9iH5gzgnFdISnh6M4mytHcR+fJLDhcP2VCfxyuroasExjrXZySzwGmqPlyNfQ06cvXH0
zfTFj27H4nmPYAC6EroFRXp+jjJi3PIgyqi2MMw4dUKK21GxcHsS4nq+I/SAx2xduoRFmmZYVQ1+
waQPbvrgSQrIG1NPhFjYR2ZV2DdiYvfXEz35sRgVAlG0BvnKvbuCotGGtbXeOyz4Vs2ZZIGNTv7L
O5hUa8VAWvVJq2G+qH5px9b25H3jcm1m24Gew+I6HrrPeQz0AbFq2vsC+gAvF7I3Pv9MaEgY423T
ozx+U+fiEoU0PbNM7/7I+y1wwF5nhqaN666Z66QhnngYaDGligus4+XsemAUOh68tI7hbYJWBBti
+Og4Du3BJB1U0/Gc+2v8mcfivsCwbO0k997w7Arq1QkZNYI/8XRQ8ws5VnuP5Pp/8tksU2ewJKpR
Ne4YcdoM4q5fWIKFMrvKY3fc9SXX6Qj9kP2Yei5xglZ4eKbeZMgIGEettxRVfluTAFHpmbly35rh
ZeBsLV+TdndFECo8K/IAkZLF5ZtMpf7paIg+uwumrwqowdxMX5/y2Bezffl6LBHNCIiJ7RcBpjkS
Sqo6PLZrY0rbPn0ZPLyIyGpdK6VGDKTlrMtpvzR/Pa+EFdIzTOVuxo1g8tfUAULGWhLTytw5+qcp
62pYFJyuL85TJ/aqMgMqm1AaJsSBL1z2qDFTOTbk41W2gsSrALQoJ4eTMx0IaM/89lB1a4JT6Ra/
jsWOIFrs1Z6POLjJyfdjGTA1+mty3aa/1a2cc2p26l+CK160k208IU2fLKeiVCiXXlA+sLKXqXr1
X43eG8fGnombJ01sjNP5TOdFPQfSAYD4Xm6IkLWcRjS2pONhsrhTXDneAw7b5oVj4jgXe3/BNFgs
jR+n+mOXdA8PUqbcnR8JJvAyta/G+Y4XI0NIp/P9JTdE+gBpeo9dYowrTfgKDKpap8sfJzHuuVnD
aztUafk4kTMyCge3jpFXN+ye4/irkpfErKjx/gvs7XkcKUZoyngyzDv4H8L4MHUvvdXwb1URE6Cr
34dKxx7vKMDUAbv5rwOZqvinbkWSL1VXttG+CieWVa0j14mlpqjC30CwWZWOiE8Ztefncsc+2bVX
o2E1dCcf2PJ8fsaVGp3vYNu5FUw4uwuSCppducZLIIzFmaXMkOV8ZS5kNmGDd32+ZqeveWc7+ZbM
DKKqa4Wpdg9nA6bY+OXPb8EGGdvGw6cKzumtY61En7AuiFgWVcUDMZ5QtziuXFR6cw1o9myOi7OD
CRzIyUWpRPMpkO/sMUVtdQ1MWul6PkwQZT19s5wXQNBqIlWp7SYRtbnzvohwUNgIBeMi0lrTd/MC
YzFrpjIhPkeyReMVc0y/oznz65OMcCdTOsvzD7imFEUGofTq2cRLLkV2yWznnkN05yILvTGsiEfv
rMwPVj5EcpQ/rxvhnEihq4vXo1m9L2sLwPzv2u1e/JwrpqgOw+3pXXy7OD2TiNRUud+V3wXcq1Yb
dZ5xr2BtSMXaxBrexD6d54UgRfWXW9qhv8vyurAFtLyNfE97pMQ3oxpDhmdLe+0YRMkcLD4NM9Th
vroYnmQyao4Qo3iRX8vbHqI2UDE2k4r4UoXRwWtoenDPf+acnUqGPlIhHWFj6kcKwqwWYoDDrnTz
VS0WwoeNhagXW1kIK9uSzeDfM+WdFcauaKNqFTEeR/OTEEHceN+VSZxEB8kd9KjXyDD5wifeiGKO
1i5vfqZ6vz66tJUp9XcKbOMu520rE82edQLnQA8+KxdYMrusTewwLeKRvzBupzaNdvFouPzdRVcp
IgxLB+RobDjKzArvHR0B0z6V46oaoaoUxtsxxJ+oAdAV2LTGYHKUebCDH/zrr50wlAxgH4OUULRP
wt9DdVbSJvsab/B3mhNotZifng4TP5I2CIN9jX86Z6aNaZ8FeddZE0AA38KMlZNCgG8CktNAW8Xz
uy2X2B0e0jxpmCtYxXt31TL5cPKrenjkb4/gyrE0RbXuGZWT99C/NuGChO0mdf8enL36uvZufHqS
xSKmHeQVYAEul10tsiLgq5TeG+AwBgpQJpXG98PzZd77P/1xGBJNDH6UN/NpqmdEImi42FRPy4PR
So5qatCb0bSTR/gnFWZC14a5jI8JXqXJCdshqRGPivrpQGWujmfWYFiwhVVeukMmmz/jl10QtGXx
vDLb0B+RYdRhpv7KP8HwNCVzPfyLsBToYbTC/atw6nwYDdIwYZY4qe2maLZasQfgLuEcq4ZplIFZ
oaxAENzmayKGgVOHP6GAtcrTRQ0g5Ta2kh403mqzkryHCvFgsJW5YHP4O7CWWdD8qeDRzT64R/fT
Cawgi7ECpXnAjm1+azVU6Y1v3m+4OuuET4+gx7szYnfoTNQVvlOBNjZzaik3oQQtbfwrS+iq2YgG
TMhLxy6dfiFQzBsC1+J5MnOzzg5CpMHFC3iOMfkaYsambJopWL7M+aY0OHT55CLg4k+ZPhrboiq2
WZ3rtAUzxFQuoCYzzRUJ/XqFChWXFiHrgZlFkJbugfNYh4804PKftEDjs1hiTkmDe+Lz4ZnrTsHp
OdV8TjWuRu181tApxj1y4SCKo6JYBWb3mYn+yqB06wt3qNU+GK7/GOUYTbfcVajT+14aQud/ryzY
8UWjpcxzm7S0EUd/2ClGqn2UV4pMlZ4gFR1Ac35/SBYu8djX9MbOuTSeTUeVA+DVYP9UBjz7FHgx
tq4QagtaQslErmjI4z7t3vFfCPA+Q+ZT07Vvy2oNPqGHesLgDe+B6HKwLnoxvbPl95galwgaBQf/
Srs+UqLhdu2YUeMuIWZlZNQaKBCOk4jt4nucXpBMEAsM0kSsBnJ9CIUwmLiwhLonGYpqSBbPidNb
LcWprvHcdrltT35qJK27kS4LU5JJyVLVWpblxIQCuDXxnzYO/tpCbVtRFOPbwqiC9T20I22i3AZx
6yjn7kODez7vJXEHAUGt6mmpSpgy7bhDA0+lSrSFBIeQ3QGMKiIfaoJ+DK99Vlgon8JfH1VsLBXm
18yn+UKRYnlRrci1x+vynYhBisnz2yBjWXsK9YleiqWftCxY11/uSkb/o9inNtx97bJKu7tnr38A
0F7+CvRWuVuac0readq6D1geayR7EpCU7TZOqIcPZi0xkXlF7nSpXGMSSWcKo15HwFUdLkzgdMDH
2BbstOo9umi8gzkgSjIG/IWhOItEXRjdxwqaqTHOjdV9f/M8LuuwZH5yHlhlNAXLwvLgn4KNnwps
dJUy9mKrvgUXwaMbs+xSmfHNTBDbCRx/DayJzyqIgySMrJnN1yUj8Q3LXeqcNJ5lj/Kxqwux1ta+
DxwjcCkxICB16K1SQLfqKXs43cyArpYGboR3e87EQ9/FoFfuK09Mrgl9dQUSviDpiU/ySHfNQ+d3
ht4dxBuGHz5m2Yj3C1H1WKE5X8WgvkFcDbCIy3uVLQzkHyjnBAFtxU1evhB+hw6JT5Tu9zETWT6n
Ti1Y9Gkgx8sADoiwKamOE2KRo8LweIYNpUtuy1RuxA/ayhJE1aCp+6YRY3dSob4jc1AFNaOkVOBW
Z8PA8V47o3lifDzEg30vN3ODIR7NBS5V4owXdqws5AdCLvPfuZ+ukDO2eVOwlCZ+dr+nCWBMZfIz
VWlFOczoM6Bq9QI60JVfg1u4O360PsnZnWkPc5HIZvnzyZIQq8XjrHJZHEDJKefCqXcFBFl/wBir
jp3hryLymtsnhsl1C9Uva1LjKg8rReU7DAPlUc7Yn3sYmp7a3dRqZj55M7BeUCvQBYPU15olOmtB
0803H14ObXoT2Y99pRySiFCWB/He4qVaTzy6M+TCRnV9tN/Tl5zfnj2+1lPwkDmmRlHyNPfIeaAe
OIGxdzouQF7Rv060zSSXlQ0EAO8AJ7reGKZCgbpp7YhN3tRUAdl4hp8wk42YH93bZSKG+gZFYx0c
WgrSyMpyXyxnnm14G49ecfhG63ojmQtCUqwzOQk7i33t3qTMcvK7lTetFxDe0NsQ9XfdN1tlHDY6
D3DLH4LIrVNE4hexEO3MFKB6T9aG3vVqgvfJGkLj6BI+YlTtSCkrfdn3G+2tIbgPrrJ6LFlVwiqp
9b0mTbN+PQQu35/NEX+RjvKxouE+5z2usCIfdUDMm8Emj/R86wH1MGajksP9u9o7gdpWSOk7S5Fx
FWpowX7zvkLWqOY7wq2kiChFADB+4yrNHazYdjA6g/KK0amitWweuCT6KcP2LXxZdCA/rpnZIQIS
2Mi7/QmFOz3iT44s5PP0Dz7x+g5D9+YmM99KgG7rTLExPk022EwUymEAL7OeO/kr6lQMLFzVWq6h
4jRE5+3JQ2j1b5TUSArcdabJWmUgcMFn92tnF33WKOlurtlIIrk82lYf7uPRrRI2b9b5SvzUlu3n
3+Ywt6a1/NoARb7JkvQuCFDt8n+BsaYqc9S/RTq0kRa1PaNQQ8e77fUqRPDoEWXuDdLea8RuQF9D
X4eyM6umN1aOKwdY1TVZGYhAQ3xcNthp/oUNV6CHVJFEKHQW1HanADpcCHuCvUNf1bW04WUfMz17
Jv5ZlqIt+fwayW/aPaoN8tJcn8yBjkzas32Uo4K8XwCvL05CUDij10QN1NeMyuM89GpfxEhi1EWy
/4ThvAn37PLaLDGQMqE4a4XUphA09evBYntZKWeGIH3JkYEd/lfuuZzQndSzzQQYguTh8CMNZc6X
ZrQalkDuKB2+b5Hg/DP2HqsNrGQffYcRBbbcNgogiRL6xqjU877Tekd4PHZhTI2r7Aul0gnPpmyg
dvLdLtUUMpxDQqtqIunrl4q3lCjwFItDbjzlt8J/zzbz9ATbh0pp6kWSBaDwjySxmqWJwkx3GYnO
jwivCcTYxFTKMVjQbR+AnANfhGk4J4nXxB+Z3QA0TRDGf9SlFy0a+P49xnRKzyy3XiXCAHTm9+Eb
vv7p/sWeZrRPK+jX+d6jokLrpXpWCeyhqyE8X5Mgw4gmVwYhwpOIawzrlp2zaEU/7GfNa3IxQnVe
WCvo8beNZShWaQmY1JwRXQ+LsGfZHcIKOFPmpyTRlNbXauQFlhPVfTCTLt94QBdjVzzGaadcPJ0J
/pODGHsMUQjNH8xcrwq+OJAlnLn1Y1bgILEwzX/R3CnrzkRHJjTtnbgJAMh4M7sfY86CBQZcw2My
e/wJt8Zbz1zW68mmw0K+rvqdA3nbRhLQFpIdAjXEfOyKM3mTe33E896A//SiFpxkSWzL6cmDYJj7
mSpa2i9tfCyIDT3QSnFX9xdmDb1g/o/OUFMFeU3CB07IPP7IMkWolthfOojY0M3v/y6rh89qouOZ
C4Ah9uN3HA4huezkbHUuJLvocz4OZN7p883tVICgParnTX+GkVyPmI2Ok83VccG1XoZ3urIUGLmN
UfWqzN+v8Khh+IZYkuEOS1cZyU6EfgnaxP+/wWMOdHkG5+ym5M2rXs/wrdBSEOPeiIa0MqDxtcSh
VmJiiyfIL4ANpfLijQb9fx1WIuzZBfod1IpdFa1UlDeLtOMU9zKkF33lioc/d5GvfgBYPqg5z2iF
Bj9G0iXEEKJzAH6evXejG9pUB2LUui0sdZPvnM55zBo0dqSUPLg6/gniDkkT98+mCqHSFpXeSCj8
Wo2Yw2Uvv+gYtI5gHF5cEnhehR/r8Sr10jdPwoEB0ShNakpgI/vAXrS0fQPO0mt1o/txp3P7X+rS
Hq6I6dYVrc40pQAMuxHNo5C+vsvq70LCO9VN8Gwm6Cvw6hEQCBtBKYdeguBmDSPG+nXauvzbW/o7
OwfMd6meKk9rrnY596TSLrRHL8f7A8i6qq+cYFPvX+pEXPhyvOreXouqnjIz4/Jm7rXXDZUZuD1J
JpOKWkJlOngOJwvB9mXNhgA1Dy9OYEaCmmdW5eWJZUfGHzcgjtFPxbI/rmdiiJYoV05pqhCJaprv
5zrY/JXcVPy1nkrCQpnJ87k/zB/jsEOAIqagA0n+lFBGEJss1K++vkIlfAKei/qYhGrYOE65lt6m
R6GrDKFbp8dcLXvx2ief9g+5tW149ZGlpdOa3cBAsGxFzwn8MP510kRcO1DmGkYhqdA7Yn+1iIJx
C6NUvjHqOE9y5h5yZdpZqHEf8LY5TesDgiAr48ciChw8/ktM5fNyAIohkMus4iIAGPA82uZE1Jod
90yYwQhX6XyNwiovDB9f4vxheFEe+ndb2rlQRWQWKlUd/21e0KNjLW9JrX5qkZr53qnuoMQfcpAp
H4nAUR7Mksp1wLqBgoxRMyw9Hym0zGKtSLvlLiHTqGSpKirDzVcL3ViqBEuRnq8MZIpagvjQYNWI
oBNPmdpXw+uGNbBalfilVffMslxwDPHHkrbGlkHDu/zm6KQ50Yn34RVs+cKEDLSqOa4NS949L1pu
3EwAabj3ISOv1amkXTeqBWwppNSC7S0CntesTWVu8vqMuhS31P4p9fYWjIcVu0+9/LNL98NB/1nO
40FV6klV65MaNMRrCn1Ln9BC1kgMJmnKOmNBaXN8ifweOc2bVRm2pjdwa8+gM+2gnFuggUL2YBBt
QjxUB7053OQXMwkGknFfKP/uxS+5Ju2wfuaz8ecG8hb/Vm5Y1Zd0a6DThMZRzG+mA5FCO4nH4a/b
Sqnw4Fbcfbzvny+JwDGM5+PnMJKMqttR/8uo9WiNCGxfNfzZwrti0A2MlGBoBmsWhcUWETYkHzJ0
mdUd4EFhWRATDktdn3nJ8dZ7SUJRrghzuP2yxdzY+6pk2doHdY0EB7bm/uhgDtm0QrIcZwwwDdrn
SqSh+OEiWuTJ+CumAWwCrMlVgwcsXvbx6mJuosrPB/4qg9f52t74QmtE7Mj922UvMaykpQEihmml
xpytGQ6Eo2j0j8HgtvA+SkK9G0Jp68WwReu6cfF79U+dUhQY/lckE90Ev81ByBUd/J7UKP3K9cUi
JshJP7q9YZxvBdjg3Pa6yt7hGFOE+HHFmLk2U0SwYwR+qETf3S876wt+/H+T56WWRw3wwST2mmQB
wgn0AbLOnVFmJZxjd6ugk6Qhag75oNvT3WSfEhbsg+aoi4ZFcVmyzBrojHC8MN12xJZ8jenot2ej
5HndLlgoKoHOQHfbkEv+RUnZ45KJb82HWsEHJCHxPDEDPbEaQBK+84KR+t2R7nT3wLSbv5k5EQ9v
lkYY1nBxqlw5hrUqJk85oUrNVzUtJwyQ1mzWudQyKxXA7RM44RznKONB2dyF5CMiqyHFQpDy7OcE
Pzo4NQeNMBVx1W1RruXEOOliO1BccuGGP4UINmaiQlyLLZWtLW2aFkvj8mRAjCl73sioXvr5xUp1
n2Q/XyMNUAAOgZkrYlFXrOG9q4f8xwaTIycbgadG5gSFRcueDW6SiucraNpzM81WW4N1rKU//m/p
Zav1ZgW4jm8+3ATjn84KBZxloRUdXQGApg2iOodUxJhfi/8wJFSK9vrM8SOaiv4i161uQX14RcFL
7Zj7prpV9aY/Ow5BljD0Chi/i4YKhYjYtPC+4kryQFySzTIO3mRZ0kipe3vvQ+X4Raxk2vHCnHSX
l6lG85RzuGc4tF0qhLFhHeuN8CvNlIxyedoO50/KNKybUI40aO/RKHZyNFGIGOZkYoAiEsS/r2Wy
fYpPIORgxOTlcg14CM3CS9/gVBtcqb9JBe2dzCgy5XZ0g5DCDXAKDkG9khcgB/mQqy9BCOhkXso0
ImS47bDczFzgHczsYDRsn0kOA4vsb/iuFZWFANMTL7mgagY4eWzwsdtTVNFnUA2nVT4EZwiZf+3k
Y2Xy0XTZWZEjTjGID68Yb2xegyEhTqsbC/Z7TuDnCD+1w+p1oBuLQ4ksIGk3VdXHnOKCk0JnHcNg
mkdRw2rlaKLK02AAvk/qoSvXdAPBCrpXUcmWDUxGp4cF6InB/Nlh2EWAPkDZ0TxDLITwwN6U7p7e
84U5s45GLHnwnwtjJvI8d6QkwyNxX1flEG1A3Bmo3CKUz2PnyUbkX20qXD0WzGsX9t1rQOTsimQd
o/PR9uH7/XAEN48+zRg+8sbP7leEviMKym11w+EbGLILDFMjZFU69ArxWG+hsjfbBQmnGMSbVjY3
/rwDgMZxyOKSKjCEfjnVHU3uWOGIN7u5j49sdd9J7huQNYHr7HtQ2Z7IqGLIIhLvJVOZW2Qn7nBC
IcZz6u/4A4IQEcIexONavlf6mkf3DweBF/0Q4vvrfBHC2UmHLEu5kI6T8mWBeUaALu7826cji1nb
QAQ//bAQiSZOm5DauViIp6LJmhe8VIQzZFBS3af5+0ZgKh1J0uC52uZp4OEsbW1+IbFSZg9SkJCd
BS7wlXxLkTw8V34C6Pk1enl9GxK+fH62BX6K1PlY2T2XHhmN/o1xytbsQ/n8rTluyHYGOjiPL61R
daP4OAuSLkZhzcFDdt92lqifefRhIItaWQu4kNNRw6zO0mN5ff4sSXC9YbPY/yu1+iYlydOC8HG7
pyULuhsauTkQcrKzs4ZldVRyRodV/FSOlp0TIhH7G6Ig6+6N8D+IEx6VxspBthBYsRqrjIAeXNey
ElSkU54JviFm37BOI/myFHmaW1eZZgMD2vTv8yd1nHCJglFWgKsPRjYFEkDERDJBYJPUf/Djyqj0
azrKVPcEW7uIsozDg6//FMXa0O9Ev9lbd1EitIKGtvHHOyH0kIKgAR8eu2dmkhdZjT5QaaDiZmd8
erQNyURnN32mDKiD9NgFrD2OEpGRRBPHChm6/JJzKPoUhwJmJhZT1VRvuoOFPLyep1XVeZMgZCc4
qgeRRqaH1GGljBk/87OBcE8KCXnZIjX+5u39P1uU1m4OIrmRuWOiE8gLUjzoRHz6PhUOmHDcjgV7
xTdscDAoETj/q3IwlDpEXhMAzC625ioWVveVp5ZjgCbbugkQ+jWIFbzQFWYSrWl4iyA/y9zplV2J
eVfDOQWVKkNugB+6jGFbdE+lgMJu0o3mbMQH09f27zz0ejk6oN6UDDbh8a9RicgsywZNmzvAQgyJ
shq1p1KLjqCqAU6HuUUHlq3iD19KSUGekL52foUzTeboVPWKtSppmML3xBy+bgc0lGJtR1831mQQ
qVgwDfLyOE2IKSupf43WT18bk0fQ/he7PACnIrXPgeJZmqpOCE004BPMH4U/T9/DFZcQSZSJNsbQ
/77TI/2lWIuAIMzP226F+iarYizAthZHQ+Knwy9ldJrG9nZjIF4kN1qhkX2FzOP8s9Y38KS8YzED
6EXsVCQErJuKLQK2yV2NUcYtb3DbBsSw1/i4wLhddKkAofRXYecJTamsCOOp1Eefrg3LaH04blLW
9OQ/F7s5oTGSO+/ZNfSRaJTSxluOc1zXeBv2lWfLZVmb7CgKP7dNeM+DfNj/4oRqux+hMbSzKMwF
yKS86HQHiEkeUMJrwYkQVtoyeLflRH22JH2r9RNGs55hM9Z+K9qEMHF9uuZFXjsg//pOxefncR3x
hGMSQ1viXFJ5n3a94QstYk4f/CNRtgxb7fUTkPkYwAIXMU/+HffC+VmpQB67yPpS/0wDlJ2/q7oK
0k6pKvyLUtf0qV4mx0KS6LmoBLB9nf+6DF789zDjmKrs9oDFAv56nGLtDUUTfXVEEwbJVDDABvou
e548pHZUwgw3LHuaX3bwQxr+HuXaBKSc3pbFta5B1QtedO+m9CsPKw4XyKSuUFMKlf7P97V7wMmW
+epqseEJ4u9iWknWRtF4kKiNZUileLNRjjXTKXGm8RuQ6Libmr9vGplRTicdWT0ADuX33GZMrQIP
duRTbS4ufDvGYXW2nB+SPIk0XH3FynSGf07J3MTGN6YHMqZq18CgzTnRSrEW1zuyxOagBKsabCfW
JkOEW1fz+TBsw7xL8IMzso63lT2mWDd3QQUryvBwSfIg6vRiG617dJ7k5B7NaRnOyuUek4HrRogv
qlSwUswD3UEc5hmmAg+BuOAzmH5Xy1c+CjD7CylxUuPQGrqTe4NCtUXBXRnZ6pjevgLqKJtqqezw
ywRVqeYMUIxXfsLAnn3Ssu8ko1dkmMyqcc26F8ZrFMQ1XWhCqQmbFg628e5ZNonJg7N1oMlwm4oe
Fpe385VGAmnX0lhUfYiBzOVmG5nYhsodvaZrx/aggC6NleNF0tIP7FAGFFlvRC848/3nYNUIvDeu
wdNgC80GmM28ftKF9InkCaBev0xhQGCaB7nc3ul16CFbOjOza6TDq2h4tbs7f8B8h4q8/7XCVHYP
hOrwl+Km2erIx8pfEfDrKthK+pDWMiLgdT7YqxHWkVmHtCAyqiWIom6GWOJYZiROg7GDk6Nc3QrD
Y+1vKJ8/lQg/v6Zfy0Z6lmsa54q5fzwBe1DTG1ewbkSu/4E4JKIOvRzbiZ/gKKIzoY9opUypln5Z
a/RU87teAVsKGM9zUfP2CPuporhME4981w/9U/tV1Y7BasiHyDQXCAnRxuH9d3EwbcIREczQAgaT
ZCb53wW9EybAlTgY0IflLcytwdr1ScJjTxAQZx4mZ24z/N4+KKLl26Mr424BxI2wnzI8zuIWiW2U
HIrf1klIq0NNPOABF2jIX7HaMnuemA3NZoCjkDH6Pl4N4A37v5jNWiaJQSfpk+/I8d4VFbEwGJTL
LYbp+/mStyg4oFo16qNWGTH29HJQE3RNNTJc4P33xx4ShtcrF5+7au4RhrKjrYCvIXnyRsoK9Hb2
u+7kJbO0/JEtMG11cRM1U9EnKbRE+lKFqh11BeJRVdNYaXIL77cMcSdLkpIDJqB6PJNfkOq4PjRM
OqODj97gTFmpkzOcpK1Y8sV9cPuyy9KN7rOhyCeusKmM2Kq5KPlJrrwYM+lKigGmCgLeiSu1d016
IYcHu7gSaS4MxhqSyWfrXjJzW153B0WClC1XDpYCXFR6VX3WRqnmkOtk86tn9U+ugMu04pKGrmyY
YnH58EHRiRXHDdyoNwuRRu3R7FFhEBX3EnW2SpGfFmOhM2+rER/1GHZvlcDOJ4EFHA+87bM8bYGH
oyYoedEbNZzdqlOqtNwVPuGKCaCm3626cXsvogNHqEf9r0ehXJUuEZroXDctc9qIj0YM6elhqgqZ
IHiU3ycFXJK29QlC+o9wq2kw3gYte75IC8tlJYVX+U8j/BaN9hCdjtDRiDwMNsbnby+3+qEAJnGX
bYNIKATLGpizuHQ2+SPq/sScmRa3LnSFxqJh83Ek2Twe9CxP3m8wf14eX5qmxVDVvZdCmrPhPUmY
+T0vIDyHL3C/zC/qW7uPmSZSVMMzy62cC2Da3BkHG6XFn9Yg+3rUEx1FFZw07v+LZRYkdr2765+f
FB90oSYLdpLcCppXZ31rhiWqmCS9CUwODSZyg8VOd+p659KlPpYYrpu5RekcUl1RvmvJBET8upZD
9b5WiyRHTHyQS3GO8AQmCgWplqJp/1GMvunA5NFqmvV3SiLLpVFqKKcEKuxoYVCvxuf9UnQN11cE
jQAaBoi1+zzzaQ+xRWDAHIxKgefTO/1ogBtWUjztuib/sFKHyTOj7U61XdSyROoUfr6FXhQwyDys
Nh3ZOxoDnR6kxc/XQF39x61ClQarsBc3hhU02F7mdvFE+KJ1WG8eXP6JnjBm/0C3Tk5qPLsD2n/J
mot6z66oaDa3Vc5vzcNweZfVRRqC+Sof3qPuJs+83M4xNnHYjLLS+QyW7qc1rav4N07iLz89ldUB
oSG7F/ABbXSQN8JX2XDBXJ1AKXBLWt1e3XRmctm5YTERSWnXWnXypALCJnImQhPY4mF+BHMTtu73
HLE0wMR4F5NdjLDDUiIfiODbzuCG/0Q8eEhrHr/6CNsCBmM6BZDCArqHD/HcQH1wl6fJQbD/aGsJ
SC4CsUJ7AsZAebtwxR3yYM9Fv34hjbXfZHRnn8X1CxnNT3KZvgfU35hDncgRA/NerfB4dg4pqThP
5pG+c4uGUBa5FgcWSSsPaBqOoPdnFp1YeR5FTTSpHABJoYSVLDiJKp1OhnWPMyk5yzbYntkRA9HN
qlCYlrYoSx8M3W+ssvG1U8kf76CtlrdEi5d3bzBBckMgS7ugjW2TgjZJjuueixb+kc6eZFD65afT
o1nNq9cwIdYBTgvi/YVU5GBB12mMRD7kptKkuLhqaW4H20Gn4dLoEk41fFwTg1hTtLbKY69KIgXW
e2NLdbSegsbuzBIexfSFYqJv4CjyrDCAGW/Y6xyNLg3qqQkkiDP/Bo6h7ZHePlYmzNNMhGjzAg1q
/bo9mtWAy+BdMaCavjmresldmaU3F2iKbbemH/B/QxFLeBXBCOln2WbyrxQPt9j0ezOs2HLOz1dL
bpWPGjrDhvV/GhhNPjjcCkZf5o8hLiLKsv+N/QTYsil2NaGgfJNBnNa1hTObrvhUw+MM3lA/4XJN
OXxO7EkOBg4caEiXTx3PF0/p3oZrI/N7FZsg95kJtvEQxeCgtiPfMgvnSw8J4V9mvQ8ImjxTy63H
P3J/+rHX3r+VBEz8lPxBDflDTJoPtDFD3cFKwxKzkveNeQYTc6XS2bfLZ+zh8qty6WbnXur7wy1T
fnyF1HGcKdMb22W0xm6AyzFlL8oAy/ROJfxyHej7Evg5Dv5HsFjRQam4Su1WXBxSMFMRwGb6IUfI
VihEkbk2/SwonkcMExebAtxsyFkdIMY/GHnKNlzMzGxFBSj/JEz1tIQ5uvwcdWMgha80WNU0/rvF
6YtFv2jt6XplHR/Zd2vm8zGXsBVE2OxMofQAq+YDZa8/pTo6sFbtxVlIFA8e9b3PIXBu9bF2LwW4
hR69rYatR66mKHo6eZta7OnYd8GCwpuUvrxemBNGS4Dqgwu4eyod9eAIxFJAyaxOjXyNKOUGFJdP
XYcBv6N2lLTcHqeVy0NnwY+JlbuZWj86nMGkPrH1PGSrCDG81nnHIfIs3n4RgV+0MsoewT4HxGG8
FXhHJkR8K1YPRTzi9n93akTU5LKiI92wEdjy8J1GVXaTM4/mdq0q66brX7NPBl7ZUXKL1knXsED/
RxVl9+lHeLI3k9lro9VO+BopaXMrxvZL1d3hBy2a5aS//p9VUVmbfC0CmZYRg3WGmWU9GSlkl8bx
OuYfuA7s8akiLvfN6DLMI1Bg74QH6dEBerJszbBA8IkLFYRFDLtZwDuQmJA6rIciGAdgGVSFTxol
skkxnGmDaxMmaC7fwXrpoTt/r2JIPQySpS59TNjjT76emgZiN3A+oMqP9cGesgX4EyEswHMUaLVP
6R0e/DCK33o/yoQfgoS/IMpl4LvsKUbHpRi52t68qyIICfuXvFR0fwfbaOB1H5zCpbXomx1YA6Ug
HcviqO8lValUtgCGytbrhkMlTq9xYk/MdPq/zZqhYMuvb4SD935KnTVrknUEezpCb3EZ4KOn81qt
Vv26y1BETk9Ya7DuHIlHR4VdUiWRxOKPIFySF00cSow0ehUayx8XDlJYIqy6fSGjs3aZjL3iwJE7
Cer1i3FwQLgePSfmEDKt9wTQSLQb4aLdWptZvkpR6Y7uBRwN2IKSgXGcUAsvf+ChntgiShJdCUpE
Lm3QDCF6m4Wvo/yHWNY6BOvhT8WrHcscJhh3v9Nk66XtG+TqJu4YLnplaDXtL1cM4Gu6q0LyACCf
TkpxDMJJitKxdBsgtZHiSDJ6G+9bDMqkWt5l+/99lEruBDuk+xEjpEodiI6Im1VXR04fyCv8yf+1
CZVRXRkWCjbiN3dF2DAbc+Et2IMVG5vW/rqrNZtAs6yeeixPEto51T8ctiIq69zXkI9464nSrmDk
1m+pveVTZuIJRBCTNE6UvaGokjMUeA1yByg8xxT7XMAyKJfu+ol2xgiIeJhR+DPRM3kdJ9NbejKH
MAPKI9qix/4OyDYH2xkiC1Mjk04yD3JWNfLVowfP7FBdBZ8KaQouuBFck1RfVOCe26ctSLZ3aEiH
kDeMKUegPZ7XFk3zeUu9sJJlrQ/+6usvy0ME2qXJ4Ao+4/yVJ6bM1Blg691sWHxqskbNTer6nDk6
zdi6mLECA5Hio5EpYPntCjRZPpNi8RH4nrXmQR+7Mo7ij6g3evKXZLXMBJ0chp1oL6CpGLYiC7EE
sNQNHDV/7He7K9F44qURngMxXqVXyllBu09ja6XCOvu7cEinoOel0C9+gWNDIQCoFq6hgSWniRKx
uyJfk0GCluxhoYbFAnOjudVB7dNq+NM6J9bW+RzrzPfN8hY4G264UeJ8NCqiioWgIA+3PgotTFXb
zsxCsFErXmyC8lKsec+qji1idTlzXaspWMmEUFt4LvdV887XrfNR9XbGPcYfquT3R6gheS1KaVWB
UA67Eb3qOyLnqtW+T84Rj5+jOxnPazQImkNuNzjaAbU71/FhDbM2UUR/E50J5YarBtqUfJMhQ8Cz
Y0zQX9WljP3sqBxCPejhD1LXAR8Aigr3gEviwWf+zOyG+Ckwsfu8KlXxfZeuYd867jUpFQ/TsfBk
i2HnMWzGld6AIjSyF+BpGtooK9uPDr4xB4OzPhfbsU1a/08iiEnfvJ3lr/UY6E4Ma1bYX1cJyDBg
giUhwUS4M8c0nNpSDIXBHAsBzKL2Pa5iO418LvpLfLeLv4cAlc8h1xmXLCDk99k2GCids95Sgh6n
yTTIzSGxQJNNacfzHU3exzI0OBHvZX7R9K6AAF5vGSB3xK4DHt3dytJWQcRusLIJCxqU95OBt82i
AIHeu2CbkgjUbHSkByRYaTWTYNBiXWVisIusZ9upsMRJR2Vhi5jtzotEej5FAgaus6ytqYQGklv2
4ZkPQK9Ym8z3C780NxYctJq2b1PQ24HP+50XhITm9KyKRaAdun1bXFt3o8kibcupNLTMP8EHl/9p
cnMtxlKDChKmR6LWC5HSNim1rpzNaZhEycDfIcmv55EacIRUBx0eFPPDNk3JfMVd5YXPYoTtBkB+
+NTHNqJp5J14/G81PHLBwdM6BxFk7cRgJINBFuU1JVZTD+oFak6FNyDHv8ZLO7Q0ZAqYULBxXwvp
SP5k8fhVCq09JD2Roeypg8ONBBxRS+0P6/+Jdhp3KkHAN8TILIemLZUVaabHe2Ryu+JJ0CW7cFEK
ojJ91IKnGAIOZX8pY0sRIZlULXZmH/GkOiwR4SyL8IZtK/zutftG8D+gE6dr98/QdXa5zzd7pNfU
SyV2zX0He+NxdsOPvdBYezY28bNv5qSr/W5GM/QfyfWHm4OII8RGjfo6E67mvmBT+4IPZrcT7Ukg
lL9CqLy2WVZCxCcoTAF+zMHsYSd2qS8ITH/bXtwXpwK/UWlE9/QzyBKyBPoZdTVP92Mll+ekGSj4
z/bGGYnFI90GlqYxzFFu5DbSFQ5qiAX9PbpVXRRHZ1a3omR+FTrgj46e7fMqz6d+Z9+MiW6+Onid
0SVboxbHnxQIZfeao4pZfzmBpB+EZCm4niZ/EhqxGx3G2puwtuatWqIms9KaDn+QjqylVehrNVFS
C+blqRxfhBghC9wDc3Bg4FgDiZSsKZDGK6Xql3kepQ/u1Cil89yvjCERuhtZ0uD3s/4rTvVuu6L2
xW2d7RcBWyVhIz7MhEogd6GjPQZRViKcdmyFH8GAnEtHPFIzjIvMZ0xI26VX+p7cL3qpVDDzl6iL
c2yHHT+Cs/FDX2Ad1n1aynx1CQoAj4tmMCWvgxF4UBbqXwQ6WF1Bx0XPuA1p9VwzLIwzdgClNBmD
uWUDmu4edkYpBiS9BKu3uFY0rzkPagKGANUWYH5VGNCXo4ze3sgs39zmm82SdsZS4I1Zu8B9auf/
y6xAljaBgoOqQyRZDKlQGNI6dbyApEdLeYr6RzpgyhS88L/oLV58cCC+vz7ozS3rrkeXoKZ7UVka
cej4nvIYxgrk51pAGhICLAohX8sIektCwNE8jLbEFWVqnT+jD93fXT03KLqvHU9Cws0JtLylSk3v
1wOnk64orgMcp3O5p2BdfO5O8tEztAdvSOZ58osDH1E2r2bmuMv640sqUhYZ2Z1po0rea8hH8YcF
Nf7KCg0orG26Dty6ejha62dNQddZfjfAzNI6NsU6lkv8tlP5xg6njiUNtG8Hz8vf4vnDwdeYJ1rn
XB1daFEoHv9VlPcMta0bSUKNYVDC1LjT8plSrwKioWNEm3bl1UmQMyzZW9h7VqKV5MbjWmMFFcG4
NS/wKJPgCOXwK/0+WUOgdH+lxzY/dBvVpNWoPIJHZGzLImN8nhGsgUlCjwsU8DY5xZBZfBwR0Fml
qz0ZEP+7YPmfkCVmtnLHfkH2i4j+7JLcu6lzZdjigb0rcngWRMBB4tNuaYerUX5SPnBd5dSVxA6Z
9ptBccD3iUfJoCUr7Jz+WAj4Q4pBKRA4wb2XVL1q5wGW5zji0+I3qWebFkBDPhBfNJ6Shj0e/BiX
ZoILho6L8QrpTOd3eqAp4wrlCu4/gg0SejF2F9xZ3M/1P33GYkekQT2+mpmLXReoPe+bhooDoHNM
oE6Lybq8tLPBT1flNuuulWa1Kk2ka5vpLYfp5VUD3goBWp5vkdBVKW5FspLLAeFYPPARCcdV/1Ri
uoG+RpeMvMksdShuU8/YuYQEZIgGR2BuvYM5QO3f1aBZBjoMmZWR2zm3LVnnfC1Iym8X2qGIytUy
5nPrVt8lEQ5Yju9WcvMGD7+Rj3iQL6tu9Vm30xxnBo9rCyQkmIjlemE/4vkQUl99lB+N5R8AXDtS
1JuREYYp3Xy5k47qFNWSjHLgQsvCR2V9Phh8AdTSVoP3sJ/d67ykvfT31O1lER6rOzaPw8l6tqke
JgFlcb4Hnzg+1dknoqnVB2cai4soI85C4dwcbnwAUmIKfRBjo/JID96JSXB70q9wi3yMvInOYGbv
VeVmFEA+CNjPRFIhnDmousWw5ouAK71cPMW2FXDbHKAi97uwHTErjlI/5Nq8pp0kXe2ywAqaEJqr
oElYZETXI0pa/LOfAYD7dbrqqss9nyNLvfzD0HYhEe6sCf5cCfmvJpiDdl9tBMMTw2eDNIUd4Joi
Maa2HYM5/7nnYy2/XzBfskOZIJHUKxTZdMBISR7/+DxfPYTeUfomNlRcVFF7TJGiSvLNshzosE5G
Bva+IaMo032aoHfQ1pgKzdRIsIRz166gQwdObhwRJKeOeEjSSIIvyhzUxnTtZYZiSFXOqYamFBlx
voKUSr4MFTo0UjMw7G2WtVClSNdPrkGRnczT7ZY6pP929fIrOvydPpdYgHvsbyFEoxUjBePs33xu
o6A60d2xilqpv7wCVccmsO7pFDRLRiCILVOvIe2d+Ewuyne1mkPhPUAG2nlkMjO5AETv9Oz2khs2
LKaUCZwgMyXKY0po1d7AeQAXYs269hNuQl9lExm0ARCQ5YBG1XjjhflTA98mCdiKZcrZpQgBMlhH
uMTH48uhOB6+NBNuy7+sO8y1+fHbLzZR7TA/UmcJVt/tSGW373tiD37SzqQzM57pxFzGay2UACOO
9pk8vkeQMKxzdJqeX54DGLG21Z1fu9U7AcUY3gvPZzUrkP1CLS5AQIlhzeUkDuxGlI8D6ucBBFih
6WdWMFO919fiMk1MNPIOCNi2u0F89LP1a8aINFy3wkWIYULayPW9vGFQ0uTxa4gFeUnsBxv1BWje
bVJgTGgAsVlTsvSIj2iH9obOe2Coq2JLS8EEdpXOS9uBAoQmUEcImarE7Yqoj0aKVHYQCjfrZBaI
oaJuSIC4TIW+xaTes098BnagDCJSlS6KLpWJPAXKtt0+Oq/0RICBUhN4hkiRM5myhg/wpGvFUMJg
WJvOwWZXiiXxSZ7cuXMWPqOuqz5bnyn3x8p1BopP3zJvguMpMgS1gwTrSU3YHAtxtdPsLhLRZpaF
UkKSNYr7XKQIS/fMuGFa9q19+9fpG1dcLTv7iFlirCAfiknHBmXaxqWKpALAwoq8N/6Ls4CyQ5cf
ZhFh2ye4EzeIqWvBwD3MDUsZYetKv5bkoFmPQwpHPa6js+6NqtJ2tpAxYQkUhO4OQl1yJuGlMqxF
jkNWi/lfoSgT2KJ7dOmovOtD1QmH1MWVJkJ3B3SW4mr+1CozA8EO0n4MLnKll3MZJ+EgDZmmG2XU
zOo01idiYW62W48zhyBRxrP05E0MnIuc/k0zyP48/+eff5T3J4JlZd1aLFnn9K1pGmam+iX7nMTH
aDRGbDQiscrDNNUiHvEQvcTKLiNjroi0s70s055rWl7cHQfbUmYhEgk2kTMa92/4iIEXJ6nAHqBD
yJS88wrMdjerhZ7VET29pp3grJi+Jg+OcMvKgILeCSsOAr/Cr2msBs9LyyaOnruZU52MjGvqFa8l
VhBnQHBcZF+pUMZ8kNOGUPDWSFGSix8B21CuB4VcWFIGPl1x37K0j86PxI8DDjyCe6L/mWMr2uaU
VQV5mO4meC23eqVFV/MggWassjOBUygPWSF+SQJE8s9kZNALnTj9RP7Bv4qId8ZnAWCQ3xAIb3Vu
K5Ee2kwaZNiDViGqUBLyYNfDjEFH/2FIZQV7iusS3KjTcCMeikhnVzzBJcpjqBYZnljGLu7yg6FP
GPOugyjzOeCAgC8+4GVsXedsmf7KyaO9VL15nRgYl07oN8/7PG36KaQdZE/m9pawSxQH0bP2Zuwe
7EBMN3bYMTrn/06S6rE9R1R2g7vGKH4KswsluYdf5q0CZOuffipJldgdiKqbiZYxP40v06Ez6mi8
lfyNFQuJmd4JdbjNAUjcpMDHDcTi5nPa+PbLb1t6AUePD51RppfPoKnJoHVEVnSkDyBY5KCOjLd2
UPFEiUump/SDLjeN5OomOOBPUYsqqaOgzMRYFWizOoWnFZOqo+pIM5LqKcPk30Fo6bI8RXQvBY3R
EBelocipYd6MNJtx1GpUvjl4vOkM6P0/5n0bWWdr1Xs/DKnwLkttEDSTZEq06RMocobGKPDOT0in
VqAif+P4dfvtPZVEb+AzMJj/rw+rjGhDOhxJrWfj8QOH0VaR3Zipd4CPktj4RYziJriqPEhYDNvg
WzBcpRTQcljuN7X/0sNHkZ8CytkgewBuMx2MFx69TwSCmUJQ3P3Nkzt32hu+GIYdQSrVKjBvQz+w
eQD9cpRFM+/45hVFhujiw5e7aH4j1NkY/u05kuegB7bGVd68avNHrWS+5A8QmbaseMdwbXon/qaM
fuf4iYG2+pWdEbbImr0L6kLpbZelnoRKlh6JUhrnYfC6mmUxo9Tf+RWfhtANGVAfKbf+8TlqCX6s
3iOCkfpscq64UWDtPXLJ1DHbZJpGNcC5ObT/ik+ZQBjX9WDANEpbkfKu9wgR4DE6xo7rQsmZHxiZ
EOtpEE1GwLwpGqvWfJTLU1lguBnqlm+UlbcElkzXWqHMtmPxGsXS/x2eO2mFf7Wn8BM+ZVu0oNcM
SYHyVkGrFN4gB4IX6yujDgkDa9nRs9oN/cGqNGOzmxla988jmVJCe+eu/NnLaVED6ZxNkUt4efB3
DyNQ8WqvsEn+d5ozMdDV2vT3CK3y2in8lA23LcEycrcW9xUg1pJoL0yOUaMYcd2e9TD8ZibEjhZi
xgsxR0/xbVmDK9cKxiOddiU6W/Bx/YPJphQzAZDAAX56AMl0zJv2pZmrwx3LDxmOETtu/h9grV64
PjL4kdrlE6yKc2yu2Vi4tp34/StP6qD8cQ/xuqkhlpb+7nbrHNdEH1ngN7cuePKu3+tWi8eqH5T1
38i3w+KsxUqDenCe5jyy7hp1g0XGd7BwmC1R7NQPh5gxbGSEwZtJHztpQH4oj1pEZ55EAMHTO/DE
43U7q6o9jyxZFdDiZ3F7rt3OJTkCT8X3gfI3r+BeAWjGVHOhoDlYn6jPF30TUgs+s4Rn7CkJDObo
R/9Eft4GPVTB8IGOaeX4hCqujp2pJciZr1dMUvVEl3yEHQ1XkIt6IKEYcsTETm7s1RtJwQSx3sDr
rrdY2azZNy9dIxIJFJ81nvKZD9Bup8Xu7/ybaeAami12a3BcSNxi1hNfss12BNk/Qol7eUJvUO6m
RifpfivAKZaq7W0gVKt/fHahKdhlCdSBCjKimAC++h/N7Vfik0HtbiPThtZ+WYpIKctUOe6xan/e
FWoarGwrO3p/Ve8FlT+o6EiN3Q0Jt3WQ5fU8dEmw1kCIMPFefr5VooQqLVGF7iJgsFqHNehulgHB
xaRY9h77AI6Ewq4vmBSAYYto4/6K5orN6EJCT33bKSo4WWXNihpT7jMhBXfZ1EmnkxIVYi3PZCNS
mv9HefFBrT+2Q0XSPWkezxF6TH3PuDhAn3vPZ00iCOC9l/wx5tnXjbQiUMEfMtlQ1pLBDI1RUD0Z
FOAIPVZfenKhcMShg6Ny42USWUmN4K72WQw1SPF/O4DaE9iwtvoFcaxyz9/RGLVc92P3ePGACAns
w/fusEfFhvAuU4o6zu6TiVOMorxmqncq12ZYCvOxWdVOOvcJQcD9uOUExipY/ZNAO4cy43y3doyM
dFfy03dVN9BB9msDFMk3rS04OdXLtrOR0HatROl+aNfNLIj3bNK+XdSHcr8AH7TRsodF7mr3JRJQ
Z+SOcIPyC6V6jOG2Kr8uzxdmjWa5YkWIBT1n6VbW04LXIXAPlgFP1o+Owkm++ksVN5k33b9s/FEC
Yer0VAuC6an1wkRfVhGNiLKeb0aFgESA9OzOo5tc3pwYf/m/TI83ER7qoWoDUe4OXxm123qmLciW
mBBBjtIcBTirEgOQPmntLDEwc6A4WNeB7wAVRyw+IaR5CHo7se07RAefVoYNuD8gcmu0ADNpqozM
95VSBy4umXWIWvrWcjrNBBoS/0D40Qn+fB5lUF2vTfasthluynjl56oijcwTJnMHZh0H9aOGHw4i
47elcNsfKdKurW+ietKba4Ec483cRgweDgppBz04GElVGggoPBW3vRlTO/pnHwvYLLVwjK2s6wfW
iL1jE9n/x8ZskFoTTHwIMYVAHOy0n7BqJ4bDsHm3h1a4e4Pebe92quO5P8Cw26eQk1nwKvdi3V2R
XJevZvm8omlxSDN4XQrZsUakPUNm2EQHLb6DRXMPZhC7hdRuoUvlA68/Ao4/e/Bi9gMiHFHXHXyd
Qa5XapirrqRcujGRMHNSo6LXnV7CbX72SeuYIcBMACDE7l0eceZoUF3tTSOgDO0kDtcUvd7DfbMi
ZBM87NSqHhS0uNRxbxblO5VmDxEwXutc7qfIGpYN6yIkEYEUgB9lnPvlxkFTNsp5aYRaeUS7HxgY
kZU7co1vEg3MXQZ0whJi3gIjjySqVAN92RieCLRQ0J0DgcXT4jhup1VsgbLf1cfoNANStTg0sWnr
+A4wepaPZDu2Bg4XEnSOGfSe0dI6be58vBKoZUyxeYc8N+tb5g4oyueeTDgt8H16ZfFlkp/2CKqO
s8aJstBzwnj1RsLGYPDWRpWMH+SsM4sN5NXZkARsl/cbuOHGNnX6YRe1S7XYxVKvvxEqQthP2vRP
AqJhiqEdtf67QypfIo09WHDBY5zHJECj6OsPjVmVr/+ZU14q5czZqeJSEf66qKE9GkZUXQbcTuZ8
TDYkgxHXIVgJffW9brG563G0CZOErkvahnzrS8TvqzGk4zFeCxmm+y/ALUWaVY75oiJXtZbjvca6
KR1Mkw94bEP1ncL3QwoFa2HpZJxdiM+p1Y5qNHmfgaLKg/xDqxRpLHvM3aVlLL4Fvywr9HHI7l3Q
0QIExaNn4DV8gU18MfO7MdYyXKMUq4LNVvqqd6j07lfWVvaNCZ6/6uoYRaWqElIpb9rcjSdypaNy
eqFW5vMK8O7T3WtYiE5csoyIx52Xq4Vg2j2yIqkmSd9Q4FeIPZlTH8er748Pme91fdtvplawE8YZ
oxVAk1GQ+0rdNyqepkGmfvFcoPQ9ulHQvZtUo+FAEs8/cFq9OkGwdelU89V4oc8sBpHgaFXmZVt+
l6HvTX3DLc854U2QQuZ1qgdOQyuJdJ3Pm4NsddSfdR8KeSb2QCh/rSC2LC/qvVVIBwtM9egvcXRC
JedLBbuEljNSCRiQjtQ8ccDVssZaiK5ObSrIGgfwdfCPqiQIP2u+D7z2Zg+Pzir3xgDWLRDfdm8A
LpmcOvFuPRt887s86aP78x1QovAUB+7SzSo01yF7+gtqXViN0vOrot9ovOiUU/+ngIxqSOqaUkaW
v8bpta1yONcIIBT5b0CzM8Uapr6jES2SOnA6uPn/vBuImqmC8gzdEYvCncnWfPVVueiPn6j05Jai
pXcbcnm/hjenuBFNMdwaRY7b6lUVm+LJ+AsyjbZtRckGa1poSuh5NvuKVe+T+W62F85sB78CiaJn
R70aRbTKAL6fnA/Mpx1xh3+HJyCTrSE7eNtohMlTxtQXDsU+/+Y6pvwW9asvuPObtuCeXejpwVxt
r83DJkOGw0n/ij8EeVoQRHjWEyJRsAAC8PVsShK/a2vdW7PYB6+9f3CXoVv2WQowLxafHk0kenrh
U0vR16Q7nddlAmr7aJH/NspY4kiacT8Fklz1JMfd5Q/mblGjU47WC1TYVtc2JGOZ4hAJ9dzhxd9n
zZojlkX/7p03qjbL9STxZlDGC7wL5YAhlna0HrbFTDYDSvf8CZVSk5HHbC1wtdAsqTVt4c1FfV8D
ZwSQwYitrkt+uLBVdAvcz6CKWd+qNrZXuIbzJIXqJIFPoiTZDzNJG8slzbmNS+J5/R4wX3Bz40T0
2TbImxzjKhFkepJuHJHf0I4kz/lQpGbdINlvZh2rf8GUlPc7zqJe5MFlvml/8qaj0vduTCaFZ/Ot
dx1U4PnXO/cUhJ6wmDL3bvy+HLOS44iPb2hSVs58pkD9+F88VO1FCS8/L+ht1/6Ztbn0cKXvxnSl
yPoMy8/ZHdBTWrrDokYzgl25sbMNT1webuCiT9wynVuD98tHBPIODmQNwaeduVVdQQNec6lwdZgw
8SFtTHWSA1+OG/89/Xem0E8rskM+Gq4g/Ilh21uvaccMyE/wfpbLWRhtG9lAvCjXAJwL0f3BLBBB
61xTKW1b9HeBwQUNDihT2Z77OBZtXoscIUgxdtHU6xdK5cnhBS9rd+vYyZg7EagBd7qO2QGdp4y6
OUnEG6JhTNo7jDGuXDKfILosvRb7oU4nZZ4Wt5ACDA74tmeZpmfWxXll8pvBUy5SOkmz/owyqt6j
blleOVjkmf0e5d+yVvpJrZ4va4xpXcxwovl48MlD4nKYvV/xbYUHGAV9SNfH/hOaI5mxeTrpTGNy
FTo1JbphlOJReNtLSyISe7TIdLq5CJo1I+R53t34y8bhhcu0961nNCR0e/89tVdvR+dLtEU/5p4b
jvN3fhI8JNGEV7Wq5aa7k30fCHO4JSYYzjJN+BkG3EUHNiOQkFhmAgVlUXbBhjCp9yLq9YzRD4Qh
/r72uGTARMj9a5O8L0IRxloPYUH4xfPTai0YiCl43midTsVrQ95Y86KNrGuPnrgezzi75/nH4ZUy
t0iWRPQzlayWmfBi61FsqPnvgzGiaWbEVf00dPGBavyRpTOR4Xq4tRmOEWkm9RaEsurgfloB+GDm
KCftd3lcoMBrPNTeO07yIN4jdXCWpeDd2l+6h70HPWXSoD3PyJ8NrQ8RLFUtqCDpDfClVuHS943c
ump1mWBjQapgP8v9yFE2nDyvM+Tq89bTTdhY+eu+vUVnZPF3x9R4p96eFHqyiLxq08kBCYVLvDtt
ZvljYPbYcskuL2mHxS0iAxpUTcLGtUhf/xdKRqonahY7tyuxDa61dHs49kTEIKOusCu4Y5THs7Qq
ambq4MGYpbAg55lb5ozywOGmOO5WYqowqDlKbY4QaIyY0yq1mqp2ttQ9ORooONYDi+vIJrjSbfHH
eTN8RssfX0nQKrYiWorb7LDTwsYKnIQMcYl924xx6g5pOB+DdD99SwdpIThUjIxvVwkUnHpxJq8M
9IywwwDfLEgRs1u35hjpzysVioOHKFOTdlNMcEFFq5aIcjIJhnn/tA9xBfeX18d0nALdcFQLqd2q
sSKl1jcz1BFCGD6tRARUpQRb/GTfnyYjx59hp6sx/jucuApscr5KV1d5wWMaXS2+1DD107lTf2Da
29W4hXnmkFRr7SDFMPivUNq69havJnBXtK760staqJmPf67p2khmVQfTGSc1VRLFbfFhiUZCCoLL
8V4MEWhRVV03onmQZKVmwJCIPmwFkYIZ6OY36BeJ3nz6ZGXOummTDa5IBgda8c9kyC3q6kTOBTBT
A7OHcTn7fei0GHvQ3VSvrwhC9cepXJ7cseBFfgr4zFTIeRAIUMPwV/OajcvsyHStOIkaMMSKSfW/
Vrk14UG/55YmBED1SyCD0k9AUies4iCPNekgTMHWY17d9Rlq2XqdM2naXFQJt625aTmB37Xym9bF
I3aw2b5W02K3BR7YpFW4rZZ0DTGOuWxuwqGsHN6+8crOZuhXQafOJj+8l/1/rrzE6TTrMLsFKVcD
65/hw+ykl625NLOExHn74uZF8Vj+ZjFMMR1Z97rBYoJOl2wkrWWPTFOxsAQ5nrgmPI23SgwbepPK
cbnLATNvK9tX4YBz0HMNJVrhtpKTXKEw9ooVd4EuOkNn8rBDT1zAnkQFXh7zsO/KmcMWUnhCm0jB
lAVDQaYq8gQOxbZxplvLb52EFHqo4G/WX53TrVpyBZAHw9npSwceueWBuxwdbjb5xgcPIHez1yX+
HV83BHPukauNuV+t/rJ/0GuCE3gNe8AyQPH0Zq3NbA3Xj/uIJMr7WtVaE3QveP7YXgnHSP7mpjRn
ecGfa/LKwFaHCg2e3BN5qbyOTtCoKTMqBUjpAJX56kWvFBNGtJafSk4Sm5kYfoWm7Mgrj4ybkT1t
TBxOaqZZhEkPnbXFjqqTiycwjYSWq4/06ARLxWtXlO2dKff6H52zW0sOZPBg4mIEqVNhFgjsf+VV
hL5+oqW5Yj+oTyrrih8KTI/MxEjib9fUgap1dg36DoAmxmy0SUMeUdTl/Nf5YbKDIISHVD2WsmDZ
qpepAVDBC4Uo0YmzAvGx9zPUbujbGk0LOZBWhn4DrEv/YUxAk7MrU3X0ZZMnR971+VjHLoVsI7Lg
/JJpiJdhvkyhi4h5q/jmXZEJlV+R6Jffg40CMK14cguUtreH07CthkS4ykTU8dtGJjRtHVoYia7u
gACifnKIsQzUaPAhKIFT+cBlPayICXQVX5ea0IXLifXCXhoA1eRawJKgtuMBU4O+l3WuFUHX+rPq
0zwEE7QEYEovEhDit9E2vb2Que5rGWm6vIJXUoJ3BCyJLGQLEO9JINm8AUm5Rn/MyXj5irkzCrV6
/aArcsBGbUM6KaN/ThRksAzkW0Fj3lsB9ZU/nQmaPAWv1Rtk7aK04XpHZywO9IZs3mZr3GuBitsL
B51TS1GzaXPSULh6W3SuwMdexAJ62oYTBoZjZVcn7yOm8x6BBwbBqlbQakTMJ+b78wAdNz7hx2zx
ExD4Tx2m4qq+UbsaRIEEmCW4mqZcsePX++d4KGCymIeetPvmZig5Z36ZWcJLt4PcU/LLsAQQbP21
1RKj6VWOsjsLD7bgvA0sJccwrZ9OJBX1n1ujJGfmmHmVNLrlzJ3YKcrXfNRpebjCChmi5mjv2PzV
DxtJerid/VjqtpS16X0RE9HhUTBrtqFE8MaykZatQSCR6WVTC6R+wP0Jt9jkzaAa+uYpdXgJImL+
uUHvv/xN2HjCgR0WZcn+ij5xwAIPkgVxZ6yGcCH3q+gjsxDllNJEDr6j/0HoLgZ+0Cu9VUcal7Yq
oZRAWiQ6VzE8LUNbjeeCbeTiIjytb/KyZZgs1UXhltPJdhSxpapgr+2bQiQzimcl+I0qTLjBFr+B
yNLhzwJoWFvLRot1dlkkrHjOzLFjnXUTpaalKeDIDT8BDGUSz2slT4c5yfVFO4xvGM6xk76NUXBM
Ewh6NhXc4ra7DJTYoK4MjsVsJEKXjDzvVDzV6c6ktY8Kietg1PmnVxYrSIuxrlUe/vV7kGcl0whD
GJxB0ogyqWvAK56ViGnheOIwscleL8AdU6la6b/MXdzpc4nr/1JfSBLmX0kh+WC5kN/1GrIdpUG8
siJ1ijZffQtgEjq5g6c8Z5M+KGxM55Gom2RXF/wEx7Jj2DwiYvGzmjCu1XmDqCdJMyTtAI0rH620
asvyIeORUPoKfIg5ut/Qt39Lx/9Grbgty3OAAY9j4ukpQGwsTmnDRMNBAbrdkxg4Q32NGmkQz8N1
ijEBgjOXP6rQ06AKOEc3kVJ7/L5++nSrzHE94un7960OCHHqrohSmDNmBsl5PuezLb5Gevjbm5np
2Cml9qeuXeAWT6Bczm1Ag4HNdYhhsrhxh71WFrFd6aKjgmBAAyrR/J0T2yJJ8XjrMEWRmw0IgAVd
jtanZ1pc+0mjeAxjyKVtlQkuigB7TrA4o7J4AdBfhTEUfVb0vwfeoRXiUq04FlBlIjVVImyYI0R0
8JQ08pbO+GMPH3xcOTq/TJW5XAfBl7PP4QIel+Klk5jp4u2NxyhO1JbGoayQRxO0NxA1k1beu0st
1ANFRppOqENLNMh734nFBVmQ9CYH/GNZkd97S0zmHPwi5YWLL/A3m0zyQxw9V9N/88v9u/jlVprw
oLkpIKgf7VC9efr4ad0BxTzQmDvRp5VXnzAcLSmpEGWj57XmwkOqMezT1eE+zv725PSpvhWK2jkH
ZT0zYCEXeNRr6LvUb6ehTHR2OrMuXt9TIh+ZxOwiLTVimKuS+tIU4FNv0CcgvYZvXtMHnyt81kEA
/TSk0OGghmjxBnw1l0/AUTqb1TRdHy2kZIejj7kESX67p/JjnUAIl49hw+D9r5HsVgJmBicLbBex
8VMLSuY62O6OEBj3/XZmdMI8bL0GARvf/JqKtF7csgTHQIXsoljhR+XqniQ0ayUWL15aWLxp2wzi
CJ9oo/nAcm0NuUk6blnkwn+mLpskLw2trHGPjAALChPUGgWOvqpnchyRs2AN7aL6a5dnRaUqLPqy
K0x2yShKGMdlu672q15wouMp9Munt39bW+IjPt0SAYrRcR/2L6B9HPwnf1YYs9sIxCdX1mZJ5JE9
xF2aPo0DEcZDcMbGQwTrju1fkuu1wYKwn3CsWXf1bv2n5klxah/mWqJxcQQPMBbXEqqLoZUSSqO/
oXm+i2OzyRFRW/lsFg13PvqzUUcDqf6I7UQZO96+1aUmLXIZ7/RgwQW47GtapDEOIrboQslg/1Ov
mlKyERxZx40ksSrM25lkTpBfjRaaOsbNMhigbIKk8PlMFdRzxJnPLcoRR5DaL+7Z6BzWLKW3URcw
rSWHF/BQPDcbmMOd4maYOOahYdRZq34sNAATu9u+po6/iV0PjUlqAuwgW/42p5IOzbxdyCcPmVYw
qWlZh2LZqy/otWtNyOLtXmkX5cKuZwnpuIjpiI5qnGhU3fikVlFn41zeWWd6kBqtlBQiPkWGtFv8
Wd1xZeUXx7GrCAcNZiQGcc+1T4KG98IgWiPbSkPbWOaQshQUzxunj0rMdIZLwXOFbGY0GR/VHCVk
/NzpRI/Vn+4PuG+xWcZ06UmTi5UCLW4W5HKjpQ6F53cdDimZR97ptXGuWFC0AjeQxvqXjXuUNjG4
kboBpWOFuU/U/2UW/xYjC3KO5fionYQDFfO/oLKoXcYmHbTuS7U0HCaay2A7X6ezrjEJqFdX2SZy
bXfD0H5N05TwhjVl/uB+9xBkDgD78/Vvs2zaSiyWjSC9h0KxFuxA0FA7p4BdosvzzPMHr3UbxXXY
Z/Yly7EiUs/deMLhaKhFZK7inovU/1HsLKB2JMwE7IcBaEKt9Ypip1Ly+a20aCH80TKhNoYjjsEx
OY08ErACgIVlctGhLW7gUU+CCKN12sTZ1Iothm7UNI+72m+mpWkluM6FFuYdnf1Uvs1UCdAJvASE
upv4LpZdWokZ2i+c7r7LQUSqQ57/1naqEvzlQggW3XMGGaiA88G9uNTRCnfP2FoVwt9awSxtdBhc
IzHaMihhH2GfiU3uu8LEZe2wn694wt/I2eTSDzPsfAuf7SA9bvV4SYhDm2UrXhTv8AKJtfy1guYf
u3PRHz7KKaCk9YZLI2Ab4j/ZRC28akZ2EiiPQtF81egw3p/QNE3OPkH+Gxiav3L4WAVXVFEnjDW/
vsPtZgwEauKbq0fbBiBK5NdjQqBPr69lQjhA5wVUUhL3fQXi/SenWT1r/Kk/luN9gg5wx+WtCLxe
Zbat+yaSgCPGZ5+9laICCZ0X5ZTmGw2wkdB8nWOYRU1hT8zccx1pC2L8J6eedrTAJxace7w6uz4p
7VUQhijVmuTcitARQw3Z2/NkCFRf7w/Wo2cyFuzQVRrX6xRYkeVLaTTJBM+8n5ujZbKutuDZE18+
SDEThFkn9IxLYCHxmH7ItGSFkF7jqR86zpjj6fM9bprxYsZ3foDP56jmTqPKNNyTe72fVhJIrLmc
iS1AjefP43NuNSrQjL/JdFsKp86LwIGXdehIKtINeAO90w/kF6703gT/z1jxpz0p7GXJJPfwjF2i
GRin6dF4fQMI1pU89oZ4r31pUJvgKMm7EEIth5gjLFgqgGn+lkzRVzZAQlpgUJjCSFxjE0UAYYzZ
MYsdExXbIZtseTgBAnCNhvQ8rbZ86PGoTc14YRhFDijDC/Qnuhv/vR2nbKaRX4FN2IJkjetniwpJ
S3PmP8DZzQX7xYxMdoo2QPf0AEu0Gwwjpjzb2jolsrxPcunGV0wt9ImUxlOPIcWEQ7mJFJ95qE2R
4j47CI9aGXnda9dzqrIHx2wiHL6NtEQYenpldNSa15/9SOpAqHgAlKIO1PTV3xN57JS1KOMXf0on
d5dz8BU7FVMLJxHqz6Fz47N/5EaAkkrzk0Tb2sGoErxcy3p8MbjpE/TKNLKHpBD0GsxMDN9VrQmN
X/BC83YhJReSY2FfteqLGt7aAZsjs77prdSNu+iy4pjFxfZAHgetry2UFswY4UJGKdt6rDSfTWd3
EXpOhd0x/iOmd8rXukgGkKb6C/HE5jvo7r2/cGtbYgj7zUnSx+8jS1+SHdmP+RVYRKC8Y8wctIWy
wuHr+Jl/qXfQBUuIPDYVUNoUCAh+hmE0JUWoYmfM8KrUw3LGnOAHkkSmoqa3sgWWcDGKXkuCLl86
I8Ef6uS283fjlAAGu6mlMZRmV8aC4hg8F3EQOBMV6c4m/d/TZvS3by/OElWF2I/KLtqtZVfLfVqK
W7isQGfFyiN9fRC2rETDVEIWR7+s4hYuPRaFkdpnP9EH1J+SL/iRJjikmVA7TAImb+4YmTnWNsEC
tzU4Q2kn4mF1t/jtJdTSCdAlhigXQms+8SlRMb+30DPwJJswYWu2Ig6wotQw9alaxd2/nnDJOise
sSnXKnvc4e78tR7wBGxSfnuo1qgRnPSQUiEZA9Maf6eX9Q+SYiOj3KXiNt33wOWPCqi7BeJyCEie
VFnTADn6zpbWgwVDYURpw3jAV2d1IJA4g9Z3NcmrkUin8+JfIZVSuW6QuTx4UhrhO1pfWI3LqROU
bY1OiOXzJTSzD+T6VeoJ68GeaFHsGXVZZR2zHsfV6mzM/gGGnPDbO2NCY83TiFUwt/4YeEg+v5+b
57uxydLXekJLkO//S2iYzeVQcnQIjR5I8vLWN7tzXfM3jqpPAbMx6eOC0aFhQHVee9APGtpGDEHa
XMWlKytpTPJw4t+PqCWZoEwI0y3ZXEL+x4fB4wHkedkQN/1shS4MnbnLi1udbWpO9gtT4EGD02bB
N4TsxwZr06LVEKWBP2PWD178DabjS8S29ASlSxmcGuMxr2psrIqywsFgiycUnRkYgyOCpcMkR9eV
i4Ljfp7tZEWtHsjy6abjj4v2RjQlExtfLi9ptntOUu5aIiMNU2RLVxc1a3RI1tWB+vf1+agV8Cj1
6+QyP5ugtjhuIiuBKGv42tb+sjoup77Ukzk3iDmoPXag7mtUhBbX1fM+izhfzd8PTDjzOc2HJ79u
A5wwo6Bwv75qovpgdqJpqu7ycEPg0+/zPt1kzMAqi1VfNHaQ9BSvHcnqtAjZsqg4P4iv5p0ijaLO
SmPzroZdnBtbrFFPYYyNfqJ6PBHsxICX1NJfw84q4Awk5IL7P82ekQ1qqHPye9wWgX7q8/3rG/E+
o+U7HbOVxAiGfmr2lf16ftpAPY7ve+BKoLmtbBMnqxmIjhKvnfFXUXiDzYUvcTfwnbn6SPY2zs/u
M23wWcQmNAmdXCBN/YQq/bl0BCqCVi/poRec2YrA7IaOkSRYbA7hKk540l6E7KdmaQULx7bZ3rKc
lTEqnknD6d9YhLdUwasDtPcGk7sr7Yb4oSmB3ppT3+uirjTjMmWGYLVhyDG151IkDFF5VsDBpBG7
xEvXUn5LHuTIQwxDSYanup0nxmTAgU4Cqb7iHqEyF27h9Pe6hczPu20tOmzZPccsH5HP2xhHcM4C
mGF7v1g6biewurV0z8vhMxNPkJ6A1At7ya6hPv0zYV8RZKaPLCaKXldzMCz9RpV59Qc60op+0Zm6
1QdyrqivuFSOGUjuSXuqJ5jayViJN7K7Gf277Ngxbvhfg1i2y0nR3MXdV2Jhi+h00gR/6yGO14Xr
BiB+tjWWYEem+IFlUmyuawfgQ3rPKjjESDZnIR5WI/aGxx7JJyTdVWoU2OK9ZwqBuyATmAirWFdU
cpOQ7Sie/M9dcnJd6T1qoW4zxbEYIQCPd/plZKSy8iE8260bfcxd87iSpx9S9fAbMQMUU5n+gzw5
wKuPVchgLUGpdlm8lUu7QTczJJozn6PY2dDb878ts3KrclTsU5z5jgoV+KwJk/F8UVNTu0vOeFq6
hcXayBMOEE27G1ZlPgx5GI5EZQVgg6xC83JXFMiJjD1oh8kkuEZY7oUYCrIZke7jAxkq5zjAy7hV
88SmFrCcESQQO1kajLjnXc2aWQQJGOKR0AXYYxi3zQmGseX8GhMY05Ew5hhOuwThEqy9lOzcgiA0
YdBUufxwCjxHbqIKIjmXI1yX5iYlNGD8sUPJ0zUhi6l9izTLh5A0v3uX9YxJlL2QXCEaNs6vZmoW
K/BpQo7FYToC7SPg+0JmQ7SiwlLrn0eZV/HuvFDChgMFLAh+VhpU1WYhjl+o8RqD/rX4KvnvkVyp
kgLYp5v7DaHN9mfKZJnyzNhfi1GJROc3AzVqY9u7RTeFay56yY47Q3AFOW70pUiP9Ov+k1fGqY5X
t+upFbnE8bTV8Wx9Cwx26vK5icmLlkE0Pz9lg6yl2vtyoVUDNeFG+g41YiqGUvDUtbCrixbNJgsl
HGanfJIq1jD0lZqogkgxclTIpUtyWzOMkfhmg+xvwAWNiBpMP4ct/7rfRUM9OB/jWxYc3cReVkLl
WRiz0sb4uZiA8XIgdfyp8CQhgqayoN0ZlFWzueB0/g9nXjbHtCQ8cupsZ48GIrc8h/m7giEd7hEi
FdfgIaUKX8anz2j1YUEMuV1aFOhUX1ugtwCyyOJiv0tdFjaEUH2RU6UqDwJtwd7HK/SLF7pEq9+R
B439+LzTaleSgx5rW3MWja0RQI8zJJTjXWbth1S+sPCzbjsoudXS0EkkHPZz3ZUK7geJseIya70x
S99hS34BJhBCsCT52E08lnbT+WNviGvTAln8ZpnWm0KcAvPs/8sVaeU+IPdOWYVsQtFCK081p9V+
vh6Cj+pQ4WcEOJX150GzZTYN1tUAOo2HZPva+ztHUYws0rUmd/LB/PbHiHvvlUiJykYoOclpz7sF
b1o/3jRJs2AryFbtyrUgoziMtGLy+8HPS1pNQUGcXeuMdzjwvn8MZm7fDqq/PVNJ3BO6DdBL8Ns2
b7uGylvntudN182bAorz6izLFxIbs4BfGxfhTbIypIUXkI1tlw7ZVe2B3fX0N7gSXHL3sSyld+a5
Cum6E/YsZ/Gkuzg1Zh1YwJQL33leTrvAVTbToLJFQih18WDaRZg55vSUgrJ1IhEMT26CIg/O3qhH
LQ5I5EBEwsIdiyGoWgZGMidGQ9jBzv3A/1ixNZRDBXU8aj1R++gQd7Hl2G6QBq9jHMRQQiYmVFFR
JQf5rJG6NQeIijjF+pp3kwZhVCuWu597aOW1kRVDWhGBeN1fo3jgjV6wjApTfoy0TQRRqanXL3Qf
7m5j3opyOfBNkk8MJpj3R+lHQS8hsR3J1Y+4BnSwmTP/LA6Li/GYhcZpu/BkD44L3HT/kDgsRGwF
7bsM9eRw5vS6jh9Sdx+t5iWDBWgFDW8gj8JSr0d7TZC9UGH4JxT1PkWHEPeCbH8YHSVpSYVlFUW+
zBgEOdQVeq6yfvV7Rxy0anCeJk2OiKF/jc74AOulqrnpLRr8b7pmGFmd0h9CuHt+Zvm8MRI55eNg
Pk93XUAIQHmWOyayxRMCqe5UMGlEAgAQhvBhYPxwWkn58Z8DlMy7TBDdxJQXlGowkAxxBRM4pOVw
Ieghb142ksplaV+L1U+m42ML1TOrVyRSOCC5UAYsW7ZF5MBS3w+Y3D4qdpd7+/ZpHMxcBvAZiont
WmiXFKucAj76dToJUHFRYRUHsmTRprqQ4kisqBwv1NKnLA5WDjH6PjVhJ0YlWA0jZEbPS/qRU9uz
mQtGiFsqguHP+Upw7Cxseq5wXkKEiiYsv8XWQL9pCbWOQPmQiLNwZw4g1omLNTs7rNQtGzUIBKA1
FWwrsfhoj8DrJep3JTAhCGvuI4ihE31XZdtBBX2sa3EsxmQ+40xYJVgWfeLIf0Ll/Z4xdTpQOApW
wyfZ9RaxXWY38SFH3aSWkR5NQrQbLIlZtk4GqiqSOJtkGJ87SjDlKiSnGtAR08+Us+dQHnFfaGhK
z0ek9RX3RDnLVOnAk10B93VV6rwvAKKNhQV2FGAv8OrgNOePzu3YQH2eXxcW3tQld+Wnazup5iXS
GbcbSqrVwKU/Xgoj4YS21YIyf2sdhQ6dHeXVxNvvzgHXHnXYOqYxfejjjz8z9U2RYkJiqQfs/vSd
ePqNix3oBAWdF7phRQvHAXsfDAo1YrjxVCiNkRggSjH6FJnfVcK6bDD2YvF7T10IsbKyFswPBsMP
8naE5MRgj7ICkwzf5bj4i4s8+3NiiJ+kO27ETEi2G8XJYcHq2j7dBWeidMagFvbaoNXkdo5+vvCQ
SBxuTdWd5D3byepyyPXLgBeOgqv/BYaedDBzK42VDdZ7Q6F59IGjwWC19ubqF/bXv/iUeWcvU+7M
ciPWm+0ZtXdCLzq4ZpvKrKrPkBD6VgfhTcfHrdIeOkYRABORDgAB8iJCwuuEfZ8ZgOGXALR95dzT
PIoZhfMcnDyYYj5UPMKm6DpHZ//FCplU0y/BXWp15cn25zFdvLwTw+HYz+HOo3w8u6yBN/+K4slo
3GRklopBYeW2tUdWYAhnP57W+IV2QsFpa9EcjGAbokY3fEE6eKVmgbsj2wY9EctoqvCH+zA7Xigv
r79vykd9jaapkr5QqesWh1+D0t5E+vOfsPh5ILpoKxRESwCzhPzvvgqUT38kzPJ4lh8DTbWT+MFr
5omYHqQdhGIjRB/5mFT7EwXNd4Rox5DL/s5HT6Ga761LseFjxMqJsLAwf9y2Plo/IYqU8rma3ZTP
PxdC460WGscPtb/x7h86WRVilZlTCnzNndHAYg/Oblel7gO7J0XWdCN7FijsB7HFX2GRhGX4GdH3
Mrjo9adfEqGD92Lvd+tJIrD0EVgjpLgjyfIk/Bu+iGB1iVv8zrii55+K+iNyzHiyynsKJ4XNa1Il
7zXcemqpm7Z6DVy2jF+AEv2W7Nvp8OI9IMMiGIKtfim9zfH2VjsOt8T5W9JbSZavPUJ9xBOyRJD4
SWTctaebFQVCkQXzbpNYXwntNpMp2HcTPAeI6zXHKh9gfjr2KZSFIsLBWeoQjEjg6Ko6iuLaQdir
Es2aj21NpceH6o9SMw827Fr0oy31T6s1MqOkgDLWnTqROn7nJfbS6mUQFla2wv0p1vT2kXZNr5Dr
09VF50GQM9UNQljwVrt3YzZyooWq8QbRJNSOsPcKvBXfBrXqdBwyajUShLfQy1/i6suGtvpS8kY6
ythXnKn4/8dFd6xZL+t+Vhq8+FOzSQqbnkpwdRscvz69UdlcrGX4S886gwWKmd2DAZdEcyS5V/aB
1woPXoClxoSeGBp61DDRr46oxoFxIyRTIPIcoTAA+G8MYtS6n/s0Jo1Iye99kIudX97Sdi7lHo+H
XxgIx3yEYu1QinGe0jFl9JcCKOhKfD23B1ouqNHg6WZSd+PE7RNdF+GnqTtDJh9fGuiv84cz/VtV
i1N5fSPIxu8MEP2Blvv8H0tMNeEoXyeTDkySyBMMlji5c/iiD3E1rEynVpEoQpRyPKLSnXCJarUN
tXjyTUw2qOqcFKZOiPZoMRtDdXXpcGGALcg02CG1QEY0suIuPwwakuC0+K1xiHrRqCMq4zDRWOfb
5rBPb4+ZuI1+7ZKqiimgLojHQ6CGYQMGHyfjlUL8p7iPwGFAGQ24srbudC72wT6mYXuX3UwrYmVt
wPTg8m3n1U0/Lz+PtkMcd6jtrWcP6bxyu1nkXn6ys1tgr7kuq7v12vTv9NTQTVfGKN2/BgEWhfjt
+IVM4goHqkRw8gYCNwvky53mmDifYEmaGMg2Crijg6q5mYg9/BHcAeQT2dPx8N3hcjccweg3Gjtv
0lltlona1PVe1VURu1vsH4eiifV/JHBoJjpAfbhx2xfaCE/W2sxJkPwLw/BnBDVLP4TaTWUNzmtc
kLRwPx6ILnUS95vAuGWiPI8bm5q7CrHgUO9o8reMu+74I1Cv8bu5olAzonnt8XOY5hzBwWvbhRMu
kDP0nPWmQz2oDjOpxb0MdujHyRniIAnGVN/dIm3GTh/AUXuCntUbwwEwCM+KGeJ25kii8+s8NKmZ
YVel9MjVpzIm8u2KXCwFPtRfoRCSfqkJqjdVJexejjEbUrw3oCmXK6iGDSm0aJcw4f3hlm6m5fs6
kO52XDF8kE3jeT5TkbLBU31SaUpjBPB0Jlv3mr66889v7cayoaVrh9XHcHsue6xlqB1YnQT5k49s
8C9zs6tT4DqJ2NYHvwvGBjF810zf4HpgN1z0BqIQ0bGMrvaE94r/IqFLy4q42bmLaufQwj2skr74
Atpbg7WMw6RTKl5NArODNtRBwIkvqkWy3GKpBFMT4r5zh23q8FAFR7kRO4UYU/P34hZWyOwBh4PV
EPda6SqqIxcL6/fYgYBaStU7MC4gyQzw4jQbOqWjplRhQJDQLHdmq5rDt1fq+vwu7OQ5KtqJmnAj
upCsYkhMNQJzYp0Xiw+FyzCitb5gvPlfgIj6Oj3yjDo7Jx3QVTaMlGVcWvZE+SvKa1tN6eprQuj/
7XO13YGLUWZXhmvx0KuHjXgNaoxoW8wKH4Mh2QTN/Rpp9ucSWv6qSGKHK/di+XT0ZW5pKC6aFjfR
hG6EKcBdJ2ByNQShQvlIK8vs7AQbAQnarM+uxV/COTAyTIQR31Lp+F4Wu6gWa1yJ7iSCgoJgYS7t
necpam5x9Kp39eTVSRI1XDjUntmtStN6VixGNCBHmwE8RR1eWzgUbCy183D3p6fhHV1X/mBwFNWH
S9ulO8qhMUS7mEliXzw/2lNzxvJM/4S0D56wJqY/+t61gyORQ1VOHIyUfuhjyvF0/sdtc71IoflF
Yc82LFyZ9a4KUlW9OakzaZDOvD95qSKLxxkXSMH4HwC7cMIr2BcUr+2XQaduXO/LUIzZYfKR4Amz
Vcnazd4i5xiiVkHaj9v9C1jXpWbSeUHfR+v+j7Qg0+87hHQRRzdS8+fyhxjq4aLedGhkKtPaw/AL
QzN/bWXNxncoZw5201N5M9X0kmBGlXmXrsWeGzqn+VsxfdWN0dkTF19i1syn2pYYdbpTJAmuRJam
eayQ9Cc2zM0ZNEmwk9haRLMqmfWQO5CfRpKyRSenBGpE1FvL0m5/8AARdVqIOcRHeR2CPlvrFUBR
2TXSp2RyIrcil64E22PGz49f64CVrZcKVyYqr3hJ/TPaLkzpk39Lebkh0V+EEnDwLS5OolbR9USN
7nBjUMgd5h3oCAG2Y5SfBf8dYymzPuHI+Ezaf8OecebiZepkDY3CIr6qgnBqaX5mEsyqdFT8BMaG
ljbA4zSV0UD7eAVFj4O+HsJzYjOOI3B+ez+ufvBPC/Npw3GQHxjh9dEoOD/AH0wGkgcl2LjDnI9G
1v/CzKANQQmNWIia3JxLDGxggK5XWnZo3aaNEOjPbdwDIrDaSqLrShLGjlGhr1Y2THSRtpDrtsrD
OgTJ2oFzLxhufF/ndo3CX8CthVoA/7q/YBsQFg0QIMzQSQ9/ernmMyI3TiBzrY2NeJw7qG2Fj0cT
eAXq0X3Vn18llEJGJ2DkH7exA1xUbGT5LgnCIvneEfWsJZrBy8g/XsQeaiT+ObfcxnSJ28RNU2w8
BOb+XzDZwVAkrhf/4FbJ95S7jptbKq3lEp46UDOkXjb/D43I8JNLYFeCYL12gooPi55OanX2J4+G
KLW7VwiO/29wi50IP6PNklTa/Y/5QJQi4+Uxf6IpDSs8dDgyJEVLF95TkCb4xBxU6aml1JzlVL+X
c0Hny4ddfOPG8DLmv4E3hMZEY2aoSs/e6JcJjUtqqaHj/6FiPb5McXfOekmwcsNzcf3doQmWgcw8
yZmgoT54ZvuSYzJ9XZv2UHWQkuf5xm5cSculcNbkzEQGrL5JIYbzO3A1W+12iPNA+AKerN1fFzz8
AqPqLJIZDFWZvRZiP52vxGFwO6LjzG+Sldb3/kA1+oBV7ltYVh84iVVNySUFnVwMfIwE15tX+cpT
G6pDGiEMp/hRsYRiAxup5xmGr4bBer1HGqvUeY5a34aL9M9442qkvPqkAJMPgrVrYKKBX8fVDUZy
+173PqIklcZLkbk1MgHXF6El4+fFp+vLKFgvmN3RFhqseGOfk5NyP4AiXyQn2UMMA8aIh9xwzeKn
GiYiDMwKwaS8jx39DmhNSTwo1t6O9xRKfDJKJWDV0luN+v9CF72HiJFOhUzYS5L6BzajKZixrV0F
pqCwGCm/8zxOHclFEJ9UXFe5URj2018DmBBoQK19/w0eks7zA0wcL2FItG6z0MNyFFBOJ2uRVY8L
BQvNIoqoXq2F7LMzQ+/ZDwsFZZYTA8dFJNuri7fKT34ucfNxQThKsga0S3hHrTVg+gLkzaat2yh3
3jld0vlqYnrNUnaHSpvqE+UkRVHVwXI7G3sH4B5uw2ffvDoAyWFNpilUIJol4W4qSZ6R+nyw/6Ch
3uoHJ3KhWiy5XcJsY1XBCl2AgECQ8yGLG7pcJtXLv65QlkLiqcB4VD7pJpCnZSUHJ/Gm8dJaVH6A
djzu70hsv3sBVXOR3dLDvkYOqFLnas2rNcw/fc9DT2QV5EoszzlcZlG8v+ncoz6jF+zda/lW5NA9
vft0D6ssCDEiCbu2Vt5aDQey/Xbf3c6xe2dZwpuEa4W8b9mYsyWtOW6J9Phva3NDnivderSyv7tl
TfXCek7Vw645KR0zDBXYHre+D3pYOeeHrzoxanvlvmzPTd/TBQXrdVrND1vY9CreJhKKARNUZLVr
JqEkEUsyvG/BpfIIXQP9I4RdeDAAByMJBZbIWTM2ZwmF0427n15hpON7H/Uej4i8j9xgRLBcqIG9
Wn5vyuntofTxnTadnIgzN7qDnN+aqSu/j65+F2DrhCW/beMHNi/PDCF/Ig/uBqbUTcxPUeCWfA1l
n8ShyZVHuJL3jxzfLUTLXJEBXkAZhPUz24Lfcm03qO1HAXYHKkofcaC5S/pc9ob7aiq++QBD3d6v
V79+u+ZVK5n6/bEgLQ3pZlEi/UX6o5LqWFKAxcwwO3p5shmELincsAQ46h7aBAJr/MTnFCM4Ccgf
HUqMFcGYa/SOq/LnP7m1lTGf8Hiuo9pSw2oHHyZsAqfzqs8cy4nbV9PhbdnLKiae1XF+5MeMfDNa
uEnn9htCm0UGgqgfBb/JtumOEqyWam8p4qBlSTS+1FybqXDlmA3+D1z9JuQGrqQlQaauUWhoNtJP
1PYfWTTEN/lQMu8cVr/hCvJuFaOJbIVWRHdZC6wn0EiEWygfeE7P1s246gHhIibCrwDhkacN7250
OBirc0QzPVYn+pPdLxAOS51gRPLBPbQ4FDOik2QfkxrJ3GWnccEfwfX0tNrqrsR0IvjP9hftxZnJ
P27sRhPhd2Uno0+l1SkpGD5K5JrBXTTXCe5zZZYOVrSDh3i7erThrHlqNBde9jB5h7Q68Cr4NhDE
/pc8fmMYVcng8PN8FB1LxY7R8/GmhtWqAPPGbuAn4AmMHhL1lQ2vL+x+lDJm846y3Wwzq2l2nMeY
z0YHV7XLIHsjjiY+LAT/SAwY3xbbXedZcV1EuKuNBUdcAMU2EGBIhQUpXuokGXOKzWdyYZRLtzhj
HeEFrcUee4NRbdq0emRyB5ayRyx0Xze4juln1Te9wSVA8rdnV9QG2rifee7zviw5FmruzLntbIDd
UNuxZwi/b9pnmueHlO11T6tGrXWCbgQfsBZbHaNq8PNDRCe5HQ2/AnOuwW9xeoLkSQvcFj6pD0kq
IE07rjkB2R3ddEAEQLSYFRyVLtGjtRPBZpX4UyIa9PWQijEU9Yn0bq1XsoSrN7u1G2CHowtdEShR
qdqfTa/q8qVAdFuFEAuC2WRTvoj+dxuyeL19zlmkrmQB0iHg95VYhXw8bTLA7YQ+O90MSX0peulP
uo9aP37z+TBAlDALm9udkB356VwW5sH0bIrlXef/Km0mQMf1lj2CLglCo44HQk4ZXh7jLFo7/ihX
loYxi9+km/rwwzKAq0S6iLmow+lpsEtIXw9Els9PJ5mFCF7TVIVhXiQ4Z42cooiDJFo+3G3tr8iu
hLdsCWGz8iaCuTjqYmvLcGgsLVkwIFI8JwKDj/IEnduE9XdO8JGkuRlbryfhXrIOt8rxtLnqFyNz
wIc62zCRB2sdYHJaNPgSGBgBGuWQSqNWNsYmddOKC18N+7z+K8S0t384HZa5IXsIgPX/+xGuBaIh
KI6/YfRtdT3/uZL+b/JoIcO1/6j8M/XXr+Y5Gd4LZBY8v0I3wJjh6WbwKJBviGnu5RrSuEZWk7ky
HfAdghWD2XsKKfbSx9NAh6mx45aD5qaM6e0KtIgeP1YJ4SAQoTBlpw1b/NBBM5DUISha6rqLhgse
PnytjVx5V+s0KAqcnArwtcBJk7i25icYfiHW12SU0qlyjuYd5bu+pfhs9hEB1hhn/UHj3jCwLkjL
joyYeiEfbWv90bkeKfmzJIERl3D3JruqSOG/6DosXPxGuXBTE3ZKlsZdYH1KkqpGcjp7bkQ6hQbX
F5V6tA0gFduNF9gcxAvyWIJ23Yxdp0LDlcEOcYK+OFVhBLL+foGwsy4j+CnLuvKngPhY8db6rXmC
VH9C607Y1qBmmcc3kepKWS+t+S1Pg0M9hbUInU3NC59OHRvmyal/KMQVRCdoV/VM9h0Nh4ALNoks
N+IsKGRMtvrDGBocHdFJ/TQETFa9tWdD3WDPcqF5EaFIQQSy3l4/73hqsIUJ5bqlELYgfsiztyBf
fSKL88yq7w3/Hrwig5cDFRZ8sE/ER9aM13hwdVQ7uyDW7ZP5/nU8sEZXCmSNn/5rZEMjdrIfaiZg
VN4B08C09fvNfnI9ojF0SVG6PcuveRo+oELtWFA0n9sBLVkgG7GmmQaBLtgKsTdpsb1maLzyLCyb
PHeNYUnm9bAQPTFDND3dAO/5RfUR9qXWv6mSBafLK0Mpj61ShasGQ1dbPwwr1tB8bwyrYgN/n9nB
qiDbkBKZG2ZbZVRqc1TsDopv7DmDcWnYsrCL1nXNE4yX7xeD+64cTOSvhj+4totXPgfsGD833bw3
LhJjgwPeKqb/vziUgrMc3cpoKkH+Cj+JTvUNgMZ+dd8P6+wqCPUoRIpnzP+SiIC4/f+kE+NBDBuc
pnphE6+uN0mEqdc33HxnkFOLulZL5MGgFLgW+xeJMuxjFTnGuff33QOk6fQnCsZj+BQmVJNnDO4j
3lIjb28MAklKrMKkLrWZqRTGDVBx1tTUpFL0Iv6Yxo3yaR4XHoBcz9NnYwYq5cK0cTgrexkuX2E+
MeLCUUZB/GdxMVOnIbv8wQahbd+8CNpLTrqtlG3VuGuYUwo2y0Bhvnef3ZHQJRRT0IH+NaG1OByS
1TqbIorJAoYhofVtbAH5UfzdK8AObloVBMSolFlulTft+FgVC9s9fvRyeDpcAf3GHiHaH8eJ7QaT
lsFFFR+nVElJ7t0leOOCTwyhLTggy3CCOrISWudI/wlVzPM8TjZ9+hax5vX7UXpBSjDYjQJ7QQ70
QIAVVWVvzK8tO5pFQeoLfQ/PMKcvCv92oRYNj3NbateOI51MQ6hz2NFH23KNY066p0pMzIyN9XSO
O1K4CegUXpj4B0VjLFYlX3JNqfTrPSbq27jqfGEB5r9Ztej5Y1ukhBdeXLNsyOQeUZqyvIv0R/HV
2MmqAUVnECokU8uU9xWOXSx8zLKwCLNBfqV8Xx+dlXX7fNUUMDcaB589XEaNAs58WDlNs/gOtc27
cnPBBjgZuRLP26bUkh44dSVSnNCZP5lmnZMHSh9TgazMXpFWKCB2cwHKbyUwBvRbLo9xtdJR1sxU
dUAk3UmtXw+J9S/Uu9jZvCv0RqrXJ0CshFlmEcjY94dISlD5rZg8Z6sNTMO5Bltc37B+isYbcarz
FwkjxrTlxNF3W1hl66huTProcPjSEbH4erm+dNXixwJvbZhxxYvIwGbaQbV24zgjERK21xz2KRNl
F40WiVWeFpEPVt5wJ4G3yxh14C4IHaxOYM2JO8qnv2P0Wtkbee06g2Gkb959Pop0Nb3m3tNbPlc8
HdBiR28j34FO6kg9SoS5ak5Z246vt4OHbF+cCnYvI3V8qoLWvyuW6d98gZgDjGxyi5koGssQ/7P0
0zJnpo2PfoDIqjyyETT+GSRkE4JdTJyYacGboBh+54aQXhfi6/ubes5FBbIjUhpXFzEvwwWIaGP+
kTTVPIO5v+k6+46IVEchIJHDRxveKIKOg4Nh0PXQxChU2RMoUfSF1hiASKN9cAtXkft2iaBurQy0
Q9ZDAj5rpDhZszUE0kOgir4ZFXOP30Yyzezogv9jfovdBUVhV9wvlzgcXz7xTYyAFJTeY8i0Y+sZ
eWmNt2iz+mo8YcwH5tyiLSm3tmK+pxJyJGSpC1pGnUwze3YZEz9iog9WHYo2MXcGPVIVpMaKGpxG
4gTS2Ul0KN3rGoP7SplQIbzyK0xmDNiRTH7/+5lhbgULn7sETdrc+dgkNDXEZv4gXK7mbpi0s1TS
K97N8WU8nXQ7bZzLpgY+vNgOEUT7MxjoYZ34W6fTUoAL5RLYtsz7vc7Rv31zUvo1J5QI09zJGBHw
VFZXqnOUDsI/joiQZvydTd0v0Cr2aHgJoBlrdrovlv7DatSVqwIJCgCrNHs9sXBk336xAJRkX4nT
vzaPMXEwqotHlnfO4gccVqBhdPomK3RDyRK3u6OxSyAdiGBZIBLjwanG9QZ2PCKwu+tyjilOBbon
Z44V7cUneLBChB22lMMusxHHmjjePKHfnsTlzD3tMoffjKx54TcYntsotZCpgqA/jQxkk6cTK8bK
HqpYo0WapiWL/hvWE0n9Ob13I4GrDZ5H0mZYUUZ1F+RLAq5/qGysFlBBMPEe7Ip0TAaTb0K+xVSl
OJhThTY3dQbYmdSCldYsNifhAh0qyZqfpJWDk82Y8lrmXsu5OHuxeOViX+lyAmcCkuv4K+Pm6pYn
ZhVXzAF+fmeyYhHf7YztXKWbHWBxWgO8+ftHRb8OL/f00BwqiICDtQhRArCDrF3Ye+ey40J/SOm+
k64K79rNkMuTIVHaDuSOiPxWn6S8l+ueNYtBV5JgwDG7vEUFaw2SaHkXyDpaJ7rmwJxOiWeqfY+u
kJrIMMvT8OrNPtyb2XFeE0JWminsTonCdKWB/1/QWjbJ8fkArgGTH/6g5Y9pEU8eF/zOunzbvJub
Jf/ayY6c1PVq371EB72hdln7xSwlaOIyuJTiLjvfzuHkamvHMfLuPDXT1IbY3UtD8IbokmKla4u9
TsmvjjJ8IZf6UBXAMN/PASjVWkqnmUGZct08ntwLnu0xLM0YcSR0H6bBnDDzHScKx4xVdUX2eCnW
46FDyYP+EKYa9unm9bXSkzlc5wLZ5oBvjmB+Vlw3hjMEbuu7Ee0Ef6ns8UfcGOH1KhTfm0yIX9+W
ne+jl/ShkYyDesSgntA7YsCJ2saEdDws1osgmlpvXRv1EQ7S0qRxVTwd0tjdczHQWQrFOSGyhCGS
En+TFcbTu2PaY9h0kRxldrQP69CD54CEAMax5sSo/7jSkp4iJoMScRfS0VJQjFAMc/rmPpACY7u2
+FNFBrrEWY8mg6vFpA1wPYM3XZfsXPc69nWic8/3InE1giRP7s8i28TbYlDFMNAF1toLGM0xdWa6
McKhGx5lhHL0W68RIoyY2Q/lc5Tgh8FUQrzm04Q8ENCh/rHnkJ1FTVEnVj0R3/UBWNDOc4BcuI0M
ENqDAOHp3vTjVGkpvadEmoONlzeveP6H75tTYmd8L/FVKMVAYAKZ1zwFRIM5OBpsC5QpwgwyBEUY
F+xv5H6iKjUGeKM5lnoLcfnDn7p94ffusid9dnm0rDw8xsqMZdceiJkHshi96uq7Ml+nd65na5sQ
8KJBSLOmlqHR0Mf2Gc19dHX6L/uvHI3FLyJ2n1zH7xy4cBVRckMJ521tjiqnF4waCR0D1UqOJgfg
GHvCHAyhbMT/XK4gtB2AZgzhD2Wyps7+6BfhMySVcKbUuWU9YpyHKELCkaHUea4ewF86suKH0PFK
Sh+54IujGdRy2g7zXAp9vaPJKykLaF8Z+xRP2a8Elum0nhOcRnmdusONoGofiS7ogtvbpTlM2DHD
3WSuuBS48gSk2ufNbrG879xrhs9W04OGYkdXDqpVC1JA+EO5ydWfaFSKxbezgQySsh8LmDqG297j
TxzUyZfC5MAs5zheXAeTFTsnEiu7ayo9SCf7KaFykjw20H/HmdlZEY2m0kEUp6F5WlGMvw2/1eMS
mL8WY2ZcYZYXSjyNWDhby3sgoQ6P0/6uUDrdjE8N3JiZlI4Iir2T0oLerDcmGeIJP2fTFzJnzxEV
mDx/Rr/tWORHhmmtRqkN3+iXtfyKwiQaE+6HIqF1EnSdKaTeAtexcvNAATJ2BB1iND3UmC97xeA/
/SGW1fqHb2zRmZ1OL7xleNnDhMG1+gc/WXEKFMUB5NEs5M0N2RE0X/T7mCjUMl8dcYGd/fRB+6bT
lrE2trnPHq/aN/tTn/2nWSkq6hwn/7MRDuO6DrfuMDN7cAOoIi5bpOsSzZv/yMWiHOeSyP0+j7Hm
e2kt4lKfgEwY0Yb+aSLTYzL12gCEzOO9Hdo1LyeXSvWmKQXsJARt/n5DNHHKVR34QnH91k9QvPTg
Ri5/wlt5Xnuveo0BGvHBVzg4D5WZUnOWbU0zxVnwGjuUCM21HRNH4I1UWG2xEkj9JGxIowaIdKSx
E8S2NoS47ZSSEGM0/TafdP/ItBu30dGqND+QtrstkoaQL99GtzRP5Y3xjsZ+KZVes6XoHD/zY+xs
QpEzKm/SQFA2y2CfVYzC2GMK5GBHATDe/w9tlotGspQaZNmhOa8P/XhgNECFHWzcOKb9ZynNb9Mq
x3jiI1aN1Temx4RrZ6GwZjQL234FCOSIKcFimwkYouLYyKkyh8xITABwwbbYdBT51Fplh65yHlPF
r/VDOZR4BvTrZZdcoLWXycNtmoCjR/gahh1a4rvHfQlIVP3EIe81uRq/xUbnZItAfwm1kaDHMOL0
CapeZl8S1jHanSNnZWTCdIrzLzGeIRjEYWlgVbUYqFHfSd9qcy31+QgdMRCxs+tIMqqp75TUCHaj
iYRAYNrUlrWaPCxHcEZfH7snXaxTEx7uUAVkznuABGoyuwlyxJy1p1d4aFJQ9bta4muLFn3aKATG
rEEWbhAy0JGrLt2Gw9OrjMJnIn2wUtswsva4z4LiitoxUvGoHdOBKtjd2h/6VBlll7bVl9XWWFln
42BEMyYgHySpSQ1g2lUs/zjiTRB2niLzspwAeXr2rqiYu8jC3EWgxTN010v9p04PXXOjKXuGxN9V
qUZqf9VTL9BAZ7JdOBfE05ztLsFu2ckIhB0H/s95Pfqez/NMcriVjwsdsCxSqZx5LK5JzfmXpMBR
ZHxpIZxZ0z7gKJnRqawyZQoG4klnX6CiIPGjQb6BrhhIiM4ysZNGmQDDZfEpRFYqgpuetvkhKsfx
Hb2VDwhdblsrWu+0Pn15oPfgOY+KPmX9anBCETP3w7qo8/cyvHYu+ljFFlwS5+q3Gsq6ZcBUDS8L
mPyq3yzMgcajRNu5irkcDmoQBtniNogepJd9aOdX5Vj5bvzFJfXbAS0wKFpwyX53aH7JfVn97fBN
F+1TtizS6lwQfiEyD1wI0rn1ikWpb+E5oNuMwiO2MpaXSTv+Hx+VoOrB29U6IS2ZN5af2fQXyIRK
yB8ZUzXmzwP0TcVwlJyv47vPdKmclr5I4134lhN8tlZUYYo4XywEkku80PbBnoq3JFuvp5A16a2A
LtdFu7dvscwuIK3Yzasz8e9aRyVCiFox7oLFYxEZZ+pQwE5ZKSxaMuM0+QFqtPcNNl8Js1/l44V9
vLAL2no5PxOrM9MtQoaoTNtoOnujkJhvo0S29zHoBPJOHDnUC+icKpzWe4YbO8lUDTFAgN/JCsZA
mct/o+GSnjDPN9Wc8VWA8z1y/uyip9MuXH/8GgeFP9psi7rlwir/UEasyi53e8EUQuW4+zJNQR7N
4+XI+KrIYGSE33F37DPwacKAoj04S9vrg0CyOVYk9OSSAuxAi5ANCjbuGMlPqhTtUknxZ9VrAfaU
UgDbmd6GL03Qfx3VH5BtRUiBgXUvveUy4cKENiV/BerwVWSCW3ilCLWyKrKFzwyDEp8uH6b5hhKT
UYnPiiSM42ycFJnRuNrLDruDNLrk2bNzvb1+5oeElxjSmwwkQv+TtfxrcGoGOSDOx43OuAn5IBAm
NVK3maPReooqBqeKDZ6m+DAVR0bYO22mlmYd5r80TrEU6pXwcffWYP15eDvGApj5mOAFnh/qAYl5
NbtX0p+jS2C3y6oIUR+ZmQbJ5jUKDeytRnrZc8o7JVsAplqcwq1yM57VzK9VilNh2blerFvnJY3E
EKpZu9xQjWDRiNcBeKKhJz0r55gjXrEL7bxbXeAv4cogIXLvyU4R8cjH771HDTS/Bzg/vmaD+tPr
TmL4FfWEzudhmCo/IxXUA1WjJD1ekqvo4Kvm/OMn2xdNuOUXJo+6Iw/FgUWPbpSbb95dYLjprYKa
/zLMV+S4h1/Qfq0suqumZ9cAVIadIRfudBDZAIt7U3C7ucKzV6oeWQIZxrZCOTxKf3tXt1RskZ1E
HHmWcG/zWkfjRVhFfKcFLsOdxK4Y4RzGua2kg3oopXXq/RDcY5b9F+34liNivoJ0VvQYfLIPQlow
URzhXRnVsVuuEDwsArHfspCXqyztzdAwwpJ/hqSdq8qSd8r3BthuRp5iy9buFZIXoZuH3rzIkVHp
0fs4FCq8T7dElYRBbGPyybwv9uogJ53S2alpvTdD1nI/VfU+c+7O3vxUU5BANOyNGHAPKShCkYrr
pLumw9TdMoT9AAhtHrrxIhbFzIIzMGT1ZaLYl+wLuCQaVXjYThRavqDklpMVDj4LT8cLPaa6x3dn
43sJTFpG5G6hdSJVc+FfIrqKb/63AvRxQUZySZpBcVFP543o50pwpRnzZPcsXiO1s1TpnvUaQ3se
0LD/q2RK3BChPBCnzKghLxsKbxtSVqKtOio3pmzw3g6AsAWQWTe3ky4LzPqpKuYsSFUFgMyR0YT2
dnTegfO+r7Mnbg8BC/8b9mnExLuiciD/gCfcByHd8Veu+yIv5hH03Le6XSh9OxLuR/AuS4jnrFRj
90Ng8BJ7i0YCtuRFFYQ64g7NTi0dgd42Uo6SYKLPCoFgIndHvRxIg97gUrp4r/aMbn+lfAi/8O/x
AYe+KyHr0SKG08pPjleDHoqBH/XuR9IyPT8WR8ArCR00i4mJKseLTvayxfvRtI4/9pAa9c/4QSAg
p/IBXGgsOun6HVa4ooF5w/zZYxGGiVAWClHhgsaA3MWUQmaws7jDFE6W5yqvSrLSFGro/z1lP7vb
NtSOhZz4CSBQM5MSURQRY+ulfFv5oQatb/Qba9wygAI7qUX739rDLNaEcGIhT+WBFA/vBPBK7cRK
BPYkd0VntMrkwiqysT1Vso3mr2tdzcEuwLM9z5xMTS7WAOIjid1lrdgdsg7UybvKGfcJ0gipVbcr
jzQhh58jmRnLH2U9Q7tVShAyxvg/FLqtOo+piRenVs/8X2N7bMXdXZbx7QSKOSuv10rfEWiRbgqu
776FBilT9OSntdBrwTdpwNKMnSsA3M9+cjeHFqy5DG8E/m2IxABttdJeWCs2pnM00L+9VqUHQ67i
fD0Op1JG+7eerXN8vQcqOH5fJ/7R3oYMvdjdlMash9CBJ3NCQsqdqEG9H1lWRBZrfZZtdfTc95A1
aMQqhokp/yeDUsTUy2tFedxoPx6UeoP9esxAlCK7I9LZ5Zo7Sf4c+aTeYO+o4PG7iibKenmiKhct
3fd/6PJiFotCU+WfTrwMBy1NS4DsLA1IPZ79HhC6mmYSjYngXOUPBnGPqusCVUuvb7QPUKDteAVO
QQOMtJWHgIOzngoJOeKqC8thVZ2xVBAzU5svdH/g5QT5ILgLEqaBD9E7wHt22h+kcwQ4+VwKWQ9S
strjz/vpYZDbXYk6qgFwOa8/WJdekUOUHh0iJMvRki0lyUy27hABQ9B3CEuhkRcgmx28kNoqxICZ
sSK3ojIIYxsFNIyf51rUdJCQAmQRmoeUlxz06CNNJbOTVgWteFgra79nKXQnVNvxbQy70IpCnj+o
fvRzthxlcGBOQV0S+NvPWMdfUrzUeVy78xd2lUEWi7ztfSyDhN7qm/cO+eUVr6mTzvuxYQdTARrp
z/OkZacB8z4ZmuHdjFz52HT+AxvbYP/oTB4m+/FMsNDbNnk/quPm4UyEePpGGoouhovGXv3nu0+8
xKybAD58GxivpFExKKG68I0N/uzjbYNskF4S6oibLJgG0OM2siVDk8ntA+QKJIg5poNLo4NeF7AV
rhXFIhntAGD9pe2jukG4hHxrl5RKnX6kwPp5snSEbS6aRN8NGn/RYkUpeeFDKx+STWYmTS4eHxAo
wjw86cUhlkMN09dlQJiRdI3qEfLRURaRPBlo4jBb1GgIpMq48DAGhVXEHhrxOXllWSJltYbc1QcK
N3M55HQOWibqkMmqhjtSOQqLV6uLYtEMT2LPgxbVjsOAQM3sUDmHMEQ/4QZsoVqoGFsmEN73ZJ4V
RXz2f36cNwC125GlxcIwyblzBcXMyGjNQFcgHTZTDESXwzej3ZwRcGwxzGNsx6/Xzvge777+tIhY
AeQBephAahuiB+ik/KPd2o7Y40Imd0BYZzZpzhQG/COTUnCOs5ZfBbG/S40h/AXIZZYKygHA/8yx
fkVDBrst+u1Rv7wwy4ohWCHGewJwI4/MzqbY7NXL4rQ+ezeMyeOvwTGWzJkvbjWA7krTEtOXdffQ
+7JgdITWfCXjbi3o8fcNUgtTZ7IlRLfmj5Djsg7oC3MyKC1IVxN5lG5TAGf+IuJEJLeMKwyflqhl
ycqvxeubepOnY8HnRxQn2DzilmNvQIBHAMbxIliEAfrlK/e8mdSLZFVo5BPZYAdOAOEJaFZDUgf6
N0A10gYK+12gsCbm7vTaL03rPMWevExS0NJLkdNrcbEt9JHX3IddnLn3at/wRDSdtPbL01Gln8z9
fn6QgZcOPTPV+FSGSvraa4AAPYeS/Ak6/X8C7Jy89IHh24zRfDXcnmi71ImBY6s4b6tYepRLFMum
j2dO+AWUne65wKsyhP2HfDAeBxdWzzAS/1GYmR0GmGOajijA4GwiQR6G71Q6ixd3s8eFVdg3BWpk
SbcK3xLCCn3bIoFKmLvhpEhPbunVQ+3XPe+MPpH7s8TyObzm0tOZyjgKyAJDn4Wrgbxm6OLCKPBV
wH2toXhfZXuvWnB5wU8NYZf7700sKkUIsy09IkPGjT/uJG7lbpyKnisXzivvkBSNRpFjaaRMHeYj
+GKlEcIrAJHgaL7FRmytMWu5UEz5d89GRTbSPCiOXZmXcl3g3QFH9Enq+8LqkM3BLOz3TfmcEcoA
BxI04gyKeI5EInxqpzXIe7PR1vl6KD5dxJmFn3jB9jcRsFpAUs9JN57/KU2yg+E1BuRCFmGgzNrE
qV8Yngt8ondlAvICOHy3okeyML0dp+N9R7PzumhBmMZgZFFFSAHY+BSKfkRWj08/RbyD+6vWdRRz
fO3atKk5MXJJQgO95RMYdbGQrnvPNo0mZfUB70OfJwjmutpQ8KFWJgpk+O21PAZ22xr22rA5/X1e
vOhX1/0OB3DKqGMAD90zSrWnqn1Cy7rJpO9C2ADtOdDdRdaQqmlLmrsyeT4MqGS3HlrRf39kwyDl
qRJSxKFegJXpIullrtn1hXX2mF0HKfJppfQ4Acn5eJsZpSzPMWinufZojBkktI6Dtx8qSwDXqEPr
xO1r1GlTHPtzFRVDoOmEwe25YNbH8I1uIOCMdWtE5WxDjrpia95CwhIwkZMSDqzVmKEofVjAeVIc
ETT+znMXr3956rBHOgqKw1eedieCWR0awS0QLBHmwGPdnEPhwpwXuGJDjFiOMElt47ihNzCLbawl
Msh71Ly2sISVlfuxvtjyiRVIr83hIaDVQrVpLqXjqRBWcpQHf60iSH006e1D+vYvHEM4oXYz7wh1
CItRBi6p23XVn3wJMuajajcvjrKm8kvr3pFX9/UFXcdwToYrNw+qvcYMeGzw0qaxLcYd3hRt/+vo
FIdO8T0yZ7/t2EcoNw864k4kOpFojT9nuzsIAgrQRUxtro1G6haWMyArVVnexHJszADh/G+yC7kD
NUJRv9FhP7ADBPJdYad8dEJ0p2ZVImy8U2cBCmt4gzM2riKRiQJ8KKLkqPCgmCaQQxX8y1vMft3Q
kwiy7hWg+c60YsQW5odRngexyfspxBcpM67gaZ3v+YdL0yxyNt4/VPFABA51XsveKEVFDOPPsYPs
Y0dhhmzY5loIVBCRTgmwmqx7l933SPBtroH5E/ES2C54ef2NpQVi4z9kG/L7YIND5US3sMensfEq
iYp6S0AP64jnXY6c8ch7Jsf0PuMlhu7gynMXxcd4ZheQYMzkJbCZeiyahTPu5aY4BWHE73FlY+S2
WLBFVJtUCkPEgfZpo7B09nbsAsEqn1KK4HQe8Xcf+uVLqul5hF7/qP94/TcO2s6U3hvfhhBgCdgO
Kz0faqDStqtVS6FGsHx+bmovtIEQmuSCe+FQEnxI2wZbo0bgyomFClJz83qSd8ypT3aFqhIFW70u
fMJ+vnwnLuPkllqutqWh5lLeOBnNpVT8bXDDMpk6RY5zMt6+RiFPOjjHPBFXD4c/SE+IkFFZGO32
twPq3z8eaB1k4lGv2dTjrqyRMyzFcLkAEhokgWUf0YMvQAgQAE4V8D8iSdQ5pLCjGhyz74anNF32
OnVVEb9kY8Ks1vjihq+gmqEwz2OtVX3Wk3IlAMdpzWTXGzFNsoLdnYBeBo70a9BeAe1BOxl71toy
J54gWyrw1FrRJS5t/l0Q6/VBDJ+k9H8uUBjgmycB2rXI42h0Iwq82/Eg0H3MlJf8u4tbil1OGhG8
PZFlspz2JLzEebL6aQnN4MeoKo3mWISU+DG7SjnuojHeFAB/K2TsLSbTYqyZZlYOf6eHpBjou5YJ
OaldeocjiQfNzsZ6UxyimUbRNbxG0Q50i3MUg3uZEsg78aQ8D7+LhapDrfNLPp85EFMgjEd3TM5b
mYYZqD3W0UHIHRDhnsjwDcky7uCtwKaaCXNDOVk4CC+P3zhbpVH+rqUdV1IYrYBEe6yYePFUw17i
az3IdMbkc9LfWMOqNPVsoxGpB8KtrZaVfGQM6JfPODWlBwpx0nLzTlr/ifQVJChAZHGFl+Vth7V2
Bo2yLuCCSkQRYpOxkp8Jig/UN9Pq/FMWAaA/FZ+8bt1MLUOCc3Nd011A+s0HRcyhJspbEMDb5piZ
P+dWn+kx/FOdnvPtaY/hPOzfeyqm42b59UlF81W/4i6EpbtmtUBLNpxszKWYgcNMpXztgax7bTnS
K0v/e6R3yFqU1G0wQNU1ljnv90EeKsZ8f/Pi+MlhcrHDGIHBKYkmL3os9kCgxKij4RO8BZdlc8XD
uzQbxxUlMsV3s+ILserPtf7PIbGeHhsL4HXt1eoLKjYtTpVOqa4SLpXUVMKi/fvrBJLXmkQM3ICT
5XZH3Ly413Rsj+VHytbK5LtUh6TnOkEi4OYLiyRRbbdoXf93o2U4FZ7ZQJljpr/DQkmGeCBshrfJ
GOM3DBDJXRgAIhrgSGy5a+d8Z7T/SCWL5q8vaB/LQan/a/DasIy62IO3+7uTZZghFKY5fPmgcOiC
ulWtzP3mw9etK65wTzviR9LmTS8WwGkdGNbbJHCvbC+dIP2dTY5ao+r9UVQGRTgTfcoY7McrPluF
PojDPTQC/a9bOXQ3weEPOIzscpA4ppDmDLaZ2zFBDgtiOVP3UgfcVy42t294dFPYUQmbMKbLfrHr
hSfPJbVlqsf0u80n8CWu7ecYR8GmH8WMEsGKP08vaWQAhW+DzJPsHE5T8xYRorhjd+s4z0Sdem4k
+/7d0Tx+Jjv/b5zbz0r1BVrJVLEvkzrwDkn985QJhP9FA9BIb776K9/fmaNplDsOrYSIw/NQxA2u
noAIi6bDi0dBdleA8Q2OhuAvuayTDL8oRddr11r9nHcdSL8RoVdnu893/UKcmlkN+S4YXGUNavzy
KmGlapgKPI3Ep4+NVNQhdOf5b4GMguXXI9cdjZXiH+lA57SMV98bZssYmzE7rZhMDWOxaOkGm4xJ
Y3Vspz2LLa/q7K6Rplk00tM5LqYdfURvBLJxXRqWEh2BDbdB1nVN3A6Q91T6g2yQ+q+qKybLHUK7
vdhMpk5mhGwi2cb7td5E2ASU5dzXyVy9RQG/TSCT13xcyp0bdFhpLqU/Zb3ClQ3vQtmtrk38bhGZ
ZeJDSI3cUQKt4DjGHGGsootd0HoXYif1P5W/Jb1MFINaAFa1UaYEKgErBYr4Ss0yucD/k+eKC6Rv
aoO/REpu2rYorE5HyuBYRMNfuS/C3zQf4IXhthG6CVVGUilnzNwbQzKB3AgXTOvlgJxSF4xErgFT
mbJKgIUsbTh+5nzT+xV9lYY81QQVmlCWWefrbdn+HHiw2LHZHbC9nE0C0jsNND0agBxTqgOqGVYP
lVUp5m2ODyKjRtmDDBVk9To9PHe7ZY4VuabFLS0FkgXTpwnLhgznD1bAy23PfWTueNNR4nK7aZ6n
Ji3VGL3HfLj0tupxAN2U3QVfSvz1XRESM5l1ndY/sjhmhQLIJCAxpq3Wu+9GevTdEro6H5yuH0k9
nijQGowN/n6A914XGTV6am2fupqy8K4EPCfDxKGUuEYI35TcIMo3JFj1xciP1SlWZZDFRcZeZkN3
SmhodBaYMuHE+4mbAmAVOLU44/tLqvAND8iVO9vFdSiBhnagRxwfWPP+80y/V7/U3ndFDXm6V6N3
8B4htwgrg3TREV5y1fEVHlBVCoHP22ZKMkKauOcDdM+A4/eXdVC9Fj9NSPr+7z6L2z1BX9xJzKRF
j59izkPWEJPEBeL1/M9eU2a5UhrIFcJnXVepCQEnt17PZYDi8+EfxH0SUnOEMN4BOCINBvNMew7n
+5eL/YhwENsHWX3m1uknWqyrGeL68lxQfaSdU93gqS6ULJ67koYJ7VwOyGQG7qj8pviKdHnXr23k
fR7rDD8q408qQxt4V0TIl9x9Bg3U9PdaCkiu7oVA/UhcsODSuPnQH/7qq098BBpctYT++OTHLSEr
RmixclP3nyYK1D+V6XCeiFCV/K5E8TUe4qti9KD/r8/lR5BAHaih8Gjva9IWbYOprzpzO886xd9b
OJYANbD3JzEiCZLCbsT4TRV+7sTAjkVRsVrYrcgyflpcWt9qI9ZD01S8IQWLh5lfpJ4QVQUwaxOS
g02DGp6phmXJhSTmCOA4Nh6yAoPTQVxRSmSm/LJJdvlKzbp5EpEp3qquV1MYBJ+piml2BJses0Ex
bcvF59qHeFYz8I6gSOhKa5asVxVt3Axe3REJ6phFe5/uarHfLwktMe0fBUaChAXhzuVN0PqNB7W5
oFJGvdwEH+rkj1CDQxFP3V1sUsfwd0MRJsrLqL4WBdbNHvRoGVqRYATxtz+pSnjKyo0VW9bJIY8B
A7sQUpqCqpIMSiK/RtvCAkTf/Xhhs/iSuz/1gDC4r5EjXxiUNgvvosubw8aypSeA3JpcDg1RTlOB
rZXQmzdKrKhlSl5FRLTUcDe4V984R4VoWuuj5QDpuB3NFtKtbE+Z507KzqGYKRxMtwiwjEXcecG5
TsUAK3bjycBSOJxaRUf5m/8/B1BAJEe5NnxvPKbuZWZrOQP536NL0dyoa7AjKm7nbytAQpqXHT7+
OmuOWsUQk7kJEjvgHhJQjy9u34zFfHZTEULDt/h73aJ8mWpgbunbh1l/r3QY/O2db2ellNkBOugh
JRgGl4a3eT82Ie7Si8RVI5glmwc1uU07aAn6pjS8HXoircbFzOptengwZ4XrIOmuBfDsmO4zKoT+
oZ4XTZSC0Sr8sS85vJX6XbVF73geKWedROi7spHxLeqI4eUeQVoUd0MILN1wOHzwSp8596aDq+Nt
WciuMfh5Uosx6jZr8q58EIwaR6ygLZ+VqMuW3HqlwZ8ALfUbjTWRmJQnP2kZ8m9EZSJSHEobJ/9x
kJKv7L5zX0mWsfm9FUG1O07wAeOf5CcO9VmJpVLorywH34LCEpYPRs7Hkb+3lNf1fa7kBqkQeQS+
r6sg+unocpUF7dNmA4BHecFNPpd6LGoCARAFM3sRpiQ3Mtbsfr8BizK5v6RSIpt7vBU6L7txwAao
Ezzp2pwP7VoDM9vUDuHH8kWo36XttVBua1jMg3REnO446xSdBT4U9zjXHBzGVp7QbgFgjKIGMF2P
A8fYqWv6zb9JJbwO4iMw8Jv5S1DFIJyKkNxpHE9H2BnEflV5uy7NNXRQwMuG5RoqAZT/bTVtz3RX
G3UN9HGwsBjWV5IlyLX66Saz3nN1FWUvXIXyitu91Oi43kkwAUd7wuGuEiDnDiEcxeuuKLTqaSZt
RvaX/oAqke/m7vjKBN7XBC14S9sCmxkT69X1qMrJ9EO/nPI6cEjmhVYqwIvWPx3w4DujxRWVfmnT
x+/q0XoFndHViOiUQVLSUhsrnnJkkm06Ux6+tK5FnKayaVk0EChaqu+3UDxNd3tV67ujZmUgqR9k
fbnc1lrAOlVARJL6tHzRovf28+dJUCaFqaxWvvoJVnZNdWXAJ4vQbjGPZWbdb8XVMWxaiRHS18ie
jrCG+pV9S6qcDPSC0WD5n9r3m0jMn2UkSNqiPm5FiuwKAgj9QTSG20pGt9TYuYq7tJrQjKUntxUv
iwr/5+t+//1wgYt8UAecbDBi3oCjpQ80z3gtNMdIJ5xljA85Lts31RjiaTEwGC/afQJZrF3DqB7d
8jlF8dOQcBI7aR3pm7Ofmt9Bv21B0ABYIQmnqmGwWhlRhcFUvEAD/feJFFuWD6n+VzSz89Wig0I4
+W4/VrFR3T+amRRGfo3srfnx82N8gADXfWhgK/Bpl513YhPRZQNhGEgamg1CFjeWrZ7M44W1JnFt
AEOfksD3yWONDIGr7i5wU71uvQA7t0Blb1/v8I53uEd7EmmiNMMlbiJOGvfls+5J6izHR3jD66uf
WzJjthQEUVdE0Y/thPifT4Qan6hhA0TvrvZ+tfcxyp/YEDIlREmZbY27mAxbx44cigEUMQ70fesW
U6HHT95pEbIKWYLAONArnmRHt6g17osAd6pyL5OFXyPjNenclfQw0y2MKgrk5vhI6GG0jpdRyNCb
QAl5N4ii1uWrdQwbiEf2iEU5Dse0FFfMURcCcr9jyyveg+gKcF/hZ1aZOwC174MAkbQY4513S64N
Z4SP6SOUuGUmDohcEP75kU4mNhd3FerLfKf0EXfpbsCY5GQNljyZUrFBy/kIBCpWIJfAmuYV5VfO
vGmCQjLZqzw/u+PbOEaUm/opv6aYbjPm3SHdDTH/oI0cjRnFrMVheQqffGIsnA4sd8KvucHpy7CU
7qiMcQjKBS62iHbGPW6RYrD0qhB0nm8O0aswYd25hkSq2fD6/EaN27tuNf+yVPs3yP0veDxuZq7R
uXIFFKQF1JecIu3t+pfhvY99SvK0e93HyQ5mKC8Vs2I4GKEQKK37YnaU7+Mcz0uRs8v8lPc658VY
0g6ckuwi64OblJj6xt14L+v+F3NL6XqCiQWBtINRFEVe2pUD5RQ10ADTiXhr1iKGbtxrWjLJIc/5
RooA4jdcGVYuT/MqrS8Jd9nP3Cp9xWr/T1UEUESPhT/n8vb/PG63BgNW6/62DpeP/V+vPHF3ZWeA
R3lXbTrvvZrPHKEDIIppFuXktfmlU/SxmjSDjaYrwJlyDbHtOosgiFJVx+UZxy4xj3sL7pNPftwx
2Ox8yShGufv1HPRbwTwzruKtwQlZJoy2dPJ3HXrtmdxgiypq5Va1e8DSDGKy5elB4SJ1yec4Bpgr
qp1mLMpTaXtz4CAom2nbNvn1Ddqupv3oAEE+bnMYSv9jN35or4VMqylapDvzocfXjGTmMncdsmWg
cj+LOhUqE0+GF3JvvCMgZWz3CHB4Llwb4JRK0R9OycNnDe3HB6kapCij9sV0nePpER/v0+YwitwK
wCJYfVkWjlMy0Mux5fNODU0B5FS+4Jw1ah17C3b4CPl1rlxmMPKfBSL7q7VhQEU0doo3rrCguz1F
lQRtkZGhF1bn+T1d24iuhnG9uIi/auOmxM5RgU5bSw+5eoixLQIUse8uf3d85/4MoGkZNzboU389
zdvOtU2Eu72XqdlZ4/IOa0Q1tzigOr/dUsSjG1fOtMd85vCFAbomQm/jPnwdPp2gKYmZfcUe7V/t
HG62bB/1wL6TUYv+Rsalk0KEKSLTkUXmCH+A23dVht9TlAvhELNcjRtxq7R+UQmOzTjHu2AisKl+
0vKVTP4XmbDwDjF2ynjN1caDUWoptugFzegrRhY0QGfcWSOFh/AOL7kVSo+Y9SL8Sgfy5KIu1dY4
j8iyHwLTp/k4S8jxIDyGma0ZlKMNZNLWCEh4SOr8iA7PPY+zPDwnY2mdhcpayNP0a0foRutz51pD
Xw2Y3coL/wk3bUPz82f22mJBj6qjIucszJWSouf6aY3uIJJlOSF5R/sfahuJDdR9BP7v8G2cz3tj
02LweLow5F11BgFnJEzCYhv1EaGoA5U6B7KZyM8oWaJnFi9jXwlrsitSxCmJMQ7Wbdcp7opKxYtc
nKkoEu2JHfrGN4XPG0byB19k/uIUqWMMzMbuydFR3vdvHr5ZdkdmBg15bOtpTOY7ERZL0zpEDOlR
w2nTGDQPo4V4lo/s+cmrAo44SOjjrNh1BYJdJb4a3RUXjRZWy1tJiqgYfPaBYNGY7vblXTEWOi+d
dI0gXM+hshru/J9C30hT7NqftQlulQhFhYHmsv9KnqHyIdcbQJ2wuwnnBAlQlyggwOMDUrpP2XVa
H+jizmMbgE5KjdF4A0BcWBuTJ3HZk/tnKdglbSz/lFs+aaskS7joXkzp2C2QgDjUXnPhxjyHkoVX
ANAFtxYPKc0Xgxd6kmJBj3cPxVVD+LHkhIOGm4+vBnhQEMkb20pxolAy+X7YBbWmD/LPCLUsN43n
yJvcVUFLml2M0Q9TqxmExJkwuBX/F2PnV8ommspfD9V3Md3Z44dGk27gUWAUsmIz3019e66Rg+gz
FALlG9rwC6AJ2dhIuQO/5tXbz9ppnm3dvjVqZ69HeTp9U+l6bUn+719Dkt2RvxmbfZZGh+fxLyjw
FExlwW3sotS1yTNJCvO6YNTXIGiPXJITUdayNCGghrTmTTRlWAyEXGzkl3wSU866KpaMjqgcOrx3
lpzO7H+cn9QBZ1mAhqIe10BYdm+e+UwByJFKsa8oeSwM+Z8UZ3Bz0F2+PAzut7Yt5XXC9qTw72uw
2Dc9NT1trT4anjyzY6F9MHiidtTYLdSGI63Z0VAm1RoczVLvBV5/DllZfrMpeeuQTp3Fp3qvpjIC
iAcRve6FHGusKbgRGXOVdjrbLsrfhzL/BITifA2nWBnJzRIXTxVXwdDmNZSfkMXFA6wdEXHwOepj
SRCBsm6hf4VIpZbgwXSdMhUvAWeyzMvDqx5qrAeyizOV1m5aoIF8XuRoG0vHoXMoye3xC8lYOb+B
eojREnpg9Chb5bw9vpiqTbKKIcQ9/XIkQYlptwb+J1KHxnFmPB1o/ZSYLK0qIxBf5SAAmEihPgPT
+lT6DjMKb7iTAquQpFIgJTI0XpI0NsO1r5i2NR66hhpGxqGxryiAGlXiUsnL5MN1JeEIRqD1oL26
+TRdPQ97ZOSAm/vv4bTPoC7jHnSvx2/CTF+Sk7hNU00bGJT2HgVTa8HDrCSu8FKQE+VY02EKg6yb
gah0WKSGdrhQBrL1xgoE6Oa7JBSJqVWkGsV7N8eTKmd+qm0iwofWOl+d4VX0Ooia6r1Osuny+rKk
pGhK3zOFG/7tz62eZOiOf653C/Ct/UdPvPuwaR8jg9YYyHjGCokVdxEIF8cqsSA75nK8r4OS0yJs
LbGVRbhEWyQyM+bQMVzHYPVzF/4fxSs4ZIx3JJyvfr8CB1e0z3J5VxFO9z0qVfkMTsWkNhNh9bg/
39aS+QM0OTmO9jBgiQoDPevVtvc42GZyOB7j5+5wF58MIhsqenQTAJWMUl9+SLhjfqfsTaAtNZpU
qyXmsqHQm+1rDVMugERQ1hUc5rt/SgClrGg7PwF9NyJjXIBWj4yl0L5nB2z65BnrvWdVd/nf4w9s
PlGGNSWEcsHu7QoTErqgUMDUvioNwotUKIOEloqGVmm5SVzVp7InobG2ZvsLUzx72MBvWQVq9nPp
GfHM89Px1AANJw5VO+tg4dABIfmseDtlfMQqx2W6bJC4RUsQROy36s5UhAANO2J5DJyGPgmAQqL3
v+HDLLFjD72fJqgWnwD4hu93G1lcEDUO1MwDS5CCYKoDVt1acrz5dgYmrH1BR7QoF+mHXsWVlYRf
FgshMzNdv5Tu5llW52wpNaWGXVxR/Pzu6BrxYhaCpleDJ4NbOs3nQH/RSsDFi8eKkJDTMB9iJ11B
UpsbR23uTtlIUIoF4FPJ0m0P3Cj4ebLaoy662g94zx9m8nwns3vMakkctIh5pia2fE6a20vjQVos
Yd0wkgru3leUDXJ3jcLmW5uf68NYsUhv0pak1f4Kz7DzgUWZUrhSoY43uSkpGZLQ9KxOGTXGC9Bz
46B2woEnXH1Up1Nrhs9mIX8IsZXid3lDGUCpjtsa6g4Xy5B8iLvdkqESyhhLBmlD2ND9cqBJhCFi
KTX69etRQyedAjfjphRPJqn/JGzBuC3VprQRWbMrxPShm2Zptqr80eEYV09WBpWoXQHqgsWNzlec
N5Gcbc12G+iZ9PwRNXsJVvEAnVbZyIspTP4T1wVdl/OBan3gLyFeB+4TlB7s35Vf5UTtwFhIHSdl
z21nIVXIW7JXTkn0KHAZMX92kJ8qAxZpWRa7qo+/EYQOQ9XpT1heJMTuGz+U2Qosf814/hevMqFv
h7nzQycA8itwmlYQ8MQx2QIyRQNvwetPK1mZmQML6rPEt7nB76nXf9MVASa6mjVr7Avy4bZ8QuXZ
Geu6j0RVbbHcdmsAMBvOGKs+ekkCBeWWkHWez5FbnmvfOT5LAi8qPMgQpZj2urpspGC5Ee7RHlvO
NFolWZLkaCdSfv7w5zPoS0JoR9k0toZd1uK0b/Vybzo/34pQCaOvVTS8XJqDj25UJa2QDuHt3vnA
vA1DMYbvMZT7cKcocXgME6mbYNgTDSyz3oTOcpO5DDfrpuolwxfhs6q4IJELVi+dmZ/h6q1Me01z
1syHRqu1n/lMnxFhVLM8pOPpepAU3NMrXDg4aQhddXSsSkzHOeRXrt+rRD6BBMVVqOPDDh1GWs+v
7WFGCdbAeKF8Pbnud2vktKzQ3e6i1mbhsdODIYyN7rz9u4MdzWjtB7yBLDcmQnZrneojOXgVK2yP
WXz5oxOsczFWEY1wDRb4rYLpFa09OKmIS/5Fvm2b4wktkmfBFm+9YP7hm7vUSofXyOUW7tVHmJlM
3vXHw9lx2WMepDymM+jEtSMD179E3dYxnQrcBELxO2ahHjlwgg8e+RE2iwXng2z1t4IIVLRx5XtR
xt1B/5JX5uCvmRzI2jH5YsyrqOhv+OSn0UMSFudMm9N8NmpQbCkjn0pa1ZgzvnALOGVUlhEvJKYg
lh8U9ecVI4s4LBgM2tpXNt/DO0aYuNaT1HxEAS3Akj9xl8a38CLDcDrZK0x5KrZvVaIHcAtx6yfO
GX1KSliwy4fyn/e1I0Ct0cKpf1+dmvMGRkJK/o8t5l1orNkbwC+/vjSVszpzaywNi2aVOgtkTiLw
A6NRGRhXOsaVMbz/m31ZlDMuYiPaN7o9bpmveoxafFIvkqUgtgEQwiI+NHmmjSIqy6HAh8rx6tr4
R/iokS3Lj0SnmHSDFUJvGsjNnspK0QZ/i+MRFs7R6tFa/GIKAna+Zh+joFG3Pd0qKQxPsR1FNezi
lVgMR8cX2jsuXmzjE9M5F5pZ10kc7XfNse5boIDiMAwPF5O12YDVkkCJzc+giBVDc3PVvIgf1+I9
Uo2Whop1DGonvjKhuCY5tLfi6tQTSqBD2NgezM1RxsVdhe73fjoEilKH3AJTifU4siX+Md3QNm1Q
mm1HZ/JDE5UwGMf2rKIuFcklmWma7QetRW1AitXJgKU+nsEm4kpTLEEs4xUCYoVsDmVmIt5UrQuN
+TTu254QTLPqdbqQWVCbNpI9ne/ITB97DHuj57OEAZlZBuc3T55OncRtB9h7W95n+90Wegctn4Kx
KNqOtMIBytxSfgoRBC+m8QTbBrH0pB9nUQOASg+9YdnhAS1nBsCL5HXSisjIfl7MMnkimBdYZnYT
/CGv2Cgd2HrbT7mYJTZK4cU0OoZ1EiNfsJGwLMr1L8DAlpfMfgTThghCJQ3llGUUhyjOPEiDFOd0
UahgyGSBbj3nkU6GvdbRQEwpSRgoNylWEZVAD3Yj3RrMppmd6sG8fnYUCAytZMp48891KkYGG38h
ahg9l0+c+GqIsOOlRc7GhI/YWwZGRs4MEaSa7epB2pKqUw6WfRhSQEe+9sKJin3jjGCcRLafQMIl
qye8hYeX1ncjOvuvyjWRUxlyY1KLmRjv/J8kqhfGOkAmVepMb/Z5M6JLtvziibnd6aQYVSjAZ4rX
usFqGKfkGIcUW/LbLmZztaN4c59bHGCyK+X7DveEsF38DJGBQl9YuV0OujC6bZoP/zDwr58/WrBX
D9BAShZu4EtdnUXnRiqz4e/Zm9hccYRK66sfWjoZuIlagMsUYiEEiEBWNAiUCdVg6CPW/u1ZQRd1
LrvaArYAdgzAOkW3OHPOnqwslM0NBAsRyViJVXiAqKqpEN6+F7I8rY72B4rle+kvobKqVY8PsgYK
aCR1AkX1ErMhyhWvmoldSNcNpqS80BR5a9YeW2Nc+Tm6ilk/jptRPr1idNcbLOSNXT9lYbeSv4O7
6959kX8Z0qaCHwr7qGp1OAckP67cvuNLBpbz4hDxTe98P4LCMUw8x22xFlwiOXyMQHyLD8znzM97
pINpsEyZPeb0dXJuiP7HgaMW1szdldwATtrZwBJeWiIf/GzsOP6pb0y6/g5qcUxhfE1h890f3Cmh
KkE/H1j/EQl6tBqS/QrkHW+1toG4bBeeieGOWL81qe5ojGWW+jmKb36/zaORKQs82P/Qpl5vbJlo
sOlNprQ118fAE7cfdh++BysHFcNd/9l3Jdunza1absbtDVvyVnAk9IjzPaBgUlPG9MpWjUTHpGtD
Q2k51A5zwUlehVHle6lVKQ30hOfz0+aU1XhiIWFtGD/aZAdf6kqBP8Q+4vIjSTa4kUuL/KH3HxN1
qJczi6b907Rat7NKyThSCuLYkOiuqhk95O1smjmy9H36VLZ+/RANkWQBobbGoo2ejDxeM6wzhOkr
x7Ap1KRiSF3dQgajsBANXoZAnAd3xym26NAUmPqNZflx9kswlMWLO9I2iMQkUk/lc/yC4K/Gq3cc
82AmM0xShge/QjAta6hR2JLkd46FSydy9xEXYXz5xaYD+downhf2dG5Ho70YFol4fJqLOOKq07kS
eAonBvekOeNb9rn7koMo+obuKeP+nZQsnskPSjGarM8VYhUG+LlQJzmebzuxRfVqzLWJhGLxHeGy
8otauOEVG9Epcc1oIp4QPdbdpneRMep1Ha8BFF1AnCoCEdHTj5znLDglBOP0K4o73FuSP8m24sJy
SoCM7Izk5TyVu3WSCFhjsym7jfLbOIJGxji5onSoAPgaK30C+SdaeFypp3fjNVYqu4+WlCtw22Wz
mDLdf0P/VSZXEq6kOV9h4SkAMoesZUxMTlmJOM+981Gxkku788eqe/+At2n7+L63zLgAAYyJulOt
FB83B6VCwopRaexd1xRA2Q85wCx61QM8A3tMcLdPqLUV2st0DQOrIIFAxStAs+03TLAqK+eOhLx0
UyKg4MbjmTd4pv1ncFGv4r2UYeBT0F0gIg5XUf45160yhC/gqjXWk5AqRzcz7/3ilqzuQmx0Rbm8
FdEyvwG1jLKf6W4j2CoeHteJhueH5LlG3wkihZ7vwhA++UsOtWFBC5KeKT2XP8hOMhM2VXhJWvaC
PQS3jtI8yUsLs5KXWObKSG1jFEPoraaD8nJif0DMM0DpLMCaRxJFW1UOAPRVRgu/J6WY5vKkfs1y
Cjejz495px9Mr8thM0YnKeMBh7U1Gz91KbkdSEzztqEOTUhfH14CcQjqvPgbHCNi8OFDHDCs7MTR
qelXRGOG1NeJx0jwqSPQvK0NkfNxHk0KxDMFaeY/3S+UAlkX202pCnn7jdN8fLQCzX12VgrDU9Kz
nThjs9Mi/+W1QV99G/xDYPi/n72uM+sJL8xfWRiI1mKSg4x1+IM0t8N3nqBG4qWueqazvRmJJwJh
qLDfTgfts3Arc6KGS2zb/I2NaTmQsjJ7J3YhpHepP1vlNd5bMViuyDlToV2V7R92/1UUbLgBt++r
XhHqKTS6iawKF7XGeU9gsuXh0J08P1GzXDEZjrRkA2Pg1DWgOFt1mxoUXahSa+tJB2By32MuWz2i
xz15VZaZUPDv2e+PNnz2dlMLsiDVgBbWOszgvDHTcciCJPTR1DB8PLKmCy0Uz0nBTu5NooT10kUF
o+UVnJdBUQ4gXfLYg6vLzJsDZ7LbUWs5TNIBy6AUrnyCEybKIWFJOkJ/iK/5sbOpNfa6wSDP8QS4
D97Bo6mJqyM1NbIO/+xsirGbhIL1O5ilVlBvexxktsfFWa18UAOGSck8M0Y/XV03YOhv/lU4bFP9
aVSbbCvPxZaTBPbcxKfZAd+OFDSyOou2D0NrihrADr5dkWhWPjYkh7fLQma1C5A2dWDvSDc8i8WX
4kHzsHnluWqQbniAmwNDeylY2SbabS96c26FMFBbCLOdr/onhOCuPGZSeecKzGoE6r4DJcnYaUvO
Pq9tk7w5i4r35kvSMqaNiyUNDEtutpudhEBEWzZJilSZ123BPNTL7g5+bZ+F4o6sELHnOLtp48ps
xHT9JVQmzOm33YXRYwJ/j+DLyU8Lbj1A5urPiiD9SXVhKopS2do7T2TwuGCEYyNbe5kHswsRyqVR
dqxb7Fwmqbw7dENfbPkPPYy0EiPhVp4yCWPi12NyMDd1j2dD8qOD1YZEFf9n5u61n9ihiLCAD00q
b0UauCUUJ9ws/fyXURfFA04ABH1FVxMtsZoatJveD727HNJPAqa8Rmni8eDaWnKjZ5bR8WKhGhB/
wT2tzdqBX31EkUHNZ8yOrMkhrF53Lmdokyhkt3Hjil1RFMy2AwH6D7VVwMYPLhGdL3yn6ea3bBuB
v6l1y1cYA+TTiOuvwgYmf3ff4IV//n1rjnDb+BWcfRw4Cfg2O2buapvTkwRQ4xvdp01uGkWqYMK+
wXvHYPCd19NGwESz+omom3KLuV4imEnrQWKpf09oyjUJf9DYGPygaOvG0uq2nRkJ+n1jR5/R4kzy
bUeGr757JP/Ze2Ht5a3Nt+ICAZ7ZTOhIqCJTmZqAWIn3nAqEHp/s+m9eQSe5Bal00VM8iH4SPXz3
XM7LvptKjoX+2azgeWPbbAolDIWbQVF9TFApXViperKXx2Jo1ql5Ed96cVTWbnIc5cjE9r33I7lK
oeFsGJdpvb3wPg9YkGjA1ghSns7QLCI18Lzk2noPexdicNa8rYpvP4d1aeFRM9ECOzLpIF0d5z/F
eEam0M5CyTM4YCt/dIdj2Jv13aP6Coyr2aH+8ynf26JkKMIuUmzfE0P+GjGiXusuvqJRg1I51V0x
AQG+p/7uwRXQugnFwJbdHiXTh5Hg24dlLscp2Khvig1YMTfCvIBPnidqeMpXw+ZN2cMY+N02aMTz
XDWwGcZkoIy/aS8HY2qdUhVMnKGm4e7fY5vhx15BASUYgyEgnmIqUEw+V5tDTuuHCT4+yrPZFwKl
Ekc0DxzJ4tI3+WK9uOXNOJKRmRApHJ27Ft2REXSTWQ45rcZj2RH+Cpatzznr58rMM19xKXODzn+i
Q3OuvislBzzx5SPwPkT8MslVwrESqyAURHiRzffsfQV7CJiUWAEozjL9Wbsl6VzP0rQhB65ZRxD+
ETbICekRxK+Xc71JIZKXmFMvbr/Jv1qArvaWETqEBngyM3WxEUtgLwPr7dTz8tj8yJNMD/uVndx5
JconUmW2+GhDZWS7tGU9aoTIJ04VtVaKt/YPaAYBCXqEupAJLgF94QD1dpO+Zl+o34Ip65/Cxxvr
8TR7z7aH68IRwEtY8YYKvWI41mxEggKKdGn6J8v2McBf9KAZnz+9QPlbS1Y+GzaAATX0llWB+lUv
gNT1ql6WVtuTUKHxJ+NTB0YUFsPdNbUsZqrugZT1CZSoscON4tRXY+pQe5u3fiLXNSRPAmhXNM5p
yQ+lAdgxMJzW8SEceXwzNDsPhizQ6ZJnbLcDGblh9azKQErgAtGWjrpfslQG5ItrN8mzEX3rb0eq
4OhEyHquwNnuhRlmA82uozltaSMaLV4AraANfq42g2TBBJolwPYE6NnJsJskASn7rXcZGkIk3pzH
q3lldG0Djhm6jFCI3FMorQ5YEz3Di8R2V8LD4+fhU4d3bb4IYm/jJBdObGOOuF477EVihClqckG/
du+Gl3TSggfJwXGRgPRmXevzs+HYu4KsbD013Te9fBWA95uTwUlwIsu/cZMpD/cBZqG8rkKoW8Of
UBoezzorzzx9kUnJK2pYdiyfNDM+IRpOVbk14vcNAIp8M+KSVX/ObMvaNGeXFFBGDGOtzjJLsj+6
fr3DNW1DBSNC0/uPHPHPLcUpHatgkhvkKY314+mY5TUPq6jpIfCZmfgro2Hh3PoAUgYuze0OJxTJ
RumP4guDiWJDVExsd0L+JS8dPDw+p2s5nNVc2IV6d6SoDyzizUIQyhVbIFQlhyHnzf+BwoGb2aU4
zCI7VkSRZcqdOyTh7tdBGka/VWBIjZQFuJbj0d1w+OvTa0VJb/n6Bzil0c2MpYFf39XhHlLxOYTS
eSdoDWPjRZWs2LnrGPAQfy4guJrdYHHIL3hUZ3uIs7+1Jx2Oqkza9J6o8JhnivYV3/neuLStBRTK
w+2Gyi1BXx7pF+tMmDDo2FA/+pMOn6ljTn0Pe8QUddSX9AdsYSJgEftZMOyC+uFn8Ac+ed9Ee/pz
oZgTpZfY8Hq1X+8H3CZd2tOvFxLGUUwB40qx1e2NLVIzla5BCC42L9/djJYHbBM0GFwZe3FcvMMo
jT6p0fOTEX+T9HLo9FlkXvmWPiJjzK89n2VkwlMwh1qqaEbI1ol35c8W32S+SOJLbFYpqBlvLKTW
zbr/eSvLtRt+ZG9pjaXairesdBzfB5xFEPHPo52jR11EYCUjaZp5SJmOmA1uIrPdN0wGlaKvL19c
WNth3Hr23V0rM4vkubA8DuXf2mcQGtKG/P6+eM3eMR4hl/JJPe+bQjngJ85BPmxXzIViMo4YFTeW
IzlnvZ6PcuO5ck4KGTmGzTOHyU93hRoyDWAwdwTglAjzI2HcO/jyufWB0msa9ICqTQwDDQ9/R4Gq
nsMNMpsjRt5U+j+Hthi6GEhtzCFtK/SlyIa2JYR9n/J/rSYic2xKjwDFq/PpKNeYRuE4SSbDia9+
2osG+oAhvKS/0zIBFnMmn15V2yLJ+5qEz9fWMiHZJy56QBl548UCSxHIJdVoofQie7NJ8bn4g9JD
IgHQPGvpXhhtJzRA7AAkS1FVp+goRCBi6RZlCBFOv2371dVuoZ7DOIRzz59fOKL4PHQTVhpCQTGQ
9iyKZTPXbMFoeKqXES+fcndLV1irz36ajZ93ozsdUtGVHWaxMHSa8E+yivBiZEHja5f1Ypi2ao+i
dXMdTuWbHq9L0W+dphgRS3bFNUnv5esGRxTSXXsveyF2e0YHKFnVF1rnUBjSbq6JlOLUEyPuzbXN
6efWP2YF9Tclv+dQpNjmInVwvJl3/5Cc0Rv4kwd2wtwQj12j8OP6K6mRn1sJzAme+Cr4lyqpMwnY
qZbf+Puu3Q3Pr74sBARx+XCevSlT8FR/3wNF/qQ24fYiUq21eEkMCvCbwa3TZANlm4AYk9+XyvY+
O4ZoaxBd2fQRyS3CXb6WTgwLy5+BKCQwThs/RKKWMSrV4a5y7RqpGtSCzeXfS4FjZar+7ZOVE3LB
rgu5hHPKbymit9SkjAAdTfkFoMsBxHZRtXkjphimI5hS975ZQ0ns/GT3wCv5NEolP2p/g16n+PN/
p0NRutGz2mdFqALYSC17X2TZIoxRsgEAi3/PhufKXwZzk/II5eBJNS8Tqa4jZjJtll+9fscmCBaJ
rVY3aglxAJUcshqwaLTboPPqrxiQ2kP7Mwt6Xyvd1YLz/9PeEPeQ4jnrC4qXTT1U4HEuJE/hTt3f
SmC2N4fxSpHbAU3hYa+W94K2Iwv9CEDwBtpCtCXjalX4h3DifW3AvOx6XZ9MK4KQy3rAvmK+x7v4
SoG3VROgE3dwrcR6Nc4b/LnG3LINlrZn5CrlmZOh/R+t+1x0OU70yxCsAQznwjzNOVmBRO6O55+x
ke9WxY6udgTdwL5dZ/p2ntgVdyNIDpiRYSC1WW9TQKTB/ODkmiqHb00Y337X6e/PBk6+HpujEl+q
CM/MyUXsg9kqbst3e3Hd3aYHEFJGRtCHryXc8Xae07RFVgf7a1b7+hNdHgVWeoCgZnMGJrz14ZWo
7qSz22WvKEA7sClsNCDVyrEKMbaIlHzlFYkcxapnFcpNMOZOSoQv/06oVtwAyuC1g93i7mslb4RA
FIJRVpntfffvfxHjSgJYqXHw6QXQEL7tj8pbR9zCF/8MBTbUANMjO2XiW2sSQpGeVFsBckZIXSup
SdoZ0gnUdEG/JYsf+mDcW8NQRmIC0q8z5KDmfMgkNPCwfioAFiWtRILq/AhlqbvurVPvN6mNZDKk
mQ8yd90lNOlZbHim1Ls48zILi+ybrRmv6BA4wVGWjezbYmG1+lEHjW4zSZeZJc2xza/XOPtVqsza
FcPUlmTAiNgBY5Rq4JVtDEkIXNkQI6h3lrJUzShW/EA9VFcYYBQQo3clSs/2SLskyJ140ZHs90MW
ZXG2H9JuNa/64JhnB1GsyQ/wJGcmttT+Ux29Xd55DO3wST9WficxhGybS/p8BEbruVmOQTOYLjZN
rS+s88fSA0iY4liqCWclunxQuUL32at7MayNpDa+09t8sS36qIWr95rewnDPalgSEhwV9IN+GkVu
BrRn48fCIRsoMO/s4BNOV1gmLLy9N7BOKB3oPBcKAr9PptFEeAvsGFAWOKTy4I1IM2lqObjjSzbR
hNlEVxI2aMCbt1kT6w4GXRCkCZM/QwCok+mt3hE70CPSCzEx1LnfPcBnzAp3pEp1xA6J0MvCIZ4w
9Go6F+zi8jUUK71zgXieMOq0DgJelZryNTQ+2yqQFWzhs+uJMgA50pt6fE7HyDNKT7zfSWJSwmGW
JD2mO0Kq06H6MyoZWQ+30zr0L4EX3ZMAH/ovbB5oC+HHOB1bu5WstjfXuLpVgZYaCw1H3Y0EHnPY
+ZTvf2rkYcRT/X0CVg3XInHI0cYEbO13iB06fVQWl3YFqXLeSyYbfKnAo085/M+cOE4m6UanZ79V
2xwKPv2ESoXNKrCO5GhqjUJO/qFmOwT10uDqvUzL04VR5OP6DTpTTsPtRzyfqfUkksOydwcJhZRg
npZmbzjXe7tC7/yJko44tdFy/VUvNxGLUCQd7rWkYlEMw4I+xjhVI3BXOoDV/Axn8l/7FE85h0NA
xrEslzZM8TBsRdsfBn+xAyj9eFGxt7DJm1w3XNonNZfCsOfABiFS9O2dmeairYBf0Dg/Uz396bca
EGXV376mEVSeUvmNnVDL4U9YjUaYunNR8jz/INQN6fHPnHOZ17eiYR7QktPOQM+tGlyjVWRfnulh
o0GZbnQPqF/4SFfBya3l4AO3pOAMuzf4pCUAcYhrM4WJwOxF1EcauAW9u0qRrzmodjyY5mnqLn+z
UptoZMTSiyXYO9I43ts4KBlxMvuLIpY6c8T/OYweY1DJ/UtPMVqwV7Rj6seWKDLN4g8B5/XUm6tk
HYXwsKZoWoYjW66jfJmeQ94tvkQ4i/L3N/BGOhnXMXZ8WWPPGKZlmsdWP4ARJytVBBnHEVkOpaHX
/UrVE972CJa6mBLwhaM9PDFxjcpC+fUlNIeVbMxbMzpkNdpfRxPa66/mqgsOqOMDSFQFfpwOsJmc
OoNBRCL4Mo+r4tO9Z8I23G7l7OQKoBkjpcjVQYISCFNAi0bZss7syhC9YEsEFIfkKJT5g/DAajHQ
qk+KDS+nZ1+5HE9lxN5smFvdhdfjU1Rv310gmbD5YTTH4izS3ZcieSvZlH4BTHwXSvg1x5o/dhjW
OWe1DSPgS52x0I672J37Yp105xx1hdqPfJAGM6V/6/OpUNmFlvU/ZO3xWRjuMijcVXOV2IxjZ4Zi
JYemoKDarefBylZKRulxsvGHZUMrWy9k1+8zykDY9xZIXaFCq18Uw8O56azYIm4ch5qScw8DE1Zv
Qv3Y2/0z5N7Uy+LZLnDT0qtXOg1H3WMLXmIvdLj/nUt9knOrPTlBzRjrB5CRA/aL6yQrQ8GWS+2/
vhBcmrbRQ+dichrBG3X2x74myw4gk7m3O7s0cQH5OeZQFFNxeMw1DKLdk503d7bspmsRfIjPC8GN
7ilv5SSB2frhXL/BLjMKVZOY6K5h/MjtyUykNtgBcX4bqjcf/unTX68SkL98wJpG3gPZrKJchXwp
Qug0UIk952ozK//daqBhGg9rIxLVQ+Zw4sRQ62L/YKBraabzj4BInA1WFBKSX6v4/ztsutz6EyaS
C3em3hCgrvhVYTyWRbpvAMMpgeIrOrDVUt4DIsB32lCwEV8TtVpl5s+C7zzO9c+R9PqUm+oYMrnd
Ti96xasF+mJb1GerTh48W4rxhxbQJCFiQKUgQzD8FYx+vuoCDiplGlrRjld0+Gm0wKF2ymu3elZQ
eiCrDRl9GjO9XA9wGaUjdvt4ZThygkuJJ/JcrrtRCRfN9djX1m2xTq/2r9fqONB67B0BugBHobfc
905yQA27uaH/KlIyrCDdd6WYqSTyZsVhMCB6Waifaz/aEFGe4AbWsAYnM2Gjrf1KFlwFiNbHQCX6
MMEgKqERpTcT9aP13K7PG2hoXZe6n6UhxLkxZM36XuAPREGbvCKH1EF0TmJkGWF8EtTtoJmm9sDr
SwEu9WkI+u01Z3Y58Yllp5ANsnBRXizy2rAKTnKc2v1k6Ad83U/S72lSAluudREgjaveyPYd3gwK
yHCOcAAWjLNKyT/hcnqaUMAVzA78mFE6SjxLUQ6IE7j9tPcWc8Ry1nhXQ8ULc78A4sRq43SZJ+h4
gp55jJVSTWtY3Fm2NhCQkwUlKRLJhnBZB8XyPK7iXj2N2vdhRsFnhqnUl5EIfWqtNhkfjOc+c1Rd
C767J1awy4W5Yt+CDRxwiIvRl6mft4z1pqv8ZUrB+wm4TMfPy9R35mYXezeQNgsZaOyXhXzbxBLm
zScrgQ0zoD/CV4XPXEr/VPaFxMj0de2hJc2r/NmQh/NTaO5A79P27Wl+fwOv7Vx++kSQZ2NO/okW
b1wdp6AdA6fM87O//aphf6GdbL8+ltRBIf9r+D6M3frTPSjvPayho66U/o0FlZSPsX1Fr0WbGOvy
3GiFFb3h6XZZhKMZV50cTNVt0G91Y3IV3/9p8fQC05jQCrcXUu+eBwIoAN81qeuuh2XNI+YpsccJ
XOEpWRtJwh43at+Sx2CAsdorBL9KbDLm/HaSmSSSzzGdCDBT0E5hnUE55pd9Catrg7SO81dwXaF7
wQFhUfLprkEjBhUkJAMOX7tGZqB46uUMEhHIM/hUAVWZ+O/KA2MuGSNgWQ4pzV52notwFDSemVO3
5C2ZaPNfoweuCHvvsp4DaEZ5D1F4hehx02j2qRfjw0tVotf7/Cxj+sgi0Dsb8Tm06G9lBb7KMmkY
JZejXGddgXbPMM+/Zsl6QoLcT786qH+Jw2KqznN0cLEuCHboig8COdDatVJerAaGLlAnSVVCQj3t
rTKS7qUQZaY7j7Gt4jZP6uJe5hIcrm9CIiP+qsVea59FqtJ0socMnZXVa1CjdpzREtRkdFmB3gdc
lNxczr7FLy02bN2N6A6hvfqsBxerKtmNcHruzVdTTDW9nYhd9GNeSJccTPzOvtfShne+YJYxS6TT
HA1s3249AcEiryKmL7NGn7NhRElag+kB0JWrWwFM6MLlKyfGyHjLz7dN1PhPZUX1JxuVL+n/alN3
MwCyU/R/Cdo0OI3oIuCs4kAAyXA6vytkgCbRn8Wq9MkqyLbznhCOvUO8/URZvWZjcHxbKadcQw4m
Wgq0TG41mX99MlwdnyEF7WJJpwby1LqeqnSxUns2rceXFJLiiaIe4JjXn7gSi4VgFJU+9V94BEwF
FSX3ShfNYMGbcp6zaqU53pjWBMmBLIVuKNpX6QQU1MbBfxhACcjZ4qJ+KYvc9VcPgQIq2jK2ooJ1
3NHGw40uO+myvFZQa6kEoDAHGM8VwW+MWFre5/+Exh4w/mITAgqOTpLh1Dvq9+tAuoLLzVbEoAA1
nkD0hqoshvft8QTCkULYsv9Q+Gkj6e8U+lmOJxy3K3eYqHJ7mkWMetH4jtfG2TwdM8WT3tglPnya
CJD1j+037vjKFqdBw3KGPp0+clvYvF8FOyln7VEkzzRb0pxxdlSiaFvsGMRDlmFMmsBF09yr35qk
AfBoosV5jxTaFsOEcuLEHFOQIPBZWcwu3qmP/VBFICbz4CZqja0yi1Dfr0B3A7CP1uiRdXOXmULS
Q59hPeGagFx2wc3F3wsbrr/HJ52ls2hIRx8Ouaef/2E2PY97pp8hSYLtxTBXHPxlL+DS7L3/pKLO
SNCsw+CzOIAFo5TToS8sprrt2JIYsI3pcKs28tEvmjBcdrTJvcq6US1TrQJp0mgpYEMx7M5k3JpQ
BoKvKHawFuTgKjrHBtOzaUs9FsXdwU7dK9A/im6f2KZo47bqWvbIlONCHfffWP2Iy8GDby+aaEk6
p2+TYkcC2E04S/TX6YC9/iZ12RTaCHM8HGTW68A10aGTCyHpKkDPsJ9eHQz8NiHMTDnpEt2uGdu3
SwpRw6rrBqW206JXyUafjJBYrAnpuiJc2FKZi6Ww37f5eJsKiiL91+++CAM8YQYfYSlaYapqMgc7
ylU7M2H1654Bth9p6xruWLWGBkG4TfoGisOE9yMcBrWAdM0V1r2k6o1SHIKhX3GiSY9kZlPp8gXQ
OjlFNC6q0/zeeEM/P8JRWTsXYLTiu/13lonmsPs9sj++j3IeDtkowh1i05JoNzVw5CSKus56Jb77
GFjjWmT0ArSixcf0i76KKqtQ8ieqevcYYfMRqKibOZ2hbeIwGSMHt7hGWXac7pbHrtIRuGRSu0fv
6SrQC+VomRm0V2t9aSws2FavPHza6Jvt0xrMLm83RfKQHAfxqzCTP0gM8GocbuWI7tDPHjlYFQXB
ltYOLKRofa1AtvWyJkGjrfsUn+9n9VdlvRYAslLMYMnub2nqBeYXbBpB/oCOnWkQb6Fkpzl9cznI
8zEzWBrfsz2Mfru2DyPNiFXDocn4y4Dai0L3ZQR4KS1IbLKE2xVC2YKsV8n9zH8HhwOdBxF3tbZ5
I4f4fhH2yEVGln14rDJntC+GqZ3kqfRPEeQjQf+ye7uJDErx+cRZ/EGqfidDlqm2rk0Q7dUDnzMz
DiK7Oh44CTRmeBy4M07Djcfxh7Cc74yPOnEtOa0ZPoa8H16j/NpOmQjnopW3gLz2EGWaOxUswtmY
qIl41rCUmLN3Ar3JoTZZ5gwPjimcFbUJ1hwS9t05TsMsDyrtv3YyK4O/y6qgxJz/OlvwZbenMnrO
kT7l7fb2uuXVaXc55PtvO6aowQoMaLOiZ/DXbMpQjSknmpNOuRZRGw76j3S/zdkm0UiVNzc3Kv9d
edX6RqMxgqgTYzsqyzNUeHBxAyHuOOPNEFh063fviVfPukkap3bXzq46V5qOTSlSu6gyt8DfRO+6
CiAXxuwbdz2l6fk1JwUVdZAuR4SnazRS9V/CLTEaTm9FeHr7pdDG4oKOcBecMrLHfQkcQPkvCFgs
mlbJ/y2UDFqYneq3A/eTKWuFmb3uk90kxiN1bazBZqMiCOf0XvOITCwqCcWkJLmhYZmDj3Edj97i
t2nR78LKLX/lR7SReYAX/Toy/HnvOizFL1FrBXojlAa7000hOG9ZSqGTUOOl7o0clXobyOVtVv2X
bv8Kl5lADg6GF8rtHwa9WUwPjPQ4DbVEthAL/F1POSH0Wbg1LtE8HH/XD2nVgdmjbl8sgTnBqAGN
ZrvAHqOwO+AeERubMefB7VxkFvJdm7n4aEMDGWiCeakL/juuR1Z+KR36acXADJOXlS28s3KVNwOn
ohAsprh83nqeSNciOCQngpMGCBEuIE1ffdquT4j8zoekUjYD1ihFV1sjlqSB+LHdxUsjbQPY0iOK
QD3UM3vX97P2SAP0h0mKFAqVS/iWUqxjmAaDTTseeNPXKVa3sgVrxekrpazXytI9xVaCkzeeBsJ9
5NQ+uGTZX/cN4quuy5oFcp8XGM8qKUHxYntIvHYh8YOtQpsMgfITwd5zUSOyYfy9kk8Mi+q6vgER
Kdzj8IU/yhrqyx8BJAqMRzy1kcQeMeifBFuClq29qpp6SeOYghdfFW3k75YeiFznNMT8Hw3moXgr
7MOTcCTipPX7H6qdH16R5AGlZfkT0yB27agehetHI5Y5Wj2aOaPzOKUBp7v4hWq1f6MD8CMzX95b
AByC6c0Y6iq/GIBYpDNXojRh9ZZMSP8DTmmkMZke+8TLZW6ImRQrK7bzQW6iD5YUFfWijBDNAo79
I6e3gs3bu4jezIULhjWHFHbmMXVbUA5OIQN2B+AqTn/cIN4gISATeqXmBToQELCSu5KfKNSljEcA
zdZvgRMiSwnRdkwIIlTIE8+0WMWkaJlNfbbCmimspA6lyUvDD0FhAachJTmtGn6GcPCzgoR2Jw1K
/J7077IqbD+CLhtNoVdhgmoSg+zwxxhwlnwSDtGOt0ukyqirg5nY+YCda1pYaGitmLHgNEqcnp7e
g8Gf4wUrzuBDuXAt3tcQDnEwqtUH3Kt/ZTWmPpNvWRxgfejC6lwA1LOCJlJV2FV4swLjTgYvarir
DUd9Sg8qygCyRnl7aEMa0kIoUEXAG5sgkblOsGbY44RjnbIfI0amp1+HlbOKAK9JbQilDawvspEC
sdS5PAjeKHj9EgowwyJsEQBgruJMFKTU4baeu/T0zcQTpqJM6UUfexAOjL2EjdjU3ENVSAzl6vud
DNKuLuQfy5sxWPqgTk01ETdleDflSYcHhNB163La6KQtywm9Yv/RJ585lYZUQ8Hzeyf+33cp8SE+
8p0y/TkVGdnYFWUwQx9Bivrt+PXOtLbkWKmVWo3wF49P2gzzkTKrHu7yAofcLipamDZjAWFg7Gct
lnnJolpjcMNxwCF/ZFaWHPYl6KVtpzFIz9sMH0f2xakZNz+N6T3LhOFRxu5tXIvuAqY0Tdvm0TCa
AifzGnweuTL6vUDeyDkhyuyHaecUoyoQd4/lph5qE9nsx5Uv92iO21wDqVc5iDi/PCiR+IWbgWyO
m9VoIOuJg78HDyqYUqrzb34qtKKgKU10bS0DQtxCwJjU0HgTPJ9QBuEp+cTJrPMBobFdYlYhjb+N
6kItaVtMNAlRx9zsOIiVOlZ1cywl7bz2oNy6r4NL0uvauI+ChE+/8HZOi+a5I6o/N15symgWKlcx
o1MbZp2jGhG3U3g91exVqIfayeYneqjLJIiDc8QUs3pfL5+eU9PYt9H8zHRcOFDroiETGHFJlKfH
+CuwhMVGzsiwdLFIv7rVQawdb//Wmg2qxNi2DtZPrVSeL5hOxdDSFxCWrejT4CZiaDFcL/tB7opU
Lu3h4ijA2EwIAcVCMxWqLjcV7fSny0NTQ3u0/vrv9an9gE/scbfMvxgoSAYqkq2jJcXjyTK/4CjI
O+tO1K/i3dFSC5b8vHhQwuouTiIvX5pw1pnps3jOECDagn7OH5Dq3q+SFUrUtD9/Ty4N3g9Z+16A
PMypKTlu+9MygNXsRHgmj9dtaSgyoBgO1+TzSwR2MO5lsSQwekPOCa2+VRPMhSWZTfK+EWKIF+2i
3lhD7poQB4+QwAmvqwOlpoZIgxFXH5//I/bO+N+vlg2/zcwTwj9DSkHRSRLG8HiAAQuMqZWm7hvm
UVbewA1b07gED5c7EX8TFh7F93/oHJEv70f9J6h9DmklwtY1FX/cud2Qm0fzsq2yukSYkBoC1Tf6
T60OUAG6uwEpTdTwqycJlvkeoWsVEcZRlLtyTjMJTLgxD1sxKd/Bg3YeZ3c9yzAIM1vER4IAZFtL
nlCr+YTC9LvGhWy7IMxVYVFv3GDt2MHY70GaFB26U9k/OQfPsCYJVZdj0UEm38TdSEFnkX/Xgkpw
SFssqujSEqhGJ5nPIySvYLcuSyAsIvo7JtE4sdcabxuagBSr8ZerG0RSIVioROmVUHXqp1tNIJ5x
KtNAYGgckGyNeo+ctQV5lkfN2zwXS1VUJzP5OYxHIimSgfVSPf1N4+7f7O/Pdgn9hltxsPcHHSU2
gRbQWKtcjzKuU1IZPMbbwhXwZoJ2MG2HkFrJdzcYPvtDmic5nVGtDvhpgUF6jK1C4U6Vmc/nN1pL
2g5Lb2lYRr9wytjWYLrfwpNrL6mLw7g/Hnye1Xsw9UfAIq7piV6AtSDWj5QN7MDtZQk5eEOAWxfo
mUbsK4/rQYedIXBUD1B+MfMnomW9U8isE+tEhGYF/dttFYImXEM5jFZypoNX1Aqp3lGFLYiWMxcJ
zz4vW6dMJ81AGgD9kLpxXMD1LeSExlV14w9HuyRi+RmjNlJlGeHpf8UnWYVrRQ5wlE6zNTVXqPYi
HzGbPMmLc/FgoryStBHLxNrZVJ/pqzLAK0sJt1DJwUHEdz4dkfSwKMyRE3qpliRKw9RohMFjL0XT
HV3CGDvlnSoGQBijIXsy+NpalJJTdGQ3Aer+/jA6T0M8y1KFNL7xCPCymO/npS1zQbOldHwD5Dpw
Yp/PqRDzSZxDgdX3AUsZcN/F2x2GOyUvgI6d3KeZkcKmeGX5bhUsq3FPNObZQdJ6gKz9SM6bxfXe
LfGqS79gmwuC+ZxPsG6Tyf3bIbyHX0wCagrVex5cCp/8+AH4ENHF3jVSHfYW9rn4b01UewM0qSWu
/bqIQP7LWcr5/Q4CzmL6vp37mjh9lO625W7AXiOAvZq340a2xohw/OsV0GLl1cY4A6A9v1Z0Kt9c
Aeo9xMrokOFiCq/6cWd4pRulvlNDUA8Q42CziPKp6e62Gem1RDE6Zep6PaVkeHllKk8ghysSDEtK
yfsKBLKhfsju2esNidtZI/uShGjs32n8vo1Q2+v1vtpRszHz468QVuxolmX/XjbHwiPAT3INLszN
xmGt7cdUhZ/GdGfM4RxMF2R32PrHfoHJ7S6Us1EJEg8Orr+vUi8lVB1jGI0u/edxQTBAsPUrcBv8
/RTgoXx0FIfVj6gjVN/ESlDwkIAjgLzM92KtxIVbVVhr6/NPWcuNFdYvbxrumc/3Cd11a5RgpsRP
Q4rPI/2rI13Dp2H8DakGbrswZoeF9PhxN7uFvMOycEzpGxHHmK0NBgVgUQMjB5w3FRBXy7l0MUUr
t91M3nIM11zERwNAozBQsu3nTV+nMsTEffjW14M2EX00dsJzNQQqaxUW33xISps2WFBEP3jfrQQm
M0thR416hMghQNgSJbCLFcIatvOfOLbIQUFNaRPrCVSuo21iTOYIeD5MS6CFTOA+WYB0FOCDtX6L
YipDfZFMnw+4NkdcTklFDnlx5KVQdb3yNrcv/a4EyLloQB6uDeVLzfmjS9FriL3VYCt215CCPf1P
IwJyOpk+RzXONil+wABZCHe6twrrswCQQfb5Xjj4qKsDiueQEZJZGXS7ZJhpuY/orZ3W/92nceW4
w8vD+HSAqaFe7Pt/+ePE5wr1sEVhloaO712lSJEpwhJRNAZ4r92e+JpHWd8R2ertWg0/GYbJYsUS
eQrxKrjA9xpIGl1MUKjs1KksZWT35s5uM+Xea+kklL2lLqQyyAWfYqp9CiiESjQ+B80adQ5n+Wad
7gg0iOoX2VM460bgrVoH2k3eoC5aXmXAU8xiN2b/zMvJL6meh3eVRnmHe3FciHpqyWuLBWrNWZNt
04hqHnDkXfgFRRvgukeWSfMkMAiziXgEDRB1LEaDCl771CDYUKHwgoSL3J+evnmWED867J7AOfdS
f93IFPXYCPjNqf9aHaAmWU3xgOSQfr4xucU6LE2OVL5WLRWsZUM0HDgtXaG0wXObP/9LrtQtWTly
bdtKXj9XXPCWCxnvg4Jy8Zr+RCfgjhKbAzQ7lOf06UX+RwwwxJxpLKH+zdx4oqXe6dHV6XinHvSC
tNZg7qrd+L3CTfT0uCnQVed1VVPDFR0pmlaM2Z48+ur/DKOor1eWnbPJ9+y/wZVYY/pIzi7sh0En
ZHGZPuhRh1lkCxU7zPI3/jGRmp1VVLTRZgd3tAkAwpiZzFdORBse+W8OleitA1NUP4pmQaGHaTuZ
qgnKemGVygoPLeslCkWnaaQPhJZNqahuyEfvzWbGTPUX9uXJ1UVnjRi5BNie9/wiD1aodTw7ZXS7
fy09LxkdeM7tD/Ur7E5CvKzzI1FT/Z+FI8Aag0s9uCWu9+uZLmEh0YEwTsKnyJEVJZdq2v5NnKhq
4r/MDHaQUSKyhV+IlDvmmYanj55udz2hqCpdFS7Cd+lnwhAasc2BH/x9nWTcJHEt57+Qz+Yq9HJU
fcK8wciYVRFkEUdFthnv17XdbNAt6mykSvmgBRTlezCXHqomMP1wUemzD1a3taES+HBS0RvedH47
U9vMron08hjTNJCxGfgUTtjAsx2ldg3muEg0Sbxn+AbSjBUoxzpJFWnzVjfUD0L/GMibP45uMzjm
1Wzcwe8OfsNren+hs4b2W/vD72xgq8SUFIWEWPXyeQE7aAC3IdCFJpERpNXbv9d3LpCuAw+TSeB4
WQ3A7g8K8xVbQNtfeZZlCJGWBgHdFAEVrTagBUgQvUiKOE4zTU7vvPFtI1or1lh4o3G+cS7MUlLt
led/LRUW5xhTlv2Nfpzc7d1kw+2U8EyjG4nWUwMucOf0a1OGJg9PZ394LLrgYaZdqGPwLBakCYhl
2CxqIEnrFRGb7rCQWDVW5on2cAK1l6i5rlVcwY39gKT2f72r/wHl5jI9kx2/GT7klujIXubcw2gF
uuKlbC6alGB1EoBZMil9OI8qT3HuhFoVNImwQhsPqyfjn5Xl0VYxwrjBf2UepmbXS+Qw2HMR1ppr
45mNcsG/w75tDgi8mm1INTOJquGTfl1eTg4o2hZVkTIkAlvOXH9Baj15J+TTEiilG7UVkxmTvoI9
fK2WGFZV9NbziMmARUszItr0HJifo8wBsXhOzQju/v1HFiFNyEtPclEdwH7uYuaUI+rrP5V+vJ3G
6N5cuw5lscq4h9/HyB3EynjSEwy5as4rMbx2yKg3Mj+DVL71B+XuYUGGYQyBwVqcu9AdV5tGR/SO
lqckakNcuQqZEFmN+JA7Uce/VlDtw6GvmoeVc4A1WbKP7fgxM3Cz5rDM0ey3blDT0Bc1J80IQbDB
vAQ6vYKzn4FzpLJS0myOuYIDZq1ReiUv2JUGgZtc9rzk33/FqX3Z/F9bNjl8XV6j7wuXHkRToj5b
ARzhRfpy6riNeEUiUhHfn2GJ3PuA0z72s4SWjqY2//OSuAi+qSpKHdf6/iVb9sC5MCNLknu/vBCD
olquyrdSYpov2jN2eqNYYk8+cmzrSg/h2rs3BvAAmAu44PEPBw3Cs3U+iibLHbVX4B4pkQK9pWly
eD71tgIGh51ydRsh8WeAUqEozFX7d5kW01IGFkyrHH4hUQrAciv3qZieyMsVHyIc/IdaCWlDHNVO
/2+CbJE7+sYu+F+Mhez5ha+LU2bpNNQGqziew/8CbFytgymEqLkBTSDUUqH3D5Oi0VYhtkZz32uz
KZQgNEoEleutP2ZF67oqQyOaRZhnxck51co3pcHxTDuBSXrBhWhJO3KRcLc0ydyovuXubegR6fOs
gfWN3gVhOdpUfl5n5zwzTrjkZoeaNTj0QTDP/1pvYF5sYBZII8Ov06AlxFRo9mlBrHjW5LEEe22j
Hva8gwxol4+l/bX3lFBMa/1hxw2wexEnkwHZSoiGS6AVHWa24GULCFFvC6NUEfb6fr9fH344w5UV
w5hILqmxpyZFFg7EMGHrvoSHJ/7p2N3A2NbB7t31O/5d8XjHUYt+Rnvj1PmP3Y2fqbBEVfVUSg9n
KCe3vljPPTSkxg+h7afXcAzHJEWhl2uZ4oojFEGACj0TpeSpfWfqdvoVnvvHPFn7D5MluZlpUM0q
iaBF/xFvFZMLrz6H+bt8gLeDvho56Pcp9XdBporVTYwVPtS8yRTOkAk5SuQWLHIcrBEj/VG0023g
lu80w7z5GnIyakUeMcE2FsSQOR8shx+Ez9EzM09HRBaCHszVGfy0izXpjj2X+H0bpCX3kOO3Q8VW
4pImtVosvrMfvTT6MOYjeKKnsE5Yhd/MkLrL6mEpNbHGc3vOmIY/fOfuW+lpvEXskD3ubnNhh78q
iPStIZw9pa6XmaRm844qN9iACEXCLmK13cGZA1uTN6lBVuGrGMvJ6FzsJP8xBb2tgss1ncyn4DPd
xXvpZkZH2nNfj+HmfAjoGbo7qPK4hfP6S5r+YMBt02npwV7Qr4AHJxoywpp7dXxwsdR2KZJeTKPl
u5TLBlBmD2v4sJwpP0kQXuxzfDi9S3yE8hg8rfs/4/jSvEGBZyUEE+toL+Bab7A32UM/uqrCMwWP
b8MwunxoBtXZbwQqsKmaJ65hmtvvWA5vM/vlpdFTw/6iiaawTd60Pzij3rWaS/R8Q2486RZ1wZuL
vF9chV7n3yC140gvK2SAOIvn9LAGXOosNiB3c0UowINKMus08S75AykmKWz+DRPKFUNVEpLowCrH
iUin0NWMhoOWwdZY4pJu94NklonswFxh0PxZt6Zgku2LAhXT6hu9mnh7djEiNsFNMUcW1APeL3s4
21MTipcMdOKBXZ3tIDqV3i23JVgeV+WpZPmaDDKFdLqynhRQW+ULeIGqjp2ROQvoe3V9RItgUnym
YT2v7viD0s0B6NHDp0AVUNoSTvk4m1JKieS6uB3sQ18Lq7LNVLH05HqEltSXaLHR1EwEoJO7iBso
cMtRrN2L+bRW/746W6aD4mEFSblcDf63BgdYcZuKKJvI8aNMoYz2fxH3Ukkpb9QwQw54EHca99bQ
TKoZm/yVPPCzlYx8ykqvMxXYRCuJLf4HtuJbgApPYvMp4+WJs90CwWk1DlFihAXDzk+qNBnCL/Xt
2HGvn5u5KW5nrXh2kqIFcaUCIP6P6nJ6T5QQdQp850Yw30XQEUt5zBVTFeFWSgGXJv/gs2OnxPiX
IZihE8cXtxkoQSbZkraDtMbS51x7ljEMH/LLMvGw1YG5Ms4JNtQ/WlSrk4RNjET8k3u7c5g1fqcT
kyh8lhvUn7zytiLZKLPWBcT7mVW4tcW9GjMNWaR/gpTHtbUsukDRf4tjUNJyQaFi56maMf9LlSGm
MnrRvvAaTumzf890/oxmMj/ctqLr2/NpzqVPhjETco3uUz945c9cIIbB28h5gi4BILE0cFGGM6IB
b9UWojLrOUNjQKnVJ6jhqw2iQEXKR2cbQYvNSjs0PFb/BeEajpz2tMOU3U3eouRErSDCH5lPZFxf
q9S/PArlLjtgF+lMCV99iTyNeDDrLf/W7YwbAXn+aHSCxaoKjiyWj8i2+1BursPx0RLCKF5vt1gP
fP4hSx7KF9skelY4o6xEgXV+emAmFFQlqQW05TeW/stfcGa6l153F55qnGI1oTMxfhjfb0G4K8R+
s9OizbkrWFLyegXh0Ivn6VkYt61D+NJvC4mNMzlMgWB22GgfEv2JWjIR7HDyx0JmlOeHXww39JB3
qkpx3wuguo7tJwdccGKkKWKLeTEdqyxlZa8KrX8ifadv8TITDVohyO+pB/5rTQl089hU4b3tsevs
mEWLAoWb9IzYdy4DKbQKEQghGlXhdRwDdFLlEHtDzQ5YFiPEkVpPsphDxKDF4SLbD6J84DES9jq+
YWtmHwve/zJevfm9VFtwbmT2aa0YhpbJ6Dg0mvkGjZr3BVDIIyBH5YErHSVqGi2JZC8MrRFVg2fl
P6G3OF5xeuT/vQOuCrwAHAgTIDBFc89lsOUPcZZ0gdQ3/KLKyCP7sOtXRGwqngOcfcW7iOot5EGB
wiyl+5/gezrEg2YJIUnxdpREEmhA1p9L8aH/FZKTsZ+/IXQWi/nMBPvCtl/ceT9yAqs+8wv9ERfY
fiytfhLjU2qBTbXWGdfvgMFZAy6qu3En431F0jPM/J0XEI5wbh2NqOR28NDhZ5QKy+qwvEnLcx6F
KG+eDOMD644Dk0QgyfX+ojjvYQ8OuWVstAHPVHEoOQVJYay7RYQfE96lFS+J/O6QNvwQg3B+sVFC
4SVaVkQuDYVb4gfWJQ+BRWzzNxmV3+2+pItWhByWf/awrjQjLufG9S/tEGYR/B8nRFpdrnoVbsGD
fIF6/+Srwz5bN4eNH7G6eu0RnTVlbC6+3NHeAOn3yF50SOY1xwimiBqlsnNyEy1TYg8ugyUdHKm8
LqczTheOgryC7SFDAv9gonPcTS/ZIRYlemtjG5Z2nOKYEgr7ouI4uJHfX5Ky2FPwft4xclkexJdl
6jxR38/cq2MI9642LWb0+Ucdb3yAzFeWwn8PRFj/YzlPycnWH3Vub6wbBybvJYnO7yekbtXmStrD
VAKk/mkol+Thedh9yVYySwIkad+uP4Xhms6s6cPVrTkhbQ57sAE2QkVua1cPpC0VPpcCQlhVtyNl
c+JsviLnxhYBdt2alk0niNTSYsUikXWZivfVSdmrzdrUgZxgyL7AwVMcjYd7S5bKc7vi6YviOYRo
SjC1HikXv+OSATmNWqzxd4PaA2BNFYWrRnBhowvJPDy2knceYLH65o38dtFfLj6F/Bhv2Sen1KSu
vKuk/SI0h6Gn0Ng/azw0fTfeoTIULCo3k9XujFNDJQbg+rVkgblqBuHyie6OKFMlbcyIjd/z0tWF
D4196oO17V4s6NAfH0XfwgE9/FRYmuBwCbBaNHXsWZLSRLMUJP2KhN9/I1BIFKlCaobs+GWuA4Ah
pJzAlqL4x3wch+sA0njLJTxZoz1DsTFEvcVNwi5TCixweHEh2YSzBOveUccphgIESa4Q1lqGh58S
0WXf+dtssKhHHi/NB+zWHZL//c6qBkxSbuWX+TUQlUiyHIzjIhwWRSGwcFtAaX00cvYiw3tRSG3k
DWUZf8LUZ9wMZeFnadKiz0ABTEPHxWIdPShjj/BrYPuW01PmjiweQ5/zXYhkC6Dhoh25vQtsEKQH
7eya5WqP42cDQ7RuTjC4rHZQ8g5n0UEqK+BGJeZ+tTDPZ+LQzNMW2lW7SjIiWmTDO4cPGXRN2zGV
+ExPz+Mcw9wsCDdmmldwYMDygYno6vGCWNvMaHyLRM1VsKg4oBS8gV1RVwchZUbvfdPEETNGm0kx
83J80zJs1/GA48ovWeHot7trsBs+8eLjXNno/V4sLMX7ASj0tVaBlGX1OiyAplf5ra3Yds5rZDvq
4IMFn53oXPcqD7qVSw0wW2sFbpB0mCyHQk9sPs70eRdffWh82GJNFWhxQfcQ4rNyrfASULHoLIJb
wxcidZr7kwN/83VZ8MKWyrnLF3jrnGq7KPELfDz5Opj4qNppIlZzBu+Ui6bQb4qVsmPi0g8N9HTc
g3bigbyJeGoV16PCgV9FZSqhMZrzQBI6VzbhM26xhSsPirwr5/CYTjcIXy+G1DCuzmk/uo8L1qFE
WjaoeI75qKvLSvo/50qHrXCVmiexeHcbvQPa9QLZlD1w2isJf5ppPH7ozw6+gBuXgfxQFpeCHR6M
x6avmaT2JNSasBgm2pfc3iFPGm0nrK9Dt3LYwgQioDPMryvDNWILvVYP+nL+LOaSxy1YQ0nsjkFa
FxS35DEf6fNXYHSVIAeGUqRsG+3xkyobpyTns/9HdzKpC2/TzsA0casihgNhQJYq6WWNmmF71+5t
uBnVk16vRisF+XKRu6Gn01UKeX8lZ/yo6m1RyM0L60jzqY/d5iIaMX4VIPe7/CMDmWrbD0JIy4iK
ttIAbIARFCSNY1q81VzEx+1fOsEaLK0pIhVJ5ZzzXV+QNL5FNXypqqZYqudyd4zOwKG7/og1gF9e
hmLC/mHLJDE0lmvm1o3YNyWxZXEtsNRB/ddD5orw/s4XxM9ITzfOVf3a/bzTbmn9awBIvnqF08kN
EVduduck1Jh0471njwr37Wb7okY035j5ox61uhF8G1Q0w27WRumii21dzRNEVYoW6ckl5LORZ/i8
F/kt/gh5fy8IYDX+EBO+mP0RDlsEWvcdjbCJT93e/NtlSvWBZPF4WiMp/ZlFvldy5SJPrH0BfKyM
0gXw7if1wSTREUcjg/M5PC7GVr1pPTSpcftuvIBzliS2lSgbR1izAZ8nG07GTS+6ITaE2Zsfwl3/
+BHSsMs+4R0d09moqyebRlllwbmMIvru/HlewM5Qh7gdje0X7qq2PJ7b8QavTZZtg9UpJt8B0Ct8
IqiuBC77PWNUcZqLe3TNuEWW6o4ASXOdy3y7vdZCAWP1gLwlXrlM144LM0PdHbaTRd62s9GqSHCE
ulOJMGd//LDCUNdVVpnb9vMVvG8l9HTjmC64KJ8eKqnl2v4VHDE10ohommZAgleee0AUd72ATZmX
R5TKVIRaKt7kPzV2xUaOl6LNWYF85fdBHmA2i75MzZertLzR6Uxvz2KsQpyMsaHzARD3wAOkDEI5
lfqLONUFNKwO/8StZKyRupONprrvrKrIfworlR33fOwIIpYuPY9qmRAgxh7UutM0x7EY5vcTFtmQ
UCwUG+eRKfWA3+ptE1YOxIAVsgAEWSAPeDjxmyF6iH8B7QRl36/9djFahVpNC8iOCWDLf6WTQyVL
DLN8ki/xT/cBqJZyzKyDIQW6RKTmGGT6YrcnJ2h7EnoOqRpHJRoWyyCIUtzSUM4NW0KVzHdsNejj
Ksrdd4HXZ4S4va99hhnm8/fqy0+tiR1TaDHo9NWHM7CIO7qj0njW+xGEvXUjgaU4bYR81Oj8+9PR
C+NxJc0Gmtsft7s1zCKs1hpCNPg2goSzD4dpdMmT+sVUWNLq5tdfd754I5qdyZznMbQc/SeMUWHO
8gYIh1vcUqhE8VjS3cbK/lKeGrye1mykqMkvTxDGN6SSaODy/T0jDnIz/mAZx0rsaCjzRZn3pdjM
fS6jDHUR4Xcry22bZcAoNxsm2Sua8jJgOcBJWyFTjQ2dWsmoXN3VsBACh3FPxBVWApRziIconWNn
8D0dM/tZ3KpNMo94lUdONqJemPzUHoOIu/ay6be9KPemif4d1eM5y26yFk5TLaFoC3ovhyshjsOR
YIO/XQpJMiK6ZQnkr9DLpEAEamJATuxsVfkPDONjZmarHq/5TqQEGbTe49OpqE+SP9unuCSKyLHf
VqAcM8igefw7FrLAPX9OLK6FePYlcTsEgwGTVu4LZOZ4X9zpLY8FDITbz6GJT6KzS7LMBwdrrMUR
hKTWPFmXFXSf4SDaVfvxEMVEALNXCH+DDtgkplLD6i1GE1/903bOJvZfDJcCOBC7hgz2mI41sRlH
XQZCT0EzvQ/VmoszuRJP9LeAVy3JrPb+ApmlaNx5UtUMxjRhvtMsO36lvFvM7/6q8ub9WbZUuqub
kuk9KOgm0uyTpAfuvWyPmoGReBSe1EFnIJr+yxqTOR52cGtJC/wnEjm3LYFSrCqVPpcpT5EOELdg
sLKtRBbsNYBUDLwKjZcBJ6jOfH7ftl0XI19e6rzsR4FKQrVAbzvQ31/ZtsIG4nELQYtv3JTiBE3X
6/PGigx1r1XuOhDMC2zIvdxNQQcEOxTKke7Chb9o5KuWpyXD9nvYYbcvqrlWxpsW/Yfl2G/WHXYe
O4FV6oWLVzPz2JJWRkdvWK6lPwB+pFDiXaXuuIuKxpAKl0Y3twrnbnPJh4f32mDHEqZFxIzfrP9x
GJPpc6yIQ5hX3yXW6GGwDsBNWUQIHSGZXT5vFo3D/oXT2vfQg6/BoacZvzwViW9iWqqNd91ZtPXC
SlU52CwFswO71ojM7stjdA6x0llmYJD3Vbq3M+OtgqpghI17H+WGvPAnmtD1raLP21HS55lXhzLZ
PXFAH1JVUxbvwL07BZPJi6Joi1cF4CY6l721n/w4jRNitJ6Xc1EF+MnLNgCquy+90wmxbkoBrT6Q
Pi7kYtw0TUGDiDkW0GsvorVdMpn9bwWnH7LY85CRTQjLHlfPygFTP5uYwuVOMQfjUj7reOyCnzjV
JLAXWRq8l1Wnf18NYbDa5bmK76rYCKtmD4YnWJaUjFf08g7CDr7xrYHMVMSZYW0W6W9ioHPQ4wBZ
w8KruxA+lmxZ0VFxhlor95NCQWGhfKErXLpaEEaDcn+xsFemyhX7znDvq9VOFF+LnmuAI18wrYdT
/AwbBIzwYIAbu4Ou5+NL1ewGKst1p5fAmfJsM8Fih1OKqmj8zdq3kGOgjqwbSDUPU0m1f5Cc53KN
IIkbYBBOpYRpBCcbZecilwBBOopiCZgdfpjRVaAcFTMw8AZvPNA87u7gG72gy5vjHEhkOauJmZHb
LijpiNdutr8lWz4ddy61uWlDvfHQoxusG1CtLY/eP4tUm3JYDuyHtBlHOjtHVNyvXYamwdmv2wLO
N1hU/5Plm0X8535XhQVKbYkaH9+hQ0FCstoDFTqDSt+tmxYXdLJsRbei6UByekjq0oNXr13Rkj4I
weFxzkZiqp/I1av+a/QfXwzH2PrcgY9PnqcmPDpp0cITEaMdL499M0Ap3K0K7EWLynR/DOaQIyqN
ihYmQhKyoU5sVAdntFL6GA/HHFw/hCgcH4tmEFRJKXNFtNAzA7bN6gPbmENYhcYWHBqaw4oPtCWZ
Zz1VOAsHr0c/aaqDlrfyPMHJutWkQT65QgcYK++FnepjzP9hbrlQyiMUdoJMCfNs0P9bHMdmPN22
PU25pihUNPE08G20hkpzFnbQGvhnymGpNkuFpmtRSavlHx8sLFXrJwZmvb/yPMUvda6oN0uXRGer
QiM9j8knhTXpvZd1lksPQXbgNUmcD7hps8Q9WlE4sA5Z1SaenquFn8uPaU+W6NqXObfrGOPUHeWg
nDc4vq9LwaGKKnqs+u3J8y8H4L8iZ2/nqivnQ5btLFIlVr5xv9iX12ZLZGMUoCvhW56MPJTDI41y
l513DrIpo/q1OBkj9RoBtOJn+AjWNhuPU1528q05bFqBobCzCpuYvU1hNkeStZw0hyfGeZ1eyuyM
tkLRtlW+nuQN5O/wv6aOrY6AT8YsFWE9AHq1xRA42Lu/ZE5KgARECISs8rfsMdXmCY+NSYNe8ync
w1xNVR/XIHpCdT2gzk+r914VJMqMk7o8S4UMDHvj6ROCV5a4O6X0mhrfNeWoyXChU4sTIvzo9mj/
VKUVDUMHMmmbSEW5C7rJau6JpREGmxXa+f2GS/GLD8FXnM7ZVdgwAdX+sXFpKoaW3U5ieTitLO8c
4DKhE66FKitMqUUTJJKws5RMf8psulMENiYR0OG7Y3WwKoSSMrwsZNZ1KhyIlvWvj4ENo++Ori+R
AOg8jPvOWwvNzl3H00UzHi9kThFrp5x///T9017rN7tLVc+zp4YEeIrTgogIezVaUhWwHeCJHv5o
ygxbh6ALOGx9MqHDv7DwFgT95a0kAAH8jFbKwuOiNv7MeXJEACgBgAK52VnprsQ3nP0t/oSQEggj
bv0P2hWL5OqE22S7xdOMftpW7z2Pm7l0oSqocw6cNlFaXdvgj5hRSUjjdDdBrdZ78MO+843L2oAQ
ZJnALTd4u8vedaDBNrpG12G6kBcz64HPxdXQWOmMUlVwJMOsnnW5IbTSotXOGhoWqz0Tjmz8AvzY
7dW22o+sYUqSgPkZtzWnfMAuWEMQSOmhjScqbkdYUg3ymBB96trAccFanpy498MEBTisOcQ+knCF
R5G7GrnZl5+Xje5bo0havea4ey3o/rNCqtqhwSLNVCv2yooi4/JZj597j8skAJh8WlXRa1w4Yehq
jRXKf0lWg0u9dEv5JYc8zUR1fLyqDAeeYRlKugrMY+tOuxUeRCn+AxGL+migfmqEGjuT5jsie/Ij
VFrrEl0zN+ZHQCRkeBn4DJzlVLYEgvsrRczh6I3xXbTnOmDOnGdBLx/69nCUWhtcRF/V3TUlLWwy
jlglNOQsmKr2MaAGM4dQvtU3O0qaPeRt20/ys12jUU9ebDNP4tQ0nZm1BNr96upIgt23Kzl3tB93
rSWhBk5iRJy7bS/Y3jYz80HrhwCg5izRnEah5Ajo8XXXyQtQnyDTSw1+OTyakdB+VeLT6cWXBKw0
Qm12XJtN+oGE1iMT+J+nMGkh0adFRAKoX0bpFFoPexjjQy4kVBPxFXt4nF71SKqQEXHm2I8DJ/WP
PGr7bMFzOng4crV+BBmKIEsOR7QM8L+XFbmI0m0m2ZfY/y3HlxbHDiKi464fndVT/bxAwSiz9At4
pKbHC+cJWxNr8XOKBQa9vc7PS7rhW281MG7sWwJ75uR0UgtzxFQODR4ORnKLYlVJ+wj7f4OrBYTg
a57uXcSXy3BzixocwccsetntezUOzhu0dq9gLu2OPuwDmomU4ktpWgT1o4sShlMx5dwVtJB0V/Ed
TGDesRlDRze1WhXV8DLaMBuIUL2UqLiTUIBWxx5wFWU26xtTuy/yDvWvF9ImtplB5Kmdly21ORSm
FrTHqbvgrx4JIdPlTr4VCHdzqnFPoS2aQBlB9xXdUPVvGnyKLlHZqvXgHNSo4gIybNSYe040+7Tp
URAsgB0UVLVGv7LnPmDgaf5pzKKXkOwnoQEJOqcpS21F2HjvlRsvqchRR4Wnsxsc51Zb+3x9gsbO
0Wgo/yd8xREtlA/0YfqK9R59IpNeL920Yz6aSGyJV3PQ2ayRMIlgKamoqFAy4IHyE8/bgJKVrPiM
xoYSEp8jTfdbqNUWCg4USQdomHmSHvP3YGJ6D+fw9fPUKcGlO8HXHPk5w8eoSC1EaNQKVLiGIDrQ
7XWSvDYI3BVy7P/vrpHz0amaJAnMq0uV1giaIkrPvAqCdU8Qzk9353Bcc2A4k2KcxZNn/swyrWx4
FR6Udg2vcYu4H8FUr4D57AGkbUGTnF8wGuwlgWWUOpkj7n9+0dnAtUqI709meX8osZpHxNIJOuYz
iV1/ctrdJVxx2Vr/K70t0dapUy1THfgtDyGzzBgtHahe8I88KThjpxN/2hONg3AB0F0k6+qZu1Wi
CPdGA/KQi0YsiHIvisB6mpnQmdGm89a36Jrxydfc+as10vcZX75ImjrZ+963+HBG2oudEIrfzrsL
FquZaAEnN3E1qEmHVQSZA8lNYX9dnD6n2w+L23pfKgwzUX+nlTR4rSSXg3cO+KPtBGFXSrk6OpLW
uFdr3FIz7Ge1tcVJCcMARyo0JGHHhBWb/1mi0gRJj0cTZ1uo+VIdDOWAa8WvDao5iM+Z4nW4fT0+
6qQ6+gQYMv8z9mSdfCjGleF2pMF2WC2O5f9MgBLJNNLrAOSgFSdj6rdCkfe0cdIkEneBNKvjkhoU
uxThvoyIO0lT9tjBOFeQxPbY36mdVyGWvGaj1l2iwZ8avB6gLL8t93CG53IjTnpZdJGbo8rChj1s
RJIiUX48b6jyxt3DwS3pC8l+mgCnIsam4LuLvbCGWdHN9QXS10DtR8cSWP0QyT+Ec+h9fJJ1SbEk
dxUkeCqfpY1exeYix9wgpv9Fx9MxdaZT03+NQmBq8c/xStOrV9Lnrojyh0+Ju/9ftYbTz9zGoV38
54umZ+j6B4YevL+2bm8ewos4k6nP3bo0sof5hZ37e1bEoLlnhncMw7h4cPXzMWYRMOIXsi9dI9Xa
WvWgEnxb7oY1U1L4RHir3aD9AIhZ2BPwfCA6vDFb6I1cXKpWzlk0OUhkCB1qCU2VwPrLXQ1chWZo
1FGhp9MAUxACq0fkArVQ2iTXJQV0r1MuVvBD50hfWoIRpNX6QjQ9HM5RuG4PfiZrNtJyNPQd6Hg3
HLRKXaQPd46ADlTY/8qz3qv1UGfhlMTvwT7FF1ZYWdYVLLHIaQrR10lM9sqfJeE8xjPHvZjFim3p
aJp/4zJagb2LnMuP8YDj0OYgao9VU2EjmsIcyw6WMiKFhBzphC0+LsthaSdt7h6kYOZvAC52qOsF
quQb2WKIkxFYzguF3Wp5BLRUwTMVXZemE1RQe0nDByHjNQgZyYhs0KQ/7/j353IayodmQumb0/Qc
LbP8KY63DLjl8UAxg7QHPzBCr7fAQe6gYQFfKrGpbdXmJWh9VkFbLuHUVpsrImmIyZAe2+gBohfc
rpw4S2YN3YfwwK+vjyPgc6YUeS9ChBjf9EtQpqbGbp9TnRVrYghtw8P/p+bT3v0+D1nrFZUuxzpz
jmSF5F40tGQS8cNUswG6abLVSG9QwoIRbNQjPjUFNKSPbIt/KDuDQHXSob2kYOjaBMiBZCwd+Oj4
hsP5vs9n1Fe3gfAhpVJCmOkkHbP0D58uuA6dwHVMrFeRZFQeMiHSnhxLOTEwzNHk6XvkyQ17sgrG
QP51j1SxtO8V/G8fCZmNdcXqNGa7uAVlcEj4fzPCmUwTVIDtof11yQRaVBFkBLtAo2aqn0fK7z2R
hntss0VQjpotUVYKNkwsM+LZvZtOULE0cCDqEiJdLP7rBu+nb1BS1wnaFBi3LutJ2pYslYyEAU2C
9wQ28xrg0KQPWai9ssqiVkSH1MG0ix9d+KuoKKAuiILnmvpm3hZl8TJiFxb4DzKw099xqgtoygvV
SLuh4FVCp8YUR7oKcn4A4RfeOJ0vKSc3JfIs5Jscz6t4YwScBJxnhtezuJpNE5aGMP1Qw2e6EFuE
XHujKEHSqnEZm/cNQCN0Hvi6Sf5rnT45mqbTvwAOPOtewUy6DOiIFxyNI0WPCPjLJM6cTref0RkQ
qyD1gBTj1YfUEQKITjBTuAJTi26dEx1VbisKMfd8pOuG5vV2+Eb4+hRU2B0u47qYXL0li6bDcad/
7m+n4WrUKhavGm90PnTqo2yE4DBYkUb1+CaKkOegF03tUjLCfhLWcHFHGbjHsir9km+3ivlo3i+m
uqgjpNZk5V0h2uTZ1QSLB9eK5b66O37/Bt053TXpmkr6sY1543GPU7+0j4rYiRGu2gpqnAgVnu9I
0xElAVCGYtZl/PtNn9T1Kt85Jr7v4x5AGsUN8bMIaYR4KT6ZDWlt2MfOAbigHtE8e/rggqh49b/+
ivi2YwRckn6KAnI3aaQqEpRzHLquYU2RCFC24oi7b8ZQfoplh9rcaV9QREzSqhUTrKL+gKYp4TeD
YYJbwAJ1ww67nW8r2HSGTtPo5QlnGwRumj9xrJGdWfBVsZv+cMSFzSWg9RlOh5njBeJp9V3OoHur
dXZG8ZMvi8WtRE5Bcz8Ha3AlUTlnrRPtcAnhVEJ/3nNg6/n9/XPtby0S4ztlkSS9LUXSfOIDbMi6
NFVCR98VzzzMTc8gT/LPwitdN0N2J3JvcVB56RtrqO5x/ydHuv5Nex+lLaxSqcvl9OACktwiqGlr
cZAmYbxWvU9u5PRzp/+CvoEZCteb8PpZkpqP0+VPuqUP24dJgRELvJPozyw0VmVjNY82wloKLiZ/
dDX0WfKclOC5xeSwj6yhDyXluo899mVf2BdtZaCr2PK6HbA1aYwNzSXd/0YD8ezkppP4c382XKt8
YI6E+6C6Sl6/xyCDXHsN5u69AMKuHxQ2lXvlv7jZi8APjE5ml5Jz0luDWCe/Dcv7w723lUbFGcBi
30RMMcjllnCdCWNwK3C34YdSGkiTejYBKl8bUt7YZVdRvCPpjolGeqON6Ot91O5RSP4Uit0/zMTd
ktDsxBFJdZJXdoujcj/m6QzE+ClF+KYahJCqqXftpgi94PsGLnE2aW/zA0ynyPu+wMjTL+BVmTfl
6l9eQT7/nvLFxdxXmFT4Fm1iNgRYkAzfe/7UqZhAp1XdUxbau7DaE4+5o3vge3IBzUmex3Ktw0Tc
jY+FPPwsXmKT/Gy2yvix7+9NoeISQ8glkirRyfXlMXLiuiQuCemDGm+mGGzaDDzInvIeSiFS6RUX
5PXIwTJMST9PkLj98UbdJSHME+BFxmvaXjMtaaNh/hufKBJU1I0kwwNcg6l2vuqJJ/xYgsINxxre
yWT36ztVYpX0MyxJdLkRzqo5aKMQt+3ykr68L6DiHJgI3omMprpbCn7iL6dVU1j6Uce2IxhVYXHt
iQcKyVGhJzuN+ylaltEyFlTbclzRw4KY94OQ26MUYdkT7kdyZmzvhpKy4U6bhefes/jpCHBv1keN
duH9fvMkmRuasJ0qKNB9lE+lB3H38LylK7SLxwyy9vdSxIWY8+kZjd8AeKd2lS2qdtr5/D0h4LGI
DjG1oH3j6rhBkb/P0JfH9n8DjLnhQCLb6E8bNHPAbCH1QBxk6o+4YsCZt3w6JSv1zoGzcSJ+gkj7
IRMgm6b6KCGWDsm5+fnMCuDwbCLb6w24fyosS7Q8ubcb3z1v6SuDMfM7ajlPpzt+cMJRdMoR3zww
7fnkYOXgWdgVIBlbYFdcTTqAOqjEcGOG5XXOUG8tbZM5CoGVoSmOmkyEUhsY9NLaWrfRbvrnAp4/
jPR63EVvh1E+dQ2qTol9VMrfycQQoFd9GKQzHzevMtZCfbyYTPW+6nrN3skt+kaccmMHLfkNPUka
tR8iQMKWRinR+uKFZ0uQl3Mob3PXdN2scbLH3/XhgHKYezDpmEDeN/CtS13hRUsb0m9va16QcO/0
bKQwSVxCxdWZLqGk9re4U8jrUppX2oOxPGbYB6gwsiZiay5qBF0pN8RZYb0bnkpWxw2gUoZ1FWhn
MQku5BydwWbAyzqDq3//ERZJXU7ZRR0pDaqABeBim5bhWNsGFwGFFa648KaZ066Ms9j1TCA8nUO7
qDhrnLPK6qDyKAUV4tMvbr0F3nzx0hz0Yj3hJTk64LSHNpvOEalJh1jwubgps8UAzQGnqWCReRFk
3H/xZvr+VLyOzlA8Fr1jPKEfurACSNkSkUqmwvtXDUuPqoHgsoumJueWRu7yiGk6DYOmgaHKQTPj
rm2RPJG7VfvSJVY7hg1mddDmuKjxtGTnEWeUeDZB/jDziVTeZPaApFAdVRAaaWh+Pg3GIt4Pvw9L
SKRg3bYSHSe9DmQvtyY0o54vWB3+zHANKtzzurLWaft57ZSGtA4quP3I6rYOozDNLgZfYdLXQAB4
XQOYIMME9KNht/7BzMKZOUBl4fDhe7Kx3k9b8WGb2X95qf3r8Baa1ZqzDBT6brXTfjsudLBU22M9
MHxGwRjZY4uMfVd4+zLJJBx71JiM7XIrLpqKw4AFZeFJ50t9YbZyTs0O4NJJtsNeBFeD+wBAuhe7
Zk99HoCuPL1JUVf8CF7XEu9SRqoUAcBzdqjhqiNbCv3jYsZRd+TpMUOYSvL4E+XFE0QrMuBOZThD
0aOEJ7gL0l0xjv7H1cdqzRl2XHI3QkA3bE8x/TPL5yma+rqKnSUonYxE6we2vbClITm/Id1EbfUA
uH3f6nh+y/USodvItSrndEwykg9/pPN82txJMK6aeGdtVALb5GrnNDoOQrILtHKLbpHFT4Iw61ky
+tmmLgkEByPWekCdn1SiIveh3+mzhyxf5y75rYJSuhtQjrudvAib+ACFnybOUr06FrFXBXP26scG
IVIfCxTIKAsTseK+PXSQsPKqr6g9h5i/8+aVL0gaFykP5nsrYVqYd3W1puO0dQVqdH9lxUYz2zNE
OXu2sQMfz6rMQv1lPYm4ckVJu6/JDywp4CV+hTBKiHH0ym+2Xwl5x5sM18E3eAjG7epVSRqdZAuU
h4jsyUw9eZd9HBbdRHj6A0tWjcjX3lvYnmfCNaKms/xeo5DrcJvKNjjc9ocNOUAj+M/GdQtSDiW3
P1ysnj12je7YS9j/I0Rx151HIzfSrWzlYCQ4scYVAIN43bLvahqTtR+lY2xj4g6SP+A+ROYkiFtN
XjrACpRqnidLBWX5PbBt/y6XYGn2kIMHr+ok7DjwBcxqjsLqThtf8szwunvz6xVeDUOE737WMqwI
m4LU3ZJbfgqbfFlYoO9RxAw30NP7IMvsO3xCvtzNAdxl6muMn/vrILCQ+vp9TCoqX/yKUgt0lj6t
Q1W/i3Jj/wAhZKI2WphbDLPSj355LsN/mNlQrPNPoBphSxmPtoZRPWxh56Enr4S593br4CuRxepX
rh/Tx7EuQZ/Q1psygqdZNj3QkZHL5mbDezhwx2ut4CMpStR7SpGXK1R25+nfANhld7Ul8HKHmwdN
vxm+8zjG05R1kAsdmiAZ6HRQmEuCib6xUMyNGKBGmS41uagjWt8eCXdVSVVZe0xTljODggo/nvI/
3zI25tQCDVs40OE6jCCPMD80/C49PmQHvkzlqO16xT50e8ZE+AuX4sJdz60DBmQEK2jY/Zuj/qLo
FUt9JkFDnZOpoXYuJSKh+n+JFKmdLJEbxKmd76dr4I6AYeYn/tbBfaISRsQ+nidPhQdRl/eZrpUM
D3FsjnHdyQ0CuEsM66tfDYolO1TbKAbJ4L4jfLXOTfNFLdRtHrzsfatR00qEphlNLulJ5J8HBXEy
yKco7rNAm+XSVDAUeV7wYCvi9Dvd+CVjh6Q/XEl8Y6HNTFqYJBu/G8rHiviqePMP2U+DQqADSqQM
SuTnlrYCRANXPn+/8qy8MsBEFzVq1x1wo5RvJ9zdjMk2MtXwB/GIDrakuN2mlLyZEezdtjHv8Mmu
ObSe3EfqSBOR8aaQnlvt3SXsPwRwW8Pv6RsOtTjPCF6jhm+e+knjmT077b+cLL60ow1CBiwDlAgl
g3VMsIXJMyuqoMqZqxYjFfXokTR8BG0PQOtlSEN7pEXS1w/shuMSU3Knbl/9p9JvYmR0wL7RPLlZ
FXdYLsAhiZoU1TTHuTSyjCn25fdXcAuCLteXgfjHOWErzvLYWlkerIXY/h6IUX+diSHgq7F+oa3f
h/22AHnXdE8No2mCSDipg2WHN6724ewI5B6URqgx+Sk2Q70FET5QlFbgjOzkNefuHPS29McqJUj4
GBXc4kUQh/Zzc0qyCGLJ90gWCYWTx0JI2kk5xOBi+YvsJ33ii4Wosdb2RzJYePFOm6mfbx43SRY9
BrSEypTI7GI+84CbEIEqO8HdnNYJitC03QghILq9B0yqqrXeTY6cCARHDZT73hgY8FKteIKpwQsO
pJFx4L3+1d6ayItL1jnLWS8gDLqsx7oeUz4n5eTfUB4K9eAz0pgR3tYRKAtjqJXkzFc1d2Wk/pZI
oHQF8kkp5t7l0UO5Jbpds4rKiUVLGDM0k29YtSH+hg1UHnLiutE5+Hsm4Sq9ROOKG7S9RUNarXTv
qGZOLP1JZ3BAdNETduQwrU2pMh40UraBU+ora2MgRwCaNocDyFL/oIwYi2OFa2EimRlvoIowNV8H
8f/qHhSvfAoQtgch72JzPBjvzNjGWPPYDEj5MQXYGs1Sr/R86GH3iYcEHIvfwytp7ifaILy/BWwU
aBmzlRefb5tN2Ps+p9NY9IE8Zt65sxWI1/5WU8Ed9x3qZ7focYcyrQVuj6k6XpwrabFcP6EJrgth
+YOHETUsaQ5e4rGUhMmix1cccYZ7wSd0PvYJbZpCLMeWAjZsU6Lsl7+pm4gVRvRsrjNX6rPBc6YG
hXZvTDUf0C3JNx8iZArCjkRW5U/w89/aYTzRH/ZHzrIM7cpF0RXvb5SJCIrM2XmCJKk2AK4/kgeq
FQkeuOKltkWxvLZiwmSAlyVai0CmRkJs3rqOFVUF9GOi2Vl6SH0QOO5ltL8D+pxKPHDVu99cxHT+
huDv3ffYJw2ZYtiQdawF0bux85KDxaUbo3P18WF+yx4hT02fNzNEFAmtqq9s2KcCjlybh4oTmSct
Ho/B7ceFqbW4Wu6ybLjtGpdimgbfm6PO9ijCSEvgKkuiAOpu2G7AucCjSnJacR82JsSOiTots0Yh
oghdoUx6a+yDtKeCrUUT6OR8rqbVQGzQjo//d9G4LJRdWhVj4OxYJ8K4BGNwSVpRDRKvTXMFsCS7
hg7UczVP8jQS7n4Jq2HHogGeqkpgigWyL/HYQ3tNx0CuewmHd5bgdpk6YojK0Eq7kSSlfEtkMzRm
6jDLPDENsJceUZmcVwe3teIqnGIYDUgdcr2mYMZsTQyVTB+HfbTxo3c2yXm+ScGqFrAqc/2Cy9OI
+hxCqeq76eydqXW+7ZYijz5QKVZ+LpGpQj9NyMHO+ev/+T9k/0v+iJxjA001q9peKGDH3E5pNT54
YlCQsMa2IiTi2sPCf0qT5rF4hyLMvdFrCMylhSbFTJRNNCJoyNCqODg8GBHV5vjMUweZ5pM646f1
FC9YmCPW/Jd/RXfz8yeaNGlyXhkV6cDiCjAYD1b8Ow+2N9fPST2/XtsD7x+++ObF2kovBP0go7+q
Im9Xt4sLiDOVG8dzcbVgyi2/3yutpkSewvusXyyxmE4AITRhvPph9TSdeI4SUPWaUkGJW50OeLm2
iWoRtP+bufKhWgb8Br8ORH3CLhy4cgqKNhuADzTMtAxB2l9aEUc6rJYXfH2XGsZrnxJkdkY51+xW
BSPGA4cgs9nbVhpkJjBNCtu0/4qDQyLFHMDXAK/l7QEJZkyBegWROfo6Ad695oDREDd5drrkVJC3
Jjti974etNCtlo758DyrLyxwQALf63MrA6cqljpz8Xn4UZLtdqQFavbyLoBxoHgJavg3xN2krF55
5ZzOv9yb6ImeWnIC7Q/o0VBZoWEx97LhgrMWVts15FDUoMP3W7ockx2kvclAtYGKaOc2xPGVS/NI
ySknuzTj3p1IsWYE4/mgst6fE7fZTRZ0wIQSnaDjoDZ/k2dhI+AlQJryIaHlPenYxyHAoc99+sMk
vY1k3XZSnGzNWL/K8ewIVXnnjIc1FAhCETWmfqeuPiafC5viiHKGhLfjkcXFAAKZsteFpgfqmOoy
BaukjVBtq69tMXDVhQupV2W8eYP4tCArNKcYm2Crp4zRR1Q3/ClFxJ1hmpCHUshUEQLWsjCVYg6i
xeZ2avSebhnlXOdSJlyqSymgz9akkkQFPjuMhvWch+FxATouak/ouQkw64lV0aDIE1dvThCF6Lm8
pcIoBuYQH66AFloSObyTGG4ohiFRXaJI0bPtmUocD1g6POF9hvHi+Y7cTHQsgWlaYtvcc4GA1v+8
9DowN+vOQe0XQA+DAk0aemKlqrJRquZvzVXvuJMiLq8h+tXiGJfQIqBtUKbWFSsrB53dTibPBpJn
Dlojo5oyV6cOJ80YJfKENlapHT7fDa+7UwJsvjaawDLdPOD5EYob016G7wLi/52ZhqqF7xDNlORL
u2PNFAYU1YL+q9oxkHSOW3V+uYBjQo9IjF2h/ICpahw8dx/hDMtRuIuGFiJRt+FF6IJCD49r3xim
ZGL6A8du6lTzoUFQxK2lGReLXMNuEdorvDACn8mX5QagkmR/h4aQMoptCpg5GDGVVDq3Lhqklraf
AKQSGF4YHP5HOob3c+LmoPUPyqW9Gf/Se23Rwa/L0uJ4STatBmbKiMWThZyTrdhjxadurRGR+PhS
dfpqvHEHxmYhP+1AFT7R8iB8N8cg4+CJn0CGw6Ko+UPPeUYYCqerZGYjre6D9Czv0iSzkIWeJ8Ai
S+kCDPxXyqJh3pWnXk5MAVc2cZh4wG2mZ3kwPQEITetoe9njMou2gjVYNgIPl2bwT0Me9G+gLt+R
MR0TEjf5zz7h4kmwBi2bstdYzJ52UqV9hN0jBs315gWbX5Q0MJMPWvig5ZL68dqRhl0gHZLyWTfW
1lHpeNQKy9jeYSa7kHByno329ykluwKrBkgrr0kQ2xDe7gXnBX8Q68oqVqnD1c7dVpzNTD46qat+
WhThptE6gfyMPbwzq1B52MedXKXmHdO145eU0wCYSgFWZ/AJmnEX9B4oQJe5ywlLvTQvSdZFcpxj
MTHUxx6n7yKTASUz845ClQRDuQSZC1Z80aqvncovI39T//pZuwzCsgJGvWvfTkBi9LwreI7Lld71
2dCVeQomiNfmo5/ETqGb/CH+RmGSawdVUr6h6AEpH2wvRzRsURVW7PaXlmPk4c8VwEqO6sWWk3Zt
n69niOm+Qrf70dI8c0ChOrtDQP+Vzp9657QQSztyFkdHIoCnANNaLVNxe4KcEGO2CXgEK4hj4rV6
BduSwvvG/6VSakx+b9eg/NMvPYj/ue5ytoakDoGIpPHomSVNldwr7nJ+FqwHfmCmbjIF/uH980o4
CbgHyN2vlVR+wBaFXjn2Q9FSqDtLH2YNezSsDUWSImtzEnFDdPzmUScXfzAnULwhir+hIaR99ae/
BZkT3uKLgP44boCb1MRuXi3mUeFkwN+sz9AAvtgS2eK8MGLpWa8Yjo+LT8+W3POZM9gw/IB/IvbY
UG6JNraU9+4IvPyAWdNzaOKUhSzijL4iJu4IJ61pyD24gDmC8mcrq0AQI8zycOw/D7jZobrFAyVU
UXQJwFGqnbPwKonBK1FH6qa+2m0rdZfwpQCrmKlUf4q8xkGkjGTf8a7ZzMSyVa34C/wZpCzqKsDJ
bWn4WGKrQ//h2WmDyvQVuJJ6Y6mKJGuTsiYUwfW6EBEHuztPJ7FjArTAknH2BPuQCUkctL2VZXZY
wwV/yMaRr23uJjz1SEWUUkd8Y8xuiOKXlX94S9WUqnBiHaNucSaw7DoUQrnlzDLI05kTkDcBuc/+
RlUi556QtYqe8D7uI829AcA5Zz5NXDmJ29hzUoj88dcsxre8f56ZTCiGr3GzhbWv7pCiIFZrqCw+
hsNagQjER/daB6QyLIuiAo4TDA9vgIEJiSS7qua95+5TmvWrofU8R7mi5Xw/8THoseK+rrHEkrY1
54N9jSr7Dp9KEPFsIu4CX1y4ZIooGV5PdJn0d5jC9+e53XnqMP7nmNv79wbjOFarCMM039ylootf
WbMxKyYpUx+Kd+dvxmuiuwfgKpS+hJ2eKjbrvu6HwQjWLLpotgaVIGbYrpDB8kBF6hpj7dgDNkIa
0Y2i5Mza1LdFew5Mdke9YzSLYKdDJTnsn/YgOYg+03yW7GkuMPmsk7S0xmjURzbbVsjjUdqmcy10
0H1Wu0ot6WIvBYM16xwrkUyFehRE+ZiAHSSirMY04feRBg/k64yX3zCo/br2UI08ItGt7xZ4vg6K
N70VhzNZiCSuP9BsvjXujZhuBiKg1jg2O1GB9bPNCMiOJPGWQyanPH+I2XUW9toFmFSngeE0IsEe
wf7cJ5APQ+iq3ig69VLrkVBzwXW+z7LqjkRFTRZS66DB+hFzA6ErHeTGckSHYtvlzcRC+DY61t/c
s3B2jeZUkXl0spA8/57CAfOacODm+a9NmsWLaNem87kj42a0Y0Djr7Mi2TvZOs36u2VXuOD2oHC1
2a8ONhyaBsow4hNdazq9ffb7txSKhEsS/6VuSkvC2av81xusESDhxy4pehFeB++tmHC8R7aEk/VC
8hOF+tmW0Gx23SdV+OXArXEUTznXJo322IA21sEl8343LWQm/mPmtreogaMIA1U5eDS+CC6Bdump
2SL+Padhdhf8w2zJlNQeqpdRLN4UReNRXinVN1v3iN7VjhWYx5CODmC5fs2mH2ZNKIa9TjkGnKet
UNTieM+uHYnFDKX9rlIULvWabLd/KFvhkrhj2lfpiEhjLwbCQ/qtUhcQGXjkzLy0PjmI5UDxEGr+
AIG3yD4d3gXYZxnNnjcOHIpgufE40AlMkvew5Vjo8KrM5F9H3D81gEcLZTURzKpF/vdqG+z0CJ3Y
gYficuhenAY8ZnoUnaarpkcxi4JyUEVsEY8nY/Ai4qLol4wNezWhb3wvx0VVGiATy9DvsHyHEFjO
Ha0UfgrbkAjRon5Q3S2xgQY2nd4WeijoxMUqJ8BIZXs/1WWRqsIwLlDmN2zEfBoEZIfg/PAv8r5W
04s2xle1ZinlaHh204RxDObNwXXqrYRGDpTN9TEQ95LDzpZj8vcIMSmg2SacGaWCD85S9w8NcRIw
od3AbmllXPw9wEz9ibFh4kZBD2GeL9VxN0yGkHBfKNltiIuAZ22q1jJVoxsAwauHcJBbgNHLTaz1
Ul+TVJFD9SMMx7KD+IrcN2mGw+iUslq70N7GT/8GUTGFCweh9yaeFfiQCvF63SzsXGz4PSEMAGCU
PavDBZTJRDhCqeuY+q7Qqug3lCayNnhyR5BLDiTsSMeq991pJ5hmUWtl7AMU5mYMXOheCsczHlaR
++w0Z7JtKUU7LvkqqmE3a5K9j9VaCUwIkbAutztr7CvIAWeOXLN4IOY8y+6COn9fqZJ0tA0svhKN
UqkXJNPPuPkMP5qM+O+rZlFekVX1IiUcooYs2ZW+qK9TjiR0mV+5w7G+h+g8F6Fu7l0kj9uSE+A8
DsJz24UPyaMhs1m7QPjCP6jNDj91GEkUFo11WFlOq7AbSI598p4IV6j30QoA3mUH+vxYmbI9E2Id
HKvq+ALrzlWhfxixrQQECyjYl11rW0vBtxqoLeHD8X8NtJK76AAXT1QeG2cfweSmBqQlhVdgMoF5
rdxnzjbvEtY4L+SlPqSJqMWdriJbNceaPVczyff9aLKfh4Jtcls0GD6nGuQzmDB8n7EZsYVeojt8
l5KoN/OuquA59vlfn4FeztuxvnO4Kh4wWtahkENRfPvNSsMf0n+31ARhXhu9GL7G84zZDCLcd+3E
q4McydY8zYlV61Yz5Hz8DPkRZYDB65bZ7SxERJLKdd8j7QFglUVia04oFAb58Nhtrjl19/slcSCw
JVF5TG7Va4D3XVo/1XCuL0hB7KZk20/j26sVqXM7yiBJ3PWhfkPxDbWxvb84prd1sFJS3U5Rn5bd
ykW6hGQFer2cCt5nrjMTTpBJnOoYoFvjRZi7QmWfLJBXSJUCI0wWQC55YTei2wpS6BLE4UwhZ4Xv
i09jPaeFGTussRQmGuJF4Z3PgHGyQAqcspWtdf5Yi8nFevH48C73dmKTyFGTgVuNqinMn0Nyi5Eb
s8UlU4tt25pp+d30rxbMVUgR9Xv/Bt6e476uCPqjrIOPnSQC1xp3Ge9p2Et8Djt6XfSH0HENWeR+
37zndJHT0k5IB+cJM0Its3OFjaHZPidXacKa5vXOvZHWpjOojscD+UGZxJesQZtuHMneB71UWrHg
uvimsk8PsRxGaFRkEAKJB+QFrzB+QlGDzK3OpCwmGCdY6TCoQ05tocvocbAsaO0dBbVXAB0p9P5l
2n457SKpuOzRR9B9YpddEFn1aY+HHkHYvs5FnOMG+HmypmK3otUTrnxyx2Oi9MmI7JcA3FENrni7
lYlZ26vS798vUDDMQPX/5E+XH+aIP8mwf/5vWgLsoBHW+f80Wz8UY5hNPyHEoZIPjo30J+C4lYJi
1DNTj15QXR0Q6rIb0IzEPFtZFKzvcmTwhnU9tjpBxrKuPdUO6hQI5+j4m7XcSPIMYNtgy8xA3ywf
URmZXTtN84/XNqO3L1CRqMoRc5kAHXxic0WWcP/swoV/doMx2HBoKKWIGpjIbgHyxQC6oSA1yy8+
b24clgd0yypVPv8eB8HB2ZGWA7w0zuFwCXn8+Zmawy/1YmHP4B19HxMBPD6K14t9drEBh+86RbkY
nN3GIiKjh6F70Xh/OyZFGE9zepNovMGZR2SIgmdhyZ5FPnbXnIwKA5sqjfU4V4Cr90A2tm8Aoe7Z
vwAMq11jhcrMNnHXLeacfATgHpge9ASzA0hCvoT3AzudMUXwypUhw3x/hMaLp+oFjMW+QcvbXBm6
B0qxU3N43+UWmRl172A7qNhMCZCUUbFli1lITGDsKk9Xl/ZJCRL1LRB0Y1GMbdLmF8vnTTbKaNZ1
jiKiC3eVPEq9QupjlpiEP6riTC5TeOUcnRbAus05UAdLcEMd9qvp1mFkvQTvVJRlfzQa6biO1+2u
1KRJkV+XbroOLBDJEEX+ZoDKnCl5ZLEaDrlYPsg5O+bb8jr8gvghBtuU4HLoJwssGNoE39DbcYy3
CJiCJbB4j7anW+abV3CXVMpdWMpHH0anTJHv7CdVrrTIl8LC1FHCw217b+yBNtBseKAl/d4oGIlo
85TWSsSemWsSQXlrBgedvJE+Fb9BPuNHvhKCuH4XEsKZzAiq0z1IfTaO7qNATGzBNt/suJh6NS1p
q43qv6qI+ZT18iLskXBRyc6YpngVbk3VmyIju3z15Lphf1zxNgYRj1sMrJdnEMLDOtvvG6PyUtUT
5a14EY3SWL4jgDrAaGXa7q3i+X/YVF74i/FsWFsd13EQ0RPyQ47eev3YVFy063OxyN/JMAbWtFft
PhqB1vFA9Kb/fgsRKfhPdKaG0CR8MTm2Uhk7D6rD/sUHfspECuyqp80LES1W1nOPImCyTsfFlOVW
f/3k6R+G7EEycuzbQDT4DArdQ5FnPmhAmhLCtOOuuqbsidxUOtR0p3ez3xzyR5+b14W856xB5NsR
GD4kVLDCuCE9G8v5AH7Vwl93urp5g0Mzc/w9ZiwtidifVpO0O/y2f4KEQ4nx/vUAWIjPiAG4GpGg
GvAJpJohcGPaKHuOhKl62coE7T/z4MD3zdZA3SNgkkO+ODbyTgcTKoOI924iO+G3Rjj8LYmbJE03
ON43T5DSfEe12w9tfbclxZ1MKq0xKEeS5/l8HCHgrLSe7EicT+GPFqO5UsXtjP0i4lnDsigzcOH6
TN5Gw8Fgfu5OZtyA5PN14BrlmnjlCoBZjHwjK2s0sFD5dRrjhdLyPJ+H3VLN8kXWtiFHMdmsgQFO
B3kVJJBhh/enGBsOQrtM/YlgeWyWmBwGCNL6waUiYhlQGBNjePnhNXvs/tRgaoJmprJxrC9Sjfn1
v9Skl0bljdSeCeMUC4vP57Um9sPKDyhwjwz7EBt0Lq/JriXQxqid/WSS6xucrESwye9ZifzFkCDl
tQpwLMI6K7S0xm6jV2nBh/bFMXYLNL0ZArUJG4KOvEa96rkHVTUlkPH3DyZvV1P6TYdxdOwutDzj
b5IaMSQdCChBhATm4IPFRiwfYxNSAyzQbVYtqT5wobX/BgE2gEVUE27g9HbUgNduxWumc0QJTIv0
3u2wFPJymEM1VXPyh9CBpv6HCDOWBUiPdigWDLUT+vtqmDloLJazYbamZEVIprPbD78WAsq5HOAJ
W0/XiwV5ez6AJqevFRqGNKwNIeXKdKEsihQQyxbqpwUTqjOxSvTzwvUhSOcCGopi9DAzZu9L7CNw
asat1+ggg4iPlREVr1iviKDgK8NSULAZPkDD8iBXxZU6WANCyNNU0kJbuc/ax512v54hh2tJLsjw
YcxlAu06ItrLqGkC7gx0jRwWMEX+WnUcVVXyol2UIedfADigyvn2JJe4vZpEqVdUCYaSjbXTeSKo
HEblkjMeEqhpPrd8gelg+MJKukr04otcJJ6AVp5TJyzK+PvrNwnfNdJ6rGPccTnjXjyo9/5RcJt9
x8rpK+B97iISllqdUccx8r5JK5DtNNniofM7WhUZfUqdT5LtOJsKkuLOlXeM6bL9X3XrLTYMyMeA
AePGs889lYC7zfUYciO5luYnz1DYYZbkQ6YV5VBPQxF2VMKkAA3C+cZoZakPjGtzUhOZZaIvgtWX
R+u7qP4t6aIq3ZoKSM3OuT0h/98NrvUbuHYoS3WrdjEjCQ2WbCVJn6Pc/UaLqI8fwZpY5qviTHwJ
jywjksghY5sax8Jl2HACHzyn6knbwm8wzODACpDGHD1VJIX5GSF9saR54Fj1R027yFJplmTh/6L2
8LymOOJLYiEHA71jRRpLryjoaaiOtBAwCdwkOwrpNz5IgELF67PI/kh9OzP7gshOiHUwGdaKaPal
DsvcSwtW3qCyi3MiD7uvLYxvMOh+RrJj7m0OJrLt+OiiAaF8KPuFsAIJviQjAs279vjgv3Lg6gpD
cjhWBaBZr7JheAL4+XZMhm8Yzd4ERMovEoScOrHTjcGOJPMUMiNMSqIkx+3K2lOSUdUq5YtqV6Pq
CRR29gd37hyVGIGSwYiFV3wHcBa5LnqwPixr9kv77n0lzui7vozAP1nwQWzQZxUVLmmURPXnIf9+
tX/o9+5R3+vmFktwIIPbCPTd31WcgCWBoriLUAW2ZS2dm9JOihtb7PdlGBHxq6xGeNNaHq62S6/E
G7PRBWmDr4PCo9T4vV0oxeZMUUWsfy85eAwLZx6PO3Dbi23idDDGyjh+pTIZNCcQJ9sNzuV2cRPS
+9RgJuRTphErxs3SWZMrLXfrQw2zp2y3FOwMB//8+PnTp0XJ1CXMR76M/M1Rt5LenBJ6OMb204Ei
hm/Dxb87tsba/f07yuNcKCFkXqf3lSC2l0vExqwGKprzjbfxwNfgYYf7lMPu7eFtq4z2JdUJGcE4
fp4IjLMNxIFGVWbduDNzPhJa6ubLmEE3IjohAqDOExs1tYoyEuXhLPLMuH+RkvmQC8OLc9YJDfPP
Ejuqi4Er1EFm/ZxiBr7Q1gFk7yVJkQdX8+R116GVLn2atnqpCmUDyfGm6u++fwjWEsfb1/1R+25y
CsyS4Zg88fOMJyDYzpXcRgt6hR1Gp1yclyVUnVOWExmPaxUbmfSDIBWKJemWlGjpsU8msBFd1Jof
qzm2Ruzu/3z39X5u4IXN05mDVs+fLYJO2pB2miL4GXHtkLxSce4dc8Ko5C5Lt9B6sWuzXlY/nTel
nC6rBE62gH8xNBmxWDiLfla8QFwzvYzL/0fxM9Fg9rBOmD+m73y1oGMEDyd/pAudKzHt8WpkRTJm
Z7YotrO4vaEhj/If1fIIVSv9uWMJSkEXh69qtoNslj+AIcFU91fIJCABgdrryttjRwSgA1q5x+GA
gwmqYfaYQvQdkFjCzDk6KLSlNI7CleBMR8m9yoALkkQmUT6yw7SjCducYH1erXAA/m4T07VMfQI2
t13fSKE47N5WkEzGj50thYZO3ITX5LcEkGmJqo13q3bMQr6l6edVhByReqsJpK4G+VkGEsK8Eohh
oHpQ4GOAqN5nhcWLz6BS0ZziTIkTrHXPsNVqrx3I8q8lDb/c3EYDRRiuCHOobdMPAgzfbWcBFPuw
Yd2A/jymgM3RRwoUXwF3iuBmxWDSJmyd23zrBlwodLl0eajqs/otfqxus5zPWLCtvXl6eGUptzkO
QMdh5CDqp7MQmYz3CAQBTRu8PBWlGaZ9WpW2tIEOZKI+1vcZd2nYv5gOWnvzWbB+SbfGzZD6WyHN
MBe5+QBlp7oGGOHoioh42VlfILJTAMv4o9WEcE8OwHqHTMyat3dw+B4xJGaKeB3ACQVjv/+UDfR+
p19FcZHhWmDRoPujKfwu204Dkol8Tlg2gwaJZxe1JlLCsKkYBV7/KfCsGh/KxK4J0WCbGSlxkVm9
1GO2i0ZTTOztbAhqy2HzcrXF8TZ8fAfNGCTRCd11+k98nAuWDJH1qCTNbRUZ8jw31UiDGPc7dAGF
RzYO/JymG4fQHMT0tK74a3rPGseD+OksANqWsB9lx3pAJ9Ns7mzj4i/3R26j2AHn38eMzps9n7rS
B3CLlQYqrMUjzFiKVneTOg8IIyCiBkWWJ5Uz/k6dYj1iSb2BBmNTasgZNAJeUep2p37fcum4fVio
U8wPSZ0c0TE2G/xbHebB1bqtAiO24qhFRyDy6u+GVrlPAzcLeX3wAO92tPhZ4jUH5jvdk+EbcHRV
lKlMUCfmyxrh3UIi+CEcue9/R7F0pXlFiXDTPkmkYujvvfwwF2AuMrMmbE4YQqb/J/gM9B/xmc8K
Agfg2z1T1Vg+6PmYYLVfr/XfV6m4KTwRvfC4UNh+REciQVb24QpSuxDyI2UaRHilUviw2ECTS4v9
OTaP26F2Wrt3136L/9xbU9HKSwQ8k1PsUTudI9QvsHiIhq+whxjZyDbYKL5vpEHsCK8QX2N2JxEo
wpolVjaIAYXDby6zP+/sSKJBjoBC/ZBb/6g3ay7pW7e7k1bhMZjv1+KjXEnmkLq4x5uADlhf+WwC
oVt2Kltx9qZ5+881Wr5NYzupFATDq1wg3rDSYL71mQKyZZ5zW4yyu8YeuBAkMc9MDkPJe+7+/3Pl
Kd5iYNgVcb1c+517xw118ynpDtpqqHf2zb8Bs153oqguiOfX6lzYM01YzXStezkdtI25boEG49VD
wGan3EMUkwzQTOzfoRPkvF1TDXOKOpXBdZz+HHZmMRubnU0rPkvoUAA7vfuaIEwX06Dt1cq2WwtH
nDCo76GSw7eRBgR99UupjNBHKFcDakJS1t1oCjHQ4Pxe7zOYhR02H2FVpa6EDvQ71mtSKsJ+b4mY
Ny4FuTAPGpfq5niDfuKUsdNN4od9D0c2irRbJ+lx65eZ3In49jjQ/9LoMN0pt/73L1uo3VBou72K
uEZdF6LOiem9M8tXTvoycTT8aEVaO0Qf1C9cwpB7vGxT8aHwQdpspGpJRjjZVoeDQKrHKa8U00xt
yndZdoDzd+S2FPE5iS2CArbfpMMLX7cOCjfvuEIohwyG7hnM38VlP/cmDuxL8kA5DlyC1oolD05E
r6fB7igtOHj9xkqjefZCYKIHelMzCYm7iXQRCJU6gyRnDHcRyEH8z9bYJ3oO0uHmfJcbSoJKnCf5
IZFAm1Z6533J6muCtXEy8nTnxextYGIp+eJjuRhnt7s8GBUswP9BIxE/5Pk/ZjGXnN7pnm1J2vOZ
O0MzMojPsXHc6YlSnBF+2C58oRXaJbqhdXaIzbMeF05HdbMMuzSGJ2lckzQCYA3Hvfphzlp24SHC
t82tOisbC0Rdbfa489xZf8pOWXiGJpMQI5BEBiFEcWmBpMNe85zJhZlRmXxEChpuFbaKVDYg3ymo
gb0snpQAzmEJdIacJtV4t6qw77fRbynRvA0KnBfSVK+P5ZmlxPAvQbMlhAmpedTqBzx7v8t9D7cp
Z468oFXLq/HWzosrCVnCgfIhljxb/ZACr7A96jx3apibVuAs5jcsMDd9JG5sWL0KPmsw0sCrLLJX
/Vvotkkiwez63hRGlQ41sDiAS7UuN+pyfotFldJdKMAx86ZSu1ZKhUVV5ZXsZ8mEVpHThBV4B7O6
DmTYkpMGgJvRiXcw3BubxggFbkU5I2Xffw+2ztaSmHxZ8KETIPeQPIvupsKrshS20U12psFO6m9L
TQd6DIIUbp7Nw5f3YirpSIMQQ6t6cqPmrTr3aC6Oc4ESDSorMFr+JbOOiIIdg5inwpLoWhPdsL6b
UfkBSvKZdZLSSU45V5Hf3t4/2yFGEK0DR0rQ2B9N6TXgSdEMNJ1+8MGiHDARq3cwCP/pCyFfbSRe
HI8B5kvmLiKtzMdbRpuxBOL3xDbenQMni7tQ/0htlLGBnJPcw+PK0FyTgpBxp5C6DOnRwOc+4V69
CTSamsIjp/ThrsLRVlLTwlDr4OU+etJl6GjcNQUvU8DAAKxiLladuknjIU3kPT1+7keuW1K4d7CI
6mTE48T4LBN/dD/axUVoQZ2I+RBWvFGNLoj7GtJiPkZYBV9Olt5rK5I5R2LUeYg4OTgKvKmENdB4
qL9KN/pHEqJFUkz5pz5Gy9aRVTB2H+9PNdLIP7AKXfRA9M4BeR8dSq/mjqwAcu0P1DFO7ktELBc8
wAez/fWbGC5C/kM3UI/aVohtTOTDlzfZXV5p/rm0/Jh2+YNXypuB1tDVrvbllSCqa3QT+gX3GfPB
vGJhzsQHeYeG8MWECiC9jYlbWJNRyzgrMGAGvNGRvqxo0Z0xMSb3I5YeHMTaoNCYMFpwQWhF6XIr
VHaffh7munpDlQMC2myAJ1i0uV8T8zu1GrIBBV5PLXvWoZVbDY0SzMtOcizOgQ2tldautsf0judI
tILBLfa6aZwo/kdx7Q51MKD9PXYnpatPiwzqkmvyL00YICBa/w5ARifH5c5eiI7EVgGZMo8w/CIz
V30VZOz6iKUTqkoz4AWMzItCNwxtcPRx7JNgJ2hNCzyNKsZ09xB14+veGHyUtrIq7UvXWzacz7zI
Nu8hmds0aOhgWpPmYgM0ybfxfClxEYXlt9LsxqvUt8F16xDzDA5RQVidNieK1ZE0upYbokM5AxEH
ohc7tksKeaCnPsVVnCs80WaqVh7ah8GzY9MPVG89NP4Pl85DB8QHsIQ7dLfGntCcezYKel6OYtvR
+3M3rLbWQe8wIx/vO+KzLYmrYuSBZ8CfwSeCOpUvUhKm+bpeAOwnSosVaxUa0hizAwBtPSWJMgJU
CsJGvmfrRt8iXnA9FznAXDHQqpWwNNCGctZSEpSewygXV6TFCOKfF7CPLHagpfB5qoDDClCQ76nS
6CGW0x6gNa+t88gaIZ85M71F5e88+P6dvnmtkcDnDIqdCPheIUqXcaxmCXaNMNboUhT3u3N8ssXK
YZpGXvEk33adgrGXJHMM7gLJZ7M2qDBzTKS99/sR/8D8JwECHB5und1VubbdNBMiHlCqq6Wr7b0K
GQ7sT7N/hvEkrko8cykLS9uQGTvfzRH7TYXQ077xVyCccfKqLJSb7WxbHLhRA0vawQRBHNsEQHKo
/9w9hqgMmduBV1sm8LQw6scNdKExsZO659J75A/vdefbpfg4gB969d98ANcqQweNaGMfOB1hLgQP
EaKvmC/8CaIBuEyeryVcJm51WX05eub3X081fQSSH07nL1sCxODgC9ZESZMD34y6p7AHkeKDE7vL
ylc+/2dpYt7Kn7FVAfFnzf1/581AlKZOjrh0PEFyH+0tLhHRwEQolB9IBZel5/OXOGKJbA325uqB
G2dXvWlKkN3vKaCYOfLJcCv4A9UM7VMKXztwUqQdOp0n//YU30YmNOzpB4JZDFMpFzY1Bs2UbSSs
3AgsVNkRmaLOS8PUwzO72lMrnlyAdbJDa1a25OXTzaVMJ3byvfvJRsxjNx2qlS0vUbCo06qP5Oxg
LIj6oZvMCNY+Ma+m12WcqJkM0ZgdAB/4J3dMrHu0FaknhnbfcWRoUrzcdEhiZcA1PwsXfEg9/HZl
MVV7MbulB0T5D98e09HZ4EDFAo7MvLnenJYxRRSXt7PsOrn+teCA8ypY56NqWIm2Z3EKrNp4PO7e
c3QXISIcD/R42GI17XdQfb3o5MIiueEP6aq3toheBZn3nwaM9tBCYXR5uatR26q7PTgjjDjZyaVX
GodQae1Rfr+yXJqZU2eXaJ32c1SsIHqJZbaUw4nYmiT99ouJh6cdKEryGqw+RbUSn7D+Vn8Lb359
V3hBek903Kxg1/aB16XxNphzbpV10u/U8ss0wfhfv41NfiMB68BlqSwIzGc+0M7Xd/pMyIMx/pqS
AWS3Z95eO4onPfyjVz77jQCoC1xHHi/wJ13lXfg6YNl3eiBCuv1T7xMBP7iGJKXVT+75HMWQDVQ1
TCSy0/xHt4LzGQMj3as7o0ZxG7nGQhElAimFo8fV4zPi/1vNR8GUBP+rEJJXAN3HzQ43HLu2P+1h
W+q5+RU/fXzFyBiSkdiMrPUellKR+t/oB+sVcT3PvtToBRl5ygniwX4AiFm5eSyMBiTstJPTHh4b
zCiKQC3PLG9IkspePREvQ2XucAv+63qhB1qmLC/H5ZH6z40euOXtK+PEMA6gKk1tvJhPFrKY7RP8
OWuk5zVRPCR8n8vyASNETV48J4ENp+Iw8KoK2oyekpkUP2mm/N5H5sRom3zizu7ry/tcf3xz+cHb
uJLJvsPXPozKWepBcQ/iftCno1Uj8KnR2L9Dvr2hxw9U36yzslM3qkPgd+Ziic8vzqvUVj00tfsL
Ae/fgPrkC8hIB2+d/5TrmYSMw/Dm/aIwTakRjdYQ7IEjZY8E+nEufN62C1V3tSLpIpJYqxdWVqbg
hkB6p1qXvqzy67tjFADceAN83uDkk2YQMaCHPu06Aco6VNjgn4n/75U/hHkjBk6qXk1zpucQOmGx
IXnX3qiz8sQ4+oOh7L00jfA52TR73lfmIBQGJytsEMuVZuRfGo7R+/qfZAFf3pQYA+Q+oLE5R5DG
J4qy38TSwQwaXrdWOFgFvQ9bVlHq7QMhgKS/bk/GxjyQg71hRT/7W/Dg5qHuiHajuK330eGTOkae
61WspwhIB+zTd2SwPbBEgj00yiZJi7YSeJaX8t8qfezieA9cSMbgDlQlmr+oXp7G+ImclmkaGj7d
29WILW/08e+2/SHvkWK121c4qC4cmUn4/0BeKg+GyBxD2vC3nlABMVuCCslK1JxUPvP8AFuKMcFc
cP7winBM+XZwQzcN5a1NbXI1A9pgja8bOEuFFX/8Dum7rsM6LdnKsVSHWuO1z9z8lvOLmT81kFId
52lSSfNWMzPHccWOavCIoBhEpd14/M53EXFb9xzzXn8lfAXEzeK1TB16MGRlL/0CZtfhY5Bpi/+1
NynccGdb4XajtwNGFCTEJ91Ba2Z2piY1CDp0f1v2AeAxyyPJSd53GrUWEhoN+HR7FgDtOpvu9xMb
hH7x7bHBCrFUAyfQLwoPjAPaIMRRU7niFloor4/qaEArMbqLWoTCKmAgWgPlANZu3yFzswDvbjCv
zfip9I0neY6dP/SPrxRhOwj1r+qqlT1KknVF6ppUhZE6we/m+ENdJbr6RNI0Kca4qHAGFGo+UVQ5
KkqKEa6mJp64uqnCCrOuMZJ1eKDO48MUiSXx5a8ignfAy4mrpf9BFacqnHAZeoedevq7Kam+l6fA
TqnTLuGWsWqsnXd0zq+1mGPf8OR6XoCzpRi+o1iZEvcH1e0NKV30gCbvitVU2xe3irGUol4WLws7
Q9FFhjyR77eIgX+Z8GLabbR3gIkYi5ejR5zQV35ajvwgNyeFOwQCjpVBjcm9P/NTRcvj8jRV9d68
mDWoN0iEPF4bSSImiBCgeGptevq5k/ugg6mfSZTfxjLhct3OiY8EgjTMPAi2k6ONfZ8+0gixo4wC
S+ha6ycN+cgccK4qobRQwoNiqnvC8QFA5XTvwlYOSoAjllAF1y57uaUpbCx7IzE8ZIGkcsKWz6e4
M7u5KlwSXnoO2s35DfvhFros6t7+j2Qa8SmCp9HCsx0OQIG2Z+soVbtwveeYYnnmvBv+ExxI2B3p
GQ6TyLrktyl7V0+94m14nhKnnHXuUyFCAS1FIc8XeuSThELio8Gc60VpJCY4RzqwqDjCl7Jg7jPN
Sa8/HpWMfgdVl0TSR4+JqlXxg7mYyxoJsExAsS93YzkZTEZMlOzyRygSLHNxdko2Gphv9HO8UTF3
d7PNsHhFyDlJQIMkBAMWzQoAW470oG9eQl/OfcNNew0s4s+0YP1HbyXUHLHmzrmlHgwN7zVuBYlO
G2txlzm55bTRobKdUc2dwBVfF88dFjFBWJmPkpnxm17kR/tcNcMD9HPx85pu59LZomfKSaXUYsqp
Jnwd6Cd9cLg8oCoX6x6Iy4xSaMmxannUst13kf+YeGQtwzUz5bM6rlW3Bi8xmVHFpIX65o8insy4
8P0YAPVEB9JmsbxNYDdnPeRQBMu0z3YY1S1wNnxNfOMhAgd2NbQwfPWTSmuX9THnsNKgQPP0JAwZ
hTECsG23fpIj3v0CubznRk0r0AsUYLiN3xh6edIv8xTgHCAQyPGgJikNYMHT4o/mRVBg3EWLY1RP
0gBNZ48/cN2NQTUoIPA3uIS4X3PUhqB+4Ic0iDNrEFN/0kK3xhmfUbE4CTKFzjb79g+fXTMK52QZ
J/1hLzvmaTODfP+o/5gFL9VRCtyo3eQLeiaLxZ4miebUJ6I82JRUZfIp8Ng5r4oOnGfvhwnohXCP
3ha6aeUtbHePaDS4Ews3f+iiLX8DA4a+zwoMWqN3ot6QlKTxsxsQBNA0vy9dGOiyzYkIY53dVHLk
/fRzaF+4mAgmpXQJd0wmHxKqI+C+iicU0UNHKsgD0saNKnMdZnbXrobKpeuUqQdlKRUYpn8PbVRy
XjJjMuPrUkAPFwYD1T2R/X8w8khhBSna1yEEUN9AAkKaRQP1OM4sJOZMpgCdoS7kjOlEdeqq1WQq
LIc/cyqTcbda0YvFUg2WJoC/hDCRzkdvw8BG8lQwI43xtO75iq2iygCV05yFUmhzoUuY6hjSdwOG
1FagVM7F6USIArxwOk1LhUJ0fC1UtSHHtQXqXtjiU+5B6za/bO+Yl7jMdnhbBgLxDPXzCyTi5jW7
S1+Mqs7E16JuryH4OSBd8tzJlaXfzDihgyUxe3JugnIcgrTdWWEJ8/qFhSAhX5A83MsQ/l0IAdrt
T6hUyVkL9NFWr/DBGDTqUnEbFGd7dRoyehDjPa97l6Rx2HQDq/kPg2RdADBFXp4wcgRe2K9x2DzE
PaicUXibs7tQoNzRniEFaZFTGbQcAXpHMEW5Y4KcymneosH5FKsllbU44OAZSt/2VbjMJd01hJcj
T6M/WichSnJS+6nE2P+IhJxdS0l1zHF+ORRe3PNO6iZaPPV1Dca5GUZ4l1VTFa3AAggoF5fmYARm
bTEV8J4knXhCZk0nv1XWgw7GYzrAphYTm1VQZCuC+lhkt3XRVJcBu0sDDPx8iYUkLwVa2i0OY2OT
a5twp1U9Mb7ewEwqocoxlIETlDEHgHuNBYAPGkYgHXQ6q6GP3Tgz7IT6mdedY6jUvXjaYyWULjdg
LdkB4Au6RdCDTRc/Txmgv3SUBoYkQAOhz0sveP2GhlP8/U3PNn7Cp58ALwvCDcKl+hMQyU7huwtb
ylZa96S5YBCY7sEngryXz3/XHnNGIOYEKf4LKtvOj8/NKxKl7koT1qlXLtP1qxWfxpd6VoABkAGQ
GUI7a6xbcuKfr6fkn0ewPSLL3ZdPUrZkaDG/m/xpZhAAyNEYuTfU06SeqvPtqbatw7Z09Hcw2fU+
OYpqTqyGZ8XR2p88TLdEd1yqF9iQF8ht1k1qBQjNl7c7X9ulWUY3orjVmErnK44Cmu9Tsu7lGh6z
4mG5wWC5jHh3V8W4fCKN+W4bX5XT83Exme7sft7OBFI1HzpSPteoxNCKu2J8KzgGfaJH1lXfrDQG
SxEii0x8UNedOUbYk390en1P40QKahhj6a7v+jAp8s8uuJi+Wd4YJmS7+MHQXdkGFq/NHW4hIeH5
FZ7UcX07yleCSo+ZMWHgvwOsGNu14CwhjHs1k5oKN1uQNa/S2L9pdkag8WvKejU1V/hIIIn6wW56
JmQnEN6uC3jR9QMLmMkqhd8JM07oGKqv0JATlbAgsmnaL1L8Bzz3o0fNFB3Cj4NgJ2jzvZLmJNVX
1d9dseTjJFOVeTFxVKUURZyktts4oQ3G7L/rhK7A1CDXjBvJr/aHVwOe2dA58fPQ3Y6qK3FI75qb
ojGmVYddFScgWdm3X5qdDPLIguYdt5triACa9QyD71GlklKR7hn1MnYrbTkfvW8OS7h6Xpa1Iidx
8uFxuvwQrdXJE+YMj/AggWgom7lmDt9O0RnnEAteptP9bYSmpVQmrXNahmb2wgVUNgduJ04gI/75
ToPD77Q2EtuuXmLiYM5U7AETmg8wXunsdRSUUjPZu0sVvlN8O1e/8hkcR/7jkpJNN+theoIp1Wpa
Jc8YuhPxHD91ZONLI9ypBUdJ2sb68bh8nHg1RF5sqZJwBgoYjEwTgk+8I+Hv214M0IEkXzX5jV9N
FuORb1OSpct+A6W8TW/J9OPiYiskmlr++QePTJomXG2Y5d0pV8QnXN7J7dSEeLiSQVwNXvfdy9aB
9OE64RxDskzpjkP2YTP80BQ01Vp81d/ewfNZdu9onaSamqlXaPhxmeVy2gO+qXEdPf0/S1dCnWLE
NHOTQBIXg/V0rwMsxvucBH+JJhE40U1FEfrewCZKc2FpM2fJI7gRsBU4HDuya1msSNCmZDfwkd/h
UIvfbhv/rMfBE5tluDGuabZ4CsQshtvoe7W5D/XhtkTkKFl4eYM0LUykb0ftPQ5IPNEO63MTYR4M
6IBaHnhbDcFIMOGKlXGJ6ez8DxcQ6gdvT7fYt45AYl6veB92urmcVI47WjNh+kEkoOYLLOorAOyF
WLzBzScP7t75kuK8myBlRf5Ua0XwmQsipTAXRZMCwYjmvvLkqlqC+QJF4XPocYvurQ4jffN/ADGG
VLUjDIsk06TZgRp4PAwAVgBWjAyMNgaHtQiiQTWzhYwLSmw/k6ja5SRGD4cpK/g2FiEbJ/xirx5J
8lokkA1FIdDUPJ986HIcfkDEWY/BqmmYLMMY4SsCBJTmKt0amN2VtccIIz8UQHqvAIV6uQU6IuXJ
z8e2lDnCKTN+824g173Gca32iyFfQxkP//KOWqJLw/q9he4R730Llr+hpeXYLNeY48K1LZ2uLpBl
6SDR6tx9DFdxx56r8W86en4dlxUg870raJsp76VPEzp8Dls1FLRA9RhChPLquyywos0IYrAFTXb8
DlPQubp9PvSFChWU4RHSHm7YTpkWUKojHkEz6B13QbQMgE2ygsw+v988aWf1/6k3AW2MukVxlUcN
Y4fLrqL1mIGKD9DtfrMKaFd7dH25VKP44nN3NUbbz2mbV8IRrp0GJHz5z1NUiM6sED+p5ZAIKq8v
+cSw0Tt/w3U8Qc2K7HXkaLSfOq1mQNJhXFxtR5Kx7a31+fdUpihhUEJc9CxHjkkl2c9L4pmlPbcU
beUtu1lpgc+Rogcw1MTxqrk/XbfYiL6VRLwtXEiqjwQ+L089fb/mROgj8g+YtQrLVsFydy97970C
Uzvp2jRGn9QsBNWuZZLN4+ZRPH+c16FmrsgNQnt+VkTux2NllcBomTpYNbEPkjwEq5kEXb0bnX6g
fou0ELxnZK/lP/4NN2XS7d6jZLFmj/wmHdyRqFMmmvYiJrt5AVicQ3lWTy37AlMOYw7t1dME3BGL
z5vWQ3Ze9ln9k+HjIWgLySZY07uDvFU1cokxr5yW5x7G26mtAgG7PLBxnFFpnmUb1BJK0csNBXBf
cHYqLg5KkkNyDNSpss3Mwu8gw1FA4zChY4rNXtgcXaC8tyo1M3P/qO1A1k6L3XGwDVltgbdJxD3X
DWcK9jxlJNL8Nj5rGe8WbD3QvItn5r92vrhRBISywIY3f1Z9WFJpAge3v8P1er8VueBSmuRzbsVK
0yrH50NnP/q5VrOM2OEPZrHyiZDorMgeWDf5ZSXsu75ooAeosCrIEElbgMVWbccrF4hZjOcbRttn
mcH/+AdzqOdyIqqZ8/bNCjP/riJqwE1srDxcfQwQVNMi9C0J6kex63mgI1QR40VJUO0cEPHcMSBz
ueS6m5ApOx1lfPUsJ9Q7ocaP42vzN1fNgI2XA0zoCh45b6PCSRk5qILobXj7o1cSCBAJ0XypkVxk
1DzV4Ed/X+4a230YM+q3A9WpjoADP4Ruh6YvEEnFbWbcFtd/D1iXf+7nHoCBn3D0XuMXRPy7Va8M
4BFbJJLzE4b+eF567yedlw/q3ahb7e2zXxCfkmh7OQzR8hAWm3zyBwu+clqjOAl/r4UlMWCzhvzc
OOaJX2W2c8UzxIcklyMuRnp4H5LpOE9YFpxG06FSIQtn7SewhR5Ljg+kGPyza5NAdQcpO8Ese9Zj
NbgEseNA6cZhO8mEI2kMeorNtRVV4asZffb4d6pWBPA0mROrKTFZVEMaX+N2+wI323CkqC/KAu76
S3dXNfVAGn50A1xmMJ3mFVvTCaXEaua+UfzTdaUoa6lv+J7z8H3NDoH333paJRPLdD0fwkW7YvNT
GyVeJA66L2Ux0yimjZexsyhC4vkm5JttmGWNKdsF3n/whHyOV0FEv6BsCEQ6dwjIShTOxpcIqQaa
/pLCAAWJB2YK9OA06lMo/auZfaD10X9UOFUJf/2ClXOM7GBoWA9N75zfY6LY0p5bCgVqNhZlVaNF
dXOjDDYKvzJ5PePSGu8iW8/lLOhuDrkfsahf9avYpKbwaeU+WZCSgCUV4NlfqxXkG4qIGtcM8GU7
TplrVeiMEZQHjrPBA1gCBMpxlZoxHAXle2+9PPy6p20eIGoRaGK++qlB2uqOp5LZBWN/8uChITGO
NhmK0RlDjwHhPVvUtnVSHny/7O0OnfiNM7OhSA6uldBZXhN7+SOG3aZyDFczYLGFxfP4a9yBvoYU
pfItJ/H6/BIWDsqvPeXWRWX0kMGzdBHXPcUa22w+6GJmBGSEVUgmdlUQluFfPayE+Ld/614NE/XN
3jJiYhoKpTqeyqZCD4n/r5Iq4b5nXo+O8TSQ42tCNkZMsQjOUqMXl1UBFkeVKj3RQXlh/goqVAI9
Lej2Tr8iuBKK7sZtXOJj6R8Pdt9hjwkmYYJ9klDIooa+CP9HFC31ox4qYEOEdSlVlFMgIQb/VCoz
aPZi2xcx1zMdtHxsBKV2G7OTuL0/bp91mSrD8x44umy9YsiQKHpOXxOzCvQkAhJusrlWhWXLwlw7
V8tjtwIoUbnGwfQx48vPRUxTs2SDpDtXfcJwca2Nj9sOLYwBjq3j2TQ51oApwtIk8i1I3HVbXkO4
uJPzRVrQhTJnvGUELHfV/Mk9qAFAot2f561FvyNTfSY9FSzYqi/+SdT9CzQjjOCjPIO8vyKZVill
kvWOFVd8j+Pc6qu3vcQBHIEzJJI2lcygM3RbAl6S8LZZVL20dl81mT+NOOyc/U9vAGRdekGaEFdc
2aCox7T/b7VGGhmpxISfNDyDc+ieKUx2v3m3V97iujXtYOYqF+c2We2wZaCGEtLEPWikBAg4t5Pu
+BUIAUMldd33R2tI0uzEyoX/qn4Iz533VhDM7FMIAxuwOnLtq2JfvXfrq2YBEVPsprjip4l/+67X
H5MyHLcAitCZu1+n+CECF4rlmCIXv4Ng4tYlIGGtN+yWEj5zYKIqrnc20vA6YpSCTowifxKgrr3H
Y85zcyzpGHYVZnFy1Rq0kl1k9l3ETdPjWhHc38dxC6k5jZvA+7IZLzVj53mrsFskvdrVpy79e1h5
NWwM9HgC/dmnwa0aW+VuXtae7TK+D6sx++MBhaWzNfirGjaeqx5V+xNtOhs+Um9dnNOP5ndgoOom
OEK3Rexg5bHd4JcCwrAptImhajrGRse7/cLrRpMIPojbOVKP5WdkY26CkMr6a0s4wD98vptX31pW
dde8uj5UDI74KCHzG6fUsvacqb0ej7Hc8skL6I9mGWo6U/GJagmrILrfg1osMNBFQODCbU2aLlIC
f7QnKJ1GNAfjczA9IfISgCMJ91AhULvek0IjKfQh727Hr3fC7wytXwoCjL++fkNC1272J2YyMIvh
cTIobSqVF9OsR8fBzNXXgXnIR2NkW/QNuMHLXvXD/1YejSD1BhPtBmZ16hwF2+hm1FBcmrxn9MVU
2qAiFRsZGQ1lNSV/RM/6znBjSQsRyiafxavpu75v+mh8aFHVlZHojblIXbdaAUWdtQGijzNgcPKY
1kks5/LNMi9F5/P9G17wnsPj41RB1IA8VmDx/U3nWKn3nWXieUkPpjNVRrGNTTsUNrW/CrltYKvr
QfEDY0MuEm+rf/tC5NhkCHSyDWKEeJPBY21i3w0aQYkgO7Q2+DnS5sEQJlNrZIGdtVHX08OSe4RK
KFx6SggiG7FgnqrjbztwbzpEL84Jj5RsXDrj5YZQFpkgtP0puY+70aIlEGA8aI5lTtsnJUf9aSAN
FmtsqKTV748a3IcK+DKaFWvu8VSp3PQWQP/NmPqyfKe6kskPpYCo3upw9XMTlFtl1DLQd0ZqpmvA
Re9/6cCgnPulKOsOXKD2tr94GDD7FK61h8Y8dbHul1VbXUp6qwuMVBvubhzSK8+31uixmlg4BnZh
GSC9tfExk+4rPXDBY9oyjbdZjaSY0JLiv/ZONj69SKeZiEpm8t32u4bRxQysh/yrw6ktWF2joGJa
U9ph8jy19CxW409LVnoZNR9iDKhQYkhbXeaxi3BMXSNS86FKjSPrWE8wt1FXU1iIp0cCtxIHs/DS
UZNTuPY2y784nVSFdI3/wxM8jUhyJP8Z1weqIN+6vdPkU+1M3+HUDyiz7PnamrQkpN8arp9QSuIp
794NfhdEm4IxNOB8iG/H2Fkh3BkaJA1+k0IuuGz/n1ImWt0jbWxGZLZm3koH067W1gqUibX+1S2w
ghlZmsGXN0t/WfEQJFklnTcqH+bMA30vAg9DmD8iq7X5zGGZ5v3CCjUdr/58uJVEjYryzvBeUv99
565vClV8nCgkqnN4llsujqfgDB8prgb/vPnrdf8uqWRqMi81B3VTXDEb7oz8V47u5fjoqjcBQJgR
1TF/iRDIXgNdgsdnGMZagnq8vsEv0Bd8p+taQkVEQPC7x78Ueg5c+ad1aAIhZ4QuslYLdEdLhFYh
PWcTY+LGJgc/BkGY7b3vyxc0lafLaLSiyKmW6KfId6MPEXo+Lhkj5HMma6ZKAT0g/gGG98XhtpEG
iaLtuMITiXKkFgDJ9CmuqyEF1lz2ElmhExFUEi0tCLc2m/3E+/0Kg2eUvJsJINGXxQKmS+AapmxL
PYTVLECF+O3h29zO/AjbcqEP+rKcqxYM5g62l6TtXUApSXGrWNYooz8oxKGZD7Yo3p0SbHImCLi0
QMxCTdmvp1CtqjbHxDe9Y9DDjQRUH9czXj/0JNmdgBoYcKpDaaUG7RZiq/W6x4T0ojXUbaYo4+r5
E+RHt3WzdDkUHXvm7yzc7ITutDsz71LYbZfFNhbW7edVrzUhV5QV4UDBA2pq7qym3L2ddhbZtM5F
iqzkgWwt09gMV+4vpkavn1ffBFnlyO5akBCfGQBO6taFspi63J9dARQdm0ZX56qHWx+3ib4GpswA
+M55dIQBL5lCW5Z4PNzbWrv4LWMswCvlUzD5IH1VyVobGFAreN4aHuGtOhPAH34khxKsq24mxVmt
0NP3bFu4voC8eMQWrASpXHM6cg8jTkNwOpw/OQvc9MpeeVtWikbB9wAGNIUH/V4GpP6nSd0FSbH7
AKz6Vir+2PNOyc2VExuAd+WKUp5Sp7+LFewIpCzNSdXqqfYtFnyZ7cjJf9qpDuweNO2k+mQkp4Fg
4Vu43zZBXwo9YH5+DzXVrkicJBaVEmFSl8JRDT/E4eGHNiBfaWSojwDqYr5eiqe6oYsQttGcn6k3
5q7V21PKMMGZw5w9A9PZnC6NtFEuGKjAFpbQQVy4ph9F6kXkInCv808XPXhKFymOLIiiBZcSWcLc
dEwaRHXLY/Mgj94yCvW9foZd0oGcdGdM5J+/gJ691rhzVr7KwQhIfPQP2TwoJf/iZN3OvsRY9hYN
FioaJvDchBH2L5y5+R/W2tZzOXa56jZuMONzu+Rbwurkuo7tbvaRGC6MHRUQfMNa8dLfMofvpL/7
2LgTGdJ8ni8tqXPIYNK4M0GRbDCiVD91pofzSQmXQW8/uLlmh4efgURIBlnlsB7T5iAyLR7W4Ei2
x7E2XSvA0qpwRHjtQJLmySAV/N2T2HE2HbTMtm48cJxVeGq1Fj9cwsg/Qd1Dn41FsK8JY6UbIQ0c
70fTQDEBzXxGwytua+2xUCetO8EnbBSlHLOOI+CasShWX1ZB9gB1wHkIM+Yp/dzCMKlpWtj0KnB9
pVm6r6xmjYVK2CSS3vh9TU5vMXfHOcib6p3M/dKbiyxUqgiiJ9jcqYGII2hrJd3n+oezghKl2vGo
vtbBAbb0iIo4zEiYSfqELGx81amih0+4Bm3dvS8TJ7SGsFsOhB0uXzepub1O0Vvt9pmkkE0JdvmH
L6zfDTFjlcIKUIV6DTk08Gzxtq9yd4xmnV1ORBFglt2MxUET/Qh8hNpge49NqGBJDPxrAkMhV/0l
qvsNS6CqdxDiafaL03ct3cVRmBp5TRoBXDI5LoyPyo+f4NkNKKjuAaJenMdwfqCeJ1/ZwX1RHO0w
Um+CbSCUIAuKfJEady29Gv+hOj+nFTNYguYQyq8zjfXOjSNT4bYjzuXpkKyXGHGG1/xeUk0mfc/q
KPasuW9f0n/5Vt2Cn/9yINc2+CaODQTeZF5g350BS+mEGNacD/CQCa6hsQXoczRKtYT9ZHFiXe9d
XQOmsccdxLlRn78GutBmCjIjoCpa8DJCo06VY79FPFR6zaVgw/h99oISYX0TgqjEBiDz8Rh+kEf/
xzzhGNjA/N0GPC2qhorFAzQNCn1OLuHKzqo04NCn2Yi2vDOv4p3FX1ErOcLpSZGG7VMzmSgwzYZw
gQDkc0BYOydl5gf5errjV+upHfwedZvnrmkYNsGX+UkZAkDeQIf5waLDTzSAA0gE7sfE50/F3dS+
SwWc76Mvi502YMe3GupsOjW+9L8tJRLBrsCaPyuQd/SLUQ4T80n7+NUY2h0KpX+wTxRVh1Y5r8dX
BpwBMTw6vYfJLd+08c6GzpHiIlRipn64HuT2WLw3BwM1qu3QsbKWatuAvkwF5C5RMt8U6gV5d3FV
tTxQSTmxEssmsbyS4UWZTtxWi5DDQdFA1MVWyqY7kuMO22jzUs+7yGUoKSeq0Wva4T8SiZwQxzR3
PgAlU5GGvtDf3CdpIWQ0S0vmjL6pG1vYhSzBEf68Z5IMR7gu6qcNVNt8i1ayYDQJ6BzCJ36eTEsh
1M6iPklHBsCzIyaGzj3Var616oaTAi6Ug8mihtxm1nNEJ5HWZowpxdxi/+o9vQwGUIae4QF4aoeA
UoXxeoSYUC0d+bF8/Sk0jDQMzWG55n75fTo4Hgr3jowyOi9LQEyAnTY/KAlgkqWY3VfJ8oS5ZdlC
VoAur5M0lliOCvsH4Ejzm6YMUtju2edjWbnaumqt7+pvnekE+hEos4VbBhCECn0AyFXVcluDEjeW
oGo3AxBzcJe5YNIh+pN/7+gOiYLjIMWPYt/9gmK0R8g0xqt+uaKT7cSdqSTChRecXnNf48ETC9qJ
pWo401qZMoXYpzXwlAb+aEVez25qbFiuWkaNvyqnTD/iqubKFXvNHOiDdSJHuHbwOV54edaXtkyd
R501EuhT2vXQ+jeBLujYvvlj2DEQHWe+WTfIVJ/TQfOZUgjNA1LJyyn2GW6OEDj7JU+E+U96bAVM
zVPvkywzssdPPlt1imrgrKIFwAqnu0lQRcZAEnIHAV6KLXRwAte25z9G7HU2LbOrpsgY6Xlri4se
wnvdA9KQVFfWBVVF/rmHVqMnHbD0NYT70p638CdHh8BD2o/sc+YiPW3Dym5eZXP9u9NMb18K5NAi
pjzjbFmoTyGMfuKBWNy0fWdLzdDcLlmSKkB4jba7DGBo4uFBe2upp/eo7BIuuNBBO7Y+6waoew4r
ERlgB432VJyppiq8ofk2XHKU0RTjgGme9JEwt9voArislmuH6+zQwpAiTlrLcQPcBMJmvbpxyDtW
UpIWdhTOtKl//9PdMgulrZQiDnfkL1p7qfwp4aMPUtOGJqzRsRct5DzajKIiX8u6FtcxdgbQ/Lq8
l7u7PYQej3ESfTCpfETteWYRhrJaYMdgnW/G9HT/O4C95bUriL/yZZJY58g2SRBZAVH7KLAmJz4V
Rq24ZiFnVQx5RO2MdmxBYqHavk+TJJPNpfoDqEDZUPCIgrwF5mXb6Jfa99l1yVjOTaGQ0tNvjeiA
FHs6O9U0lTIr88se73SIrZlXQlZISDtkHYIwTaQEN2FfqWnmqLS1hO1qijrvsqjt+zYn544Xf3iD
E5fh5q7e0mfgKjU5zwi80N5tORd5loGhIjhq+PRKT5l6HAN3xVmXVdwfR+IUKFM4cK4Pm8o+EqmI
JfN/bIGwVBCkGuX3JDoaE4nfb2ROoIMyBfs+98UgHBeycKI2fwA79mx5bxH0FKatWjM9LlCWFjuq
khISbmCK1/vA4UFURRDUM8D3XBqLil8R2YUXS07sWS9xFOP1ZXNBmUBQWcjDaUMUwqN0WQqaNJWW
gNMUAHlEaqr+tBEW5gQOp1cjZtPTkREiNnThSqZe/eVZQCz7osaH0ITce8K039AuSGUolBd8u33J
t80BRbT454Y3Foduo5+wifoUz1Cde/jOWGQ/3oNcRS0KhZahJ1Q3gYLTpDJTZc/hG/pcdIbMOZgf
AyOTLU8q0cP2fvF27wfTCligei7agCkSJF42R5fr8nu0lKO1c8BEWYBCUFmpbS4GseRvzOeNRVsG
HCGwT2lmdONLw3BeNGPHoImno652sYAwDvyycar9pYEZ22L5//BqDGCoLhQoRQRnBxfl4/+oH/Qk
QqOyguIw7Z+uq/NwQCxgRUmja1Nip1k8QjvrHnbhtWigoHjhQ0n3p9qoD/UqLujVuE0wE7Rdkkdl
hz0gfBwN9ujIxQYKTz0E5JThm2q6FdNNDEu0LiEhl33307mqJTm8TNtc18QIe7R6K99Gke3aBFxf
ce210CgheOhN4YwDkYQgb4h0C/+2J5/J7IzHtRUBPA9orfTKbIbLWVePLr1m7x9zz1s8KYzB4jdq
zfRUH3JOhnDYqxwSImPb0etoMreNGWVIX+JzkPTaVWdnassOVzInvJUZNxCkeraTx1G/I/su3sL0
HtHXUMw67U3ZWqx/O7333zvqDt8Wsw6zp4MboGjatVq9Lv+BSWSg+UcjFejfXGS1TccH+mBUeTBn
Kl7huKtyivfCtrhXnGbQ1Agh9YdGjlPaUP7OadbitsW/TnClDjRkSHZcFB1KsUmRmuaCGo8QPu7c
ebwx6wtrsS+basz2mG4XabL/xJuc2Pm+Vzus9/JGHYYFgraMztzcA8Ll8M1RbbEJEXxNyEt/8NtQ
MJPcBYcIsxXIIoqLEs7QAytGkvqJ9St3Puz1nk8Yp6ehvUq1R7k6IynMELHlaZ8kKXn/FEzD1w4J
0G9lfcsDKmDeDqWAw0YmH4WpVDIVA5KAa6NkA4P1xDbq1pXMABJmrdzfn+0mRDpGccodHUgoiXdt
eqnDI2qxmqiX0icxaEckBRobhsramxxK+4m9aZbjtPzh1I3+5rZCKIbp+tgfJltV+tJsAllY5JoU
HOkp92kf788UQp6JSqL3xqOuXdnHuBSwCmJiptVTt5dDDr4zaRaj9xsg0juu9/0sXrrvEOqvCkwV
kCoK846rKIElIbk3Ke4AAyRIlUY7WluwwVrgWNcPY+6jjXgylyRmvIFrEsGHTzPXab2aocKUGv9A
xS1qAe51/80GCjGE8OfJshFJzX/nln4CDn1GuHt2uuvc4Nz2vaiJscqV9npHGB3YJfpCTIDg50BN
sPLniWLM+MlQAobR+eakma+Ra0MEyy4450WCNin7sbCKXpZSkDTsG5s/bdnu3YlYZJPtnFBSgYey
l21XgN7+nCw6c53W3D+uyCgd53d6tp3OmjrHeW/USe0F3n0lJJPY3+PqAHHi2/5OQkKvfK40I/vx
ypHtr/lylKUw3A3/Uz3SGGSIG4ZDZbyXKMg6oESQYlI27yoV5QbL3+Q5Ug2ZNPOVQP5PsO8jII/J
Nsabmv3pORLjyj77T1met8NsRgViYObs/M6Nbil/Sj9/JEWvDDjlMlXtq8XwHP5ZkWb0yPhCOYm6
D3IkaBqbOJH433ux6xta76vonAf0WW7n4oLDTDIsCASn+X5z8yOfkvLd34RIoKRvShoiWkL1YQOb
Go1HsjseUp6V79oVUqPcLkhPIJOqUDcjQdBWxtSebgK+S/7VwW3qwcpb2sE30d3h3lWIRXp3PhZE
K7YxnM0WbS144UEFMWriCu5rinsHxbe1BwtteMPN+x+rszp9SPbckHxYeC4CccHuUpciv5R23KoN
1NKovYpGCYOVB+ZYP7++bkhZW/xgxbFYAEkOIZ1zgj85Z+ovSDz22tpYH0tCms/zQL27QKWCUsZY
xdAHw1C2g+nYLWbS/ynQbK1IKyFDZl3kNJRtFME3QQtOkNasOwkD3Bk1ZYtBUYnn5qiilu6EtMap
xStgq2Vei2oSime8VDn5dqySfqIl9q5YgM2xIRSXCN1pGg8Qr6E3cJ7ZI4EHiTJ4hehB5dfqi6xw
9ENAkvGfHwobdZO9LlHi+rLEk0ot0D8wlLIAT9uoeCKghhPN0E+giumCEZcVfmCVKliAghHdOMCU
phc9OY/kOxzWyeFhUTwj6ULhtGUY7yAO5qQfIXkOpIIwEQg+U+/HhN/yFTeHH2PuY9ONTAoTWY3J
JZQwHr0n+i+o6kVCKV4Ff9AdnC65kNILUblayB7FNvm6s04RY1GEk1g7Zr5Sgp5oU7JDwQHOI87s
22bY+efawmOxiCBfZ3gSqliHDafHnCcdd/Xo7AvFt0dpiF++0lPJoMESzmIdeR8sWYMG+hjFNy9y
22EvlIgS1d1P4d2HX6Z1UkkFqYbIwlY2fqigdWtlFHO4ARZ2tblmMO9bIGX36NjfFKkrdZc85VOw
XJNSV8FzxebDyFQextiCvLzyUP3ExhSPyCDpe+r2pEF/1N+gqRgAe3o2EwdNB6iD6uk/KonMW6aJ
+i25e46hdM4R6cbeStBNYxCrOqSrcmqlc9cXoj2a3V+d7A8Z4wCCTPDuGUuTS/ON2odlFg40NQau
MnHpcFTgTep+8ObpP5D8OD7x5ScAtQGxHbWHCaHyGER0aKlneKaIFBoGH5Vt6BiGJOK8RRNfxTKH
o7h5ioEOSEhHGYF6Eu//JvC58vf9E/4RI1vmD3IsXEgIREoMxvl3OWkth+1pMLKjR3a7Y6CdMCK6
K5RoBNYAO3aAneomgm/xp8eko0945VA3GONBRsYgn3FenZSLo03xA2VTPbbCkDIBKH0CyNjwZksw
y1z8v/ypPrb2VjK+RR00Du/i1+HJmAotfthKScfg7ENnI7bVsVNmqRwl33AZGcAe9o05WX7gURwU
hKYr1qHb+B2lxu126ObzaPh8U9MQAwhMKbpLPPOOaWmTcrwia1UT+BYwV995ytT9HFe6OqqTB/Jy
R73cKKyead+5jt/3j29+dTLzCLPFYe94RKe16H1ka04scrqpgLPwMR4Koa10mLN47EcQ7sNLgxf1
uSC2T0/xxg/O44W50UpIBcAtF1xUnrC29DzNZcTHLp8FEh/1rYtE6Q73rFaDoKKin2Wh6YsqP0ox
VhNXNd5j3CGbQb8Avz3CSzA2rk69TKQBAKGvlnY7OKa+RDciWFW9H0WMmyuzcSFkl6TyLsL+r0yw
r/6/UOwzq1p/pOP3t4E+nvMJxG/+CD7n0Gm9E/FZdjhbIHRjkI7ESx17GWPE8LaGmdP7lcBHw8B3
yNvXIm4KIJ2LBnpGpldel2zg/NXTP6c+bWptM56DKgRmAM+cvTnx54ZAu+APyeVzsbK69yk0gz1d
k/tqQvd4lnSX/DSsU5vwu0dMncEXqchbtX41ukTAgKr15e9+c7vAYJ3z3iMEu8heNyKWfBAipHZi
dDjDKWJMDWpGvCimmikY57HZCkrnITzWz8tpLJgM6b4Kh4gBbIgJRsRe1VRq+MVcLXiL3xNDEpzI
FsR7kLWxfbXSuwYPh3uzNVHRSTe1xrIFWdccUAXSkqwFSVYbqRGInAnLTbgVB3Pd0RUyuKR5ntb3
YDgweFnYksGHxfsMjMpDGZnOOEnaMPaf694jHoJmt0ji+YoUA+qZWoSuaOBQ1gJfUVsTz9VGcDAT
z2nVeYvmOEgmW3lHQEkj+lh+lTGgbP65Usf++j5mELVWPrL03eA/pDPE/5re8vCcV4Yccg2TD+k6
X455T+p9AFyJxqEYYsrfTbsOLQkJDLchmwcxxTeYWnljxs/Pcb8IxRrTkmwwRpT3XN+cA4sI6FKL
uM+cgBhzIPadlTjUJyK6dv2pNMIpN2z+0S+BinAB+7CgRT5p7pXMSIn+4e/NHQggZtiDKUwhq1PM
iybQZc6uDpYxE8BuZnYZc4YEu0O58ky772jSZLgXVkOuFPP15IrgbQkhRcDKilSev1zn91JK3gbv
yFt7Ctupd2UyMFTWY0Fp83oSTGbqP+q5sGqRC1fCsgDYmAdHCWj0sNou5mZxpDLrQRUpljcByWhq
OBpJHDHQJtu3TiTPyNeQG/G6GNsK79mLypnGZK7x2x43fJrJusi6eXtb2cnoIHbf3wSwru2gW0tN
YkVDgjFuupLqXe9fbXrsfS1A9bfZ6bQxAWZOV17+EpQtdoCq0d/zs/d/233lgjMHEW8tPQE6hrc4
4/vkIPXCfLGPTNeS5u+K+OwSIuI8zmLwrghXByHR/Tr58UVJProMGzCkocOu/2J7R1NDc12xLTyg
MFTR8YOW2US7z5tXVW9A9ZGu5iqLk8FrtWwdUQOSxoyfD7a9Ar+BsTKu/zT276juP3swRXA7gvlN
q94Hr4uuMe9gjJSa2b5HK4xjZBxZkBstzm1k8F9reZWGDixAyyWLqI9i5Ks1SOEPXjw0r6Xdwcgg
XnWErt4RKmm3JMvLJ0QBwoC2IVRL30TzgkkxM30+zB3GhJFruHVx8cHc6v5syzKxqr2fs3P1xHoS
e6GGUpOwphixfX8RDi301gjh0Jj4kYNFKHvE8PjUWkHludtbRJeLv4XQPDECHDbsWHezGrHhVVQ5
7PWSdkCGm6oYUFZXHnQTLkN/E5J+Z73FgsL/ivT/zoF2mTXlo5F2Ln3r5L0rSGfHusqUyaTYdbk9
0aYkyG2ssGhRL0YoiM5yADvk6XUfsofmIyiazcrVH53yrKjY1npL1fcN1h9bSZO1V50Z1u+KRHWb
mGRKcCTg790CzvvbznTpGSJH/NfXwtEJWtd0PIMGDGEtBiwhYRs0Oka0r3NOqoV1HIEuF7xT/dbI
qVZ3s5GmERy16YC1GbAqCpQUwcG4omlpljsYHg5KcKN1nI5QrtXYTUk3JGg75gcKloFJVez/JI2l
tqyWD1P4eIw4myKuLfve+BZRpTJT4X95FjDi15HnjMjC/5HLPdgwPq60adjI9bF0JGLTWsKC0EEE
j8qpD2oq33SmH8I4eSECW0DJihhZipcFeu2suajSlaXy3jMAitOUJLgvp7bDvSJAC1u2u5QBOYrX
a7NQBaj4Xx8l6mipyeCT+mvBBIYVqs6HsXcrojGaA7GUgyIfpcv7fBjJ/uwft/pmLFRpsPxHLk7V
MJyLdy5wh5EdtDkDOIeK5rsluM8hwTaxBKDPxJ70w80W60jAxhFr7hDYXLJfRlz8IYLTCUrLPGoZ
yzRUdcmL+N7VnclCxjttAYjNAC1C6Ww/r4H9nriOZnlY12Zumg3WB4nVAQSlzWguQ7iJhQlZVNsW
7GEnFm8KtucchRqvbni6zpSBZOKdHQZU09EF1kSGYT6Io0GeYdo2gFdW9w4Nb3+9bUJ63uIX2HUl
F6olYTEmE/PZ0bXVG0x/PR8CSj/usLu3xWB0YmqNXegKkO5IwRhqBKDA4eVoYuWG8G+eCCP+1aCY
FI1Kai4/hiY96oH0EH9hEUunNKpUsBrpnlaX73zNLKzBeLXPubT3KA9M/kTnzRKGfQh1vHyqABf7
boTtuLB8q5UC4bAH4eDXCqf8xcmwHyOPy0cuzGVh0eRB8MRBq+AypKL0/xd/A0tJIEB8YZURSeRk
KSB0sM+9vnfyu4xqnOe2nTY5mxA0EuHDWxeA+z7D4NESmvRm73mYVdMfuJ7/4uYYTNCT4e4Kk3xD
UibeY18zCY9kYqFh2SEgD18yuj/cCWzFvyiP7E7P8mF0AHrv6k1/RqFYPaUUJRPjVABdFWZnr50v
jcbHdLuKrJbTqjygLdh1Y7jsaz1EaWJmlglUMxmpmETvHNux6NrtrRVvov9TRXjNagz0aNZDdyRv
fCebrb/2QLtnCYDj68WPmPo1wGzj2xL32ung5Ipu0esQ2V0Uzd8H5VPzytQJ79UyYtD1e+AAI5dz
sQTv3LlvaTPeVIDH/UxIAsDXk4qZ596K/+wR19yvoKAsOKqZ7JO/zqjDDcvjLjNP99EYdW9Z4XMR
+iv1w4ydnpNHc273RaNZChzFtpWgZJbypY4Hey+f8EKh7n7KeuceH19phy2DvCTIhBGKXL+mRjx2
KEtMwStFNCUJzdTfO8R79cX41ZV4nJ5Iv9u+iTw8y/sd486CH5u+xlDlpFuAAxOJ9KwDiwtkwbEL
NGhYwRTI7tdQZy6XrXy34PCmb/78Q5F2v8IqBg/rwYOzUpDLUEvJ3bpb8ILUbt31Ve5EjSjeedeQ
qDovjXm0OMc47Nt7OKV3RvyI3Npd5wCyYilKprSkNyLeXqLrmy+RoL8mhHnkqNzkT9PRzRxUWPsI
4ysS6cnpgbEWkK9k23use6h+KlHKVa3hxPv+O05AzJXTegLZsl8I9Gij1WwJdq1yh6OQmATG7T7l
3r7i0c79aeaA0R6Is5sC8oTOXjgciIT2Dc8DuNargFVUMbKNIchYB4BfcivSgY/Me4qp2FpmO8w/
Ix5eai/VKQWPRDGaAixZO8Dz8C00Qpa1hsvV29r/X8mfoQ2OMxb7kp9kMgvWktMgHiVrBVpzEVY9
UHo9+LLm9m+GpPS1+USjaxwrurpoXDUkIeR58f9r1Foas6s3GiYJpsQVCel3E3cQuQEcFz9t91zB
k4qkzi5GoTGqVfCU8vDe3wp19zVMxYTyf2N6YuRj+1BNBdw7Z2m+BW33GLPOpDLPfzsrbnsBz+c3
HkE9mlPI8AM5tE6x5C1mVYb/Gp6SXhIxpuOrhhfKCTWZsYxsj87FTVs6B79axzt+LKh6ANpuUEp9
Z9E9CyKKemuuEB0nN1BmPGaMPsnbgckETC74PjURzoBN38khcZuitmil5itMXGD4Alh+bSZVSd6h
jS2QYlLmzFOj4qcf0xE83XPbG67ueRqjNe73IQh2LtkhZb9qWadrXDNUwFat1UYaMAJxrgdcO2Dt
rxBc2mxqPB/aBVqbxiUvUi64RvH/Qnzll5KNyBnafF9DoY9QuEp00tB8bCaeeSaM3/QncJzXq1/r
k+1JoAhYmih0iS3rdVhdJcu1Ttqgb3Bd4sfB++gA/Wpp59ZsF25shpmoMLC9d2Lwi7yIWcBf1Kta
bmZpR9FeWWhdfHQWJqEl+XCuW45sqEaL1m2jAPPio+z545sytz6q0gwsi/MpdAVkN9iHr3d3u9qW
I3cOb4R3arwah0Z+AJhR0jsN15FpugjdGkV/aTQKvCf0/wWFXIFA59ECPPHZwFszqxm5+sicFf7/
x+wv/K1zTCrjgI3jzgcjPUC5Iw18+g/A5V0Z+FChXUX2dFUAPqOYNZPhJba3AivdYU/lcXrrDFJ1
Wq96ycyK1EWpJilShNaWg8GmvPAX29ynoWwORkyRI878bqB1ycr2Q0KO3W5l/ol4wJCL9q6TODLW
kZRsfxVGhBtdupdsjwxpBD3zubC0jVSsn4A+os6FAHaqK34Fz911aN0SxA/f4AU2OgYRS76b5B/s
jHpm02iTWN4eQ0gRT38Jkd2UyZ/45iZX8e2EQb1WhjgC5E2H/UyqWgRMA5lzwAoDcwThoXA9G+AW
dDod3WLhjQi4CZMWRE3aDvpXS/hZ23XStAiSnUMkP6J6T/lWnTmTtE7iYxOfuP1Gons/L1/AXs0W
VaLBcaqUkfF5SQAtmU76mcl7K53Pq4uWt3ftDizW3nPC92aJtYoWI6XipvaC4V0/N6CzdxBqr9wh
PcwsQ8kMnX+VmoFlUmVJNZfsgiVQ2iNEWfcYYA7nwnCXrF6SqNunxaw7tWoPqZyMyRH8K3E+pein
5de//w3MtePblXBzV+CEaGFH5GXItQPtzYElsI9av7VGYFx4pWF1nj36sjVlDcN3c1v13fwKaI5l
R27j5lVBOuiljxRH0grNOa9bFTcKY0zK7808qRzYRrndpBQy1S2cPnzriLjCZ06hcrwl6o42jxZq
whatJJUhXQ0hJk9sg6AZXrWZW2blacicb7RrIIHwvp90ai44Imbh7wmWzdS1/GdKrlChHw9B9Mo5
QaEKdPuoppbxRCSCQz/dNVYxUW9t/BQNV2FI5uSWccV+1mb/9z7+ExppE1UEycv6bKTzSf4DfxBh
rXrTIWz33ZM3ADCCHi8oP/ZrtExjg2J7shzfiVyxWWX6xBKzLcPBhbsCLTGuWqOlO+ow3/yaFdbd
eZysftQWw8Dt1ectNsa1d6/XvsCp9pMjmylruZHvKPmhOm3L6j7+er8dHyfgljm7aUG8OKoNoHjB
odpmKxR/xBQ+JtIBammb9Ah+s9pcT+UkCH0U4XEh3ZJ8EnSPYE5/Z8+9HqOPx8csVyKk6kM9PIQ5
ay76CkrWaFkOaksso5dx3dqloXnsR54PpCzR2OASvLoYXV9Y2AVpHQjQFGZclfN+6uSODjh93+9X
Ok5L/zCSRnmsv3MifwgXYqydA5l8V5cZ86GQ2dDnaaDEEW53DbV8vYftSL0IuPms4VQ3cKggl1nH
UcS++ReXEKNUNnrR6CdBEqRv/vlhEHudCTExSKD3D0blQACchUUIbaFelQTnVkFj1ASzOS2cBdLF
LVCWQE3hOmwZmVXPtpnU9ZVJYrXuo08n5nE1TQcCJRfJkT5D33UDmkSXsVHrCXgJ95w6QzWJkvHz
jvf5GNz1wgxDZtDeljZWsWmrCxRfPiwIYWVpjxxbQID9aIkv9KPlVHILLgosP0bZkZIZZ7xdf3fT
cwHq5gM4pu21+5CZ3rvMPFauk0UR8K5MBNyIFmO9MM74tzTsGozTvMBKqu2rWouHFDbtHdcfAvYU
IA85gcq1xCI6A2wyGN8jHdbHVlh6moR8CTniyV9IwRkAQBQRyDT9DuPX8CX6YpmLNxyKk5MK3PXf
Br5tiwSQiS485DxGUU0RCwbtEyDr/QUM//9gJfsvbxsW7xoKjsZ6q+fPl6ecNMMlOU7ywPsJ0YNN
wvkImP5KCQvul4TtnZ8+Kj71hhxIqvsfmasvAy7cANgbA4PkXdKBuvQGjaDqW9ajraOxyU7nrp2U
fUKuub8jI2XRRrpZe5xmPTfuf+ICN2t+MMf6rYhatEjOIda3hLx5Y9UMhgnXHehu9KTM+MRxcImN
eGIS8kq2fZhGctnPOlmX7XbADVy4rzodaWHKFHnEpKOqbbotXTi250skEyBd814JdKz992fqlCAD
rvBWF5c+C/RA6mew+vmDAOkzqPWAoBPhN9v6g6EN3fofomCu4FvzGtqINeVVFN9sQd3K8YhwWMES
ocQqx6R84bNEYj+EVbypLxk0HMnTmOE7JqRur43W8EyKUD2HyJtYf7k4880z58sO0FkLS1HUA8Up
KbgNNMj4fi6KhfU90/Nvi7uboUe5uZogMbGqFVw54mf/YIk/xcAXigN3uOSo1QJS3hvJbme+Kj2x
Sr+O8LuLZmGo/rTC+UmVp6ND/dDBeC0G23M9TI0/oaSTlv6G3Nf08IuH8m5ExV1+YBEo29ZHD0rG
emGDfK8HDW55bNwFhMYg1XplyrM9Xw7BwhxjvaViq0d3qpCrhxveDhRmD8nIYLiY64F50TmnqQWm
1PFfhbJN3QiZ1FNnHAPdN0mBt7FToMF4Qdea6ckeSAclqOpJZJ8MijFIxIU7mAL/7DGHXy+0kuzR
i9boXTHzC6lnICeUnLN+WEvXKoe5Har2Ja86R6wvJGt/a941HXy9daD3V/ViKAutxj8CNIzTYuP7
yKrLtrzLNXKyu+A6iMmSXMZb432hm5OnoGjDJJb8fjQ8Kr/YVXqoyAVHzAr7dXCaqVv03kVEutxn
CBEMsuIjR8rKPIqALNTGPjW08oy9bDGI6Xu9jYasXS2cgGbGLWF91blzN9LdPdgrVJmjjfwE0yjW
65kg/i/KAvmn26m3HWa9AzPhBXNGmQyCrdmnhUeh4M/C3Oswmxq9XdcAlFVP0zrcjKxyaENTSoAD
jnhJxLuWg7ZWOYMDmIUHNp/8bj7yRA+jM1r+6FtyNP8Zy/72Uqm0mEIvuoPzv7c2YYRLiQDWd+xQ
ItYmPR/Ey0Q4XlnhSplyRSiQKq4CyFPMK9D6SEZeUjsNyXKRLtTjZ5qAFjAZPMHxnhnqr0KZb/yE
QIPpnYTi3vW9YhaFITrBlXg0QqIti6xBqdIQ1AXIaDVIX6LyzCAXeFwHnG8QUOMHewV0OpW5CDrt
I8IQzeF9+vY8stQiMmdQjL7lSGOeMVjaHtEs4UJRl8wTfX8jDO2Etfo0C6y/rd86AETkDbsdJOUN
o5c89RZn95jst50q8+80iO3E49LVsQpZWmYKBx8tRBCTzn3moZf16TjSb0snSNidV6YhtAHoSUjl
jJBFGYqZ/d4qxWbBcjFQUs/4TJwM9ftsduP074o7u2Rigq/6d7rFnXsZObXFXezLceYVK2r1UBos
/CPe+J29PqrbOxHMtcfsX1FsNpqMiDjdC0NIKITrQEqlEq6IXfWmYkXPhQWIKQLCF74VGvJYstsk
jGT+fN/sFf4HkFAXBns6uew/0RF1rEgKtUT5ezobFipq7YgSmx2tBR5M4dLRc+g4OiIbk7MM/+Hq
4S/Z0LrE31xJR8TJgfd4c65+cbu/bAXQtpl+Gtlw2qD1yM8oKHlVg9sEAMACRspI1w1tCuMXAt6E
OHfv2dRORrHpiasAs6vAl25Mng7WCUb7QZgwOpH6ad8kk17OtgrlfiE1iiTovAChX7brs2xZFa/V
DxncBiC02eeyO3KTXxDiVgxaF3mCbrzrmjwaCvcx50TerR+sPHylyehEHJl/fX37lsisK7eln/2M
N8D95Uf+FhzYm+bHl01VSuwyHgmsEdzq4LuvHhkb/iOEn4vFn/SK1vButb8l1Iz/sLGc2lfuK+iu
lQ89mVI98tLDm8ESb7Fzi9mQHeSCNRYgJ7ch4i1B6R26v0wDE6I4j7sX/Ggkgokg6WaCz8NI1K11
IQcBIXYAkrmM+Luo/ydnIEfxF1DePLC5IDfSuy2BioUyTYqHefbIUIrniabDQobWoI0JKHQywqmQ
HQZhBmCYYPIDuLcUrG3ZnClmU0rqP0hfn4iXCGUTu0vElyvbr57XehKgW1JnfO1gJPJlBCH3evtD
pesEE2dHn1pDR9k6L9wxJSpjcsC9q3IlyS27U4aTWqIGhvV4K+jSR0TqtFlZLxzCSmPbyFSJytWE
a9KbM5ImgCtUaqBB1DsESfB6h6RVBHE/NmH9PjlYa6yh/wgiag2BRxJcOLo7g4Kt00g8wZO6wTgK
CiJDVQAxlwnSg9ZD59gtBD7i0frKxEM/MFVlgKz6plYw6CfNkuZ6J8EKx++s6MG5esRvxRt2PyHR
iQ7RT+7qFI+oPo0xZp6O/WsJpoBp+ILBKMujaJFCZBAKGdMNHAvRudvIpm00Duffe7ewCreEUEX6
IloTOqi3jczAwR0xw7u+5kN37pwAz83EFvfxVC5m0XcBTUnamSFrxxwbr0oQa/wBUtizIRx4hp+c
ppuNsGlUsAmaLrWdBWx9mPMOFBnD/LvtadIRBMgdC+xnoqjGEPLB1TRMo9PsD8EJHz0PNRnMKRkQ
o7xWWh6HQkjF8KfJBhah7I+ExQNTQuRl6tpihyhstECqFxf1cgwgTpc+yvGSAryY2D6+m6CfP81D
tWb3lhaG+A+PchUH5lixfaxA57u+B4czz+SHBq423LNCyHpS8xGHL1JHggXqJKZnOWSlCI6Kij3o
5RQfgwnDCvq6uUg0/uT2z9S000TLzsDHipUFTCu+PpBinSzPGO6olIR3yK/uuXnRCRfiTiQLV4Ze
He+5ZPRJunN9jIXUf+uY/NTl7w42R5/o85QrCTgsC/u2blQnhBUpl/YotJOIUqaYDl7Sg+cmRcx/
R6xeF/wCY+EcG+E/SvNZjR6H64MiJalO/j+WVdD2UWMvRc1AcDPn3D7NI/cYC8zjhJjGw3Zk+0nV
JnxUepn4S0QQuGGxm7qaq+M7bFuCz+FLq4ebANhQKVxTK8zW3izfT2Wiek6W6CGBaq2nTZBDHufB
BKbuMzfs7Kq4OZckJKkx+39CVljQqiXDvRcvdqlCRB4nXB26JpQ22COzH4QIu0FsJ5DDcLsqWtqh
4XTZfFSEePk4kX7ylEIyhHOU2FiCIvyuKCJ06FcerhSxTGVv/T/LVUdpKQ0fC0XolwQGy+fyt5ib
9aMNHBXbupKnoeYXWD/eLZ8WWUkJ5WNBFfznSXijvtvXh1wuKod00lH7yAFwKvJKwii9RuWC31Rb
vh33+JpX2uXvuXxztpys5nO9Mmpteq73hKpWHgrBDB7c2DMc4sNscCpSTI+ACv8MLCIkobpirF/l
B/xGJj/P1k1qHpV3D3A07xxXeIs6GvqivibCo6NhXI5zLZS+Du0ejYT0LzFWWMsPKK4F/WB50VP3
EuSSHkX7A3jiYHYrPibjUvjKkBO6fSD3owll5Dvt/lse3dm8LYGBDkEkzypHcrLfFY1XWpxcGdUl
YWljHrVri6QT4F6DXUBLAdXfmcUdrbXG/cxnVyBoJjlq1smwosoJ2QAwfIH5C5lOVrxFF9biZAh3
P4yNi8zZXxBWz7nVtxUYTsTvyGkJ0a8lmy1fA4WgbbRqZiSz4Fi+zRPrgk0pra6D7qFGncdz2Jey
u4n+A4YvxBwlYVujyOiPsp5XGbbxeyKVoZNVff/hpwwL6EPkz2lKwkGQpmStd+bbPEzGFUY35f73
+mp19mFsxzC9bqDkZ7fYmFHFGaR3W/dSnseCYvW4hFN1k2DucLUDCGs5cW+Q0/wGGs0G4bcK6bTu
EGagdIyTFhCt2jDTo2XsSIhi/+U7kL4QT9d6mRaZRC0FMN3YQJD9VMPUwBEn5K7WRX1W4rQwvPs5
n5Mdp13vn+ghWOsIGfjXvXi+P059itUeYteITIEFC6yc4ij8ZLokPFDjLqupkR9Xptyl9ISPV1TL
gcu7AhJ3/l8IpeCEOyoeSXQe8qBZVKJKZ+twdmwg4ZuNwY1SLvEM8OvkWjembEbKeKPvAYHSxkBO
8+tytfTLF7jPegJtpXshCTMfyk1wCAewLWmAzt9RmbxlBYpo3X1yIIzcQTRalrMRL1q7DiMPnq5q
W3PMbDE3rgqgi/KzqtaZ2s3I9jDnCYo1bygTZTmy1ibEpzv6EkY9s2de6wNSFkM+e2Ejm/TNLJKb
Au3Fl3NiHTGb7djMFC3JeJOEaBmZ3a4A5+jv5zx4ZxyefkDMRfPToWXS4358F6/GXXXemkdqjNu8
wDbQhmtI/+nzsUZGZND4zwyrVUwGmLonqLuEwR3IW4RZmBcQy5oD9sCspF+hATaUffY9qllERDpf
KDmQKfBxMGp03HErptSepwczBsGhErIdeBorQTz3n38uHHwJhGZo78zjAm9mgyxpJYfvCOWCpzXo
sA8dYIWB8m6tF185/XiOLMVPcT7bJOTTaPJ0UyVQfOryM5adAdzvFQXAfAtPzu0DO0Pr+l2geceo
lAABH7KdmxFiwR5d2UP8kMe3YwF+AgvvYXUiycPTrhSkB4FP8UocDOzcuTsO79nT141bNaDNpF35
YkrYYHELbOBWW6/gt+j2lsG2/jjo8rBExf7lgOlydbmI9U5eajF20xUyqUtvtPrv48FqVcyp2PCr
+UnmdAPyhyEJLVHDyDrGn9wvLzXxl/ijNWzlXnua6y/JLUJc7mzZcPvXpWdcSX/eVFqn9lHusToK
gHdcUkUrBfoFpI7sAg1jmkVnZvLUTODs8mWtch0bsYnmYs4rBC9Vf1g38+xRoS27+27S2UmOr7Gf
Sm5f2WtqIgL8Rk41WQjlOEJj5sMx95GxtouA+oFhJV6k74OtLtMMjR+LS8ym9/4dP6jaTAUG++Ni
+a6SFBMg7hHSBxe1YyPng0LRJFZ3Wilw0WvRM5eBSKKgSLu0tggNwSSRnC28+iqxAAMP1LI5GPvZ
opMZFgFSBFMAI8bGT+Cht6/8tMO02KweCQbAPOsLqJjT9wPnec8QKfRrYBc1g/tnY6NdEDjv9J58
uAHZnNfC6YQpgYoQK3X5+xD9QC1gIouT6654sr2nDE37bM+G3W1KRCidOTq/yWLq3MlxTjXtKIHD
Ccia6zYphXsj76zO1DlOkcgqD8esfF9LWy/941tc8zg4VT6IeS3top3RMNWAoi+QCrVD9/MnTqYW
AQi4qd3S6DF1hJVGj94iY5wPDtTH+xxYErW+iYoh32/saczpQhIqQX/8/SfWSezhsYoWVZv90+KK
6V0Bvk+ejYL1RZp+M7X+KMHq1Tmpxh8IHUUvDfXZf7zVZM8bKInB2wuATR9/hRNB0yRrGyWvVe+0
DKGVItul5hb/lBQN50TPblzYHf/OF0NpQtewl6W9kujHXaJSDyyfFmGhzWuhm+FdHnWxmnpQHlmd
0nfv34egoLY8MJ+U37WZgClyjlxQESLHOMufFsJcl3CVRRIUWHWtK5M+HQ0n++SBWFpF23xKSak2
GF4q1Vi4lRNrqtvhrKKFVezz4oqWTaK3Hv4eKVqlOuQUKCrErSJ5R9tnRpxpDGuB1b0qVIRsNqUr
Wiqljin32EzZ+oTvyd1pFwvmC0oVzHeTka83n/LXFn+JFQYRHEZEOzQDrircoaeIV+1xv6L4k61F
2rd8RPH72Sn4d9XyX6qJ26+zXdnZa5F1U+4gPoCqrzY/EBbko9Ls9KRDph9LnnW4JMHiFYIy5T+r
QowUcZtj/CN2ZjetBbWyEIpvADRy0cBTfjgY3De81nslYfe/cWgrZes9hHgu43cXdxhdCBlXUfAz
myeztUhKmSfqP8MABtSJ9KqptcWPtIOCVNoIsdF459t3hQ4WyPw/F51FN/JF6Syzo3QtCjc2sxRA
4uYKBINNgeGHQdEw0c9FMZDMG02X5WZoaMovn4vL4SARM9dJ4Lb06NYs4avow85/qH3KyHKVxphF
C3Z7N/gKojv3Qt2sCckDKoy8M6eshYkX84oAgsjoaj78ERqFGZ0P/xMJVslnyfmMQiYRA4wMV1/p
Tfnpx/kJu3Z9/QHEa0mhm4LkSBOoYmzM2Qzc+cvLEpEDovAUcJ/nYWbHoNchx9o+S3FlCO2CFgD9
KxfQZBAH3Du5X5LJyWHSXP49oNnmJbRs5LlZcaOOUR52z/DnFTEL/pn1WRxshNSflTuQWdYUaC8R
knQc1PxcGqk0enZkOmlRvRqoDFP5kN/vLmoDpC6xrm+r/lLrw/y78Mnvd/fFOtEEX9R9EeO0qPgj
6prHRZNj8uvQaZNXMw3Pe8JZ84hq1oDIEFF+tnhD8fNdUC3UmS3A3f+MDqNz+MtLD+57loBXw+E5
0YZ0U6WLqn6jhRl5gWnBpSCye8tAbpDtYtdc3kFlki/s0boBgBBxs5PjyDaZ2rasQr13P/ZexQjH
ulMDg008kdxNbBdp44p16P1kDBE54bd82P6X9vmI+4llOChT4Sh00BjwQk5QWvUfxSCbZPHkq8ia
eTYkTT+dMUx5n1wJYzHcVbUu0GR7RndFlzZ5iexkzbitb6HXdEEp2kucJRrhstUvhGJOej67epRh
cHX8cnHgDHBTYzQdzOvvU/u4M5zPRO2fqEHdyO+0GRiStAwB4a3fDlDhz6iD5yk0sRnTL/HWyNwg
ty1L604Ufb/AotFrjj94j/Sam+eOKlvD81JgrA9ALMMFKxhh+ZnIsdDPvO5qBV8d2pginYRQReRT
2+cc9zhsn201qxjLnhuqKtY1JVl1erdZztZtZLmhfvUqsoZQTIG9HFIuXmXVC1hpAEhw9CeFedtO
Owg00lRo87uh8ljtilB3+Ggks6z+B+d4MQvnOp2Nfa9NYhPjphDsn2iGEJoAJ8sHwA4IXysL2pvm
t10h5S63YdMf3DrlhoV3L+QzoxBhoUMGh9/Udwv4uL/vJTEqKWuYK06+wLTOyVqMHJuOLQTGnlWS
QigUZojhxE7arAHwRZMe5H4X3i743xJuPA2VKaERQFKpypqqEokrRRHBdCAlYEZ5zvvire3iUFzW
srcinmEBmHGI5sLcuJu0/FWVcOzgd4eyQMHTr6DpE4dclNIfukjtyge6YyaqTVFUzHo6i507cREg
D0TwS/+N5Z1q9cjZDqZ6ZPt8POjnigbRWujmV/vprtVT2W3JK9f+i2RCU017u5wL8kWnV9Ra4Y7F
mndiHZA6M3ebaDHN7YMwdrU84BEzm2xrrIe7wW7eU4DzgeI5Pea28X/3yepY8yl2AzuWCN5hE/TH
WvdhmEdvCrejghf3yhFgsqbimZ8nJDY5UmDsCXcK2qflfKMKTnF5lgpn+9xRTq7b5rKXBjdhHoxp
VWfZxpmDNjg/3wrbS21HxPfxgII4eZoCiNT0hpstKh+M/64QXWf7DdhjR/sY8GPlygbVPLzjE3c/
NKAgc0m/0YCytZTF5fAHU7M69BHDsasiji6OLZEVrDR9vmjwyVPAer2kS3cs1Q2h4yMRydMSZNYM
pfqcGt3spTChJN9Jymr4hkxfwfGowi+D8YK7jLyIcDrJS4mQL/LnOdha9h3WmKKMzJhuuJWbbUbo
+uCQOaVbNJMlYMHiZPNssiopDQt5i+b0OvpU4Dt+BpzjlNwVnKl0INsOAA/IIc7zej5xhg8GVs52
4mIqLSQIAm7XKBDoU/XMwU9jSlkTWEpSZ7CwTnbNzb+lP159KkDpx7tamqZ0kCn4kBGmnMWSDOSH
OsqkHCXVam2Jk9UDH/3UqmDOr3+Wb8Dj366qYpvpx2zDSeiEHgZoSb+CCQX2Q9szH3qWkl4DTafl
dv+Mw8g6u3joqW3Wn3MxkH9gI36gn6OnJTX2ID6ZgvHuMO3vxaiiw5ga3+Jpoq2Qy3gE47ROQkJq
FCPKgHx4kyZPKR/4fRxksH7Yaz3XgucG8mBI9VCdnVY2IHm+cddVPY8fJEXSD8+i2QrGLL9wMCKW
4K3D6t0HImFuExQ/h453l9eA2pyXkw4lcXi0Ek7XT7W7uhNqYYKHlJOlZzN1TJZHGrNooZiDY3sG
QDUSrRO3xbPCuFZDT8B9LsrAurJF+jqGWMO7/OCRTsdnaRvWKGmaWHI0GAZUYg++164CcMsI9De6
ZkfvLoeKCCGxwBoOCnoLFhF75PkXn5Ud3z6PhJAyDQuUZxiTcRGEVLGIw4EMt7Fyuwik4XnBm7ps
9iEZjQDKpZtjcf3qdG1d5In9kDHeIc1VLZv85grVDPPUxslPR9D4sC1E6TEGytPC9vbEAAq2V497
v7pLXDSQGGvm06hoGZe6pjoxUBlu6z+i/zrkFKsQatmQt3j9PyGFBC7DWyWEGmTljzBaVquOLlnI
WbrHx0o6c0bnwFRrvU/l3fiRITqyszdSQdjZMysxAhn6trUdIEA4iIUpUnkpKnDLtKuq8gKQeguQ
7BE2SpuQpZZohlyxVg/mzOreBemXgv6HgQY1FLJqvuBxTSG0QLYKGii/LJpJklBDrOoTfgjBas8J
3wtaxnHAuzzy+ct/cVTP/U7MZ9QyJbIWCXr6K+fuyxfn/4+tiy+mHpy3RVTPQTC9aRTL+/hFIPAC
GlPNM1BIFMUaJNhQ/lCLIVR8Gk1yatm7vca8F+8ji89xMOlodFkyeSUaQey7nDOzMYNkagw60WaR
t6Y/3DwEQsmCY+St7c10E2Uim6OWjsJHmOfTyM8wmiyJtSs13Nbn41G7TpFzjZZvOLSCcrt5zALB
FwB0LFvjTQQ4iOkR9/SVpYciv2/qX3369hhz+OKQs2bF1yGREx+e1yl+nuh12VLC9f3TYIC10azX
vc2vwqlwaMUtSgOJSjQTNnWVn0oauJNPFuOU74sdLfLDTTrmi3Sp+RkRHOXGMiYaRIA80M/maFd+
SnSnzWj+unB7timPlmpwlDyHXoW0dcGAhPawC6j3x6UYUi/K5FkNwjcLRLrPF4drJXfFb+fZaoLO
9z9PaulXTzrX+FjBNGokB5L8H0k7/72gDAE7DMswQ1gNPrvszaLlhJ1yBRQnB/h8V0O3E3vwNwGK
hojC1kq10QomZPKa7gQKu46IRUP6Iqpa+JENPuqsiU5BJQKo2wYSpIgI0/OjTJcpMjW7XgDZGNgy
/MxE+2YjGswtzRIspCcAlo1/Ign3+I1QKUyy7E5w0PyteeKpMrMAGz42nPojDhIFFZXMG8VtncoQ
wtMzQUdP0/f2nvg2Q3B4ZtFzgzjPWCSxv1quZecLH142rtnavapMxB9FEdWDdjjI+yA7ARR/KakW
bdVnAgNcYXb1HZKYKTxSLUE/HMZR4euJ7oB+4ZB9IJSbiidyF6FzJY3jGBx0VhW74kwMWcRd+MqM
PTj4pTybxux+pGbxuCAv421lhquQipYpdpvVRug6ZmzQFiQ99lN8RHjttP/Aq0BUdNtaD8Q7geqR
r8/6IcjsUQM5ucxoDmg56OKgTaJ7Rs9MV2DnAzSmCsEB+fu0qHkhDmprFN08Io8O/tXfXckZNEex
qMVAnkNUUJAUBepLuaNeUxBkON0t+i9/ibHxI5npAaEs1xf5UBRn7T4VCaQjLJ9aq0KiPtHzIT0t
J0pk0pAj9HdqXVhw3Jm3JaIyrFfG5MkX3250VaqlhvOHPLMioOYb7qDWfnZ1K5MYF3ALv13qjJWF
dgd6RsT8EM1MFHy1I6tMa2o/oFE2uQpaXprE01lf8zkMW4eboxkOUAQt8etV8s0HgLLwdpSjUNhA
Xllx5t/KQrxH4XAHOxWDCep/MpTt5WTaQMnLBs9vuLGGp4PgrrYxDbY7M63/7Ud7wcIhKGkWgyXR
snnTCV4iO85tEXqGhj9pxJrcPDPJFdWu9a2mR4lmrTapm0NOn2iTatfBGQxhsiv19SbnTtcyEshj
WnvrVfeiuvbKwaRSj4t4nNE2+0xZwVkcZ8xhv66H6M9K8Nlsk1VucGAxlEQRcWfPAKyLaNe84IeY
3RU+uupjJV2A7iQ8Oiq+Uj71QPlb6XtrhjZVuOpBusO8giJOHPFOoRydhfec1H7jCXsFzez6KUJE
g7MAA5BAyv+OAD7LhIfDhEt/dxn1ylmZq7sma1IYB9W8AMKkBpKKSwz3AYVtoy3HicegItH7+a0J
3oaVjdQjCJ9K1yyxgui60V/EAgcBdy/avU/WH5z+rfRrUn2elNsHCKYjqg17grSX2JkGIt6MVtSY
8mz8Cu4k4QsEvPvRXB9dGQCqJ91J6FgohmIUcWQQN4ktpTTaIxMBW84/kxf0A6MsPbCB29M1BP9H
woAacemznUN4sEdmTzXxE7iWvwpKNypB71ed34TzH5JE9y579i5f7wnZrPSTl/zQXoiJaZMK6NCP
H4iT+g5v/Hhn+Js1KrzwhT+eY2YbST1jPtAjz837PGvaEMlZD7iczp14+6R3+2SNZIOpBfjWQpWV
03yVlOfUz+NknHDtuMSxvxyKyw83lMnsxZaJE7n24x86rHFIweRz2evfpaywPCb/pdug9PQHbNpf
Be1ha5dGX5kOIZgjxyqr16QC6J9USObEd78ajRaf6dRARSCjYMgKLgNchvgC2uSBsIj0RlPf9qGO
/g5HKSGawVd2RiFMhhYA4kylzIHuKNcNmllHkvIklTIEOiucr3PNZGy2Bo+o5psijAbov/Vu8UaB
ug/s/VupCH5+8SqsmdZAeozLs1t/WDo+G6wohjBLPOvHOb2YiE/l8dAe+Xz9jXMCEXzt4xmsvGbW
LReuRwOHtyna2IInD0CK5zsRpE9Hk2EKkPhPM1pq8/AqoGnEwc2f4QMb1dI8pNohfnlsQ7gVmy//
BFlTvA/HNsx9zRb6nW/FAehUV9sPawInOiZ0qP2VoJZYI+frYYKPjmr0J963SKzf5291Ei0cL0Pf
UzAruJhU0osgSTS4HfZv1UvhDhjCVCYhWvu8YRzavWZndVByl0Dyz/7J4A1k6mFZW6PPzX4h541J
P6gRIeBigSCImU0hqPPrx7OxXx6P/HrJgzKnEtnANdyTSrMHS51HRDiStvP9ODI+ImOhoUC6ScoB
XwuAPMKrJvRoGG+be8ue2QWzCarR4CD4N5SP/niqKsAKIaxr9Uk7aSsB14xgrBUCjTRzkmwMNl4g
zvsz9KXOwk0bA22nOMfaYB+dxXpDf0+ntNAUsJrLkd46WNFagj6KetviELnjVos4/HjpGMzS6t0Z
sgQqe6WLfTnsGG8qAaRYzELi9E5Zo6jlldXYbb7F+8hY/loJWGN/R8jzcx1/UOt/LJLVd52Tx12f
bexmx0H0WAok3MQLrpFCDgjudO1OM5DvmTIHhZSHRqxt1clRys3oDHcl2rGIdzdMNDzYswhQasUd
8UhD5ubdt5VKGlnvAeghXhjBqTK+5mxRTab51YomLDWVzllr2hHBVtXJDtqjyEXuAjiI23NBr/qZ
WyaxFwVGs14j9P89QrEpisLVFjsG+uMe/TfdBRbMS1Ohu9cUbEbbhbbcsUfw9Xg2xcXJbJC23/0u
9r+L0wzZPy8PW9AYwBEL03gFF1nmmOcRCkIZPdLjom6om9DWRcTviFirXNoMLZZTyNNfQLamcG/E
mv0nIOedQ8o/kl5voD2RkbeoDhABHL6oajBj4eZT0I9r7w9R2KNcLmYSjkX8Dd/CnUMaPiIlLPF8
eyoOpgg2yw7IaDfbaN+pWdokO2c9bwimtbaQBXWd59d8Av0KuOZSCyCCwt7UBzKyx6BOcEqjkuxH
DHfPA4RilMEQD7xL/ELGz4PwMz+NWSAZ37crA8m0ezprERvrJqD0KJVpWBKnQTLD89zSnV4zflam
w40SNwE4huhxGsAhmccc3troPp/adH5bjjQdJjzofhFrN6nTYLH05f7GoZX8V3uNRPmWbB2+X2hS
HMhurzEjRjBn9w07MvcZdg4lrQF4WfxJHVTdek0obxkjey+K4tze2N8ppxBkzUClAWGtBf7VgrBM
oipOSb726XHb87ryQdS9KvY32WEJy0PMrpVzWMvAPS22ZopKu77xJ8/mPGBWQp7M9w6k0rX1l92r
RnTu7NMFMDikD6qKjBsh7P4fBpHIgQXyGeQGiX/HuiPpB2oNJlFyxwYp0cKnvWdwmEoCsZSBIoFC
t4y9Hm9JRnoF+xs2ANx20NeEG3d1CY6BwTrUAh/iSE9w6MQ+1Yn/TokLoZ9E+wK+i+5Er8I0I+U6
FrcdqjljLvqX69skqDVttOt7RBdeVG8dF/+eanWUgCwlX8Mk+cfjmNxXfaCMzKbgUN8SIVniuIk/
bTspKFU7i+etI6E9aQGQohZfYu0DY/in/rRX+GVnQpH+KRN91k9YAreHSkjzUvRNZr4zlWBfU9FN
4P9fxmOjL6+v7AMVysvidjuvU8EPkCQnAT3mfkcwGFJ9fPnAwcUHWChl8AToOUxcvrdeHVEc/5Wv
w3AGFYz4il6CRusI/Cpl7kvcqO3F6N45sO06yiD1L3w1JCdL94h/YRowcuuZA9zJKR1fJ2AIWPUR
i3ap1wJki4amTglzX/NNZWB2xFRjxSoVy2h1CRzbrXoUNg4lNXsOK0r05pWiX9NU9g30S96Jz6Mv
oDeYpeG9upb4TEWK5VMGU4t9GBCtXp8erJuaaw/GM0I0rlA+uo1+gCp30ztkxInXxVBzGcwByY4U
zUBb+K+90l0w71hL835lx+z+MnumD9L5aC63xIM4bdg2nbUZkVakfGi7m0GWtQm6ok+VA3C6AsN4
b1N/FAnM9e0hK6p+RP4FuhgdeuP1K0LcIM1tDKSB+fWohYpZeg5+08iSAWTmwPFyErp8I4Imt9L8
RRmE0Lg3rgZdvgPtxZf/YITHzlHU3t4v73RXLd5YhUTcWAf/+vUesHIUixePtceXg0AmWgIFvmMy
kJcWayEytYsZTCLH8Uu08GVp0BT0qSfEhC7h/c5giRyAB9LOlCmC25Sqewbt4IVThYJwRpdbLbiF
/iDDFG/m/jdY1PobBZZmeYPQ2C8jFhUdDE6b2AzPjP44BQefksICb+zI6cwELBly8mSN/LkGxnLf
s0GrwZImBVlYphc4pPOLaRvTgkS7RYxvcGxsGfFulrAG2bdlJ4s90zHHhKx3drIcc+XBGIPSqyyL
lW4wCmmLM14oVt79ux49xocR7qGxmoTgoBqyXaDoW42LyJnfpKlJiT74eFyDrI+EVp4SaRHThKxD
jJKbCzspQvRt1CMM+RB2qHQwIJicULCgPijJkwBHcCY8Fp8OCY2pLBfrf9TUfJMud50exMQcK3Jp
N/HC4IAIyya8LK/o486v1/GVdRx/hJm91L9GN9IqYVKNXFB+Yt2eaG52wFVqY0HpmGVssIBnfPl6
MP7ASExLIHLXhAAwrrbr7MqXg5ORZzgsVjMembVjV4W31+/d3l1jC3QObzxgdle6Gk8z/dtTxlHi
jDgTkgUOPcFZ4jF6eGV51OExbrK2D9NcbPKb8asEgKnf0rvLju4gQie5xHMfudGRcBncRb5q9saC
sXJ7a2AEeQu/VMMv7298iwK3Yp3w3cbAlOKIC/S6rZMP8wDC1F08ZoDX1025G9tZWYFV/xGEZJQS
4yCviKAO8XvxWwma6l4Bj1n/lhtJyB5jpo2o+v7crIRyLkJlTivJy7YKM7OsVRyx+A0dP/7Q8s8R
FTCqjyFen78I4S1+tuU1TVIcxklrWwYq71bWeW9lPf0ugdu4vn30MNRHFbBvjlZE8QlySUq6X8di
DWjwkkLrtcu6Mibbu5uaJ+Jw0fK0686mbzDEhYk2bN+YqzgG3YtgEiaF3nUaRn+vMds6LlYdCwEn
ND1ULp5rAQo9eiNlIYN6BgfYJcF/Q+DzidtSVqrTUB7EuARr25PNzQQhoPlyxAHVtXmhRaB6EGkd
6s6MPjuhFSSkBPK9Y1xxCs1PupkgLXN0fMUged6rxePoqX8GfxUKPCJN+ENNw+DKiuhArPMbOE1f
LsFtTMPJjdJ3wg0me1eh+MmkJUVWBrFYjUntlICeNm3rNBlBO+cwk4+4uznJyADmnB/bkT9ZPqUt
bi4edse4dNkrC3DKjs76Q/WbkigoYnWMzTbOjsKHbppkFZcWQ3L4BHQ0HgTKWqIf+uWZwxX1Af4u
qAsGcb0ywEGOmw0ph4z/OFlfVVhOmMmym7GpC3tvzJWxYu8se+FEtU4RXwrd1YQyVJLTIDzlz4iQ
CTbjkcMWlRqJT+htmnsuU8QmkMGNl+z8nwyX6AeAabXzRU6AarV0r/StiWPuyVd05mliyunUKj3R
tNOpx+jWXDzWvyUK/J0TCxgnT7byPmZMhq0JVr2m7iJKxEFKcXEXNFgqo+SpmLdXZMnyrhnQnltw
x2WoYBR9z2VI1HeIQzSEwCYcQiFyvSBEK9T9h2KIYGydR1640nf7OAQd+yCJjK25GPEYBU3Vh55f
+oTTHmY5EV7zhde5vx9TyC9/c7Ls4JPgzb2pkn7IMQvrcBCrEx1bzsqueyFZnZuGAsHLeZwniupj
gXQfbumZxOAQWoGqgrCGHHC9pb0QLp+yc2+S6pM4ZUNJ6fVSQf+slIpH2HFonUHcJCKnD5J+HisI
VnOblJE7hY5LnSswER/dFZJ3gcUTE7XqkFvlOKn0cCzjvuL2U1/cqzOBWuBUGHs7XZHa7F4QdoSR
+YMTpUSi2ij+H/dWz8FWMIFSua3Z2H712+DhPX/K1TPw/xyb4OX+PxjUY4w68DxFuyMQUXlIkTG6
Zqr7amBGd4v8gy7KedivQGSNk/3KeerVg5/P+HXC42q3MTjodsf7MarFpHoMVN8iKlozpI5TlFfU
5WkH2Lyuuo263f4ZEQ9Wj96UlXgF/6nD/bmyyAWjR9Elqt2KNY/V+s03EvlrHRWjII7WhSlrxYT+
aJrPWz+Ki1FVO3ii77/kB3tAxFdpNme8GCgyGZYOSSJBVBN9PIrFAYU4O+AKdXNPt5dD46AixA8C
tfeQJTXrVa2I0y3btiUaOAgcF3GS+Xgolc0Jkg9uWRopjlIEmCc3bxR73FfZBfEliEL9727DpanC
0wCFr0UAHdR5BhnnU4OkyLsA8AbHEnbKsuNfHPz84Vni06F4BPBOg2tHyMY7t5iE87HoPKzEtS/4
3qcK9lRpUt2eY86KfRwekT8Yw2GDpuvY7PwPJaFa3l4Yj9fI7gECg+xX1Nc4zUq3uCLDCwJEZ0Km
ihR17vEXRSTx7it0div8t41QVGBMtpU2S0xDK5rtfXXnWtJndV9Pe7tvkKUWHoCGiOEo0BOlvFDi
g5L74V7jB9m2JiNTUHkr4UWZrWNYinNA2C/E1yY5EixwO0s3jfBsp+hYF/0fif+cX2NUmnmxC48Z
QgV3T4Ho5nhSgGnACd6dzmnF8vgSwlFD2VmpiZ2WwRCtGrUwDuIRlACOZq5rY9BuS0Wnn7h08QkF
byxjpFDI/KeV+NrHuvZj9YWRyUJKWeFzd+Ok3GAYoQS2wsK6VabLY4T3OG79HTCo0F4bJD5Xkzjs
EPXfKdVA08cZGbnq97pzv/gbFTuFy1S/QgIem67SOkPk3tRSL62xDFsMadsdUBVLVlN0lVGIWxPE
d5Ha6kEMaYOLWHsgeC9fKRb+RierlvJP0vFAyWoe0KZ7uYBCIfL66DbbxsR3KeXt4aJfALuMhwWs
pJdO+b0GyuI1XatVVb4/B9c0Z6LKkYj5s8W0ymirs3ydoU3AiIfalDGLNJV8haJbTeUlUdl8y5kV
I6LJIk86twm1E3+uBxtjGrlw9M6D9qrx5/0mapyylVvVHlyH4prIDF3F6uuOprEhGEqisXL+UbAW
OE5qwAHOcAfV5le3FJbmcCCpZ5emSS3//oSzs60lejcC6CRZ3morOo2G4vWr5nTK+k82uk5tIEfT
pTN3dfOjh5byYfenh7S2UzX1384Q0o2H5Q0e2qFC5/ysRsOW4V/1o8gptchj73NOoxMSy7LPggxJ
5yX2RbAW5L/zTt+HwXyPMuGPvzIObzb1ESH40K0aHsTVtQSsFYSzB/tT4FG/ng1EzFNOKicscDpu
pIsgkp3wOShAeRMXPl++DSfL0rsDgXbIut8AcI0t6xTDTyuAKJ8KvVPhd6NFi8Gk2fPviBKbhmCU
V0VCtlux4E4tbGcTdmqKv6/dnSIaPcXSMMlvSlr6NELiQwePo4mwt8VdzkNdbkcy+6uscdHz6R4r
rBvQcQJNwqyymSUuGo2HK0tWOvVZk2ECPuGc180JymnmonOkB/kVbpH6pnmvNLFmaWzR1OqzvW22
pxqhOStk0qcrpZVaWdp68Qc2fkXOuAfPA1bVo0KMU2k1wox+T/2uejPR54PVlVGyq8VUNVOEQbyG
EZIIdaqATGfdfV5vAvt+4ETZMQFC1KfDSrIDP80Pxut1mtHIc605TxFrhS7mOMqQVCfI5NNA2blK
0nGSiNyNVO+9OxkZhJxKtL3yPFwO036WdQT0TIBA9BHFA3qM36rtC+f5Zyk9e2GdbnlxTZxBMITG
dzyGZyAlUtOF7nziQVLiEkXg1eyUqmkMb40uHDNWNeMHCH1Pbq+c/rMRRpd43f4R9mre06IBpu36
QQtBoaDUfbXbe7N+P48mAZO+DYQritwq+5mZMtovZcne2zFUlNJuXnbOXBEZwqDMoXyeSGx6f8MH
hyvxnFbBzP1gcZVlIOM6/zjrKiTVo3zjXnqAT/Ji8/awnedfJcmboSCSzqRs+xB1QttljfFBJK9E
pPPa4wv+6mzVlicB2MVMsemgtcgtCkpvayAlGH9yqRqjgZ2DmBNEowVaWPC7tL2epJp0/WoCOt6X
r5TBwoDU4B6SHBHgQYXOI4JyhNmH2KQw63bVucpjXJtCouXPl/09oMzAMxHbTyyjfxUquYL7qawr
5huQB0JMI0PHyGPMyrCgiuXqNq2FBRI9+gjApFkDaypjqyRu9cdywIGhOrH651eWziXwdF+nzdnN
AGhcX+D9SbZSXhOv+YHQCr/l09On4VM11WDhUbJSpaGkGtW7GyTtc2gmFExcq6NLKSt2SX0WTtbD
mYj7twZFtQdULOg+XTgpkAx97i7wNRK017C/qZHGKNSiKaPIh0wYliC+TD4tRsBCMsB+4gcZrKmO
UJo9ds4cgivg4n3u3XZiCEbPioe3NFRfOnLkUUpSkdgYy7poF9F6swuzCzXQdyoA+YCJkRI38l2q
nBy7Lii7fAH34fXCzRLUvgukLtc3esaCH1PSehdVcRfewWNMevk+XYYxDuubw/Txt7A9du1YHkpv
Q0tg4kDOEpKLjIArQXWeUWoAKOlURJV/v01pJX1TimCXrI0vaMODQuGETq7AGjiHY2F1hEtAjtDV
FLJ3WXaDO6zNZVI0rjumRysdoWOF+ovO7k2Qv/kSbHpFGTuGjU7dmuk+rbzrlMnrLWjWGKJ0mNeK
yBwPazSICt9OeNaqvYwQuHl1rLHkjlQgLfis4WuzqVMZnI6dQ0ikjgSu142b/nT25eI+cxUAAF04
MLe7sEeBgdP2hgLVTeTcA1ic55RXQ6+aOcMlRqx0/LI1Vnq5GLS75JFyB0NdJBEbZKgG8qMmwghP
+e/BH5DdpTevXzEgGahuk32v2Bnf8o8NAIDrZyuK/lziagyGw4UsafhFG6if8+S1QQVwACh9XnLr
nATnBGzDlRwEzLdNtv1Fi5qFcW7ngks4mrijBRFbddO4f/mzRFkSwYn51GnBKdhpzdrA1apRccW3
Im08O9By9UzKOKSRqywYm6XpVskrMtmHxxBa+/lwk6QaYp1qKMIrO5nhJzYPGtM7E3IgzKogli2P
6lkm7XlxLQ6OAY19Y5q2VDIbl8Y62JQeRHkvjdvWJeMCzbPrbsxy8MRcX/GwMIoBBNxOBXTudl/P
arM3Vi2G6XiZKkE7fApE+ot1Sf+s8D6Gh5KEHWiA0x20yG/7QwZOv8vBDQnQC+0LiDi69SAzHnS0
PdRcuxzXpPUR/gmmXNgC25Bxat6IKMbagpIC1kcCIIhYnL33rGMwjgK/ZU2w30Bji/sosJxHHTFN
P/r4RlA8V/yzHZGuSGiowcABQe6Q+1U/AZAkwa8Lh3pSlRmDbvpWGf80a774JLTROJ+uMxDfxM8f
yxxZb3vTSx4rcqgYA/nva6II2oC0s8e7/eeQYpnReqfD9GGtvanPLnDdBizYzmBbqW+OumOemF8c
YJnYNc7X1H8dsDl0H+mAeJMNhGkqeiv1mChTIQjEqGmxTHMNtsmsGpvsKnaqo28TXg7TkgyXvZiB
LMKWOD+ufp6TEhlCWtt87IX9le4leS2PA73XeB7/QCG2GRWFb+ZPDXhPxgGS3hyCMXsy6UvO94+z
T+jpEdNUGpIe3hJlkMTboNA6lyqzXJCqvG4lzYz2a4WgZ3y6g/CHQtJ67Iji0Vh2aNGH1L8jJIct
28fU9cTBtkTbpCeS8HpAt+fjzQebhdLZYFh/LWupgGKIMCIgKeObdnpB/+vFVrsEvEz37znDfgGC
biPujhIdtzqjGzwxjhEtCRC9qFlSz5x4Aa952+XLHt//+2o0yJy0PR8JOfTAnU9SYoS3VpdjQ0VQ
k8E34PgY5WWvRoHPgoFmqviXX1xszZ8FUmCMLI2+z4Pl+yaiKgnAbMZNiQl6cGKPuKO1LIayti+Y
vLFsFuGWtq8lnqoDwwQEAOPNy1ocwkO+nbhOm3dv4N2OKlbJ7nbNsaGbPP9R+0FTztvHD0Qej7wR
cSiIU3QZtqkoaGMuOntsgLBXCNGO4xeaU9YZ9Jsn/uHSkjdXZpSA4F7K4lkUtTV1whSNqjc9Seo4
qAdA1HTRwrMKGvS7FW5oQrT1PMmASzn1wSXc5jZ95QzcTn8rBQTzin69bU78N7i+52vED1f3QeBi
cLr7WxwZgLyTNTVnzl/ckYO52q/9FrHakMYhkPq7Jz1+T3X+63Qvdpsr2jt7nLNwOsBY9UCcGa1O
YB/GScqGZH8DiBive43RzW7EB+ZyiHwDhkp05M6/V2MZY7vdaFQIt+EDbKq/bm0v1Z0wRS+jkf0p
3a3XW9d9Fk46yC4HwyxZQLs33a0wXeuflPak6ddbBAR6cTvvoMYp/Wa3WA17OJOrvgnKYg9G+OMM
+8AI2PbmvHgZwQatgFJMi80drWKPD1EwWPaXkiRrZdB5tn7CwieggvTWdrqBpbm7UmY3Bn7RLxYH
VWUfTgrLe5mdtbmUblwCNX3Uu+MxbPvbkkimLRdaSlCwFT0cJisL53SwxorjyL9tIdlVoU2H6r20
mmrkC/EuWUbnN99AfQnWjb/3l8XW7+bO7DvR1hOaJtqcZQoiV56lOpETmusEzZBuvZMPKqYlciYN
9BAllwSTT+6JyyWR3bBJ+5mZJN6yHZ7xbFxHEAX4YU2Enp2Rfv/PVZsngbXHsK6IxfoKL127/E2A
hwpbAbCYsIHIy2z5/HQpLWIsOi2SY33gqGKIwa826qxxMHTrRIjfb1bTB5Vmcdm0dlcG4TCdbha/
TUz58oaaN4oirVHgHkh5nqHR+6Yp0ZSxefY32Pb22sIQQJzJqOUmwLCx4bPf/VFRUc68KTkhcIVq
kSHUhdO7sTEP17l/MlasXf1wxiIAhWblOx+iW4CsJa0MXIgzXt7Fndtp4vrZGAM2zsfPBzwdt2QK
uY2o7YclpMnGOGs6l2kqeuQ+oI7nld/40MW/pSpdsd95Wiof1simVR5ve3JmPlpSipln+aMblbCS
bSoE9CTjcY3vBz5Da2moVGgMVE/dgpW9waYmdXfoQBdBNUYCi6/eQ1QMM/5glrmVpWUPGu/A37Jb
m0w/reo4BrEzH99UCGD72a60RgqovOJEkfCBlFOZKAedLqet+j7ItAQ2AqfSGz9+cjyNXu58QbzO
uW4GUlhb+gv5qktqZvVynpxnkGkDjgdWzE06m+RDaqP8WBa6EEKmYDfB01OsgtwS8jnzj1suu95A
vLl1hywCb8EUjWWCL94gvEzvydenJ7DaGgGyIz+vGRU0MgrlnUsZ8MbjT8GJTQkG9iLukcW50QyI
0UPYeKduyJJkczw6e5zvUahKXh33Fd40qQzmRPB6T86Q06/GhiGrusdzvnt0PT1tVxhBVMtLwW0T
ltiD56Y1+6ybwioRs3itbwyG0bqu7fB6oRmpS6COCPuqTrHtnUKf60BPjqlLuRo/ckilaVHwI6ds
zkjfOiM0tt7Go3cW/j4ynSn+kkXfjlJ7RtarsZyuPWultVZOd9JJwpfiVaxOVYCcjA0UCcgSyetP
ouwbctwACYMi8Za2wPY9YJ2dA9HBZky+9XpnclXYKvUPsNoWSaqx0fchetaz6MDuAkamHvuGkJJl
HYNZ2iNAYJtBXfxXJpVa4ZTDiF+gzlSd9xLxeFxFCi27LlDpO/0by/mLdungv4BAAqu82ZttTDOs
FAru5EH5mNp93DsmSSEHSRcGy7C3ULDYO5CVXrW5saG/mmh5FdQ8nnjJ8fCq8qaL7D4VJkaTjUHV
wtGGDYv1SlkhU9OGZRckgUghtWMaf93j2XmWm6iJaV3EEozIlJmPtn+hGQuB704gqqUQxjgaQwNL
qXWaCIyb8t35azcPL3AtBKVZuvQQYgKcGnLwtMRTKhuJ+5nko1YHBK99xRliFK9qnHnZX8a084QX
WVHUDMom53tm33IB520p4RoFvKT2v3Wgrev3Y95B0xhMrWr1UFiawTXx3znAAn1DgEIBWzYqtfot
Okpk2rEZBDf39545GHqmOI4kXHctbLB944XVFDnnzSQS7QqFUyHR4CmjvDKE5MhAQXFZmh0N7zlw
4uxC6jGkpLKF/hsIzN+ZhbDaf+ofR0gSfk/Gh3bbR1JFZTKqtGlrIIXoQaUgy/OeYNwgM+Yeb9la
wWPqkVi/FVbnSFSgEFMjmhIQ1Oghn34EX84h35J+GpC59ItDQm9CU/Bs0A0QrkhTh/84Mj5ZgZIF
LfuAWYvzj22N2RD5CyaKygEYo8ntz23/peIfVmgcTwPPthMFhq8QbBm/k+/xbCAQAGH3aADW6Gto
P10HsL8te1rGIWPT46kTwv93PFenG0Y7oC7vsnVIjbvRLmPnn4uyi6pUQ0onNm9t6V2mZqzPICzT
hfgh+h2r+tQhREctMnh9EDmrZijw+EbJbwwbDeLBNYR8xWyXKq+02uyZQrKZgXvoLiUFSU9EqCco
JY4BTAxyCdXADKaRAncS+7Al6kCkcKh9bSX7UDgmtkeR9fMgVT698YOVo5s7iOBY7eGGktchNoob
OGgf6HWKFQtzPWFOL2a3bTN9w1H9phtQJu/u8W/gqomNU1WJuC2EfPm4Y6UNoyuyQO1Lc0AML4wP
7+R9TbWZz0ufIwlF45SBWHLX9MHerUye7YkoFYI2ePnXAZ75+tijZ+9cEnxZ12PW93mjIRo3BB7B
rxHVIM14GeCrScsPrFqm+wuQd7Sjuxg/QJpuY02e4iygJXokBzPOhmm7+dAk12DMB+DaLBUJDmKs
xcGvVhuc7SvnafgaxE1rZ7zljkovZdojnDzx5qBxG6To13l5JjmZVZOk5hgn/LTx0xrxHoj2VhES
wg30P2NmPHnX0sM+IOnKPIyiqJongh3AFD3fmKbDzd+saNd+uuTRKtnOlvzriERlOtlEUUuRbbMN
VaQ+Bror6Tf72Uya7z8vXajFKTCJserVIHCNtRdIekmN+3ZYxV/UUc2Yg88j05khcxRXmTPddTbN
OP0UxxY/akCAt7RMq9XGLrDzDpAyaYOan8euuSPhXritzbuv00wrGb4bwmeCwsiMXdV/C2cRK3y1
ehfF7mBeReXRhUfvIFu9N69qPkcwRQvjAIRY41AYvR4kbbotLvIAvdOTSPj7laDHMpQdaXWmDnRH
9mgP9t6leyHHXjHpUZIWw0S72w80+xZcwDZRlt97G1tKZXgu++tcFMtFi0juhf3UFxxLZ2/tox5X
jZQVzwBQwti08zfQj5rWekdsY1EUxHjyasSo3OoY6vAa/f5qCEpYjr5O/9bT7teixn1hbGeHaAJW
VQD/9OJw1rH5zlrWF+apHV6m6uPDHNvBiPLQ1XQfCWlDW3FmCM7NFbXf7wby+Bw8Ncsl6Vo0e4u4
YAh6RQL8AzKrh6a3M5iK6fvgS0bluJJ9k3osO/rnr2H578GX8HlpC8cq7B9vshalaH52Nkgip2IN
8hd44OHkO/+qgQ3VpcGsASq1Fu4CyJSf08T1SslUDB9bHKf2WW2XUprRRrG5tcLYKaVNHoZp+MwM
yWvsK++LinIxovizRhex3u+ZREo0C3uPbNHkylbB/pIcxlz1oBFYZGMGrRU9xUUXdsIzoSW1cE69
HClVQKlN0H9H6nlRgUG+4uX+wLCOwDUWEVQTrJeNbHxyEvbaVWUqlUKzeTO1Yuv+KPOeLxShYZb3
VKrOS1YQc5R73ufnoErjtqZnYk88dIuS24pJMw5PtFFnPg3sspc+pp4JwOh90lqISzR7obUTAneF
2b5cwJZpeh7pa4GcdgiPYvGmoCBa1q+A+J24p6s5zbKSaxTuiBuVa/HQ1C6wcQ48Thwkx6oiVFEt
tP/YQU7SJb5dX560XUg/ODcIeDyQ8krvB3v5HOMgH6M7KznXrS7vJhmtuwT7fMJAG04Iszyzf5yV
6a3NTfNxkXNeZeT1yskvO8FrunOxWtN/L9vzh9GyPA0xMCgQJn9RmJQvVHBK1WJlpe3I7oZ3G8mY
Eg1aUbwRRtEbI88bFfbeaFA+DZxWJu57rmCT3QiJLitVs+ChwfHHFEfBquAhfD+Vd+FyJ0gHLHyy
MiQWjcgg29XjG0+b68L+nSxGeSolFP2rGT0pPDNOTXN6oFTGaq1kBWJTz9pXZ3OwtO/ISRJbQqbE
OZe4t8nYUAfCdmV/RnPUkzywnVM031CAYuGVPZq787ybcMTiF8txrhCl5EisxiAN1ld9DQW58wUf
MGRSxz93EspT7h+p9Edv1Ycv2LuZDAYLnCr8M3QLlqGJkUjOBJ10WfS8P+38v30YT0MQW42ZXlUb
QGx0aj/65D0edb5tJeFvUF7Rt/W4xPIAtkE6eb7BCF6kTMMLu5A4HF2B/AE2cLaiTtbBJLAjtY6+
EpkjHotkKUTqkr5HwxYpUUUOElNxZh9MczwrZo7ru0hslU1HusOnG0ZhEJmRK6jNrSHFlX9PxNMG
RcswctbJ665fE+mAi1UYusQA/i/yhgOD/sbWGvyO6hE7iMDeZR02JItogHwmE9MA289WTRh/MqSo
2kKFJFmnYKqYVf0UUcwJ3GN2eay4JDpKIn1r3rc4BirV6sfLEWDqSP72UNng2epbI9BWJQ6IPJhZ
1c5dT0jnE31FvkQceE7f3r090Ef+z+ESiCeMJ9s+//A3GZewg5rX5bjlYPbJEFb2xe+bgLL7y0as
WvfPzU8lX/v4eJRqV21DEJVSJlo8eeGMXYDvB8LM5O2PlHO2X2KP+n9cL8AP+SG4g8elrekZgZMW
CD1Qvx6ctgD8kd/1NVKzqO+6MrADTQMU6Vx3ZFG+9sDjt3g926k3ezNA9FkVyE9L0u750fqHI2/c
dX6iZWgo2tFz3ThggHpsSAnnbyyK3Dl4yFKy6JyAGIHofGEKN+vn9UzGUVvTAn5wonm/mQt6fHQr
u7V2rIyJhMvmMHnh+EY6L4/vFXr2o3yPxc5EhlRSiwD+y143oNuEwI7/KIU1qFoDKvKk0ZVMR52m
6N1mplyDc3mWM4omlJ2eUJNUa2VZ0KaTTGKSWKuqjqNV+wBTk3rT11P+A7aCPowItWosKnNK0ndU
7mLmOnSj/Gnjo9hTVpUfGHYqDcHMTFlAfb5fnuteqF3pMQKLjiOOHynsN6dzXQ8Cmco5o0wt/6ct
9aUVeTIq/GekdIOlU7YiUXD3a6t+AQjlkJxAtqpDiXshGF1Db9KZ1OrXhPR3Lqvo3t0yPk7SVJ9y
E7Kocx7CjO8XaEuTdttgUQXD1XhK2pFvGdTUdy/eE2YdsH5xzExmfOXF4VYXqcJ7LQwCC7zyY2dC
Z8o9SsDdlU/b384fRuBtd87is2BJCCvMi6NRp8TR/1sWQLwOXO7+6q3b1Pk5xmu5CZdU6KeaIJXy
mHS0kq6BXHoYNpL3UeHQ6AaBwpiPWzGftKWj+t1igfeexvDCdabHxonUk/GI+L9pHbQ55AOOral9
HBdJFijNtIDXe9foIlDb+EtSg17DYkxBQ8RFotkV5I2HfcJ3XdcxhzuzzH0tg8THk97mYBBFrj3Z
ymwm0vzmgEtd61+11mSfKGojewQIMnSiTRDvyl4OyrYN+4TgSqlp8/0DnMCK6/q8+xKuFAaaylBK
dwM7HSnLQTv72evcVN3AwuJONwZQ0coBgrNCCyBCXhXyAJLzOY28BDauUWhVMgZlASl3jM0/TES7
VeToYjTytrr0PSDrztbn40bAun4Yp5uoAlQS9OzCFZuQeR9Eh8Pm8NAl96TfFUHU6jhMb7hvD/G/
0CCWwYSZOG0dPNirGN7WQJve6B2/smfPlrETe2z3stxkyhWanxlRATfna8IAojrgWYzg+nLRe8wn
IFzJ5fZt1zCMqIDjWECMno8FZFMR1vPR+1emcRvhaq9jl5/h9WP18n0yPywkNsdtZoo1kXKkRG2w
Js0YBM08oWDoluTx79N8M+ENQEhx0zx2MV1VVkrKMr5IIccNmQU83lJv6SOTScFxTIip+rdcUb+P
SvmLouBHdqeVpCXct7oVv4OCJQCw3drBycjFj9N6DbMsEAAd/vUJjJTVy2pc9atXPgZcGhjgfppT
g/CjJS5fXS6rqx7xAktyMEdP3gr4I1/2Pj9bB7YrSgy5boNjmaaiDnXr+br5BqdU1DrxfAxULSlu
pzOolEq0nvEr3elW8E5Y8WJgdQM3fKIL5p+PqKFiryTBPmrKnsGG3tIIlFYhAYxPFTrPi6XeZauu
pwrwKDeg3pm3bKV6eg33VjgO1v78YPtaciTFS8Pnce+w1OTLvLNDhsVytHOVqeRrcivTW+ibQ5mg
i8p9cdxGvq2ZVTlj683/SD2jtZoC81J/kSbEzgULH9KX5in1/MxFmKgfzavKeJ2iXt8nJGZXKaFc
URnW0cG9oUZLNP1P0MwISYfApNK+XNssyXKc4mrLBJBOMqx7UoBXg1Ap/FyMC020eXwn2rv2qVEL
OD2G163jkZb+as6d/x2Vw/w2c+mm3Wggl3/BYgahIybXOq+StTVZ3x3dmxvkTVhaEB+N1U8jdwcy
SXf64l578+rrLkQK0Jsk03jg/WlRlG1HgewWXZzRGS7Teuuy8LQog/Abtb1AeWB2+GDSSW9O2J3x
3EVyZV4qvpuZ2DflEWMXDwqCCQK8Bgea/BMMxAdmxBM4d1dNnSB+xTjuSoGuZGLKqt6iJDAUDgTQ
uvE0KBFO0owY45uK6FR/S+hLoMhsk3F3d3oriTdba2IUzul5VJO8obNS4yZABdEzgKQYr27QBU8t
YTHMUNaiZW5vIQ/PV2/JzDQUwxhyjAbW4EOT/LcOWV+FlHv+eWuGreqSjaON4GexWCYxOciX17r0
7iUyHw+no0zw3VbGeEAmGvAOwBtuBcimRO7UIdq9je6fpfU0E9Ls/Nri3K6Oo5FmpYBltwtWmSVQ
w8/A04It4jAWuwWfx8j1BwTThAhWkfU2Gswvg62cNJAhHfva8Az4qG+ebzK/+UMiFUyNcDYTSTI8
QRUX9Q/FbPWmtatXd85UtwW5M+8YOLqJg1Zu/MctMd461GmSqMgU1buiP0K6W94hLJvuE29nvhvo
YZiPPEjQbJcGWfAJozH/gmheOmswTi8/D0LDPVF+NftXY32oZtI9po3PMJt0Fm6tL67d69jZriub
YK3txaGRcwsrVraLcujI5Crh1OO3o5Zt58h+xkw08tVc5ZQlI/P3EXtHYmIxs4sA3nIsJyCtOc0w
fOzqmzwECFmKzVNNJVodHVe8fZ7fqhYhG0nRxTUDsqIw/f49bwQ4sVLBZtIW+x1rb5PwouU0vPJw
0s1PFXt5xjBeG8FfpjxKImeS0sjtZfsLVP3dTCyICtPX8Z/DFMhz1vEuWnN4rKpX4cpfZQ78ZBj9
fQvU7KiKEsoa5UHbUxATl4cO81WhBnsEv9yL0Fbrs0GwrsrGltz36xlszdiWa2mwt+ErY4NuMnKA
7B1iRBRqci4qbgOxd31PPFIutdv8HT8hIiGDD8O1nG9WJnhtuOujw1/a9XjhJegrjmAw3xtg9H+S
0wHX55sm5KqSINJZBPIeex7CtMyWP4nLGeNuypZzY+QHvNu0Z0XVPH6ANzHrzy4eL2y3UertJZOY
0OgYxlpjWSunEVWT/Kg2QJ5zLUf6QOtRLsv1wDYi5QR2/1Gvps5YIgnQkGtlMgXQpK4sWzjfDnRg
MwIvxXTlVA0X2Bypfag9hOFRMKieZIeYNWlnw2LyzO2z5E2df64MnVYrXQypb3MkWkgbEiE479Qz
dMvjBIN8n/rlzEPOXaSOMQIQd4wb5BChqkwpunoBxQ+p1xwKyYreymDt3gmHmAiKBzYHn/6GY6PY
n86QGYoeetyw0ZtqNp4Cd/nm7gPdZY9jSaF2TWScETfC9iycaI9pdsNzLkofFkxqMrk4jSGf29fz
X+UhIJO26ek1x1xeTFH7MPv48dKJ2kTsgzVvNxxDKtHU+xzJvwed8j5H/sF4XUn8A2JAmiPC9zRr
0jyqZbXzVCGPk42uIaEU+w++3+xTKAvb9gg04EpDktvXNmmUJ2DDkwvMU+iwTzrNSfbCGE+WtUPT
JuxjoENQllZGVvTyfMEJrcTNr3WKEktQC6L9Cb4V8Ez2AY6uP/vAODjU4T79kQAyRg/gsjxCtUBr
pGZVqKSQ3F+U56OYfbshcO0HpWnKErR5j4B4pRPy6IHUOmF8sehOCNDxskD2LbqhcYbGSkLTFaCn
4YJ3yrC/3HNZGk/aWFXxzgoRmre4Y4Xk/YYkzKD4L0/pzWBb/aM27EHJliTcfMl0bCDaaNU/cN3L
6D+xtWQuITWEzF2oE2R4NuRXFB+TjG9jLzti4JA4HteXltcSLw9JmBCXBMz51CSZgArH35iPzUTg
78hidqegP3llOYFyQWE/H7kmufhSAqw1x/9NR4ZkHcwxhhy0l3W3J5SBe3RDEAJ7AygqFo0m7ia9
J68+HVHtOJVIhNyM2FMVwmA2r04e9blL+uZbUoSSP5QOj3u0VzUMcJiVJ/xgG0L1krP9qBlPM4Sa
iRqYvAtrV8hXJVki+VhUn+QNBoeIKhGKtDBfc+JVTvP4Gw0YcYOQo3i+flTMrSlhtREf72UQTMUZ
Y0YkzC2d+famxMZRpnEpnc1JvUZ9JEyWqtVMD/BOBnm/XVXEKxKlhQPl5B6KDFQ4fbZ89JkGi+4L
qs/2h3Q6yBrMARgbGewMT7iBspIuBe7MUDVy5KRaBp0NIThvK6uvZt3yHOs40B+5IIdteMcLNhLt
ezXZMfZIWg28uomVrNEFaYKX3Dmc34crVO+LfiuSqzVAfb2rNk3lI5cCfY/IUw8ak9pWn2lm6fJD
A4W8MnCWlAe5xNfCCaKxgLm6UcHJOCCLf0WLLsILI749OTGVWG1gA8ICQnyzDFx3YtwaGIWC6hdZ
r6kArydwghWbnC3ahr3/LVR9F8RGpwTuMh2iV/m1PSJyGDx8tMSCIcx8d7TpER/vV9wCZFisTKxe
2Sy2E0XmwlRBXo5CCtDHVTP9OE2LalqAoykBI6sTlkSPjkQbeBDIY/w4195DUbGeHnrXwu3Isy7v
MCfvpnUZA7pfqv2LL7KSpC9V69b/lEuVSTG+Hj22qPO+hy7MHhd5tg2M9qMoveyEd7tj2FmzxIZa
+J8cd8Td7H2R8khn0SiuQNTmeiCvI0J5rWQgPkRXGpeBbIopPx26wxxBWoUiksy72W6DyPLybQ52
/10+1IyTrjLXXP/jOGMMY67UxeGM/zPeYiSCOtLdWyvpH33yj6zKNcaxseGN86jqgvf8anaB4DbX
AceRo5WAN9DlV+Ji3xqdNxv9LTU+H+/yyXd6DA0NDfeyt9XFydIN9/VG0dufRyqWNxzip+ZX9E7Y
8I0le0HfbSD/VeUZunk7ezBpfhmWt7W4x9XgAlFP9/OeH7fWWW99Wk752wrmqdmHNAtvB4Bb2R3U
xdOlrQLaF1Plv5pY4k/uhtjncsrkV5g89DSAfWYcS/a4k4TyWuRMlzIxw3BhtoSrDM0qm7BLCqhi
vGlNL0ZKmHTcGJ+5g+pg8E6gqZ7GpdJ+Lyd8WYw+6sTkTr9CkD+Kv0+/L76MwFtRIr4N9hKerA4l
YSnA0tfzKlQs3tv/P7Xujerrrwf+miwg5x5X1vUB0rLSzi6TxjWkm+wQl4ySStriFE0GZE3Nxj3q
Dazi8+nzEwldzielqT/MtXv4txdZra0bi6RwqGK66gDe5TF5vvRc/EZDSrxV4DqwrXzxbai2wCuv
Ovu4zczLDHxT0IqpAofC+go7wXhboGnzRJxWVBzxl3GkQ+eBgCOrMp1uh7R9DEoXyUKNzTOE1U/3
OoDlJaVcjbL5+88zjGpEaaWAom9KqqB/HgNRmCHVTYbQ5TZCr0BgnNj9n4sJCxQ+LdkygnyDu5cU
IpA8TVGPcWdDNOBbr16Hgqo3LODjmWc/wD9qENnQKTzOzmmIShLyUzpEPpTfx8NM1PFHnZrxLRz/
yO8+NKbF4ChdQC3EdKdTpCk7omFCed09fiExxXhP5CdfOqzrWiM3lHLpLdh54QA7kZCPc0uKnaGr
K2wseBgPfSJX2cG1mn+0JZj7UThCwcsT8EpMSr3mdddqGFkEHEkqmXItVPeAt/hnE8W0OR6TkilM
9hKeZW5WHfWreFxUwlmLTCs5m2HTiOK+zOb9X2r/VV3pX4Rw1vYMB+Iiha4keKTfH+ZU4GxqhBny
zWGEc4n9rKGSO2CZUmMvPCUGCnqyaJIKCpOEeFjOHz3jWsB6aTH0Qogwi4059kAhntnemIKUnbFp
ONauiuil0taNh9xOWR7V0c+B0+2mj5e4X9tDIHi8eRxpFlmSQLKT383mU9UtXltMLMFDbrawAgX+
Jnhf+1nbUva3ma5JnsRrUuUF9hNhk9pkYFflYmvQFolb7D2W2eDmmnrICYif18agZ3/e9ka2Lir+
RNl4/p884Gy5WEostKA2r4nv3lRm3H5+QueqTEFZlAM91yJuZmpph36ixYZbiqA0RDVffyFc4KUD
edyqvRYpqs/BCONQEdz4y4JPojNmorlt4S8wWXn2hP7fwQqGr2aqK+zSAZ8jKQ8jMtp4fDCwUsQP
IFfWQsJcoi9Bhe+U1Ols402CuU26hSHcWaNMbeWhFfTn1zLDHbWlkAM+80aVkk/yNKIN2AE8jl65
qSUBaHA2ptiIs0Bp6/LBy1yMEqxVo9HLDUWDRlpMxl2FJFDoOLKqbFy8ZHFMrAin5/g27r37JzPq
G9OJCr7uOcei7GFjsQBVeol97LeVfp5IVv6WfbhrNkG02Vk0BD5F9CH9R7APNmH05C+5H6eczmzy
q1JXa4yzQDHo3AZ9LF9rqIbFftbg+oj+SjPDGFb7M5OIoAZjVSg8rJiU5NgJugmzuGLxFLU5rPme
aFNFLzd+E+56nX2w0pHntj/RSOiK2wZBeNeusjCRhQzsSUyMtL9N6M6mFXMBkZqpGp8y5nG/0y3/
fvENnw4mOnih4J12OdODg0KA04wjIvD5kXK7Mru70o1zZK2MRBb0iYxfCq4uHhUSrUJZ1/Ki7o4Y
7WQdFoCmBlRgc73toeeoTZTq1gWRtkjgy4BiHgQn1KCamMn/B/NrDEXG9t3pRKVtw2EztbdiYt3X
w9azdIdvxMoYRmWi+ClJhcYMRnWgLcOV8i5yKUbu90HhvRqid1WtIGMpSFLX2H0qtLs4dfG9jiGj
Gs9OJuCpW98hRcQq2GQc7bm75EEfN9K+JFVs8z67Zz6/U/58fTsO4fUAfEssaE/4irG7G0UF7wyV
iF031i7B3lTRlxCbNWMXWsxl0SJsHSs6uxQ/TzZDIznz4hLolR5zvT0NKM+H423GiFJBB5BFAxYs
ppe2juCzNFTvAxosND0duuAV8aPekUQILwzEMGcr6iDOZZ6YUCw10mXLPVSy3xqHxKeiqUjhCE0y
J8IhraCsbjU8UrLxkVYa+ZHyURlD546ompZFI9DcL8VmHyFcKx/TD+QZ1rDCY7b1sdam6YWsPNPM
ia3sY3XT8+LsKwtQllatWAmlRIrwmMiI7Oughjkq8xIOn4TtvHQ8BWSYOiJz69m0A++jQRul9dg/
k+CCBB6pxNArt2vV01joZBtpbAdiLrvfk8SEKLL4RvARuSDq26kMOR1q4C8rHMbzjQO68Qxdv0nw
FXm81fZJdE0avjQWXjoPvknjEYQQWnaPQrl2TBa45CjQNl8La8WZH6fniLEvRPVXJYfRBlkosTX1
Xr147MclFwW6eOlk0ekXTuevsILRexz5s++URaJcJAA28muxJV6fDkPmkhm+GimnFI/XYnpt6GuO
/VOq4V/myp4OJWcyFxCxMvWVZIS1wUTwfMmok1rQfV2OABNPUZKrbN+GOFXKTzTDxx/ivqJR6Oje
LMVJhFoT4iLFgZCLTzAm7errB67Rm9O6QvCVjiJOl3J2Ukif3VnlqrdhwDhjiY891ynsQZvJrgTR
snNAZAYOE/kKLLwXRhZCtk7CiJnZjRe4JBA/rhyfA2nbTVx3/pUtmXq/u3yA93PZfNLzvHlfQMOh
OSjAbgT0T6QLRXlcuqGdro+U3zESFL3goWEJ26mdYiybgM8ahaws1vP9WMbkf8drwyIteR3uHMKH
HvnOMi06OhRWyltY4duO0HDt47OROjow3fn7a1AJKlIWdPR9SZ98j/2HUjEr4O9c241FVDDOiF0V
zOOV0Bo0Ik1piMgIJRVYZEhsGb+gfG8gCtN6ymrUD4zrjYCfblxwyFYk1S/Vge8E9HOse7dLW8G6
18fGOLMFHTMHsduZmhhu1cnEO8iVGo05hYhXCEht8iaB0vMOpPLTUdx0j24xbft18AMJdda+LN3Z
J86JHBBianfYAPP8tEW4rflhh7GveGytwd5RvbfD4tNGiL2HaiAljRFIUrlaaWAHg+f0D5cWnXe7
G1E2whZC+qPzq7jGsZ6AeKsDD0gmWUJWi1E1FX6VGdGGR101BDTScblVy0m4ZUNUBNDAnWm+gGI4
2gkclC0amEsYGXTu1lgfWJZGPHvglWNHjCaQbdAUeB5kMTHzkWIiV6w48VvJKWo+9qpUcAH4T1R3
ucaqD6zRfWSzBgJUp9vhOUCjwURI1CEv5S8zYiqqP2/Zy06lnh7lvT1DGt6Q/xzqhaSMYOeOwJGB
vrXVYIN3gyRo03mRBH614+eHG+0umeJCnQBlEP/9SxaydOXlR1nqqB409YPgDxKnxICSXIn7gEzF
gJ9+wbnZt+yCzjr4z8fmrCW0fDqPyIsf2C4s1RuS58pR0pCxyHgsJ2sha254p+g5t5tvjelJncZD
0WLaMB2OzkGnDgydIR6jI9rPFS4G4CYaddOj5qprXoJA+1A0Hhvuo4lxHSXnc+HbVJI8AyV1IsVY
v9UsPY51MLsnvM6+7JXerU80pL5Hd4cQBMTrIQBtGVHo2PSulDzfHUsx/TO+1GvYsjFDvC/+TEoo
eXmMJ3xoY5RLjKknQIlDUFlpGCFJqaUIkzf5OwtkTOWSjJf/prTcRUkBHEGGq78Q0y37NVjlWt+l
9WhsnKq92Pvb1+9vKArL0ylqZQpcgvaAwhu57YDt7oC7c28V4zxuJBo73kQLIUEB2akyV39jq47D
b8Ycc3UqfPZ9ukqnXChp8rz8vZ382psW2u3TUrBF2HC4il+GP8B/Ol+A6m9XJih6e2/lKGnPdUmD
v7XlI22j+Ze4c3z4icG5bLyiHTEqojJlmyuOTLUNGYzhrG0UENQ/IVE0jPM+RwbKjDCj7rTFstm4
EuY6lCAy2oc/MxPTniMDg+JxacZ6apnpJ1N0V9j4sn8d0ICaOklgufznsV3PB6wzlJgeChzZQfYM
s1MP7u1bCKLxNp8GYkGA4C54p6tFeemLen+nVL0fbLOfJpr/BC4Qy1BsAh09tPTKERqdW/iYB3sM
BgZgwczReS65+lMmg8Yi2E68AB1TFwRKfuM1gLtW8EsC+zJNogVw+Zhfr27Kileo6MW8BXD6DDFH
uoZ/iDx2V1cjv5mIQsV3wZ91VLPlZjimB8pv8KfGjbn0jVo0yWPBRiHotEdRjIx/xwwukquzdUtJ
RSkcWWYE3I2KPLvpvRyz5Y92lZCeAXtjYTU6hgPVdGilRN82AnbiiywNcteG8DThmPiJa9FGdZsb
10oaLgs8nXwACCjt0jbiirH/3q94SZ2wSZgzUm57s068j1+MzCv/J/n2dNVV1x0xdntoRyO9cQa8
3fqku3/Vmzi5rwKsTb2HBX3XpR7Cy38GWFtDPLKZWwgztxaRkWD/PUXFtu2cCRQ5jmOsu9hqyhtJ
e9yADZWvgq/I9r+A3cnZLBiHavFTaea7PDQqcPRuJYfbHRc9rQ1e8kXMM45ewIBuiWeptHwim+BE
ZlxkBnS3uiW2q1IRgIJ3Jxfj+Hg4csDzwoiO7N1WTgEpdMD0QVgRjGVEDUNud4pRhkBVazmX969X
bBZqjcCCwyIweKWC8uD1f3WvFS3wWZBkXbkvBYsB+1hQLfItz4f/Ykf0suVjteYATxzc3cFeMEe3
pW1YKjlMo9CmVPx+oOAbiTbMDJQjQE4DPByULqqwdYu9DzE+73QtgI6CxiY/VPl3zvzuflZrRJwo
4MBgUWpNdiWIEsoIEv6Lr0YKN6Ctzj3tluVfTP3+wwDP0B1ELsyU4vhpseegPCb2eHjgSFKOYBG2
GLpXqeGwtN3DFzM/sCOZdrLvIfnZ9Qtumf7VeM3e10o0qbM8PDcUl83nQQjteTm8RE2qnOoua7ZA
o41jxkQtYLCCmls+QiEdifJ5F2vgwVdTtFDaQpaXXdxOlDcpM9q1yGwpQEaAq4UvbUSUHSL1IP/l
vzazrLarhH7ToWba956Ge0d/XFFSWrkgUC3hb+gQLHnDDcW8x/2/C1RFdRIzoGBXgKVNpVctdaKI
h0MEv6bluI32UUBjRLgQUlm97qYxbjtgzSIAyJ0SmKR42EPj7UI1F9TpywPumnh6bSuqbwhRc8Sv
d1gUSHCQzp3lmZQAkvEGBlNNcgEp84XGsfGnOGs7FroXabITfF4v7xz0anZBwTJdMekJRjKHrL/T
E2q7yzr+O3nVewb3iX5uN+45PF+Gsq5Ka3//mO15Khu6c1+gz/A+fa3fLED2hRRBdPERw0fhT3td
NFntjbMZNYI8H6b8s9S+RcCEzegsdRwceL251hTc5FnP90wfvfKEN4fuzySdNPAaSwObXMLPSaxx
6TkJIAhjMH4rksdmKTRJV88z/7T0FS+FCqNBbok0MD2MfL7wzfoP5gNemKIJgmM8QdZ2HQMqDbK9
Ultaicqq8SHjbCqdjwQGLs0E68QfiNkOlNYjC+vp0AmvDVGiNb54nLpRBXbipz5iQx7fVBaYcuNc
+8HPTAZ0L9i2eHQztme13q0kzx3Ld3hfhNyM4NI65VjEsieZ/vOBm9FYzyea4xKqhLpyMkKIHzZD
+V5PLHSMGQegAIvIpGjt9zNf47uud39qbV1/0Da8rvfhb07MX9GJdEQK+fFsOpZwl786bFAedmVx
4d6LCGqUipaKj1nvkK6YLxTB6J4p34YxRSUOWVqCncIdL04yKs49CvflY/scN5i7GOqwW27zDbOO
Wl/d1O8KLQnWOmiJEwh9wEf/MUYBc9uszxXh+BfXpjJngKP6TuK+OkmDkMVu0UqBNn92VHJ4SbFP
h0NHTjn9zCVpHdcoANHjTAuXX7htfWK0m6qxWeJHaWNd1JHIH01SBWp0utboVGKm7BHpDq2jvTXH
snsXfzHP+HkjhlrIOy7XMn/FKs76GoupTc/vPvfHwT1NW7Uk0F0MP3QPldDJjG0xoN9yNiN/5Gmm
YzWZfboYDmQJPml1QWsWGQTtOdCZHfCoR3V7OtbjtdUblmRH27ayKGSUwOpSkpb4iLpLsS9ODrlD
tcu8F/xGDs/du+4K5gtn6IGgH5FZfAU4RuDhC3DPZ4hctkl0HujerlknCSTYpwVIR0XG2m7Y2LbD
Kdj0x3tGxi0AdmEmSc55Szftn/pC5IeC6Uoo/vjATf0BzwdbYMDoI31pljSjl/NU/TWEbl+i4Aom
HTaTuJqQ8HPm/bd5KCiuXVvE6o9d614qAT4OZNqawfKGyiWLE7GssnhNowOutdDEy0LslSyEYKaH
HchyXMUZSjk/mG9T4rrk+dPulbYs99FtjDCjnhFzxVKlv5S00wcEIVNXSWHkIyXWVpnx1FuwjzbY
PG0jIH/QLyc2fke7JzZpIhUmKgirKn3FyEDbTmw7YyAugeopNKchRC/JbKiw/Y3CZCFtt0wBbMWw
w7v1cpJ9HWDQH22RPULvJmYkU0rD+lsCHxWfylXrvC0M4rATflZ9rI4Z+OVQqhghbzoz8aytAJHy
iXRLIxK5Ax3i7+BHijDxPmrkpEgsLdwPI5MZNJVWX+RWPur9eT4OQtipSWxVQ3sIUyj5nnzggaFp
GGFwGec9KMgwZakkrvVPVoK6MLgsXzBllzTv1MMypZvOtCaaFN/jg01rbPAV1bIOTe8bsHy9ijgW
6olInXmzUT8r0uuhLKQMlgG+DUgXShKkFoHO+AJM+W7yQK7YFTxQFY5qwooSMCrVNxv4VBjLc6RR
Jq7yK0fnuNK2IwA/aTyLO0o2cNsq1aMOsFPBBIFclGojVa/M+jSpNQj+aiVgH1odN+QNGYbUbW47
o86/RncJXkUR55bFPAC/DxYPYpnpwMwXjw5mLBiFp6VedNY1wtIFhH1TmgzHG6E6wyDU/BcrebK3
FxFNx/ZQ870uddmeHxT4B3G7wgjXFMzSHd35DWmwRia3SUBmdNRqwB7DUZeF8FBMXID3aNKuZfbE
/+74iCDewLj4/pMuNRoaEzLdtkO4nu5fwNyuJvO5aPZZWk+cKzRorVUnafseYZb6vLxI8uhe5Pdk
UDxp+1CVDlR1oxPBWq4kQ+Rero5l9iYY0ptcSjNRhCr/nadZJE7q6sGgrToTZkvp5o+JqOhuiUne
eVs0/gLvRXuzPYJ4WiqsV5GLtJtYq4QeMNCfQGJPxow0AGnNcwVX6SwkHmFigi0kgjkMQhTFcA/K
enjvtpeMwGcvtUvVMf9q1SQ5QBGmk/k1I2AsdFVkPY1Ft8BWAHZg3rt9U86eQc702mizlLOGpeG2
d2i1PwZPcBCBGpGIJ5sbaN3TLwbPrkCI62WKoZGvDZfxBWldbBavnghZMlgFkQkAgJRLYHBtSVjT
3FfTbTtWwIYI2/ACHDbl+NMndzPogxBfsedtw6UPXvlqMhFCzSL2N1WkuJBZZaj7U5Orn7xfBG9j
5gJ3YNgkLUKoDJfyN/d5EaKJUaJhg3GHXeh46yAUNbE5Oo21icmQ7i1boFODijlTdDWOI61ujdy0
xTfgEtqvUXdWa3RqsvyeF4kw/SAlchY6dn+N4GXS6ADBLqTBFXRxkj+MLOIsO1ks9392Oc8E/okS
gZH0ZrfucZVER0FxtpM8SAAU0tOAIcArYXybZF+Ca6bKLFx/2WOlv4iRxENvCLA4XT2pRW8kCNdS
NFv3qX5ntKVflDnTnNg8+hpnOfPX5RotnVBQHs/2KHQK335gB3xykJVSR+w7UHi4Lnqpk8YVcwaI
v8snybqIhGj8qah81rmT83X4kIdL/zlZp1asgZgjqkhf2yzkNAm2D8VFBxCTU7HtudCTBzZJ+L/C
EStEGQjBDTAGV2PGrq6H45JBLj55eGYiWqf+yEd8qaCEoPjCBf5LjmAarB+HoM7Y2nCkocwkd82V
y9r9w2vz0mgM+dsQBjYYtSzH0Qo5Yq7ff7y9kLjhImGFfTyOo3mkjH6309bVbe1sVBabU2+IiDDs
C6HaOSUuEfw42i/+pGJIsSLUd5FhL5zMaWdkeMfQgoKBlD0v7Mia3r3r9rwQFHV+5YfW/KrOkxBG
STXsK05vbSPFFVPW+uUVclGFAfBjZWtmX/KU0jgj15uFhg9sg0EPKltOJM+H/aqDfGJWn2ypUEoc
/biX5nDN7hCcFezwLxjmsy3Wg0v+ZQ+lMgdr66h2KbA6TNmXxaYDdeTVtO+6qadwMhx891QwySZs
OWSwClhcs8LolnLc7zUNhykIrQrlYQhoHQObUPq1bj9zeDPhLlc8YREZCdI2yO75dC2x+C7slCSg
20R6wv1lQDdCw9kjDEPGTs/HaWpwgcHqW0XIGZ3hgbBPAp1OB7JAo7VqmHtoVsxQCVyuI8t8YVTc
hnLrtexZf+n5j5tbxlq20LAGv8Cnc67CY+cYMYBpkt0sn9ZibJVS2vD82u80nG6IEswbQcKwI7nq
yvWA4J8LxH6Izua8GZ79OyjpTj22dkP2yItVmJlmloN85dzzDSaXF+rviKQeUKHVcWCHK3Se0pj0
CZsUvq4P53M8xx3MHfr7K7mT1f9o129/k3+XeDi3Tsjcnu9LbYOzvbylVkmZNYb6CwM3bGN3iykj
SO2QSiwxkGw2SLoVQIoR+96mqweU2wv+bi0vcPLWQr0GMVqcMTGKM5h62kWfDHnmG4m9sfMKEhmu
j9WSF6XhQPP1BnKwwV8PmmPbtG8+k35YpJfKKOaBOK0Fxixfykuz0KAuO+PDNlmwhLENs9Q82S5i
8V0685IHsvNo1niSGVCZ8l/cyEImNyIug+LDBXxVsjyf6/j9UhxjRuj9CP6MNljGt1eyPnQ4MqpM
ERK1lHpWinoh58aS45AWVj0CnnvNd5hu8/De38+oXFrNhMmna+RV1Xm3gU+jaljFiM0Wsk5TNQUC
FhY3XBc1XEcrU5dg4MD8RivnCIugtFML0Pohi0sIrWPSevyZonLylv8iO2DJ9j3NqPZYMd/OEgnb
KLI/yldmLzoninwM7wifyWQXt3wUCVJzfMwjwdLTQgi0yyd92l56zsjKqy/1nIqqNoNmljZprcEk
bmHw/UbwSZNGJiwHcetLywPcVtypO7wML7ZAR7271e9bOPo/jjWuQIqDY1ZI35ah5XSvotq/U2yX
jGq22NF2npS3k2iAGND3ScHJdCePYXMAVU7EuC/SaPvl2s1Sd7b7HzyT/TOOigeviO9e3JlJxHcQ
eckUoqohExBWiVay9YiwJEuzD3gYZNYdq/BaN1M77xLgB+jNHExyctgFztd9P3bgtZe/uXqIGNkN
rQBj7ljbJGip7JL0gT/aBD/JW99ubNGiQs7rc86UW88IPcD6Y8MFnGi0JTAEtYdul9GRfSuRZrSi
xTlo0sywJuxJyPke/Fop5Egg/L/pAJX+OFUqsJwtG3VRjUEzbgXx5Ep+poKJkMO4wfDuoUKgf9mY
S1kESevRxspcGHbGVyK5AZX/SIlDnP51eouuz1RWK7dKiCQpk0OTymneCxCgIqEoCcs2DchDq/9i
SnOU+qO6mBbRpfMLj8N8JuF402rci6ZY23OfzolF0mz0+hWoFLqFNrvc64qBwk8XeVSnZZzvRw8n
pTHW1n/E44XmmLsiTCbQgdh2+KBi9MLs61xdxTaEMBcaagddUmQ7QrzlXDsjlrg8z87ZbEsvEpop
LmLgr9pmWSg8IOwaJi9cTlfGKPpYCDhcUhwHHN853NPNYmJTIoKmkSvc4RzdmLDTqjQ6bkVNAH2r
IsWF64YY2cXmgyq0W8ddprkgRZwa0Gr9vU+qKzZkG1cafc8nqjWUY3I517XtNYw8SxpfSHUWS15u
S99wlF/+EwiSeeBI6lC1vAfp/M5SahLRVYAzEVYWThBI4iWCILVFLYkXGi25UazKe4UJtZvxYYrG
WbpybQJrhqS82NPjd17nSfT6CQDSblvIVeS4Ww/v9iSZSSwYED5gjYOzO6XdPjR/wGG2rfaCy7bK
XRZPl/JH7KPSyZPaUuEiuwxdPy9RwVCTZtkhbCJSyJzeGmPOsx7XfM15/gDUd5VGZZ06cHBw/4FU
w+t0J11DGNO7A4vDFPsIL4GRk7186XxR8RJTwP3wEqYZcPaX/LqDRXLGT+d+BBGWxSjiNkiW/YNQ
2Mym0WOT2Trch9Li9pg0zJOkD3J4WWbf8n/vPZmv7By3Y4qaQwR1/t3rgT41BUK5xqAaqk7UU2hZ
jryIZ5yGyDR6dvFkLgf7VbLkBMD9aQEsSGRztG+g6tKcdJiL+Ge8grPuyu9hru2fTPBf9dQIEK3c
/DljtVvPsQKiW7PvfFAuByERiBUO1xSjrNw4sG3fLy8jNt5cGCdk51y8R/NGG/3QeSoaYYhdCIfC
S6otAcyuxu5CjC1exwWobbPsYs113dy8Ts9NYEivPAl+zhHjI9vOD+kBz7v2IgqIZrPQwpelRZnv
jpkIJhmgjdRyvw9glilHO4tWXABx6zuG0eX+ojOT2hDziE4pGjdaE/Z/fnRMw0c5hWAE3PRlCHKD
Tz9KunkLf0mvFTqsjEyN9C6+dJefAY26HDczNMF2YfuknwiD1TopBcGOaOfhasp2rrNFjyAycKsP
us5rwE6avIQBy9rXzQfSW8pjfuWLFxofFWpCd0t3SeF5e9iG7h1m6okdtCSj2esIv9LFsjIkmepX
emMdur60m7LHIkwAepwSLDulkIdAP1cJouiGe/130MsdK05KrpKk2jVENAe3tdxVNc1IPXJ+VI00
uyClm4zigE/lsjccRdnb+NJ9cMzIEYmCj8CgoKbak5Lq1/OIV8b4t7N42IjiKQqvf9r4J8p9u2Ku
L+6feRuu8JYS8CgqkydhpFDP0VXeDG//sLdyJegqMKG03wApmjaE47D4n1g8Z6NnednXsgvuywfk
FRKuLmBOfnPxsBllmdz/3z2yySfDoxH0tMnmWeD3x9kYNusQljnacITR6v+w2+JVCT/D3rIkAf+d
1Awjq97Hm+Xut6w+EdICF9esTpeNt0Amhwr9i9rUPe08u0BWB7J5fLevardGThQwP4ZbVVQ8A16b
CaL7VP9SGgDSpFjKcwoknQVo+rEq8fTMidighJvyJDAnE9/96uG8uvgWGRmGx6OGg66bP57Di+KY
gO9WGiky0S5NXNkAPOIvXkvlDeGuFmmMNZ24RTGDhfsDhVvTMJ7GlbX8ujrLDwauCMCrrv5ZjxQR
r1rmDikPPx5MgLxbvOlDCaXuXI7jFR6a7zhHcLa7OE25elZFzpIaYOpHWpVY5EXMkK9CgMR78MRQ
bqubMhdPBsJ88ala0PzvJ5a9f4X6Eqs4vAC5A3HOH3KS6uQ3vhrp4+DIyy5uTgvtrmxh0hXj5EzW
AOR3DE1ZJ+iTV3OdBLbmhjymUtYP9IdhFV79DOV+dOCoF3KRN7L7hWRMkqgr6bP85B4J6GrNTo1o
pjifN97ZtPU+1Y1WP6XT7C1FIWYFTI2CIEWvcO8arceFfUNjdTS5mja7F/kOem3pqoEdV5nx46H6
le3tAfBvyV+wlSVlG3kfXkpOzgXGOcIJ1L1rcAMxTT0RHRepBF1pPHz0Lr+r92HiNU+rhEP7RwqM
gq/7WZIdMHTjmxssvIsjdrImvOW2KcEiyH9aSALIple1MJsLJUtfQH7YqzQEkgpcT7x99eNQwnuk
vSEJTneMzo2rgTpJBKBkTgqJYTdUvtoB8F9uExQajcYMAOsZwYMuYAaR5O7gw3DtiObtosDAKS0V
xkdeed2rMldZ0Wruooq7k8/EJ73AoeDQz1zhgSY13VqJ4JmIXEFIRxpGJfqpdjvQBkYQ6vzVlhYQ
MaCm0o5xCDTDnk1SwlQAFV3vZRF5NElE1DmKTKOxKCAIo0IIV6Z+LIWb2x/sz3sng/DG7L7Tm3qb
dxyTrCzBLeQCQPk5b99rYGN8H6bnah8bZFrQhrSLFD121h92tc3vGxt/iY7In1uv6WIyShNLonkg
xVCw5YAlt4AFzprkfVpTJ36I3biUCzAe87lvUnsoQl07DJofgSpVciOWReWGkj++JOeAFJJZc2XR
QbJ8hv8yU18AEZtRMlUKz9cMMnydPmzRph9pwRZkzO31c97vNFaiQ9kSiuYYyyLaYHwpxvJJWSDC
0FZJksKXaUom/fqbN6tn0687KXP5wn1dBtsf2n7vgQoRPbOJROWEO+iAEKFOhNBc44CTC7n9j5yj
Y7yPIwSwg98asm4NJ1kUJLqPFMuGK2LdNeQe/DH+w6hFVFRZkUT/9sJEzn498p5mcfmJssMcGL8j
htWmh/Xg3fBRT2ydQsVL6K9MuPibVAfz2KYF5cGLbyNQMPB+Y4pOzfzR49ZH8yndLJcgmeubs60e
h47FpmHBY7kP4T5hGoGwvaEjbBRSQIqti1SbrTM0DYY76TPFyjw8w8TMWlz0Wy1WTOTOgrUL57eW
yAtKq43HkqlLDt27NaV+U9gwqs0unJd22go9gUUldfMNOqFJqunWSTEdaGSyGc0LOIkLwNyVhLR4
mgWUqz8EoFvhFNa4Hj+zBXKRm+XyBUMFTGggkmKntg6CpZe2CyBOj72QctVSJdIaOzTreBJtu9Ny
j+TqiwMwkgqEZU+XzLljRsrQ9xfxm617VfRTZ/dL2i1P4E8fXQvGRR1H/xyH8VTocKMmlaWJFgdU
GfqhX6aCuxjuv6qDwuQLIGk7UU3SYRK+pQdcdrxnSDmR6OPVxw7pSkdGffx2iD08KmG4SNfBYhGE
h5ohxpacyRC/5syHgeh6/W4ACDp4ikxLYfHKjINUBAnssgv/NA8roTjYGVfToDMoqtZgIksWOGqB
xWJJt49JclpTrKMZHy0b49WqQJ7//WdHClWi33SU8pdwFMm6yHfUFHTZ3z4MrZ8Zp6BtzdLEDVOL
WEN3j+5rbfrdPggQZvDqgojnoa2AMDj+pTyj7H1zdYR0EfxAbyyim+B8q7Slu9rS3iEELMW7ET+Q
Gq2pNEgYcLk5HoDS2FPG9FZsoJsllq/i9roAWUeA6RTTiRbeIkc61bbHe9SOB8G+CWSo+Yb7jlCS
Xq1O2cIdf2u5FtG3EByMsczXJDhcGmaVjTao2U+eWwkp+7ZAPXBJezDhxYbK6aO8HEwNuM1ys6H+
vdPGq6LoMsS/Ty3g9bM7GUC+BS/7+nPviiZRcyqt5D4bs+M3WiWWC+GEPw9wXPNXmgPkZiIzpy3Y
61VTBoEgjXYjeUI6BpqtKaodpsGUg+wkT5mUyGdBJL77XAuASbJipMSw1+69rgr5SuBqPlVbIzQQ
VybXUmlsnqEy8suzCoDJAqWnK4xI1RNp0qLFBE++PRcRf/S6FmxElZCIJOfiLy8YrD9q/jVcN2UO
xfJWOuKQsY2VtlJqlVDUyKfp95DU1rYWKlkOI1lb81tsudIYzMKaLh6YbH/HFunqmHpM/E5l1QlR
3xx3Dd5sqwMy46FirmVDv87GeVY5BR1YBkZHvvszhvHrp5fstbLRt7zZl0ZgSK1HK1D7l8IOsraT
lef/n03CN1mNCHHpcTjoqyLO54lGoPQhcV9f6AXlejJU3h0lqLaQzAKoPuEzLLaty3gep3H2fZ22
ZjdPjiRvpI/KNGA+gxXXQiZi2MKY0EFIR8aP5mIqWkKC0Jk6WRH9u9mhNhXsDDK/9oOrHN2Cn7uS
Mr4OoIMi/woemxUKgz3mCtkRgcO5uOFRzCnROF21ZjyioSWgI0/6378zvWlHRLfVNpIwkkY4E+bN
NnnvDH5K49P9HFUOgoflEk8UUCmz/OWtxdoNUJ0GoMJpBCgxqyVqZxlWMCLPpNIkuIHLioQaclZr
Wg5oEj6zcRHn00bIFHg6GRg8DcRvl/M8i9i/JbfFJtqRNs+r3o3FJDi8Hc1lQgs/wUrHUs4qNPZS
s+hbgZX+MSC3DxuKcNzy4+qbNQhJOTNdFSQJet2nr1j30exB5t6FRG5HOic6LDCj9VQ7+Lxrf6Af
62k4Nw4IaUxR3mcbrjRby0DcyczUkPsVbIGeldH04SMYMvpOFE+EQNorTOt3OG7xuZcezvHKqDg6
LtZiTHfHspqkZ2CEWG+kdUi/oGJ66z7f/OBkyOnENKt/++UIya8jo2TZZaeTeMFC6DnbV8sV5e5s
UKssvDL/g8ekJLNtSZIzIyAwaKFfsMJfmn+XIPSRYCUonirUQZTBp4zNUzYNr+p/TrYpNot8Pzmn
3m/x4OL17xOYz5zL3DZw+87lkOjKhBrvFfhoR6IhVLZ+e/c6LiXUBfsBjDNYUuGQqvKYE4LXC6y5
vc0RAV1JLuttUNoolTpialq9fkWYE+YJzmneOIbhNSJYc+eUip87x+wfaaMnOSvvVg2WvgEp4UyK
JwBgeIwaV9qytikVd2pZyKEO+vzAqzkU/BxRw65596dKpotC9M3Ab+LCtNUOBTw71jvPFWMUCvag
ULKRB4Oap4XMwhNi7X0rmyNkO31r4ISV0ywc+fT8cdz73QFbAyaPft+Q+vIdipLwmyB3KhuFjj+m
uHkaS+mPic6VGa2FmRv4aUrHZ8DPAZXIadhctBYIvEeDV6/PwJD7ig2tbCpVN2cbKeYjQYphZK4C
TudAj4/9b09EC2Lbdi5gABmjpR4v7y1f+R9nr/mOijheWzfiJPoBdVBzT5wjCpPkWHmImWLcaVDn
m10noAQH3E6YAUOTlvigGVGRuNmTexvVPPDJm8thxfBrf+iPRFayxOH5glnKM/lWIfir5GbgUBuw
tGKBJhxq4vjmK4uNrq//508QxUXTYYmuXwh/wZngznVxjlS8382/eLt2xVUbTKmuNb5U2/Xp+5cK
B0n59XFuq0IFI5/BhR72sB/ai9BAaSfyakMC7OAXJaDA1TAfbbIYcFW7gq4Knje5rtwKWhymWakt
Z75q3cgh3hlb9o9/9g0AOvO2cxl79wSU8HUPt47/CDtrUss5nJRDRROcXslfOMamYP0WssPGKiFG
Ad/bN7jkWqwdPcyHDdZIiAlLBCvnpN4tpVbmtFrQDPifr30G5pnlKZAYKvtqjh4aBR02zu7/NIXi
Mfk7GBV7kWRB6LrctM59/N11qP/Xnc3EcVYUThuUb6tus8keeZhCYBfzHZecdDwlRiKa9elTdBeA
Co+FROktrqTL21Gxp1a0dL+0VSFEv9hTNOPFW6W0mapjE2qqNCeyt3pNaTwdG/7nWK/5/5FYbhSp
tNN5SPyqA2V/B+qZcCSqSgt2mQa5fqg6jgiey0tO5K1v3NRUYSSlT4C/BFWOjf8722eK6hPxpluX
ocGdNQ1xJXUL/BOpxYdqHyUG/HZqhekG/cpuQy0Z8eHVTxu7blE+LMMQ1yB4ilkniXxMJgnZXV5g
mCsohleRI7YxUAYxlQQ4uukbuGZlgBkh4DTAaWXt1XZk924refJwzSdgkHka3tXWs+O+ddfZ1oA9
3SNdGCIfXbY0rZeeqQazEyuPd1hxs3fLYzURq5VU4pBn7POIL6fa2U7LDlOlcTjLcYAa0VW5RcHV
ABsOE52Bs+frOLlajavd6pN8lNaM8+0Lyd2sSPENHgWhMnD6QqaCwgCnbW1TYDkjTx9wCTHyii7G
5MsPWedZADruJaoi2KaMbm+EPZUMBpZyfQ58AVcDeGw6+geIa7pkzmkaecBJxJe/2i4ihB07kufF
RruiXRjgSNKyU2v6XFEdFY+xp0tYHmPI5J0tdSF59aOCXxUByoFu3/O4dl0Nj630TZp5gqTQJAr1
cbxY1W5o9yg1qHM+W4LMQn/1ryhYNUVFC0iHsfwmibnrCkQhw6dGilIKqH8hraasY7hEvgMoFnRY
jX4WkecL2lyfWBwxPATqk7oY/RCiSbaDtOufScyicr4t+aXZCj+EIjpCsVulM9yZGh2CkFEwzHfl
0Q3ckl5NZxAj9LvcfNNcAfhFWXjQTvBcwn7aGmmj2j8tzuNG04K3TNdqyk00ZVH+aaATIL78yDA0
1cWx3em3hEygXh9ueeWmc/wHoh6QSaG+AqGfJT5axxgfmwVYTo2sxuocz9OdBYH0j4/aJCkbSbkv
eEB1Fr0RWyy40VRv4U8X+Y/fDjyXzK54FriBqgs91pDo1ubdqWSPHHFOd8basSfITE53QnsAkdOh
a4WLgG1+KbCaczlz0dN5RW9njFKtaXcwbe9gUZJpBDer1Oh9HFOFJ6CH2VP+iLDWV9LeiN9e9l8h
x3ZnPoc6NCIZ+pLR8e9wgExPYpgub9UdrQPyMy+R+8diFC1I2Ylpcpn3ovowKgtHFRscc7LyGkuk
2ElUvoBg4nDkt16YEiVqPqT5ZyMJII60BbCM+Cx6a62cdVBlTkxXYPOoN9+/wS0ADEhz1p8jaYDa
aDtetfp2DLdL1l4r5MzOUumbiEiXlox9W+4cKfht9pO6xnaHbyvDRn1ITajsNapEp04Gcvc/hiK7
KbT+YUunqbBp9fCiIQPZbZE7rjQBFXwAlSrTPewYUvQcbJeeTuXSCcnHBB6PYUGbFRNQva7Evs/9
fYZDXyUY/EJxAEjfpx5V7CSb+e16k0j1MWeWJIDHJaPFimKxh4cLo99My1//rcuARLGrMP5xfEu0
MNan8753uQkFzpFVaF5PdsiNXT3XkA3lsH5r3yG2wx+b17qUVmweYHrOYX2JUbnZH5qcmXCd3C0/
PqUUUCsmiYzB4t57BhT3xAHicHINxaHDObEZPp0AkD9OLOTDwdHNPLCO/C7IU63S6IlWRvUWpLLz
9GU/SuLEzLrxQnEMNEFgrWBTA03XADKGPITlazj8WeDipl54LwrJLob89J3/vrRIxjl59y99l77M
mMyZ1im4aneGDTQ9LNfMKnP3Yg49IotuyCesO33trGakflEZfbYqCcVLRxuzf4r17Vad3tf8amyk
mbDN8GDdacs5wZ2/Nl444nysfRoUPcywfN+NUlxTlnbxbel1gIwWpu3ckd1006UtkkM6plITfSWa
d+BE6jOQEg/p8Ug82zBpgU7OoD1KjjpUOtqlk3r0/k2xLxRtCQLk9xOAvDKaaO52E2C+I+uar+Q+
Ak2JPHwl8dgAkJofHlMDO4tzKdA6WMWiXCHRpw4KKNx0mbzS0rVepvr2amAaYMxh3t2rAftVnBcE
hof6K4n9T4ZDbBSXgLWt2kcSvag0XCFJGdSBVcJMThiIyTtuyn3QstU92LHOOK0EhljORkP+5wWX
9VoNm9Ho7A1e6pcT6KLATc7QfVbp0EbE0tZtORt5A0MJ0zT6uuVijgDUGlSFV90czwhZj9y0lb8O
4QXtzjlnSPVOO76QlqRFB0ppeaxX6CgbCapu7MBrzszm8r1+pQJqIYeKr1Q1IHUcxm1j2DIPMKhg
QTSeVsiOOLXCS5nhXFH1ZpjFwy4sVUrL6mUsx49MIAPl/ZB1gLXkK1Xz8PwjdQJeHe4v7TB9nU7c
wJi+VufB8l2Kvp86UGimtzJn755DLLfuYbQFf5llkEOLQLJzSRMY4vvlz9WMi6lMeHyX/Xpha7RB
w+S5G3T1G8GU5Jtvt4pweKWElBKgHe49edh2d21d27YHDdkzg4ND3+sZrC/qyh67T2nSa2DZi3ZL
oxgrP+jbn4FE4Brt8UeJgCqsQuU7Hzms+gId2F5qtib6/SJJ1spD0IreHUS3+iDNlpHNgRJ8kqC2
7vX6Q8+vie7fM2xMfFBngwE5fQPoL80s9l7ONOp01iddjfN7aD/dJntpqprfdJHwUYHiLzJI18Yy
UZ8xgjJvjUppMlNihen+rWcqybxwdtM3mOlxARLocGNyQyWG0aoyj+R3h7mJDPojhCBJZShym9QY
K0DpQrtCNzUBR1IO+AbX3PX792hNUXUAT0wOjG7bjflI1KQAdL1tw1XFrwHgo1yccZOXw4PeOKaU
y5rG1/l1EMLycvHVPeVLOekUOxnYZXn60Kz/51tL7PpZbW0EhVA2pt4pm7oatfgkncOmleP/Gi13
8VzBdOHj/TzC0sb9UgYw/wvvDpehvlYWKdWFN/KbTwUrbcMV5PByAgneOcLdIBa8+921YkA7CmAN
eN4PQb10h3Hm0xZm0ohvK94MGG0O//TzIDsKQGwVGO3ny7TLN1iHSznFK2OHUVqARzKXqEXXUpcw
bMoxTpv9xri1fsX609FUU6uCEfo8HwP5lZ/keyCyNPe2Z943mXF3CRADeH4sLY3SRhXTPHe2wpLf
++a3MrmNUqwBL7wM9yrN5w2PAVf+SicuygD4x31sIE1FDR7wdjbLdk/rozZreR1nX/YQN8fbDfvP
2lXsiBZbkclLmj7EkiVduWw+oAoS0vt7G8x2qzK3AdtVwDnZvefS83CdRfyaQujYcKNu+FTcxxzH
zcIQ84RhRAP9m53YB1zsJI2TpSHGuH1bAHX5Q7ayIUn+cHskuVBVx0eGtne0nQoIZSXU2hp+VUUF
AIEPssDmkfukCZJGW7YR3qqZU8uSB8hh7GiR7F/D4zJfLx7nRqyxhn66sC5O2y1T764bNRrVlXmZ
F37Rrs2X87Tx7otVxect4wNAD1sNOA6lYPOD59sWZFBcOOaV/K1Jt+dcUK0+eQxAQTt1F58WpndE
KXfdsXr7F9K4SZsP2DX7UHdBKVJ8yFx/5NrlsXvbjjSKt2ATGO9RpcSdVWUBS5Ek5pAioi2PBR35
1ugE99hKq6xlu5+09AA1FhMc1KsrR8F37dONtBWmZR02eBVY3ELBTbU2zJpifQjVGEs5Bhvi3QZZ
sTLX4XmQ4PwQrOrCZH/HrWbQzOj+ymNHoc90gSFK4bjz6TThWSFfZkijM159ybLcgaOGnPSZpSXj
f+E7pjrboyyhzHRTrinAOLmGroGb0WItAvZSE5ycaRBI8s3gZAO2yRu1fgmiNlnYET9w7EP3Mlju
Qwa4lV5ZGPAJS0NeiFFvaj+zLH1Fg7WQjBt3wb69Ncq0qak78AQa2UV3odTa8mCxuy/Sm9xl3JVJ
d5Vzf78KTqLvrOyPzYtO/V4pHZzN2xtX/ab3hDfOVaGRIzb5S+6EoDjlKd4gRMT4e/RHufbr7UgH
B9TZtjvvjabsYnc6cjieRoknOTo47PNyn9u5YWSE7HoZgeVdJcR6pevfWbITh1/VKX4sWbMKm4XZ
5a8JPYipqmCKSFS8mJ7+ePO087ruIewzXOMIQFUS2EP6XqT9cIkcCmiIS2LECnfkVAXK8eSlUJ9/
ZW7Qko7y+qcS5iXRLSLAP4jX7eMq94Jzp4M7sOtaskoA2yYxSsrPXHo7nbThoUv79wBChtVb6Joy
tZ5snDySMKYJVLx+t1FK9A2yi9iomLph/ls67REVkbXWvI2JES1sw3U0B+bib2cFvKjwvOBh3Jzp
xNFjloGJkFYGl05dtFEqFu09vIx0NO47ey7vKqSiJ6erny5CWVaJ3rdJHue6DgqQcGbtE3UGmZsL
wkmcHCNVrPN4gtNYagtc7T0Rqm6AlIMOuFGhJe5sx4r3ZVo47nEMymCYa5YkoFk6DZrnVjJvGb4v
TTDbqYqXck232t/e6qotzjMc5PdgS3ifsQTV2+NrvNlnvNV92+Y5WVSMnqlnLJPa0F39KwBnGkm7
MH1/pJ7+5WkMc4Sjx4DJK1HJhgxQfu6obK9n/Kqmt/ISPlCii7eXSxpajDfK2i0kIT0ojRqCQrTO
Y8/cEj66A1HoSVt2VSlTWPXV6xbqzT5/S8LPUH8x00uxt1M6amtSivihS/0XIBuVof8XVFiGhsGp
GpATNWFqCGjO9Tw1+aC3kATYQ5osdyr/XnVK5AVIrTT0t2OWOhHUGG/gb2sQzMhoKwrtEQaSerh8
qWiqw3WwGozsWt54x0RpeIO9Jq4jx4+fS95PT63D7oRK9z93wp6qvKUP/3zBGDEoLtYh7caJAQOa
T8VpJTyyplHcfq2oHvX8gn5U65oWFM2hdENsWLRLNT9q1ZHqbFx0wVAtgwXtARD/k4QLfHcJsAFu
upOzcWC8bCM9MsBY7gxU0Jrq7K1tr31sLz7gZxFWKQZ+kMHi+KTBuTfZcYQX7MlIAcG6qRkFrqda
wLpuBm5BwOaDatbvbdvX27hmTv+us0mwAQhgjyUI5KXDDcZV4wlCw20UKkVx6S2mV4LARdPBFe1E
5PfmgFuZALI9eTIr93KbuUOWNznqUvURu+pwRT0bzOqSdVacUZsNE+2zMgV21rrUqKg0813ttvSZ
EYePBUlWXkL7NcWd1XFNjCYys+bvDLuamEhgch8iCuttvR8ABHo1AmgBfSYOPeRuxlS9ExmG72t0
oMkytRvPGuy+qTA7Q+Jl9rzJ48SgdVoNXiFNzbJoAGiTZQADHDT9c5BE7x7ePDSe0k5a8cRnNNol
BkXuOjv4O88h+d2M1dgolmSb+cMOfmjTSW8wpjkeJ84HNReATW8igdcs7hrsSwijlcezf+3tT03K
AwG1uINUmIh64OW/MihLlghqqsGd2apRWOdJo0UZaGWlUmmCdT2/3229RzJGxlFOeSrgQQNqoqle
6CNettA+xj9Mgz+pX0dm1/vj6GZpBr9A98Zhq3Gj359nNKr5KNlyeRS/oCUY7L73cOjFJUnz6BGY
0SWrZwUnsEQ1LOCesaoE6BQOkepqVe/SrXoLexj4PLumESMMGs9ed5WXlk4uQyFSsx/K78PGF/Es
yyIZxn9UcaVfdCk0JgyLG0vlTSQmUTe2bUOEVSAWlF9VpAaReKI28aJLzMfwyndrKQxYJKk4pxvA
aJRELsO5CHoHRotY7/STtPEOowliYLNinj6qjdtlD9yyt9iOEAkhYoNKUcnapHDbFVjP/7TDC7iU
dH2e8DHUQtC/ad+JAWK1/NainMjeqif8eAAxIfQrev5haN/dqNOqYPYhYaEqdwqmQ1TJgFlr7lsT
yGv68gD87MN6HN8mSaWKeCGf+nRL2XLVxTM3tohsqbOZdEgzrq0t3UtkhxQhI+s2kGleVzWQ2n9q
D/CcIGBtb4KAMCD1jwI/Rw0TSJz357TKBbL53OrAOWifDS9vNQ+y68B0cotPWQymLvFg4s/DivM6
6iy5VF7ZgwqFhvLWOfh46rbxa8Y9XdLa0cvmW9fZjmF9j/YNYEHn/42gqXstyh5kwwiJuAyxtBmp
2edd10DyOg/ZGVvVG+lzq2fH2+3HYeQLO3Mb75evLivlCuunVu+b75eL+hB5kv58jbclbO29/c9B
Mh3PBGY+m/HHnXFwb9BIAx5pDZE4UuXNTGmpbOTzwTsPf2xxdLMi/EjFlBdnR/ATiGBOdPhq/IWs
tIELKFsCREyRU73fCabxmkx19RxPN4SnM7+fBdbE3cybBEcOstJOgYd5lxjwiq+cBAnb24rRHhY8
ibpXaj4Y1CZhsqgK4J2DSvDTehtoqolFBugfAVq7CZqx4nIymscsm4/OrIQdHHNVlyUaVydsENJM
2F+Z8WHY3r4rJyDoMprh6eZmDKVg/R5HU7G97Y3aO4+DfVk2KhWI2kt0zmyDcdVhAYFmQtFkUkuq
I38zA64ud2NvXkktxB7gMEmZMDU0rKMgswcj2znK2U9EAZjP48NhXxIHo4yWytQEkcDkN5WaTlk4
rZ1USfON30VmZ6W0yaIOgSObOTMlBD3rMXznebmaH0ZwkN4DcY/Y7N+m9isQvDwBNoQs7jKw8tHW
KKXykarsv5tyuTEgMsrs12gW638SsX4XFfl1A0XxQkm7iyCRQAzgg0KapojD7poNdu2JHgDAe+lI
m80brxz1IB++XHprfS3yv4FDwNEICujTPTVILMxIuaw3LqzE1ETlh7HIBVLMB7jnFvB1z1KUxA1O
/967QQ4Zu8UzaSBq1XO5PnlIrjaS+GPuoHUEFRtvFcQkU+DQj2VnCNBY+VviZrf/W9Uz3UiH6Ns9
gnjJ9hEaqwxrZEy96VYPrC33AOynv57ZxJCwVvqQ/UQjiaqBOvFHqgRWUs1J1yYTESw3Zbj+hGHl
Uou8CMagAEmAc2ebtWd3Fi05qBoI1ftBbQ3qmbB77cZxzbv4cSYN4i1pvtuOw5jg68Ja93a9RU/I
TscdpEulPfAjNU7U2wH79RiPqIsGJezPM2etha0u6EAgQ/Xn9FAYgb8um0LZnZUDB9F+dDxO+SPD
WT1QB63oFX8+pAqBrrVtsusOkOFG+2R9otWCHWVdB+/LoVeW4wCIW35TUP02jjIZBATchkpgPiTk
njDcxRgsuzUK3MbcWwdF6cY3tFIaZ/8mKzlJLVQgmSG/VjSxYD58fTLCiMGjsYbdb+k3EJhm/cQ6
kCnhcWr+xh+nVcHN42sloqi3cvduZEeH35OmC/aLWIDNlFNPLnNBDg5NEwbcTdLhlx0uD0mvj1pf
l4WAlBCKrJfDI542MnMUkcnQ8QwUcScPuArwGJsAV4kU7cKdIbveYFzBnQ/l1TapQRczJa8PlawA
IxY6HbyLE+a6fld7hdej5FPaOSidY12XEC2fJConLyDTpnx+s0MboIDTSy1PDBuaa9p/9oo4k5SB
txL1B+sL8K6jc52i0j3IqfeZxKLb7W78hM3XQENtpSWagNGYmsNttn8Ap4hxANZaGijCtRjV6lNn
wc4Tv9kEHCTbozV9NJtktBDIsRAiHBuhNXqO95vfdgsj4dC8b7X44+SH98MX8YXfSkPSIbvj3LbD
nZ7qweVqpjV/7NMUJuBgrfQCY6G1l+QRf9vhj9Pl4t8QEJ0kGFri117LqP1h9OsvKqQDE8S+145q
88WsyH3vMTkQU+vBNOrzwZWAJpLm2i5wA45CEQwgfc6miS9Wnw2rMgIpn2BmBdWnsPGua/8IxuM9
k2MZc+pER8ExcxsNQEo5ke5hGSo4IRR1y03Hmlwu2WvwDyWm6Bm+219Yi3FNugbmoYKWqTbmHQLM
ZF+ORsfNVXPz8f/TSZXErXvawGRzX8E+I8SZcuIpuOOQJwrzi0idr6o2YTvClZpmS047eXZ2VSYR
nIR+hXZomqOJqRZr2x2aBYbuAZtCHbZRkBELyW6kY5m0Qcjmxejus/WfY7GQS+h6j3/4XSCYJRlh
Ml/Pi26Sm4jnQYYl0y0ahybZXXPsUIZnZcNEBYghQmvZl2QWLCBD+lG20c9VscQLZHJ10E6kO9Zf
Ss01bAsXbSmDL3mKUy7uAeag0sAyHouZHpf8vdcM32z71djuSlhs+mV+OtLwGzKSF3uoFqBVrcIH
5ov+mkZxRrdRUwifJujddtiPSMOKzthrh/x21cTfHkIIYoJie5RFrzoxqq0Ekh85zNIsoNNZyFjG
ab4LD6EsNWwRc0v0YJ2sYv144L687j3CVxF5zJgZ8Ysiy+Dpbp/ub16vfnMv/EJ2u/2oxwxC/iiD
mdsK/4zNPVOS092cXX5DX0Mg6JF/KvzMmrWmEJpMRVGEVM6GFQK18IwrBTbpaP5yDQsrx8gZDpew
jD+FULKEv1bAv9HMmBjCssLV1V542bX4qB8hRAo4P+QRxepBdLKSAOhRlH40ylMBoSQv4XgCaT2M
MVL9E/hI1i8mFYBFT6J6PSBwVs76w7YU+MulJcqIOHMh3AhPNxDRU12C7q1L41NGf8dWDa63q+hG
jE68qyjp7/tvuq/sUtys8H2WqenWNIt1Z86vj5SH4KZsBdiqGWUWNGs7L/pl71akWzp9LNtKxDPE
I6ewuB/1YNKZP3V2l2pM2dFQ0/4S4vGx2l+TkAMat2+DXP9HYizrF1PupFh4VF5m0K/fVIGoiLq9
JDii4fKHJk9TwGZZwHtQ0kZrtCpmAEQAnQpJOxc7LdpgSHjMpYA7lR3m7dxMyjwVzIvLWfn3+IA5
LInDXuCQZr6ZHTiCZ6wzcJ0ViQf+sWplO4lQo97WAkuFo6JL1WGAhZdiiOIAb3hR/f1+vr367ofk
baOHsxj7PUcEpHRtyyi5H0aiuGdrTtKYmW9umGyHb+54dW/SWvpkz6L1NbQ756CFhst7WeDWLXND
4kOUWDoNHoBztxu87UOJ2HNykYx3QOdx8fq6AYuXcpTtbBSMnPm/5jELNQMswUz2IPRBouhnXHO2
MdSA//IAHUUDcW2Eh86ONOFGkcXSpK+Buj9ZEjvGtb0IzYNHKzjg951epzv8avKLp3Oyy+SarXs/
Ebmt0VtJvmLBTq4ZLUbSwIkDlAynLcRDSdygQgh1df0WZ79Hrfly2ozuDLal6QeJyRI5h5eIqJWf
6XPrfR9VCogyRqzPFa88F+db3K78CWAQmCECgt8kzThbl16dR9dUyUcU82ONr266ssoMubsHrbSb
1kizk82R9YhW1plVVCXwdNZv5rBd00B744CAVbcjZSEjTOEORv+6i9Hj9pHf5aBmE+jfjuqlcN5F
P7IEX9PBKmU1PkMboAVko6cnGs4b9Q1+7gqgvoNqsve0WbWngSMQttVMGoBkz7MkMm1yIb38lvlY
LXqvFpyjvYRoXe998Tbjjwf7P8dF3ZmhxLWDb14/6dRlU9/An59thaHwC7PV5H5AmKrb8SVQjAiR
i4lsOFBZ9tXCF801BsDNB6UlLomKXl5h2Rp+v3icb1ruVpfDXXoHvDZpfSF0r9MFUoArWagIgeJZ
ORjnjSx9heUFZMjeAbYitZRzlw6VURCjrT5OpTkn9Srf6xTIIES3NEsxeJgY2iFG4ItMCnRfbSB4
fAWaq5cMdAtdB2cVwqOBPcwxqsmrpeZFa/k8KedHquYUcYAD1AEZ7pF7g9qutuVGjHgZt6tWxJPs
R4AYT6QzrDW/ciewhppO1vpCsm+SjiS6GCEmVPxEMbK1O7v4D+AsihzSHmKLC+AbdFBZfdjvQX9/
+yfr1XQaZnE6our1WMASM1J3cmAaYjBJfLeydqNwgMi2zUYulosLf7v4Xtw45rX5lwvRQFaDqSv1
m8kwKkn3JEC+aFlsz0rIm6jIAXkxCIe8WtwZOxkws1NyQBEHaL+JlMJaOpRoi+0EinmbZcbtLi2f
vmfVQ4fR4zyNw1Jr7iLnFGSy6Se1c7ioYKr1ZYMvCU0wTccmlE1txrYiHwVzNcc0vtwqW9MJORq2
OuaOzBCUJ4InIQ6L0WP6NJSW7Q8Olg2f+y17b4xgNvjn2aQ2v4PJrYDzizQ7ZeX8GjWlJoswP5Dy
m9ddPOb6+i6JdSYcT+rwFw3rXMK4hSJNiG+RFNumZt0bDjkn12lA/v0ZpFHFY6nHLppq8MP6CCmb
bvdY+YsgfxuTqqB/ALyiybekbtbH0L5uKCutkGGGt7tPNAgfJ1R7Y0g8vrIpXpZACEg8qE3eCned
Frm/f90dR+c4IhL0jnPGX02Rr2orDVa1esV4pFLpBnmZECUZNmKiYqYJU+w3XE8yBx7ExfjjB7jH
imrjLUCayXS3mKcz411vGyzPkJAYUO5/adOWh8/0diSZpbFEdst6Z+o3dbZCe1a0lXpBZYQU8rZF
6UVasdQ06u4rAZg1vHUgDCzhdc0DrO3nqaBohdg3c4R+yoOn08EkBBfHR4J8j2wAujUfQQ2tOE6p
l8uXIrUKmw5DBtEOoJlXoXf4APf+9gsz/rlOdqsr4Z41FyGk9FDx1VfM/tLQ6+vzV2IUxbUjgqSS
p034WrtD2k14SLH+f2zFnbDHP/XgqsHnvHAmYgLUdDs9qi4hAzFUVuugDGKz9PYX3VSJT4pdwnxL
seeNiejoM5BeKWMmvbCsGkYhpzGLBb2lbRYRHRmdVQnacrZtUc2XyUj1hxnCV+XuzJTRTGoYqU1t
FxQ2CMYz2+JrEUnwUuAWZMS4FxaayWMiwcFv8bvfk8Z7muAPnWZGCUs+e7iVdKyFgZmM6eYpYBxv
+846i8jKUdI1MDJhgFXXZuWA1uRTkTzTnyV1IQ6/kPkUL1SthXmIvBz2vDeWoAVVAo+XugRyd6to
LnzWd/49n0M3N0WU1Z05mUbpmFn/uSGrvBeoSdZnW52e2L7eAQpGYzqNiVDJettw6sNGym9kYhVg
69xZAbx9T/jFOWl1OF2TH4tkMNsf/TqqyEpNk7NEo3oiKlPp+S6TKyPbEl112tKMKGIu6vl2uFkS
oJxMVM0oWfv7RnjFHDPpSwsVX2wee25tgobGHVxII07Dd+nFUjvBPCpkcQXjtMy3opiKm0Z5tAyE
AJctOYoRor/J5/+Mc9VVgz5N8PpdrrHtOPlZlkWryOHtcNYrYpeThkOhaI04IgPyVFc01dAvaoth
oXqGr+5r9qcUWsmIUk5BtOy7Hh8QgNg+jpLK4xOGs6RjxB8X/iAZ85Jd/vPEggkOpwDhz3K7YVWd
UlmOM2UA9XEyaywHR+zwUd49mdcrbWcw+Afatoc5NQsQ8y5dIU5Qb6ItfRhvDnQ66YswDyc5ADDj
NgeKPQZuWo51oFwtA9Xjdj/EHEk15qpQXpwhZa5sz6ZAaX1mw7BeFJntiQMCzQmaNA8gPdWnG1Cu
3KkABdCHeRhu+bTqG/8v5jiJFIqjB1ZR4hSU+/ofDDez98KWLWnalZs0t2pmkxyCtUXCcZE1MzeR
oLDX8mKWszByfZxwAMHAmuqiu67ICk92p2cWwzE9qqcEoW9VNmh4TExszoyQ9Fm5Xc5oOoW7K73x
eC7dqLUN7B13bSq0cRrKd+5eBb7GNe8kjxklOrUyOaPs7hukRcgPVZMzbxH2fU8bdBBD3MfipXf9
FWag5fFuPqTO+0trBRG0H88I/bI2QIJPlD9uepcROuLA9nldlvl2an/levmym4lEmyI7sEW+KbpJ
dBG7IURE+xI5x8BBDq6//RK6UNsTHA75CagV9Q7LwC/p3EkDdKynRzrni21bxeTW3Tiv6gq6i0OC
bTqtnrWY5zd8BLuJWQZ8B6yWYtcJrcQOc+Td4QdNB/fNMy+Jkjo1FOeBkyEMaGSqvyLM/tScrmP6
hjO9mCGAODQUGTF9A/nwR5rUMwrMs5kJBz3lGwiVsoiQg3RRs2diK+r/PDZKEXAvJAm8cBqITqE4
Fn4J1qKC6EHoDHCRa8JLuBiLixJB0cOHsfDCzrbhYCxaRMfsB7kFMlvwkLa9YricBQWiOdXwQRtJ
jgYbXi9h98cH+iUFWw8VeK0WQYGpfw6VIBtE9J4qAaRMgeV1XhL7zIvl7FHatleiaIxyJxvfgqKz
mKsBsc7MYbvFEKOZfbqN7BcfFsDJcQ3RhngKWWIsoyVeG9eWt7R0Uug+0A8wNpHsAAXW2Xx2pylL
FibvvHmaHr3J+jbWTBLumeM8qTTLoIb1YPVjcsFtsrYXBhIySyjSWOgFXGSrX9tRQSvS+qXmE9tK
syxb32Je+xzVMUDDVIyVlj8GeyxObRqU4UdYxMC8mYxEf7LWeUvg5PdmezIUrOHFBssooRtAJUTC
/ucZPIA4JydYpq21z205cJ073nBNT2z4wVLOp//dm58V+S5gBjBDzh32J4opvmaLQLlbZ2fk7Sz2
AYRF0oui+wN0Lnv17WW7wNdcy06+sGP5pazRnzNp5CG+6k2O8x3w9JrktN3R/b45s+3F74swxNSs
hnXlAcsLFpYKJD9ouhAXhnAHZmsj1jNF0PqCrdcTe2d1iFV73cHRP5znX1lGoTsmNOrtgv4DjxnO
Py6203xoQNBwY8MaY0Xx5RcLq9KF3ZOUI1oR9idAoAojRZz2HG1gPl47d6GhZ/fappG4Paeg+bor
IV9zgvWy/XksSExmMzqt7fEBxAVBnhq0sIXAWD4N59V+lHJcu0mjMqgNPiGJnRVDGPdFML/g5J0Z
amVWDZ5bYo0y6VvDfGPHcgrozhUdZ+MuL/lkjIYcmCGcF7FW3a4ZzwCLz6FoxUaGI/0l6hk1cb48
OBF0xhxG+NVOWDYuSpaQYlskgBd1Fhi+2Xbn00ePoTe40DfCEjEnEVhmdTYGSbRx3K5S6t4lUG3L
64lPXYr4ZLAyzFJh+dADq3zaKfwlSJd/znpmUO53FdYvdYhwcKo18bLuRpxeqyGyT7LFHtJkW1DC
KHqz4qYv5CN5GlSE9AeqDp0JVwhn56qolqBN+FFdSJHdEeam//DjaaXfh4gQe6Qn6PtQ3GapFdKN
Tqma1nBfACL6wexCpmkgcbRJQe2wep7uHxqU0+3mmXcCndM+TIvVbjxuYC1azOn9OCPzdI29TPdz
4H8C7rNP75N0ZTmegF1gM1VOwoq65pTLAVrJN3VEDLWlH1C6cY0O3o5a6FPatomugFqa4WXxQIlK
DTFj7IVn2uJKR/8Wg4IE0BriUW/GuTjFUt3eV+dxqM8VM5nXQs/pvcYFd3EdCQ2MJNHuGBUzNHlA
mssUxDvzOIL40lvPIGNMHCogB2ybsy/KTMg9FZ0vd1oAIBFFkC0xFvsWWTaYt6LtbmGL2+70dayP
2ibmkcQFMKsoRensi3j8rAfBcN7P1+ShpqjTjxaW0MB/Dl5bvaDRJQl+7mUUT8Rk0rm87oB3XJ8z
jv33mDwmSZ61AYrwtVVbxcVrwlFRy4xPb1EmwGbvSo0ntU1nIy453D7aKHodIHyBPtRNTXJi8vYJ
W9UWOeMSzzgahKvi4NqJjvr8pBmjWmSNAt6CyJQYnOdMNb1/K2WA6XrJIVM8ehtIYii+QmovTq71
vGqXQWE9YvEBYUaJrjIO02P3uCs40toPNunPrAPN3IocVBMoxC6EsE8h5sowlH4+KsdwfCpyMoRl
UC/oNohfGu70raRJamKJm/rt+welViwr5MxFv7mpeIqnoMp0PR+OHo3aaPR10iBktyggLggNrKNX
LHdar2htGFHB3PeoPB8PVI9K1VqbLVjAPEiubUvVIkbVwNFlRr6pA7x9WlZ3tVNOt2omFTRxsS8j
YFNh7eM3iVfIIAGDrjFuEwwm+i/PbFagq2pVCL3U5yu6OvWUlX2nRDwIJVXukIj5pQFw1MeEzsAw
aI0BM2WVBvlJrqPkgkys1gqVqsBEk4h1rTNVMbuh7rlyV4S0oDGqpi6icrqCpl4/ZyqwjlrEW9La
leooTsNioEiiK1r9NyV1oCOqiQY+pM2UWIy+RiVk5MdoHtOu0Fu6CO633eg0CObdqAZMuY3ssqSN
/5thoJupAp7zBAu/JFDSHC83IBedGEqYfn1QFstGYzw91o/kicaf4Yq9aFUsCuEBF0kmyAthhGP1
+lm5G826TPJYgLFu5rqC18ZOIcZ2WwrMBE1fmEal0rdzduTxVhU5xRg6s+JY7khMKouDEhg0Qhpa
cJkJkBPPrOZUJsfOJSsN/zP35HMcDMfA/vZwifTa3Hp2uHm2wRWvaF084CZuyTXEUPbthJUeA04u
E5PhQMW+tkk0vFt2lCrE17/+qq58AUYN2DlsrqKSuqHwGLM0y64B/3jFgizeUyg0RyJiGsmqJI23
Aq5uCqMvK3QgMebyLqI00f7gsVj3ct4ZwZM6l5sjzLg8/gy2F8WYffMu6ZMkYhVWO2aEUxSlWlml
b9hvbzOK/9CyU/1HEzeqOGuuGTmafh+z+0lNRJWMOj+x6pu900dVoAqW2m6F7Vn2gyHiDLMY7gRk
4QiFxVnYUfvBM23UxN/aW9+VCGrxLQ8UOnFhKpHZ7CESpMF3Y/Q1PrmYSokVyOGNAGPVuIxq8h88
/CXolUFZuA95aYNZXvLDkUVQUFfZETD/uklfxaw+qVXcE8NyWcvA4Gt8ru1E+pB17i73PzedT9/d
/BG+r3jEewDxJn5QfHBcNGhWyaSITLfbKXa/aExkCDh0oovPdWPACCxguKPrBrMVTXHnAciuFZc1
Li5QyWr77SPhPF3zdynSr9sM/r7WHme2abazVohLqHTTx+lxtmAx2adfhPnHcsaIDcdjwiwwzNdt
frrrrgUH93+cDX89lADC+GuzwrsES7nDc41eCeKbrHtfPHXn3w2aWJDpGZCdXfmfmeWfRMY7rpGs
I+Yu3PEkUOubMrAQZAvRW1UCQYDKhASX3gi6fNVnHC0g0YyVfX4p10SP3JN968XYd7dtRU+y0b5s
L+kuLv7TnUoSJ1wexlDT1Vr8YpfN8wFbxKFOuxqVxxgQEfK0O6lX4Xxcq+8S8Xx+7R3WqL2KWdWv
X5VRDX5RbC+2KIoqZcoZGF4qi+906Ob0nQBYhlVj0sAZ87lG2H79pI+dOY5LLSJJkLPg/MUDrKID
g50doy+KPhW1luiA8zDTWGs83gsvR83VSmChWUMZ1EReu2l6kb40KOaKUmipjsx1FBW1VUaWvcHY
uiDb94ADGna5aN914/eQX0lWY/lLEqPIlUALi1ORyShp/+VRok2vouM0dlda5HrTo5EQ6JWGf20J
jNaX+IoyFWb0JdKGneYXWeptDZ2F8Gpt/Huv94BnlPzWTuq4sqckAW/tIu98yCk2nv1oYi9gwCLh
ostl5am0aLBvc2EzDvE0dE5GchxFuRzN0C4itewDMZjIivEBud78eAuWcmuIBHgwIGNVfFlZKnYu
ToJAL3Q1Xz9V1F8dlWiJK9iLKLC8gRKdeO8XRPvqw5RIKXlgiNpdo8d2Vp6BjMMV6X6a1/tuTcKj
d4Uujr7NH6ZYk9C7RbYDLm7LScBX+f0HkHsyMkOw3vpDLqfSf9jgHzZxOVC7CnohpXZd1zuvAOxb
13TntdYl7p7a9NLkYFR9eg9Cj5UJ7K8L6LF07THwSrQd4ZUHfCd+ICY36CHX2eOSooJSiZg4tMVI
ri0bKkOorQq0rSskNuL81+Y86X/StXRtbOof6bCWwgFm70+KDKLvCA04BEo8dDgZup3Pt9aaUaOC
0TaGtsfMpSFekx+jLAMSyEhuQ68t6YKEMAmbLyP0oDmm7XqMBz+/nJ+uSQHaJBNM1Ejeu5r2wdT4
gxayip1Kx7yRuvFC5/st3+CRxj2fq5RTj8d0qxs1OO6UmFWoqNlrhETb39LirdI9wWRdywwvSFow
ZfZDSQV8BL+5GzPkMn4zO0Q4fgjBDrRdEPygiWdfcZj6ABKqpL2TRsxF9etrIF/Iqz2/ocSP0eXS
VyXHC3jD49VzTweTc7VcvBAF5Nyczrm3eNh4NkEWJ8LZWfcB/LhxZaXH9HuyHi+SeCACOo98ufO1
Ja6dLfz6mBaqYVrrUkVWSPb/wS4ePUKDdpDPmUt2C4OfMZM+bZTkkF+4bj3+dvA3+Sao1sLIqry3
vM0GYAYfyNXHZM3c9D7jyKQloQroOR/uIefg54/IigSNj9ciVXLHIZTkJ0KF3/jXL/Mmbfit1AdZ
sR86yrq71ZTsKIpVU9AZdyN4Td1ljkjMTWuul/ZVo8nQOmuqLKQvM5s9ycxrhNQScUSynkm5cto6
iPXxgnkOvUnbYNTGD7iORnnhGFyo97vA75wYl1GZiaXViud3nndV5DZvuE5/aKUkatR0r8Ehx164
ZUigde0H6VLCC+QlYzZTko2xEhnUfMjlSDFAwlyDSWRB8D454Lk/PmxtT1A1YyPDxTtWnGH+VCG1
xY2pumi5f9ZhGQs3iFopDRPIw8XhJ5uv5YbqOcJQ7i/+Hg22cfVc6y9LkqBpmM+6lIdze5514C4b
mNVLTgzXK7x1WFZyAJzZsBf+lTSIJ+6KoN2lsC5/Dh+BEL1c/hGlaA3AxNwB2YY5gyJE5q6k/dS+
HtU1aEm6y0jkmIUrC5CaTMc/cAnwZk8CHRvvETPm5OePQtacNW4ttzvLOwlKKknKmnzJqkUGlfau
DV3vh8nkgHx+zqSI2RPrd8crlDHpY+Tqgb3YdPjiFE3KZxTRPyQKkiNMwTNfyGzXXeoLIQXHf/iR
I9VRc3459RBPscoNUw5JviaAx7c6lJUvP0HUWVSrtevPvhuRlSPcfXri/AQdpcflEZ8sCMwaPgq0
/Swv8VkeAPd69DB6z9N11bARKCWGJeTldJkgvcaTCUetj06HEmBi9vAXnmf/0qTc3Vm3T2SwfLaF
S+Z91GpWrQQbLjLWYPQMutDA7PEEWpLQP1gVW7bSkBR+eTBf/ugL+Nd4RbUtrk0aXSTZ8aEa/JWT
i3pCvacD6f4EOulAiC38OSFO8/eOJmrxPauQ4RXv6IFffGUrHKJrEIDuvnED1GnDRZrbUU/Dzdqv
n7LDskXKjma+5p7soCG0pap2KIlbBMpiMyP2Lgi9dxBJjo3pSMOZVaRndwZGEUIUyOjvHolGlqhd
+2/IJ4UnoZ6AKP+4naScpNOxdWK2nAeQweYhPf6Kaetg3EFegMjnx0EBOpNWTwOc5g11lKENTmNM
WvOF/6Kdl+uqhdCFwR/flhDaeO4oqFjG58AuKsu8hh8/1QXe7F8Htinnia8SpTYgo4hn2jSyaM1f
/Ag6SzW++ub4V27Ak8T0dhjsLdFx75hpM5PN1SyqrWUQB2vrhR8PKKZsNxrz0XAgzuo/XJLhCRuC
emTWGqmsQYYcs7ZaGxtFIXce6ok5rk9zbtBzfR0h9Ol06StMBAFO32xDb8FPNMFXzoXYvqkfkqoB
sOuRIEqD4/hlkuk9QubXyt4yQ3jcFQKybWc28rxK/LmrtrrqHpf8cdVTTJEUqlXrAW9vH2c1BLCw
wOnMYt3uwE6Y/RdLbkcmIBnAbJf1iyWFoGYYiTZG4P2XBkXthWg8R9AWyDp4ebXZTT4Xr05m8TPN
6lyA2OitcqLMY35XLxCoVeNEKpYOvAh0baVa7CP5n2lFh+/NyDoMekQ8KyS8lxuqyE1kgDE0tQud
/wtrw92ay2pVnN5GE2hZCaZPHXyXvZ2yWQ69c9l+ptElGd04kSsPrt766S7Iacn3ErL5j2t5z+QO
W8EtH71xl8fEH1DnijqHkN/Mfkjvzz14cUwoY8j1zj0d5PjcB4bSaEN+37lTMYAdTh2SXBQQ0mPM
0ySWhEgflNwKOKSIOE6Z2HdrfOqIaNNLpkIr/D5tSqBH9fMZ/XvBl2OaOGUfgnZ2pX4LXy9VA5s5
bcw88B8R3hMxc9VRtmoWPsHnvv8QoYOCFbMu963yAMIP3+nXfCyxgYV3RyKgruHC+8PU2LTt98Ed
O41bDEhG/wwhsBbTq0++MsqXZrW1WvMZxAwsXOAK4+F2vA8ESAp5yW75KJGRUkrhmR5Y1/8TV7gI
5iKuWKydeDbJ8IXB1Tcsp5yQklQdEPC8V9aqP0dCC4Y8XpX/LoDHFk6PXKh/jkIeWEcWSZtMQSVr
kaTi7SNQJROqqXQU4tC9341p8tuS6IMdXavIay5t0NxGm0S68fDLq1bf5i/xhvAmh1zEkLGCtQTk
lflA6lg4OEpD96NmFvtaRc3RhUmjKeksXcyfhtpERk7utt/scBfXggj874fhhwJrIhnq845Sq8eI
uPqRO7dfrYRz4q3388UTEl5mMtDBb805q80qlkSRqw8++HpNjxnjZnBXDBWQZD+zHKqtKFTKongG
f8Z9ow4Y1FP2wgXI8Td2VSJl7Q7XZM3FV+XiIfR7Rmmu+MzweabCkYPmojvIZlrbWRd1lyN14sPU
Z/dSDJfe3Wkd42I45w9qSvFnXGWNkYwVWAX0+izXQrQxjfkAzJWjEeJAapGLRYPKTKMxb6CNiSGb
hi5DqG8FYzwcwzZlxU51pTv9RTmVIl7RC49EvoAUyE1lgflJVez/I65B8sspFnv8PRKZD32YLHYw
5qYRtSDeeRHNA5OhTs+e810uXunCoPhUIyb6H/SNkj0GHYnUv52vRBM6tW0OvA1E+UfcjgNbd8XM
OKntUkWB2e/reKoTsSTO7vdU3ZyRjZVX1gY4Wwx8vcmQD9XFo+yPckm01/2tt2mOHNtRqnCxiDQe
3gvq2KgbIkeWnCJvCR0d3RcVhppRl/otMpbZvD8A3vLNhIAjsy/XYooXUxRi2OuCAM/ake+Q8DTV
2MQdT5o4I6NhsLBLynu7eT/r5bhKmfWENYG1QvoLH25dyNJUAyt7i3SrgBSaL6BYG3svrqXld5gi
t4igN31H/J1ogck3Ta9okThXC6g1Er0ZI0K3TZRunPozl+j8XyhuDDcEZ5JjE9k4mv/vztvlbmFP
/+rDWdAM66jX3DZj/5rr0mCHXzE4YQERSYeQHPXVBTY4eq43qacyxfkbefV5Fwb7SIg1Za4mijTZ
5WGWUnI8dRVerSBu2bAmTcsOgBZ3WHN6gw7naYmpRdZk5AYBEQSbIWqGP7BMsZz/RGF0yGlJZoyA
WTykyVP1pp4+0i2PrdMF6rqxGE9D9kG1WkoOtP1S9cbNHb4dwcAjOxSVICfqiIAN/cCfZdGKLuEM
iUsnyK7K7buzVGaTGr1KDpA60lVsHkR0m8IVswSKGkCsxX15ooU5p/rViouoGN+LuuJUX00Tkt1M
c2jxr7R5zpxY8QHH0t0U7lp2VPUqtYbkJhIPnMdrbmepeAZrlLWNS4T2lBYRZkc0p0ZcwXfAeYpw
KHOKAx/TyLS1kaDeEdd8NrGeHcJFtu9q7tJ0YH+vLsUTYx/e+7T0pZM4ERCSBYwMK1ReYZkIgxMD
bWQN5Eu3f/q211uX2oqUkX+VsO4bphI1A+lzb00q6vpEcfAsj8ccir7UZS3VDrToCUmyVPWQiI3W
pZd4VtjGXdt7yZWwZ4HwJcRMexPDO6nvLoywYwqPn5AVm7dHabcv1qmJfPRGURiOQLqPla8ueaoq
nbnehDFQEVqgJGZ2eAW0AjGebTytUne8bRSPv3mkPVm8GmOfVrfF6nirbXWwnqtSlI9GXLSJKiRS
7U/PagdT6giauebyYhE37CPdZWfl9E5UXKadz0DnrJg5ZM0NbNiAOsN9bUF1fjvScM3d8OWZPBsU
VNHxEHPxa9eG21kdXwJPUnq9ZAbW7Si0VL66p5+V1D8FxB92Qv85cKYRnyOiIWAyWuj9mj8fdbOF
ML1wHtVDFhmJZrSg/CZOphwqruBWyl+B1yySYB/roLYdkcU96e12l+mLGk5sSx4NoRvlivI3yvtr
bM2J+Yx5+/oh0+0q2jRxW9RYdugf09Tv+lX3QQ0FTzvvh7XHj6LDtm1ClnNsJzQTLGbxo8NNK2Yi
zWfGLkGMVTfEHhS5VswZEvglQR2nIrVO+MLyflP5T/eqY9ZKvTaGhgdYNSbJwtXy7KABu82+3aFF
I9HUe3pubgHP8NBKI2rfvpJVwBCWELmdRXhRNcGgXY1J4ufXlKCJjerXSBdRu2C4scnV0/8lXQEh
mu/GU9ip35ACq04u2jeQbG1nHhLHUj7sUbdxoi4iPHskSCuwnnW0KHkJ2uqRlwQ7TJxUGKmJWH9i
68Di8IGqhvF6sHMZxoo2lC0IRKExf6JrTaExiyJ3FWkoPrsmPl8AcMGVEXksi1nS7VP9vQb++ufK
rAgjSVEwVBCX91YemUC5SHxb6zTb5kGcG3d546mXqC+P13ZdaE4zTLKptH60G5998WnXHJgvhj+D
Wud24mRb9XR8dTFVo1fBpR6dgastB/UtyDUBX/UjAF81FF1E3jsyhbaVtXS/F/ndgGkx/lKEb6xw
umVWJrmGE+wyWg89izjOyvrZETfxnN951tlyiA5rKAvwnfe9GP2b6/yeEmcRHxpDHr8CT4k7jidS
TWCX4DdgGUDXFK1PpIA/VUQJo4JbWBcCZX/vR/WUOUXyzGZZoN0Vr5IitELIH5mJeQ2SD1jJP5pY
buG71DppjdOpTnq8DHm7bAnFeuVIHMcy+HSZTpGvLVDATDB3jUCJ5Ts/Flb4s/q/u+tdIgziTFq0
ha37PQGoOfCServ4rJCCQHJiEUfJvEAoLVJBEGnQNmBm6+FldPZV7EfcVJkF7ZlDBmxFDIGd3nix
6k5opYPtD6pWfMMFztNYLDyoduc6usY2nasha/EJIwHWJDUwk/Y/m1+fLRMGy03yVxafx9NyM3U+
Foe3X/0dULGqm312UvhJaeVczrr827Rp1/n2oaTUHotehLxoJ0ZUZIYfLhWSxGbBFhrnWRlZc3c9
FXGant6SM9WwRKLx0Er4n6C1B83ZpytxzMXl3Gbo7rGxaXumU3wGKxNaLfode140Bz6U91er1XQF
4GBPSUPQinIZ/8366F801Z6K8KPID8MogMsY2CzbANBtpzQGV4RzSwvbBR3Da7EwNzHHhv6lNrB1
M55dZS4ThRUF649pdtSPvAvzGVW5snTMqPDN8yCqP3WA0w3sf8EKNGtAr3YJbFonbH9n7P23Exgc
FsT5qxwufraK/cDF90shpFwyAoX69qvjaI8vQfua8k9MZpPme/bvMHVk7RSQBoxj1XNP4sNMpmhN
8e1ljFy8EUDjre5K7MgQJheLTjxvK/tzhXCKzL2CKg7v+tlFzWNCk7Z72fkYEPFEBjX5RDUc/6Nb
jVfXkePvV7A2kTRbsJh8dTFXkUyMY+Bs/Hv991r+uZzUjyC4Asoz9VkGtwiu39Bud7ai4opceLu3
0BcQe+HLVxF7jj9tGCJRHkz9XXY4HH+pBvOd8BnIHQI8kPNwRHt1fbO06t/4sXTWYLBPXtwen/jT
Hp3yJtdyVb4r2wX040EWBQdEqliQvysF0zxR79i6Ox7R87DvIO6QORUQEhD2vHytl2dout+9+l+5
baGoSAHL0eHcHQ2emQWtg1NJOsjk8pM7jqSigu2bTioym4DBDLZjcOuD8nzkoFZ2yolOG9dWOsc2
1hxcoynqIELMu6kCasKAiOjsy3CeWgwNjFHDG0+sZvIIUqRkzjMiApIQpwQ+9r6kYOk/r9pYWwFJ
BOJZ9MCAus0dS/34ptJSMSqVeSE1ogcbOolpJkolhU5nu8pPWt1XEBpvFdtOHOot4Q/2ukQtDMBf
h/boeBe6kZnNEdKi2aGYrwvXeqJZ/WM7mYHtT2Ev/8obBhFGL9fOm/q4V93PSYFQ3Z3CuKYnHDD3
VTo7naf5lnALCOwdAcJgEWdMRq1eNZuSXyFP3ysbYPENYrkmTSwNZL8GP/Nc6V3FpWJ/CyyICbs+
GtDgBcDu0fAAeplBdIqbqbJwEs1eCQwYhkyY5w0vd270ekDgBqwHginRURCfWaFkSzlrdwhewqju
J3DVtXBJmV1aWIcRzDyuoxOXR9ljHa53k0UTB0lY4N98iZ1YNZZwIMr2CzWO01XPN+oTujzjOrru
YrvTidMzgwUN/QB9v0Y72sB4oBVnUQWrbVlrvWGBaC9YkXnk4lkigXBiQHhHpRE2XJsZFELmc8uJ
814UFEA/jp3TxcmLb5JvB30W7tgoa1PXzIc4KueiCRtZAn/FHrPUS/bPlsvp8TjsL8YVXcysgovW
oVcHyUqinIPqNxgESsws6BURh2fIknsQgkD29NA6OA6zya/Kao6wwki3Gq+5oYJgR+lHfgar52Q/
629KpmPNd2x7AagXBu9aHCg4T8vuBoxw33MQ1ygqk+L4jY9mnFwvYIX1LMHb+lZjHp2WdbmmDENF
ppE8CJV3vSffiWK7tSJL0+yYLdGVOPGyanFJl47AtuDwM8/KQRZfJq6BxdqMxai/tLjX2DV4fRIl
r21FBtTkCevUKBvjKA2dcN7memOy60zX/cnuGmjbboU+PAOrMczjuxAxreY6ypWMAY72+ps8LABj
6GuWo6yt8J/xhUH5seduACV+CJpU7YwUtrUiLDSznqbJvbZKR+umcTLVt+kBZep9DSGEE2j8F8eI
p+eVUeOtdtLTeL1aNqcpgSQ6E02i8pwUFrTdcNI767aXBSnsW0lRdENIYDkcWz1Phdslgg6DE+Sy
gv9GDZkvgT+IWeroMMN6DABBqM5DLAxVwzIiuis72kD7P4zqWc2NQWXeHOFcLfTIpRLn11+AN4/J
PHvR3pSPBT0I2LgTtUzerAgfttlUuGj/+Jjv4BRsG5wrdx68oS2ZejktlWfvdE/yNU8sfYT49dHZ
AKh1v7wjzj6Hi9g3VJe4TPEaEnDJD76qSZk/KVlXQ4oq9DsuLpYujdG1y6CBrGstfp8/vVWBrmZP
c+XNewxyQEWirW+kmuSemlWXQn5kODhwCKgMKVWeVP7Wi25abzEbYZrK3y9gRh9baFbapqbJNin1
eh9naI2jtuxUpqCHblvVDpyVfBsHAt//5D849dSUPWeSS7PM/ozRumMUhdVXP63tbZYRX8HJ6IhF
bdM+SDVUdK4Hb8odCZembowGc/YwJJc4VUTy+fikRZM2Ep6mvGSsEb5gcYldBZIxU4kQxYd3eusd
U1yeMIuiYGGHB0iSvjPVNQnOkvcwHaXqV+cd421Jk0bKlJ0u2uVxgOi9Gs5jGsv7tRXUBprm5R1L
2vcAXB9R3jUIc7Qg5zDJOWkEVFtfSxXDEl/0cqDS69v4UcWZgtDSY8w8Jgkjh/lPaB8HepYQ7shm
pNZOwv/BOXhZACaETExrrvVfuB2g9dLnOQhVvxWeBLqS4/OHyaQL3Rt/mA23/YhKVdLZs+h4mOBS
5jFjhNEqqipXoB9QeT1HqRoS6HgnMK6HTu3w/YdrEli0nUKEQuWrKrE+uUID1jJYzg4wIP+bLqRO
Dd99R84t3WwZDAKJ5YYsii3YLl4L2eYqYgYsllQhlv1z9IbtsImfL2a3aQj2WCCbrvkXQlX55EdO
v7Wfd8fCGYiMb2bJ2g2bPoiI7SHrAVZ/CUEl1rtcq3ARcBfY17RYvsAoqNta+6KdtZqvlf4IblMF
592fa2CdHsrq66OKQMIvGX34nxAtJHVHBZbEROymcCa2QMJzkAvtvjHtR6z9GJM6Plqu956y1a0/
qcT23yoq297huEyA0FEbN3dEk9mgRBiMrJU5+7qTmWiVOjKFBQYxGpvmn7cIAMK+Sa/uyGdKhpap
h7wHSn1+S1mlAzV2qbFWEo2HgegxwwKxZONXlPmroZbcYjcSOGZeG1UDgd7DqMflUx8qvpewID3z
n1dw8lBYeoSymsncpufUbGNR9iol/gKdplHWpYHc4Ekh/jf+9ytqAlHhxNYEzNcfpThJqBaJdVOU
tBUSeIVAU8jsW48SRh/D09jo4MWfiGDB+dMa3mTrpfaqk9iwO5xG4336p5sd9jIYsfV55b9Jk6ya
dxhc4qjy9M/Zmyi2Ze8KO8J1kARw0dIAlOZ2kIFA2jVi1LUvsC+1mqI15GpPUVmnML30GLGCOSnf
bkBbDLjTgKeLDh17mC5c48GC9bsNltzJztMzKj2/ASjNffwvJolkw/VEhM/PiAPHnkXurWWla4W+
QCXeS8ofxjVxFQJW/3iZnE4/I2XQ2d5AU2KeIXS1hQjS5IISdbyEFiHzLCRKNqMP8qKeUD/djDEZ
QsCWABO2bXe2+3u9Obifz9Nk4tUB+yoWDcglxxaRrbzZhH4tzt+F2kxRR06sQQDzcq1dQnJ0dRZO
Exgzd60eac/8essWXIjPEvXgi0O00y7xpJbRxi2HIbt1CahaG+h4XalmNe2ECQ2VezImeYrnTGie
jJxjR33RNsb19I6umO8GEGwdT6W4aRPYc2G4dCXyWVUcWZqT6Ql33QK3jjLMLdoe5GYpu86Ri0mx
BSbtoOCBWjAUeP2ivHyqf1uPwbJlUYR3zRGqB8hYfytu9YAZmjNjyu/XWGXwdYAtQW8MEs59pB2M
NLlmBy0HCYPNm16D6Pv8sUHit3M/xWcB6Ddquhwm3ND0/yaAWc2UK9Qtz48Ve9a7EFgdhCW4nvli
KKQrvHrQggOxVVf/fvXm+vDc6FZiFzU8WzLbGSFN+u8Pur2oOiIlnwDxaYcfF9MXvFEm0WZr9n2j
gLYiRZzTOftsZME6hy0cxXZwvnT5D+wb+lS0m3W+N7l2vVk01A03vdNMRl74cjT7LCPucxY/N4D1
DlTmm4dHkMXHySz7o5+kfe/WlgZKQ5JZhl5BbThmqc8ue43YTq7WK0nKF4ahIgKVPAXqQWeFVm+O
ZXpADg093BHQC4A61uHJWLfs8Xnv2Gj1/foL5AL0n/e6wzOA2KFAb+LmVqsIotTEkqikZc/FwfSm
gPMr01lHmToSATkZzcUMO93BvQx2dVPphkkhWkAK8bpx/xeJ7NNPllz6kW4UgFIJUwmQtJEo088Y
eVX5hOgtXsAofxBpXL5W+KXdkyznkhDpRajCXyhsB8EBF+wHAp2yW2Ur2DTfGfAs+BwuGl7JaFgU
7Q2cynhCU6JppICfExAVH+6AEV+J0Yj/UJfa6W5vBr699WuyZH66xqdQ73/Md/EzhCgmKtTGvVqz
iy1aobKzWrIWcanAuh4BkBuMJbdOOeoI6OF+hcPKwis7cvamIwSRDoFuR9mLIDmvsOz7PjPbD8Y0
X4w3ljxGiYiaTNmMAovKY3ESiLVbisXCu1PZZU6mXoMc6dB8WvN1yk28x4kHkHlHaaVyLDTMxl04
hvrmjDV3v1BBaWfObBfmr/XDyKXiskB65EKKkMrZAyHrR4/DQvR4KjcqWCIN3tcKxHlTcWN58EzO
ivCP/tSZaELPG7Q0/jaYPMVUqEW8Zc6uC2dP79nMrI3oD7WXYiAbTKIgT5TNU8XJx4RtibsxfKYC
1vzAO2yEWwdWsQkc6RITRrLn3LyPeV+fwqriljTjgcVyJlHg5do1zQW0IZpyYqin+J5ssBcU9avU
iua1GcxWMqoWLpLDlaSDDjwm7YncSoM9i8xyTAKEfNJFzh/J+1wgR1LtbcvrKB3bBDogMOCXc4Yc
FY0BSrDJoxMCKXLVkifLuayawX7ETYHERMnPNc0L3UZEDP5Ownkp0uex8kjs2AWv+CJAntQzz/hh
441CImUVdAE3+xmUZx+qT3Hlu+p8ujOHBaw9++yFs9SyKbKv0N+9Pk69WyqAkmJFkN2yaDB91QIe
APkaSUvu12anBCnVBlmWTPP7TP1FUts8Mfo9Ec6KzEklnunSaeV+A018l2JWRsth9GakyiXeUTNL
Llyb0LyzuJ3FFLqDt8seMwY18Cv3BcuYTVUBC/J82FpVjKjOG+SL00j/yBGaNK5XiyGqL/JVGZPx
PtwsfzZW7Y/2eNOZvBbfH2Bwf36XrBFh378cWt0EIY+lQYZ9iMa+i+HtcsA3j0J94M8ZAtj3ko7n
AaGla8APBp4AYlGwgo8TMG1z9WakFNHC9NLaZG+ka+ES/+jBoGKYExji1Qi+HeBNrlXif+R/cnph
9uUP10s9ggNkaO7ZV07//U5sdkKIRPDAeJqkkyuR4vjEu3HbQGfSz0PocwhZvEc7pr8Xq3UZPyyq
GpA5/N4ESLHiwomNkI8n9pRyeJlAzzUVhBm8g+h5uv/zD5I7vAtUYXglzwg+tS14lNFUySvVY0Qe
RynbupyDP0Pxp8p0OR1JiKVCpqpEZujAG7v1lnG5gsLSznQDFxxZ7eECQo8WubvXFs7wL189yrmv
QFDEPogH1/s7t5ymqNKnrkk7NzXkqSLmQ6Oyk1KYeNUdRXN+rEg7vZIzcjYJwqKm384xyN0rD9ZN
az2LwJZ2Lc4HI969HCRux9is6Ge6dm1s6i4E+1gzO/1ej9NKmf2R2O+x25E8SXb5TjXvignkazby
inL62SukLYSbk3lrlgNN453wPGOAF8kPwUfY+l/58BM4RsjNOxmMMbDtMoJURz6NimUg4eKmhzAr
/MjEkyXqtNvR8iHG6czcNCLeMR3AiBdVvrGZL3Oql7nYQyRJvf18aSqnzDmRQk4pO9lCdtGmE4Uh
sh0GxvMcrO35LyKsKWl3iawr+les7wkq6N5RiSEZNMuPzGMQLRmtM1q2rJFRJrc1WMGvVfUnmgmK
D/BUXpXjnwbRETEmxToRBYsvxjuaK+L1jMa93aFL82jMoLcMjtDCfGjaylUCMoxfMnoIeoHutIRk
dxflMrTHaLGAW9cFBcKMarfFBm0vP8AybcgXOmk4TTVXJ+jVML+kybDEi8inOx9t+fp0m5rAatlP
3160zclKys9P/0UdYcNo9kqUZ5J33Xabz9WWCYHikvuTJo/0vDWahIr68hRlLc3uk1Nf0HHKJNcn
Nz1XJLT1arRqSr1NXWb8+QW6yo+KSZjzofppMivcP33IXDUs6+DnuGTQnew009MSt6PkxeI22qKD
YQWnc9wzfKFgJnoKioBpROAUUeEwCqXc9EKNt4PsjcEgEQJMADNPpph/ZP7m2Fnk6NqukRAWsfFC
Ik5aU+o6X6AtGnOlqKZf4eoIXOyAU3zXXNfsLev0FlCjABPTbnkfbHV1XdZRDQJAQ3sRvB9luYZL
DsdkoHjbxgQ5rVBjGi7Q+fcHnjLMQgQkkM0aHxhZyWvBcKTJNYGhmT+973koU+izbXu2Bi0PYleV
L+E4gYOkCLAQmYfAtwod9hiKWb0Pg4FBXGKRdZmCLZFNJenfn2QPdAz+L3424/j96PVxhgCtjtih
0QlNYyuZy5WPNAE4pEQiyhXZ7BB+7dpPNNy3aPscwoKOe97OOeslD8B8cgphosFTq01ac+qoigYv
aEDwpbadUyesv/22aD22Kdab9y8ZgZ6+8fRXCEaO/ziloMTcdZPxuk7wyBgIoOhwV8jMy355nhHe
ltvXLLCfWKJhIM+2VccJdZUKKM303afXvBGKWteQ+oN7kpT74idykF5j4YGY5KaKlEp9Ry3TqwG5
KqugVOapXg6exjb7dctXbejMnXgYpWumPlUKj7FnTayNgpwl/J+ft5ui7rkGl20+Ee3ZGRKH65Pe
kRrB5OM4YZOcCUptIIaQLuRolzRcvpOiypFZI7eoq1xjmYPaBpaNOi+oNbcN2hXzemGEuw1b4EMQ
QdAcWHHCtmBITy2JVcRIGZQJ3xrvq6u86APCd19tZ5MNqZFKskooxbJokBJDONlEZmLKkwwsSm1P
iiREWqW68IAxtA4MArWIJlZeOAiCGLJV6Fv78X7ndmxUv/bCAeb8R6eV2HebNVNTF94C/xRyQZoU
wLF7i33My6lsZWk4bQdnJDfidAwYDjyZg/0hYiPmcYtk1P15dZHv33uFCAHKsBA2agq8pWHTxacg
RJUW0+9721FirfPgZsu7QzUGJn3SotTne6ork1UiAkv2pltNRPoKZ/++OFx0//LVitIsI4MBN7aN
XI+iY6QtWLk7n0XMicsADonYgmwY+Q4xy8aXYx5mm+QTsOThO6vbYmAEG1U/zzqB1FnHoKZ1LsNw
b0AGCrTA/PkVruMZ621P7MTseUgcQowYfKM0lssZRGWSsOYRj/BAK8QAhOR3IQZ+iu2zqFUiY5pv
A9UYySLmypHJkPgnD2sknzUAwY2vjNnKg0Naylr+BrUaAQkotoz7nH73Km7/GnDAoN1ew0wp/zOP
32WL2K6U9ruuJJ7cYbNuqITogSPMy1KUl7RyX6GtESxyEEOx6AO0EeIxCl4aRIILP/Jdkrv9ws8b
L7lCQBll8tykS/AwSNvJ60WFaaa3OxqzehvHVhCPj4WjD64q3pNFJOx5uLJEdx8SoSxOUJQQgPXe
Nurv6vSy6WEf8clXCUy9iw/pZzemHslNcZK7hrRT4PiPwJ+80vr1goOZF5y/ESMq4H4EM3tQufys
YWcsmH89bsqFMTl+opuuG0UtOOVItW8D0E291TutJjk6kGS4cGXvwj0kDBYGu4gIAeruZY30wqZH
VmKAB8FTncUu0TD0TgA7RYFZr8eepV6QmhJ4XcnWULeisBS8/7udqBSiov3tEltsqlhr3TLvk7D3
pnP6zhXmB1mB7KLfcDW7yg61yHlVGISKxppg64bMW6V+lvlqVMIPGtbOm7tX+whiLX2Fkzhn1/tT
oo2tN6enpcsdSv+aPJzh4/7yvrOyVzWyxv/ymdERPPjlEqzwJ41AwxVzdaox/sbCFedL2Mg49dEA
KdosdDbKOZ+LGFvTL64735/y54U5OaiNl6XS0kCAOJXLPkorM1f58rBpWhiAXKw0LGDMk5ontRfs
62GybLPn53vkOmNn5ecfTzMcYohfYwme4thfoy4Ht7OVUSXtJ+uFCObdYbxbzT+6PNqfl7xzS2tG
YWwEN6oS6JTa4Coc4mDahDR9sQZ06Pog8vrF4ErARBIvT/ma8SOpjWQNs3VmMm2ofzqvtxV0U/zG
RLGl5OMQIrcBKQceeflKiDYCJrh5jbXK66eUu6Ws4gFItoJf9w1cCZHTwSgnbrosJn4IWUJvHaJB
BivdXg3TELgT607mVwr2rkIXBbAcsuupMKDMZlE5aVvIIT8WQ6+aDWS6+XHsVcFRwzVmPUXx3Xwx
Ybd8ciQdqdC6KLh9100+InDQG74jmyNH/Hx0YYoqpcVzm/5LbMTYA0Q7HXAlpjsMXNUCs4kGFlxD
epkKx0EUi0mUWRCkFKJO3R9hv0KNVxbsfY99k8qziAFc6sma4yv/qay4MVrhUWAyFP/4pXlxOaZV
MhDw9v+4/teMPQg1YvHLbX4tAgJAiQcZmRx/q48SgyTSlYHbdaeMwkl1U8YZJTQU3Jnp3dYNDS8E
2okfAOMPzpfSRfPjcRigpZIKxupOF8NAXHuW7OG9EJWWnSQ3DQk6SFg2tc34PMoKvgH53A+b2Yco
uR2apW6vjfqSM0uyH3HYcnaiQDFZrkMNfKFFABT+QtDumhiLTRIXwseVjyGskPIwQWg8qgyR6rh2
tLQPyVTX/wHaca4eELNY3AoWkrHED8UjEPyoW5sBqrlZooyjRQO2KLl2DQW+7en83PGYPT+xKpVh
W+uGEReDx42D5HkyNoFpYOjqpkdOqRPEVdYhkWLQ10LtsBxHtbLyFhW8G+GhU/3IJ91532KRby1w
wygokCDCKnpmoPefnWI6cNn7GAWiAp4oUKcH/egbyOtq3RBir70yJVMfIvSiS5//H8KjhdMn7gcF
bPG4ilE9+WLcdaa+FFQe9goW+w5QbFrq55wCfaJfvtUtLWkWriXOkoO0nrPTvD8WNqtI5GjAloKm
QSwgg38t25gH2Gwe/aimwwoMBRk5scSlItmpwqdNv7LDZXf3PVD0gZ9FMdreKtZxwCx+YQdxPnBg
mXvANRMVbFCZRgNUn/eZj2RXvxJBA55FR2ewEqdXiAAPfaZpcVodQeey7j5l8FWzSORr+BoiMImK
TCnH2LIox4g1LeABp726s/SB327xODlYQNbHw58MyWUnkQzsSu5evqwkEFocPuegi6JCOIorlHMe
/lwxw+sgrQfIaySeN2Isq5nUSa2W8cV6BwgQrM7odmu+yBMXtGkB/VtRbAtSrKzlRcJpGlttGUcO
2j6wpTs9yRg3vcU2tAtHAZQZmjDjTew7nUK+oknwj+qMksc1gGgmKkcaI6gc/lFCeeRHN0xkNz2Q
lor905dB/pjEDHgc3E05EGDSxE8er4JNJwAGO4zfh+8vdFlVVbXmab684iA5zdDHouIV7hIW9k3B
gueZXzVU9aEz6jA1Dm8qsZTXpaUuDlB1Jhzavi/Yb/CKgonKw+5GfoHIhyrZdm+ISQ8uo3t/wvdy
NTjRSeNjUqeyMWPceOcQTuowKqRJSvEiYmJH9w7wxc/r6ydRJnAS5JG3JOofcpP32ZFBieiAgIKk
gXJfGXZmX+eO3DHYkE4SA/a8obytEOi8aNlERnBdQJnywqOKN8iVGiadVdRSGM8tIEppvHKogpmT
kGh2YTz/ZY7DtxpZSp6Dp+zNVgguN08pUUdAYhl1KRY/S+Omx1xbSHRa3PqpDbqw+dgiIh/XBWd0
KijitAqD+8r0fkHnwxASG/yd2BH8AMVU4Nuquup6zByflcpbQUnvmFIkqCW/9USBXmw/02oGO+wB
kszp8GjbTJOtE/B4D/+x8yBSBbMzGV9jv2gwC0TZHMa4vkvBud6X8Q1eHGi0V1+otUQay2P000Gg
BJYbpKO3Sru95jmHN9w0Q5jTI0A3dAtbUeRMygUs3CljAJv2YY1fRr9oh6BJ3gwjXGtEDuUzOYbt
WWJWzCONxoO5Ox22Rgr4Oyf0x6npy5zYQcRUft3bkD/BTW94CgnOk3Y5lQcCEVxvfrcOPzrh84SA
HKD4huADDTNC/nMVGGBlYjqxS7jq0Htip0qd6T+Mj150ngzhYZPjB0MRiw1qN2zLzJtEY3C5rEi5
2Px+51BguNX2VBu4LHZorLaDKC59GTLWZOJ90dwt1jPtfP1iFCSYA1a+5ToS9Uv+n7F0B5WEDJO2
bfGfgphAKvd8hAyqvqbYdcfe+UTqb8VFwVo0oC1rH2/9pFHWmqRV1JpkCu5Gz3ay6INxmXmfuhNp
LM+eY6LUToRU51DKru73akCeS4OKvDt5HMrQyzN0vbwUve4mbky5GzjjL47lMjXsd4r0rQ1Dohji
MgP04e1vJfgY946Hlpz9MMUr/FuVf37o2SPHjY7UGDd+irhd2yd31vDrFOVY3ZDvVHzLht9lBRao
aQuPUo3xSmb7Kaq2LYLZgtowegEq+LgjCjpTQSo2rx6LSpkxOV1iroZnC+Al+k2U7KyWb+ANMHND
U8xR+IDXBIy8Ts0JTdyQmngaU71ryBGSWiZ/l1JiQNIYSY5y76RyZ8CVlBqv01hAIS+nlHQ6TQF1
cVMygcV+NKIbKkTSTKyyaiH/vxdJRBGUL7CXVd2bByh7q+LpnYsdyGQb8EEgNT5x2I4bEa9sIkW1
hpqL4cz7qXP5ixSIxOJvu1VtxU+siSp/54PbVN+NDRGyxLBc/emgsZSdLSvkvwJQ+TmxbZDtBqev
PENLaQvdP5U6ay61Ut9Th6QBQcPz24l3GTq0yN8D07L9dVYjQTwDV2Gu9fnnwzOCffNVEBbjRjqZ
U1BMhYBI1X10h71GIZS2zenQ4VCS2YarId5I53WKm5PnFWGwc0djl227K5u6+kN8nhMBnmDmn/UR
QC2ehSzvKCiBEhKSbPm1i3E5ibWBnFEYT8EWBpVPlSWvbkIE/tGcXRXunt/q681Qb1LHAzaQEPej
SOd3Q7LcyM06DWrPH/c9hTNsOJUpysgQKT9qDqEVDTin6aJllUUNGvLuQTtEyHVP7aWIb3ODILCs
dlrPTB1XXtTjN3YKvMETf/iyEgdnd/HfuerRx3dhWXQJMpjIi0DWdcXuOzQ0pjgzRIGyiiiu7+5O
2iUyG80/kurjUTIWLYmmF4HemIqtynB5qL2dToM5AqG5QQ46NNwO4UTsPThXvHoTEM61WODoUHNG
Wt29cb2MOzj4Y/G4Vsp5o3DpHnjQVSuSDY0Rkz54gZhQI/OP4wW25Aaraj5vL/aUdtTEB3FF0U3t
VBkX0qoA/TRtIzVU604Xjz2NC0vBaMPm1h4vt1kLQ4gGviNZSQs0hFjoM5jno0LLatUQQotutL5f
vFaIGUpgefGZwhkTwIyxCs0f9gzUEetjAc2FhdinEpLPWjYOZl3oZYMTEi7x98Z4gCIBPYWwq1bg
Jn8E1zXeWoV/LSC1nvRo0AJsA+GmAvUnzzmQGDF4MyHMXlxFzWeobrbOTtH4J0ugr+VZuou5Z1X6
ydqIONROsxdBE6uP4CLYRQrrvi5Vh4EZ05ntkcBYMMKMprXQvG8zEMCNAeYKm42eIEgcrTGJ/DGK
hJ2KMy8HDwsS3FQkvEOesHOW9nW7F2CgaOEN89aN3AhFL/cTp8dnFkmRV3mSjotP/CglDjE0wJp5
LF5LiLDjZMlzfYQjBIbE74hDgRkkto5Py4o7HDVmPGl4F/DJSL/0WhDkpr12cFGWjSycqaMIOuYb
k20eQhtcE5+S+wGcJYs19zQ6xshs3E50i2sW9aaaqhHFx892g7S3M0dqbPrqeyvO2NoyiuqQmrRV
2ROYBSQeYHpvQLktTd1N/32VL+MAsl0jBNCmtkTol/ues0FQgeu3Yu2qk2dQ3rpdDZcGhDebFSAs
e73+uFCR4scu74o0906cLWll3nIiQe5KQ4ZqgYVqMHn3IZmcVEqjyPOZFRL0DWCFhE3zgAwxrBDi
lwC8V+FH2WIl3MIQ6GsG0GupCkGeP2Zjye8X+6FJBABVdG9GJyJJ0mz3p5KrxxqVjl7/G2avemBg
nf751U22R3Bew1QN4unDIyubaj6hvHxlQAn/dRHdVpFQk/961rf3ztQdRXHjIV6LVjcgSN/OTC+n
XyAhMx7QfcLNQ9RfOrBWLd3ULujIRlKrwMKxxVr/3d++Cuta24stR/qJlxIIzupMb0Q1evyqgUbx
T/kvbbP2A7ajT77aif+/jnNqhkPx+gUL36HMKnvQqwtos3Yu3uUcx6IeaKGkmknc+XpSQOR0aRJN
kE8s3Ibd3rhVKRbnZ2r8hy69zd1yDnW8RYZhAfVA0cjpwU7Xafjf2LtkCrmwQSy6Or519o2dCpO/
1iehck+do6JYcwCyujK32ggFvnE6emuAOSDXBW+8pVH+duYIMAmCCNwtkwoYeQ7M6cm2srEOvkzE
TenSMChvT+aj0Amnlq0jHARC8TxKG4ruX67mNHGoVeP6twgvp57R2NgyV0sRhk5sJDgdzb0uR7A4
eaeNZOUGJHXqM14wIo2AmWhqdoWP1m0kuSlvuI6ZiJdbWkMBGIdR5zMGql8cOiy25CdkZzBveQFV
iXU82tm7qtDf/Xt/TlTMvX8HrdmfKzfCqgkZXAfUtZ0COxYVNAn3qBvQghhjwVtpctxTfzvOPlQv
csKcBUh6lUXIskdFDnORAYeQIfFZetdvZ756ODKrwliQVNM4plVajD/Cvpl5yyQMN6Jz7JKR682d
pHkNuuFIUfjxNSBjdBIubLoe3qKlotIY44b79zyF+SLmV+BGQlwaRunKNeA0c23XWUpW9oqMYApV
GayrDl0MIXsGhkYAjjjNEzXP0J13jULS8tIawKZVLCQvFqrlXidAJbdxtf61yI4HsrMBrMgRAKW0
FBNwpGE2uKPKEqKda7Oczc+Di99uR+MsPv0IwkdwdpT4bmZZAmSlwKzDRqgeB3RPCOtMDUBE6dGA
KZ9Nc7d/g9BCIePULrLf5IDJgk++qYd0/k6sMB5XYjPUsHD4Bn6iEhzK7UqHgi8XjgkbHBTADe1I
39sw8GRKRRhZtr9lI7elBX7RE2gU04a9WRGMX+BwPOTmjJQih38YnZ2Qx12Mk3WwpS6HnhfeR37i
AGy98IizY4rtZgjYEjw3tCpPGfgSWzoCe2RDhmm5hpcY2UZywXxRD8XCTgR/cUIDGorrirRWRZyk
KgIYIXPegnlXAIQT+CX2H05MDjRI1dydDvMuFmpSARa9HK1MNixze9ySvEZCDhsQSzBI78xgTTu2
JUR2yoN007W8kVFF5XEtkYMr2c970InQoNP/b/4tjbHBnUaHLDRS8CVUgjk81ixHFUkwpF2cm8fD
OsNC6rOjUdLzlm75kI24D2XCROm49LSjxP5zwuTOfMTmSHEurFXya2nLhokvLOQtBJs7jEt3nidl
i3iwkdOOM7KHIAI0ppo205zv8anQEUAXn+gw/Rcs5C8Q8wW4mqYR87DLRfVtcQykYSyK6gmbQnEy
HsT3qSuHVMk9QkQdcwXjTWLfJMZorXYG1fGxw7i5SLmb/eWOEJtad2zOWSn+sWZ4v3ftZz6ZB5v3
Efr0vnawJ1Ps+UTucgZNa22TzT+Ma6+LxEZButH1adn6I7Ot9Sr1Uz2p+5zWYHmBD8L0+YwcIIz8
KQ66t240NHTqID71ZUNuoillrynN6gyhQ09BAa6co1mqvEdMKpvO3l3A3cErxMUENq5vnanH+bz8
dTHV0rGwTKOv5DzoWLX6Fnfv4QurwACEmwveewJcJX40jr+EeQWwjcnZh7iQqQVTClGy9uR1Neft
kuwDtmOSp7JaVdnEYMQF+pna690JqU5AW6mKhM7bEwbmogmXGNVe2TW7/SVYSLiSPzy9w4eg2m7G
6NRe6c/8wu/b8KXub/Sdsljt/ays+gnwIz5X8USxx/mc0MUbsd19v4W9Ib2VGoKV5tI3dJy9+lrX
FyNb+CN2lXervGQoo92sH56L64Y9E4A7KV7Yju1NbLAF1Z9Ny58JvDZzzvNfhWwf1olZ9Cp7Em3T
SejXIeVpZuPlwFkDMfqFkXaTh/Rce3z0InbRTfwX2tSuY+5hWQfV39A69/b/5o4N7PAv8Dbh7MWf
nk8vny1BpdXZzMn6TGUEImGRybilv4VQpr0ZlSBOBQdKYJTPyOSzMNzNEyhEZ1mOz/vSSJ/U8cHo
0nH2/q9n8uRgpeXoGvxuPp+WCd3QadqoXSHVv+vh575ENkbEKJM6z5QHW67XO7WtL7349Zdw7NZS
tPgk/4BEmDjKpMSoxGkTPeSxiisE6hPvo8Fy8LfwyyFl2ncvIQMMeYU83eiaiYgkcHN/idbz1Z+m
g/6+62R3QHNoQPhG7Q2tZKhJGupqK+MZmR1ae0Ou1wWeAtcOtUjA1AvXQuru4WMUvdAhc4rnQC7v
348MtfkPJAjKSEiCOcrUzs+RAOfzBvOQAUjxtgml0+bgzc8ORXNd6ymitbsAcxFF02IlKGTJJCIf
adlN6jj9YirxKbu1d5bZpajaGQMALR5ne7+7mgoqrxk+oRZ3+3tI4rvd2VLtChaRJ5sLIP45e5bC
vuUojZViL0nHh1Hr/mLjYwKrDrFFPnGqq2+ghgdfhIv96a2XyolObsywNUrOsmpTnxIo2WTqEmzt
UfKcCyW79P0iSiST5PNg51NJdLS/qa5Ne4SrKIx7xXv4/88fJzT93m2ZQ+wJ1Mcj3ZcBZxJi3006
8bJGl42FK8hzga4h0tsM5p2L2LlPa05UNX5TTan8tfRh2KKfVQOZXYBcG6ZX2fj7tUFDTKt3zxqX
lRt803IXQ9wa3qQmuZ0s+17Czwxk5AavcPj25zDJGRWVHRZfPclmmvIOxdK+Y4uC04Gd3+JOIRTJ
P6erM3/6UWWcvkkvLuJ+cckE0lwvqEUVq5h8LvDzu9I0cMS1riZCG+DoY8DU6jK8MxtYnbDCBUB+
Xxhpi/Sm7DqjcTr/XER8xWNRk7d2eTt4zjDrmKRS6mcU+zrcGwEESTzldhF7BNrEs7+SKWto+he+
2S83aOaxtlmfW5GCJlfedMoM3ypTrkPFn2XkL5FXLSpeo5YYHpqgKhG884uLrEqd/Ejdv0p+R68r
WEjJeiIg+hmhdolSCFrEAgvL44mbhDcCeduRHfzHDLzKzk2UhQmNqWPLsiiYy/2ApAoS6oedPcWD
HmF6SEIz3ZCV0BcyUN4lSmRZLAuCrTXMyLSiItDNVRH/7yCXJ8zheBPPk5ho7sgJpunDfU30NfSf
2AdCnTwRewGZOOEg4miG2Gjx9/zxUD8rqK3nqkCch1gZmcOmtD3fKZCbbaya9xd5jehKBipzZUXY
ZbKtjH1m/IKLLmVt3dGOgbKQoeMg0qj2BblRDJnF5ylFgncLS7BTjVWtrbwfAlFMvKi3oVV+UpBv
5K60AfrdNt6hoBYfhQVjGd0iex+ycFxUdhn7LNnBA9wATPRVfUMA2pjFgPP9Wh/pljr3h658PO56
6TWdB3Na2kcE2xVTbDeUBI/UoF/cL6x8iBQsOVvEDE+91VVcWV1+k8KbzJGVq5T1jp3gWXGPyBfj
tJH7pFjMJD5BgoRxx4TkZYNQmI3MJ+Tct8t/d2yK9zDQP0pqRtiQzwmi92wy7qNzWPjKtylrZ6aJ
2F4S5dKNuXhlpBm5Zbo4TdfdZu+49F8uZeMRNSXef+4iDCHQr9PH+QPTunf/b57mm7BZMcjW7o8Y
cwtpZmB7xuYA59vhZ1VLFvGogaQAGzhOAXp13ilYqUPPsbgmEZ1qvpswZIAJRPpAoy8dhtNWVGoh
SYIGC4+H+p6BIqvl0EJ3zOdcD7lC9yTJfVZiJ3eaUEqLTDwljIm+fcXF2Ft2Z7up2j0gCWEFunSA
2+UB5UI0rOj9VM/16gnb+wei0BkjsWMCXsZ7T9sAsRHDMxsTOA+rJ5NOkYJu/3nhrEn95I0Mtqu8
uyyFxBaOxd0hxUjBu+FZROQ1px2K4fnBAdet2bWBhbW7fyIbNZkxYJycTDIRU7fZmtXK5UZ/tIKA
eA4QteunckehJZpKT9SvVQqWeiS5y1HSN8MKL1NdQmfrgwNxzc9WT0Qro9nFIieIjSIgbb1HOo2t
znItyzH+ndyH3ZJo62Jy5BR7Xcyqbl0sECJzM3nLGtbVsYP90Jj5xD5Mn4h/ofdwCBx1Urngo5Xx
rwcz7xv8ISVHqZHQbYkJhuQEfKa7s6qJBGT40JM2CmVm+csJTVw1PslV421rEXq9TWHdHSG13/Vb
hUcMlYagE8CqD8cWOkn/rYSFoVkWZW/6+LZT9rn0ZGfbA6V0So1GYYazMAK3ApRwJigzMLWTfVNi
8GaJEj36xFnHzVM26lq8d3YtULI9MT5O8x9jErsZ4wjFhw4Bll+CtyTnCn9qw/4dNrc9CUBDtuff
XmI5x3IZ8gxPwsW2nHRW216Oqy5xuCyzzFrvY5yhFjdx1lfnf1jlSgx2ROd3eW0ird6LATiuUjg4
3zh9DJPY6bfCeVMdta4DYi0uv0tIBXSSV0PcCmeo0GMhVB9Cw2Ha10EgUfJb/pgDwPxx3DcC24PQ
gI7a1yJDCjWYYuwWi77l8/stJgGJ6b41bvWNPaLq1h/s8Eqcixh7G4piOrco+Q3iaFopa9eto+zF
60t3JZXhleBGodPOijtqhShLBySh94XoFiApTM0QI0f1czKvQeBD2FTkyzTvN91dOe/VNo7cASZc
3oo50yXnsVSZ/h65cQT6BZPMgfbSQjwXblPfni/OjfXTd0Zy7B/06Ofh/7/HJjNYbIvqc4NYpb+5
d0223kDkc9ozGuar2oHFLiqcIyrRj4Vu+hgzZoP6qzPIWUHQcE6fE1iuW2e+bL+DYwcE7eV/57aG
EzTnNa6/5cOHcM3ngiWg8VPZpHADMULKN7WFaUUvejeVf3AQUO4zmauhaGB1MvVx9JW2CePhrPhj
ICdNjcsZAYJxCPAtalW3wHGp5AbRlO0VzDoY/NwI7uDotQP8TN1GcjHOse36ZbBS1jUl3ktS6XCy
XrUTm9sNBuVwupuVykzysX4PCqFZHj7ZNDO1uFnXQm8pPSUoAwHx4Dk9G9CNif4dMjJH64toIxkd
HHP3fv6eYcR+jqoslylfsXnGK86pcVfDQ/KRk9zO/bdC8gTXvC6JDQIYuL4/djLToJlaeGtwa+fB
8TeET+oJ6H7sILKLOmCf5BuXMEfSPoiswbBtVg2zbQbvZHLGYZbPij5cF8aJjLnG3c2FcXa1jNfl
a2gQ5Vpx0OYDU2OlJPaTVt/jCNJbyQocTv/0R/FGFFU6LrG4wRDVwLlDDKZAGhiaT8NEzLziFiwD
lDq+M1/Ve5lYFcA9RbK64NZxv+lmwc79eU/qqyAqarkK/0b6P1U2hmg/vqU47sPHRUwpTvROKbyi
qxFw/X60tL5rZu3MFVEPDf8oOSWCOkoi/pWaYO5bot9Ph/zEDIY12g9rBY/By90OtwPlq2mac2Z8
ciZoPRZFEpvQPgUokycUKzv/NrceNhwrKlsL3Z+08BNvdmHIx82CxIszWV2pubfkmao8l7R17s6K
OO+pNATaEXL4bTZOOhoKM4/eSOh6VJFuW8HoSKDxR8yhpqB1BDZTozcz03PUgEccbbxc84T2806i
63el5RA0MScT+/c5ET4OXfwpZlxR1hT9GZYOOibF0I0wSB7yEjIWX8XQ0fszgmecvEgmLijAfnPB
7KSeX5S6aFFSirLq1uejpbGG51EIE+C7lEWOytnpSVurkfVOfjRhBbnzxEp2eNWGr8gkhmOU2Vhx
qz3P9MmREffdOYnt94oLkM+BpcMwwawgeui4yFBhi9CneNBMqARnL62nMt8Q+kPWFPmTQPZ9h5Fo
KTMcBdc9TNqBlt3ZqwrQJZmUbFfxH+dwAcbqfYUwNzUwHwl5TcW30Z/vE/67RMJSbzfvFvW1sgzo
3M30dPuPnRKK6QlzDc8tVDCsEi3j7JBhWJWuAijGfl1oMU+njyFiIXchgt/Mzd9mBYAkzgFuGUVQ
DLTrmkM1OIcoTQpmgABcPbC8u47SNXSSne0n67J7sJVS+zn2NSoZsNUGrIf7gRb4mvuKXc3Et+wd
2eRWNP6zh/v7HOnk1IMJkFwNAEvzBSmRkxDsnVuTRqkKn7YuTyzuHhqArXXmZp80mOssh9RKD+a2
eMPsea3vBjxs3ifv6e0ee77Ja/XTl6A6oLozVxcLtkPwa8mtSg8zFAR22Riv7vsiB0dUYlm63UxS
+A9mtWJN9gI4gkNV2CkGTG6omvfXnLxnn/2XdVbi3QDHDmf9V/yJmlPjtjZga9ysy8kZ8wb/9aAV
H79/gwONrFjQC/ul5UgfN74Xi+4wOBOoA/S900qoOzEXg4Yjbd4Sy8JISqi/eQFEgqVkh9BMBQZx
EtyyRZWJno7RXRHJM7Ug5OHjrulS1rF/8+mdi0FbARgHq/I7TdTY3qGiqsXTQT0nsRjYRCvjMkSf
mGu/Pj8KvAn7xeact2DOyA9jOkg3PsqV5zv4IdMJI83gdxeeO+4lRyfaA7DUbNk5Pc89S/hErfPW
82pS/j5+mySIPD1AGvEs9sfP4TL4G20R5Il+KlPwI4ePw6l9PG9ncEXSq6WHntwY2qVZiqKzEzRk
KPblSEgbQpxJxUzXSiVIpWJsvE/0CS+2RPI8HBALY6AV393R9l9a/koBq6P/5ZC4bOcsP+pqhFYR
U9j/ag7QXKKsLN4+lbjeB/oMrO0YRPb8ufreO5frtVblA9UOuFESqUiTAvEf0MQx3LYSVR6TNBHR
AZ8/9cWwoYgCoI0aqH9dcgms5qyVEH1soeFbXPIlk0embPK/ZXj/KYDtcAcS8sAUmBf7y5KmG581
C14JSmztVt5xac5UvcNmONJX+CCA8pFwR6NCItOuyIAXpBaqve0lth+jT4dihPN6G3aFg7DBL1S9
XqVIJRjraGSM7gEHcIv9hIBBGOTQaKM/rtx82CunG0MtVcz5Hi/S733YHrlYMgA8aJg4FRUqrQUH
RoNqIv8JphHqPN2LPOAgyw4D3cwvoS19gnimXkSnxODvOqOayT5lPFGS5GqiicN5k/PxgrzeIsLO
ZUWNeMU1vYlAMPbSkyrevnTki+MIfjWjDi8my6enIljR1hvWQpQDEASyewS/uatuNga2jQxqIllF
zgI7LAGd/QMq6/K557L7Hu49NRDz3hRyaTiqFkS0W7yO5skpg2C+z0tUjwl/00EqkaNIP9aOWHbO
tTUw5Ez6hrzrd51adLgLWflfMXkxmYgwlADCxGtB1ZA808oM/4NomFoj/bCxO7HOxAnqNs50/vcF
Uf3/tUXIe9yNygRQPQhDXYT1t/53vv5efkWN5gx9OVW0l35c4TxUt+0M1HBEpGGiP1iG/X+CbUST
J1jhsCKTPoeHYkJjBEGH8JRzIOiLIPqDXuHDLd5JpkVVWsNSMz1vt7YVuw8TPvUi+EIYpO1v6a7q
d9VQYwHZLL36CVTE0l2k1gl1sz7Z3EbUGN8z0bnQVPI9anzk+6OVdO9zZTFBRpMJPIp/C4AzXP9W
21gWRY3DMz/hS91XfOVvkcwa07Jb0FwR4UBeD05+qIXyuAFiUz8emErAssJT+zOSIJyCU8tlh6ce
bsOESaSwuthK5ivNrkV+aktxwp+amJmRZG60vf61Djp6OdbcCK5nEywlUPOUT3TbKAsKVUJUIuN/
xfEIo0cHAphb++VyV9Hi0Q+xaDSGCYWaSau3g+a2mjZ2tcZP4cBAjBSkB+gd429AwvoEVg6rvFOk
FhLp9Lds8pMd5qUXbejdTtxjFq7l5P7xs2qa4NN3YuopYUYhI7rTykiIdL6+n6B9H0nic50GlkNW
eC9EVxx9XN6Z8i2RZZMv02dBWS18Nzr1D7rRrZVE9+qyz3qsS3iRcIU2ipUrHm5xnfdQFqYDgxSp
3VhZc8XxAn1GIA35oPeQcDJ2pXPAxBVBeXyy/ot6xE1LD0uz/BalxMFvC9l+ZynImYLf9xzmLf7f
J0zjPT3ZWr6Vpr136x8JyfDD8hg1FQpLIyqcReOM2wTael0NsZ3nXbmzngSl2HTn0Dzs1+5KMIG0
DkD0NLoSi7cQJ4wUeh9fcmIavFX7bQXXVu2e9XJJRMDD4+RS6kfAEbCq+FmrADq/Xsdu7K93s5Og
omRjVEzh+n9VrtpLGRPWWLXJAuHn4Tv/QbmOLvenOvcK9o4r9+Hsx8Rl12/aYMc64X6tSFJrwuEW
8f1TsXjsmABde0zEb0UQ1fYvKn2bV13rhc6y3NTICKC/4HkonMmZ4zhiiP9c7UHm0G+Q2FyNZLV8
8YqYCsHvsxi2/skrdKtIRFCi+7X0F6ap1ahdLXlprSx4c0Ozy/tXGE/qHJlRi0mVGCx5QmEOExQv
X4mWk7izcDWHcKxxJu/hXS17GSxjNFpvEw1YZkyPZ6UIHqaoF0u914RALIibvJ0kj8keBq+hQJMS
dSp8nYTcP/0wQgzGBKrt7AuVr/iWE1zvwxdNL6sHWYJ9rkJbSETikB7njfyqfzeGGU8LOPBezKWO
xYmT5Ysa3A0H6heUVBCYvkw2DL5crtT0Tyy5lDZZ4BRXBW/gjtmDxAELH9tFe8GMpjNBMafF4sIr
flpet/H/js/ujXSCO56F3hWUlK4W7WFi7UJPYFxf8UVxz9HiUUX0ZaOae9atUl7V8BVOF4CNxvUs
cxcME1pAweA9jlJirvPoHHLrgNaVItH8DBvNy3Hc8leEksJKE1fRIjLTEhpiJfxfnihaddkpn90V
AYs3o3TPM6kwuIWySxawqc/LKkogJq07T+e/knIpTX7XcEejeyAGuQ4r0VdU4uCIonAHB8xnUNd/
IIC2PSRdbHxL2BSYONscCQ6sALYnhcfVPpOTeqtYxTKzsWlLfG+H/PG2go8LwasuLrcBOpjg7MqA
ZXRPxlH+ywt1VfmvxW73j71UtswqTC9F1PI+55HRF1Ckl56fs1FO55zXC+rQ9ztwwb0hLFTe2cFZ
ECcf3y3YJfjzWXJ0i1eIn0obSbe9sDUw4cON5sWoWa/jEzXKT6SrsnLwotXiwnZYQn9NqlYC+S/6
I6zuYrsXvOtdw5sJdPkI2yjYVJIk7A7kcLWSYuyVYQ7oUwt/iIoeigQ/hNHWBj7wMqyQ61dbAf3g
mrC63iUQ1SG2c+TK/CEMuuemdw3spcn2fOKiTAD7UO/c1s86zsPcJLnzSMg2UfZQ2aq9BEx44lO/
uWSQVUtIlbAXaOTSdWBQyJbvex0d4UAXCkoh9bdQw0d9/VA21ntvV/g/mS/ySg1iFAwia7wnmx6J
sg+Q815DI0gBtLg4w/3CCcaT/3k8KjaQnVvB9ROWyuTLdX5E33tpvAnNEE8S4H/u0ssxHShsM8Eg
3v5A4a3PtyF//L3K3MRXQhkbEBoJftULFqb/uRyxgLjxX6Ul9oeXKyuVCYvYz6zv9XJ1kI9d22Kd
Xua7u97DD9kLVFyIJdXFQn7xUJs2/IZv0Wx9eYPzuWmhYJ7EjLxfDoFKE3TQkFmKwbUqqV1dEa6A
THMw1/FBuEqtjfLlIbUXYSaqvdBdugb10/P1eSYoDjfn1I+joNXSRruF6r1JJn5XSRX9RdhjFHe+
sBXu/GXH2fLUco71yXvVljN+anU5sqLhACnyz3MZL++tO3nGQXGAxFNHDGDY9m/g0rdkZjsCwbpY
p70QGTWGb2PncML8hilg/ItHGg7DL7z51RJ9Oa6zAxCKfHLl1bJfID82M5Jv3UyKhW1G13Jn1fhW
AjNCtP63whlqcv0OyogURjMNwOrJAnFMqBGfxheAbbWKx0HVrnIy4zPbl47ud8V362JbZLZn9Xdh
GioRgXmRoOrGotAIlDHTVo5QpZfoNDqqcw0CdzKdy47nuC2A71jmIQvHIb+6UIpgCRsxuUQf3LWN
gZ5K50SYE5Go3y0yW/JUkrg3TDlXn2wHWfTwp+dGyZ47aKK/1//BubAe2f05ZPm1njq3pyrCNr2h
2HrgaY4Ocm1qyBMdKVtNa1GzeY+u2w3gsubApAMmGcKfwNR0Je0HBMRQyaYJodcAyqCcK4Sa6QwA
uA8gDieO7aIgfQngRCgQFpYYC+MdBFsLHLZ6lBRiDxUS9PVoX8HfFPpqzRU+NlDfaMXyXcs1nEL6
gwxe6vs+z0XqLmyscsYUENNWTFnl9exNUMPIdpgp8KhX2uA9O4M+8o5KCX0HJzYft59ZodNOrLiz
qO4KVYVLiwH1D0+cEc+OyikapwyZ+ZSnpZ322nooNWxAVs1jnNGKsoKmSTo4NTLiyYhW7F0Nkc51
rrJplCAKPznXKPZjKC69rUUbkRnChXmDXH7+7xp8Y/lwLW8uzabnaBK9rgVuDGZZ32Ia2GncZQMe
4lVHiQ54tgR0ggEWnOM5wMjzF7Yee1qGoSbQ5yRery/MrYZk7AhxcO1khBqDIQ8E0kbdxoZKt/rb
Y8DKs7CLnWD5LmFhDlKeAYjWAwRJ8LIF/ausEChFZrKttm/C5rNDJKb023ihKfl7RzrNATEXucfb
L9pjZGFVjNrZXh6v3Qgwocz+VlKMKxKksWKuWFSZYe4R5W7s9y7rSFzr56FVIt9z/S0EKt/JNUjb
J8JJNKNZoZb7riFa7LdIm0jxpcTo9xaInPlUnTLXSGfEusuhOPBK3iRouWJCO6YcZlKOq+ZaY31R
INkIJ29UTuuM6R5GVlDDu+WQN9MOkR4AqWeyS1X2t3dtIwei2ROMHQkZlf5Hh5Jpm/fN8Hp5ELfJ
PNGvwIbKVmpR9fW0eOCvs7Uj4c+IGib1M7hD85us+iP6UkKdG9FzeJZEeAv4ObiBwBPCNxY2vrP3
yND53z0oQlIcJBUvF+JAQ9n93s5cg3P0H9PAVSMOx0Puy/QxfhUlvJqYZ57ot6Q++d1XjdwzDAOm
SzgpKYysb1rBl4hw//cBLFLKCkL9FvVZaFFgs1z9h0WGFQJlxH5DGQDDvMKu8G7m+vjLLNkh53xI
XhnTnHVtvD9m9VzJ1IkYTeOmFhLSHu4Ubqv098je9RUe6pm+aj1ix0xW/GBxBEBgNwGkNiv4o2Ax
Kc2NaYCn0iEoR2XqOWltXIa4qUzG/78ZYNsrsPM/yq/FycVUtp3uFxZa0ezrvgKbMVrtW/Q9FCNv
EupfIEb89+U7zniwKurNnm7+C2OGfsCSGMfVRArr/8h8uMmB+Hb6eGD4CqBlDPHMUZS9wYySYYvl
Z56r9XS2GdXaO8g+UUc+fePW4FbiobadzRMV/SZPaghc7gGT7f/FZRVoWEWlDGKdxNUlP7BZH5wE
qVDS/FRyTnDSALAIIyi9SpBH17YjndHkuhKy9sivwfD68ZjhgRKFjsuqa8tw8DRcNKe46PkOLIH4
pmmcGSBj/YvN6wPqgX7RawF0OlieICvEQA0EiKaj6koKj7sASILpJOmaZ0dWxuCLM4FH0R6b94tq
tn8ff8jCwmhVElDE5rvthsyNimVOme+FyOtUjSoTGRp48HpV3fCqV8a7s9aI26UWI+ik/E1mcKSc
09pqR1OHnxewjXIcrbWLDBjkG7BxTmxpivd9M/iVnDQ9q6AR25OwP0Hp/xzRNwtdFeERGsv0Q0uj
BSudFbD5vN6BxgVqgvFbpkep+v64qwMzqavwy2iKZ3M8dgYqQPuxmpMfVeVSu3tV4P2kmgWXqy9f
Clpew6QCt0Yc6arWw7UPzVaWI72wRkpT5jcSxTP/zrln5KdzNsZAzkQws+btMa43yg4qkpV26RuF
xXrRcKtoBN5RCVgadiqdCItBAmVTNokQGX1WiG8yQKmY93X9nGFKnPGzM5nidx64Q6KV8hrb9xft
17He2nVOH8o7Hi3kNzI3QT4YdipH3BzpGWJTaJMUL/qeLlWyzBCUoLAopvTfklTxLNuxfRjoZE3W
tXoRUBknQag2QlFanpJLnuZggGOoPZ9sQw3pIb1UtFKNiRiwviz47/9cGizHIhXFOy66znFyQZtB
1MRORdzROcYXrkTONFzKE68btmSJt9EkGxkN+Fq6IsYZfvop8slonFPl78/iXlgdvPvDMqHHWRr+
6NUGpu89PRsg2Po4poiRzyBFYylSYOW3J56X4NeqJknrKNQp7UR9bUVsTY50oM0bNv1Ga7SMR1nx
HHf7gvelegzxlWCFT19FF5Q81ExpqvI0DL9493vd2grP8Jed5nFygkvs+bWdlBInPB0iy/vli26S
DudnD6lPcHO5eyaW7xmsRxHMhiPZLVAMPSO+J1ENCrU3r10lgKZR0pFvBz0MoWJt5LlN7c/fx85E
uP/gVnTUIxafcouA3oYPhHSiX4vWrVIlHEi3znw8/gdnVrHK456w4fjDciA0qAxu/99zutEmFKVn
RWr2Y4rgpGWLKBg96smYwYZQ5i4IgDC5uSCajO1h6pB2aAjxqWUSPwM5dlv1K7EhoRronk7MXC0k
vD572S2amYCLdefGyjTD4ERJL+B43SLqA/kvKEnqHg3ZHEg4CqXQTneE3SuQO8C/jnIyF0dJVAU7
QPBMw9q2Lrj5SpcFDmrREAq+V/bMAu0h0QcAP9Q9W3UbECTBUbhskDuKycSG4WKSb93eHq10qPYx
ZeFdRII3fPgx1LzLrrFbV/uwiHxL8H5niAQmAnML4sZ+THo+3cOjelrWafm3l4lWhXlvSUTpXcOo
gqQNXTHosjDylu2YoHSZGndeH6mnLD9YFhO01W6YOdAnL3uSTnScVC6uVxjV1FfIQ3e5ELFgK29L
Z6RQpatfeUSgtbRkwpZ9o7WRSpsq7S9M3QzFLwxi905ZkTMpAd+KtzDNg8grH8xyEz+sbxT5CzLG
0CEjyrfJp8krdf+rg3+8EXMjoM10hG0Oa5wVXy94szmq5xWEPq0t7bFZYjHkwPiEhVRcIq5gUtK/
o1v8C0KAq5ie8hnGrQNkvboifzjKxOrsw5f2p5gIgwXO6pYH+5NZWaUdpfq2mpc9rP2dofZal4t3
jGJQs5v+UXZ3oYQxH+hnXvaiGYlYGY+T0qJrYx5QUYF09ievgemks3GkCy5RRqTs1iOGQpyOsniH
HAgIS6i0rEsjlMmu4HM53/80Ofsc0nvsUAReYf/G+nH9TrVjjGt1bY1CJSCaBlbu1LIhVw7qwJpq
nfZm/6kpATZ/M/AcNKUKdzCdrsg0Z9T2bN2hVNCGtrEP2xkUWR3RIOlJR2tZjZnOW2dj6XY3aD2m
CXx+37pGtsxv9ECmjUyHPKtM20nQ57BvW+AzoV+uOdgd64Q1fZO2OLhiPExWWkzFEPJF1D2PTVMO
LWBDLSFefwQN72XMOAFu7aTYh82poZrRlTyV7rvdrp2xPes9Us6RnRVh1r1oGokuI1QMCzxL4Lax
2m831R7UfFk90kjksyJptvx5eshgIhx/zaeaDyJFIid9oxiCXEtZD+N++02x4dwkufJvNDGMi+Aw
1nJfeQ6osjSvHP0L93rwOA5rpuRRBUjgLra/HHYXbxqUIZgopTQaCucm18093VeYjwwX0rq7D3ZJ
ASf/0PxulgICge6yoZcLhyK5LVPx9qWF+/i+MjPUUmiH0b5PkOFQOih8b6uw4NhVk4J549UkKoGQ
kKbQ6rLSpZII08UYFESYJLvcr3b6Bn0NYNJapa3LCU9I8jXHEsCUqZXP+hKyb9RWXtUBXOAiW/1x
SkyaU9F3U6ZXmQ5d3XEQ+cfdtpOMSsjzHBgJSYnF/RTpY3JLhF0YBWWHrb+QvTYtQFHMbmIUxbeR
WWgu1N+kQMqk6zUym5f1CCnn6qFUVQA5pJicit8yVpbAfLh0Q1hPO+2EUpZnmhBTNb/+1kVRLi/r
h23IJK9iqZAgR5nN0kDVbTUUoo6hBBSSO7w0n9WfjBomKR3JMqlqKlssVESc45Smqgf5z9mfOxFQ
G1ipyvKaAePlMZAQwPAy6Ib+5K/enNHAA9Hi1vPh0+n3jo2HfsHxSB/2PdxM3eBBZZQqtT5QVTuP
ZDEe1QcPRGJJ4G8O7MlOGB60AgriDfsPpbNH9iM8pFQ+L+8Qamjqf3DybNset9uxbmOWwikIrGw8
fWFHu/65Vf2exW7vQVHmBApZqCMcz+wmO7jfAJQsJ60anoLjmU6uXk530RSfocbq9GHW3uxvXg94
HEUnZEJRfJM/i1OKbHH4oog+4r8JGEUnsTx2XtHhCEG1jac2jFjSdaHNT4c9EEF3L1rfgE7vbO5O
qLcuJ/C3pq8EzxgRFyh4tdz4pDffZRqvh0SUkrPqX5h9RyQ1IX/BFG3k3cvlN4LPZnl+UFHqsHbP
SWr5lv13GbGUFc9g/klW387ZfCK7bg5N9wW/tInLadywQcyKn+lR9Lhqimv844inY1ga2NCHz6q5
5D3JQvK/6zWL5iT/Lcf0Z/gb9MIxJVzy3up+CU29uEXhYftDfYJ3z6SDP2LoFCtEpay97HsEOmZU
22dHejmTwOXPB+UOiemO+NIu1SX8umUElBa8X6os0H3qq8zsXmiVnhQ+JdOa1sbLluAR2u+Q1BRB
JiRZ2gt+82dAvS3GToKBuKiSm0ItsfnV194/Ht2xFVFp93r1t7mZcwF7+nn8y3OxKMrlBm+J+79G
v8lQ6pRurWjWzzrsfzQQ58NNkqFQoOmcvaBTY4Ueqcq6uGbSMWM05Uz1Lt14SwTLUSCG9/B833fb
IFU1hAoG+5yYSPNvg4V09ayek/Om8n9h50avczozBGO6fCKBVVFioPXZwElFnnLe7Juaqqpat648
9REvaiaVMrWhWkcS1xjAU+F5DQxoxLCtskBfCRZVHDJIttHb1pMAfiU3fGC9tvpLsHVeRo4BAmJ3
p7PYJ0EvUOoeTGghuoX1yWdFPk15+4yXxN06IL7TBosqKmi/GvhVE/OKBjWKqaROcbB7DFGtjTf8
krcsXC2ecZh++9dcdPvfTDb13vMvOnnCiyE0XBc5+iQdbnUfEePHmTjKi7A8xkEN8U9uWah9F8LZ
Y29N9Hphk0+SiBSI9hGGzQTp+QrBFC3JpKDpomCO361F3qeOHOc0xVLnKhYCgrCqx/S02D+wch4J
Pb+Hy/hat7fiCYa5nOlvf47nWy1zBGq7QIqEXE8Abw3Tj3RDGaLCYmdyzgQIRGGhTxLsaFZj3SNS
hrEqeFSKpQvvHlpw5MlXK95E+LhDJjTRLOCGBzCGAHlohAGbTu9/sD6wtBqHyYmSMOmBFx97JCXt
M5dSwuemQ3nPPH73ZL2mKX8/KwvpwSQ88xZ38OdlzB6LaFBzquq8Xu8YQ6vKRTvyYUEPwOFv+QD+
3Cec93NJVN6EB4gQo6A+ryt20d65Tl7n/igYxzlCzoENbPnHg4yoBTvB0GtAMLIZxYo7ae0QTtHb
gEIa3B9NGAGlFVEVoH/sAIzVsw5NyzPiTKeNHuhrkIUa0cBQYvEcPDXmcqr24oxXBNh7wM2xASxV
+Ij1hzcnM76+WQNWhQZDPsj5ungTbTdbVYLfPUP8dl0fpCU7hL0fbXwyu5B+kNr7O/72bnuWKnyW
bXlLr37y5m2MBwVR1v9ezB9XPBCtkBvJi5dX4gABz1h7wB7UPyrLNPxNoPNHoAkI5FzRCvLb7kh8
EiVOJojNu74NNfCnb0otQmKmLzE029YcKuYZwbPl0ILPfpaTcMMz+bLKoufTVS2OqpBghrxPHaxZ
KMedFQb7nW6APTIFwvHN7wNA7UfZST2Q4AE7J+a9DudnYF57wrSmPt/cp+eSsfata1c6AoDwJ3EL
Yn/B6wd6LWgb4vwnsRPmAUgdvsrb0cb1murUspYMCoGNB1mAMQJuYfQFuEyebu1IWHs0DoprBvzW
XWHJQuEEgeIQJiv//NGoEkcEXC+1I8wkjJhV+fKkcGm0jsmk7DHfGmDORpg+dKXQIWyy1mO/oDUP
XHaMZmSh9TeX4ObLm6Fm+u0y6mahpjo4vJHgiF97vpVlAKZlq4Ws9ua/tUvaqiikvwC7j6Hgx4o/
5zqpCgiwJPQFWwIRNchE9gufZR0QRvDGaMT7b+76huxo98uhQ1289rosvZs45VlmMoDEJNblJpWy
7WqQeN6E3h2NRiceOzLFT22JxyOCI2IoIvDf5kFzMj23x0NvxjJU6NV1D51NARxuLyGza+D61R+o
binufuI3qUBeG64bvBkc+pRiyK/EGRInf3eTjArJPRzGwVCEma0C+syg5ypIrT6UFAZJj0mrX+oB
gudmWpSMviO4H7Gvy6y5KdAneOnJVwo2TISO+fmJRhLbAgyFNaSd1YLzr8K4xnPZFpY/r/3iZ/9L
eRCvlBeCHGLehs+2PzynkJHbhtaR7D/hgRi7qYOH/GYCmQ5XXAEzJIHzTKW2Lel8l6NUdnqaWXDY
wCUQCUnIPHaEzv9q+g4i1DUmpSkYd45OTol0gkQ2Z7o6Fvskhbz+J1bfAy5S3RGp5QZqdXt/cRiG
BA3o4TP12rWawCgkgeK6F0OtxlmlmxTA+x5s0z21SJ7C1w+5iz95fcDBkcxw2/KzAU7pI19nPUoo
a31o7wyYGa6/nVi1aMtJn+BMiT+q2TKTo6xmHyQ2pT9poEm81rUNsamlqyDdb8dlmKtUZz0NhnjQ
oiAOIUt7UNnzvcUPRmuW5LFjwcJCVN3Hy16gEhgTpWH19NzfY4SHW7cSOPnPGrGS0aoDLZaW64Gb
HO1PRx2doIlI+JmSn/y9mRjdXprvfWY0K6TFqOoKwg6vNgFopzh7OGzYSexJnb2/o3HwRn7y1bD/
vsdYdy6NHMKXM0vjFLEdB0KLpvbEGu0V2IDd+lSuorkMKbxbHXP+l+jW7XWrsULnUZmke5gJGzOk
BDddJEKY3OyO1nEmJqazbs8DfVyJa/QVAp/BHVvUY8gTTIgxSerNpL5jtFRiW2EI6VFpD+0xydi9
55lg7FGQZLm/FwRJ56UXF41I6E0yUOgoSsKaAnaZq6l9KDvgO/smQxpH+W/avrzpUo8u9p2CNjgY
09MOAcK1Worq02w2RN3qe4G8p4v5IfpYbxVKvYbgioBdTzZi6UZxN+omMO9uVQmfEfmxZq7FpKrF
eAF026uDdhwO8DuWXqnel4XPy7DkIDGG6Uag2TPL3x5V/9eJk3kUrAVviCdDDIL30e6cENWAZiwY
oxEA+OwG5mLTTP3YeYSXmdXAKbir4lMAy/4EYZwNMcaw+Fb3h7BIj+9t20svy1xcA6oVs93P3J/m
wd2GNdU6EaQKyo4s8uiTRlLcHfqqBB0lp/A7Dz6b8sxfbttP2nqTT3thQERPKUJEshQGk39c08cX
QMoT2bdkquKAzLSHmh/yvgj9QEOv9TWtNsGsxqtbxAGUPmCds6EmZzUVgvzhYyNnk+UnZff5Ycch
pnvNqlYqObV12obombv8qBnR1TLMLoBy8eh1yV4KdeXmA4uELacS/mb+TsGcDygkDRpdPXp9H6uM
wdLpX7cTWnteEXvJomWgxLNmNjnvltaCDO7t5okXMsPCmM5JuNMdHq27dxqcOhYipUvIvEIQOX3L
uq0AI224aZKJyWLVgELgqjUyS+b1hQdaegykShB99LjUmw3cn0ttitRnVHpLmDtd6OdjNXIHAdut
ARn+3dflzTChV6U5lJgirLxtiEfHNQG8iYbeoJBdF7hCZrTOTnbaiGdQuQvdEMoqe5xqSVB0+cyQ
yS8x7FhkS/7SmoE6jr2CJkjyHgEpjYI0mEl/6cWge0F/N40oRDNayd0zCwj/VLMCq+/rKqHL2RTx
vmyMbdc035PDsyYWmR0VsMugBOHCzuXMtYpNzLLYuwV7LxTXLB8lh09pfkGIDgYrChFKYazhe4m+
T+qaiTnFqZWTbyYMdLzyVUKL7mtWmOYhmUSpzPonrkvAUjobYfAeXRuEu1DYAKknjlhURqk6t7I0
x5WiVOo4HboF8NAcBMA2qiQVcqQN38V8JQ/JhbkelY5K8+XXtxcXSo/9MQ328lqTkS02WIOVnpyz
NFPFnGKWiYeG3BkYPYi1/AJ72NICZKwmldU7yNMbl8cv9wnXA/1r0Mq1SWy9H2i+VpXPdX3K4Btk
ggr29m28ige7+iC5LiCIIQrvCn9dXK83jYQM4apx0Si2CBJV5y+9oHpwEfSRJh9vkKcFABxJcWJu
FFEwylQKatdYGe7+EWQR+p4p8ZeFdWGGJhbil3i32f4qatHPclwpVZ/xQ74cxiJqhTVQZZEYYvcW
bvQcPGjxZSTVXCiWbHFMKHYmz+OsMBsWUDBqiPTnhwgaF9kHq1ycB8OWxM/CgZ/kvyu/Tqs6lnhg
4JEq4A4+kQbhm/hXBs74XJYPg1gd34idJr1+xRkiu7OiATqWhPd9nHoRSbWHWwQOJ18TAQA6MDe4
gDQGut9PwOOb/nm34Sw9cWoFH1Ptw8GR3Wkl/8ICrO7ID/KleLBnyUHzk3GHGONif/gWSfjksYuT
vVyXGxc1YhV+a7KFqCzJ94E6mezl9dou0CwxUGIDpa2CVUZ1xXn20+ilM9MAuvYvKPMbdjGtTdzo
ZoZpa88rng40hmur3/y6X1ueR8vjDnYXQnON/+SVcPcEVT6r6cT+W6hnScLa1QJ35hsr9qQkH5wt
3ZlsaFKMZa5rRsfcsmHzYM8plYSYwD4GLdYTy/LyoqA48S3xYCjFzfZjwzlp0iObnb/PbNAx+tQC
GZcGEKyi/joLP6p8aX/Id3MyXaMIPXChzMTHNhwm6WfqWq1B5aTxNqU+BEfJaDqEZXR+1Yc6R5XE
5TNrl8q2tDSgM1ee6d0iNMoIsDGZeshiKBeW/bbT6lJPDYgeJ0Jxgqd0G3gCdaWM74eF8BWU8FuU
m2Hs89CNO25d9MCHNW6HdcWJRA0voAn7nr4ozssz4AyzKvneW3nfSz79p6jwtUZj2geDeYMXw6Zb
deoyK0Nvxv/O8cQNh7AKcT539espmDBqwi83vnXzY2kZu9ru+QnO0uXWeNDDCuiFI5bB4YS7+3ir
LNEzvLa5IpKeI7oLQ9+0paUR+121fpeeohUZ2MntlE6uNMbVoA0BnmJcm55RDVbMRn3cQfaI81qL
Gv7+9702LmaLpmyIs2KtDONces8OmPF3K96aG/fQISoUZmv7y6SsSjhYWaghRP1hisO5OjOO1RAC
lcBa3nhp3a/BQN7AEI5X5F/ReoUU7MOc3rMiPxx0uVjxWrpVYOc/Hv3Avj6pO/mCkXlwjXq9SFBc
x9Rd3C7mm/OAzywgHNXQ0uhfR05SqFjNdJGd/tYMoMN4rUDPiBUn2gpBArtxJa9FG3aMly3bJ/Xu
9pK55Ab4Q61wQOutkkSqnC94FycrZ3Usm4+cPjUDYOkiCgFwVVAHZq99I+4FWNtm0hF9dmiBSaNh
nIUirkKGaOu6gBRt4mCJms/guLVhsZtr5SPhFCsFfTkCV3nvUA07kcebihc+F+3g2GLhqqMSrvJf
ebLTK1UtdX5xKnUjf9cczJQGMx0X3rzGKRCBdr0gS8aqelfeNPLqhiw/DKw9Pnaw2Ls8bpGwJckG
SYIiwuvUgqmRuT0u/4PbYih0jJidAHQgxbwXLDIEuBBzatePk9tZhNbmGxUDnEeSVbxybLKcbcLZ
FRd5CIJolShaqJp2y/efrb9sZ6aksdpe/JFl5WDrpk6tMY9SkSlfg0kxwntqwsXTt/GUa9eZLwEi
5MSq6xDe1X10ZOwEHZ1bL0PZoiekYtgHrK+oLYVbj7+/ILfaZBXdbtfiNIV2UGpiMOC05Mg6eB3e
UKKm16DTZuWXhsQ/i2fk9VoJMpNZravbIdyhqD3th2DgHzQPOhJmMcLSu0Wg8xRliL+BwamLGc3X
csOTBHEHG7kiqGfZtA2ly0uIABJ9l1UWzLWjp6mk+AxGQOxmsYCjL0ce+Std9921qQAov8pH1rAJ
Z7YR+tKmqAmClFP2GR8JnVMOIyWrnrCbXR7MpvC+3PvCLJn/m11yhv1280GD0GoHQPVF7RYH08bg
uOlLVpi82dq5NYYxCVoZd1pNj8ySLRpUftO+9nQTl70PhvSl03qp5jxcAZSv5WPoyJHw0HeVhsao
r1D7y9ziW3Wul352oHkUY1XU20f2X/H678V0N9xiS51rB0N2KlPQ0VOn29sFWrApG3qNDbRSce2Z
HtNnfervG3Gs9zGPOu9FavTP45u2xYHLwhQTCrwHAkKXvcNjNK6L41FbAdOeLqd1KYFp22rpALw6
fZ02uJuBm7GIRa6bzlToWXBvJX9Ok0UZXvNYZOKv3R4X3V2/6FttVajkLrlhXaJczAP6FsSTF90W
Q2eZAqmayC+xxnPYNlL07lgEwGCUVm/pd7ifCosQiMp4Mx4k1kQodtiM1fOTRugNqS5aCxn0yltS
nfaGVzVCqex7B2p3mwdDw0t6wKoF0lbjwDfaEwyV57r2qAWKzRfLt9ovMvbb03hwkPHGoXwmYBsd
8MZuUbcD0Qxdw91bCPsbUxkSU4FQC7ytSZQry4mHYf0m5a2FEV7oiX/dn6/eGiCWN/m2d0x27QKk
blacV1ulfFmL7ekiJuvKoF1VpvODrItwLtr+QeacDZJ7FXjtuyMIODIjfXZYPGtnZc+Bht2CPySf
v/yD1ZBInOnhokss/2+BbOu20+kqh2bJ4h6EoQlNDR7Zv4x8RMxroQ0fWnMA+sUt/TA1OhzNlg/4
r7Cx6kjPApp/d+DSNtKhXaq+IJzr/JLlv5c70GITeov47+dFQ/ezm5xadZ7W4jB4P1HMtCQAK3Ar
o3jXccViNFpauGkqGVxMUth8a8w/gbHerDNRkkAjuC1VojmJ9oB7fnYaUuwku3u+aJGaStUhS5aI
bN910LQnjyg+ZzwxHulesxTtSVUHVJzc6BwuUlNazEa4QGT1C2kAoK2FRnDQq/mqfD6sZTSQNMnW
CNey6dzdJzO2Qk89wXoqA6+6W4ok2pdOjROye6Zo3y5/cx5L0v8kSd6SefEuDrvLG8XxK79suBdi
TQtg53Fi5ZtsgEWfaTajj0eohQpSP988yPPNgWy6cjDfkrsyh83raezPP4VgUyxrIr56rKOLZohq
5zSZkm1GKeKh0cMja6J7W+glIgMWW9AHafLW9F1m0WWg5JhY6B4VAAkxKvJkWDo8Z38rtDE8WkLq
fvJYYcb+Uudv3j9s22jphfvBmGqaThzaHpCqhSbL3KyxACPif3AIxqfRl0Ued3ye8jiovva12mQy
4Rv90wReVMolZ7gvtD4EdP3s6lZW4MUHDrpvzpxLPFsKfs90eNkrL+Ky5shTWwS6q0C/qAasgqzR
Iul3wxg/BVoR21zbB111BIC9VXySqpP1j5REtpfw28a5fAobGOU4XqBVTRsZYAgk/7gYx2BfFIbq
qOnXcDBQz/dmY+exp6dMWZcyCJfduojAZ7sRBIWgq9LeaEX8Tu7P8dh41otaXHdqmFTu5xw7K+Li
fbF/eVTC+jiLFQS5eQFjGDLEqwOHNZ8F2z1MIvddUid8L/570NKbUVwdY5Ji2FfOEHQcekoyKNOg
2W+vdA4Uz4hvbLiXP4+xJkxuagQIFlUCJSflvd5HhYIrpvWbYt8Hjilid+eIExncl0EKbVw+NIRo
dFTJmxGkRWM5vXAAtpjG58ks6aZczbStklt4KOJ1Ng9C4uAh69shh3NBAbZa9JqoaQMNJi2BoF9i
EiZ+HrNoX6i5lXJ30lA4Y3uJekWkgyFlaYaWIM/QjS4IzKNXFJKrtTdltTlBL6nIfV+OpOffyCNU
DOqBATDab0WzLUSgNwMs43q1JfDmsNCNGJzS1duigYTGqehaHH5viwhVL4E0taCNXpGzT9m7Uwkd
UBuzwyuaBfCW9spU3axUAvj7QViv0jcnPtwgJM/t0kEFKgOooUayeuNuVJp0Vxcof/J+/IOKQrZC
Xt/F1xTnzF/h9DK7n6Al9I51d/FdaPSm1bX3Xt0RbuIwd/n9bZWXzBcMJw6f+ZE/9J5qsHArXlXC
3kr58VRbIODksXD5NNuADcVC5WisOoKTCPqdKJUl2T0w+e74GP0LQHW8PV5YyYRC5TqIzv/84GD4
zUgBa5aOCWfidcnq1Lm7S326jdRoWX0T0+RPretIZO+LsylfHJLzpZ1EGI6TiKzCcbjZ2VBmIb4O
7xrd6OujeCchEy1VQO0Jq+oxquXV5MgmJ68N9sMwa56OU17ZaEfaeOtN1XKDK1jGUxwpSNgM8CRM
xweUPJGZSUMaTeC5EzxXa7lLYEKwUYutOG52onBrp4dyAs7J3UWdhUlXisncBsuIxilStXEwtqHI
Ldy6+c1mDNMBKUL2N1xsNdfof0Ay1mRwCAua/JP1qoPX/07Lgd7INtvtg5NH7yetajqQM2I0TefM
MEgO7lP3zqQRN93vTiAAlq1+T33sh5KhUXQYNSgOMFLCix6rLYkLaLy5iuW51C9cMp5C/EL3b5Te
gThyPPDIJL9xpg+j2rspmKbscbcUrDV1zyroYu72HRjZhM26SKCUzlOF0WgGwo3alLPSXNujQKTQ
ky4hW3wIuS30Nbjek74l4uhYSYnSFbuVSqNI2a1eQwSNGb+ajaNiPd965ocaRF7cBvQ+kZ2eHs3e
AW4Zr29udCEz2HKze1fFXRbh3sJ93OpXoY1JL1ZLiiH9U++g7BKnAJRfMYysl1zQ50i2l3ez+FJy
vUeDHOFLfLuCzWkOd/UaenqI5LAZzDSmbtwF/uFuqh9FJRA7w194G7Fgy8Mne4iPFcIZlEnfgKFK
KFJj7DIDjj6O3/8rWUdSlkKhjeZj3zOlVi64wPip5cMXPmoW/Do9zC3GgeenwnxtnT3zmqcyvgnR
MR2R935p+dS2rYT/PelX/UNGlSUC3WT3nLc6Iy1mYQxSJV+SOUv1DEwi7sO1RXyriVdOARe8lICw
Nl5wKQd1ddpTwvUTgPGiuTGQGsfmDn9S4TXqFr5QdYLqoyP0HB03Vo6invZefNQroDxI8d+3STv2
pjrzegC5n0XWCHzQv6XyhzPBqzAnIfnQwJeQHJp0Pk4HgTw2/7HQENDFXVf6z3KT456QJnHKKsCu
RFsUeX//J5NfTWVQ8ZJCfncH60B+HB3Z/zhhjEbGUiJze57d8ervulm818Mua832t+VyiN0gi7Aq
g3PvS8iyIoRCka/0fEEjxj2sjWzR1SqzO/EWGJkhU7KDKaFNFzd9GlR4C156HGMBaRMXyMq/0TxD
8ztPoDvk6u7q9buWFw3fmAFy3DpsHNJWEMKs9gaBQoGM8Q2gSDlOWhkhmXaTQ13CmQ/5GtVM3aQX
jD7hia5oIYm5TeHu4A/bF5YPH2TllNhlntGOVStdjTQSkAsXkRe86a5oIjnrKnySUOTaNlKY0Te1
pb6HMuQpCL8tC3twwxFjaBLbGgKLcLMU+WykWHqdOXNxmH1zRf8kpPFvxpYx2KQ6EXmi5hYPc6rF
618EAqLobVYxiqBF/KX/yuVotTsLB8PUautfpMZhOvJ1GH5JERYuA3xtFPxduKB34oH0SwyyF5IN
6jK85i8bdqNr8jD0Le0i885H+qSLxO73YOPIIy/5RdHHDEAav4gjjgkuvegx/nCNuy0vOF3SIhDT
ym+ZwDx/mcL3WOuNkyJUIbJx4vS7C77HsoJ3cify8HcNpCBpgf6XAGTkAqvsAxP5biPe+FtC1FMX
ajDyLqVu0yApg1VZocTKmZHs6UswEcY0ULdcUuD6RjgUkT5mltLXAcXybDOJyKR5CItp4QMa/oGj
VbVrlx5k1VP/gfO0PhoFL5awUCF70qWHLMxayiJLrp3QY9Sv/us3o/+esYjyK0GjzNnUMxMQ5x5Z
FP5lxSase+jwBtf8PdimSTzemzL7z1fEUZkhDG4vHE/QX7iTyTj8TINRaow9t7AS1s5GX1G3/HVi
Fqs6YrueLXci+yKOVkh857o5OJWruiwFhHhuo5FLyA3fKWbaqHXZOTYNh2Dg3uHu/PbomZAJSTv9
1bcaARrVvkpza9a3bKyoCc3ItjtXas4MquMcaTJcpjmlDUU0KVCtgG3rSis+WsVL/N7ogUf/QIOK
EKXx1/xqisGctIKTb5Sw4LhResbIdv6SGoQoGekdlOUwRlIFtpahvwDrRmWjtJZWlBkpjNn1BSwv
xiF/1mKYLSSWZDLIMlMuAwzSBJNnXO0aYAq6dDnyr0xW/iPDaupjXxBpRN9FRyOPAjgNcElAMuT9
51hOjY1eyvzEjlP3uuSJ5ZR0dbCnY8PyrFgp4oW5tAniZY9D2u/UglIUhWPKT4mIya4cxlkLvYK3
MOVu3aaPoCf4fXadDAbXmnidTcJoIBxtOlFqs8dBbusdZ0TQL27OB7MMG/FaGSD/LprIiTYPtpdH
L1OQUAwnK1v6P7KEYOTjnqiRrJAPS6UiYgi/8S01HrlfGTjEUu/zZdgmF9x6EHrdRvmCTLFSFBka
d3lLkkOrHp+DxF7tc0E9hl7v/3JwuQ3QAMa62qc1gpuxUa7zT/3v0hzImDJ1/Xj6RbbjFj+45nQV
rB+8ivF8R8Z0hPaGU1Fc0wOSZuxOjKRO/cMpwwByy0yC8As/C3sxFTmEKzaSKpxZl8nv1m2d7boT
F/Y6Ais8BZTQSH0cta5/YSHziN9Hpy2uk6IYkop5h0I91wqJ0nU7q9ql5ScxfhLPlbBgAsOjeoH3
cA6WPXetwcg+ssLkrHGcEKp5nNrSA5GDG8lmtSG5KJFdIqGKfmV0keTlgQaBFrO9kCUcFzNDbiOn
i6XXdmhhn3n8SSxhSR7sTzs8bBS+Opv2cDHuUVoYUDwd7Yqt8rFIuGMum7Ojurjkrz0G42SN/Q2E
xl9NhTklAV0uVl1UCj8PfUDChS52zpx9EyH0M6BALsi5kLu6lr5Xp1+U8A74enEsqGPQ61zD44ik
/5qoYXmb0/qtbN4L90Hu1U/fylbSYjD9gtKb3TjttERo8cbZmdx6hFlxmN2gGzUHvrVl6/p9PAjA
W6goYTIHyhpq8adTgglm1p2Z5TrRrIgOGf4TZZr6nyONkE61iuDgiXrKIwMnfbw030yzaUDFoK+U
gFN3xRc08W11edfO4h/AcoNSOdtDyRRYypVMdGF6o1CWlpbLdlWXmGYElhmcpJe+8SO9rBfeWGm2
o9bNtnGw7z5K+LKf6u+Wuk2w0ePdzKJRWK2mlzoy2owi5I/7BPJgAEUx625DwKy9L4+pUvxDXtqK
A12ohd3/0VynORELILCWdKicTe/yJeWeUcpR+17CZjNIcfwS2TSUKrQfiyGoMTgQBqevLvWgCUuu
4BLB2p3BOcXzrBdItyZ1e3hZnibKXM1AqCPHBqgeOXBewqoWWETGmSlzXFumutcgKcK/UmtaUyFT
R2hYWv3/x7FdwY8w7CUW23bh8LqWldSzu49VeAOuzGeidVRnhJdDMo7LtAmftwN8VAskzj8AhIKF
FmAuOnTvMj8O1QCXtiIF18G3korbiDrd6s9/N9wEiBbwZlIYRG7mcbdBdt0N2QV5y0RdKNbKwTnQ
4YKHdv5c7IVk7KliXL+05gcEjq6vWM+ltwc0CqymZccDclYJ8te5bFBbjjJXPBlQ0JgBhfOyOC/f
aJwyX5WkgsC9kkIk6Qz6BiWAp/3MkcOk6U54ETbtsQrsj8PHgm7BGQt0crgf81Ph7OAG6Na4t6OI
YN5bQsFlBGgNpCaVZemWHX1rLt6ybaY7ov+C3guvH/JwvZgjGn6/gSnzUkYty8Ss3vTOJXcuG6C2
KHiCnsmEhIO3K957OGzVoQ9PMAH2YMsdVzb7SaNA6uSGplYl6lWl9j2WgddVe40hRlN0nTaBYJto
NNphWtOYYvhbIW7rtepLy5um06obcPQ7gIDZEaYZGNwaGmHmgDtzUzezL78nwZ/WHX+lcOCUFab1
hEL0FOxJtCxmS5TnY+DJsgzv5FJ6wrnORd7eFRF0cHHRmCr8cHI6ecRgka6SzYHo6tM2oLq9guNX
oy7I2M4V7YguG5UoZQcm9t5O/iTdPXffUVzUQ1Tw7y/bctMePiWFxJFq9QYcCnNmAxPhVz/zBoAY
DI9cDPVefhpxRzJlJGHgkS2k+VQOA9ufCWM+wEa5viEIeaFGhF4Ext8G7SlJ+CU6RTI7djxMRAtb
MSIdAhtHC83yxXtMjjoAAr6zX0rQVHJRojnSnoWM/Jb3wAI+Q6QQVemg/6oBY/mN7PslSsFK00qd
NjuiYGRGzA2wnn0KpUjOCO1DmbQLxdg82DAxIx1Aumw+Ca1xLUykfQVCJzlCezOfnsREV4MiiRuW
wCEYOKsHGFTuqQQBalVusyAKckKky/dRDegsGVb57lbvYQGoHEhBOMwQ1+pobOchyfD0Nhk2aGSx
GQcLNGAIVsIFtNz0WupX9+G4A2WwrD+Fxu0lt42AQ0Ue6Eb4B1Jm3JlwmvacWNgTuiQQ5XvvHvvt
i2P3fNmOLrIPyWBqcm788c33TelEomlJIS6SEf2ula2z74Dz0CU3bdOXrfLqe6yutv6cDq0ySUMc
ZN2kt2XzH/IU+npD948LO4aKsGIE6buPcO8E1IwqPv6Gws2N8yyWiNITbwq+ZWrhd7VwwBVuGoi/
La9BFLgILU7Qw0kb4aEcwELQH7oJommIG4WyvM63iK9BePp1m+H1DVOVzxV5y5qw24S+ae9+XoRw
8zh284w1T1D7HPtXtWNE4Ff0QiJo7xop2p2r1rOg8+r4X+r3CmTO2MWKw4P38+OSkbVsOWoJSEaA
BTvWgTRUpZfnhwFWq1wm1EnBArGnHrpdxIs67pCWSJ9lz73bJJtGPAxMJaiz9kYkAb8H80mfOzck
DhhH0iAUaGUWc2I542aipSZX745AXJQNkFx4hLEcyFHPQOSOu17v5buAY1xgv0z05fg4a0PYciK5
Cf677aEtS7TrQ+J+CHzsuKrnd6QY+X0TAKbc6jdqoJdLDXgd/9XNOUHKFiLUU158t8sVxp+XPnDz
D2hULN3Mmxe4whawtkOCtZaNIu5ldnmNh6t60f8cUyc0GOHAGngIUXTrfmGPfwc+e5rC+XQpQJg9
qDRABMW5eIrKq9HzfWSErJtOLYbD3BnP3CjY/mtONoWTdCO+eb3uzT26EFKj2rJxXGbUcfjnMDQx
4ZGdwphhTyeZ6It6evUm0+1E2S+R+IErwIxmGkX8FXtOpV0sotF+c0dUIcPwOPUtfwQNumVW+r+F
tywrP36ovfWgTDuctoSIwKA+4YH2oOQz6mrZFqKSlPFzuZn7P08qrJCAm2oMSKr/xOIK7JbV3hX2
vPDvL384OSS0appT42EaHqN05eQrYkYwfzVcKTWJpDqAItUFj2kFmfGk82BC3jPKf2awsmuGjeHI
fZ9nQpSeeDDxNvZ3ZaC2eDjS4U5eS2gom3U9p54+Gf1kVEnSxqRywvWbNTS/x6V7rb+Mr9a/ZmFz
jNnNZF8a8hI+FzOVkzrGzxFkDHy78X6vt9lSn4MPX/aaKTSOury9qnh1D8HtYk+cG5fgX/lO79aA
Tg8li6po4IeE2EiGKhy38IE5i33Q+dlocdoMZtq5GObUNJ3uuGuse9oabJmo9VVLXYrBhCUeFnxZ
R5z1G7HI2wEX87kUG3PuK25puur8k41GLq55q9jag56C77R3cuMBA9oqoisxlGu3zvPO8bEE82UG
wy5tgrkncJYS3EyR81c16Trffqu7irrZZMz6h/a216SmyJBj/KAWEu43/x0yn5+BMOs9RRR/ObIM
niG/LNIOA2ghzameCNeG+1+i3w+RLoadEnK0vbHok92jTsRVlVhee+EdppTivPSRxplXX9RMOtU5
rMdkiSNJqFk9dSGdRchdCUcDGOmYRAX9Axv5s+YzluD7angjL49QpQuExi2jraMrGnsbZXcj9KwK
03Yism64Sy0DeermdHPwTpJegC1gZkSbkdSQVnznli2K11AvPu4zJuOScapOPhAF+k5JtNFDYNoY
jQQGGT/FOyuS40LRCUtfsx1SzErcq1hEy8sZwVCHgXmCFkICZuIXKOSl5O9sKYLPwoKmC1A4xuDd
9qDWn8V44oBvd7at17zSB1J4iYZHikB5BujC+KR1i+z7sbBxW8ZwjO8Fmr9v6IEMaXfItGWz4be8
biQ2IJIeQUOoaYaL0ABAxsRCiECqEE3+s+MlzEeUdSo2wpHgIJ/wGbIEfAsJ4ShxOoeL0IGwuus5
u8ApWZ024MtqakX0KRJKJSB7EDyJ5XeOhkTBQutmWlFde9Yb2pniHr8v6J72oZnZ4tn+gqwEyTV1
sWes2XnroldKqTBQ+cv/Nw/dlxjRXA6dEt6Qb3NuipIqMSuQ7eg+kEESsJcfy8isAmainZpfCN8D
6gqAzImUGdqjC/6e699L7xFx1nKybnZrhirYcE9kPnQZ8Ni/ePqqEEH1NQjdNk7k4dQt6FC5GG9O
otnRvs0/u8YUq0M2IKkc2a+pQw0ckiawL4IFxHD+7cr//A+fSLzBlPyTNQCy2JuH2GJQmzgUo/ZE
5J+0uBLA0nTFYYbrhSzwO2CJp9lXvN3q0Zxc93vtRKYec3x4CdiE+p3bMjrh+hJOLlZHOYYLCvRT
/V3Y3Ix1BbDAfINg+vGNSQvCIpJhqVqqFymTyF8+/F7Miaj6pQkakLyuXd0nRSt3F0ynIFWQyClH
khSBtTN352GZuB8OdWb6hN5NSNHJmWPxpPncXpZv7afxq3yzeX08cG+JwXas5IQfDweQmRsLOB6w
Lz9On5xGpaCYMKAbba6uvzgxlYVFnhnY5xnp8ma7RBonPJfwtAsMQueX+3kcv0HwNmW5djPYy7Cb
1LBisVfobrXcz74LTW/3QS1zlSljqUX7Euz2QBDittjfV0EFa/ID/ioQ3OmjybWXG1u+4hqCKyTo
EiMs00YprkYRPf1gl4Shn0NaZ1v24MmsUDZClTrF1BZtXiLL02lyCm+geKQkGtOXWZsVoD0y57r+
bSSXg5fYZ+mSn8JRYA4tTsIi5UFNhjREKtv2ycfjEXxg+41midxk7DUz/rmFloUDcSsL5Zoj5oyp
OR/NfbIiHliLTuTz2Xwpf0CpDp3+J7ha2THvsD7gHF4cxAaabG/ed9bsxV6JckWif2CcD153G1Q9
zm8LjBWsyeFlViLmfw/1pBBGqy7bOxJ7/XHetcC6QnqhHwTJAnIneM8bRBOtlaJFqrrHVrvgcvBr
LfMUH1Kyk8hE2a5o3ViMBcuy4auhAhJy+LLWf6mokFJyMWOStP2/GuFRqtupVSO5zFQtFe8bJMV7
abUMHzXa8Gg+mxO5fje8xQpw0ifeQ7xYTfegmpXo7AcKS8GEX9CLJQE65UA4Rxsf0iW9hPFK10Ym
0o1BAkzT3OXE0fcRpmoce0UBPZ33YZnjKAwe3mk6ywZP8HHQJxOxcVP5DqjMA+kGz1vTGyq4sIpH
AGtTksPVsp1zqR3o/hoEUCeGGIGL7AgejRyc5ioO6vPftHFN59wairLvepUvGikhw/mHFWkfcENL
emXaCr10iFvwcshry3F2dK6Y6jx53p2L5k9CW49MtI2dYUehlalNScPei03eP3iETjiAgS4Xxppk
+pk+ASDJDSWQODyvj58CWArvdJr5gu40ARCfkI/HZdDuO/xl3QFC2OmtDehP7yhPTD6tZZJD0c1r
k40iZZ1Wcwtjf0DoqMIzTenbvQrdIK2d1fVHnMJkt0eEtlVRir2B3Fj4S5Aw/XJLVjGDe4LatZ4/
DqA3pCK3CiJK0L++zadHSB3xpPiatQ5q1aXJQIfHf+GkmvGEEOjqTk301gVjCjfUT1k3qGgXtSfC
FcMPLNEibI4H4d7RT1ABQcBre+Q0OZNGnhok+dm202Y8nGyNir84qI1o8Qs0cEcSRzWXN5FO63Yi
PGvNd6YNwNTCaAP6KSevkP7mJW9yGaNkYyW2zJZWpgIWbHZ9pvani4esj+pSElKktsyUsLgzVot5
uLoGe16JrH3SyzOwIt0Sg5jNVoDxpNIhz2ucUDxDhwHba4u3bk58Os//Sxyd1aHL7qH+4kwl7R5i
buvnJh6HCcxsbqOYTjBYXorooKJiIOZGVI8ErodPD7m2cN1z1FeZtIAuG80uz7MALqIbAKJwwBcm
5IYcu5PlYk6uAANUy4Pajf1nrRzGvIPDM7HPdxMW19P0aDaVG7qnzNim1PCLGyz2dJ3QnUhN5X7N
A1tlmMTYAbMTuN2UrhPdxwGSi7Q1BpLcLpVNp6cJHWYRDJuNl+uEejXXJC0YqKcE/QNBurHlAJly
sjs/YqhSvw1kRAzOcFmXgshoDNjAhpNCbmiqfjlw9Xg5NT82CPaEnkd/5aU8mn2pRx5smqoNEI3G
C/BZXZtUA1nvcUJiBy1NPnJTKBZ7fx6L+o5gFRGDV0mIF8qkXhCmHwMrjPwdYswk26IK4kSd3Kq2
sn+WHx9mec3RgCJC23bw7CYJcjZQaeSa//BHLzbDqDv7NQC/FdG0HP5IJWs1/6hB+JfuV7YPA02+
q5NyNtgb4BRFmVlmJVxSWJf9OmkcElO1hzK1hnPYmZAEAwcVrhOXQzBxQI1BcPd2DB2RvZ15WRLb
Dvw2PBMFmG2fwV+X2Xn/Zyn4Dnc6oCLd5j2M3H6QW2xV3iHd9qybd7OPsltaDnkAqZJ8AdO4zU5n
XaZ9WtE0Qzu85EpsSZBp492cM96AegA0jB3RI4REyKc13Ddl/ESD9DETgfX5GAv4TxB1rOEA+QIe
nPzIfj7OcBBgINWRJRqUPwiWJGBvGJ2ZMwOZLocYDEdaB3A8Vn5GisyHxkZvpWCqDCwENeDDMhth
luF+uGMm7SQO1gBG8HYZuTHNPm8tPkKGs5r973mnKUrn+SPLzekwzSyy++pKBkYSz9b0gXpg4SvQ
dv/zAGjDMI0UUiWfMELRJkKAan1lQDhuulTLzvyhU0Xv7BemR/48AGqdGLZGMWeWMVN7xu5z6cQy
ib2dB/Bjc5ypX7dUy0bCLaCQhF0IYpsksr6MUsheRQcj74ywBn/ghpa8IzuAJxGQCfbCIcyqzpKD
1B0zfRS7o3J1T/d7+69oFdsQsh7LjWXhTbUfKYyjcWkmiEoypUOYLQmFbXNJUSQcCddbusyq38HA
jmy2Scj7lAHP+/Sp2Vx31sfeBbNKAHOY3pSizfxagTmPpvDt00u0dYdzLf/MrzbA5C1hE88WCFiq
BteBEMjb5FUJEHQKtVevshywb1XPkbkA10U/rInVkRYx0ndS8E5pXBFB/lxWnP78P8hGVnao/Y6G
PCnNO2+4hbgFtDWip3P6xV9lCkX5o8DHJE863uNJimSqDpD9u9pZvPrSulfr+rAiQwqECzXICOiT
U7AkFsYwly/pile7BUqJ1ny8Aa9lrvKw7qVj1LDrkrXJrvIb5UeClMojv6A9VpRjHEpZi/0AZLV8
0RIcj/G40duanE8Sh1CqOg4w/DIDZHXrK68qTCJ/E85mAob93+HylAvst4N07Mbqj0/NVKgvKlBC
gxGJQy8dlhHeQarCBRVBpDllSawuEgziapCB19r4rjWJ5SaXKs2jfgyGGqy327PFyu0jEw6VQMf+
QErZ28nOyWEWyZyZ1i3O8YwV7cklNviYa3/E5RDmlr3m8IsXkJMkZCpkiY+naAgw5GQR+Od2R8zm
6JHvUizAT5RLBDkI9vrzFoFPe/i9rG5IkP4/WNCfsFKjlHefT40pl9UdfTykY/eAOLbQKVxP68xr
h4psMdA2u/PP7nmneUWqvdkD5zjZh/HGHopA5BfEJHPssv3xEr7ml48cUliNF2tv0h4Oo+DTDKUn
E/sl/BM4qY2Ly7FaHO0sSAwpYDHwYQJUOL7+J19xnjxdgW+gkFYKef2gXuWI2hs06+nciAsPN8pg
vTMfW5POOJ+hcHbRJ6Hr5ZnpsTeQNaxTYiYc/xyJgLMtBAn4qSCT1WpUsdjGhbVcusZko4TuXekz
XgkPlbWtjnzLPKQtWiy45o+lBVMOVeBqar3TQEujgxoGaxlm5E49rmiv8HqVGGltGEe1lFi3ziJ/
L/iPXeO2UPnnvsuzTcC7XEmCh+gP9opDytFCAMeYR30HmCjENTNzM3YCNUa5jHxPDtW1zMlwnmeN
/dbf1MA7B0hSWWDln9FoEmto+R5okQ6TXSJHU9QfUlSolTM6IRKwkuFsWVn1fke/OkokfkqJnO8T
Ha/u1m7qqnqlf4uE7+whjKpcDCXE5PMNGXPvSsWl8CxZ21x1PUXMUpWOs360uPpsHNtreY9yxh6G
edjDR2d/NpsatzIl9ll0ULLLCE2V8Z8ZEBlSBnQEYpnpMCmx9cxCx+D9tNFUa9n3cG8EtwZpO9PD
TYVyz3RMEJrHIKT4f/tSW1OsyywZlEUTn4yg59gMWIoz92sr7D6lue9yvgex9aNiIfwQDULmpfFj
CRpe4iDzB5vP4K6OPM0cJl9tSWTnuH9uRnm5zf1m3TDVOH2TgcLQatUYlZO+aZ6rg+pPCzaufzy8
1SYIhVC7/l4l7Hm1CyiYSYetLidxTME+VWk0NizCJ7yfxoKO0JW3fSYML05G3o+CLbFzt87+vi43
JL9w4i6k9AuYK8P19riUv+L8/xC69i5I/l5BBJ1IuPETqeUyiwEa/TKKo2QiU35Kmq65SKA5pEu+
HPk+z94dkzZXEmNhlMKolaBPCPpku/4OmNisx+ZYGuPl3kvsTsYZhftKOtwWlSlUKwRwDWVd4PmT
y0jaljfaAmglzK8z08SIPLNAg8P/bU3OrL7XpxzIk3mXybeyU+/Fi2fkASN1i1kdpaaA+/F41ysn
UvHGGBkxnfhdYDF1CEFaEXi2rpDOPdc+Uyj/26a7y7u2CVeIVJckVNp5BMVUCGO4YCRnQ48PH8q+
nnAIByOou0qFTx6Mi6wh2QxyHxfjFHm/mfaqE4l7S3dzCnjAUkoNNcuP9AM+Xr3Fd7goVFRc6IVB
oNV1B7KeCSniH0wICAn5pjmpjsaw5ODX3QvS2VDSiRttOJqgkaVm+OlVE1Pdu3SVla41NBk+vAoI
omPePMYhki0cYcKS1EBQIt9rijHyBTdFAt2v03N2eLyahLZykm+sgy+Sy69Aj5xHmEZ1dk3jfsj8
TpmduMNyNEWGGriljgSOtzqGG1qOv1TTBPC8l5TimbpeSyq+TwVn6wsxNadIiwH0QE3/7ddhs/1N
PxV9ehaiBEbfpxp2HSbc6osF6QJ6j4lhp19CqG2kC+hU3sXyuBo7/rU4t+k92ml5+x/fsH/D5ea3
HuGXcuhpANchzoDDt2mw1zigCjtSCgCG3uha5V/BMH4fT6aheBuHOsQC2CCWDOiPVk62YGD8ZNZe
4iZLi+4x8VM3q9eGFfoB9bo/RQ5PSUXhXGcTMfcxMXytIiwX8q8T75WcCIyKOK6Sm+WSJf7XK7Oy
31j1a/sd7HUU0m2LaOL1eNVTxqJiIA/+UYE8NJJmH2pRG6tllRdbGp3rOVimMu04ojBjncF7M4yA
ScQsUVF11Io2sA5WrMk7YsSK6ET7mgbdZJeop6vt36aWjmUmUJimcmBv5qAmMjJ7d/5BeC/yk6VG
rx/KORJOX41fywWvVslCZ+/S3/k2FtlKzZ/2dXv4Mo4mr4Ar/YqI1zwRDA7ISLZpQeaiONru5ral
yy2uPnmU9lGwVBUbV7BCddRf0oXMoKWRsJiHJdRw3KTdcs1hXIhHHYFpldu2WJ+0FGZy/zfrNxdk
7JzguFmoETYupJVhWWg5pLIwmBNYsvdC9R+8B5FLDfJBgMmjaQ7x6tjt7w5rUEqOdMatjYkjPyjo
0Woi1BRc2H19NrGyQ9cOjYg+lxZEtVttSh6BFkGvDftWOT6gQBcM6GK9/RavLuJHMwWbnXWRFBUD
z0www/L8C8GFr2HgroEfO38mchfrE/7uA3kLRZpjOJb1ZzYf3F3wZv1fDUQ8I9w+wxhz8/qLc/+/
RATB5dpnmTrjguqd/3elSk91jXNlwAzXKENFS9jv9fvEYXG/3larCxqf5xX784O16XeWTtO6xctj
wf3CgMbVaJ/Pc5Y9OJfsdh/t+cF0PqPRa4qTn4+ILN3wvEtQUHixbVWoepBFgKGeOZyFdO6MAgcM
t1dhIDBLxss0xXFQTWWJKC8cdr8ITKzTBLi+lLu48DS0Kpj0OGo8A+6ZYnwmzodv7/yui7Ym65nh
QxQ8dlOMGtATBN5qomNLzmrnf6VsjbtSu7YFkY+4qrrli7oAC5luLWzJB40m8m6psoj6VNLqepx5
CNvGbOb2YVvP6HVKNvLaf+rowXeWDhzRNd07HJz8hPqYabDHZf8SykPrLoLuaPqBl9b1PZK48jy9
BsEdnjIHAP3mdc5bgRw2LcFsuqGZL9t+DxZ2cZZeCP5dMHyR9hxg8+1FV/yp6kd5CynbTrxksyWX
ufS816hTRtF8grxtTftYZY/veqkMh7EnZHrNknwj1/HPFSZOnkP3Od2fN+QP78XK6pLVZ7LDABuv
32ZMfu0aBL4l3nT4BcIaEt3FbcRvY1JJPGUNtExjPJGVkE7aPqb8fUEQu9JMwcRYood0nZaLpucH
4hRx7xH4SHcBvu76oGzteC7PC5Y0ZX4gyxJYkpiZ2g0zs3ns99qUVQUYrMa3IZ4cZULFXJpgTY7S
Mke6UkW83zrcliJsJM9S+XvYKoYxaxayqUiv0yO7d35+Rgq2r8/JCFpeZ0uRlP3APeKhxdnEENfI
ukBlMMek1etS0uBn6shAY9eOispVJswhePZFTDKx4GvcX/3PxoZb/pcMWJwRjxGb7sQHj0kPWVKo
D3lFnU0p5kI4o6DwzJTRuHLIHP12Kn8hmcwV7T86BnhxoNvknPFMKPHOVEB0gCP2VmoBPELUyHep
4ogU/JRTKj/zINqvpab1i+yH9mTtUk3LUmaBklfud5rQ4CbEAx1/+sca5+kjxH2770M2ChR5dBQO
wPN7VAhnjYcFLuZ7BTBPuwUiRUsxa47KQ2btjwUQMGIDTQSv415oBPZNbSePBuC3F3qRoleyUKZA
r2MBFTfxvTfjB83TIiob4qYSpYxHpTJKBF/B7OoMSUV0TluglCGKxMrROJVajJ+OJLrKPMy3N9Ft
nTIrO/QYJ4ggdPaK8RWhfseya9VAnBG2sG4w09bIg714RR1wd7PKXHeF4Wua59FHQasgD7Pjc4B9
//w4BoioirJ09BASmMV8DopwKnjCggkgbBiMLXLoy0Hzo2vZK7dI0rbFikiwoeW6++FbapjXYLeK
azN5qXj9O04yLgBUKIN0SfJZ6sXrLt61wCKqpklYBkcua8HQk+q496GRn0mXrfWVoQZul73ZwJ2P
ZboKS/g+zMGScC21ryeC6UBEk2SLVNU94UMGrBgF7r5cG16QkZ24aUuVOmNONYeGYgwv3cof7xqr
VVJNtBSsz8BmvxQLVJv+2Qp6QJqBGsDG1AtmtPPrbkNdpUWCjKEoXXDR9/kCmqCxwIyn9tw8hCUw
XqyJ7XFkl/O8Wzr8bfL/PKE+eIGiLtan+SXpR2Ok7hNPpzbtjOrBLsWVjweQ2sZSaHigqxQZKEuR
q/6VuWEkM8HN8rAoqvbKdI2Mf8GHevbvUHYISYhMQ3ZwMo1sm2uC9KRwjUNTtyHCNsyATDq2UNuY
nhYkLTaTkFeGvoF9EVqKSDXAGRw+O70NxTw2/+yqSlBtB+PFLugiw28+NC1Uux0D0uSu70A2aJrn
HJ/VYqAFpqrLx06BaOhfkcbCyzQJ6RnsmfS67i8ig53TWsJnfmihLAob1YM+OgyT5MnJ5JaoIP3b
MguVl8JpSWCXcNps8kPiMRV3da7tvKwElUCiTzDVHJ1HhYrEkO2rPPXAKeew8IoDeUdmfR7uIyCi
hh59dwlUu8/xB8Oox9VdABay/Z1dwWvsTyycUpxV9ATFooDMdyxLzDUBhRQeWItSPGfRF5sQFR3b
x7zo2QP6DAXk3yiDB6JR7HV5j4qETySYqCQYGsz7sdsh5Evq7T3Qzn18mvMjTttEcM62Eiu4oTKW
mtpKccyDzzH6L0P+Q28Wv92kQMm0kUF6PA0p5oB3mmTbE9Oy20/bUGHwssXIrqgyk/BbXC5GxqSQ
q2n1NDiAdiNIi5rSKVu6Ys5IJyvdKtdD+nNpKYK2EWeODwyLU+axbHRgajw8pLfUQd0O7r6VYc98
uXwnv4A76DCR3xEd3bvYRfFrKIcQBo7qEg+Ui8Wq0QgYBT5VRn6KlBmT7sH2uzWY4/f2lOi85PBU
sjNBkpWR1m9Ewc3n73Gv+NsN4Zxmnl6ImxWkUzfhuJ93lfSUtq+Xtij/1Fqi3+MylgqdtbXxtv1s
VddqaP5c8o0PVtLWwTqHEezoiZyv24kRkWnkQHc9lehxL4An7+CJg3kAnRc6Zo33qIWfCcWR+CZC
8gool5/SeOhr6yiOzpXQCuWbBUGCH68evA+iDsXjEE+XLTwB4+1wDkBsMdf3j0ir3FcL0MkQAyOQ
zIvxIqSC4nZErg4enYFOJYuitVcAc92Ko6PwC41mR/KLvRMsEMEUmp/Ak4OuRbKhyenFsvlL53yS
FmX0EU4Vn0y6PFNh8WcDSRU6tLm5dEZWQNhxotpqiSoiHQt+E3BhwAZKZH32jerZSFxz97SA+UD8
HyfaXD5lJrCejSLyR/ijLoTt8qf0eI/IcSwqS47DJZqVaLzk9i+ynl8+SQMa4klhEbvUKjxwiHKz
+JGin61CUA5Ut1opg/iS4Wg3wp/g0Hd6nbqTDM+z8pYaGlb3bXKZoW0y8axxV8mErr430lFBL897
4WYgx8Gu4RJfRDoc3Nkp8C6RU8DFsJq22GV+uKLA1QcjsiMRMdB4B7nX9YRtThb5qsVBxwo6fXOP
QIc49Vz5gGOOiwrHOTyDuKEDd72Pc+pFwI/FiD3BilWAKF9unAjg722V1gTFoiXic3gXzocdRRCk
79yCpMPCfjgr0/7lMr9CjPIJ9bUl9G10LNbbr5MxB+ZX+hjJgLOdOc/J5TyNRS0MtKWxxXW8F+2E
c8DHORv5SaiZdPZKgM8NofIbbu0pKLeIETo6z2N24WwOiBS3WKcV9ADYwHaVXpi4pn4iJaPYDAVY
COWGLLLZIOr6/eQWz5tGQexQn1QwRlESQHQV7FaayDUEEWcAy5+YieS+K8OcpOetbOW3o+P2hXpI
7Lm4ceRSYcVmVm2kXfE4S8FEuZ/c/5XKmmKAJdeSjkFIy3Uy9plrcyamOjGmRD4xCF+UgHbpIxQX
SfwShMnR0pypedlKziISxfEAP0Py3uWTRtWcD7SR/uo8JS2o2qeL8C1KO2uLjQByLybtfeQHcDdw
C+Xc3I6yBkscfkZZj1Et/V5IDYq9Adv9I0FixWYNVUlTL1f5lg7NUutLRYffgJwsYyQpoy6Z3A9c
vFjvUIgV5dok/AbY8knJXzMIeKv3H52xyGvJix/NmuTtKd0LxjcKLhSquguplVkQU+WgqhmjsutO
qY1dED4YYh7hiLV+5pydwWQS6IHHq3Cy1TgQ/3ezymPCcEefK5taW5cUPiVyZKO/7aj6jnHIlFs2
q4CCepuAeJpmFt62D5i/TDlgKkBph6mCXkbEgv4IkchIsYA7npMnTgvyOHS77LcisEI21A13xBCQ
d7lZDArgW0D1fb4Eef3+JhqztpW03YiRUhtJTI0C4t8Cv+aUdb97UACBBjGF7Hb7vkP+4puGrqxZ
w3w0j5Ww1R741eVUJeZ1XOmhCYCuXtnKqSDRfrjDcSQEdWLrALpeodB4zLwZ6fdr96odSqUVcjc7
aQt0mnAEn9Byfkn2zaGuSLpbvScBeIFYE0/9O+Q3FY8XsGOC/Ees7O6PXd61u+2+6mjteh/4wFub
UhfJ7a2pEeZ1Ssvjx3rvJkPW6dVo8GUEAUZlYg4APVmZqjEfVMghKNboGAMzbL9ns2mwalFQUN4k
uwc3xoMcvZdoWgvY5a1q5kSkoAmBGxTUk1YitKwp65nII8PEyBjwzTomBs1H5fEfIY+zxPdauZUa
cHYL3ujCAmqsPjnsjCaZ/Lox50SxlS4iQzz3CNXAhRGLMVP7+ETlDdUit7hqZCDlwKHb1TvzVLIu
gyHL8Bl7/t5YUgWZcC63OrkGltSVloxmWaaKbkJIogJyfB67J/Icoxcnwv+FK4F6nXUn+CZIbLW4
iZ7BkSHOy6AXtJ4Tf69qC78+vMFGWESCzNUc5RWno4hjyjGwHNjmcqHzvs8IFXTWGH+dAus2BXl8
ej2FIbpxOkQjR4k/Y6I3Wb53jVxzTMXla/bRF9ofQTzQpPkOydvZDadlzvBvjP9c1osV/ntoPZHa
J9NpnuPAW1m7r/O1yukSLGeVTsUL1CbgKKPYGEYgvPWXKBlumObQkPRqz52jKO2MlEzQrIfe0jbo
4o4Wp81zjmYswJ3BtuHQB/5/h+0HiiuVkuneCQPoeBSxGqJT9ZMa8R4D4BCJtWBoTqbm8lZEW+3w
qq0nKcSlCz5uBIZEeBstdL4BIi+En5mbBqT9hlihYFkxV2JAf00ihnH07LAHOzkeBz14IdIkJ+i2
ijI3M9ufbODAxHEb2IouMSqot6BgHnBEcSHW4JQ0LnQmgB3Ew/pNCTLwHYbrTqU+ncETMm59P1zx
5i3eG2WH5IR7rcT3YU3f3eSMRM+jqfTVTebbbFFno3uPWwa7pzGAVEridKVsBhHkUB36VB/vJfv/
2PgRTYptSh+5xpfJQNiLrQyArQPMmgWiJMvHAwZ8Ov8dEvWndXk9Oq8kUJJ85XCnRTLBDfCDFENQ
FGpwJQ9Oj8gtOFQiv2RDOg3T1wALDO4T+psOqWT0jNhXfPqVlZwpt4b3fFyfMqTSLrfAjmgxOk8L
K49FrFSfpJRp/LKgVhQc7NgajBQfHUYchB8qoY99mVU7lZCQGbR0cImi8o17eyPIIcm7qYH2jdUJ
UM1IPCWhA8oG5ehXxbLB6mUx9fVz8CxqggQA14w0qeFbckeQfbadC+65NTWV3aqAEUaf6l7KAEtx
PwFtg7EJ+SMAMztqYcnbWp9QJXtFfOU8GmUw7n6spMKYUuP7vMO54qRLsPUXBqtwLIvozruJM05T
hPU4ROCpbJxs50NurAvTRDBm7UAQGjHSLP/BcoFWEcERddYED/FM3JpG1CWAcnKXOu7W1acHnPfI
An2XS3moXaGnyVDX89BycdG9EL1VI2uUfRutUjQYdIk2PqTj6I7on3AlKktWlV/KdXbehL5AheDh
obxpVewmWfd3zoAQtus0cAnWKYYmRRyy6AQiAit+TpYVaRNOhgkTE9W1BHaJDcLd43UNmEZ7vWCg
NsD8JsVgzGRRHYxrW4+ec74odrB6a2YNvLZvUmVYod8J/sume7i8W6UBkHUITOqG3WAsvPckhJcp
OYB2wYu7OdPsrxE+U7f9WOvoh8dN5gEe/78OkO6Vkjk4eHTyyackx7BZ5qDoQ/9Ex+PN0Vvh7ws2
jFN8XBm5Wytg1StS7HdhKF2uzv9uflba3dSwMgZqcaU8REiHocMecKOhqA9bzSOUy5rp/6A2qQV1
BdOMlBFv+5GKdLEzsREUkNkhX0LKBi4YZdcJqddvFRYYr9mS3bEdot3TQUHsb+JBw0PB9kKNPAKw
lQUWO1bxT8Kglfdp4iqw3m4i/Pfw5w/slAhokGv3FB9rPfy6LfUSIe5/lm8LzxNnClz5jAR5q849
ZYXW8TIFwztz/7wZ9+GygwBrjxTMvqlX0Xz1Q/6GM3V6NDd73/bnIw/boklRd81wKIuoWwTbyGzt
d10xJG2EA8awFgEu4v4AdkEu9hH21gG9XhVmgkxWIn96/s2sQ/JuAJS63ipFFfE0j8cZcnA4nVQT
wI54+7+V2T7xG6WPP9ZzGTn/GCGqFJXCOWhl8cDFDpfFePtNN1bTzvlT+TT9UN8N7d2bOtr6WOTw
W/Weykq6vCtTABrDLEUJLF5uExCQB78HZrLFmVQcRSb9LO4+uc27Ip9LmCxGMbkSlJnQfjMwXlrU
8vVHA47IpWdi2ADb18j1WFonw+bNkYyy74BEdXQpInJ3Z3SYyRz+fN5TYFVZ0+AT+9vpRNy52duM
OzMqPc32/iD8rVWWLkSRFbmZoawAUm0CZYIvqTrj0uW+MJGHyg22hrgMyAvg61/7XOZasHnQiWpT
/j1gMyIuoQCyqF6CCYQ87idOIyWTsOviVmCNX0nG0ylO8gcmJa+SgIx4YWzoSpIakkxAHs9K66gv
XFJZZkJZP71Nz9SaGhK0EuLZnKpKv0wSpG3ELUyrZ4RGVqy4OGJUwsq75Qz1aqy1Sjqkh0x1b+h7
tUv/PcoJK3jJxu718EE2eJSkpTbeJiK9uTMby1G6jx/uXobu369aiEpLOI81+MYoTUWJur7mENXo
ST8HsgiXWsX0Wl7VjztbmeNUYOqsHIJ02sXVq7GVvdbZ7RH5LyxtlBkD4ounXNlo7SHaE4cAaPGQ
6h25WI67SfVTE/Ovg3P94B2B2JeEoS8xCdRj7pv8ljSyHj2+uUb8Sgp07Wp7iOmimzfskPPDMlA+
fnkC7aojnSVTctBgHjLPle8PhrB/IuD/qDXiWh9bGUuPfQF3TON7ZiNOCA3+Bp+GB/XosfK011tp
UM+fy288wAG4R/eUFJ69bhwD7GSq9Xc0oBNnw158VqoB8LtQe+e/BhNouS/i6xDgKG6DONSCMNkq
z25fy9sid/giTW9bRRpF6eUGXfJuSWhvrmVvX/DcOirca6BeFdnLhEaA77cxucqJewLfl8V1L6d2
GO4qH/MAEgW98NVQhOTF6JnfnApxbj8th9DCTfTpq8+KTlp7GsWwn/opry/lBjJqEv0wYDXlZT+w
ykZhOYcmCTY4yzd6wB/I9nfYnjHiUDkiL2Wa1D54i4qY/aA5lvmRGhbWTVga1W3iq8tDO6CkXCkk
uHEayX1K65t2wUnbAzvJDaAQsWWjPsULGmpQsUW26ip7Q1Ko8UptZUw6TjCXZXf3YvHOng6RsE1w
BQmvz9PsQLLdK+YWZGIqrZMjk3w09RVPAAAJLsApXwirWnLLNzSjYgwIrD0hCuifZ+ScPR1Wd8dm
cYxFKmuYhqN/wArTtLHl1IlPFhP0I7qPeBUQDkcI7LjeCEZiXhXNN8l3IVNak3oioOG/PCBsAtfY
sisXgopxv+nx8xSnBy7LjWn+Dtb/wA7w7i4Mu+iuA5psB0S273oAESY2O6PwknjeND7DptXB0gzI
7zTMq7h/8FSfNZl69G9+CFveWbPBPzAv/GZskW9ZPuZaN8vN97qTIn9VgC+0nb8fF3luaz32JKI3
nCLmG8gTFz1btNlS/nG+/9XBkGR4O5KVCjgJKQ0lAuh0qNUXSEVRiifDQdkMSx2S1ajkFb+LsuWq
30KFBuD9sJyECztmUBFWoU4giCVEVqIRmWks1eoN7hu4vv7/CxiBPNrrCQAM3O6B5X7DTR3za9uL
pCcR2dPZpIndFuh5bpotb5IV58t56Uw05XPiiRfkrRK3tKjVLCW+bh3d1jWi7gVJcTC6hViNM2f4
ZYRWWswt7t2bZUb5eNGTI1bdFRJaz3WabZ+OBIYQNcGqWgM8PAYC+W2pX/CqLbpbzK87qgsTYf8G
Y6vK15Z8LxVIIKXawjYXKGA+TpXom5frPdl9pvxrDPO/rp6loRxsuYHCVtsDRNBQgHuenwtHcrXd
YBdoTbxNRloodXEPYYKbYLpyAEOyivC+lkI8fi7hHxAvx1ghHnPfrZPPOSN7ETFT0tkqL9KMeH8a
FwcKHV7VTBr3caW8ox7TbZETMExD+qbGV6oJrm8N1A/8X8P/3tooa5dBG3gwzhkUZRH5ajlYc4xl
B1fc8obROXg+eKwjczejN2Oa6Rn4lVV5i3EorqKy+xkzti0rp1hvVlv2Y93rYzuKEiXhIr0152UC
XXbT2cVR/t1vnw4zX0MHksshTv6PGt7fAF187kNsW7IBtN47jdv2M6INXEq8+xNmlwyTCQmDsA3S
gsLL4aqpmRhgdRHDsex5LUtfjTjg9CgXw83ZBuN5wR00shRBU1Q3sqlxw0TdUki32AE1vv8wmQim
mXuOhsi0RiBUYFzLo4Aic7X0BiVWFU1TFkyn1sJyj23oZ8dIuxKLSsX1Zi54u0nIho3vHV1aZ1Nw
+0gAqqtUcvXWSacgX2N2Aywc84DbrArZYHkzQYa9HyJCzG2GN7nMgPDqQvXxF/vom3/hNuXKRBp2
0XxVQDugch2uNAMeMhH/auM/ulB6n6tPwUHPJ6YHo13gYek/STg/arFNh2EowbQN5UaU57aqlvA+
QuNB21yS0M/PDHPpYBnK4Y6nBdYXSmzCwNUwRH7/6Y8nghJ9gwJ5fS8b3YNy0tt186nGQgMUNjOG
Ngmy18Qol95vpRA5T2pBI2iqa9zzQATjsFXgaQHRG7MNLcvZoHUgVFgSTQPRYa1UXY45WBZuJIp1
LGET9l+11s/C5SrdS2l4O9ypO/nGF+LCN0c1kxPLSl9Y89WW5MqKSGeZ8zlaUQ4VZ72+MFIPbuFF
rnX0AIfEU7+2Uwc949YfxMOm+dsMcGwVX7GZ39KCV+vRCMGBQQSwNad/i3pLjBRDWikRmbsEuZep
kByXtWdmVfnGs/AXA2vjJm8qb+n0tHVZP+PkAW03pbIC9iGRUa+dFEAd04oGQCghHcEtqqmD9QOj
VDZxnb1tyjzZQvbGZIMw0Lj6ItzV4MmTDJC2NHXJlrJ6C2jdTMVYxjLGhSRQX6nL+CaciCu8I16E
BZdOq1xAgABfibEmy4Q7C68k41yTFfViXQcSKTGAJCcBKqe9asbDwnonjuChCURHapY7jykpy8z2
+5WdegZcb9tRSz9QyT4tnfY7Nwkx/kRP8dq8sQF4NKnO/j8wP/myLum6aaysCj4YI7Hdq1JyHMGY
yeIWBjzEZLEevWkf1R0hr0NRJkbnsR3pKIM/TN4z0oz4SSKrqd/i2f6bdLF69SuU1wpbtKHGSv27
S8NYpIbvi7sxXKquNRJvhjmlUFxJIrJI/YIfpCteuaVymTelkWe/txeMucvlsY5nDKQ1TX9oZqKz
SPBs4tTcfUmEcMjraQ7I3rvm98Hxvoju4T/r0GK0dm0rukti8NJjxEo/fPEHFgmdb4Fwa33qIkZB
rjSa9vrrDaelWFTbxO8yiSZzCQZg5Eo76zg+yLbA8QY5utCjPgIwMBKUyGSxu5i3LVtm0J+k6R6g
Lek93yqzqameXFQjsq8DRo8wEcejLhZoaR59VovEnPE/x8jep59FKpa9VDoak2nggIeAEkolTZ4h
nDKYrcd7Qsug6+PfvVDN0hq/WJlWMjTQIonfwaKSsz/sY5Wu65Yf308hpReVt/Hwxrvg9JxE/WKE
3dX8KU7fcBa0S5k/WIz+ffIKgL9n72c8XKOVTLo2d3Q+ot6S8+ih+sdkXT/pkxBYVfWIvzvorda5
O95OHHxdCvmRuksdf/hxFLOHd8cBiD0cJm1YymocCMTeDejZFbZxeQGWf8eplUMrfnLTGmsgjyzH
Lt89Lm892Bt3x9fIZ+J36tQxTVXVXOI54ueh9Ah17WXBGYwsdXluBdeTlOX2ICEtPOeMNQGM7ETp
n9O/gvi6NxkIRURkh1UCQZbd2pAeYadlHGVqL+vwzyvN85RRii3d7k4sGgEEcTxuqwaXm13+t7UP
S6eKxceE5/1YAZ2A3wQFxOv7Jwyp4M2LkJf5zCBEVmL2V/Qu2plMF+rnbP5pdxEbJjiNTCYvq+XZ
lLf2l7p3oQGVV5kMkRUXAiA2mwsYYAC+0yZN52s+cn8TNVfCXw5K8HjZsovSWrSf0hnUTUqnC7Qa
67gZeNQyU9wtCrL94jg6jv9hDv0Z7w3U0Rt5yDkValrLhWNgDqwnlCn7QEcBdBZXJK5PffOsAzaa
eIrovZRrgJNQNCQeKk7aXva1/gtOgWDQXXOK56vFMB6gAcr+NOOcfni6z3bfviIKzFcn8wKg7Io+
ERk+2FAfsiZVF2jCh8V/dnKtuJJg2vEDwVO5Jbz02Jse34rjTamHzMFvKF6gJCmII26TGl372TKf
q0eMdfa6gbrqo6ZjqfQCxWjXZjTDRTHcJazFvpb+tPJec7F6fGP/PwSK38eeQM7J4vPz6HvS5ICW
9kMrklYzqh8e+R05n+vD0aG/rmSByQVVd0keaOe9z+OzpCSO+GBwvbsbUx0d1s+cbIxmVlCeuwZq
/FnUNTq5D9YuKTFJckSC+xwTFbyrf1vlivqX8MKlKlRjP5M4ckXWHJbclM3Bt0Xnscwe72mRXTXx
z9nG9jBIXAjaoSpo3Tf3b6lvTN8n3zY8Wlj6m9X9WcNAWjy0y9J+t9TZ79m+2GTqN5lzMm9N7TvR
LKwlEr4VUiXgteJWMGBUGhGcqki47dqB2kuBbtoTeg5FdoV8XIcBXgj5NCY8YeQwNQdHgQCdYGem
JNPjjEi6NDBkB5bC/S0oc3C7jjQ3jM2unL2rvP6HD7NOEsDe9yBe1XjDBfPZZFno3HPsfcaqptcA
z/mt9bFvLQ0V94ihDzMV1Zc/9DJH0IFxC81YO6p5CXKe81m4W8EYQV+P3oibJxUCwff66dO7Tb8g
XYwBHCPk74aSzsUsnuicjUi7H16twY9GjmXQX2yetpyNATs04DGNXRKOh0jiGQMO3KkX3cHvE/Bp
7yKdH6ey4K86KYu4EXCpt/B4dLWEOJSiWaJYighyLxKLzf+jjPu4im7DaQdRglmIZetozKEJS26q
/IXEl0xmSd1C4wYK7QF7v6Ztj0cFZ8ro4zRxTZNKcFhT+N++n3WDBp5BTRvtbV4auzG9goikid7R
kMTLvf9z18nTZCrv870G2yH9YX68dxVUl7yr7vbafBNjg0u5gjV8Qe8x+wgKfnh12mCxO/jJ+MPg
R3HwmDMZMbaipI+ZcZP012HMrT9qd+deptSWhwikMlfclv6aMtRvgd8ZRdecn1U1litsGLIOCTnu
3rk4lau3Lz1XiWxG4Vpkh6Mn/B+Y54Vg8gVvcTaLgEZ4++A1UZZF/1lZI+0WG16iN4gdHpnrls0i
arIF42lXC3VB/0E5wfKLoP8tlA54vb7I9/FA66c8oeU4GCSoYYStwwjaaD8Z34JfOq8xKFvjhO2S
OloqPy+8eEg5OvHTW9fSwLcSdmwhnV4amORy0amWm/IxpC0deqUCn8sAaBd15iu7v9ffrOxp36yv
VvBNL11o3gV+oGO8nZo4Xf3DlckDYawHjAG0c9+Qz65wv78tnQ/Q5TksbHMrXgjo8yNAhVLd8oq5
4JWcBWckZe4xJQNKJ5XEqYqBPp/oHp+TbDHOloGi8yYKQj7suO9W6izwSHEc43SX5/U5oCq8ya4n
Nxq6U4RMFAb8XbCAta6u/6sQLAdnwsRG9skVhKhiAtKLa/Dag8naTJ0lPxfreY8zYZei/ux1MM5C
sUggZIT+E1O0q33/erv00L1DGzdJfm34TY5jdMIjvcCaWrkMebmWxcHkxek9r4X7rEVVLAV+zvUj
XlYGNqfZ1Zoo00GUAMSa6XYHDoTufzHb+hQZGWTGB5HqTP+/d/p3RQXqusu83Ee5AxyL5BArfTn7
fygShfjX9Efn1n+S3+KNxfxAFi4LXlK9be3+i5HoK0a90VGSjSKX1Yyt5o3P5a/wYUXPJA2+9YVs
suJRmmMhYXGIa9SMAVLmSTiI05mblIgpForOsQufSEU+2HCVVaTpC85VEhN9k4aPlevumAfKKC5g
5JMMSySVMlbAiosSJ7mfvM7/6TcAi6d5cbEeQfj4bT2GHahst2sQqbnaNjwHvHXvb+IYb0DIsN93
6u+7D7nm38zXiuB5947Ydya5cX58cyhDjfyfM15HPxMZaF1uUarEM2gfxrJVtmTKUmeEM5cr6M+p
bhhbACxP0x4OvKEihHkrJ2O3kHNoUoh43RN+4BmwyxrQGym+ez9aUYubpooNnlcf7srsg+1yFJQo
yuybZgv76roviaUg0/Vum7qX/mtLjUmMKw9hZE8ytThKjQ+Q/fLMMG9U49X5MDdt+k3ZsXJ4hH5m
QPuIDLX4wL8tX40Tz21JgfC7z2VDvdt8uKvcxl2efRIJxphcHHYa2FQIzS33G2/01jZnTltHj+xi
XE9TVM8m2OSU7FXLB7Xmtx0ogrgA4Z2389xYEob8fI9F+Gx3HahC979rNDw3Tw7T0difd0MelzZy
gIADtfT6S29sl0/4K7bWKKf+w6bB5cqAYnixAus+SPG27+M2lPyspfIXMZDcVCrfPDJCvocNKX7f
CEM0axZ/7vqBJcykc6QI7EtW3SGkyoBZbAH8inQgBeJbZCqfD+duK9V4V9DPOVanpsJuRBt8aqbL
8sLcCitFu3iw7DHAaQ2KRt5zY0ckUQ7GYOYB5L8zi2IrIWbLjxT0XTeUavgMXVSnigL+jNGf8oHx
ToZSqR7CRgzE6GHzzUwf9nUFlLiT5FN3juahrQxCqzfv2RxyIluPRNUnwpqMnhWlMntddSj5vxtS
/6zhLNBKcMhzNS738rwKqliLJAQRq14I4uxGDhMAQuxLCF+a4YoTYXYKufvlnRzGkpf1LoXLtPVd
H/H5Du8R4XkGk9sBVJlxtIk2FqmApJLd5p0oGk0z4zeHG7qdbfXPC+e46aqfb0fUJEE5k/llFtc6
GAJR5hzYjD3UPz1e5Qutb6DK7oZAaDEwSEYVWZ/3z82p7KixR/2wkC2NlT7YVl8EUOnHTp3m/0gc
PCunpH2fcvtILp/PvavfSxoFE+zJsLcV4Ga1qhbkRJ6Nh4N1vMGdzt2rAA/0oGlGuYTaJ87TC8/V
Lnc9wJyP4dg2VZLQOypDn8MDlNM0r2Jbb5Uza6x41T2gwc0r5DUk9QnlROlNeHSMenCWeZGZZXu4
L20oI1FNlQbYTFjQzw9T+f2NK7QbO5wnTZtd3Rf0+EmVaULlgQbMfK/4Jcpw785m/IbBO8VIjzJQ
vXUYP9wcbXzS0Ndg4t5tCWXE2tkoUsqiJ6kdAD1vuO4WwkSLh9luE+swBEaqG0h2qB4yPgRNP29o
iHnjwGnqzlHHEqCDkEaNZBU9Db4oquBELFmbEgmJveahF1FV7rGtCHohiEdjOda7YCGjwd8fGGtB
eoiiTbcknShsnVSdlmpDVR2TUPijvvHh6fRemWQLyZ2lGQ23y9ZXphgyg336UHW5R5peVgZwF5kO
dmmLV38FhGcc/AI+FFbJ/tlstd7ADQQp4FtnZ0SNJ80SoI6dka3jvlKYxq1INqQ9yqYyZKs2Klz4
toj6HL6vRqYU9f2XZoO4Fw6+uw4rqyO6III2uanL+32W7kifpIAI3gKufWSw/uIDWMeUo6/z2qaT
VE9ovEmJnksq34w0LLQypTVTX0CNuJ3n6AwDkKiWPp5Uq7qOdrnWpCviRWN7rFCKnD2jWtFpBNVA
+Ni/hVLj6cO5WVKuLetyvu7auAjhEoYPQD1H62yl5sy33fo5XQgAVVUhXfruc0nSAvmDOZTTRQ8J
T52KE7ZjbBOs1tNuZOxaQyuGqtb0K3h8tRinMdxG5MF+TRJbSDZH33t3HA+zbJm10QDbeuHv2DDg
arg4y7zIV33u/lwwoSaKzc/m+pn9xUYk5h/47G7KzAGZD55rR2MxtTXGYdUiDhZFGOEQympPVAxU
kWQeAYrkkm2yZLYos3ooLFd3g6Q85+FrDKQLx9gZqOqL+PWz22+fjR2jumS/8EnHQ/yd7t9x9VPp
3+zO/rCmlMJEhjBo+yqL4nZD2D32HYMrwMeAP+PnYbVcakY9pGQoIxUZjw5aXjZ2DujN54LeFfE4
N5+7ZRKgIOiuarKnrZel+MinT9pXkyIuTOltM2JLvOyyxzPgE8kEEaPzgOnImL0XHc2ERRR0oVye
t/jHU9gchCOQ0But4494ZDLrthzIrcujw0JZ3mn17kMZk5hbxo8K5O87iYxjHwQSXxHkKvTI6B0+
smGQyMqHYVtvSRn1kQ5Sg7ccRwMWL4IfYzhbtZev3fehl8RiO79ypbobvv+8fsbCDRPvE/Z6j90Y
mK4o0BCml5ueG+odE0WvunuKJCDqHWKCxnb8N08agKo6tGrbFTA8k2zs4ES2upztfoeI53DSVNaI
DQECSLSU7vGGOpJTZQp9JsdpwEwWvGiaL40ZHi/qzKzpz0CQf+0Yo0kf6/7PgcS2cOoWM8dtdCmR
wDqY77uv5tbYzVD/KB5lmoALjqIlH6ngYQ4V3mBAdebb0oyBG8qTccum4FEsJjmCENXIMVXxiK3C
IzlJ0AIMQQ7mjXofre938BNx53+zak1YEZWSsY8FdloSHmVfo2ghESbgVOFeMKKWQmUGy8eFow4a
Sid93254u5kqh0itqGL3/fKxY2YVOnGtR/6123zJAvs3hJ4Fyr58yR2sKcJpiQ0VmNvihjXsFaNf
gJXFy0qRDTaYbWH7iC3G8Bty0Sebwryi2upjTBOT657PXNsQcucmnHD2jd+EbABMqNMoZaJh9eXk
VwlcvVb78Vdtn7HdVp5njCSSq2Oel88vG2O7QAv1bg5uTUVm15DSCAIbd5n/S23nl51p03Dvv48R
zMjyfzWIdiv3eNhlRRjP4VMx+qX6MUDLl52tw+CiBo4EBzTEgqjaHArHWymZJAehuV9xMrSPjtHS
dBaD1v/AVajW5WkUQ3RZ2WkuqwpSALhRiJThZ3vV9fse/cCW3ymnQ/u/mrEFis3YNPId+vCT1Ini
Gon93ROJPRzVqIBAhE3ezsgI9P1vv5AQb2I9CTAv7uMf03f8Htcw6AYkaSTNX1GxiVt3QQIhkzkl
nP2uQeh8XkuDoi/r3qUQbMHgdsBQ9p+2cQea9VMYzmbAu1zJwqS65VRQFrQWUo0DtImY8csJzS4V
mto08ctp3aOm0o5zmP/BlX5l5wf3XnkLI00Kyvhn9VQ3TjCeT2N+tvpIzMjYN5GGFqfAGCnAO5o3
Cw2PYxQW3OuvDmYU5bWVyfmHONX4zwhi4yFlMYKqhZd3zBOhWSqOdaQqmZjdyunhj0OOSrKcACSN
ZpDY5llPfYHs2owgyLqAuwRDO1UyNGs+DTCslnodRnSiK9tHQbLOqDA2YewUCEpum8uDnqLQcqoj
dnLBSZfq4g/z7v5ZKEpKu8I4JlXhjU69d9Eq2qTy/y12qsceq6RFD1a+MJOXnaAD0mrRcZyj/pqQ
l4rShRZQit9gktzCvCrZ+N3Pb3WQ8OYrkUYh9zTf5ZhrWdfSQFDE4cr1g2+QfHrLzwKn+5WtUMY4
gAAJEFYwC7cwtYT1Zk+boL2zZbS6/uTAEMvToxbCxrj+Mbf2F8hIroGZkDIX+W8fhi1LVCqtto9/
zUteFVjG+MkdenIxjlZKaKmZURLE2HK2oGLHII5myavqw0+/ifHh/ovWxDq7M/+uDy9S/J8/wTWC
ZuV9nWOCIzAJKq7Xo2lCnIafBqUEuwn9CpAja5p4TGiP2zgxMSSnZPmxYPc1gHMh0drAmm5862vC
CnZXhqgwWePFnOj0kENjRDn+APlWH9rx5Boe/MIblnoFpsryBIy8+kFhzhLMfkXP5nwUVPvYwKND
qBIckGLCWiXqR+HvxSL+oaq13YcqwdqIu4kkusaYi96ZaaJchNIOJcsV9w/dQ7bldKzz7yf5rpAU
kydipk11CkgzgJg9fxNZdfhLCu6Xkr4AiFrtmSPgtoErNikJcLn8b7Clhaa/yfwZDPP4HzhELhYm
fb9fekvFmE6AjTz13K6lfTw5EyQ3VEWkQb+If76QtX7OJ83SXH7LzWb7OrgyBJ1/cHppZkj5L0TC
wsBhl5Jn9wzbfTPeyEgyw+C2WDVtmRPv/T8uiaedHg39WaVpN/W0j1fqOTpXhWGgZ/uTxgZU+8Yv
iBUufIwoOONup1pNV2HJ1E3Aahq+h82ustsClP7oah27Qn59SZnZUaFzgS8/hkSJfB7J8o6n2ge1
e5BTR9aPw8g+YGHHGg0h0hppB5GK2cNTrMzlWyZryGWSI8HxBDqRGmXb1l+qPiT8OvGiQgyz3IzA
xnaJkBuOdvVpreaV5iXdtkkm5998ruPWClh6cP6d17RRZIo9WEGVE5W0Gj++L+9PRWfujoeF0lI6
7YhDIzXl5x75VAsv6/NG1ZdWs9rdcf9MRCp8SGdhB6UyRnxBGYKM8VuLjDACls0ATRwy2/EGGXSn
7ufxCSrzbfY2LiKXRZyZBnom2lS4q50KqYVadE7b0g9M2ElriKlDxfEBHsbLXNlG13EPzJ7qabJd
L0LNLLlpOscR+btMHPWLH/Ekk27AdiuwlkE2ECQAbU6WnM/++W469zje4LITpldDaAzPR6hM9UJq
PGUHdH+aV4PNI4LdKWeii+b0l5r7waeK9a5yMtPziKMpkjHzhkx4Go0pru7w5jw563u0qDEkPfOv
lDYwViy1MK3Gb8bdRLlOzkhYaVtvZdjKCqxi/el8V6HC62m6iij/fKU4uZfqtsSKpAEw+PrL1WOp
3VXJkc2BT4Kg2lanXUItjfssqKdEOk23OkqNDsaMDtxD5FSqtzYt6iorZRvLyvtqsmZPnpVWRrOm
utS0m5ZeJ1EbBWzWvfjO+nheT98JNBPnWl3z8FiOWKxgGfawMpusZJFu1Ed7eDO8DKkcumouR2z7
lL+KFcV9kHj/3gngsH+6IkT7oD7Zrk3ZA0/LXoEaVEgWLqFy+5m7VRUZXDytZgSqdR+MnEl0PUZJ
iKpLZ3WBtW/fjZgIxUAF31lxpMhl6iCPcLqJ0rcle4NoSQPajEYavdI38sLd5Ofz4lHwuTAUb3Wu
MuXIy6lCUCX8RP/R+r75vpicB8WrLZgDsg2HPwt2VrriWJlHa7QHIu6ae91A/9n51jCFDWKasO5V
YE+GN3xdRSl1/3kNMKfFeWHy+dpsISwQwg9nZu7+I5HfAH9R2kzcu5RWJ1OMH7Kce65wKQkkiHf1
6RHrMubE9TGzigzNMhFrWwF9bzAxhnutdjG8FxeR4S8rneATp8A14sJ/Z9csPbyBWGfgjN0dkDYm
CGaoyS0+s+r+D+X9f+4iVDhAKLRQYCPVn81iHeOWrVUK/bgKW2f+gE5tIKGnlOM11O5tXR7nYCyz
6+BoPQBpPPqxkhOHr5ACW7hahETVUFnGHgQMx0XZpZ5uE1fVchyZ31Hq6VncKgyUo4RpguUhIPrE
gHULI39lXQbtqijdsVp7fx7Ne616k4lx/FJNmbLUv8Ai5DGIRT0ZBknfh36lZpHxBIOVGv0yxxES
BFB8miPnqNWxgEqGJSFGMKz5rhZ3HLatD4150q4svcLhhbkVSItwFT5hCD4qa4yDCDySnm2+U5BV
HrM7HMk/0LBYV6Xq9WsFAvwfcK9JIrChcnsGnoappx9vYVBAEDPB+gTmLSHW+8HTBsV9ICsuogUM
LH41itNqFY0ykTnG95q24mTSVAh+3bUXNffcGHnpv3Mk6HhgvSFf/3ZUqdqMH6Fovi0q66121R/U
lRTg93yp7wFe5F5z/EG+JzUjowXTz1Jf/y2KBBrWe3YAzsmEY4x/tKa7Z+KqhxWBFM9jDr5sEZXv
ye8sDqFgq3kV0rawdDGceCQWM5llT2lcPqnuDGKfXAXYWLopPW/2guTXWp1Ak/kkSlWaiXFuhIAv
kIkNoB923xTitdAD4Z4azEEQE7OQ+8mYGJB9o1xxmCkZ9SKVd+jhbZ/fzCrS64Dkw0bwvc7/Yuyl
3THvZARYRd2K2u0i7Ku/btA880phBcQRzeXi341uX698xMrxTckBKpCxq93OKbTcISQar28y6RiP
OtritIBdt3W4zrhyfFJYTbNUbDLXB2AQCzXNZj4ML4+XKUhbdsoS3r5EX9/7s0MMwZ61Har+Ys57
Q5jUGImlJ2c2DjFGp0M4GCJxcuNAqfj56dJYIGewPZHpkgs+n2f1EO0mR+rMNeMmH9j1rRv6Zlva
z0q4MdBscm0ZOzHcOSTVmFvpEnaUCFwXT1f0t5KQK0QiNyE5N5xXn3IoxQ3lRvoumin5ePKaqsZz
wc+kxg5JXGcDnwiI8Lg3NFNIteHHOtv/71O3koFqB2ytqMcbcb/j+FF1OsV2rn5cp7IaPX//yg1s
qUs7CZ1KGAp2qQAC/LwW5p88dHmEHi0mrjK3mwm7okHYknE44DCLjMfun5kLxQbzx7nO4jX8LIou
YYjB1oZ/q5DR+RMCPM268gwic8HM0NKnsNHXYh0Aw2I48jZgilMBSMMsTjW30sdusIsRHVtqeoJa
4zAxXxljt8e25A8zV3lT8pNQ1Vo4akNa29wftF5Leic1Ymi1VqEUavFT8yuKkldY+urs52IXhfRm
J3yHoNjLMKAQXcPUlM5IaW7XKko56kVzp8UHQ+b21DCbFCh1gMWQcJKdA8EyovrlKs9ap7KW7mrN
UtdTWJ+1Y4kNPjb5NlwMtMx7LV4/jL2Fla2FKX0k3tywerPYGB7Gh57TQqJE3s2WdUrOxVseTyfA
ZSefksyMgqfcnxYgMsVkQMoK4wUdyw7ckYfa6ZPfZXbg60SsoHfzBJmMu2ZCHUHguSuaB3I9CNOM
vEiy637bMuAQWKg6v506wIHSxlZc3H+6c/COdSCC3PgMnmBPF1yYPbHtzdfSfHkJQG3WN9dovKQq
E2kVX9uu9ChXm2Xo29+fk8oisxyUBTtDGcAgkoSkCL0OZgguyekz/SA6a++mH+f18iSk1+AUVQHH
vuMcD3JF7zEw6TEZzZg5RITzsQqQnJrk8Bl/nXRXYw8hM/PgfIB4cIOEKwvlCZTuTs+nUYptdSfA
P2gkAxQGFjbztLXEuboUExvA9P6LcXem2EcatgAEQ7YG3/X+qEr/XzF5z9HjwTUNYUiTBFaSSbIF
Nn7RQ8PJ5MZtAX+JVe17btwNKny9O6k5zMgruZmxVDyMNeMkb2cG2CX/z0ic5kOmdhZue1vf770G
xVwgLTvCMIGy4Y+d650njXCIf/unxmm9z4ezya52UWP03OPg9m+ipFlTzMUPVhnFUVwjw8stLxA1
7ExiU9hR6NMLgUqxAg5kTasZZZ/75qAi9yubd44/xmOs6XskOtHm3fHQ6wfl5TJ/sQELnKjXLAe0
Ne/28OIDG0z6XvMjQ9OWHOmu5iTo3knl4raaFbDOyN0yJbMt/MR26OQ+cSexp49TQegckeXlzpxq
ryuEVuPhgSs5Vg/j8ugo57aSGDDXhUZl4E25IxXVlhpcWt/zGFMhlPZl9Lc97/cbvXyw39beso7G
I+RpzssriVYxSNHW7AWDnwoEMaVsOVg4uc299Yt3AjuwrmhpK3nw83vkmRLLvh6ryWavoKdiHQTA
250pcbrmXz4pDDUti3pH7JN2aPodSFGcl+3uKwqOleWEvKFvi2kTDenPtVOa2a26RuCLiLtK6bLJ
fm6NnibjCTycN9fQQAoPpT3E/QSrZI1XZ845LAgq5cHotd1Dj5PZ6cYkYJXpcf2Ic8DUeZkQLbg/
uCEH+RTOMxM+FEPz1aiFDeC3nccicACT6XdCnxEKb5oZy7vh/xXu/sfrkawGoMmCfo7lF/gDg3r6
eulmzN1Af7MEhkLDfWw2h12FrN9gvQ202Qs1nURfbaUPs4eY+rbaZQUaiutkp4TZPG0Y7kcyX/bU
TwNVmy/wvo+KCqLcF43B7uXzybLAkVZDJUOWzenS4RP2rngq8L2O4G2tnZlJvpnMuo0yweIIvtyz
8zl1SQ12IfIspf1tEW6847ENj0k6Q3LV1YdXofq/KiMRr2cSMF+KgXKX579y2ubyBIr9EDmPOxhD
bb6eWgoeziki7T5BUCOI8pNshjd8X/USATgxKvz+FuuuxtabIjrPGpRgZ3k9qF0Qmzb//NSw6dX8
U451CuFAqYvMQgH4zqilBSCWsh0T/Wgz6u4OjZIv3jf8JG/CuAhdPt5TIl2zD+ImzYn1WkEAHXvw
rn81gAsCTo9Y1eHy+wz+t1mIV1yJym+5wLL/M2Y0zL+m0j8LWMRimzEPDvcycO+hquRHchL8NGbf
5etkHAxBWlS45Y+YmB+1ydTFfsGf5AebhnGw6uJFbCdhNcbb9Z40mUTxzheu5WpAoOhQ0l9Cq/R6
KDMXvz9OznqNzfKncfXTr1fKsHFxpgEc0TMGatEwzgq/Ii1KqjyoavtQGRcKzvvtxcns6ubA5Td2
RmplY3WqSlQokQmO5ptgykVn+G+fDP2YW8E0FAcZdWxfMcpeg6sYYAiigw/rbFpE9vbU+gjabfIO
P2f6xh36Hz8e6noA4RfjqxYkdV4Vcy0mhkkQtAHVlxfn3tSzd4FDB3JCyzfNAzSGVUSDK9bZGy5C
dOdxVfLs8bIUtbwUJISEUz91wz+P9XHooC5Cee6W0qF9HqEpLRR0ON1USzwAnabRlJHWO88Zur0Z
SGjRGqQv7cafzxz01113k0JRLvVAFR5uTDnIa9Dw/xkfAM05qglcnhfUd+QWdpJmVCLJ7E2HI8Dt
a+XfjoHaBAvNIo5QIZ01rOymelnDgWS9NqHtnWyPYKNEFkRQFWU54Nze+uVBaY3/Agc8ASiOh4ef
2Q97+cOSuuADNGls/qD34xyYYEhgG2hONwlqO0mKVV8An5Aw9I4odS76PUhsAgyZV+E0iyozNLTL
h4fWBk78PIOBtoCnmxJRjp1ixAMF+Edn2MybtijkaDYBsW7FlPoeQsg/OezRgohx++gCVMzvAimF
Q7ULc2//npkYthaJzWTriw85JaZC0SLESXyoqnexTpc1IDzLwahVRq2MaF2SNRoH0F1cFlWA7QVN
TsaudLsJ/A2vHzK3EJOKdm5pdr+WLZIdZM/hsGchcadQgfwmOz260MbJFS2YMkHrdYR4xHFCyalR
o7T1AYen3xf2UIu7yvp12m7v0iqvgEfqPoKu2la1zcqY+opuIDMQX3vU2aFDJxWnycIcD+p5+wit
iiPESCmvPA8q+6CA2jUWNC+4qarE1PaJQ3pKqFQcHpkmOoCLwej0AEgvhB0MDKgsC81iCM1tYafi
1YaI53vNZKnMgG6l2cVbjId8wGXd56wCmdlgQd2FEtLcMK74oAa8V0Upep25RdwTP2nxBcUD8Njk
Y0S/x4x68O2322/XBdJANmQHYtpjPW+f84xBYG3aF3STPkwKf1OehO8NQyPxn4F+E65yX68yP2U0
3NU3QEXIbJi2S/MyOPLyvF6DuHqUVcVgkaWG8+DHk843Mn/MUllY2zjJyxjgNNF/4f5PUP97P6yL
K0bIBmQtKc55JsT1UQCRAYLyb4tyywOS46kpCV2p2w0iClKip6HlG4qnTBJ+6bFRCbJR/XKCDITl
3a0rfbQuixJ696+/AupeZANlkIdsg1/kv5bYs7DSSxozZ44vAqBeRys0/JiN+i/PX4VWoJ+XJ/1i
a199UH5ahkd80NuKNhZDVwL0w2Ri+5slsM1+H5kGqRGpQ0pPGtzaBNIKFY9gzTwixeakvdK2xAQg
7mIn6wjCZl+h/qQCf2do4xHO5Y+53ZILNJJ18SKiZtTsLd47KmYRr4OgmaCMNiVfSOCyYkLby2LI
C7JGye1jPc4L5wDkjYp1SWa2mtFP7xm+j41dU8buyXb4us6NrWXtfbtvs2t1Y+RxJS9AZKbUSztD
HiHx/9MjFnxHnzklndFmtMBX5sClpKf4zfDgIjOEi+p+DCOTHuppCoGZIUFxghNmNvVIPZO2tDof
NuKy4IIg6MSnX1q/R8F/d87v5zlqTNCRHHERnTFyo/c2vDy3jLfi+9J6EOt7EHM6JY4fQ3j+4fxU
pm5PxGKFhn4hfY9YUVsquDHxUwbC4eo3CvX4viOaWIepng6+B8c23dzrDI+BPF924yLL9Odmptwm
Xitz4nI/1Ye8TdAwIzP9tbgI7giqYS03f4/dr4rHLJtZJM0TcLyBfVFzQh2WagJw85XjTnkJ7Mt9
BBEN/9G+gtHC2GcnhLVt/YHaBLCHgmQtcIPwe/pXBTnxysrLUReDw0DtuJUW1/Ayc4rP0Lg34Yh4
r5g3TOM18594Sr/dzWOMgT+IJgl/GBqtZeav1ztXG7GiYeLamGD4wng6wy4iA04TTDu6GfE/Z7rE
UgpL9HeYB+p04J14oJY9xYWHjCN9z5VLeGjrqCyv9Ag86yDt+0PkV+gVvxk2BnLhhqrQfkyuXImK
jhSe6fl7IZ2GwB7CM8pbiytWlKGxMEczZLKp7C3bUvBhPqf1QjLjTzW/0Qx3LScUCXtUsF5fplQ1
gYnxY+SPH1/0AY/Ibwq7ulgvX9A9s+Wl67Q6lnnTHYykGjJ0/wvD/RUvTJmbT2EAvddbSulcL5ZK
SrSuO2/wd9zSIsa8Ov+BpLdU++0U0deAzadYknn/LzQM4YZSVDg18D/izMJurwvoCvzkMsO5gQfY
FM4gbxPr11Vs+mcZ366AFwj4ty33E3h12WaLsrlGfeG2qsPB7kKmUOA4yQaqOi1AuhBEAMRqfbBq
YEY6tkm18g+32xKGe1lqpri4fvWZXdwviLZoMbHpJ1vNe/4q8raQ6JdAcxSpdJ5lBO7S4+DpuCs1
Oz9WEakA//koI7cwJb7k5Y5GI9va5c8UQclVZ+opTzM2gYImCqHgLTIjbdVSFYROv5o/WpDY4nyS
euC0yz9zgOUF4q5ru3iUgkLGX4Kh30cuUNWkJvwbTXrO81BS0ImwKDgE99O9ZRcccKYHbSPHwjyN
0ddUjkGZI8+iNvXnKIl/9RiRq71b0lyOpI2ikf34485a49N9tN4JhZ3pqb/RIofE2WtfwOT2X7Wg
FJPR05/TL6ds/SvcOT+lEnC4Pb9X1/JUkHVPTfPEtIA17FnEEenhU7X7vLC8a1keHhhycUdkxWNb
1BtPef1r80T44A25FWPGdggkP0F1PPn2tlOKTgJUiSrwdXdFnZghJQlypiy6Prqz0n3qL55qhu0q
Mc6Pra8A5kxodqqiIpH25/hK5C2sRs29dr6NpNSKV9DilROBKjmRmXBtkUhVGw2oPapPxOIeXSXz
ZktUgIgM4y/fOlhOtjZbKPSFygwtJ6PtVeTmGwhBxNjyF68XZUKiTsHGD6HMrkNM7sl3rR5WcKJz
wulprG0q0TRYRWs2MSUHY+3gd3Hk5N8lX3v59/DEE6ad8oiMQpPvLR+xXDEEtkSzLPeJlSbZe108
VkGnjs+I537iNZy0U1khifM0gdTJcRQQFqVyyuI+Oz9tOd+0JtHPsDl6O+snu3JWozKKm4BdlIGY
SnfS3rqlmh+55XFVj1xTOzQUG5ffujXBj0OeTydMrM9TgCZyS3Gh2i0ZUtXIqL0MLZr/5lozNsQI
4kc/39mzd+4dheUhFmMisJrKX1j465lif6wELC1wSvhs+6wgNNz81owamUiQupgxOz+OfwpPLT63
YavjqQZ4umx0tHRTwVu0ggb0Dpe16UI+89ZEb7n8U9keICixB8vVcOGTL/McA4Ba+3r7bIawk5EU
x2jM8LL40B9aN2ZyLIJYBEFlyhFTRpK4reOkOxMi3Rllwm6S4gSkWFyuGmywPwncD3rJKo7oX3CM
xX/q/l50G4aea6U9u5Kikyi7mvzhISpjJzotR+KDyA4TE2g9UNV0zpl+jdeByr4tWwuTwfXF22MB
dKihZLeWWdEAaZ28Xmv1xrm6w/fAYzXv71MGtPxzGnn8W7Fs3Aqby3scZEyWcN97YOOmZt5PCLps
lxmNEltnvgODfQqVDKRMJt+a9wBgxRW/3zopCzrgUjd1TbGpZPM1DrV1FmGYWjhdeRq1DPfty+Nn
f39zj5aasTZRqgXGS9ri7C4Rr6bysS/MenC6Ed25ssdwqJHEujQI/61UsIh5q4kBJydXo/sgNKUk
rlv5aJMtlJfsfS8ZgS+L3pmMpA1ESFvfHCESstB88+/n6LZdO3BlBs6C4uJacuZLk6XC4ODq99di
3X8WerAQDM0rDQ5qWP0MV0/BfSljHkmBlGk10OD8zqvqE8SJkehUyAsBj9cuLUsme+xirZkZTF/4
ma9dOYIuy7MrdO98LGb2wmbmT4ejm15LDKpWWZo3oZhAyAgCQfEJGZkugbyyx12UYhhHwMo5yXWV
U3Q5EqvvsiR9oU63qfIB5Ot6807WGjCD2phnmzlR8XfC7AkAhjvZwCw8g61Aj03Q8XFXcGZunbC1
Yrusc+09BHlff/hX2KhFPOhzL96/K7KHenZJXxtPNt9YoZNPisYEbUjSI2lM20rJnueXpTPEAo/J
4ahRWJNntFzMPLOH/qqvSTua1GJG4Bp/UPP/pnrwOAzc92hEhtEscY+B0uC61fyejiZ79H4/KBdL
lEhzvpT81jt+qnwnynCO4librfw7/KkPcL/Iy1dVl8KbnE0e8zHaNBKkLKtIh0Ly+OZw00DQseVO
fD/gukMY1e/0qnCkFjfWnSdgrnApMKEqQ3UFUD0fnspW3oINtfl2D+tk0wZqJ4qV9apgeqrcfInN
YlAlDksoCO2Yg8IWj5p5Z6rik+KLu4VQ/d0z1jPo+bbGDcwWV1WMGgSm+xRFeC82b1++HiUfSDPW
tuFEb+dsnu8wEzfQ2IWk/boUsfQ5IwOghgQAsuRP41f3CzdhEAh6oalatEiLzSeRf0h8xr1zWhWT
srWXCm0mT3HQCI1efErQgchbdv/oJN52oWBKwyn+3PEAOCDCSs6eEXwE3UQc/wVZz8EtD55+f+jF
f+PqMvgPIlAQHXvLZAdaQIJoi3aBZHyJYcSzKC0AQ2pEeKQ4zDzpSetDVtXN+yXWVbk6DZRNNyYa
dDSyuOgt4+oP88OQd0ZFkpd8/KMOSwa+D6hdpoA7FfYQJXdMwTlxDGdPSt3pxcojOPzkoN8297q+
5F1nMflfRobYB+FUJrwfBDDhzOtL3o2LDgXdj/56S7PxraCXqErFXdISbjR5a217li9FMomR62VH
MKtnZUoEivWIJFXM3hwq0YSxXCA4o2nSO/5GPM2rN79MYYi2njD636FBxf9nsArfWd5/ecytOAsP
TA0tybBVF86Rex78zbb2PJ3+7iAoA6mRVZ1/nssCw/cF7Qmu4zwh4lfaGheVAW0Zc63zQTho5Ky6
qk22zpjdA5oPaiOdPqEGnHZFm87ngaa+C4Gf9B00E73mXGejZMLQfvhp3xjkD6CXBmCGHBmWUlVg
0Ch8WeSL56pk9dRofEeaD6MVkm0mQRxo1cgiyeQkX7GX5U0lk3PRAPt1iO6cjOdglVJZuyBciBFO
r7rYg6xBBU2ibGdvSoHOn5EDD7GrjCksAcoYDaJKT7B/FzIHIlk72OAUj/Jxd+jTFLK1LOe6nECR
tUdIWWEIdxMq2XaESGk5xu0uFWEBQTgp+JLT4zTHWSRit+rrQUez/WBSMYy7ZLTOEKSyAR1IpX2N
+nXQO4s2dRU4guVY8u2NOBtRBS2a8zrIGU8chQ3qVMyWJhjCZv8e1y62PPS3Y5Yct65cQetS/IgZ
m8gs+NGL9ckXhHdXBQuiigjOAAoRVxv6mOtOKcOhS61Jv4xioVouYjbnNqtCoYq0GG8nuATObVr1
fsIbT+SistSDa857yq7sPNvBqkyhNH+LESwDfgbUqK0SjiOLnRdKe/+TpVBLcAray0twvSNSiIvj
uJ8x0t3TowWUANNu3e//L2eocV5J3V/pjlblF3aB7KwSOLRraeh5N0xLafYNOo8RKzuD6b2oGsLY
vQ+R52qoluc+5YhDdGPxst7DU2FRPwHy6/p/T/PyKBziNwb5ktHfr0jlirEXO70kaW3VkLHMKhxX
Cr1lgw9gvKErOMx6saeGkcEyvJafUOscgxtn7AtifrcZx3QAUxM5ASqqJAbn62RxAeged8zv8p4X
w4QJYSkTDL1MejNSOh4Kg5CYf10KGyhMj9OQxrbRIKFyPVWk7lskPpdJCWkbqYnfg8d76z1k7i54
ZNBKa/bW3Sep1jpt56pldgLCsrX/z7wyvS/gi8ZibeGW90CEookSZceZZbDc4/jsmy5fkiZSPcHW
WwEDvsE09IjTejkAEyRtIhAYKYG8bB+MXPkjvr0WX2kP850n7B2R76mle1eDNBugLCdjXe7lp/qa
zslxGoz53O5e5zV2LrpEXVPMFoKFf9vqw03SR4q/GNswTF4pTKZJ/dZe+/p9plXd760cvNN80ZEM
FdDaN2TSxOoRaPLmSdQpDeDtLJ2njbAsu4FMvo5lhQ8hAmgmCR9YPZpgGr0g0EmtXUVo0p5UNtEB
0lbAOriciNsqFB8QdlKrXV8NL8xvTsg0qnCsydR8CyPNHgrEkTJtypUe7NaDYVNGc64k9Lznx5hv
NmxEPuM0DT7cFh21lVbY/6WZp4KbrI6NoHWJaOzCeggJC0Ea42Lj5hDEx4C9m9JyluDrY2BWi1Sf
iALON1D8attdemPH+Ats7+gIc+f9KVsqTFeVn/fZCXjAzAQk2Nex65bcJZBGnoGElGZwFV8ROE9H
WJKb0HPJnchjcxgsHPxoPfdAZDfL0vUVVITdrHww9QFr567ZpwmJBiiSTnIuLeoq157B6dmtajHq
PbT2Yn0kLT5H7310/rQqPzpRLwx1LfGmwzIRIMfE3SfmpyvfErfaWJnmGd+T819HSdZSDyImc1ah
zz03C4Npei7sTdP7/DIXyUuPUcmbpsWEyC07vgzRPwcDnPQl4Jy69IhdyIkqmAlsKCPFSjZxNnJV
XbecqwjxWdb4MgqKQBDd9GKbbH2CcMwDzjrZK/PuK48F24ir3lY/Sdkgelc7wGenyj7SuFwB3EBY
NxZYX7TQSbOct/0IljGEgKnKNZfj72g5Nm5v1SRKt4qHOKVf/FYaFKXtBbac0ckqac0aY2JiTe16
abZcqM4x0FdnDrhFPNqxw8dnzCWeG/2wz6otkHq7ACYBUmrzHukgED9BrQU5UQ5rN3Ju+pxcb4Vj
Vw8gXlUb7GEG08j/RYSKjZr7vtfoObNfgh774Vma2hz6CFhO1ZVyKgVbbS7K+mF/NxadVKoKhLZv
/3NT0n1HKfIvtrHV8KJq+WF3Yf1G+miy08iI5elxeHbKeYu4JBls4GFC0D3q3KKaecj1B1DOaTQd
sqTCNuiPdtnZaflGEg6qJYMMbNWeAIOOBjgWgJUUzKQH8eVnNN30cl+q1yCYd0ayRC+uqE+FuVmp
tqAACKkoNkc9goaYV9Xs09EZciJUuXMQEgj+y2lT4fu0ttAXinqIK1AXe1A+58rkjc7Bvvn+iSSR
2Oima1QiZ+J9zv110e8/9/xlAnC9nUrBZ8H0qsbFZ0fu7qIOdFJmTKPqmrNEHU5pRSKer98kDpVC
6Y56mI3yeqDzuabj0AgHNycRKvbeZSpns4xxruLjIyjdFdPrwrQFJ4jVmIq3a+1nAarEGhFBuCjt
iGYVdogAKzLZ10Ixj52BsYG2L+TC6k+XXCrDmFDP3YFhUmr15A5rk2pl5qT6vk+jEdBKmvdK3pv8
wwSmTZ9Szx+1P41yonIrv7ZoI+OD8175Qw2N0hoD+pwWSF4SICZA4vYzYDmzfez+Mk0Mq7ErNxLY
qYFMK44IoI3qeYWb5EhNWofA932rA6i/dFCkKeVgFRNo2oPACahISOkBIe5e9S4DCw744Nn1B96h
obmb4y7CnSYzr7BD9ZAnJCFJ6aWAkbqWs1M+dbACOrWL4dljPZrcUmad6vy3phJRX+3pfDpYX3f4
NCtSJCOux722ecnve9MTWvDCZNdMOR1ukrFDZrH7pRx9rZ4wCcI6pnCCeb4mVIFboPL+t+Z70IVc
QrV+lepJ6rH363Ds0xwII2r1185gdjDEG7eiDmFdr7qDKPFhygdNxX9t03FRwKIThr903ICmjpG5
7lk5mPwczjorZ5hvlkQk71rE/e9mbsIz2qI2woFUariEeXOanS9RT4Ay0/WlAoKxHu70gnydiBb6
DMDySr5yuR6L2HelHMiP07DvVHk0k1D4I3TanLwUJ72/urUebRKnk23k4o1t0NBZOtFhBlR4l3s+
MVZjcY0ZL9HTkWTISeUmTelIdBi0/c1kGZvQAq/86AX0+xxs3+SFFekLg8dv7xmhsdNtjGkUc9yq
YvJGn5vmkXPyvVy6UBnpZjepnhCRxN1nEpCxlVJeIHokdjOTGwjhAEUJuvm88lxPTY1ix12M+g1a
CXV6DdnwlQJHhj85/RCFjIrm/WUpKnd40BlRMs4Vet2kvwYqHchCXC9qQXmRvTciFCMh0SY59/CO
Sm0/vm5EZ44KceDQzz6qUmZ3j5buE31QEWqFYtyaCxDnGvKxfSHVmlzA5rQEJEI+00g9UbjMYOTO
NUwYeCQza3vZ3BMoj1LY+wVkd8YIf/qQB4/87rB1j6BjES6+szfVFUhPZfH3gSwkuW9Nt9soCgKB
EHEte+2lKV+E3nBS5fSZAfkzXg+EDJFd+v4nyh5Q58qReWfcfHsf84qjlsbuKMRnjWLRC6TpXZJD
RS5oc8Exw+PRvfwSFQvsuiP6jcpuyWPm5B69cuDqnV+ZkdNVUdBBU1mpqzxo3w8e2cGfQxdk8bOz
VEmHt0oCBZK7847UHCyFFSjotEGRQ83g3pk3dBDewooDxeK30px5/RPgUgz9PqM+IMC1uhQ/og7J
aTAq/ssGqEWusaBUoT+X2PXl4YdCuQ/8KqFuq0+0tEWJPZG6UcJnWdUvXKVbtPP5FMxL6GogkIh4
hYyiNsqbd6bK0SLHugkm0W53J3whCWlBOzhGONlgZRUktLHhaVQ4qsYXqBF2T1aEnn43JgkDnueQ
ej6grFYzVwh+LUryKkj6kWAddBsMf81QvXCLSlZhqhSuA2qwrg53nbV9wmXn55mkpkRTbwbCaw4l
N3aqowXqEQCVGeYbMjJlBbtX/HwtqBiV+Mw8A8UwqWE4ZPkhMsqup+m0qGGa41aUbLepbA5mPTbG
u8YvOmMuOiPYbNMeDzHwiKGhjyArPQVmU9A1wSnNkkenZEMfnw9unl3+y6H0NCNEiREpAD9ojelU
mEIFDd1CpRYbfjOiv/ZzngHokccXy4XBTQIMxs7Y30+5z7qtNNwu35vMtzLH21uIVmRYRAWLNR5e
QHEw/Yn3r57R238xg77kuqGpGDNTAQBfVuld0WjXZN6f29VTe/2y0fCBPUzAC9QwaUMs0dQKWiS+
fiyaTqkgXEtp52G32MjWoPXOwLDKTypRfHGHC8QRobXBL2ZlsmGm5Mak4TO+Txjkum5eEIX6add0
dD2M5q7fB+WcFKMHnfox4vU6cAdskiiWigAhNKkGDwDZA+eDtQNbgfA+42p2UsdbEMtLbZG0L4os
ovB7n9G7pr1AX5xA3jBS3x9tdLfQdgAyfc1uR951YESlip9U4IEOL5ZlmGHoQjl68abyGIuKF8Nd
z+S7Yd8KCe+Y3PByimwt9k1p/0ZS2M5jGiaSDELSMj31oqpB0Pd2b+czQ+YNkVKrl275UkvmXkv8
qweTBjf1MZrKL6Hr1WATJCRVrTTpSh4eOSTsJergoHWyUi2On2Kq2XX2rfMhWodqMg5hkVMi0sUv
JwOD+bDnYOo1FL/jhDu9PPJXrOvaTGQfT05B6tXJ+FpgTpmUOHvr5p6iSCP1SFTgErKVCjqSfOd+
ENV5bfGjyULeA8Cyqmh7FiBguF5jxfnaJCiC9swEYgDpdZ9wmW+gV0FzHWiDw5uXtwW6IGcT+aKp
AHHGPSYSA3S8aSNiGpueErrJ0Qfd5aW25O4oiOmHwusb+DrpZKpLZzaQX/RHkH5JhS1rp1vqJn/w
Uz8GitdlrWL2e4zK/ls9evUMW9C5wMlg7Dn2etLj44y/JbZm6/C9AUj526PxlBDErRcUtRfvFjUK
7TOG8ddhEkvzef/hGin0d0Fwbg7KvtiHNQll6oCUUL0L2Qy3xc/Q7dR3Ud5gI5NU5XeDvQXyhs4j
meV7rkJqPiRdZqYDQLwuvPVgrwqRTYbJWco1kIsy5XntURA+ItDqHHaNmYLbKrmkIYYgWL46meRj
/dG0/Ac5yqTKkyuyLvOc7c/SCRr4NVZ/l8L/JDFMSr8vOA40hH81Jvz9mY8Lfjg8jq6j+gJdy1d0
6dJ9kV2AZjEE6/OuIIOioosY38FzNSwU7ZDZUty7gVIu6aXj4bjaFJJp3XGVO7ZcZyT9+1EEn3NK
DvsELolDVLgMrhXpbSHIGgW3qaxs34sL0Q7rEMGePIdTVdD/VLFOXGZLUw51qqtBki5u8v2mcSaS
FNJkC7f6AGDeq8lcNFGXc2Yyj90ntlzcwwUQdOpGG97F1r2nPQj5X8pBMj3plDFzqBbw2j71ruZC
WSnRyVIqHlzI185RvaohEgNtsf/l0/0A/q+g2EUw0jtKRz1g33AGZiZWsQxNBzjFZ1LfOHkmA2v6
jGAxCDSB47swFqLCVQkPvmWVmbK6nhUT+8U3mzf43yC+p/mi6Pc9JXPfSSPhN6vboMc7OaMbBf3Z
Erq170xACdVZ8gF56Rg4E1RAuunblk997TXZ8E7uVTbNFvYJwVTgtX6f2DdyxMwajvunloXTRiEF
QE/3Gfd6Vai6cjFjhlKVWrMhyEB4H8NFDSpuJI5n5QW1azmv+RePXKaSUESiTEo1EeuzMNMRbebY
BhGWw01m3BnxrlF/YkqKK7XraCXFt1L6ez5hnaUw62LVQQfztcC76LqC6Rd/s8HLH2S8uNjoUQQX
vU78MHyNJjPhRjXrsGJzCufBJwpXIVtZWMDg+jhjSA+fsfIKOPZDPt4b0f96GcM7lFDSJc1zBEUc
MJOKNGh/uzxNnXyHJCN/32451VDvoPR9auSHg+byrAvVAKjCyU+BY0/vmS+Y4BflsJEVjDPWACVp
/e57pOnfN2n04/RiGYgfuXcBR/aJco57EFgjGq/Bp4eF45Van/jadrPXMbVoL0gqM8ugnXcaeCj9
rl6JWrkC3jOG5dd8QvvHOhiF2GMpuumSb+eU3iNg65u32IxE+YgzIGzVULC7dWnWydbJLgWp7Fu3
Qeo/EjbqbyJD7OHnSS9DsYDsG5tCgzqGx7/HrNLP+kEFzK6pKyCNgEI9LvB8GTVJxc09dwVCppBO
yNygDml13GyuELovT8n9Vov1R8oH9DRPqqQ6g95QtSiLYltXx8F755y4MrieQ7+mXiuBZTxFIJM3
dPwtJ2HwYCJnVHbucu+zN1l0DJ2yJtbMK2BeJC9LNbVUxUlM0fv8/LU4LPfXru9X8X3P/0Ay99Od
29FmwLR63nTmL499vDA0juxOWK29l+2SaHzoMf3aPjERwiNaHyh/0KxsfZHN5tdmYxZL5bO4LRNL
aFdoUq4ndEjhVRgAa02PvPUwSJyhDA5xBxDGVl870ii2doHvq+XG+/uDSLS7qDeHdFE5gHEfj8b7
knIsRJZOkW6eWFdR1XXKu/ZVKRD6OcRCTu6e0VmtuS3sWG79+BX+WPMLoY7dJPkUFdmJwQJOLIR5
3dewn57am1f2k9ANiggUpdJy55yLriNvp5vEGdyphxHLnwVOW2L7iC89fjk1wuWsx+unjyRPfN/B
9/0Zjqt6ir1enN/U88vXwhIdzKReMY8crOflWb14T+p1RFJAOdtkgrf4dqyk1RW5DsRVSHa6Rqid
ZKgD5Y/Q2MCE2SRlPGFHAJuezm7ThaJ0ZBUflCTR57vjD2RzsEuVgSylmZ6/Qckg4sdfiI8vsE3t
OOUeTSdtgBWLT1uFY/ae3IKnsSqBtFryDTp5YuNNmswsYxZNTRAgNhK6oDZSowQ0YCXQ5uCjPjhb
UdhPtrFIPQrCrjtJLXvSqlEBsvvs5myqp1ImC6EHQ3RJxXzCkHWmLRhgnAT9FPr74r4YEGTyovAN
bLRd4kARSoMc6wUX4OclZX+jBns+tCkleWVEiLYRDZ4K3QiBhwA7FUXa2KnPZBq1gZedeguZop/L
NL6mR3nKuSxNUNcOA4cez3EBzWMkEfXBgQsgBic+2x7svbnadB+nZ608fPKWNnakdVl1qJYLqLWG
Vrj8+hoLnnETHrgeiDWaaAX+IU9r+D9saa7LrHVmi8K2ojNVSQCMdIPOL5GApgO0zqz7VhCVxNjZ
+a3p9vVJmmUtLsgbJT5FsIJlyf38bdEsgWVmQkap54l3XR1q1qiT0Hu4b4QoiSwBo1it49sbYuMm
b/AJR3h8NRFb8fVFMTuCxMSpZqLzwLbLU9Bc6EodwlZvyULEjWFO3aa2DU+N5uUMR8V3qfrykREv
xYYZBElJN/d9Lf1au4WdFyh+MrriUqAqcf5DhBe1DgeKKICqKWLxGhNv6hc4vGqnmbMCkWD3tm4u
u+X6dk8I4DQRgSoDly+efexQtkMOW6t8HJsuqRPXXRoTXJoAC3uWAtczFXRItBhrlVITCFfNZxBd
lSHL9ylzgtz6b2ICTYA6dum0S8R76nx52iZJzwiRLvH5PKDSjTnXZ6tvI5cXpjdLC+OJn2jiajyP
XNymoAO3aTkOquhQ5lmHr56ouNY/hPBnZXU/dkTmbC+BUmSom1XygTvO2mtvjwTmyxIhwX1hCNbH
zVMkrxubUb1wKRR6Dk+Z6nI3nRvorqqYqHwWIlWRMfK7rmgN/jhXO449OBftdS8Jddd9+aKhpBff
N19RaUtH/wvxigu60XkRMYQ3mcqjzk1m+YDqmhgiPBW3+ZOdRgF7xgtyfMGRq2W+FozZ4AiazXwq
LAV2ZU+t2peK9335rtYNDZjLTB+4d+rPTrssDbelrUvxg7mqR7baDnpBv1FOvPN4fp/nU0Dkmrrl
ePCRG3fWfB7yKZnyZPrlAk4bBm95/2SMzS8fgfsYxqG7aymVFJ7W3e9rpRoKqXgPhomIMWHd2hF9
lRgFFlHpGJK2Tgev9U/90NNZ1FqPK9Gh6XKdvkCEt4WvOkV95aKCuZQdZOsKKFCdgGuQIdyAtrHX
W4uagZq1kVxZsFj1v6P0Sxu8xHIMgIqaEfLkwQ0JivbCeVQxZh55hkThg3expxqv3Ptxb4ew7Pht
WWkkRlaoOgdQKpWzx4lxukIHsMGs/mEM8XiYSVKHEdKJ5HZ8u8Np3/Z1pEH9mH7V+K3cCM9Leo/1
T70RJdCncmrAy1nXPdPMe3k3vW3Sv1IMI3M2TujcmvFfVvPZZi3rUbA20i5xa3CkmtiV51haRjSa
8hMru/Z6vaQL4bMHkFLQ4c7XNNoKIXoFmn82Dm/zMau3sYAkMpM2lAn0K+Sazks1TgJ72VCyye7+
LOsfCOyZe6jjlwWo7GBEUGnsX8/vxWIxZCG7uTallHijHYpINIaOSigLzrqwezOXYC7ryRtRnKFT
wGzDtknxIaF9ZGhPljWsm8cW6FzvaDXTS3w0UflL4O0wcOwrLEff8O+1/3J23Z35P/J2b0gS0z4f
noKAeLFDvphGRPx8EWaX5HVazhTHm0i+V+avf6L+28ZDaX3l+9UEYcGwGtMLYqBxNjNWZ6T89iEs
gw7DN0spsZzrhqomHPnXTFNT/qd5r7UBIKs1gy9G+jVWEfnX2UtU9g0PY3zMuiXZtXhTWkgOmIG5
vvU1TXHMWskN6z0Ako0/ZfYeKEEP0iAxCtqN4th0G1cpg89sJuLKrXmtkIKV9mQbxnAk+cGZcmoe
oVfNHmVfs8Zs9wvIfo7cPMbGuiWvjMD+X81c4VvD5C646nq45dKLZDV4puN7FG3SinzYHnkBQuY7
Lx1N0H9YCSgfg2cBIRnZHpU1lx2kbX7Xp345IotpqdRK/pnUrhQImtfwOQZWVrY+U0O0KYBpv04/
lKhQcDlSRNqKT9yG+oLEsmm60c/cf4rOJLgpOMWKrt4tw7gX+TBiabNhfieRC9YSiSGPNJ8eRKxl
MoGmkLaXFkjzSPtCdqv1c1E6UDZFS2ZVXYX+QYTi+UhdpubTd3H7CRbRxcIY0Pg6gzcPu/oSpAxG
OhdUFpDh4Woq7lfrdtkbEOhZqjRRtj4xPh4rgBH4EzvRd3yuUZAttjH1PyMt4aYM7mpcvUQ+QOWX
t34vQKXpbBt4aawKBKdwTnJQSowve+Ko8ugRNH9eFjTrZAhQ8k5239eGSyOb4lkAveOzpbrPMMOH
y0lvSn6VrioOWRGX4wBIy7wxK5JezTKAx/UEb2UDpcr/TTmGJ/tQLSrNqzeVdwghTSZyL2g73WXY
SAayC9Z8J+bhRxLg/3gIohnGjP1zv6jty76ot4aP5R8a7I8YhLbg4U6DZoQSlaP28pXmv8JrY/S4
IwX5QwowROBVI0Z83iNRcwQ30aAN3Xs68QGCUh0MKIjdRfTi6sKEV3OwS1n0C2k4ps9CqcfBwpHH
Sk2WUBrplvRTl+xZL6HtzFlzUBAXlGFdxs5a2fVj6OiYmMmRPV9iMVcP7Ze3dk7wrUzIP8adIzFI
4y7g2WX2uHACSPXqtLWKj8QQLdv2Nq69IGd3A3h7BpiRyuxyHc48FSE9WkpUIGgYhMBVYEotgugs
KgwDzsnzTp/asP/jOQsntk7HknnCy4Fx/RplodohyYbwkSrnrogDnjxoZYIXTqK9zLDEx1BsJb8H
5AJyGVCxsHWm39gXjpGZV0e1SUS8lGvxiqDs7PuKjqWFlv+TIbFWU80ruLLT3q2+3BDef1Wdwqk2
VIRkAssY9VjPaYODKxpHo/KAMJQu9U0UbzFAbHo788dxYa7LCWgwsmorKxjHHM3TKW3MA486mcWe
8ww+qj9Jnhc8JPlNrefzE9ciguY+B3Ktxs97IUc08Trptcd29J+DVohjXeMkpPjd88gwHYmVGRAQ
dUeqn3YLERZBSZuY11dhwhpsyk5v277JAZWkQUpo4dVj4APbTiuU7z67wQ9mu3Uj0eQRMfwgqrqd
0yTbCihiwjDkAXu+BUL+S4jsj+2R6GTpNRBvpuFws6WzYJkGwudopImVoQeIsnqCV6mxy5V4MAC/
/f6cx6pJDcX/F7LBoke4Innc3/wBlVsmSw+cZsW9Qa1nPWnqrEaY6cddbQWlGrpdJv/DNtcQ0XZ0
Yhc6Idohh1rNPy8AoaMO7dCpvbS2oDVq2rMScsXGmbkVmu9Fcj24RI6yIGHiMLlTeyxvph3otxdF
bc0xT2fuUUjr9T438iyE0ouQKpw7IYDFnOZEDSL1YEoKx7ywTZLHHmA41nWm/bxYNg7REh4Cu8w3
jnU/hYZZI5LEsj2B+LKjK3YpaCwy/VQbUtcT/njqdu4+uhcFAgzpQi0V0+uM5dUiROvf3fU9Xtcg
BKoRKbvJY6UD/xrF4r6BdXng8kS24jczNwYY75YF9RHr8JQwkkFpvC2xd39E/P9YJPhiSuk1Ny9j
KOv5UkzeQpEHXqkBtTcShd8I2ivjITcGXWyTDooFCYkBxeK1pI45VjQOJDBgwJVN6Mde5uK9FhYY
c3lchxjAwofEehYRGcA2W4NVkHFJv0uQLybdBtXTOfOaPgEFDPknUAsKwarODY7QQlAppzfRFQwp
G2SAtlbxTGa3YVnbtvrQuHVQQoKGDZTfGTNfJ4CoAYAz+hW65ktak7HX3zCSffj4wR35S5nyblpq
dj7e+2+RfxrIevbqHAlIgbEInkK2LdEymfpi9x41HzI13Sm7Ho6BmRYIXjpuGwVaHiirmw7xG/Kh
r/lG3YyMUvGFVWdcuf1k5emWui5h8ri6qA9DUAJH/PzVzxM1NqytGO22eCCrinEQ/LZZ6Ht0m92B
p3F48jIMeWJFhdFYPXQMABxXnvw2FpEtyO4euQSqifmxOJVphefFE3bdA2bV73ymmSzhgO7ONERN
+fxLudICIJ+Jy/o61XN44DGMVvsO9rOlA9YnAY0ZB7WQVKHkrvl9Jaerw3K/ts08ETlT73jP+XiF
5KVsibkjKA8bPGIA/iZdqmtbYoV0V/GSCePSnjzLWNA8zV0NTqGiLpQMTbEl2y44SkaLsj0SYrFx
NsZNxzZ0slEwPCHkXo3KzoaslPyE1JzpzBO0ksVPExHwov+TkAVzZJk743jql8o/2TU6H4Mylkcn
JuEFon9p8R24m6tlX5qudhqlQiW2o2EFcJUHQmlpUrAZVIMUq5CRIm/mikT/ZNpQYTIEcg2q2U0x
nL8bAXe4SfGpJ69BxS4/VmZ0Z4SyVoGykOVsvraJm2Uh+MKr3rsHb517OSrw0Hq33xCJK/nyLlEc
JAWTq8141+Cui/vHJF8pINhRbgJyJtTiK3D66DX+Ss5xyp1xTfHCyr7up5mIPnnNTYi+XWa9tFsn
vTxFBa9VkbpA+zfdOZQu+ACB42LxVowNvOhzVToSDBQLuIQVoOoT2FRJQk4MwedC+ehyu34p+9OG
pog4kFCLY0XsSe65gWFqbs++gpv6Ca1G269lM4IN6qa/w3k9k/TjVbpxukCKAXuaNC8jigVzcD7T
LPy91Pw+kovfIi82trThxOdOr1FACezqUtjXSFKkyYfGDG0D5gKiMlJiiQ53ERqjHF5XwxhmbIZ0
OM1GKFRoxNRXcWWaBVUzXI2Bwdh45WUf+m6SPdvQvJiLyhqyUVtDhZapHH+IUGYI8pzgzxUUtWi3
1Mj6Ajh1rkLodgK/C5FVxW3965BhY42oGudKSQGIfMZkqJc7osOaATJa+klrpB4qitSpFrLr5dDk
IpbrWa0FP9FymLc1HBr2DDDs8pMEi3KHTZOIjzPVDIeors91P6wqZTuT3SYfgmffGcRwneNmS3ge
uierINiQDxHZI/JqWwKSMnjXhwZaPzf1r8DKVGrcRS3akBUja5/EhjsMUXqHZgPtcDOxvz3bwcEF
tVjReFD/T7Jb/RHGR+M/wJbEvrx5clK3V9sqNS/mC1tJFP8B2u+6b2Spj4yZc3vJZl71XVmmfYBe
GWFOFXzKbswRxxArhjNItbGzMCodHwgoOG2ylsghBtFrLXmjlEqFdICf0/KQwImgsSEmdNr4C7sk
G3NsjjPoj5HOTyo1804YoDyZb6Y4Xg8QQYy3BGZce+mZ2V8BiiN4yXEaGxjc0sXfAOwMefPvD2gN
D2aE3A5rLAbxOlty6R5FFMvrfcHzBFjk8yjThnTAPOw7kDyCOfCXgkfZ/DEwNeZTLgfewjJJOFpP
Cw7Izny4PCX8lRmdV1yRH6ieBRIFO76j+wTcl0vsDTTfqckqKgRSAerTXFQ+38kvgvm0yafWFbvx
vendqVnG0CBpcskgGJJSoML+27vd5b064xDnMQq+/ARLAjNi2tXj3FDRUBxrtUzxzm71irY0MmEs
aMXhKZpdm6B/hRiDZ2XWE7JoQI/KiqEUbWh1mrKoQceEktSkrjEH7fyHrxdLLSUoYAPfjCTf+7ic
xTgiSTWDvGBnqgnLd7EhJgzroczwSGWk8OeJHzZ0zt7iKiuqw6bP/wdH2Mwqpw/t9Ukzjv3NItph
6QrK50sAzbSaF1oqNdwmW4t4qeRj4rLR7cH2dK+hWju1OiEI0f1n13bp8Lr2DOA8XtCKhIOaFpth
RWO6BiKlIS5as1IF4jgdLpI06OMYMtsSKlhuejyEqyJ8vRs9yN7wWeHp3VWatY2ujhaWuSRLPO7I
994w3N5KVUvfJ9xfG02py3nwfpuovIx0ZCbfHfmP+pkgS8t5RtogEhiQP07kOXI8ygtuMgIAAzAP
R+ykv0ZawZbzaxRhoQn3kKeJFTI1gC1AkZWal95iSbDSYKr8n73FPOzL8Xns/dDX9W7CR3ecBUlh
r1OHPTBgh5TEQjwsnG+lnE/HiolunKfjjqQR8OORAdlRXopRyF1Kh287nlXlwDOw8sbnkeQTnZ4M
rK+DkwgshIUoE6vYbb8CsZpRClpkbCpKURZVoJ45UggNmuWaAckkKTDe1L051dDgGKNjxJbtTVVg
NrO5MLs6GoVMQxmmFF+5OfmpOMsF/drDvRIFCxbC+SPUQWmYuUvSVfep7YXK8aFL7FwV6silCLNX
fRK3ObvJRVQEM2G0t5TzpwrZr7DHgOb6i2pELes7h+qBrGDoEyf4hM+cfh7N9ltL7zqWKXmns87/
+nkshM1oG/p9RMrParrU/3VbU0Q6Eosm+Y9KBeT6GhGoG1Km6hPeiHYzI9XmStFhADDhlTvwAolO
6Ut+kr5Qzmi17+GVTjKNNSrVT+DY6NlL8NdPsy4b6yxZWsqvCrb4eTn8xUCcIQWNg3KMdsSdFysI
2KhLysTfNwBH5V000v2h6wWyBRkdLwiAZ3Ifz4SBjMWrUJusBmmojezJDcvBvA3iNFn7x7bYpStF
Wl2UOkUD+drIzgY7GyjATRHhliGdDp8Du56mFY532vbnMUo2vre/sAt1unCpPMDSDy+mUlld42qY
N4geNSgkWtYQlGCxeiZRhmQ3zfr3uh/ltqcKGflGVyBeghO2TWi6ylwwEZ58zKpIm79NVT8uC9OX
Jx0Xq9hQ/NtDJpTf0DtPpvrdCpi4bRMaMGMEnvHJj7yFG0+z3K5U5V3lbAqj/Agr6Z7QrFYriRvF
QWuBxutLx3RX1p1/IsCIMlgb9FGimz3uX6js5F21i+Fw2TP45CYcxvkV/3tPxE2GGa3Zmnkg90Da
u/E8rgfwRNQJBy6vIJRKwBWlnR1MPj7hBbKMiLrwNjlzZv91tnjt9W19FNahubKDtItVAGOmRiYU
awc7khgAnIUI6Fpy/+HNV5AylVGcmey+Gc4GbgqR6xJSbkbBZyb9jSyqPgGkgWvuV14fg2AjRK5/
OmYzcgJywt9J5Wb+IRk5xB5rfge3ZjaQUNUJHX0042kfMx0AVr4RqiEL27RNMWSoAVIN0vf9aH7b
fKSI1PQ7HL1UCN/4JNjEdqkHVI7AM7qqQdSevHwBqk+9IDBOrz8EkAmnfF0AG6CO2oro3EnOTRW6
uDNlrZfhmk+t/onu4qiFtOFuO4z8nUDpyeM5U3Hb3meBfZ0y4bGanmAtEHhu+MgOsTeJ+PcPtlP/
X0FsnC5CUdpj9sTfinaNBmr6cWvGjpbV9HpZs1WmqhlOe9gUuRlBNCBUagQFoqOVJqc7wgkxvWgf
ByaT7Vt0B3TLJJC/vpW5GiiHTtHEjYTM/YPCfpcg2yvbG57ctylBLPWHVXKg4FH1ay3C/p89AXuj
kOKMQVu8iFVy+yuxE1tA52gc7eeBAZ8yvpTY+tViQgkSpqXuOvqZazdaGYVrDJqfw06p9eJJI3mM
6B+8sMnnRa7lybv3aRaSBGsQdqZ7tF8zVrDl6zo3AOZv5fae8fGTpqTq1GXkWz1Kmb72Dyhvpjmd
tkgJNzb96asKXQOtU4SthkMIZXlcd45n8xuIRQFrqIJVcuOI8iLzdVacY8uGG6KWPY3eLsMZl4cS
4MTLPZFux5WdGd/xqL71FuQJ4V8UWDlzLplcs2m33rj2SHD2WnYwhCF0nybyb17KO82SZ/+0SrcX
DVNXYvaVyJfXioJrrmpVLBhNDq4nmWNXADWhTtDnQ5fFy2wSmCnE0GpqYkPasfUzxvRtmQcVhcMB
0hAmVaWCZHyANrqGQI3pHEsO3MJghDwjeIIWz/QYujwPmEsZ0y679vAwppgy+W2DadoCC3AfiSUX
BblAGfQUualUJnEr4+01ah1OsViNvFsawgk8C9NSla35vImJM+eQfFeMrzzj2gZFH8MjF4xjltkc
KW+2ozP+zFYUDQ50yir18X1giASqR37BH6+GsGb2SAksI2XsmoRQUL7i6vz3HNheiBnnFkP+/2ns
tX49b514XzahF74bGV+6ry20MSJrukjBecm56OpFegUY/wwRXzlVXSzIGPTw7AkxRE/hhAynm4mv
KELbJLoXdvw7iVFRO9dWKqz6aBrLH/2v7sPTHY6lDXN466GPwjeQXSuM28z+rVyCAkA9syOrG9kU
MjV6c0DY4wPHcc6uFjYXMUrw+7DQrKFs7dDdru58l+VREdF0WckWCyS/jaHmNTJbR96X2qwBPE39
3M32tGH6TdJqxw4UgSd+Y8Jq3mJkqejfvpKWJslVZQ3ba/lVxgcmuEX7unQRc5ijAa/hrF/VQTQ8
nzWDFTLvRxw7oeF7EXAeUuG5kWdMMlWOmoLxjXtPlMZqsymezsww6f3p1VG0UJqIqBofVsOH7Y12
RZsPtS6HLrV1DQPamvZ6/voafcxr9WlUgFJwIIjQsuRDvy0NpOFsNh5HTOwlJmkF1yrx8GDD3w20
IzJVbpB9PI46INjFEuJ58v6whsoBJAHjwpnMGALm9UfbJKTFhcOPF0+1rZmNrG8E+KUvMrkQU/yj
Bb9N/H3C2QGy8oGQuNUUb8otTkgcQOTCEPjpAW0qix0sgogQEPhFzoGOge54sevJgJPH2WIwVziH
UuITHaqBXVfCVLLhA4NWEl9dO9moDHXOt/6aSMUm4Alss1VEPIkAxaKamvbCIm9B69exCoGpmlU9
UrQGPIm3Jy1om4C5bpNVBMH0UYi1Baja+deqDjowQAjOD3W0iWRdzEb65k2upuqcCBYzLn+AvAAf
piCitGRLeKmYY85OdBAqCf8rfh+XEkJUJmZSoEW1Gp02a/A8B0WoE5tf2ec8YYrU9ypPnYRQ/guI
1ZYX+FqvBkLKgDaFhltrs+T70SZ+TePCQbHUl8bCfiY8XFSRraJjtsmAtmI876Im2UUBMHBsq+/r
7yDXz/Lb3dqJZ+LaUYu4NR7DF6IDeZDI3Fyh5sQ57Y83IFDG3YHmWKfbGDd3GpZI09odvVBEp3VS
ohiS96Z4QUapnp5LFgkOgsBGO+XHQaCKWGmilwoL0Zt4NPHE2o0V6r6y/FACe3XFXd9WQ0isJ+W6
y/niXtxufyR6AmoxHBbbz58uMQiFavJdSi9RDaMCnXgC0QMSf7VACJQ2gNHJoPyXEtKHAR696Zbv
vS6YbrhUN87erWHCvxXVLpP43B4afwOqpJp3qu23pO54HBv4ONNfApoipfPZHSiLHg8pg+vMM9wJ
xtW7EgJWxZ/fykUtxkxBr5QuwoW86zwvqdhShCCyQ0qvUuBV5K0fmvV5w/gAGQ4aJCQaP90ihsio
Rt3FDb/cdySW+Z2oU4hGAB3Km+K8/2gbCBtY4RP3MCqu7x0AQi//Zi1nmKEGhF+rQiQbe9cqE0hM
GE8Lxya5lrA/XpgGkOgaIU/ohzOMuScrIvZYWqqfgwl1HtdQsT1ZlbQTjyZDYQDlm7XM2Gyp6zgZ
3DS5anJZikHfWXWXvlyYIDcmz5jVYs9UIRdDzmMWL+Lg6Q7oVfIhGpNF9gcrvt2wQH9OJA/7y6eH
jWd2HB08D8u4zN6aDuhNfbGqdUP8W34Chwt7i4cn7k6I+9AUlSSzDyQ5jbAfJLXhO+a2UUrbwAJq
wCLWhGdqzzMQo9naeldo8kHCwGqPBuNk6KJylcXY52z0LYGid9D068E4zYmayb3OvM66WUJSAJH1
8rMNFtL+nXwdQ15r+zmzAzZqfJwAC/NYW2oemvs9ZLUuo7WJxwNC13ubD+lutzo9ocV0GlShvXez
g8SI3AjIPubgItpKRZFW2NShp6uTVXUnMkaN9ipqrI4z/WVOPyskfsbWte4ZJXtpIF+f8Up21B6n
CnmuHUJykhoYPJrfA4J6X434nZM40q6y7RwGi+GRdJngC2vUcwTtovuOkK4rRNZkUMDz6YfoQ7wP
cXFY+3YElzwMePIjaHy0fsRP/1cNMErlKuI2rTWUyZdrQ5J6Oyx0t+gdEQ1Yk2MdPqFWJQujTta1
CeBPmNDzBJHY4Wta1w9raxQSsVw5hWchVp8sxXiD0FEL73qHHjDZbKKBx83eVYveBkvlDKQnPPXa
54S7VtRTaJAN2EB1dNByfp35l5idNuEmycNKkDa3nhJJ5ltl8DGiNRQ93n3t6lv+X9CK9T325yHX
36fA8yqNDsWN7DIpHI9lC/pcyks6aToACP+dhbFRdziP9PbP1D5BOj2gh1D3S5zVrG4l7/M1mjAr
8nM9LyndWLASLydjZ9YbhMc7H92nyDEwUVBVwqO8wG+hmvg/fGHS3Q74p/ghlLJX3+qApHA94Kwf
sX/NmoMzn08FjTpq4OrK9MeBQu2kfiPbT2lt/SSl1LoDTTFo0Mvq69B3vbMBSgQEhVyMfil5+dIn
YCduygi2TQ8NS2QvAPoQYgP98rDbakvrjml/wKTuT4fsSvUAZfaeBCMXvd8gdYGGJtvZrOyahOrQ
67S1qoEc39E8UuVSF8d6DCbVApR99Uu+mtpNQbpLAmaWwfROqxpZE5gy6QlcQU31ubfR1g1If8Th
liUaaLZxNWZxrXX8WyiKyea8+FcpM/sOZvDpRyokL8zG52OPz1IHl5InluP0KsATqK5vURcDtnId
X7XTpCZ2uDj+7vUuRJM7NXZdfyupGuT0hUvNff+1b5d4cgnvGFdguO0GGCVUztSXjZu//4SH+3Ro
jvFjz0vIJ39CtbGo3yqEsNBYdHwfWC+XxeEHbLsCyuM3n0uXTBiOFWK9f7pkXUwLGn3J/tNYexow
ViKEwXUaG8liMH+gWCWbLJ8+X+IERXtV2Q5Eu9eehxDZxOg/bHpowZiwvhzJxlXXEHZ2EOwN8I0i
fjVLwAmYIF+eGIw3D2mRm9r2De95rztFmsLvRR8R4WyLPWSDdFg72RvAHEvHAFAXC5v1S4CsKLhW
Duew68F4IAUpbTgmkNkfysZbJZ98z9yM/SOOixHdd3j7hRtJaU0U2S08449R5+F+uJg+ofSnCW46
XCQyery7AzhPGWCmyl/rfvBtJI/aw9MWUSwvXxMj+FJWIoseTVt8thweDgDmJ4G975IwF7SiO7qA
+pwyquR84cBpx9c8B17Iks9gGkLXlphxFBoeWRwvMVKFmTq+ct87Oe82lhmskqOdeb4sF7CVbHpO
tgTl5ayZuF8fmyp6EcZj4Ic5Hu6GvLpAmqBjmrHRDiIjpyTJLSBQEMyebOYZlhu2IA+mxNuNCc5o
hC8zgwehYprv4jmZlEoZ28AbHV52+LEpLil01PySHqJsHpjeAX2aiXAISiXNhxmEZcSPGf1RyPK/
hi8EKZd6ireE5CrIE8VC7h4dqcWV/52A12btWkjAf+1SyCMgRp4FhgQE8/AS0BwBK81e9OC7SHaO
BVbUglJAWVDbIJE4oZvnOSGJ/PupOEr2XMSHRb8CH3HjquyyxqkRGMz7oO7j8O/kJm+oM7q267no
j6GMxIoeJ0pIVbtsxutaCMiENwPieszCu4QITI5RkBcjvowuFZcjMdvgZWt/o8O308iXiExeEpii
ZP4CrwriZa8uqexw8ag+zqw7xo+Wk+LmafmE1i92HtMXWMd5MMKufcouA2mxEsHBgvk1/gSkmzto
J2437+zOg+N8D54PheACAcu3VRrAItPYnEhjkpEIjpAKnLcJwa+unn6OzCXl/cVabFmQ2T8pyIC0
zPk9IJFylYMk0hd4KnmXIMXG0sOVQ7Z5DIsSmrkNxePYPuhKick50K8lJDMntPpkcBkD+kBCprcc
eLBvCjF7gf2+Lg6RNhex6iUdap5ZLUpw2e2BfdRFO98gVMQksWyttpZyA/+mDIAQCsOxbKLTM15l
xhyix2Yoc59+dm3cxC3ip3L73ryCPDxZkRp5jKil2p6LV/kIo/A5aM2F5P0+24vTjsCZjpfAMpMv
zHYj1Xv9DJ+Gs3W3K/W/thtTJd6vc9c/c88wqAT3ExWIm1SjFOsuCV5BFHFuE4PTq/4T1xPIImVr
dCniatQm5D7I+NERg13O5DN3azmbzIq76tkdfghMRraX1lhCRFJxDfNQD38fY+N3H0T6X6aoXnBH
CDB0f7vTSuavQtPkQ9bjuTnSrb7ix8HoWCj5H3ldPx+Yby1Q6VhUTZR6Lgln+WOrxQxBXXuCaew4
wLjMck+oIrG4llZsSptmn5OWAwu5JOs6uxzO68T5CqiISHSN0dDJWMwv5sSv6avojU0yih/3VUmm
CYfluVmExF38S0Crmm2gzqnUAdnElU16R1ZB2kSUXg+qQu3hzyaSJ6rvns7Z1c7PrKrWoRctFcdb
vyRpv5ivgnBvS3TiL4eCv2CjZjM407DRcyyuBnbkS5SrakmZ6+0KYoxa0xhxpDo8TuZU98ZsQa6t
UqwLaNETtbVijac9KPk91uj8TpNbZ3oxKOlIScsqQGQ3gU0uXFNZkBFIZd4sjmIp9mUSi+7FXHEk
Ee4owZoxM+t1mivLu47qeuEp0Z9jDXVBoypDKJhDgZaY5wYKTxk0v9UklbCpogzt1gZrXguOJO5P
zrJ1LbfFw5gw8flGp3mTCCVsmWBTyEjuGMRc8w+y5IGxDDC9J9WYUvcPNT/VRffptPfWW4pYNnSe
zW+m8uyacgNUhV8nvIHMyEYtyN+mHp6sEgb6EXPA5IY53RqRheT4QmqiIMC1tkYKZX/IU/uilIlm
hykj1fSR7Y3rXP/eN9+NWY1mORFkitUv8CXq4fcG5vR1Ddsi5OF5GXSpKnexZknUKMANAz4GELgC
DyUdYkg3IQrOTB6JsRgX/qO4e8eEEQkA9uyMl4RmZmlbzFqPEUxVTsg/8z8HJ1MyjZZMw/uHPXUa
8tcUVmnMdm4Lww0dARj0oarOCDS6nYiT0kclc3UVjXe784Y6Id9L04JS2cRKFvEqnluHwxPQUAO/
BMFBpzVHDiLBOUVmrhq7quRIlXEE97qI0xymeg5llLaM0/xyv5nD495RSHitoXXW8l32jaaJH1lf
UqMyaFUOmIEmOLbxfKfILYyFf205sCs8O19VMksGvdJsAEZJKgoBQfEiVbQ8neJ0qD5P7kJkGAmF
a+KgODJoP224qfbNgKmVnA/GXFaOYOoD6xQROuOXMg0pLiZkh0h8gQYwG9u1aCMPPhmj+oDpIpv6
8MnQhp8lj82X1HZvC2JrjIVLFlJOpBKgfNH9nZQbHNOB5XOvmP84FeFK1h1neVnlQ1XJabESrXpR
/qnTrw18fXl6LcLFYf8vPtfSy9e+RYYay3QNO36k2XEPQm3kJWkxXFuDCqeufEdkj+ehbt2qSQiC
tju9KggGCGBYhuoVypsFy3/qc+HFGLfIhMItXlLrH0LTj13F4Yps/CclNQ4YVC253uIQiKKL09qx
IEDRjw2CqgGhV0cfHy2D1uUbDUV9AAhX0Mf7KK1a2M8nXaoD4wFLauCRZZe3E3bpTrfc2yFmazh/
0q8+RIN9y6Mi4oQke/TOlNLj+YlK4lxzm3vBoY2PKAgC7hujH9y761u9bmd9h+K/lf+2hgMjINOb
7f73dqDLvnglTm73Ito7HLK0npJX1pPgYEGNXAJjPy5Uv2cJWwcPj1PlYgXO3d/cKqtmnT3jXS8P
YEG4eqcb6AtsjtnsEmxysjBFgRGeJiEZGXp+s80zM6fgBDvPKzTZETCc8zWAf5woVOGaUTWvcrj5
pLcMvMrAzio3tm9Hpe6agvIkubWMCvmTCgBcWXr1wOueGo+rQhN92LPvIU6++KivpmK5Xd5IyKG8
+hw7H4E4FRl1OCtkhsr/yLA9THLcZd3j1cE65HqTTDT1JIrDx+8JvgfgUy1f8iJ3NY18QLhyR6qP
teeqcIMUHvdZKc5mVEU+ewTKby1xscrBhpM0DZeLHTbBYZHM7YZmVNhlIwilzxsCjBiGmz8XFl7K
W9a0aIhY4OQavzAaa6zRGk5PKgOriFxYL6sWwZMh/GlZ9AiXy0tL5772R/ueQb9YjpXJ0oC2ZrNd
9QKV2MNs1VZQgtVJeE8WzXGGtxkZk/TOKnma2jkbi31enjgP3pdkhAL0cwB/l1HdWxQ0pcqgpUtS
TfsGCtHNFJ53TY/dsgQwBpMMvVeM+Bka5C3UYijN84ESndHgIxAG90LXHJs9wtr/HHq3BGzGmbon
7uVwQ6wfotjm9n80CDpu10PPRe19Y+059ThlgGXcRXc2WH7XZBFDe5Ds/ugws9q1jiruuF9HEP7+
m9aPTP98Pnd+hJeYSRAuNQ1qQn1PrENWOEOKHCtMTJcJ1//0qEl2LsT8k0PvDze1GmPUEvpUUy+y
VmPP0EPF6s9RYHGENZFhHCouI0E5a5yhZxMwip4FerPx8WqeGq6lLH351MooJXPcCzzLS9B1pw5R
Z8dTVpRS5sTbTdwf1y5zwyd/ca38Mb35oMU+ydpajklNHRgRI8ONBlmbGbh4/A8R4Eo7gbLoVReL
QD1SunpBgax2bIORhKWnWsZ02IYF3gV7wmLotZEigJGT7u6pTDcoXX+OeoMRdHTiK7EoEu66FKa5
UJYJyOcYfi/BEhk9KbB8RabFvI/OCx0EZk+Unwol/I6G1REJyBXzri3ArIaBvl1z0Ul0iWG1S49Z
07Yjwv17CYxTmfxwDiTQloC4jjZtJnlLabxptbUreakPhp61ccZMHyx1tmrZ5s8ww0DNdhBGZhJU
lw1PGB3o3MLn6Q8g22HvFBpMwXxHW5nh1Q0td/p51T9+IRtodlQiEDGc7zwFSGqTTTEDphPSWqMA
U/u1BQgU6aIsh8b6GqfZZOIce/cDet8+cocNcoAZ4yO+oll7bcMipcxoOh1TOtQgeU401/+akno6
amsWun3cnDscaLcuFVrTtN19+Hy/gZCd2P/pe559ICbPBLbkrkom8B7dhHRs5TjTkDtl5L0hRVzY
HuRbQekZf2dU/tT1v6MyeMHtuCydY0HVbMOITrmWz+dXQhHwXHG3NqVDnax9NbhM5oNKkx4fzIUS
t0pGc/basxd+TqXuyUjr6j/UzPbpybJFp5DejaverTACvA7KRskpuUGSI/FIYdshoBMRCOz/K4qI
oGlQoe3yftFlo/PYPeMviyeanbQcL6iJW9Hg2GPPgeWPOK6gXXRiSRP+SB3kYwcA15pdvMuGnF8v
4N3Ad0Vdd4F/88PL2Z0yxyt90eJUkrfb5/Yzl8LFgkaH4BgRoJoG5x36tw+KU0RGU9YAC+YI3Kq3
T59In9E1jMPR3Syot2xMhQamkZo/X+Zl0F0Cw7cJk7rpChXNxym0cd32PcaYDJ8S/HymlenhSkko
GK3lawi90gnjcObQgSqKJ6Ucb9ZjG9InEMHZ27JxL/dtGCBWH6ZAkyKDNKcnY462Z/fZ8rwgP/1e
gmJKqFpDj7vBnRL29fDq3ti7bhtbPrWrL8sm9Va4reA0Eca1lpAAuZActm+u9n42tmCyuVAL+Bls
+wgNulhZIaM+PO41buoTRnvadx+ueyhuV20cUSun575GHs9TZU/adJgfSlog113oZbK4Cou+9LJo
eCnGpf2HHQtb+A9uVe9gQMmoqIrpH5Vk/WIEKFU+1EPLaBySRJ3b5Cl98VLuMyBWTqiaCb5WqM6R
4zz71QJ7nN1mTBttxZM9BGsjIXHjAydq0evNhTPCt5RFxxK3L5fMZsdJEA3/niZ5ErPlC5Pq1ziM
eS959vsU3X0hLvZ1/+66z8cTYp+dCTLMiyyKE/D8CZaLicLUZOnC0PdLaqxGm3fEJVWX9EvZwdqG
LEZI+/o+sB/Ti2pYNb/NMryEGhmN9bqYsbbeyJ8qFQneLubuGKgOJPLgCiGZgcsT50N95xQZp5Yi
d1+vvH6e368wCsdmQb76HH+1wA+MIgV9aBmrZkGN0PNjhl+2rTEj1WtS98EninkEidhrsnKVd9HI
xHrfToz+4Bs2hvYfbE+7albSe8L5ObqGtibe15rALKoDnoeJ2Og84rAlm2w1uBAjG2C+cRI5eY6L
ieO/p79749DE8S9iyMiMWtJe569XIA7JrSNypFSiDIBpDffgr1fhhmYCP3+lOG49TQ1mqlAwl5oM
Es4zuseT+zACF53zY4F8e4vQeF2TqB4JjDzJuZmXtyE2yzNZrbqL7YcLqABIMChJvbx1kBuEDbaB
CDHi4mecGStpXmLuTC2HVzLfDps/7GKyl0tQEo7XwH5v7wtP4UD3LXn/0bMLLYukKTZjmHaZfmKJ
YnYzciXyNgaKE4+1evMZcK+EV9LUim/QiEpcATfVdjs2JtFs1YJ7WFwRk9asEFMJP18jsrYx4cdx
rW0L4QE9VzoKzq6nnMRDPi2IADMQWxL+I/pTTAfpkg/prLn1BwbcZb/eUu2ZmY3+rvNqrrGrifoO
Iqc01YYwC9V4mHtNu7crHtc7fVDeTjFdwQ+0FCdhAy+zVlqKDOGhAtwVGzwNrsXHusVqGl280aQ+
PlJFWQwFEivvdG9v1zrQj4izl9HJkMfH9yw1RnlRvq34noSC0JEHg0B9ztYvxRnXZ0K616z7d8aR
QxWAe5uFFZH49AtYQNTfd0hCRpDxmFxYGt86fKvnrsmT66uqOdmslK6iV6RVpdc+CP48D/goTsZ5
7busrgoaHvQI7oeTNUftwyiZYV86beQGFYKRcTB+3zYS2zJ/wMPhv3XuEqXJtXbnk562j+USyVEe
vgDlpcZs8wOz5PM0eviK+tulAiFKVLonQCzR35tXCTKo+7Ivsc3DlJf1oBw3qb4hGsaUVbwmEn7f
Hfo+sB3zVJnqQUFxRoe5gI6FtD7HPnlxRNXkjsGqUA4QHHjixT2ClzHK/Vi/8DjqmZS9iNc/Rd0a
ZEXoxNggwn+O2Bh70Mgv2nOBERKgb32VS7I3/vdXWvUBxy7tiKYydW9xbpeMuXFNrqCLonhXJuI/
tibTViBwZyBEFQ7wNixE1iXs7a2zGh+te1Mmq2uCH0qGb8kLH1873wwUX1azzGTlSPiphd0BVhjE
2kM+wXbGmzp5ZSV1v318eTFCFNxxQsqHyg1Ey2ZajNvW1bve6TMm4L0MU1KuSfumXbs3I2P/SR+V
ve0Ckuj1LkFg6vZq1gNGtcAMFjZ+IR2KM0/qzJ1uVqjDSJUHJ1CqvQmSV8O2oV4EZy7w2NPVV/lN
/IGBUqik/VLxVZWxRZmAu7J+q456YZrt+jhLe7fcPm/i/nByrvOIZVtq1SX020AYk9fb/KiYM4h1
sToC+h412gPTA6qPrMgnF8CUyf2vEk71Tw/qBKwO5zIkU+T2hS9Hp6T2cUpSb7V4GhTRvkyrI6cg
DqBxoYKQvjbJ0kjEHixnrTGZLrIW28bVcaWs9w4PLWVbMfW4t9iq7j4WwZ5IE2QQDkcG6FaVIV7B
g7nUS+ERyB6QAWCm5xlHEjo1NO4pcWXrrnjPkaMEXqNqImXmCHj4Sri5Q3GCLHBhO7U0SKVuMsp2
1V+/5sj0nGVLP2ThZUFo1lNOFGtZSzXFLNOkBB18Luam5lh4OwbdqR8X59ZOywKw5VqdgDMRRGFZ
0rjqZs80yr2u6MJJOplO5kg86taRqcTu2h0Gu1LcL/OSn04wjG+kCuw040trZEpn8C0ulD9S1fDV
m85HnAnic7FuQ54jDC7i0YYiFiXbrO7jPNkkAJsUGRAqiKMP3Z12+pLqUUx4+yCkC1m2vEuiUkDy
8vkhIQYOgDetyLtkmXKi6geRDszA/6VGNYYlUtlk8q/VcqPDtJh6MCwcBlhWqG6jm5yyeveuXg3R
rsyWYoL4yHQ1Dz9FklCRLm3//Y/kQUlUhwYps7cUlPTOuLyPEvxyu5s6VAqBzR4utV5Hm4Z8qAJ9
L+IAf1fF2wb/xKf6AC66Gn8s+hArmHWvFWdsTdisRy3mlGowxSAe37bhGFvvlUtlFYNoq2m6Cc5s
ev9noEc35xwJyfQxqPLVO3EbWbvpfnYvZdrQ/WsmIKUJtaNZcv5gD6OkCbKAns2+R7DKnIth1MtL
Q/n75kirn2XsZ2OwOH7vcrjSvPdkc4Ggi0YPlgoCqi0ByPFEIA7kMhnPmcHo5D0idLDMqFS9yQbd
Sh95KWCD/wKq3N472l4H0zyF/mobO0nDW9Rzq0ioscTgqAyingvcxXoO36aSlL6Ad7eFdImbWlEE
knEi0d3HjDaMY6ewUs2YkJsdipoEqVfbnDvy8oRFe1DKPg9ZSCVa9t7ZHdSEwOga4YfjNu3+v5Pm
F3stJaKT0tDGvQloBuzdGGkHjk8m19N7mNf59wxt4GajFdlNzAEumt9jKugZZYgfquKJzgsEwPRh
CVElbpAP2DxCV4O6GHezLHnNBnuzDy1Q8cc6eCldDuARTZMxJruJPct5nA8zMJVOHpuRTwU9ZYKO
klQeg/a+NcvSfMyJbyxWJpQz6+KzWHUGAFIuIp9hfeXZhh3TcXXB7nv7a7SreyMXyY7AwzAjLRCl
uQxqzUoMKBd/VxNn7e3wrTY0YqgYb9+IvFxtn4Q8XLSyMhM8l2cE079eIVrT/mFMb9hktFbF3o8I
W+iDIu7bdQaKKPQWO6eM6eErb3KMN+S49CLEt9ox4Mkz2fVZAJUcsTf6G8cLIRWqTfieLDwSCoPA
SKP4dId3Pc9VGkvECi2mUti+xJjKEaCZtUwOjcBxv23fvTNKgQpCzf1/9XlUUQqJEVuNN7h8x0EA
2MKb/RPD9aEj5Rxk0zRSjLdZywErUFFJlPM2B7k+L+k2s9HYVCAnxOf5TtZrzpoTSi6o+q6yPNfC
s4rZu0cBNk1kBKNIkJVvk+QLuAtdTiUz8G57pc9mnWQvilOEH3+oPyuyAm1iFUu2PfwsinwVNn6n
KefwiKBnJTugNY2SXG+2uEiQGCyP9O0Dia7M4/p12CdZuZtNr2vy7FCGBkjalmLA9Ldfhbc6CBtf
2C2UePdJT1Py7kqJQmFRhll7rcd4BohF2oHG5bqBmdTtoJdOOJa69bHqADrS8TexrnBGxGVwK1li
OybJARoUB1F40zlIOK9bl3xlLDZ47clMpiR3Si5DcIn6fbG8yfPD7oPTqsexdMul3vAehCfHEut/
+UtLkohTw3kyg6/omtjRhaxsh+hSGgE9QmQjWC0WntF+r58zfjHhcCrDQSgMkddZwvzKcdyY8au+
r/HTjYZfYzJkTZC27qwNJGaHsdzM9cyUKV33lLlhBSHQCOHBVNVVz8dhMLm0fkxeah0IP6n2XVK8
6hFi36VT61n9t7huFrIE0D9ZPsMkjUoBL1w/TqLWfmW7dRWMNCe5gZq1PeFWDteYnJv4iFyYUl47
gaUwGktxAabbk9ur8pQLD46nseIuWnW9jGwfgLhEH3XUL7oK5n3wJLxW8LqZ8h17ltuZ31Xf704o
G12ZevWasxmP23MHK4TOnATuTswSUofQkUzKEeO9Mj1Vyq9a1wvgU7i/+mpPO226FkjWs9nwvbr7
SR+bhwQanbfEnUH0aL1K/EtRkBcy6Ri4GYamrGWl3DM8MhEF8Mp4H3fIL88tPqBQWoBHCl/j1nZ5
N56q5kFFA5FIqNG6SL3ykmsEuFNfOvyDv7tLHndHnHRyGVs1Ryqa4SzSmokmJ3fUgb6jqstPcm/f
R4wx231mmlGJNeFPMzrhBES7kYMGUdaX+exSw2Gro89TbqTIS6mU8UrnAhHEt3GFui2AOQZGHJTm
2O4FQPskgbe3AZ1gRZRh648mmpqRF518TtzRgg+JXdcrW7D7+uOP3XOf/meueBlOY/jQWXiCrKjd
FRKjr8noMkqMpTLrLigulWMstWyltcFIpPIzQFx49s9VhsH4ybsGPDYTwiYNRMt/jnwbKEeK5uRM
xcH3kVlgIbViukGEPouVlCoqItWG8TP+BSk/jtbrLbQzJnhEbEiac3WbqvF6gm3rXV40wD8/jORS
g2yQHvztGZJxp2bAMnzyPZN4RYKerUzIgfLq5rQ3uidyapPZXg+KlnhaqbeOARxb2eBYfFx0czny
9VN4wTpBJ6OHnPraJzEyTTexVGUdavu7rp/pOJHpWe2d28Cj04RX8IsPih4cTguqnHFcewAnPvs4
1qfUUjtQisWKP/dttvtP4TmkZ5xGFZkx1GgjhJNx/1UwCluxSzoCsyN0UKXFZ5uAvQtakpJjp/Gd
X4FJcdXg3KEt2l6n3fJE9ASyx2O+eJRimPIOQLaJQf1GPBEztIPv3EUcmojYMDJT5kZ6e//PU2M3
oZper/3OhQg1l9YZBA670jY8dr4pcX/g74hB5+x+B4LCKqkpd0Tfa9CTwjRAXybiArIbZ6GGoclq
6ICOgyfmRMaerhWzt2BW2Qv0c3qqAFacnaFrHRNfwklOUVHFBpAVY4WhG7MsjQocNS869ZkpgURu
RJ8s0zka7/IK8ZuKceeqqac1zlO2HYmowPoqIFKfYs20slLJyiIMa+T9jd5r2SlkPix2jGbGbfX4
hgnRWpMwL/ejRBCoQdagbAzEOzBSS8DP8CylX8yZ3OG7ejXYdopUWD0gLk4TA9BCLsNNnMZaAUgS
OV9yX92aOVYByb+bv39HHu9FdQI3xEPTpoRGpWIPhkZe96QW+wLwIuTEzT+LIbBsRb2kQPUgQFrE
k0rzKRJt9KMnZ0Yx61ZwQwznEWm3JwL5bdT0R9JO+jUphwm24WX+FpcQYOQla5Bqp6d6y8WzTfzv
XukTqvZL9NnhujxMgpWTjKzZAfVV8p7Mhr66HaYzYE7jWC8eCtytm1uWTnH8L/bwCC9VFxhuywII
8cxyVZGSEjMOkxa0wzUvl0PdUwI33GJFyJ3frNTkywM4Uad/SoT2UKdn0gUOZJlTfBxlkpiE2n3p
m7nNHvwffBZ83Flnx/tpIxglnswu6wSIh2P4UO4xzU8NP+MFoDERjkVxzFc/rxGWKb8jmuF5D87d
58TtwqxElEQK0IH7NT8RjJg4n1IJRKRofau2L2B9DAyVY1CMILXjXGYK+xAI3XkKjvZQDF8wXP69
Te8iYCyTeN10jHl0feKKdA4tODkY7yypFF3tFoTWDFyd/b7pL/Vb16T94VxKMgipcMtN5zdFTWss
2IIJrrqYodEpoe7mTcTIooYm32dsAZdHbcylk75RN2Q//L+pMO4/WgcM/TDmQekEv7apfmh9d0lF
shocK6KVwleKVmOewz5H4HXsVchtJ+HO0yzXajO2N6PlxBQRjalNoNsCXB0hWt77zL1hf52e7nE0
FXk5UGVXbepdvQpSXilw7fI/pcib1LXgFacVeGXBTy2Dh26xCCfxvRtSoj18QIhmL+pBrHYdMRAi
U3ZNUWXdDNEUpjBbXr1VN449Y1TNORS8tj7R5pgzzp78q8YnUviZZIyB5Z0MY17/xHoTNbIWRfLa
dOsKsjux9RrlAdThb4Z/jA9NYbvuSkORyyaGK04rsuTAzqID40enk75SlcnhfdVBSB30lLHbPnyj
tKD0C4o6fWo3z6o2YMnPS7Z5QKcJ3FEfUnpIA3N+eokNWwARB80lafL9LM5Hz3WvrsUR58DlD8uD
i5MrAGibYmRFkKVbPqdzcdPrn8gEnfeOUksSA6I3LU/Bc6EZX2NhVj4TxPGDE+PjkoeeF18Xd5hc
ikntDi+vZmoybgZVs8nfW7hiBcd8ujr2BMzINry+iObk1WM5+FivRtpe+vn3+r44ZqRu25LchHqK
pJjHoMOZJ6xa72JfGj3YiNESJP2c00KcL0l/lXZU1umhYsGsgYI5UyATTcuJsWPBlrDE+dv1I3XQ
/lDjNvLrMFRC2D36zPPAj2Bh1hjTqLDQJjQAF7HYqXi71ELc83EVPxocJCuVx0ENn3SO7T73VNiw
pFrmIt5M2JQ8SVaaMdPvVXY1IMkdZOeCSqXWDeUvgeWeXFwYY4Uos9Cf6yLh2ub/Jhhv8tKs6nDQ
Dpqv0817F1cWq1poHRp7dP29fpLMhTPUVdFuvZFmo4+Fpum25kSNV/VhkcIknbrW5oeW4HOku/ll
UH2tMUz89yaDiq40cqllljmbfntBSJM28xJlFAT9/W3RdFF87W5pWlgkDGmGFbi9nvNFMJREsV6+
Lmuiot2WGNsijeSaH2Xon6ZrPuJsZ7oVLRrAj0h3N9Qmb4xq3NwaA5NeA5NB2kCRt+h0+cRFYEQS
1DstO49TPAd1tz4Yty6FFf+xrdKwXhm6q2NF3fRoF0cAXhtte0AN7ofnj7yticX/vlpNRWqJDN1W
4sMvhlJ0z4Et/tbEsyE446PJUCMMY5FkWU98nt36uc51yPboi8NTlpx1JFQK6Ivcq1NXOHklJRu/
A3nZVOZqyti3CufXA/tPOXA9oBTknuWxfo6W7AV1y55gRbSlsCzUQy3VsvH7ZzXZiiJarx43HVTX
HSrW/v0aMIjuextjtOGfRUBBZjUwOIuIpIL65mScop1czk64D//d37H1f/QiZDr4tgc1WlrEYZNG
ldPPgq1DiqsqXWFYysIXfHENK/GulhdLrXKrfKmCOLe9cPsSiAkeETAmRq6x3Z2/1raVzQnm9RrB
GK1l8OITrNJrK6GB0AOMT+rmsU2xTf76fUNd4+8aOrzmOOZB2FOKpnQLIfs7NU+/rGuae7PxPgQ4
mzgAxdOwXuDlQHjtY+R2TAKi0Y1Wyl3w8S+gmCb39oZX3WFbBrV7mXqhytVutZZQUGI9EwQfoV6Q
BYHZk+k7/GJRJ3PXsYS/XZKL09hOUIV0pFGucfHT9MJI7w607y79bYaW+PYzSmcA0UEFU3DddGrL
3HcmfKmphSe4V61viF0hiK+0AEBPBw9uoTiktWE3sor7pghqeXkmMvUy3NVM77yF+TfTrLrkar7J
ATP+2SS/klftv+5TPXeP/00uS/X+9I+5apGsv278xRgeMrMS56OE8+8nqmOJ3XzFM6bCf4DtugPq
NefPChsS/dCa/YO2Dm10TpzMVa4E5/lXq4hWFo7yNAWKW5BW3Bn/4u6iBq6MZ558wfnOf14fMR3s
QHkRNSAyAgbmKfzehw2sFjyIiVgtw8ew0YpX6kbXuuulkIihVd7EmpFFjUZ2eviHZJbfK7sGpaPS
XmPclfe4AQTyBJD3b0XEw0sQrukwo0Y9dta1Fq5AhIdZBqM2kBHJXlWcO8TAdgaSqaKXgtvga+d+
hepRxOjWMNU2vc2R+IDpZ8r7niqHR4RPejnLUqncq6kyO54QUOr0m46e5Ilrtekp6PvwvA9205jz
60eXqkuRNatm+GgT0xEXStgOTPRilM+dPzEY+P1I5JrsUPvWHbUL5G2a7SCXBQDxH/V7YkE0HqKj
gGMJbNKgyf8Zy1o5ZmCIRNiVEjKAhRyoJTsT++bgzziDePkT4FmCneVMtwUu11NGiBN+YsSPNhiy
jzSwvSc2agWgL6gTpml6OzMMxHtk2IN3Wqq6EsvsBtW6c7Fmwy44bJLT1p+65LYd2bUImkFnFwPq
EM4Ififb3BnOda25jC2W5FjKzY2H/LeI0+PjR8Vkuj0wHT+0pVlDSnok4EbDfEerPVGWVjTbDEEn
mRcyg3AR6OCWCi1Gkl5hr42yghUjlfOg5mRmZmSfAEOfj8XBhjHTYBirccNruWu5NoMXCj4AvT50
XfucJ2BXmYLMUvv7Djhx/VIWEvhRynBtlN8sLBNVf21IC1LQ/F2ReQmKTgLtEasVpR2irSElFAPR
LYtC+ehKc/q3Mp3tTycmj4+QOH3ew0aRuOspWMQflAE6LpHEcD96qwW8jgm7H0++7tGF/CL4UQMM
IiMiS0pr6+mZGuOWuWGTkabSpPpy+bGDEQKHDUImpeVqhsrQ0w6WUbr2zoS+MnPVBS7eWznpA+dT
28ZmSefYKXUbl7N2pK5ngzB1ox5TjxFyKTC01ZJqqEnlolJ5Xr2C7NbSRMbdJGpJybBuKcRwKKls
Le9MhgQZRKGpQEv2fnfkRUXZpBbt3PujiKp7jlPmo9PJkNmeAKEoMtRs4koU8QmHAPY6JO0FzNxo
QKt0pI3xruzfhVXBqRAJUjENf+1vLLXt2y++gZTZ1+vOqjiuPszr2K9fIzuhu+3CBCPFLEIEOKVy
VK8cIN6aQ8B6AOGHRB6gnDYFv9p36SMCo+1HVNTrVFol/uvS8aQuRO93uD0LJ03PqwruMjz9MkvL
/vKPjWI3sCAEwj7Z7JpMIiRXo7IXlhoqB9kDnjeSYN+Bb2izl5vQucWH1BAaFdmkqPEIjnZASdT8
yB370odZfCvR4FbaJ1H1YBwuHRfN+KugbvX5eBFiONH23+/9zIMOzXzi8iJCLFneLx1l30OYRlmd
h/f5PmTJ4+wKZhY9+KmO/h5Ko+6bFWIFFefGR+TUb6kRrzfdwRz2sLLlKct/WGh3NV769cpMYdoi
8sksI19WU59IYn07Q3HyaiS5TufwCC4C9my5FMkXmcxJgJZFs1+m6PiyFi+XZAfXryw0FVOc1VB4
ttFXLSfoxOzzy483VoCsJZqy+8Ce0lg7KYJyf2/ev3tIcyj8VKrxTfqTvZDoFVoEJ5ML1b1fbquo
1m5oqZ1gE+JRtg589Xe+lpglbBuyll/VJoPYxBV6MMYa6MhdNbTYeRV3Kc57lmXdPWJHRYxLuvjg
hXVlBYZhL10O3Udlsn5k8anlZr1LEN4oj8cyKEb9Mk2w1t7R2Z6XVDMPdsC7YnQ6U60AQSnIoORE
5mXkE82AeWAzflm+DrHmYLpaKBlG+7bobSNGkbyhI2RUzOmpEQpIXv6GB5Jk1eCJ8yhJrWhmiGsX
qLAxUAiFoku1B0JTg8ukFNyT6vMKj56cRHtnYi8vWrI9/rdWH5hK7ha5Hhvcgl3twwPBnrwWLrjA
neDVlhnj9fHqkHSiLem40QHClTOk35bwV6dz8XvU0OXDRIIoBBZla2kGuQPeyOZRV5mLCfzJQ2pW
8MyMiBW/hHqq0v4iD7aZSbm3jTStVhUtTvakI0rty4R7z28usaAcANoSlaCV468kFluxwizbHBfW
BJiN7bO3X1Tlqu8fRTMHFORtgWgfZyyZbH0ZedXw8AofcA4857cIajO5pcOjAGkocjJiNetskkKm
xf156HbcFbKwyBdVrAyqLNxH4dxd+pe1RmcqziRjYfJ6b7mMQSqBztVAaHwNywWmng9i0zTji7iu
jr2JNAfE6eTw+NBXTIY8ik1aX3VsD0KPXeYAaawpw0dMeGgH9fYl1JbVj4I3a7Bm2X3VQ5om2Fu+
Gy/2z6CVftEMUju9aBmO75Hlb1x30/1KeS20OqhQCelWjO2Qyf8eUo0iD5+uUSgwqbNUAflB/e6z
9YkzhwNhEjs89356nbyO5XEPyFN7bOWwJM+v0SXAck9gc9yLBKq4WxJ2C3/sTFnmAqlTWVxhsE6n
z4XHzjO+ow3dDyvaMsOA+ekLyvgB+VAq0oMVFamfEIQlfZSJ0zdWr/vyfVeM4CvAWhtYz0pT1nWN
7rpG4kBWKHGMAjniiXm81mSj/m7T2HHWHa2lvrQCdnBkIuUHrJI6xP3I46anM6y2PvflZDxsYMGG
2wVyd3Reh0d/H74Xsvl6b/i1tj+nn7wv4CwjwVvOyCv1PJj3Mi6WlTQb5M6hx/C0wyWfRCVcln3F
3kCkbmsghbOjjHuIdluW4T+PWh4gcqR6v7rtmGb/Lq8ToMpFcVbGG5N9I2OFZH0KZFi6ap2LKweA
XEK6L59WdxdzzqJfU/wXJyuhu2lYqtBxpqBGPKMA2a/ofDV96E6UGaEkhvX3tUII97EoFLCYJ4ii
fjhox7GMmFejJE32XOSFlbQHE2N9yx0Ug2nTOwUsgwqQg267scJZ5Z+hbEUoAWQMwGSU3e0TaXCq
0v7SnNoSgBllhZ0whB2jirqY1/8k2c2IPhm5Wrpt+6LFr8M2rpX4nA2GGXGxlmO9Kkwxy/cYuNf3
P+0cihTJHsT+NXb/QLJ+LZLi8h0yRsT/KG/IG+DdYmOQzFZm+E7ct7bcsWq43E8mFvlNZOf+0wyN
DvxLptvbybmRJOt7Ldi+jRYbIoyAJoIDvuSaQo8OtcIQktq4vC3RfrYdJJgY5TPN9chqXG3le08o
iTJCBdIJn3d0FbnLZ6Uo7r6tJ3v2Mb+bEDnQpIs+S/Lt17phsp7Up1qZhzpacwURcWT4HIeJXNCj
AobhgYr8yL741Qx5FdXibsNHurAAIWXCwXhloJftIaNluZJqjY0XwEt2QBpR2HW61s2WCUu/tXrd
F2aqEjRTARLv0lrj5BNtog78wOhibGFjYWQ0hiY0YVGOVE7lJISOxxauEOZtTCAtR5+CfZVIQLjH
+qHmxZrrBCI+S/1uP0CNZph73yiHlRVEX5DIUyM/2/p1p40Qq9WqqHbtuHLvib13B65FhfiYzfFf
7ZtYYw9JAvPaKSYU6cGw06a5yS1IWPUWRBP0ZPFx+Mmy58PJeVc5eMFPijnPbK5uB9ySHkGOdpIW
2yYRlR4Ri2NhPYFfDVmknRp29dV+EREw+D6+G32gdGUigQHqt/vnV1LvI3wcErUXgrDatmG0/821
Dhl1zhloGfUeldhIdNvUcwu4OVNbqvZHJpWdLO1Nn2eIGRIJD0odsPssztFOb63gquiPb8Tq/Epo
etYwfYxtN7ThPxt9BeJQjLHVngIkqEIqLrNkNfYXPVSOkfpuUuTU9TTq4zkmQOwA06lOpZn3L7NS
gga+JhjT4WeMRU6UVThb5lA52hgnJtNsbjFdblHlM4X1aJEn2pnjHzLMk5Q+NXqU6vPJ1NxP8h+9
Y3cmMuUbrjiOJkYDXzKWVJ5XvrqWkLs9gHm7ISMUlCxv5eibVu5Bk1B4FQq/dVGL83r27TyvSPrL
V36xyh0kKpPl1RRSj4z/4CGgQ2o7tcbng93mymrldMDlxmhRQp4/M1xlzEoqLryHn0Oiw0vzwMb3
i85+pKyF4b1DT75PRz3hcF2WwFH6XqvH3P5NpeSWTOOfgz2i0+eQ+ABr8Co/WpGR+xWmrUWkjd8V
9T2Mn1xoDfwZ3TL5FIZr0rEpbWgs2R3ak1lq1+G2woM6SrVUOmLoTqvXhV6/DyhDa065323FwT76
2Q4O9gVmJ88iWBADn2Q7/pIpFtvpoOgVi5D1Vt/wVX2Uk0MUoRda+dPd4iFgTMmSbhMKefnwiHwY
8HmmGw0iHeiImgANO9DKRtkRJj71vQa49/qnUWYEAI6BTAkao4L8OiN/vVXgiyPP9Kk6zBdcLqGr
XxVMtZDhYhcEnx22YCE0ocgc+HJuYrv9pZNei0v346rmyzjI6k8VtOeeJPuBBPIabA73e9844zWa
Z32WNZ3aki2OhdNNkyUmXSmpRaqjbt7OXUpc3tWrI23O8OgSAK4qv4vQXDfGxmpg1kTRKQBxnqkt
BL3G1DslHQoRuJCYkbeBHZgyhpNHqMOJXKB89S1Bz9faIKLdVrj/glVK1coPFJ6ngLYkjGC2o+vd
b7PhUj2rPFqe/joDe3zdgU3A89WXBHiPSqufSDdb3TPH01oIBar9ZiTYAL+7YZm5V4cjbEGRjTLX
Jb3DNwE6V/SqQxhhqa2ZIxZywem+HTUEsYubmD/PCTyA3X+cvqdI59eCaqj1ZDvTg/q7QWkRbB2o
U4dKpFO89+09AR244Uveib8m57W2G5EWZ35hHC8c91s5z9WReaKF5qOfKiga0IenRfh0S/n9l7A1
aVYzkIUs5oVCN7teS5U+SLRDkOm9Od2D0uKngp2vxUGU1DGaSVbQ1ibtWCWxhpp8hyJAKpKb9FB1
C2U+vUQCQdJj9b+TaJq2dYBybglde9jHlCeWiI59yNcci1qMgd8lZsnxnbXFIiR3T3uFsUqyRylh
PXbtoxB6XJiyUnFncQ7v1zbxCb+JqpHFYjZXSJPsLO4BOcO7zS2fMb3exUXlVrnHolJRMhnBylO/
ka+ylEnBpWlMDQjbXN1arGZcPMAeu8r5fzl5qHaxZVVpbESvHi/pEzFVtFAoyGk9kaePGzSZdOlH
2amtr9qyUmKYKtnal/Tbw1mecMrML9XmKq2BwlYCKp8uv/m0tR5+Bm6qQ0KBzfluNV4O/DKmP8lq
vsUeAoH4cADn/EcO1npcA7V/2LaezXDOqrRi40/olPFoDAWm3Uic4nz0reuIMSRl3DslsKDayT3B
SXXZq/oRrSLDaK/w9kuKSs9batLxOzEnsM5y+wZbCQyzXV5tVXYx7+l7X0Y42xiGhzNNRFoMuNQV
V/5j8mjz7ZLnQMWUBidspzWFOFqGBU7uDsjteQcWq1AGCjeFB5uSTmpZpCRA6iRq9wrQdk0rZZ8j
vDWX8+2TVx0mKx945QNceKmF8Lf/ND9uwCZ0zWRDrEqgKncsWFibNIxv+//wmsqtFS7WHIHNDshJ
ROMeZk+uhmxz5NLzz/3FS5oCfhbRUBV+zLZ0URVUnore4CTOfFwU85OmhKbe18oOCIk0TY27A/ZY
d85zY4NapNi9Y93ReXH1+I0SqypAJ1EVTPkIowg57ze3pX27KoetkTOES83PV9Ausc5/9y1iyvm8
gWbqG8bY+Svd+2wi31C+Mjhzdhnkr4NoWZj96rsAOKQ0QBexhcvMaA7pxJMnKfwDfaJDc2l7z6hh
5sjF7EPqs7OlJzwZmmFdQcQRIKPZHdi/KzWw4GF67/6APXSvK+0K87uiLUZYhZkcsnyUOdGWf7SH
q6E77XsVoMclRzz92CsyltcLJn0GR8Rp54aCVTnZ/r0/6BM5lzell4nl8iYQ5qK06yECBTJGHTia
Tl5M5vIBA/l2+yWL6aZVlUbWh/bKtLGxzV8iMtssjnHVf+yYo5vFsjyY9wh4f7ew6fQ/oLN+Rg8+
ioXXXItBztZykC+HYI7Fu07tA84jZXg86Hw8EVDSRjg6pMeWw6zwA5q4q7dlZkE9etI0L3hu/Mjv
P2e+VbNBiuJvmAdS4PWnx1ywK8H9hdMog0tG+9ozWk7WXRVPPOF3QLCqfpqXAqhVeF5LVklWpaiq
lyGBd40x/3JyuUFlKqSiW3bFD1QtMm0p0uXRcX1l+HlBHw/qjiPAOqdJWgPlADyj89CeOvlAwcK/
R/xIR4/1UGpQjW/BkZzbTKkxP7cNRkHT3TOJP9WuwYCbwLrxYDeMVZox/G/G3t/GM55DPt9lkOpJ
iabmo6lRRXMdMNGQjUG7E5QhjtQQ6u+MO8ca5w5tAszNso90jyU6H+1uzd3Yp4F8DpWE9qXrWvQc
TVlcRDX7NQUkOXmL0WngkhXCSjNdnBVkGYKfigTNjGPSDcYHOVDg43hoYVOo6Hyd3FucrbtVk0ff
i6ZGvcHgvrl/2KNmSArdBLrHZF8u8pfij+zm47HtrbchERFUCm7/vkcNHmf5VA43y94sy1++16k/
HtPRNM6dhX5Vv6LUJl3LRvyKF6r3VtpYmWG3WxwMxLz2E8wmM0kPSMJdQ6BMsz1OpCQXczApjt4a
5/xcvq8OyBSKkP9uwjK8eOFT7HrLarARuC3QVfJPcMD5IhqcaPTvWCebA9KGGVDClfjWF/pn7SE3
uMcPK3fV2ho0xdkQjCNM0pwyLIVx9HyPY5+4+uAr/D93sllflb+cO7DYZaI7W+kHgYrKptFBvhIa
rGx6Uwgv33qZ2EHoAi5C42kY9E88Fk0BsSsjsjtnv6oH0z79tQsExcMG32W2VxCaaFhNjvCxTKyt
+JHKdCK6bojpS02P2/28OwfqhlKlmE16MAOuThG/cNlRYXDQ1ncy4oOsZ0hjuSQ7KCP2utVoqp5h
eLekChxB2ltPZELsdS58Qr+NsQpjuiyuap1ui6+4Rei2dMmvprzSk8P18l1Fbv06jh73V+C4ETul
U6fs928xnQBSM882q+34RpfkOdFUF7fgR5mM/7Vr/Hv70Qh3xZcygxKv2q9L7oXD7nUgrGcgsxbD
AQgOODgd1D+DrJqu0vjX+aHnr7CbV4/Pictp0D5jC0sx4HPnzLzCis8aL9KCoLZdWVltMWeK/hxW
a5z+YoURMTe6/RP7KN2qAdrF28pcZM065tZvUokxpPVxDKvTwy/fN6hflW/z8kl+vtCXn28do0x1
8q95E3W9sarH7axp1zEsvHmbLRs+3bEViELZHU5Vh4V1h+7Ri5tPJiOv6AqpE6QMBJf+gxUESDBf
fnbCZXd2himww7Tg6YyCWzyJTkTj8G1pPiUgQ/pTCY9LoQo1WC9AoxnbIeCOC3YulqlTlICH8of5
aVOpcRbyhd5EicCLtimxZaDsnJI6DWbGOw4yL0GyMvrEaXqSXL8+TnhW1B2wOlRzHdIxlvVZIn/T
R38eglDu0Is341zv1+tsCnQKjyhDtILRf37JYwhDVBi1Ffx+xXJ/GwfLlYwocDZwx+wYwgT9VBM7
7WO0A3Rg0ka+vA2Fkd7qEp0aYfWTACgh40xCLX6e5wVQUyVEhyzzjKu2iyYWDB/AFQGrPF7TCTzg
UNuxUiP4BcxnDbtX2RBXzhA75tVxNeB9JGfAVAnrmr33Y/Cpg4CimFi7/4QkvaVZllKxYc1aqHPs
D/dap/sFREM5JtxG/TC3xKZd3zezdvAEKxKAdgzszYslgAkSHGtiVFjnCQr7vdT7djwALpnwUlJm
T77yUWrEw0eoAIueMtkaA+GuWoy2GdSiOQS+wZ+KmNbo7UCu9UXnduhPajSjREE3HpoAX/mpsTIZ
1nzSkyI43hSGpbwvHIv3TbHdS5wO5lbnT9GXH3EdjJHKjdfMR+rehTN01N1g4Ghknf0GkZZ7OmlU
+v4KlKTEiAcfRio+lBWcKgMl2wVnGDqo8XtyuaKgAFOoZWNDG2FXyTbK2aQsYpnItJ6qhr30VJtr
O6EiyM0B4F3iGcEmpqIgLAa1kKIHXCaFzdP6XMnKgF3CxVW2WziqWaSNJMWRAfdo3z9En8csv2OH
VLG+2JzQkjQAy7rzHqxcsPBTQxsSe0AKW4GNjbkuhVmS8/4aMF+g4wfV3A5NLafA79dL3RjVWjHA
Od3zE49BLMFwAVOQBbJjejV7WknKFJWPsid18uUt4qca/B6eqoLZ71chptopTdQGqioqePSCdinv
bDZI9JZ81esH5elchhnxVgu33TXxus5LKcLLxK4dIcybMRtX2IauwaGsHrcILP9hdudT6wun2Sfe
JKINeFPU4l0kNs8Io1mO5Dk1sxnA73gNgclVJZ84E6eXX0iVA8UUpy7er0kqPP4gFqG3J+VaynYX
7MZChyDT+1Ce740mwRZTvrkY6p2b1QXgo7bLM9t+1LcmbSE5zCnVVcVlsQsYlAD/ZNux8v6NxQdc
NeWess+AdDahcdlA7RINOJ11YBjgxn0gdP56iCTtC+VFSJDbNnhH5s+lvgNu5sOoNxdTx3hAkj4Z
8ciTYps6c/FU258DqR7XTgH6gV1GRA1ndZWUDLDVpoFT3FVKcZCC/ms7aUnpPybUMNykyA6/FDgB
hER3TBKT7PrPxIqrywXo0sWCz511+EQLhW6g4J77ZX3NN40f0DZ8LiFmHbGspnaxb2TH+JIKU4SF
9ovzzj+0ZWgXqS56EUPxWpLmPC9OfmbVNufZgs8t/Rq3BmbFn4BG69/5X/tbXS5/qs1X9bg4HbPS
w13hlEKHFutsBSlFcVislw71HZPzqXp/fXgh4Kliq8ckjk+ISLLMLGlhzblm3L6BmllLzEYwqCe7
EKZ+6zP5r+GGLBpleCKvZvWHZAF+Wn4bmyo6p9sGuPWg8Y0y9KyU+icZNuNzETAl4lJd9Aon2xgs
J0zKgOp0Vt+QFc5veJFdO/m6RRz+aKAA2Ew4cEqc5XhUhHWDOrDhCXOHjX1i5sryukr1MVLfAICe
BglnRJh5scVeSmzLFZ8ASa+ikRQe7lVj2p+7eDVuzT4KFUwvHmsgiENdyr1LWlkG2SCk/zBxQaO5
NIX2Ngo+xaXItHKUG4xkPlPlOci0LbDMFQJtWXJ9jwLZE23gOA3TwaiWhVAFGgIL+QWtlXWv1i6f
Tl+vEfGNaSmdplcj+3Hlmpq7dYZIo5roWHwWp34OJsbJTP1YHMWmqo4ylwuH70Cw6JQO+PNl/BJd
xvBy9CEQw9bgkFekSg0/yHny0Cj6wm8PWNoPx7YCsp+dH4OMS3PUYSs24sx48J1pXhRCRPQlykpF
HmuwWRSXCkFlLPeRIa+WxDZqSf6mkQPgNJVRvW7L03011eofoZGBh5A3wPz35MKpoS3BvquYekLU
MFvVz++bB0KZQ7iXDGQE0oQ5JF+VQZMV8n95yAnOiRqrCHhdrrMS7wUA3ckUIuIsUImGfbss9QlP
BXKPrNELHEzBmQo9jq2xSq2ukqsubVtMZNsJrkgaGUQ+LveLZflVygX80xULOFWyWNPmnGBYxXsC
p8RunvUs3NrV+jKr27WFDt7qY6T1+fgAORI9K95Ab3gU/lEYBRAGyOSi86gYJj8VmPp6z9Kdapak
gxSRWegql3sYENjVwCatZNnvu2LIUfzozUsEmgUY6gnM6uEtrClskopVPDz88vLQ579hX9qHaen1
PZ5pIgB7WBzXXMegFg/2jsIxe1gxDnKR/GxRnxBLw+lo+7GP2oo+G7/YS+ZkFLl5bwh+eiR22xhb
jJLd1KL/b25Gn5J4uxsGGGnrqtg4Na9RHQSv0VIKjWQ0s0EOklkKbOZOEQ+4dtvoOzUZnRkjDHrA
DFbCOnhGUfF3taLgZZpQD+zBAH0QQzkFQw16Qmew5Kk+P8e0ZSyMOK24sA3/0rwUvkO0TJalJnM9
nM24o06BqdAzoQkGEQAGU6hwIhMYlciqa+BSPlxd6Gy6+Z4g5vIWVwE749q2YrLHDZIbM1R9o2ZC
ePZpYM3Po+9gVjWG8hOOYYCqXYbsqOEESliZnFg2GFaEMVHKh2tqYBzYfJHzm+XReFIggZhqNy2F
xMGqMxKqMxEYVzLp0nbX630r3GZalqEA1G0zMqJc1m1WKjZnPi5ia+HMqGyhPAfRrGFmd7GkjJmm
g4BUop65YaN9S5cxOsMUm1VkC27XwZodQCHjrLAC7zvt3D9l15RkM1U0R/bYvjBd0vQoHruMNmaH
FtxBnshn7jhbyWUMD4BrvI12TsFI+jN4lsquIz1lGmS+X2bTQITEM4u7bZLLqf9bZzcc3ac99a0J
DwP8z6fCy+WkXpWs5eZlEIdcnJ07qsCQGYCj9TURGP4YrPOpA3o3i72rfWpugmsMCg82OgNcJUme
WVLwehWBkVa10RJLnZbmwktrcO675Lk1qkXrhMkHpZWyVso1+lJ+ApHdGr23VKzsZ02SgTqXRJFR
sB78BMf+tyznIrH5b9wz+eGl3S37MJU79Eab54A/W5p2EeyHpEHGv8cFLRQd4wCfHn4lJSnZT3b2
5kfvbX5msHcHDu1F9M0n8AViCHtiCscQM4meuLkmAOVxh3vBN97i19fU9pBnmituqyixBG2+ZsGY
aWj/F1XxUrpwaV1jPqtKsnrEgwwVx/32mSEoGtXuif941GqpWgsA+2h+oVlE/t0UpdGAeKmcJulU
wowtLGj8WdvIppczr8JZmI4luMjFwNGBu+r24fdC5+on1OkaDreUFUQIM5E/9nkykOVNhete8sw1
9o6SuCEmx6D55CIRyr0dxMDVbTlLvP/nPPAnkn4CesjlOx1LypiWwV6nNsxfNl3pKwLQbp7o+Smy
WL6CaxHcMjDhQ0KR66Moa+eQyuIorf7TXm7sXFNhtIwLLC0TX8AtW+2BC45I4gNnTbyRpls4IQqt
LWCjZDane5BnNcBpAQcU4GOHqMpSphBIPAyH2AF1JZp9TfzL10YjLkTfesf2nqbownH5boRpXq+o
3fFCjv13xG3ag2JBOc9dzkScWyOLAAKGEVbwkFwnOQb0jZzxBWP2sIT0rYEw0V0Gix5+f9O2KvzM
D6DRz7cS12CnJ8b2sJww4E+QfM6JtBMD3HNsxKSf027+C2DnXEduK4E0vQbgeJB6LtznhvyTOOc9
VSaTUyOufIr8JI19nNboRRtRwz0FC9EDDXIQei/uZ/LFr3HmQmAIxpf1kL1XYcokQreVeaPkS0IZ
Ei6wd09ZZb3rViyM4zmfzRg7Jt5oEomw0PXNuQcNsj5uROVnLFefzX7ZGwCi/NraaGJ16RSIhadr
0xaNonuGjNivedvdUYU/+Z63qDH0rgsAIUfQh+8IVNKR06QFJ4CFsXPK2b9JlXGEHoeYtnweWK9F
5fppB2UeCZq3AVG125LWxj4idsInv/ML48WuFQzniW+srMSfUdS87GU1b0wgWBBsRUifv4kUAtlS
8js+vwuwXHMyPnCUcHOHHQNEATWh1loX+8zL11ocFnM/xfWt3bfAmR6+ffXZnA93mJ+/RBrizkGx
tgFOwKnZYR+3reeuCzpjLbIE5VCQ0KQLQpOUGaqswUChV6ALwU38HhcOgbk9K3qqNiTXyDCt4dhL
IZd/yKDHux5BvXo68TJmtjdteA+qSGER7bO/u5q85MLbNi+zs9V2iefhxZFs/thvZRNmUMGEsyNW
sazS0JnwkzcnDFmVPyDY31xBkUUjLVvDDs3apLnU+Fna6MPFIkSkPXqpl7bQnYiYmc+/pYx7ivUr
UKBnKuzhncqH5xs+CJYMxvrIjLTEAMkse3klgDRU6twEyLBbIjaxyU4+3+iNjOyTA3KMxxyv7/Wx
drGiOQ3n8lFTg+zlmV0o9ck9LHxJhHDE2yzgbiqVz3cm9jTwJf2W4m/zLFkPVKx1I0UqkFts6E3m
sB3FpEv9QaJPwlHIvrL4rfgfR9CSzjIErDAGYoORngO91q5ot2XO7Wn7Bxj8IVNZQz7XQdh3M8wF
8fECFC6q/+gi8DN/MVmb9zive+B0aPnfj9ygQj6XNWBt4e+/DZaStwil4jLT7+qP7EoctSEbfQ7G
jAI099Raz9K+1g4py88B0sQp8NYe0q+mVc5tUiuUoWqu8yh9TF35wOQnVOGb8xXWx5lrqFeOiLYW
2VRCezUoi5GKdHDyUZLlB12dYhYxk0JeN3UK0hkLYtvYzsoQeN6M23d0D3UbaPG/r2kUFOgcNmXZ
BXTN3KSJ0Npr4chHUQWv3FsfpJ04oTDABR8qgjTHQkw/YHSLssGOsZC0ZFyrBnrF8+FbldKMYEJe
Y5EjiX10+B0T8muASX5//K/puWUpsXh25lASXdO8zXq3wfq7pt3jinHJZIJbmQh4dbYkcd72yh7+
7VzuFHkWJSFfkJO+Ho6noSmo2ShQBcXT3wtMLmIt//zEuhwCur+KgnwbeQUGMp8EnbG3z5F1RQlI
ouHELkwmq3a7bXBNIh4OATrxEOS3lxVpTUHaL7krXuRHdGTRf4UtH/NuLUGTzfhGGZQtIThps0SC
raFpAE5K8QKte2hOOV5thn5pDVEokmTJZfGRVYuId6m+inf3WXQQD5GToVecCUXRdULYGUIfRYZY
TYeASNHGTjFjBdnRbZWKiC2Fr5BP6T+A7Ww5BC3EhBbZJPDh0lA77ESoBtlkKdN4BVCFJbot4PUQ
C2pouKLiJ4WNNNj0DKDmNolyrdE8G94fpeEmbQc/6JwBDdz7mElh8Uoktn+BuPSyko0yORUF/I+f
i8DGwHMcSk6thpkjaka/+4h+jl3rLTFNnQgU5C7pdx7IFeUT42blyt9n1WBdBmu/a7j96RqPBiKC
HOM7hwY4kFzXsX12CPXgnE7O0aJ41s097Lt7TcobL0vwcD6XxFPEHQReOSMsKPgQzsaprh8+iIIm
WZ42L+OiCM8hukTaTAT9ugx1nr1l7FvWruZ9F1XyTsNMRJ5ZBB5XXHv5hUFCp4v/UrFR+Lg+5DJG
sOOdlChoXlPEKKDumwAPHUHQirSjAbeWAUGWyKvVP6C8hFC/tov/AlHk6covT2NnGCEGNqtjHaOY
0BNw910YTfBY4kDMO76vxYsay2h1ag39GnrTG3xDD10zqpmAqlxJuMrAczvTRd/eQNyNahf5SUly
nP7D8P7x0iiDICj0mDrMj6avdoxtkF2o8cWDn/D/SoLceCGje1eUyQlLR/dW50loluz8WtxjMf9k
FOQO7a/yzyJ06AjcnxsCZ0qw6re0l9QXyhFSrlbWrf5XY3q7qhbErTncqytp9IbeBoZBwaLIt1kB
YFhYdudl38gndeDD4Pat3A3De+yCjL0zb62qXoRrbfluvSBkCBnimXLVZGzQXoQpCCUwE39ui4lM
Syx9JzkeSXmbocuLcERjcGQ6OUp1FUth1orhs3X6yZrFs4qqNQrFEwPiFF+0d0e/Sos9OACgN6yv
SHkL82DHQtUurBfnNCZh8ttXsQwu5vfvpFWBvwYRjrbQqXw2SD31qJQ1Y4XsvQYqEnbdCvVW+O9y
TBfTt4/I2sk6sVbSeq5N0OhcyCfH1PnEv+V/93sLMUYPBo92XiBX8r8C7hWzqdRqOnew+qGXMP5z
gZ1wKFq0z3TMUI5y46HSvi3RdbQOnTUFoWK7Fb0eqP7YWhgvTODXQCkJJpP62fAdiqjxZ77XU2xW
H3NT0e2hhBVg+WtusNUI0wgfiTq2Q/6DjC/c/Iot9K61spvOc25I2gFiEVuQZ1pc87uAu8mxx1Lb
J+z6TMlCjci8jotkKlhzatqPCydfNX/iM9SClY53h+7Ww2iEz9vH2Y+NUD8wi4ADOWtQz2pT12GY
9JXG5WoXfB1CE68C2/+hvOGB7kP43TzLau5gnuW2SiU8yv/cMx2xz8eKgHL78LvwUNchtPXl5cqW
f2LY1mX6BvPZrO6snb0xPQuK/LHHG9h6DS2mCJSC+7PQ3LyQk/3YaC99vEg/Pg0xtQ2dATOIodPQ
IWKbqtvPlfYHjDlELdYHNza+fPLQPbTvypWl+HV/ecdjNNJT/CMbyhM5Ky7VYNkdijgI1jUqPAHq
IXKIk2RT1BdG4e4iX8ZO1GWrU/pJCgyspaFWiIm8yEzU39yUMudHL7GIejVEiYYP2NkwqSvHe6ff
dsbSq/VngsesxKsmexZMidiOi+obP0FYpaF0NLZvIeik9qfbLIkHFOVu6Uwgl70fvaO7BC2/kUtC
eDGUOfizCsyngjBg/hWop5ixAkPHbigHuWR7I/SQ/Xyc1elRRHpwBSkQEev5KZYWB/1w2Yk/tE5Q
Rzn6+dO5wcmGnRC2HJUjPJ6bN6giKFYJTlEpjIftauq/Z12F1Cqmh1jb3/OBYDJYidOPJZQw7SI4
G/oZTe63C9apNzhf2KW1MmCUn9MrpVcA5x44Bg9nZUVcC0Diq+BA2lDI6+lQODU1PwtJTZgBNFzv
C8Ce1XP9zy5aERzo6XaEMja1KkNsyIcXyeBjrOY83dSsyz2J+Y2kpR7NHm46w4jh9+aJSmyWprEU
v6k/ZBWsNAe+1+MvP0thS4FJuxMmsDVFR3DgfOaFNsXG1kAqXj1us4bFxD0wdzCnG4TYLmZuxgxw
+930OjmJveSIKzlDNCW2Z4c5WXeTObHGGd3dGhePDdaWdUhZkU5tiJxHckmv85r8bqKITr5/x/Ex
NEDsQWMDXzDUTrqC3Em1yWYJ5zm1GRyeh3pFg+wtT5/yvfGK8QA9H3iJcwDxyTdVLmm9xZBzJLa5
PkusvrPq5tXFvZDWBY9w/iJNMn4IugP3HA1AxD3Vu58bXPZ3FPizqvjai5ch6C8TYgiprXmpYtnD
lCSIvjtexYf8q8kLDoGzewr+nItWdXNOPzApMpGmKgLpxjsuQPODEU5+1DmQ7YvUQopr/oz8EFue
Vc0S34T4QU/J3bferx811qS1dVaYAutihdepGfTnLiPwfVUKQNOuZXtuiZcee+zDtnQg2fhc4S+n
sR9b18ihmiwttETywwHzraio+i/TWQp/erFOUWqDI/dI/BilgexpMHHIn+Tfb7SllyYLzeFmSz9n
Twz3rkY/8e1ggkjAwR1dbwgQSudVY2hfsSgyr7vK4AWJOsWf5wEDgZ4OHYkv5hZAKl7hCM0/tyTL
igQ8WoVA4l2Xez4iZHMbSbej5wai/ZQaLooaaJGh++Pm5O4wbj8qmo255YTVVtatvC6b2h91fydY
ZLyf2jJnnPllBlXI/YJAVWIQpOZElQtodIjX2+CRKhuFVCHoC6Z6mT5j7yMwMDWl0v3HOc0ufGg0
9qBfHP5ZbWjamTCkMunYIa7hbbdZD0KHcbVeywBZcVaE4xYyvgIt60b1pXCrb2dOLQkaeE0vSyEO
Mt/ljlSBk3fsSVWuToaN3aWcEd742LOU0qr7+l+p6OKNWLAlidTrqG4pXi9EKvcyvmjafW8wd/qN
K7jYH+44y+H0qbIr+/iN4sAksmRQ2eC0yTeQgjAnZ0ZH7y9cMQWbVkPz+oAdLu6YT0x1lOo5/g41
+7C+r0k5WfjoCltxEgDR/F7m9y2hh007Cb3qVNtsA5kGf7qzWdHQM58fQQXLfpnwAIKHDVfWYJJ+
ByKOhxUcFMcv7qLAoNbfE5klD0Jgg+1v0CuX74urhfU1kUy5kCxFrt//aP6xjGzWKNtDTNrET9ea
fLWjPK/JomHwx7Muc2mRqM+nlTRXyd3W4rD4P649TmdNysqwf7FGJoP2IVHXL2rf1q7ycbHqrg6l
FGByQ4gu/lIQNnqiLP+A94vjqqTN/JOPvtWW1bsnwkbJqqBm/PGXe+WcqlzNywnom1V5I3KtKEtE
Vct15+bbDFPLbRLmHMLeCqedFjgkqlE/bDQHS2hpURfodR4T/Bc1Js17oXF6nPS9OGREs01WT5kd
Jav1oMeC3tjiYNzQNLU6Qg8YGJvHpLM6vIHQKqJFC/kuV216924mYnIXLoe7KeFJ3W8amxl0CA/w
nxwSOdCHbO1ulruno9TfzyMQ/YH4e3Jzq1rEDfcchOreboEV/xOW1BC+crxdNn8yj05ZbsIGZlSE
ES0auQUqYRioQ1sYx3xgyEDgOhCgs4Ua16lgBJIvbcyZXhivTYp2fJa0ifxkaQq7ERIFGeTCsTi3
ZRioR1MY16KoQUjgTFJD8WwxQrQgu58MsK25AsGZNeshDkCB/8hczGk1MJ8ohthaDdSfR/JhBD9L
m99vrEEhTL91ukLFopr4qQkkYzyuMymQGporko+5Ga1PQ6MjuvpqaFE8FJE2eHj7//6rlxzDoKzK
uJ7mGUZj8VlMAq+wvtVnU+aE2xremvRBtd6mO61UFEgnYPVCmiXLRDGogAeULVJJ15LcHltiK17s
fMcHYO5CprkvVD3TZ7Z7B/0CPaRpPlXnyI3JxHT7N0MCfKarDa/HuMa39WYPMjLrMhOe2DrCkF42
fTkQI9EzL2iNIVlGO9Cn6zqnsseNd5mk2j//4O0QDFwviaq28nKI9+VvUs71WaIyqZD3iajX5cjC
EvUZeZsO4zHykGa2nG2IUJJ2eQscmBgZ6R+zyLb2/Tk+oR5GIESZ/vm3tMpUZ+BzUlc1J+rqI6La
0bjiZhqOizZrQZCdEbi1rjrJdLigdkcEqw7/RTMIUidO8pG1Ura/opNYBUE1Yyy/k/ZAh2An5PVb
VXyg2IUvui0022l+4zQ3oOax1T13BeTHbtmdhPLNhZklY2qWl+WeK4SKvHDYcOjb+6Zw5A2kJDrB
K0+xyhLVYTSps2W83dcmrJs2r8GOhrJ1wGMmDX8xl2qB3SGhze1qfrbmZ14LowqwczqPP95REL8P
m/6xre2gyLZetwK9acCtT6ETowJx9LaChs2KFvjc0DXQ/d1g3cSZ0B18wGT6BJmKGS2sywfuGh+g
ldw50wYdEP6pFf9eZ/mZ2inO+WJtB6BM9ZC8pLKXI+eKF/yDOFZdKbDLQFU6ZcaWg88D7w3jjja6
D1A7erFRuQq+Cr3UH0Q/Df35/gd2ifXsxf6dIeFOY9fD6/MzId1ZRHdgCl2k8TnA5WuOqs946veL
RF8H+E5WYgnEGXDd3kFyDk7P20eCnVl6y2hi5cMwnbGuHvvh8R71rc8nk+RonMkDuMXZTZOivUEf
MEy0mxnRW7nVgWOWq6ewieopGIosS8nA5MIdw2lCAN7M2FC263RHjwC5RjRkeXfC7AfyhBwzdtY8
8v8+oDCvX2CajWdNoIR2Facv8+AYmRmlpzMYCHy6pC8OPr7154AGJhJgpcP6R4Kvbzt5bJT3CwT2
ocIwjVXTKOjb4EUXIt+D+S9kyDkKIDIbR/wBSjA41ggPzke5PnTToyB0NjqDaSCluOCSBdewi0lp
V7h8LvbaT4rvvJy4NShv5TNH4/3pRpdlUbxD5nzYCZriVx/4Tua9PZLe3MMSRBZv4jPoHS46+Z8B
zxAkj/SqKXa8JlXlOTR17/j//mwGxKj3wT5xyT+1vDQF1VJr+q1QbRSKAjcAaA5Neh3rffSHYFpN
Bd4gO3NpzLHLccnztu6aiEY0BMlhy/V52PCwNz2fAwzRo27TwdDa+FFI9R4YYJCLykDT+BUNO0RZ
IMWXWlUkza9FbcufAKzZ1fztahtG+8vSYdEtsQUeQ1Wa+hr+LI8lizcb2Nb5IVF2Qh7Li9/yaAQf
ninxujO2WvaHd450Q+qhasR5nl42MpIOGKhOaj3Q0Feep16nnOPUQ10N2O+vRM6MnqvfcuWUU6o/
GJyos0qCs6T9cVNdMrBCQ+b2+/NCHiJQ9WSxCNWJW1EqY92Z7W/j/+9fBIPE3uUyuub6u175bxEv
jBQWs+/OZyLsYoN5aThGCx157Q2KhHqNxv0cHw2280khcW6d8w64T8S7i3Fi2yNUJ/sv6/EBKB1T
CageaN9U7nmG1HDq6Ez7FmYNgMRjTRyRa+ooGaWJnv1ExF6yvTIxLWQ8tUay3AspgGNFe/aBNq0z
aTNo/3XrZImQmU0jF51jJtkJKItPyba5rNDf+AVVjbuXn4LcMVSpl7fx05t1zJ4hOW5IJNZA7yQj
fvfB1qlhypglnHt8IecnuJBqNcIa30wtwlqlc9Ux5EypzAzrHeg2+Fg6Wu704un6zVTC72H8VcYk
ynhmXZfu+bmFeEnTZYG041mkCHhVlvYweqd2RdAahMWcDOdzHxu1+GnXc3GQxatqbgr6/GHWzfTG
+AIGvZkxiBe40Ax8+AlEU5xOx8n4ssTIOyFMtp/QqO7WfimyktNL5GZ5KQrf/oFfaEEEzvMqFU6A
4VGSmrXpQ9ra9wS6l/nJI40JDJ/3JgyO4feqg+B6kBB5ZoWTEvo0gsJvD9ADr3GhcgaJICg8U+36
k61STbawLzpqb7PDxzf5EI6mNVx0t9JgMKbWMApoNGM2AeIYcVEbpwatUVrq5k2Z6BQM6J17Kjoz
zAKeRdDtSQ1gI/2q1wN5FgX/FT5DkrR8QI9+xR/BA5sLRt1IMp/wCf3bxsRS66uwVxYdBleHiho0
cu8HgD7D8TtNJbqHbvfC95Nzg89pTC9NulB05A23TweTb9eEPN0XooODYflsdsUQXgURihfDcjLq
L2uKWNhZgXRRebOoNdfSAjH+q0FNeADw5PY6jaev+ZW26OjbVIFjqfs/ISKZWB6xRfJzyhT3ptCd
c7Ara3oZkikcU1J4Qhcl1+59sduR51xDG4V+1P8i+e+ggDlgnz4LKot4HcRLkk7dCRX1ia+gofP4
cl78jZwFQASG6tcmReFYNC1EK78cuXtiI2P4h6DHLPV4uKvP0D4mxTqLEnrN0n6NkUkYnPv3qtYR
9Hfw5GIpKF0UgbhyacSmCFo9kUl6xRGVA4oaZpoUISodYlEcMVwmVjWHmnaj035Tntlc8Q0chOBt
iMu2fEOJHSZyQ295vWw3f60VuEG4pJOjJaSsE0rYEXudAvWRjDY9riCUwHQ0I+LrkoBpQ0/Ysco3
IKepnS2mHIjt8NCBMhnyEsik9inaaj58hPFS+/VSA/BUlMyWD0U8rptcUBmIaWTLwc69dxrRtGZN
fiJI+u+xev2YMQI25nb41TD7/aSYqkQcDjLJjLOodd8gbUDi31GoXOa54aJDK4YmRzPc5lMNCN2P
YWmVde44ksQ+4wWIxTmLkQ/JM0FuEuIwbihwgHgd0hBOjaGFlJQrfos/uFERlWhKuuU+L+HszXek
qXygiZJLWGSOyIQwpmwyUmpDhu/puiv6ayRkmLXxr+TQ4zNHxdsPq8FebCrsFS859Ni2Bc5i3MB5
jNLuUkGWLdLZoK2PGFT2RW2p/oDzcRC4YMEQbU4USKfXqeydwLzYuCJapN/ydBiLZxN3gNrOHgeA
VAwahGHo6Mjmpji03P4Cr6whsMkLR+fFOkzBia3uIn7CPbyFheu9q1JTQj+Oq6Lw1/5TFnepQNMH
yYX3vSKX7FwA5IfbBhH5R9shv/SoU+l7ve2+7jV9W0SUzYdyKDSn12amgWuLydUDWxhxz/DO93HL
LUDrguaV5c4H1GESZAJj1drfDDDiVHwkE+2i+BgV9wdMAynPBbrNu1rmSrPEAGZ944Tdsmxg+puK
nsp+U52Z8+9TyzOSV5G5aU7m6XpQegGUn62eeMKa8aYZYejDD1sYxaiMzJqwL1zqAPuzgMTUthvG
TzRMDqc9He57CFV1jBWXA2nH0bYjl1O7NZDRytTHMcDQpjiIZJg57BSX0Alg/4vXUvLR/XJWBEeq
N76sV+NNypS8NT1pD1e91R3G2ONrplH3+84S+Bw5onGLPA44lD1JRuAi1kjLKDHs+dbvfTwlB+xq
z3Wj0Q1eUk/lVZ1il2sQCdmvoAYDjAzeKQw+R0p5RvYN0KWuK90K4r5dz/1f9+bWElj8+NK/a9mb
fcYZYVc5DEZJv30r3CglDE5NQLKzhaQIY5SM/fCIAuARfRIk/nzXFqwztFqyVdbJflnaYWqv2Xsb
6M/6GHhC049TB6IOFJzJ4Y8IcIVd3KffGJc+zYuz4yPkNCpkSLSnT24X/tJPaJyeZPvuXjVF+fQO
LOR1HcMqpS5CPjrhhLgPnbclm21PYYX/s6fyswjRJYPd+OHbGCahyAN82oSf/gWJFIDFJT6OsA9g
p+9EPew6EpMUCz68lq+1Nlr4Y6f+23GGQR2VlMZti6hPD7inYr9aYr0yboAXA+Wu6zzTfPDm6r/d
dex+9/j+FTklLCRCKP592fPPS1rTbzHEJw2K9tdltMsBzkXRmBMY1uQvtla6+FD4/Y2BhsSC8BOc
ipJf49bGv9iNLIr9CI0R7Fmw8NPWXjMeS4WR1RHXLVylq15PmwUVvnFo1NHKqLP/UmvGbXjUgc49
bYLpNQ7miv2W2lna7v4ymlnN4FWSOfhL6HRx+ieEpYt6FDlHInJ60pyCZolSnHdvAhaKvGyIDuEA
r/UMMATOxoFCavK7ZXMRQ5thXA2EOjbDeNFpYhIcEayjTr9lhSEE7I+JMW68KAmJarq47WoXivvf
qBQ6pb9JFdhFu+3lk4SqUZA0isvZR6/yGveXxz+4o5LQp46+15I9q65rZBfJNsu4I+ryCXpqpaAt
TKMCDKoAskM08nYNF+HJ27BwI/FopNVzFth5C7P6VTPU5UOFZfgi5XvfTvMxklh5HgZKW4WZ3f82
738NfIHh65vjRyEPZE50Wv8nA3OTlp2WeYbB3f9yn769dLH5m8EnwAiD2r4OB9gwE0jVYIlzKlBp
Uis+pJyGZ+GgyIQkoZ91d6/ASZq8DxWhJ+OpVBtYjHcuHYXPi5BjXp4OZrI+LFphtt02CoQbh9gt
HhAHw6Sivaxi+yK72MZCpXjcQSt2WYeFvmSm4u4nwJDTcSt12jtalP3fDE40Ie6rPMM8c5f+fw5V
R+f6hP9obKbkrMn11fz36lJWGo9hRJp4r4B4oESTL9JWerpZwLobODeJSDUlk/CQvetaY6zZbNbf
XCsb4nnRONX+l9i1P6OjCSRNVSeXA5xSclQgIg/OqNZo9H3U86QflouR/UWCbDbwTGsVRVghLQvd
afpXWLAQTqtvExQ3QybbncS0lpbQt4w4TnY9Kx5gMjouU9lFd59BbMeLKAloWzyPRIPMKn4SsQZZ
h5wEi3+VY6nM3Q3PaXZ7jPabwAXZK4dQ3OnV2gwnFmr4ovoz3bQcS11YwMnAKlyURQ1ZllkrbDwg
T/6KyMRGbtVy1DSpuMcnx/NDQ5fatrsPGbyyVC2EetMy/fcxgH9VY0L6ll9LY+WWAOsQlR5nK5oc
TbsPp5amcLsMrDl12n/Zm2b0Dyd8PjWXWsmz4rQPYk75MdYNwom77pLszDWz+Stp8zym/BCOof15
9twhiFzcGIKvYmaQnlHA8hsFIoEBAm+QCnemCbKmluFQeRwU7xoLeFpUpdiTwCHy5MdGvl+UUg6b
f5PBrLraZK0C0U7Z8OCIqBGysr2cpEDr1ut8zhYb/SSGza1nUp4Ze/vC/EB+vBs/CnVMBMDamGE2
WcL4qr0RXaX3WPlFgsGioWvQ2oj/3uaMVITwqDUITLVRUPCfp7K/CodjxgsLnbUHVl7F669LRpnj
C5DvR1XQH9DuQ744Q/0Cv3CXX9Gya3amaGibXMUjULnR1uPVMoLnyLcKgxEOHKdLjALhagKHoaNF
g6czioYRRRfPnR5l1jN4K9FUcVYmoNm3H8uuJ9LycNCyjTWV99gYbI7lPrwnwLr37WsvYLOvk676
HCGnvaStjaugJ8leY7z7GBntXsZqqcOsj4+XBVHltKpnzPLnx2YfFHzQj428ozAoYAV/wA1Mo+HD
OPQZgbTuhTpgGuYZW//8Wtuzi63ovUcgj3mKAdoGBY2+e2UHSeE3w1eEciE24TnOE2qkFNV0uyy7
CdckMJcd20KqB7BkhLdhIDoMSG5Lc08vJq1WPkZsUaxB+V+joPTJlox5t9r9nLjBxxM6D1fRMuRq
msYBZytZRY9zv1AHgcGMeKKS9uQfR+AsrRnEKYaZ3wfplVEDNCBUJxuQmsCxt2xY+l/dFtZ8HXQH
Kf/x3wrMgimUdx46UV53JBX1TgaHMx2vJUkhoDOQUdzWbI47fDtlT7v5dZglEq7wIpaH4p9PxyO+
Cs3BYDMMqST1+ezKcgwQcFtl0wvfxsxLogVctlO1/uX768v82cF1YwnZlS2XiYSjraKcqbGNz9cQ
mYt0mluh6AwXPegcW332gdcl4+sjkQLlcq7xN5K2+duQhO9XZmkOjtSYa1oSCZ6CKjYMDcubrhjm
DugLt7ThmFy+zrflHvUyxSDVkkLBnaJ04EH1SAtAuguT3wc3tMj7ZoiljSpURzFQ0l7qFCHy3FWg
wYeW/Hz6ukeDMT9B3KRd6qSG89nhgvfE6qZDmgseTt5SEz12Ia/tguCv5Pf9X3UA0JlpGWJa3AOQ
PTMWx90GuR/NbRwdEN4mPcOadmxmVCGMzR1WP/hGwJkYAsCv9z0ljtUfi8vMeDxbkKVOLe+7LrrW
Fvlmrs6rLIBRjtdyA5SvSiUzpyNFP+SnEFLZ16ioYT026WjLMrCW3SLPvN/IVJclNKByGAXejgzM
qT5Tz6t1Gd9WPH/sHXu3IH9ErJ/dZViRWwXd6Zq+jyDD3PwpPwzCaryU/kw20dgRS1vgKYcBPszz
o/F2OPeoO5I92hLzALyAn514DbT/6aXdo/nlCH/IIP/vAe2H5xdvcDY5kQS/vbttn6dEtNulegNf
7oJmZmBNXoc0O+4hGND9Q1vJQX+exgzH2JJ/IK4dirD7cMK+CA4Dj1G0qHE8E6GaYs1j0xlJ/Pi7
6XSLhwzQ+AdEq+/C9LhGGo6YLpAg8hbYkOZNFNA5rXYRDm0tv3amNDPduuTJ8Rsqft+WGq5eTLqM
u31C7Tk9DJC8164ZYp4rMUZS2ZtGSXPztHKSwW/QADpyOGZXuU+/HKqe1nEe8tg9dFcy8ixK15M/
kymaOf87lAN4QNt2+52GRZwEAee8LoAsB+MUCx507Kp/gWFpKWosYxEpw2w+adNPJSEOgqjvIYn6
J6dcd5JwWkHHtarhfZWrZIiXXEIV1WXjy34W5z0QbgNR2gqFayjTWoSV3UIXYzB+3zTqRM0x0kfu
2LTAJ433v2Kfn7jZD8dMhW7pGT2cclI5AqEuIfiD5DqaYlsu7EzSYguSbQMtO0DL6il5Af4+IGQp
XHnttS4eLOL9sgD6hRXqUd1FVhKCT+A5KDwNG+HOJSaH4+2w+7qHWiOSTTJqsVh2OlQ+0S1nufSb
YF7cd74ShqTDnsb+Ff1WipBJybJNC4AIHoBSQOkJNB2ry+vM0Al9pxrewnFrDfImRsafwwWAmPlt
wJnjsoWqNTVJDoBKlepZUl5uM8FsmLSQ+vw/c0Al4ExSBvgNvX5xgYms/TPyCKzG/RUwdkqqbyi3
Mlt58NFFuZErqO9baMd0dVQhpmqM3MxbOWiNRWX+381Lvm5WKAYkRFCmUyZFSzGZ4dC89eBSMlJU
rqaQjepVd10zINBOqmKzw/GRwHekDir2rjyRkfAetU/jkmE8WE3ha/XLnPzFjDkkryWr/adshjgZ
9BgGyFMppXp0Uj6sEsgG1OXj5bA/wEqPtX4ewKeWut6f7gFbH8oUplLau2vOeapMjEs22KsvwV9z
EMMlOHeXag4euFcPdGxsQfwPcX+V5q3ker0klzOHsD5qn+kuyp07qZNVFkEOEcV1b2lKUd6X1LGc
0vKDq1KSfkstkv4QWJ2m0kqCV9rE+t57sHngzxNaXw36F+68WpoNRr8W0ixfJ2GBSqAGU/02ttld
uI75tJSCRUzO/ZQiY+P10CUw593mat0F1PGuujsOEk3eWppZ1tOX+VLbQa0KulyY4bvvQFS6iHdW
2OEwojwfhsvavvJQYbTK9HLrDEjcCukjrMzrNBaf1R2vP2zcLLQL0pMJRJmdjk/0UhMGkoUJ2L3W
X8Do7G2CCy6OReBZZEulpvDq+PePUO8No719p/G36l+kv86dTwJsk5Odrh73A6LsFa9/idWJBXmg
JT4JVftKKc/AJKCDTYs1UOf4Cd+GuEhsAraTBbteZjfZR9xM4A8dy1QN+uwrqelLAwv5iI8MUyk4
AdfzxtLKgmVqVS+AmNryubXBLwKzDxjhi2N7ZBk/8wWXb5dj6F/HnaI7pmFzWJjL3QMmIDRy+Pcp
Zy3e3t6Pbj5s9YXVkqOrwLUPsBtjoTmmjMbgqgNzhDgJRJTMus+rzdLku3iU8D3SIL6kX4qYNx1o
n5xoNWN7pgrjCQbZEgfMsJxGc6xjeNfzjsp4VNXz4raMi9oZtJ3cDDSyiZw5P9hSX1evZW+Ovpex
y4ESEIa1S5QtiLo3QjBVILINgxFTeNGn7JwCJ55tO4NTmyCuHKSv+NvSgtL/07snlrqVfOajcBJi
97sewQuvtJ6SCDjQBUN+ytLb224Qsc9hZgQUAmIgyYJ6Hp2S7SkVR2I+pbwm/DO9FZEy6XVI62Ea
VD8hcKXcsytIhz1DGB10rAagLqBlWOPzW6SZDfz525gv99QFuO4yMIaPq1lVGb4F4ed3vPPRZ1tS
Yo/aM96BqCuTz1p0ZRLHYkz7xDGcPO7oIcJvTuQ+lfkLBlS+02Q1GnyZeCc96I6ZsGdGqvIvFMHm
HOshXFmlwjwShOSEgWABQFXN3CeU+Pyrwu4wjrJY8zsU3ITSb77Vz7SC/5MeNCFLTxu2nC8FuK8O
h5caLpJvdCJb8LNTmSBp46G1Rezjxgyroqtlf+qEqQnCGy14FBh1QjHkQXYLO7h9YGr55xc4s0d2
kZMnb+nZelabOJV0X8PWfowvC/ywCYjoLmKqlZ9jMVg/gXHTLHIewsKDgq0QvPUqwuB52h/OZ8Pz
PkGad+1QWLjkB/rnEcrRxYNz8aVn7LX6nTLrHlvpF/1eTGPsN5mM/wBY/4CjthLTs1b26YsygAg7
aGtkzDkIX9z+DkkOJduMpzp1/xESEtgdZTVF/z62gC/Oe/Bl+iYOibWVjzfpm6Vd33FeEP4zIvbw
wJU9VZDcKpPaG3KvKRKErhBzXbocgaPTpQvm/hvi3W7a2g0fGzQJULyujyhRPg17yzOsDM8ic8Wd
jPbeirjDjSWPstrGAbEhlETGc9iklHeKByrm2wuDn0MA5oHgpDJ+d3rcLSHJ7qoyhg5FTn0Wa1XS
eZ5fCCMg+Z6LAFapbNzvadIF9vMgyrkhCfIgnidb9gy+pRtLftYZYjMV90zmd2NsYFEaN6QasutE
0nzRWAkfJiG3OZTN8pvKc/63FrQbHIQyph+veysn5IwE2nXEe7qUKPhUpei+WVy1zgVbkAwkh71+
/X1jSlPMGg++zW9iprYbv6vdT4VZhgYXLGBR0VKLj7N3HazNj3XPM0BFflkediP2Kf1M9LSeuft3
vW+r4PzLK9FjqFrkmPcts/XOsiof3B1+kLMtgHIqyu6b/4VTYJOTM9r5nkRxe7GPlI4w8hmEwwiO
h9Jo5+a1RGvgGqeC8uyfJuOq29lHjiMortqINK2qyh7gRwI3bKmKQh5+D/CIQ68jBhEOOtWWpPvC
0sh09ei1woD/EkyB+9m7MqX3zpQXazglvAhiecD8aGX8dWhTGlmrHBOdSqaMiKx2EfER918MUmOr
N8uPAylgbRwddVr/i4rvFDDR5zV02jTNR/fs1W5yZNm/F4uJ+8Bd6iBhdGiMeJ0FZG8tQVtHA5XO
1URAJ1r4W0iAdnjETYI8x+O0vPVYsfyELL9RTUVkBE6LC4op7FuQrd0ldZvYoh33vdK4+dvq9hZM
mN2G4jRRaURWfDNA20x3mRVOo9GsRT+Uhu0fcmElLClC39rZ+8eFMyZ/RIC7aWQnnfcj2P3CAsqJ
JcNnuQU4bEfoFzKMsEX6W0icY+jMAX5e5MNQrNl1umR+DVv8k2ZO5VHDxgib71o6b1pbzGVSKVYJ
dQ9EOPqJTnrtKD0sHptoRZ7uc0rqPPJdRfvQUCm/q6RnFu782VbrOTMimhi5ricnITPjTZ6DnEIL
oA8PYekw4uNuld2UMG/mQ0VHA2uvQauMFZ1xygEf47ChxsTGHa4g2WkgCfkLnO+MlZy/MO1MIKHx
TFsAmrxNKTyqYm15hEHwTMTFdZsmBWnT4hF4GkhlxMb95Yx3ptknE7wzcwdCYD+ZrtlCpRU0whdm
c9NifmJRFZNbzuehoy6E8xZtdffpliCE5nqOLubt4ctlSD3e7LcumD8NKdy/kr4dI8D2MFwpqoTi
ngR8ILU3hpZuhnjWAwz1XAZuDrjor+sOfewAG6N5ZqhlMwpq0kmKcQIG7wbrVHNdg4e7KoMHl2jG
hX9VCpxn4ufNqPGXlhzmElKR7REsLttJW197GukyOmEig2t0RwsI28KHB/6hk5RTt17hsPmP1ktT
Wnm3zfOJ+kVNqc9Iw2R+DkST24PVyfvenW6rJTzUfRMklDihkXOy/PBBoPkRYIJmbO9uVKMG3l0+
fGsZVJDlwVSzNYe2cSp9e9gecQhQgRzQpDBWxS1cUvgZ7D5zGeEXDg9ezf33b0GvX3QNB0ARZ3M/
hONYZGuv5kCmYT9mXHVT5VbzwMZQJdlxCK89YafyM+IHERnhvn0pfm4LEj7Yef3slwXFiPB8b44u
5Z4Dl109aZjn6+M7b5Ic77k3ojzHfwrz5Nd8VMACsEVe2g73Sl1OvHX45dAVCXSWlCHi8m86NqXt
+vzLa0GFFZXMn+POU5pudktRq8pOwC6R1X9u14rAd+pJ926cY6XdmzMR+oApPJsY+UdUAHLxMw5s
kdLktJOXxDQztU7G482YGfe5LLwp5eAlh44zPS+oeEKcuTxWKgpz3rIu/T1hDn/KXOZK/bq0Eryb
wpSbDDjDDQWm3lXPse/i9kG5+RLe4n1I1BzkM77MkU+QZRpRsM0wN1n06kQiftadF39q/pH1VYly
wh2xPx1+dedozl1r0bcPqD2v6hLaby8+yrP/gDJtlz8llmbEUk/K5xmsh4pQFkqfkZb/qUgeC3at
uIrhneb7R+sItiNMGrFtdbak4xOi1xKRL9u9g5VAn6SiTatfEopQNYUeZhz2Gq1KIfMbmZVrGpD9
rNnthLMu1H4Sb890CfNTvboZLcJWColIB/vj2Id7/TRDCbIhhTF25oZW6TzF5B/BNgs4GC26fqHs
Nwqeb+okpSPoTxjAo1vBeMTckvgMlyqaiORPI5Bm1sam1dsW7YQ1l3gBmdxg/8ZQt8PSu61N2+MU
HMoGvltOHa8+wa+yXMpJmpFQ64YpO0n+klIAKE4l3Lo27h/XvrRoJw3HNTmfB4f6QKGpFhatAOMk
uy0r1nFesFogp0TzHIZIo/3GrwmodH0oD58RlpBbsjYzw/zkU4N7x5JyI+ezSnSrrhULJE03NNka
Hw0l5X7S1pxBcyiHpYmz4UAPBCdK597oi6sTQb58JdwrcNo2sY5q5VbpfM9bFHamiL7RqVI58+Vc
gi2XPcebKIcM9F92fNP63tA12BHXh5TZoGHM3o6JGaIzofZUxPUQCbPjFpVR0ORLpuAYZuNIxMlW
L4VMOqxHG2DSjPd/hr0j0L5d/E+knZWZBBsYv4qp8z6NJfStzQvyobX4NpakWqH6LkwcngD25dQ9
+JIdHhhXgdvQvQdNv4dfKF/LYx6GzDPBXNpzH5ApdihE/9V63qZ35FFkk/xJjsLkdd/NrxqIvHhY
UmwC0hNJ0WflPjBHAM0cOqowLLde1jI20ReUaPy1wZFVADiGJlKbO3fub+b5wcolGVL93QcajChM
2/YAgYX6KHqPnO3cgr8QK3JTosYdzmR942KEmF537ym7AEVh1DzG572Iv9ntNPTVowAKoGvofVkp
ScJlDE8obFP1RTelemVq/WkBMlRXEkOaXNXQPGqX/Ym0vz6imS1VYCOVRdrSOpjGOZtdSarNWeDG
izFJbbker1fhQeNiTpD0gidQ0od5N9rYSjU/Fn1Zmm28NwEEh3DiM28vqs65r3FOSXmI0zUYUsWn
05e6asbeoTY6JtXpDtF9R2swEWghPT7TezzPJxXYKhHptwc13QdNf7JVWJKo6weyc7Gg9nSurfjC
1onSvdSLtBgU85xUV0pMrEux4gbztGHbQT1WgykWdXtILIPfFyI1b7zvTQ2eooy9EHaxnYH/x0ur
b55/nIEwISrm4G5gvN45doUMVW0juMmuPD/vvAE38m9mhjqPLGsaQVxZ4kPzivUP5Do/660UqUle
3NP3jtE9DD77DfCJlNhwGKkKR/PyIVXCsQhBC6TqBJblw23KuikLGl+I7FqhUH2Y4AMwaOcWLTTd
QBINU/mDGiYI5T/JXSaHiNDrsYgxgbugnMvhnRYwyaRlH0e6fDlfBasn0cCbgH7lD7A0Ys3vq8l/
OU23rrPQGuQ8O2X4X2MIhjDa+SWaTMEmqN7lH6cvLWj+VBEVnvppaSijtBIX1l3Reit93PAGPoee
E/Jx0FUCJKSCsal7RL2pcXQ0hpr5ZG3fLh7QdQE9003+cCWZq533eHxSM+8aRV83WUEFV8ZHUwan
Qe02pRP7rv66avkVzwj2+mRlIsbGzTsV/cPq5z0+8Tf3AZDWi0NocFQXFFzEckLRDelgVU1fxllI
iYGhxpvzOcEJ5tkI3Fd882Ojkdl996PvnnkVLno4rgmxfQRdHn0Vc+AMzor+U6LIKFOz7tSi1z9+
5Nr3uUECnuAAcj23y+wnlKvW5rUO4/pajQ5CSmtT3+8hlJNAyVRRyt3J5oyytSEIhWBRWjGwqrTz
XwT0Ar30rWKGPFjNN/Mt0kWMWR86L8qDiJmfnXi9jVsxsq3x87A8u5C6dR3wAssoOhH2tTV5BOpO
qVB5WzfNfjsS3kfjYeVhC+8inKh7Nz3Z2/5HLiExVmHwrMwTZixIlQJkQUSU16mdpx5hA7eHa6lf
+Cc13pC2tkiuYb02ad3LFVBaVqvB7B/suHwPAbnnbg9ZqVcEt+Xu5cjHVFTFtjTvJigKiGORz/Vz
1uzKwx7kPCA/DVJ9D7xyxx4LdIYbHGJXO4EXHKtZ/BpV7vgmqAJOBQOTVubyza0l08Ck1NVgQ3wv
6pgeqst2xz9c5suhj+YGmfA4OyeynGij6s/iYvXR6C5wOpkWxSPB2JQdtuT5cYJlbKxFBy88LKRn
m4h0nKy576+4GKfXuEQT/y0UKsyA15uz5MG7SSXp+zNtojY0yJZFnlkJ5eja/6st+u9H5ernqz1O
6mtwfUtcYKi/4JoWxi5FfphD22P4Oi1/Vx8bC3yA3C6BcFFaFOPE/GxPMOmfveB6+Fih60yMXO50
mfbe6umxMi8WlGfsxeFf3d/qNjpXSJZsFRmxTtNKNqu3Aoy+1xSTU7XS4UAWD9lqHbAti/ljIDuD
vew+wJoM8FYrcaYCc7UTMJZe9ms6CmRyXXhQqz1dnJf3M9+7JoxKpxXjsSbZbJYss+X3i7ZcjmZC
A7sRVCX69B+Fsex2oJCopQPyXWKFayfODi/WckBxBRSVc8NtEoM0SFEZSRFo/KI8udRmH4IIkqS9
Scd2MDnmXr2JT7ySm9RkDt3J0llyU3De7Gr8M/bfKk2Sn8Ig1HsbWKw0cpQO0h49xIB4Pd2ZQljh
Uy21kOnNa0WcbbIn+bGfNikDT3ody7JUnLk593xKZbZ8EsZE/Nry1caZeE5MpnCckch6XOGnm+uq
mAfYHtA3ZGqB98SNbCabghC6yMGBWCXXqRWpHE2ZogveQPAdNHrsv5dKTPrXYbdoVx/vxrC5tuhU
JGcIhA6AR0J9oXs5C71ksrhFAU8gfiQcwHxztUlxLQrnB7Fqo5rG4DVTdnVMR+AwDj9Yi6KClTcm
M0S1Wu9S2Vl/fdZhenlRLaF+hxsKOBR761NSK1ablmRHGtZ6jsT3C1CVJAj2EUaXMfF/XEiJ4+7F
nu+N/V15nfJK64cnS2kNvXGmxbMRhbZPocLwaSBBJC/HYMwu6jicRNnbaeYODSY0Z5v19dyrPL1J
ZjYlLCfNAVkkdyUgj6az8epz049q6Z4oiXtBgBd6P9yU1jFbQAcfDMNDhz9Z2ErfGmg+t24hI0wA
2lkBin6F5XbT/GmdlzeG0vLx1gbpzeLcT8kh9yRSYujruyh9Ux/MtIQ9Z4l/J+WhgGRgu75rpC3I
KKgEQ8IFoL+I8MaMYHbaiwmG2mSgxDi2bxBTWTX86CH2GImhIsZWd4RCmG2cwDy5TGIqQL/WKzDq
hh/DQzJA/mxlRWDX5XsaZzzRgNc261SXHZRhsz0RjJu2Pe6lq2XVkIK0o7d+AnFicl/JQCgH9n1f
hn9ZiOMw3YakavqE0gWwALnMVhRABq532Hyfs0INlFEhNKpcekZ3FQPYW7If2v9llAeRcRBR384r
cB13ywKApcURvckyI6MPOAigC0pmBCFRimkiD4sqwg9CqmK/SUrtjUrqe/B8icavDGLHVfsDdDVf
unKO6ti2EZGPk0YA/b/lKdZmTVThVi8OJCepz9mb8H6d0XL2boJKbBonQrFOf0rzkaE3YQX82vZI
WZKSixzVk4ztf4S4bBao+WArnWEZo3KNxeYeS+osX6927ybAnApl/TrikzU95pnmcE5sLEj8Lox6
2H5d0WRwqdA/phxx9bs68ZwhLyYY4//Ub9xua+zMb3IEv1lq87MZQ0hrwS4M3uDtODZjN2fyyzsT
EkUClZPGr4aTc9N3GakHbVtnNr+Y0XheStE8LNAKY8IOEXWeLE3tDyQHU0eK8U4KVzYyvnoNTsJt
Fr0SstaO5iTnw25B3yHebdWPoFgJC2NEXpP+OLCzQoza3xsiyu4IFu49k6jCVfzrAMCOSU6hCZim
k/FPHzDjoQQHR1Y9kHTfFv4MBRa9fctZdP8r3v8LKok9XoihQTT9LiKwwZ38Jr4swqn3hzSnUjY5
+H9RvaA6LEOVETSzSqo/OMSOoyrzwVt3yPJeXK5L0grSm+W65LvBUOe43EEOfHjLm3x3wAUAcDh+
A8pOrOdVAO9FoipDP9ZnRR6pCD5VwF5Du6xtd4AokiuTHm8wN/NeIjtMLhJktdQTpTdI8ORJkoWC
+k2lRUusKVPFL5M8QXI8CTPGH/kVMyp7iFvBbM0r/n9z1YdkXp9Ot7HnOHINaY9FyDLRYm9wy708
3sqg7Cffp1LUCokgUCBU0fDWq8sxJgZO9RvvR62M0g5CEqM3iCdTFaIiwq9tLajmmjUx6aZNJP8G
epqHBnyVMaXkikKpRu5P5ZTXzoJnKZrN45ofc3yf+qq2HBsysRh3TOpVtHLYuJrp5jAkAv56VBR8
vqDqnQOKXtQZWMdeQATB0dP3voQshBGSKMH38deAcPgD0TL9RI8CrueGSc+65/8UO/oTxwTAMgz+
fG+R6+b9zUzWqO9fYSZ/J+Us7ZBdBgmYFXuOZ2MGENCUtHX3AY6eC3hmPrQNPrtMzK2NW7dklnUG
9IA/CuoZ9O1ijoTGEFVijXsv9fkJTlZON7mEvetCR4KlVtCxzk+tkIVhSY6PmlFKtoJBKcpGSOng
1YH5oDiaq+0s18Zno7Fjdfy2NKcHU+uP3Z3jvgZMJ5uDfpc1sRUIg20m4aRNSfWPii+LuNTH9axD
F4mNurLcfiPJQgxmXbHbkdUBOl1Kze1HGN7b00xWhPQatbVcUbaYPc0CAMzUPsaumiTPuKDFmGZC
JGn3GWjUQOAZLrqTMxwSi/KhxN+8W1WdCon8BaxU6sJAwgFhiFLYX1jnQjfsinOSYSbb76Qnlue/
I2OJdIMu0/U/0pNxgVGsnDDeMT/nQx2gVYPoV7F/N+2Lf9dPJZb1EI4a5dlMDm5GLWt2tVeiokta
jNRXMeHwoseBM4RuZw3p/NtHbM1gxWlK9tgOJ1Gb5Vc98JLbxRG/L4wjXwSRAtijSqYpJ+gj1Yc1
U4A5KKzK3ZPztEmQu3oUtYqsYI3vxtEi6fVapZlGUtOq/9FdFlwDyt3bHud4Stk9P7h5vJIZpWHZ
tvkudnczLskA1nSvoKdksi9rUr3UolnpnjD6Cys6/mUkxlK5mP95Hs42hDY1U5xpuCESe7Pr9IXa
ilZos8/8/ah3B/C55X6l0bLhdCsfUx337E+eEH8DCbPqVCJOrnwJWbsQutFARQ2q0dOHDFdjgU7s
YKNYYKYFKaW72Tf60u9xv5FpOAppPTOtUfiJNcdtncRpKrTpR+DOYfDtPRFdERdewVDZ4dqkFMdw
UlhachEr0pS+q14VxWsIHduVKSBhCGvuUw6VtFb/kPxfCH5DGoojQHxFEbp90L0KdzFFFoEV54SQ
GOa7wA0dcSSUHsONtnrEQnLJCw1/SKGSVdakhTxpTaZ84CjQdtKTzZeWLNS/sJxGnBqFHxrHSTW3
Q+aw8h+L1g1DSWpsi9KChmVenC9SWW6m0IjhVzkC4i8q7b2CXkvgaOsHadchcf0blGIulY5p340Y
WDBORAKI33dXF+zZcE/qxkOJxfwTnYThS7VT7RRMv7K0uWEBgdeQ2fS9AAdn/5HXQ6q1pJSBJyNr
Am6SEffb4v4jbqygeOhgPeJVVjCKXKHJnUomCqY8X2tSj81ea/w41/zEew4XbQprmpQrFWq6atM5
VzZcsASkV3c8OZm89RseZRFUrCOA/kNVakxx3T5T/Cz3nCvG6R7E5g1UrkNyCpGwzyK6oDV/+Z06
uf44MpoSBTLDp3f6170ikJs4/0XFAFOZXaJtfrjAu0r12gte9BYGbZnNQj7tVZJfdfjFJCPw55Og
KIgK50ez0QUMpWc80LVnBHkHydjEh5W65oQNCDERj5YEdrigsKsO0I+30kQoRg5DHgoFLUQkBQy7
ZNrrrEhB4FpGsWLvrwK6zkSPxORnFZGZXlKKI7WESuFsLWbcm6Qnbx3sBiZotSb0cPMpgLQ1e9ji
6ehXtyhwJp0RMNO96vtyyDc2qyRc4UVZlYOebQ63+tKrz+U6m+LqPd2342SbKoALLP1UYN2Nh6Yy
iNoB5dhNjT9+CvWQospWZ0o4+IaN6UnWBVjdlGT9HktV7PjH4RL7vcIR+EHhHfd2JgnjdZlRzyjA
J9XRF/T/sNpkyZfuUO2lhy+D51E8+iLveBjoj4RTzeiv0tayuwlqnu3LvYXSOH5ngvZhGnX0RWZw
ilqpGeJtfc8FndzeGAa7Q7MIfz0Mz7lhphSdukTxrOAfUbnJlCTNp3iwOoklRrJw3P7fE0KU3zIB
R4OSLhBUTD/9QurDCHl4Ls7HpJLgSPuz4hktwjPrcAqG5FhNM11uKScyeH+U2BDBWSPE8IewfVaO
kKHpj0UqYCB1htpZjwocA8uHyxKEATbecBjDK55jUdnmtSe0nvmaiKvk+etRmbspeOu2b46NSZqF
tLrKfx9hfaDm/O2FreJPsjreH05tZSaQh49h4K1uh/iTGiX8yj2b2MSVpGyX8mPRAx/HqDi71M7Z
XXKfx9AWHNLGJUFxSC20aDV0YLjqi3yNhSIM3IZZdZnaRkG4PO0zFY1nDiJN++n+2F7D+pZSgx9W
rBdruiu43dU/uHHtnqO8GdEmN0vuG+g7j6BwHNRb1RlRARHPaowBdNqDtJdA7RS2hKA0xjGWjZfp
PtLgk6BY86X0Qt5nTmvbFUi3iHafowJRScQ19to8/Gwc2t7oVpJydYmTenAdEM1mr2nvoPX0pUI1
RAbSuMEIfnCrt4CJ+smJ1J3c/TE4Fd2SJSXd9Tb2IhJ5903qiMqsf881hmTVCwIqmSpotxLE1lpK
8nF2jTTb104oyNR9NdLdImGjdcY5PoZ/4246BaRSnClF7TUfP9Kq9DAU4ynySvImr9A+UIA6W99G
KyscvtPyaBE92qsJGo1RIqbN2TItk4Ntz1Ma4jbtWYF1v3w2/zoFuSBoHp7qwABldmmDAwoEOvVs
bDPDRxDlDAKQTKhZ3u4VD7jKXYkx6iWK4fm8bsIPBZEtKfXGPfpPcXo2gglW6/Dw9c3Z6BPA6Bg6
BOz9ojM0v5/VAGWSSeKFXwD7XUTUs//TJ7mnQf6FsGMwcl5Y1WEYSdfCmJWRRz5nliaokFBW76gC
yXUGXvOaLJ3FMvDcAisnmlP2YT+XAFUCa7YGJK3Ur1y67uF0lMiV8DONazFBAPKJ9/jFxlqlVWi7
9y6iQ4P/0S4l7HaXp+o9JB3Xkj3YQeouPRuiGfqlanUaL0Y9n3q2uPH6njtp4FdQmwp3ubX5bVr5
hDteuKo12vODJq94aNsXDNHiEDV++qgWkkGolgCKvbsxBbVGCtnKKMecp7WjGwM1S17KXAZGIxMb
MIUwtg9FqmS9Yf3IupIsPerU+eRg/ssdcGWC4OFU8/8zr2J360VAamuQyBAqVNNTotGgBqGixQJh
muIor9FFqKwStzKsKtqj/A76/XxK2Q9DOxrxaYCY0ewXiM050LecTz7ORDLTCZmiZA0/xWL5xB40
V2q+2BOVUW2lQI0jUQixXIdbFUXhKAqsY+SelVlNqIKU3X3bh4Oljjh1SH+V3S/30rM1OI3JA3jm
cT9M3jogkK928Tua00WoWXdv8pZYte1WrKI10Ck8chzkC5UxeiLCXZAjsJq5qlfulpS81srA4Jci
fAKWLCdkfPNMBMehEIoV2ppdJbjmMP7Ql6KrWlj3eXFYYS387WFVYxdnFTbNfj+Zb/Szi3w5GSgn
SBm0ZN4OhpCXg9IkGlz83UsQngV/mxuZ1vEVj95+U0IyM9EkhCZgyv/qaEsWBdYjLHoQ07rR+WQ1
Vue8dC0b2qU8ZsBxMN2GnuI0ebryupyVpGDW1ZST3QUVAVtWpsmXfMHYw5fMS1zbzr3AYe8c5YPX
MnReyTGLenH8YwKsPvaEvKuQRmTgAO1WBdxIS4dlKkWo8uomlU4OhgGyoBKMKvveEnTz5WsA7Hd7
VZWjvz3C6n4eZ7u0srqzS44B9cfLnfIt9zq6VhHdzrX4PxA372nbke+cLOX93XdXT/E8T1/nkH3w
VeC4bdDgtpnE0vzQcERnOyCbS/xtZiINl5HlANqHXwkqqo+rrjuDbKcThjQOpxWmW8WTFJtctkeR
9YxNtfTblXpu2PZ5pUgDCn/57doixpKPubX7CuXzc3fYdSO7EfsirNKgzyRT9NfWf7zL0uUYQ+x8
0TmX8i9LHraC/NiuF5Noo4nVx7UKq3K9D8Q/4/yJUDlIY9y/usz7nyNrG6WRfuIxJDdDnAN8Gd0/
8r5cQwhqPrubX6hi7F6gtHJeywovU3YCyktBXgHGBsoQbk8lQTemLEgAEjPADyQnarqqCYlw9xcz
TX+vm5RxYZgz7daPgYpPr121piFCpxEvAMgWkt7XlW4j9V+da0w8glBN6QjGdiqsY+2c9N8nZgKD
qmz4GyQ2z/iDF0Klm+XBcdyPFDgPo4zVCGSoxOCVxu59GpftFN16fX8932gV2cSmwPnJXeB2BJRY
h5gRRqAUKfx5Qr0x8eTXP+sV31L/bPEq2ufwnVHOgK9wPhp0hNAYDQuYYGaBD3nAOnjRBxHvqLH4
gb7wT2COT0iWOeyA2IGR+gtyX1P7dES/WugKGdaYl6+pv6Hezm5JgR3io6YCEeodMguk9+BovOyM
EmxtGLFBmrVqG+uR1u7o1SZOUYI/ghVEwyM5wFnAjJfCdcNuhN2cNZxLdO5eFCK/oJREypK7H189
k3RfUoAQr7hVthjeUbViNlRacgBBHZqDtDeUIXM3yY209ioZYVFJ0uW6Vbf+2p0ibT9JKkbxRHgL
N/HT5DduQDqJkeq1eNTd/wgzGvt3AoeKmk8BGWQVnXed+eP98rn36NC4kCPv6dmAUW9alXF/oKRV
rzCOaBgZA0kVZGnCi2H+tI0oxUZ5ZdsVWk+MfhdNtLjmNMy7d7GfiEf+qIYgvpx0wttEKMrwyUBo
teBJkibqn8LahDTsErI6OfO9rTQd9cMjI0NEF2fgcsWxmYHzcgeFZGMfsd1+P8gBZ95zlp8eajUs
RqMS6WsjtW1B8vLWcCUEK3Com6D/DMDKnaN26l1kKeaJZ1F0DDScJemTF66IpPBXDuL0NDKPBmf0
fBCJMlmHUGu45x2VHA+8QWeXqXPdukGoly+n+DTxHV1W9xSd/IMkVjTBWEavNiGxw0NPYhNIOEPT
bU+RqCfEVZCbhlNF0NuS1kFYMk0uwLwUSyzDJK/ymZSu4Dldlrx3bqFNQ/Smw8rchIWBge0blgD6
ln8jBcJIH4p9HzqJUvD3Q262igGiahZQ2BpvN+YivpTHdu9nUo+lmzdnR+akCghRNwKTv9ks//mg
lRoODLeR/fwVI7FAzhFaX426b3jrl03wTfVLKBHIN0+JIo21kbt1qPYBMD2rylElxAzYkHRHM9mP
LiLBtUK4OGx+UIVSUgMpUxVehtigcmhH+G2pqzyySi2Wg15W0B6+9eI//1SB7OwhYSI0sb70p8na
W443GcS8U3nqGrMPVAwjOISvV4qdQ9cYx8isye07UX/Wk0SeSK4BwNWH+zTIEyYzYviYlflWtbkk
iwabPSIao3T0nWbDpeH4N4ckhyBbERLhfQV8SSNV+p39bSpXwCItCujKZLX+2llX2Y/LDCT00VPF
aarY0uuM0pubYlxVBGz/p9ujln5SFOhRwZZYILuScSn3ZgQPWRBjIJFx/iJeie5AZElSkRBqGxBn
R09P52Ztrk6MymXuqv8VOZ199M+kxhNayRtpzhsaKQLCQOvl6Wq6qcJWn2i+3P9mRgRCi5zI8tU1
EpCYLeIkEqXclDzknPwj/jz8GUS+hoXZWd/9O2ca7cRUtY0QyXbW9CetgIJt09H5aKW2scuLO+PS
1tePkf5QaSrPMM5n8VoP4NfmT7niEFK8IGlxuNLaMiZm4BN/hNziJGbK4eOW272FJLkANXfGark0
zMRblhUZlEh9S4F6AjBXGFJ6Zufun3HhYiLHmdwieDOHLHQQWUtloCs4rOO8/oOCTSrWPKqGLiQA
L8bm25SQQv5JdNbFexdiqapQMILRPei249BdQ3W84cXD3guc30xJ11jXWBJQR1qqXrE7fRtBFR7s
jMPoCLKRHfxGdDDy2A1B7ZQi3qcVOruqxwvwtu/x1VovJKvmYs/s2Wl1FlUyNQD8jYjy/JJl7qUz
qvRypZWJbaaiNvZB7bFJ4Fxf2Qf5vKtwNUL7p0UFfjrZJFI3S33U9vIfJeJ/IW/FWQN6lMTOqkgh
DL1q9s7hnZswFzR1Cv5U/l5sTdm62irR9OduhBE5BK42TKqEB+jhXamtPeuhveurruRf55NbS5V9
/jWE6LJLLHYOfWFii0DBwa+irzsbTdMQ7W5H5xq2TrbhapGHAhMq0NBpo8xia82NujNWlp3BMF8x
IGyoREpcm+IRKOrbJg5zT8ljT7xzlIo12alHrr0cSOpjmpYqH3coRaGNt1Z3GW2Gk5taoHVWgybm
71QAqDOzVHQT0adAkRvT4m3UqNiRkrdZJS/rn7wXBQeh/iCcsxcz72gx4kDDBuOpX9iIQEVn1xPG
LMMr7jAZ9099P3mbPkG0R9B9o11a6ciZ7ggYgQOZOLxgzHOM8MatdVlTEtVgmAp2cYtQegZ1TYFN
5Oahn1ucgK8YYb6EDd3ees3DJe0HbEsjd9W4N5WqmuDVsVYBVNxpUZJvKEAttEURj0z7MW/0vGDn
IloqZO5hIJkwnyQoPv15Y9SnisNAfg8twhFjnFTG0azf+GBLCN6WfFJJyBeN+MXZq2IDykC7AOdN
85fETQHgYSouXK3VXfUPWcwbCIFhvfam1W4pjiKWwtWGjtoldswG6OKAxqNruLi4Pi93QdaB++q2
BYSaTOGcCB0GCOGfPaikVQnhQPwHvXqWO2Clhbbbm+uk3mJ36yJ25ntEjcR9Z9/qMy/7WhnJ+1uu
8APRTodt+OifiUKJKBE1Ji/YACpjWc+fCnEfDKj312XDODYDF7lIl7kazOknMS0OsFwV9n+9x7u2
jZx9tHZcyjL66g/WjRfq1A6Vpq8lLbCDfnmYeabPj0CLx5gyjB42ADpCLdVnhP+HtVYasT80MShG
8R/4/WS2LPmOXL9RW4AlX4mX4bt2TGLFX6wfJCbRJ3eoJruVSDJU9uIujx/+w+NAEv3LJ3vX+Ss9
hTwhr6+ghnI4FPzMcmDMHduqGapYH2p/GWmqrFl2qHM+aT2lQ+og/GX8iqr6stoP4T1GGTYe2kQ4
SBIqRnNDrUCWTXNH5dTUMHbeoA3SLHwaZSAiUSFKdDe6zMWFtQrBf3NKumi9EA2iZOfCITI8HrFa
kfB+xDNXwlUsGZXDYKMM0Ybqu9o26tj7eT+eyPSY5lqMo18DRHnRlvr3UFF2QIfnyhUDqHTqPpvZ
o8VHHDdzEppB2XvLfktTY10csz7HbMwwoMx5r+IajnWBCLiV/c05ZedrN34CpdDdrVdoCOQwMlEC
9YKMP6L6t6c/UTuIXGDyn8ZNJczGYLxHjRKWFJP7lWeA1IMlswP0Z1jQVGv0kEVaArSjHjjkYPfa
xLPbcLh1Xhnivdsj+PLUEqibGdLWDOxicVpztNVkDoMgBY1yEqIdn2iuNOBDH8x9SBvyAsi9LAx2
0WAgojTW/Q678bMGMx4z4yNPJ46I6NopGfUKCFiI7cdHzUuKYWggq4c2pAfHSRW1ngzZb8ds2FPA
Ba9qV+Vy1+A3QhZanDol2GSVUOtMgPVNPsmkIUrKTjstj2AWmPy1H/qFB+IbQAQ0+NFkqCvXeCJo
FPtKjw/ib7sl/bxKxLTLBceJGYH0jS6PdDMBksbIPAvRB7Cx+yetQlhTRQDrJkwcwBBDjy4CvnRF
sbX5e3UZjZEJxpEYVZ1h/Z4GYMTJhVbiNxy2YnugObegBG/M8CAV8YcWfMnRZd0Yt0CBCf7fqlh2
NnuDh9/RN+MrJXdv0wSNuum5tXAmncidjetSAeEl2uNLVMOeCwAFrFaqL04AW24XK6i+TWHS8WjE
74+tefTsSw/jQzKRoicW8O+iXVlkEon1NnnK1nXcTX1LkLTE1KiKAhZYTyj8YBcLzbxzHlW/v3uj
3Wc7XW2Qs43hOaWN4hDSdcIjo7LiEZm0hU1WTZzARLW3pmHkmRDzRxViW/+X577cTaJoQrbrgyVD
hmi2uUObE5SHO4u6arsmMT7DxtXnnSfrByjVBt2eA33qgmWQFAJGmOEmvgZWJX5szo9O+JNbij+f
SGn00mnLWUp9FCMEkdczigR9yurz1n7cM9u5rInbsVy4Ix+VNvtLme+DDhzedmxpuzWYlLlWqpYd
MH9DtHIvDSV3d5GIKwq8ULLvM78COF5PSBYr+xrDBXTX6TxwL+rVE04Y2LdrBtLzWd0rWP3r4hZZ
WyRCl4coKsC1x+bEYlr3E9+hS0rslV+KiB4+uK/CYPEIE9gdm4Vc10FjrCx7qYRZAoQQ8XAmMA0t
2PnWiuuJrxSYUuHuiIwfPOv9pPvjaSQVvXvYFWkX5VwAs7ZFxQt4YoxEcFTcXk+7NKT9vpLFoT0x
94RutR6X2TX14JSsVYBbYMI+BwX8dI1SA36KmMzF9N90beIXBdBzbOyvNuHOOlz9tSHHkaZn9TXr
z3BmXA7dgqkXW3x/xZ7dQ8r9xHr8a/YcU1dVs+lqCOBu+/oT8ttGL3HBnZrwUNf2799MJFwwl9r1
6BOpnpoHFdFgN5JYgeIGnm/u/80EUQXC9C8kFBYhjugHLzfKR6pconUVQF90G2Dh6Csjo/mucrJ1
zA3Lyq41ABT13oISR3n5nfPW1vHutB6ZOrMXOtegnZtHX52s2ehbbml/rqVeq0w9XQxtec0h4YwT
RTJTWRfRx6Vv33NXijv4pCKzyDtth8rAy0D5gaFWmI5EpH8JDF6Y3WIVv/1UjHmpJN1ympZvUnzv
5kuUEW64u+8ePRpH750csMwx0Lgq3+6IckF1U3GAIvz6GSxpwStcBBrtPxnJzPdCJYU6d0nwWAAJ
L2KmOE1hZEkAScwLsxA+9qBg3GZddkPAHcdJgoxytyqRGDjSblaL+GmGR3iGZofH3/f6Vs6uJLCe
7X4ysPfJcKqgxSewYTrf/mLnF1wrY6JlGHgzaydRuRP9aGDLrHcXOeEJiROqE6VYylZAThdCzP+J
VydhwNuln8zRh3yUN7ovLOo4btC0NDpW5lJiWIf6jR9UsZbsrPyJ6XFtIcxBMkVqdY8B82JSwlXH
6FW+anb68Nmfu7nVtwo/EtUhPC6SDCq59rZlxmUHsVnALXZn3trhIwwz3H5xjrJNlegaZVmqh+0V
ViFZuyFH+8G4dokq0r2qv5yLn/E/Otc3Vq02/3zDGmK132owoaeGKQg/AcyXhWF2YCCiTpPnFeAl
TLmT7HBtRurylQDOe/Vb8nsGWOvB69wHx3nC9WIy3ARiyuPKaQqgr9SPQmfmC/lP+nq8BcdeenR+
hHkc/mk4WOTN3az2YHd0azLv8g4QlCbPs1udk3g6NpvRmtYTzsHTtA8rC1UOt6bpHzTOLTbUIcdd
i6NcAFEb93vs3qGDdiV8i8QIHE3kl+Ma1jJBDgUjYLYpwBv4FwNDBwdpyLVKmvNW5Rnie+84Vlcg
O2pa5y7ZerYz+f1WGTY9zXUBA1hL/lbmHhE7H5xB8oRrDO/DW8CGCwrUyjOL7bxqOaQ+2S2VTCxa
gKdmEZF2ZgZ/R0rxba8hDgtMn9OgXLqEIlHkCe4JcWyn8sYsvHa8695x0iwq3fmJgQyeKZOk9Xa9
xGxW6dzQOeefV3n+hkbk5jPVhvmM9YMnMMBHjMEtx+tBsMv0xHEHNQli5o2xzLmNebDvxRVXrNjH
xbbah/Zw03WY2WqQ0pEGy/J7vOeMk1897OV4Xyq6oc995jpFTDlvihtScF7DjBbfrDhmrerE9IlE
o4JmebNeGUGx+gNNHNr+aOhHRV9AHPM2xoz+mtE/SG/LXZiLWg6eGM5m0V6g3haGBRUkjAuQbKHh
LO/43/IIHsKFA8hzyjRTXaK/FyttmA4s/Lt4coDdc/wwORg+bTtvfWzGSNjWAoY5ZzwAEpZa2UVZ
1Tl82N7qQpE7DFbLKJrpOxEXzcZ6LZZMZmAMJXqchvSSE9J6Qf+eVV53mwluoUgteqKFsnKqRBtZ
99vyzaKMdHknsEeG72HRasShkwQfEbqv9qZjQuvLPm7JG+2R7r4t83NoDbvE+xPh67iyK1Mh97oj
IODHpMAZdJDHZt8DboG+1Q9Otu5qcW+XJHrH2B7xB3nnOH11CjeN/3IETCnm/GQzJj2oEcaOVLdz
EYdVskWPx4HDs1egCoh+WEwoL0ci6Ihv4sIqcsUuTfb4g823gnX2D7oHUxkHfLHrPPfknsyZHPuj
8FbojJe3SMIV995RYdANsL7tTjxK8mKYbC6Zf5h7JX/wUkGzpQk1NZWgWRLZb6YkeOyNj5kx61US
9ACOBHlwQbqJpheH9aixYzRgBHYgRpkBEyueHyEzd4FjxHwsM6s9yfy4V5/luBfr9F63tF/rZLf+
730q0ocELoWnmEbnFqObsLXbiEhdg29EYJ8lK/TzsIZo9VgZOebXhJivlgKE7uqk2Edghv2qN9bU
QR7hNoL8LGEQXFIBpZnAIKhYuVSUSUrl4eclemfrtVsqpILbBj9XgO9TInVoKOWneqQG482ibUXd
uavGdf/Qk79VoPudp2pnTlqkNliUNrKHpqbk/v5JgW8SQOMZZp1UDZbaiQS710dKKUZx1YHFN4+j
arbUDR4renY55rzyxTFB+rC0whxoM+1aGFtDY2Fez1x7KEL71pw51+8EVXxjV9ak5LOm1PrQZAYj
FAijOkiFZtau3J0vzlAnG+AJFZ3rnFZX2LgGiR529lU2I1iwjRsZE0Ct4HTSOkIr5lGrTKPsaNaC
i75WZ+qe6jndFkE1tPvxIuQNbayL9yas/OQQ9luFEl+Y77w+cHPVNj1Dkz5xA3wLmszFLP+J/IBD
4uloHe3DroRGTZPqDv020cVMO72dyyYviSIfFIlpi1bYELPoWlDd36G/0Li/JfGWGTSg5JPdnV8x
SJqktGag/bq1dAg0/z2SxBIIrFcEUIrJe6KST4iX1LphJM/vKaxecWB5Yv2lw62e4lzUMjpuULRy
wYbqR/+6wzBgtKyTbwJOph3LO+Tm3krBywmxzpNX1WvnLWNQNtOW9+QoHhv2KuaV0TeTjmS/o4d+
Tjt75JSDVRgCF5sCbfzxUEdF3XTeDHUo6u1lZwQjDu/8LIFKhZdXGNmFcMmH9sUUmzoiqc4D4cOA
0MNyH/z/26JL/Ot6R+bG2eJqwz+kk/ngM0OQb3/8indEHG0fC4QygQ7t6Qin9Bho0ib+GSUbmvyy
8bpDujSxFxlqoTYl4N8aj7hwIS1byMo5bFyeDHVklWYnqdSlyMdli9e4peTt0u1Nyr4NJqm5bWpC
ZjKB5zzekSyTdSMpg7XnNiMkm4YViJx9RLzqWNR03yCkVPw35QVa9mIRG8Dqr/bvFHVHA00HlWCO
ZSt47zLIR8ETed1Eg9ILbBuRBBWUJjbBYCxE8IaV8eUyH3QNZIhPU9WbIyxLqs5J5BnJCCx1Yki0
hiE9cr73G/wS4ZKHRbud37m5sI7NM5gK/OzD7hSI1xUlzshPWcNl+wDNBrJcqa8MF4XDrc0Po9fJ
qVe9Ph4lcSDe/6CPZ81Q9TTyXLkrwNmqxP26fgjX8dx4mRQUCumfmEENAjKBV2edIsorGQH75LuP
YiPXWidJuK7vZlkVzuLRE1sDMwnTHVcfj1NL1hqQHilRNRX7umPhCC7Eh3/MAyMMC+4/sN5HacbV
3Bzve4FfWcQOSJltTCUQZQJU7JC10tLwKjdfmyTLriIIlQCzmwCAlSSINqDpA7RdXL/D6armIhpw
4qhE4Ke2tk0fWX/qw2gYG06J8XJDa3Ocn7/j4XxY81YVDDm5s+y8yREPzZW9TxGvj8rFxV7mut7J
j2Y5LDse9IzLIKBwQ7Q39lcYg6FXqb3R8HJIFQgQBReZ8CvONHv6NcWCXAOBg/xDD+pfmrdOml3X
n9btQpZfn96Yee/KveREzSEtUi52/bHbMqUliueCWVDp3yKlNhSsJd3mlDAotRRcILm0LIDz04Fl
1mQkXOb3pT78zvT2e5CHjJBcEhpNUEcIRb/lYO2o1AptvzMPT3Uqamo6wVwV7VQQTCAuQnztm0bW
geBAhlU70wyAQieLG0WIHbWH3Q4kEeUCzj/MYq+3Zw39v0gIxLqb7YLvn1dSRgSwUaC0WlelhJEB
7J+IvYjnksnqibOQ6jZLFO06//hU0FkW0n4V0TBytmKzbLJl6LNllIjnOWzXJaUff2nvPxdx7mFu
MrwnSbh+4v9W4yv80dCmQ4Y0zKEauD0aAHi5B/dEfxBwtQQGe0W9Sw9Fri6+oZjo+GDewBotpm+v
F1AZPGWOPjENNh8T9KA7O9oOxYpq5E7fhjFKT947HJUo3K1utpmhnW/vgzo+lbtHcxQ569cXOgzg
AyQBtvABBqI3i0n27uJRraMygMjUVn+LFvZkDOsLAKUR1wO/5Ep8Ok9nZyPj8Grn8DCTBpl0iDpa
+8ge+b/5WpJb3HpOHJftY4v1kusmQAWlp3tdclt0P3ggpa6GMoX2OLu9QjcgRASwg8Yd2Nq7xI1H
pVuHS9T5x1eLRaifErZPYtcz0qbyKQcb3IO+N56sQp6cNlm76DxwwMUjeMAysM5swTEbEThUo2k6
jYc3dVbpK9of0ZZwU+TS6xTUDpo91P9GLnw034huqVUeR/librRk/uFOkHNK55B3RkVvhw7SuD57
B5YBmmP7y3+iEEOtYB9EaidVNxp4pOTpnJq+mB2PUQdNewuI+6NWZjUAO0+Ugt4+Ht2l5RrW2a8+
pMAiA1SgJXhtzmRWEg7pKFMQQLv5q9envi8nE8yhHNZGyN1GkHy+npl8NjgFZkBZ1y3ejeL1oDZu
Zxlie6dmHn+MjiQO8CKOj9bEWknMtLf7tJUBn10Q9jECC6HwzQ8KU8t5C0ZmxileyIVQb/JRMiPT
oIoIbltbPjM3To/HPn766R1jwUXLeLqVY1YQxKueViQc0lFJmfxN2L6B63iRJX7GpKTE8ZqytYtM
yG9tNdzHzSsAh7hQw9033znBwtT6lP6tJZm+LRyjZQsOH9CgpkwPv172/Hd34WzBXpnBr8t/V2Ls
FLEI/QoCwHyguOD2nBg+TVt+8tdJ8rnS5zU8LZUo5wPfXHBppYE2zv3rioaqm9zy9GxWjwT6gWo4
7VSrbAQpXQpM8khrkQNjrp3KStMRCpYa4lacGX0lHJ7+v6o/Ud/yHi3JktXYG/KiI/smQqJbBRXZ
QL5848Pm1ocO+K0jGjBfAcKTLhMUay1J/kTohCU5MQXffrKLhuWfioB7W3Y7r+Brz5fwwzeTMNrQ
aB9OxSOgwRtGaMA6/F7A8gIeFY7XDd5R0hMVwy0MV98yIt3Tj1SEK8ueKtkFo0sKDQAY/CV5qPfO
bBvvkjkyiM1RzodxraUbVz/lVU3+1lscVrsd1yreCXLmiXWmgYeWSzF6ptBG8IO9T4xwyrEJcW0G
N40secVBhvFT3AXQQe99BqLL4cCEUPZJpKBz5hXIzIIBfLuvAfqSPauOvTsKQwleAX5mtLALdDbA
RjuKDtX31Gjf+BMTMl5V0L0ch4kHkJ/5rl/tClPSOoSrVI7a/rOZU2tq54yL6bmMja3dK3O9kIHt
QzVcd9qGBkmLwakSVMU/sPByhLrtRNoXxBwCM/7bKWAoQGdRcUVxtsrubA4HT0baebZvC9mSjUlT
99dF627BxrVCqUeORFpe0hL33ZRmYhs7AZMHugikQ3Af64+9KumGNBJSmpfm7lgkWFoUPWAeQPQB
EtFTfjN47RkjI2+Jlv381R1BmQEKVb74Zrk/s6In3bM5nq1nX/ZBnSgltNa4pgtS/gAw4pTrctp1
sSRhzo8H7zs3KIHA0FbXob3yndH2DOLx2o018BTZCmW6/eqgUi4IxYAUhykUZ7ruwXO8/D2bD88W
T0ye4MDDUFQCtUCtf0tV4WqROEgK7FxThj633YU4+OvN4KX4WW8tfKbYmyPIL6012nT3qj0daNbe
gnnF4dlQL736as3VoDPNfyo/DX08Fa/oCsV4GR6kCfD2fSscw/kpjTEwK/sY2Facf/J6HtOiIiyl
cUj93bzm5soXRfP8vU1SHx0E12HSSgIffus8MAigPtTRJEOFLU0WbmY5hc1AujOMrNWrPWpPmsQP
IEdkcTTcAmC7iNflP6hrD3Rsg9SCE4ijU5IKPbP1t9aajSdpZGmx3dBDG+BrOBvcqqulyiJ8roh/
07qnXfe91D3RxqwnUHJHHhHwAsal0dXrA6G5kSk1XlH7xjgtfX3Jd20/fW6Wxpf90rESnQMqHo1G
oLsCngK+k5FSG1z3/8sKYu2HYgBDxEmSNh6oQ9nlUXDB+lS6d4Fi/pUAiWhwkrW4wbWIu4rJjnhi
NTg7SH70mKH/dBF7tOKzd6hFebaXpBQgDRp7adyKgeMnM7FMaEQe6It5DX83tZjc9U4aKJyqoW44
x5tiSaA+p46xbHwpDJPdtlkP/15PA00htcU/wYN4fGjTVopKLcGn7abgKMN9smSOhta2/rJlzV01
jHxaCbwpyBvMU8Ine3O4zCWuVwBLxqvZihKL1f6CAoXO2sWih7e/gv45wYXLiC3PRLRGwOViS8h5
hhi2OOXEgei/p0Z5ISHp8sskQLO3Ql0x8Vl0+WTdDmXRZcw5G0xcQvP8puitXuUITKaoIebilYNV
pGX2jHjWLAwT/tTD+YmSDWzUTO7YzWcgnsl0cOMSvjYmbSY5X0DvpxLcVHK2r/FWs0XbkdQxxnwX
oXxxljI25bB4EhD5Y98hwsrAEINAcHP9ePKXb1xheASyhmTEtTaZ3Q4j4ye0TChVtaU+CCwqn10c
R4YThO09ic2zazH4WGkggyb29XpzxpcwCxe8KIYj7aUwI5fs8UdydpL1i7Tb0CoL+heLmF1HQf1W
upKWzd8Ke3rwN0SXGduL1Any43aaIGBzAmbA7IeGJBfF2CHsidmPzPKkd5//zmk7SW3PLk/wX475
S+/mxUAHw6BTugRoUjYHLaVdokkC70wrYDaRsEQZEnUaDUB9OL86R4yAbswCGnfwgZp2ti37++li
bA4NqEpvG6tpTZ84gl5UQsLOKqtFLZnKbAoeCU/SFu9kzmR7CZFTA9B0kGP7pg63dULJDKJ/HVvT
XbfhAc2iQYe441Ys8ZEYndgOsqiT7zIhi1faISsgXe4+yb5Dd7zSOgphK7GCUiNxj4RCQ7FKTdIA
m5R8YHZdcohoXxeQq+7/qlDiR++9ktus04+D0R9w7Id8FDkbBsrkMAfa/+yYGzZNgkPGLkH9mszU
LCl7rqzbGJNxtg7HalVMO4mhtk4W5b3vog+4f6//5WERJGapRsmX8T4cCqdc1VKnCHth1neODgkt
9xytZwIfs7arPJ4vu/zmZ3sptgg7Ls0CnO81LMkXsOXD2BcmeTTE+mAwLhs7aSE9jjWOBwHAWZVd
ND/DAG0j3IdZUvbd7m2sGynBRWSUVrroP38arhrkA5zr7n3gAUAbAoRkIIzhZkhPBo0hykn29Dza
S1UhM38X5yRwNHMXQv/R/Dkf11JlKN10cHqVW7a1r2NuJAI42sNV4qejMmj9QE007yQqMtj5xZS7
bmxzK03NqLgB845OOW18BvOTG25jFQRip3wolsn9afuB2PyTa0u/GRjWcMLws8F4Q0NfiQ1Rq3/t
L6oJn0i6Dh9SHSGdor06ffZvHSvxOWrtXZ6WmWC8vjwLgERaffNwQZZtnO1gQcPa3hVU/NfkERCD
Ev74GRc6sPJvRKw0dIuDYWzvoEazRtgd6JiCSCUxwwnIlaUIcMSadQQL1QMtdRvPMvwXG0qZf5Hd
KKbwiU8CqRo1ybxjPffa+vIDBYkrQvURwiJR9QELi9vDlbnM1+HzZs8iFumca9Jn+ldshRtx4DsQ
MCEfcZWFd9LysgbL6vVstWqjj/aR1Z2eZg4PKumhlaRM/5fd2UHNbJCU5hoANvmGZ+Rramg937wR
biXlsk+zftbrX/cf5LKN/GGKV7Cd07HOGD0BmRX+HO0+48SRkTZFVE8rFfsEd6PtWdAAniVywL3v
zt9yGqfVc2A/+lR2C4J1HrhT68ufsJqEOu6Nq3FNvJSAwktWWlaBFeaGbiJM6RdX/ZlKGRHjZYg+
jAvNLK4Jza5M+mkV7C0uHtqhG4khir8rmaQXmXLH4dF6GQou7PRMK9HrO8o5TjD+hNArqTRAjghA
nLuhcHmbdW7llZaLB5LwcKCEDJ/7ArSGk8veou874SPMn7/+vYqIsHkEpWwlHRcTys6bRNKHOk59
SJ8NfRYw6je7HnC//om2uAlidRz3Pp8R67JVDuCczGS5BaJd+Beq4TB2jC069h1V1qsJWOzx8oWQ
aCraH4cmQgkdeT0N6yMdpcZniOtCoJv8d8bD2UqU4pt5E8SFukeqBLVvKcUT1Jm40WGDwvMzLynd
BDycXAo2MxXD6Ac/sQthIPwPgzH7mB2VVgzEQawox52oBf3EtU688+nKtJsmyj/E+W50eTroqvy9
kHaWlNtiChnAaWkQVPfXYfDomsc44Tyr36Wp/gtQaXlayPrb8Sw9qj/mS/jXkQltA1M4ZFT55wcW
SbExD9wXxutFHAyHOvIq7KADIdoYjeSlL2xAy6TQKp+Vh6f+OzIPPYGntm0v1f89UYTk0xZItq5z
Zj4RDIt+OA3XMlYxTVqAaxOTAHVuv+xL3fUPdVf83zS/IeDJtnmuoKcyBRMi/LVC6wr0+7/Mk4ff
PpGr8wuqpGdeZ89AnK4dOFXgsaCbF19nJT7bI2PtZePvUDx7h1srI8WckoiOrTIw0aTTjRAb5jNC
x9jEFcEyjtLf8QbW0XX01E9qlzulHs+GHa9CajAJnWoT1u8JZj0KXdxKtIQYLQgfr/TvsVU/vfWQ
gskUP191F5Sp8NXqwfLcukItRT9hOQzwUVkMGFYxhHI/mQ2kqeSKCHDzxtTsFQYoXO0SF24AfZ/H
FR39kVM8LOSYJPjnBEaWoIVhnVuu+Jp0ypMDAkhICCx7RzrSBnuu8Gnh2/Nb6x3Q8gXZ+HcnEK/A
NMRs5iY/J3TR2xwmNgeoWK/IeRgylRH1CRQmGzqAQI+ZD+ixmuJi2AUnTt4ewRMFildQ2UGSth7H
+h16NVJnQceC+AXICVg/VGlvJ9NoV9l+lgoo7BQ0y0baOe1o+U3JQw4zm/vBfqqm22y9Touj6wwm
OLueyqsYzuT1E5RAMsFaqwXEdY0A6OIWx40Mv8mSWYxAKesAj3lnOcTHioA82DJbQCz/hvNRTvHU
xxqFVotE1T0+pNnPdzB6GSozMayKBS0dgaXpIEfi8GnC2s9qeSOTeT3hMzTR9qHw6SvQ285AOHNv
jE5oNxUpZVY2pNdFuyLyh3ZYt8t57yjK5eVb1ya3RuVxfGYtKnf0Gd1F0UbW7alxSyhkCqIwcDgE
U9ms4dTIoKxMMWthgYigDoV+HeH2i5Rcwm/09ooRpWr25U1c0UmS9dgeiqlTblJs1O0gW5JQoPZd
2JXCQzThwo/xw2ScqPY+Jiq19bAhmgdb5VnkPxLzpng6di03sQI7NEUsSyI6JLhcoJzsBmJVMqn4
fNZg1KIgnvLklneb0S5zOKmrCNFfQ/QZB2zdSUQK8a15WtFentUTycC1miREXZRNgH6vHwriIcZm
+ntd6aJ5s0sUfVJNjIqRJZrTPLjugp3w8PUbr1NHdkOuG6CAiIL4t8oUjHV+iIjugka71XX4oS4n
hsfO7MqtQqMXiUCUouVk7FxUjCTKKNpJn5W8Hb3Qr5nb3kwWC0FQFDSP9+SUjr5V3Y9myfObeboy
N1C1NZ417vB/FLEX36kR4nyyKwqvD0z/pdDe5JZot3BnRtEM9/k83HnNBb5vV2BGWjJRVoLj4R8e
VQ+ZbOyyRQTrlfMeu2tPlDnIKSnHiEqi4WJO+DB0pZP9e7rnsP1KhnnBsRX3NJucxNkHe1UNJT3i
gvlouH4WulBtRgRr8sDsc9T6B3Zd/k3n3T+0UJLTU8Ap/qWrSnbPh2McEoBlqGlKd+BMcL94SA34
A9pR8HyH5tRFcF0RBDyllFXz9xZ9TwtzQsuh4QDV3UBE8bQIzMiJ99QKMBAvzihS0OIbdOSvvbkd
2cpR9mS8Nwv3/1bGeF1Ef1XcSRGhobp4p1lnsesc80Ar2D9mEvyuh/Rj282dDZh49OnDqvL4Ityo
Kpil8UDevjUsTtaEJjxRwNJUWRyIY9oa1oQblP7HFQD+p8Cgl99HXP+wiPEEiudhaMmZgcSDVlHY
UCskRxJ0AQePH9QbgEm+3nt41erTtSuwda9hd6qGmb9DgbbHkSUbxBJTl4Jyfa1ZtQhEOWan63I+
3D7DxjFmUYMMNIcUmeoK329TvkbBVUI8d2GwCKNzGOTj3qo0SAkwH1Z74hXr9/v7BisdzOIMrPTo
bsx96RPJEFZoias1dsAnxo3CfziH7Pwg8ivBhgxbijwAm55Hs7P99ZTIKi1ECwTi1ZUV/Az99B6H
bopoGiizRdf7JL0VFIFMObJ+LmkBjgr8JbnnSbhJxZGIpIiFchDY1gG+6xz6VbdpHzEku1c4ektd
tT6ENQyvwugd2BRq8JQKk2kTKRqz91BP7525jRRd7MZ6ylG4Mv4xOQoFi9ID8E851iYuzRlemIXn
nX9jCqKartWp9HTYCwZcXPCvAlarfPu3XcWiux0pBVrOydEH4r2iC1snQdHbbmMIfhFVI+I5ThbV
lQqFQvTkZTcGg4TDhBqEMtTMkkehPb/1eZ1pEYXkFu6ZNstfjV+CVcLh66KcGEe/ZxypOGrfgWfZ
18YCGiuYI5hBn8UenLUAQV4xTcz1sAKslJkSZ//bfqfGehHB1qACBWeAXKbgbwBfpHWnIq7VxFF/
hAdM/vhhXLkqAxt5/slKsF5GlHoxcWJQyHJOtZAdj/3hkqhMYMPA+GPA/IKW8XJlUsVpq9R9TFsr
J9w6vD3r0E1oBw6klPicM3l6MQhF+SSLMC+LyTIsUg6SZ8IVPU8xVS5dTpMphLbK8nd33B66e0XZ
+gqm250TfV7n6QOdBVwZIGG7wAtNE3ctMthRkpr0YHMtwNJhdgQYkAUIWgbprEP1kgI2lVcV3ufD
1khbrnmIuphaDWFtIdX8SAzlF/dLfR+fgSzs/4rN2Gn3pGN1PkwnoVJ9hYJTcw2QfRJK9NHBg3Gd
MSmQRTAo6M3aSEwq2PtTILa4JksBTDk8sgsTHNWOM5wl9ookdMYoxWgXallJhS5LuplkbLc3XkZj
gC+3ypX+7Vz92m5VxFPEyccSxTMKvBQT+Qi15NzniAbnMai/TG0IbLfIN4tIv17tlBUD3mNLBnrW
9xSOfKSlvXsDcHyUTipaExm4owxLSabYsUAvghSMBziNIB0QCbabrQk//4gNUGS9BFVpB9FYKrxG
1sHaq+gZaYw/Kb9bfJvkXgW4Z84w3A1gjb2lGmTJ2+nqNSbtOi7CBfPezdGnjcgaUOldd9mA6Ayb
RUD3MQO/3okEg6o2GVSdcEQ6UMcJs/cEfIeosZFh+dP7bIZbmRmOJZfN2Nl/NnkIPkkF2z7fUmve
FN4Y76kZZGOMM/fEwsNHIHSM996hJeZ2hXLSWbMjKyKyww9K2mX9v8NfpjmrDZwEyxX2qUMHUV7h
/r5XDPfLGFoIMKBus2FY3MhEcDpZgkX8bubj81aRlviV9/w0sjo+RfoWrAVxs9eL+jNuNDommOuB
qjz4MB855iU/8dPjjKyOpGr7UrIMlr8wnOBh2v7+HCDhNB+QcAzCmsGCFHgt08LCwF1jYATK1jbC
lWtwDk34ypeNT5/QZ34e9zRyX2VlZ068gSN/Vx+iFIkQez2+hrG4uWwcl+CVK2KdBo9dKW7mQJCS
4PDS/g8kap/E85NMR7TPaOJoN8CMRcylWPz/thcr/KZPFN0FFLTd09zLUFB9jxmCUeMYUWz34O5/
vEdCS5PzhZXKUAgknw94Cc0BgSd54iad+WGn2VVvFm4wgxDW/pX8pK332EbpS/sNAJ99jaBgT0V4
otYLll664S6Il/Xpf0b0l3xkbzSgY0Dcd1OR8cYtLFq/sIav/7waXwkflfyYRM8RickpeHG9DKZD
FVDGkbA2w+QDZi1AVNfqzcO2AsX2mt23wSueKoQBhux0BfN53N5kVS2S9PKs5AnPEv0Lt+6OurhK
HZ6YdbW03f2P8LnO7wtviX3Y40ghzAxSkF9fPNciPUkKzQBEEcxWJ5X0ntnRwr2oniPdWQxzUtrg
K6xUH2QBjMjyciXgdZE2CGVbCFQZB6s6E2ioZZLT4TWWV6bH3RrNkWFYAEKyXpVSXFgXB8w+K6WM
tBRBWycBDKinBX9acTyxRMo6lTrx5mvuXPNbHBQ5qBfLyVLp79FxHZsT40zKNt1U/z5aLIBj9R+j
WBiFO5bJDCd13v/ucx2Dr2THtbHQhz//Z2NXqiuw68NL4DN2tXlIaIc0VONxX/sW0aG4DOy2bRgE
YhtErKI0URFfL5cvh4S+8ABsBNlSE2HAuQx/BExY5DtG3WJuS/0Mv5jGdQqOuJua53htr6GuhI/U
OZ//Z9iufKm8mtO7AchE36+IM+KUOJWTf68+AwboClVOm5XR+J88qMFsCavV6Y17JE8CqfVAhRCx
fNCxp7v/vDzLz6wjmlrOVMXGe9S2RTDNLFiPS/DOr/u7aSov4yNrIXR0LgV8QnZwSlPl1BZ6vVif
ZPOcyzUP6DDCIiYC1AwfHU+0BDw9Xg66SOiMY1qMmRdrR0wVPUr3y8YRPpy8Ep1BSvJCzLNCHStN
ClrRVKyAIGIyzNUPyk3Jj5W2yVfhm5kiUt46tXKU3fcPMQfmoUDCh6qDqcTn57DB6dx4jKLdPbMA
Za8JiAiRfg+uyt8hKzrX0aDUgnjPiMxUL4hGHWYFu5hBpH1QWJ83sroOXi3ORXEvn5usmjU/7Q+C
xC08gVuNXCv0B6VGv4X36z52A7tiVDuCud680LZ65oVPgy3nN3XizTnfl4IWn+e/9rDVFtp3Toch
aA2wq+nStCxgnDyMVaf0Rv+l5IogqbFfHNFN86BCzOuuZhOXGDmRqrqgM20zv4kdY8gCuxwLJUoe
CNm3Z2X3cFr6V9v8rW0M5H3PEMUKxc8UaHtf697DQz+65OStBgJRFzu+sRv6NrPM5Mp8C8pTC32x
YdV2+pGo1H4BMko6WY8eTyVecQXiAK9kzIqIeQ9RGq5dwS9gMiE201+WJn7YfaHoNScDE9pK028M
jv/NJ0yxMkhPCsQ7c389GCM/ZlNmL3gzqwyji+b2OeWG4ob5f/Vj+nu3eWwaTwV9OuTM5s6PU5yZ
Euqdl4CxdLTSGwovyzacdMGSxc33QqVm6+PKGyMLTOW4+ZL+X77xsInoVGhbCvPthR2LP19UTmy1
U5RBoVPeTUEAQGtMBqYTREN3ohOPKmHahLJdQFZjPaOvbltYysvuKWwSU7isGq7BWtZNddVypZoz
9rpPHItSkq9hep5y5knsuJ3d7KD4Ws07HKJEJMbminCzfupPAImPUdBZcerfU4AKFwZLVOKKiMZD
8nJ9qG++T/nckZXWmldROVU61y/rP+RSSSfcGePDkW6iVSL4BMVgGtzZP/Z9vsokLBgCRL6F04GQ
yEoS7OteMn8eK26+0aKESqBOCAzuhsw8Io7PFowm4CAscl6wDtzzrYDfuwiFzrFE8dTk7klJSYJY
ups83BQ7x6Ru4cdl72gpDcrC0/8WAc/cJNbEat26JXZIYx8Pm+mDu+ZxKLFj4sgyswqS0bWBi5VD
CWMtd2zeG9KplYa7g+Lzl9x3GAGdQBxslTiuYc84Wqxw3z7joajK3O4uKub2CT79zcvE7jy/AUz6
sRe7rIMcz8xl52m+Nq0mblqQdc8091OgpDxRjec0Z0fhmiXkBLEMlqn/ZkAfvk73W93Z1ADf+TQq
ZgJU6aTCP7PLpXPu9TukMJN7ueKiWYdWMLi+p87Hfe5Q0lMwvbaki52mmfE8CsNKndKuGUKYsdyR
3goPfyTT29ic64ytfxa/o7Rh6oPIZcgFT6QU7c5X75qW3fe5zol7lvkW4qWjq+AMRfcbbIvlqpXr
4TCooe4anhjHHvQouaWgCdaklui770jWI3qvUq4g/51Cb9RyG3WSibwP1LaG4et2KIaHKSiSdbSf
oGGkAGtHmQuO4jlasI/sxF42NVAzJ32EPvxpmk/u+n3t/1olmJ5lVMEEGPro3GRIyww/DmEs+XK2
Uvn3G2Djq8RVGMiLRfB3e9BTIpEoZ2OCgpalYl16YqWe6cgjH4ItZwze0BVvUwCr+uQW9nN2rFA+
ClXafFAmBHRNIfB4ewqFHXiGhocYw3n71zxBBVox1SHgABw9mRqPnZhEKkTOGcritlVSKzOs93Mg
NKqsf6qrfFjZOWA6jnLFKRmz3rIft9dP+UluEkfK9qur3O6eoBXXWQSaKJpZVkj7eQY7vRAdxJCw
jJcdprtKclspOuese5oRvqYOKCC9GGzEmZQyUGIRMrnrrYSxzQ/MBUj18RdpsvDfIwNhfI5dcwck
e6KTqYDegzSNu1Q2bFMzYCwT/PqEr8iVZ2Am6U1r1D6Iw3CmDPOtr+I3BLvMzV8VE/B85j2YFjRj
s0H2mWCHEDVQtY15wFGKWNxU43DIOm6mKCkNMSvSwpF11hz77dIgVFPgErG5OUOAlIpkxj28LFSK
sJmV0euB/jZDkkaZo2gAuTKv35mQdHiizKJHA1wuTdNr5kA85/RwXRsUGnBPIQ0+FGETJseJxRnj
h5m3DLjciX5tTDjaBEYwO0pwNb8X9iKaphxO6H8k8PBPvSTg5bal5doo1so2192QHgQZu9AZPm3p
t4U14T6hNWQFeCE0aedKwrTlOyVhjiUK5hd339rmhUebcwmckk/hJtSq+U9Fwb54xLqipKU+neqv
7Bs6XdHe/lHuwGNSO4NeUQo5w6L85rvcL9A7SLnORMtQCZ/0xiAs4k3iz/b01X3iGsWaT4o6iD9a
e6IEtwKk4vD3wnOdJijwPIIDFIpUqPv8nY8ee3b3c20lNB10LMXs/tLiAymeXf3D9azVtqQon7gL
Oz0YUJ+mpMqaonKiYSHV3yJiXy7pVZAh0Y/ggYhSwQ78g5TVRiQloks+7lvAhdERuaYNTc6jNX0B
zp9ZpDnwRjKHJ0d/UIB+tuh45vfRz05qy9pepylRxrW5LiTozsP4esYvqsa7UkBN3XmGp3DhUuZP
2VUnCUJmK/pFxZ0D0uvmBV0bF//PlNt9X/j+mJ+GB9pTOWZ6A7iR4TwuEO4v36myVe80rzpPco0A
rFJqTHF8zcwe2JHXK95Ck23DXOOm4KTONGasPLopjL3EDc/5Ui8sIiREXtyco5C0/+oNp5IwHDVA
LcgWfOt3Uld4XqAoBr/Y8UwYVLRrOCe9/ra+cHqaRNeE306lvRstaeR6pf/ikamDf6yYCSmVZzWb
kYqzOVI3gGFcLYnMA35YIm06KlcQAmm2XYFxOemvnLt0Px74wOnmlKQMDx5cwFL3GBBJOSdetCSQ
+l4nltE7aJvqQJ+JxQzKAzcPDH9MZmNhl+NtUZuOpPvUFu5y780GuekDGt2MXoxOZDUX1Xq5E7jp
2tcMEDv4uDZEVhoMKTjlsmZUJoEUADpVc/UlHcqoHAdgz5xwrMXCWP+UW7RDtHKBF4KGUyxx9cVt
IvFPDtyTzZg6/ipuYRL6/vaSS0dQgRIXdfU2jmO3HUn2Wi5R1Y82U0mGo4aKqNAJTO5vM5wZ9dR0
fiCc34blFykS8i6o9zs90DXrUTXhdPR1c72F1+PedglUmVFldrOPSdfIa5k7SkavpCZvP4I/i2uT
O0e4YCqArlv7G0yRDfdwLG1xvWmddQXeGP3vTf3liVjMFs7WfiylFZMCEvXcqK/m8LCUZFeHkFch
S/eeKCDgZ6F/Mx98i4ieIujHGN5eGyIdnYKT/RSQp5I+r5vFeKU913BcLj6MvVSqx1vfFRZjEhrz
Pf3KUys2xNLMSL81Q7j5CLfVqQEaWptotNJjxk+jLeMpBWS1xLhm7r2SX8JqAIy6fz/LRkzZRlFE
r/zNXrTGFcK5AXjBbrHgMSRvvXl+fgFAjd5UdDIqdqtjEK5OfwmUmGXgqEjrlK+d5uQ00GiPdHvK
3iFw7BPHpt9ntbTDMdWtC/pUR6oG9lU7ZAgc0JVbiBSI2REptURKFkYzBPpoc2vFl3U4QnBCAJrU
lGTbcm19GM4rPp2WRxdgGR8/umyNxPnVKIiB6caNaw8TVB5liU6Ifz/6NO98tp75IB8bL5dqGrVE
lxFu9G/TAj3yUUPKOsNlO7Ay9TE+Cdf3/rmvuAIoak1kOMuoDb+LpRC79mjI0QJ0wltYWg9uB3YC
Xq5iyrTJuikL6KB2UFm9JRnjutqQ+rwWOofR2Y3jMD1qkxswjEsB11GCvLLf47OPKZPB6w+66NyB
B2CkLID/Op6cNdQ9YAFuZuDoCrr1IwOCXD7Fvn10Zbx1CRnldpaMSQHKN+39uk8YI2aPo0nCh2ou
rj3iM16jL1ytoSJFNZdoxh6brWL/+n2WSxUmanahyHH5ocDy5lv/HBoSceJHSFZ2xmoBemPc2WAH
zcCmIz5j041UV8xwsp5n9rrax2AaH774bsrPIxjYsIm83hYOTz9BqzlMRAd3enBK453uGaThHi8K
UpQ9k1oyQRiO0U5zXyknEOhg3wmWh9gyf7153EnroAZk7euIFS6IMFmn5o4Trd4pdf5seprxrSIA
XJJmT2XhbhvLyITP1/ABZ8gtAGXwxoGm/QezOtaRGnlsQHuMMrz1hNC7WaJQX4etbS5uFNGi6F4A
1EBzCVzylMLBBOfiYVr4CwM1ltC9U2ULRNfT9wkI+UQDBEoMcffmqGz60rFg0kr75jxen4YcjLa1
MaGuSdzEo3UXTAmVi1GYn44KFmOhbMmCr5YkKPdFUJj0ycTawubaafGfbHAxGVEfl9YB/kdcphSL
RWDAUzbG0dr6QDHNPVby20gb9tKzH1Gsl1a3kTlUEv/1Qg8fR591C1AMUMhVVYtfCBEEIXSK/P6K
2vWf9wHkPfl790mVTmRX+svhLm+30f3wt1CLe6tQA1uixitWUqBQ8tnB6OQG/wal3v+4UzcoII0g
FOY/6rOFmrR0i/OsNotOxLxPS4axPEF1NbboDOa0OA9Ye2onRMFdY0mcBbsyxOc0EHyrfSpokpVo
S3HxAmspv3537A0JbTP2WkNVR/20Eo3lCD7rQSgiaWMvfNDw6xLX1Mquf05orqmEgt6QPJguGPhF
rhtT11SiqCiMynh9uIYeWOmPXHA0PrrzJ2u+L82JS9EfLhZVPu2ecq5dmL5Pv4tpftRoinqGMz61
wRBl22hCdIZG9yKbxMbhkc71OcU8sLnIg/JRQinFPXfduPnko6+u8IQ49UpkHqWSOuWVWq94ZLd/
uIdUCtmNtO9b9eeu9u8II9/VO4n06MYFRP7U4Z/odmC25IffLHJYARA4yYtHGrzILx+fM5V26Iii
DPj0DWD4hibKkslUvVHgEIZkq8VEh1SUBXYF4hpCy2Qh4rJh/5CUgM9keSdyYM+mPJci/a2cIcrP
0+itTSUYj9ieRmK8GqWVHP4i0Vt+JdyQzHPX+imDvklK9gLn7cL2yTT6FsE2X64em9gT1pVDBT4i
wcvoeKYtMsnOlNp1dNNZ710zE2q+4lde74aa5whnflnv9CeidNBv3m3UXUD0oqpcOgukS7F3VbfJ
XFXA4MtE2cO7OEmp2hEvnw0qXGr295y4zYAuUlI1YmcIeYeOuAWpf4NxSW+3jTMDAMD4NPmwu2Ac
T4/+FNjS9vk27WYy5haR3TF5qMbEqVHaxoDXkWhjr+/56L3EqG9vE6EMjKmVV9zaFfvTNE5FR/WO
YwlhmQowABEjbOOSQvYtsnRZDwX28RCkQtzu6eEImEGgqTw+/W8zBGlG/CQHpzqALvYSQ6RYiplm
pqiwMUjA3HrdTJUY4D0sXai522qM6NxzG+94T26MTo6h4arxsJ3XsATdxKpMsqIr1LxHL+h1d4P5
5+9AYrrS5uWwQTSL+THBP8bADCLjugOyA6HjxzLvFEoTZ9hObA5cHfsSFxR9GsLURPzNAQaRVUCj
atwYvjEyGaCoaLKllyXXQdxQQleqCgeSSSxfo1+dF30ggMIQbPdJHocQR7wlc09m28H47icjfdn+
cCv4RruKriVsQV293mLl74Nb5KzOXFkoM9K9UOuGWmWOJXy9fpo+F0yP/3uXtZbfFrDRx2GLirBS
LX8/LjCZVWWqWwD7rJOtpFCby5ShAvmPn3/jmMq/aPyL9zi7/6uWScKQGYkB0XZofQ8jtzVihCXV
0lWn7XaubMAwTbheF2BEtCDHSjfuLGdErXdXp0o85H/av/i3zPtc5fX3ANSlYnp5ybrH4Q3cj9z3
8um04wYQgNE12km7z/oboNwtQOWe7LnDEj66tIdLlV4/tHx3Ix+ihTICq6JwOmHkyaIqyk3qc/hg
AupxhwIqqjOiltP+TiWMN9TImiiKMa40neZTAXl/WRfYiDy89dELnara4ld+tY5Up1bEVc7YJumZ
Y553tDWiAo1lh6hHCPEQ7/+njHSmPAbQR+zkFuUl7sFikjaySWj5CzO2peLB8U+cVLLJJepQcE74
gpBQAdgrXeGtT3G/JDp7727HS6N6HbUD451s/VtQXm/kd6RsaNJzRD1AGuq6lGjNObBBJsBi4iCS
PZ4IbE1xCYUxF57xNEAop/4QVapAoPfwSBKa//V4ihpzRbrJrfjfbv/7l+GylDm8PfzYmKHn4lUE
gBVN3Fevcg4v4FBQojjPeueSp+daM9hK7FQSP0bhcYs7Ilu2GsTr3RFj1g/2O0BQufkbIYzGr1RC
MAhA7NGcBWMYIzVfjsCPbilLpiWLEB16JfYT30dTzb4C+IqO673DkiCcOnVHuwyq9yRdjOK5AMw9
59pZw2wh5SJUQumFheC8FVhqyjX+JiRwWYgbkmleV3694UByAWQTfEqas2fsqSht2RrLrMzsGrxi
s3yIg6/YRgL68ld9T+iPq+EURqJkxQ4Yrg1R5uHMfBT5OBBlU9lpmIjYv/ohm2wnb2zzmQgZshcs
DbCC7MnU6EghAkxPKZldLsnelYQHgDBUjXdHbfscjSbZHVo/xQd9nVANIGmuuniv1KmzbS9e3Ypk
CbCSzWM3KJc8ItGXjXKyxyG7UsBhdlMybBEaK467fR4UCYVAOFSnVbtPIOnSdZl8UijdAI3AIf6V
wnupPlqPeIAVb2smQa/q4iH3JK8ylsY3wHnIJWAxdl3ZosDDsXv11Zq+janeo9lNOk5eFBPIH6lK
9TQMX4YjvOYP3QhXJiawalANe5juzJS4/lphiz/gpW0XIcvcY+/PAkUtV/NO5PIhBLa97zMRYZjm
gKq3MiXIZ2kF+qzetkrS82eX60AloG2xvYZG4I3Li7ZflngG6dqXkTBj4va3LdthDjHdONWiBXhW
NDEcuU8bzfGIRRI+GmsionRn48zj6SvOl5N+NZ0BQYiqs9GKrIUydd8eXab9eSwQ1itqnLdJcBWs
kPC0AOo2tZRdxqA0XfW2boFy0tm8p9YFi3RlZrRQSL/DqXTCQ/BNky79OneFnWzKMq+2uPBqoiCE
BGF60bUXfH5e8mBhdeTHD1jQnr0o7qAk05AIOFe/BmHcxkqYJGd59OuBacT3volCUnug+HX332u5
auLdiWPRdiaqgwAx+T2jWk6G0p8Czr0i9/CFlgjaYQFd+QNB8EdL71TZWZPSH+R3zu81ILDuHDBX
JGVvGeO3QQm4eh1EVQ1RzcPz8lVx6LIy+/XYSUkg7KtNL4ahuu5VKND1QHZtL1oih2l9/Ha3P+ms
YZigOB5ide186+wwgL/nFeFLZ7TKT1zBHh6ZnwapJSEuTEliPtvXJ6vP5CSE3NieVwYbxH1/EZ+V
JQY7eZd7zcIZuAmZlMVRqENxXowz5mX10AwAEeel64jwWF+9xp2FaZqTi9h4OcnLvqKzTCpNYWaq
hpjocPY0ECaY7qfdNS1zXRuTs7sle1/hHtQ8A402p9/UfGzcR36488xq+BFcc5jxLoxh9N4O1KME
sToXiuIzAIrhThA5GnpOSzcmVRc5jnf7orUqVLp1C64Cspqbvmln8PkkXNtWInX4yfVtcKEDnj6K
MgpgZmjFWHKEFbHvAyLb7BPHyhtYY7bNBe22DyAvBIbmuvWn1x0FTBmMurQIkY9mIgHH6uAb5HxX
DNR2mSYjke+kTDmUUb0jbEXSC22ocD4LJNjUS2PP/gc7CaS63g5z5LoNf0PqZPpzitPHHv6Fvbbo
M/ogBoLMyp1+An1fi05OHDrDtjuiTwjX2yot/7GpwEhgrPKWgSafo59D1Syq5dVToVfqQhMCX53q
x7mXGgI729svoNG9qksuHAjiQ7cL6zXc3t/bw3pU7mrTMz0YrIN/lwdOALUCHUTo7Bjjufky24Xd
UEZ4aSmFmd0RuJTlQQqLrD9drkPlUiMgSRQ5hSWZoWxPUC8Hsyz+ulvI4Z1AD8XeU6/pB3NybRqW
if/nxH9QTKv610xV7nL1kM3OPxBza37WX0mfL2ik0IN1Me7KG89Tc496EjuuGOftgKRqsHEv9J30
VoFl8JlM+peNjgeNKtFWm0aARAvcGk5lwDljOEN47ES40igRd8QepsXOeTqMAXlyTLkHncrIBXps
4B6R0xbvocf12b+gYNTdmMLsMelhUnockbAM14C7e0NNWiuJ+UTlJGfARTDCdfIZA4OVB5cwhWKN
XVqvmvfYLtR0ZZ1tVi/3tIVAYZ+yiqyDyXYD30aSKX7u2kaUZVnsyWsTIoWgYaYAzcTLWkhYbCDb
M1IelrM3774tZ9qhtwIGrsC0+Ai9l0RlzYUsgROrIvI5w1PGK6R5ZF6BOc+rPVOwSrDwViJNjVus
moqKMSjwU+G021zjEASaZv3AeSU2G1Ns6cPWv6PKl6GqVI1ABsVipX26ateupO0vnWTHOlGsvdwR
U1qMSX0geheEa9MPlGUu4EXF/xQ1nLArD+wTxrKPH0TGpYs4lx7lPxQCnOtvawBEno+aHRwxk7Mx
aWvhsuYfLRVhcSul9VNyqhfAD5iL3oi5PBWjteG8tj5eqEWAJwPXizC4pr3M59cwhwQsnVvc6zH/
luq2Q5L3vAXYO/rqVzTKEu8h3yEm6HpQ3SD2rJ2VFivVVVeFxd9oImDsSomRX/6hqQzTBVfLXoQ5
Rsv0NJY7ODyo7mWagw1K+R6kue5hqRu228RfKQ/MiVuyWBjDnzEXLGu9Yub3AImDRxP0nABHSVGt
LeJgvV0UTJgtPasTvMSk4ZMOBlSPMmUGv5yc7y4GBl1uFSIAX/rV8TybGbfZ50sCLGbQRMQUnXV1
qPerzemldWTOs19pZk+os+Ng+pD1jFYCFEOdB5BCnkfEZ8HTVnEv1a+pI8DyJvkvMgESKX10/xAp
HVXFrb6XmDAjDeogQpfiYgguQmOWdIG173LkT10m7DgcPOfxAqKCJ+N6lykCaXIk1f+Z+JGsy3ir
4mLZnLFKguwZoL8Vjunl15ESE7GzoPevWFOVG7IOigX777GX6bhQ8BgTgh+BF2A/5HrIsYgvOMAV
tjjV3y7GNJL3a0zDCF5M9deDQXBPnqWvSeg2Mnwdk6S1T8eMhIO+2kgQ4cMSZ4QtWbk2cC/YlopL
qCYqoMtFvYJOVbPRLifdPxZUipTASyyCH+N2An6ZYssfUx3hmgeGG0AXu45VnlPc3lIUNwhSdJ3M
c0EPVfpzan7Af+4HH88I5T2w/yQ7bxU/bGI2cNdakfmu5+i5ga5/HsaJ85Um7TRQ8UXo0ax+VfpI
BS6CxMrFnj3/Ur/bRzBwRn5HQh6bHweZ106baGJljwTa1zqL/DNzcZftHX/UbdwfTefpy76rwJog
QTMCDgMOTR6CjhGcAoWvfsoMgUX8C5loQb0tk30SJ/OwyvV/FRaJYF5wLJ5/fteRA/mN4M2+sAa7
1GzXCE69HNBcWO3oo8/YLaR+gxk20OVqFIKJ04SuVmc9RQewi1dMGm1SJJTH6Sk0Qc+19EYbmaN3
REa6MBO/g70uZ0c9KlKf/N3B2vaSJWsRvRWQ3FIAO7s2cbnjO4/vrCnIhE+hfeyqAOOfTf/UgFAP
7tTd0DbgaNCkWtHO7Uu/4dPObPBMfmtZGte4HtgXFPlYrGtKFwH0hWEqex2pwxqQzLPPORSHA0FF
JU3GqCPiepIEVMrShNUe02NC/lIHK7rgCTtD1Hz2qdmjy+ICFxCzlJlaXstMU4zODWnNIy8VO4Yv
yx36z464LclkPDBZv4BIRDE7Phj1osgonWLwYgZvzFAgXFYyAWL8tM5vbjz4y3po6HiJn0nWS5fC
nAj7feNgWksibwiI/VFTdHwuDvuScABcKs5AxOvz1L8m5hza//zUUEFvxa+QmTQoDMQyao+d8Cbm
xLLpDblNFjUJkB+eWlFSOjdOx5hx3rvLVIjqpujwkzTX8qdqIjmwKmI98llsOtPgjZc0V5V3ROcE
ziIL+DVojH1iPKmmxw0NRDdm3Fb4qsmNTgOZU0a2cRHUHT8TCaLSodJ4Zuo+Uk/dOdN3A9b3ULze
BOI3MvYj50EI/3rcjGnC7L1rDgK7BKcSFwyqy2+dmECb0StfyfXAHyr5o4zEDDOZr5AtBnSPHS4g
EjS4Ed6+P2GWOh/gbur2TS/2qG8ZucH1+VDtb1o19bFnp7bghguaihPXY0ZyZVHCm8M7U60e6Pze
3Gz79oTxNTaAx8T5Al+k3geXMJ/Von4jpB7B+yIChFp+4EXyBAT0DWVnlPFW5Er8qf8FPUMr6+g5
ozdRjJ8koR+Kay/Sc4W9ytSAd7Ke5oUof1hBWMW8djsxWrMJY04UlfBzJPRRZn4MP8ImPMo/0uE3
gVmPU38mXJQO1XP1BmigtZql7oaRtkE8VpwilOoCdmDG37qAon1rimC/MF+NjKjgYMvwgm6G7Fxg
1EEC5Zk7hXRs5OPLZ99SYfR7yLqgHlhY0iLFikhWE92R1kuKx2RwjauCTzowrlCUr9hdyybnowDG
O6RnOIr07DYO/v43t942Sai/n5hkLMjeYn+JAcV7FbULThuqVUZ59bZEpIyE0AT48dclBELTcfO2
J5sN1oBVIsjgKI4lJPRUTHL/8zsKsAgq/jv2n/w0q+LVlaLssoJPuojcirFHayuAyBR4uqBLRi/D
Vke+Lpxv0m3+g3+B7za4VtfblbZ8PsjydfKFEyrQA+aEVtge5hz9BdDB8mAl1wMVOgoTkomWCFO8
n33wLCw6yGZGJqfbHXwJak8+rvOAz71J7LYJoBgcSwOlsiUHOJ+yW16ex4gJfxu8yZUa3Nz6cST1
bwZMlueMx+Tf5zcWsDk/vhZnQjBMFtoxNfWhRJoF5kl1ZjLB+Eug1fdKm3nmpMYhM0ARbacAnNI3
LaLZJGfYsurVFqWq8zJ4oBymlnRVJluVNb219+I5UbAV9v5sJ3BzVY8bcDP4rzz8IAFA7kqRmssJ
H3t0ipLII1V+PVlE+Awklwef+wEeYEKBwIj8I2frIqokA5XpsHhDcCbrEKD5fGb3ONk3zvNhVZvu
uTuanpbB/tK/IRK8oqsauw3T5bbXfvJW77ALc5D2VutJEoYO0t4eHenpR8TZfKsChXfwdmn5oe37
v5S02rn5+lmehSaiRN9WRij8KfotQNK3ic2s8xavvSjM7H6ZEq0qfFdRL197PP0EejN0xMdh+Gcz
74MUL1wXAzlqh/mQ1T05lNpaGCfx//Hfp5n0bYhpWm8nJp/hX/9VsnUdyShJ0i2jC9Z65Hr3Gtrw
jORqEZ7Gf74z5NfkVFwww3Q8TJ2QTrdRUDSzbrzjUkS5Wj/molyJUJJF8CgjvcteZSgIwb19XPeh
m7ix4+qM8r3+F0/wFsy5pcSrBNlO+UiyzWbBJv47/Sd4aNquaJLsV75Kp1P4ULwH5As8KDpS6X32
At4rFyq3h7Kmct3F3vWFR3WAKuVzjgZ9aJ0Pz1MMdQ+DEiPLcvrkKcaRo9fOxkRsqb8fTD+5faQy
CetuD5rrmB+xHbpxX2VQsMTslAyNr0l0MPLsWm3YkKKPB2s3rqa54a25G85m2c40kX+Deeb7Z6+x
+/3H6x+TAYdP+0j+aPW3TsYf8lOtEHPZnRClgS2mzHDNGqCsgnY1hSKhWGWCqrrl/Q52tPtc2bOd
32jFD8rki+eC/cmR6z+r78ANpv8NoNtZzH/GFoOuTEUaGDsqs8uzZdJp9N3Z3Sz9ftG5dU6zRjC4
iJRdHHsNJwrIa1PvAwO1qG0PYZ+8xSOr8qtWejh5hFUg/WoVeALjurDLVxqzdYys6VnWiLp1KdT7
O2osNjoWl/X97ttCk2XJMb1KHZ6NHhfc1vDtQjmVUFth8Js5EHCIWhT9YHq3JF5UynWKeuTCGvWp
OIpL3U9YivU9xhvHEq0JlTD2lRtKYuQLMEPV5MIC0c95+r8T87VKK6I5M4+VZlfALoYsWgpRAEcw
cw4oAJleMDh9QwyYNSNPQSSEky7lm0V9X0fCC4giJPDnaTrUEpQd9gTnYNZ5rNFkNmG04owbY6Ry
BMpK1zC2dFQN9eZjsGvuS5ZWOXaoiRvEuEVeOq0QzvJML7cFAF1aJ9B1eO+OlwfDR4A0iKRwLCTJ
670y7yXCxXnfDD7vlgYuqy2jnSHEli8vuY5L4kG3mGH8Ku0m8LFZNiCPqoW8TLdihJ1WIB7ycDp7
HPcgFn6HQnF2LFMkA2XQDn3TZP9OZ9xDpy4RrnEXXssi8QqLSUxS4gW+1NXB9L7q7EXdSnS8UrBl
d5qds9sNi3xSFNdae9oEao5jQ1TcUgG2ad+Azk5/hvt3hP5T8qmBfNJML5RuyIs/VOfKlxWN6pDu
5soEOWMzHIxWmsZc+2Z1RPyoAqxfW6Q21zu7tIrpVebg4wSpTMILmTXv/JKK/9D1TWABpPF0DGXc
UAKmqtPFJoKXY90pGY/LKGES/p9WrC2FWiG8lJAQCtZCBHm7vpvnVaD0U6VkUtSf+AHxQd9q9Lt1
KiVb6EbdcCOAtAc01yG6mA5EM8v4J5kEAmoKrvbSZzBT8P3ii/JQ9WKd4Q+DrS/9LmM9dyOVz3+m
nXvAZy3Af83BIL5ckK8u0FwZYBlvKOkVh+iWtFv6O/4LyKDu6SezxddDq+2OvbBIk2B+1Fd3UEys
QM4wLS4x6EygDO8ZjokWvukQVZvRS75mbJJtEi5UaAV47jdlYSrEdi7d4lIL45JmWNNHtb3Xd/p4
vjITIhEnMOzetVfKCX6TPOgnRTveQ/9+aIK0Pq70iDXFVcFrs4mb37DGgvJgZkoze8kxvzkWqSEt
q3XyLJIqp4P8ouI81/xH6QdIv2NxsWZTL7LQDGO3z7Zl34hJPvUB0qE4WzmkI9d0NzLJjvkm0DHZ
7QHaEcHC7aeEZtMP0o7wDzz8tr9a0JevBdZwGy2P91zBct7d0m+oL8v/HRHGEcNRInptbXiEy7UJ
ZrY+zruY3PkJ1EaW4C9n644CHipXwBvrHUFYeYI7qIMnhrHervgT2oZH42wfeJRAUpwI7cTy9+fj
6weypE2WjZC7Ov8jrcH9nmq1kWHt+rrdLgv97E/oHWRA6pgZTjJAOEFja4jgFpkgWDxMQzWKNMGR
WOrt4uwSqvkup3A/sCe1eXINCZJmeT0VyTdnx3A+bZsiJpBqOcm4DcCBvU7yuEy1paMKTiF/05mt
88/rqEm+kTXa6SgNcLL+ihRtkYcGVT75MPghUsji8H4HRgcAxcBDCU3IWr3p6F1k9GGPdao/cky/
qt2kYDx7xae5O9lBCDgwxG+YubRgeL/rwY2Z3Lt/SJKD26VtVNCHcYueOcaZWCSEuhDJ1lrx+RAv
UTVmKamN/vlxbyvl0VEhcY3zC7/E7Mrcu41CkvWeaptP/WSXL/QxR7iw3FWpEXBBivh7ksZlaKwJ
KmTo2HefONWQ0I39zi+UB+TMbZbue1/z0cfzwmI8dJB+shY3EsppmitHFjbqSzhf1KF22eztplpW
RJVtsYJBt1aQexAdDs2MwRiUf1+hzzPqrwWdH21wJTaTuGfHLmZhmTltZ4LP0ljoRlH/xnyEpVTh
49Ad84k2A3vnIsXyxVM4Mbg0xRLiuaM/DOXFk4Y/hc4jTe9FcVeeypK3qhEpU/q6M+9jaD7Jtj0r
T8RdKtu2Gwb8k8VNpa1Gw6LsnFwymjoCkobNnLgoLMEdUoawCB55RX+MFsOENaa7XkdjO0+zO1kT
0xOncUW3oc2RsC5Nw2RJcvU1ahzjNpzTn/Iqa/b2+TyVxBGxSGPdEeDgunHBqG5qLiA+T4vidfpD
AV+yoVpcQOS+/FijXvYYuuD2O8JTpd+A9Bopf5cceuXKTRY+cf/HGQYwNdA1B5+Y2P1J4WA5DPTH
B1W909nZ4xwN2OmUpS2ZIxGhfbFKToVtu5COFiwNaqzg0M+MPKkaRidmvXjJ3ob3JnT6XKbU5aV7
X4MTJDUMLSCr1WEuDO/LcBSwRueqnQzJel1QQriwHmIy0Y6SzgEthmkhjC4jDakoFEUmeegtgv3c
NScCvxV/8JSIYMnj11TzTOoVGJjpzvqaqRCQzOLXBxJZHPEn/ho9194CH4I3UDdGb63rVkfqfJ0k
tPT90fNUyTShzk3MYvmEN2AJ75uhbPvQMz8Jgk0uE3hYbh16q/+UwDza7Mv/RC1ChXwozgoayGex
m+sc4Spy8w70cvHHFvehPAw/+NC2IuvcE2+w6FVCA/oiscjJIgebFwv6L47pHSeie8aO2ldBEdcE
VX8H+zHz5pm1GHC0fvBRJIRdaottz0HMvCIumeFW7l7YFKaY8N8yhcEB5mWEUYrEr6rqCqX/zqQQ
TTT7dvgHqgMtZv0eLCPyzVsfFDjCnDHALa50tG1qi8m7JjbKJwrHYtBtbJFxrENsejcCzHeib9Bs
EYvCW1KuVBrcG61khdj32AZXzjX2p+biMbsWkk+htiBck+DocgivWn6dwj9ef0TgV/JYXqkSpPCX
2JlObKw0YvX6akCbTeCHPF0VoILyxrwUfVh+oTMmvLBUsybqfAArSYUq7HVY9B1u/KKjgyKpSBF6
D0v3ay8wQu3t+AaezBkbrxs71vMEorfyNmunBOzR29feDdU4BJyQ+4JlmCCvsMyPaL2VLvbseM/O
UJHS9yJyPB2FBgpayqt40rBsrUNzOIseqTB+ywXBbXWpIDor4i0MtXvu/XNZD9lVMGnSBui6jVg9
jgeiN1W0eZj2xeIi7mEtR/k/2dm+IFfpxyYBY2ikr87UrSEVXdiSlO3+mwAqKslTeSklNF4X2q5N
Ls8gP6TcxEUh6ytiGYqPFGmIwJUCwIn7DEfkMbCztDCeZuVFo//W6s7SNJ211sHvxsz8QqZI8CKa
gCMzjT9HOlPLKxLy5hQk6oRw8gryDkr1nJE+8baChY96sCzW6w0cB5eCqW59jGjbQhZbd22eqLY/
l6y/6vZ+BBWVaHb8FVF4YmM556lbYW0HHXUxGsaFhGfAABedu/Pq5eF8iae8XL02BNrZcl67y4Wg
OaDJ1E/5PDz+vZr67NMkBamF8EHRBa8AhEdwtgTNjnLwPx5YtzhNhgwGtssaHrz+TzomM6ZmwFQE
PO9i5MPtTW8lS2j03BiPoKA0RXjSGnkR7rO/rT3+Dz/Ruk+0XwAvXMWQkEEV3T4JLVfLbY8S9j0I
CijiCuvQzM4LPsHihSrAlRXUPHA0QJhwEFb40mBsfuGHuVE4fJs9i6GqXmlcxET1WjJ7ifptimWl
2KVsVYmNQsYgdR9sVjF9jCzSe2T0arCSXqbLCfSDhPixPTxx1z4TQCQioS3Eqkw//oW01d2EFkY3
0NwU0sTIDS4PKA4UtC/6gLqCkPUdXRsQsiGqRYaHVhfSuc+gV8MwbOZpxo9jFnd6IW97JU5E5/p2
ABMKQwrRw2IJ8xBTJiczU0cZ3dqqlbE2VNHrlXVrLY6TVdj0gp3EoHh0sQjyBL1H+7qRZ1rMOrZP
5YrZpEgrQx3RplIH3mIloMPP8oEvEGp5L2N3eJZvr6tegQaq99oWoV5ALbwW3O7Fh4Fup5rNEjck
M3uljWluBQ3sxFBCccquz4WtXxeIhD9xc7bMcTXYnT+6RJ65hL7e8xJCKhfAQT4uHZm0Vjh5iZBx
eUVbK0rB6q/ktWpNmrfMMQ8ZG5PCgZLbXEYm0JqZ4tFQX2Ucgh0bTtGYqpz6mtr6RI560a9RkeHF
otFZh6tH2zZhsF1laUY0ug8ebeQJ0/UGIT3BRvCkT/ekHLHj2VDZyeHk/eV9QDjdNGShvCmennJO
tGPraSGdN5UzfZ8e++Mq1ouBw2A6FX6Dv8rX0XjgxU9xbp1OXckJK3f2ed7L2h5wdXO9MY2efcpO
4D28FRn0dNRwuag1cADv9NLK2dk2TbyuN3UaNTAwg/45Q1WvecKYIcjr3/4pkMMpY8Ym+uxNlN+D
uXzjs25/e8SP1usLCxDxugshQT+u8oghQLQEb0ah3jQOk3vPr79WznMdJ22YZHS0Yc0qDsACvWh+
sSg/qv7W3ek2+LcA3c/GqnY5hlpIOKUk6hBfNlFtdikXh9sOovV9KAzXJeOXzyPpTegZ9ZXbQOqU
Qq5eXfFYgx+qzk8oGPPxa/3cwY5zlrvLnD+emplKeHFgLl3R9X7UpZRk7FKBcb9/SLnXXnYjq3Jl
+bYoVBJHyqMJ/92s3FQrpduTHTE/q50oJlaJ0t6jaEo55RiLzn6SfVb9rKqBErO04TX3MSyyRWav
e9x4N2dyJ1iHm0uMTTlbcO6OXqqlOSowSNw5VGSfuA0Y+L8La59yGPaR8KzAQsJ83IZtPVc3uKvd
0xbS4HHkQsYgVbKsvQnx3GfhDmwpq0oLAgoE0LlSecbBi+SeJ8DSheWuo+sqQq3nvUw0NmP5LV08
VHSzq7YvqqcdFG+F+4cFvRpuaS+jPcWEKXzdjkbVEchqbdkLaAcOAsIo63/iAwE6ig4lHR14zK+n
Ray7lyddeyz6RSpEhzUGFYMbbQpmcEUR3+hWSPvPWH04GoR7lfFL9LSvtIVYtulGkCEny1LUC0FD
N7b+zYeLlNmZ7E347dMjD3XiXRhR/cNNpTXmw83XJQWP0OytC3T1FrCFg6xykiWhtxvwTWdVwnhX
1k5n6dgbTXcpp44JcTVNi/0ugvwGZZh9wy/nvKuMElsS5RO/KgeC0rmFHamhw/owWjsSKcLMEzeI
MWAiriDajtdCZhj+hNMapBGlPeEqGO+TXtwSOjY545XKr7Aocw9jWntDiD9tXHw6IywHL2mK04lf
+YxXjw4aa1WIkI2849w/vQTpnALy0+3micWlPeicaJHENHv6vMAUFiO9tG3tpEo75YqNuOIlLPOc
eVLJypez3/0lmCD+v4HTv1uNDZCWE9Hw64/g+NXhHcFnopFHO5jd381HGhCMiUiQmfXAaNYYMOPD
+/Q4Ic6DqG0clciaDU6DQvqImahrbNpaG90dyRU8yGSTxb2gEY7zTDP2dAAhPdxU7QJxmDRHxMMa
yWWnrZcCaFDL8UgS7tw+kcbpC4dWVgu9mNfEWFXJ20cLDQpQ73bhjtf/QQS6MR3iqLNhWE8JNQmF
6mGlSYSDct0u0Ip1bTOAVKxtPjhIK4cO9FaaOxvXFhC6lEYEuKBN1n/IQJ24066y0vXUhe39/pyc
HPkTa05wo9fDOHTc6zMxY570SIJgkL78y89umpJZZTdAWyb6QgWgsBH0JlGk9cSrMVGyWdX2luu7
QJs0iCulf5Wi0Dt74KDeasQdP7d+ZQyZUFbVrz+8M4EYF3YH7I4oM+s7CXPk9469eKimL23EPPGO
gtqh+Qu7YJSEoK95+FCqKHeTFYIfZ49+tSpc1Uj30X3fVPSUJyUp6uxCpcWkh2IYBKUr3apyMpDK
NpTTvwSGffgQXQ5Fo1QzCCAA/DvVT0uQ0vQhQKMuEFr33rpoUG/1Z59tmtp5oAy65mDhJJQMQFBN
2PniIzFbSzaYWYqkaJVe23EVFVX/QCHmVRszBa4u//51wNd7zcdsdewh1j/o2NzfZfFvq1rHrB9n
Q+TisPd8lpyAHc+K5ZnYpLvpgBsE1h4zMAdCH1jIcLMpsmGQdQxkkxG9vmGmeJnFW9NkY9a0QXkJ
n2o4V5AwXwuIswBvwVz84z+moGE37qhyVvk5Oyd5vzI5SCS+YLB3aguttadABCSGSh0IKUWNbeAF
CJy+FJ5Kl812Fmn4QaFu2otlTRTiMXY9w3KO49/fMYf+QSpLi2giOUL2Q2txhLgeZFRbZ6RR1t1b
fOweLg+yC4t3HDe5NYvMeKafkePH8oribJwJuYS6MrVkYOXeolDOEmrh9aB7wXSBJomTfMMjHq99
hR9F2YpL4C8CU53n0kOmcjvIl7At6hVI5lqjBb05d5WydjZ+pEDhe1l0Ovf1kfRa+ce5443wbhNY
Xi9d7sXmQyATiGq2RX7iJaurCETTlXhTZnuEioUZUefvsqtKdaBHBI1E60J/yPtE1MauypY6hPWB
3EtOdCzMI83t9VMYMsA5vKY8cyCIzj+pMtomvxCpfPh6FjteAJyGQvhzmeGkcuZE+GxQGv45lzwm
9qZ390zOPscNImfrMJv+QTC3445msc3xXQSKkFGlCEnNfggaJqw0zxGBp5InXg5IDiD0KgNKbfmt
j/QngW3kIegl/ceManWzw6K+9rlBNnQBOzACnrZHB93i32QzL4yf2Q27DDWmSY0Fw+U0ApKJlXMf
JkScxtNMd0KlrOD0mWvI+U3quRHiXEMZ8lrIKfiadck1rxSV+eGzNvCFio2MjvoFB2PwqRYc3eil
/Os+XzpoEP64T0ivcOEwKONcfRBtb4RbwNklXAAW8Pp9o4yz6Z8Id83R749Ey7l08ZHX9HlNOEyi
3Obb/LZlOOpqOr/ut5S10iyrhQbYBExS4W36H+t6zwmMReyc51s3XmsuNcBwD1keZykfUOOalbEa
KQ8rDEySyjbdQZssStggAZl6sWbUBCQvggE6pOCYKe1/P3/ZRd6VgORcZAt7N7QpWslchPLtzo3a
9NNRdUkvXKEs7Yya/nV/4GDzbNpzw+bys7y/iGSY9aSZWnxbCs7X+yPa3CpKFw0HzG/iMLuXpLlv
ZctZHSnzsVdfHmlP3D2jmuh4cuNuRL6UEhRNoh5wCeFr74rDErHueSiDRCecZox4r6Qq/aJQq3Xu
KqHDJMOh7AAFIGUTK0lUd2K12Qzf+3jZCxk7DxtWiv5pjFMSIdNGRzH60AlPvVoTRq67e98r5anT
ml0Vk/ooq7KeYt/ZV6qjpxkIOgIjBICAUj7bguYHepWo5ThJnP3utOQ+bwrx2WtMhk2Lyw5voFYH
DZGmVryWM3apg3hzaH4TxafQ2rKyF8/zsLQIVGQlwBwACiPxm00lTKiakKoqM4qPKXlxlTEm6zfq
qxEIclX5AO6GEGN4H1fKN2XFJ0Bbm0C2FUz1Qjjkd72eudzbzv7hmdqJygrbQCcC2RN9NSL6QA6d
5Mbp7fIwBaeW6LSKKphyXTwlw5m8j01LGEgEfWxDRscuvOE8hyx0TTZhLnXzkmVztqyUoYOhfJWR
vGC5Fk3qwtMVOzYHRjbGolOhpTNKthZNlHVkUAvVcY9phYLsQu9FItat784WgaclrbOKX+qMeKgl
YK8U2/pFcQkOWZ/yQCd13JfwZyDZ3HepWGbAmzoUFwLmsN6SyLxS+OX+S/cIdhhyRk5q8Pk5rUVv
OPMH30Ojp2aHzYNTmt/JDfhBSmZsRlLqXlXhIXmbdxym24+raB3PCoDTSXSefidM+/tM76j5yEaR
LSTkM831VeeukqgxQucosPiW+z4mVTZmxlRZnado1MLj4ViTDnntJApu+hYILOaFPlqVjY8g9EpH
/CMtkwtkoKZfhoK2BK4cDcb2I9k3wG+lP+nFM487dmj3el068yhu1HIY+PhxaMXl2NgoXJr+xZYj
DXl4tUQ1Zt90JrGeSs4B2/XEdipJ8aRVVho5AEuCyzfJmXOIZM7WENGr98eqvLRaOVSEJgTQjVaU
eKr8WLnh4Q86bJjgpGBBUMQn4AgZNJRNudNLtwywHTsZc2Olrex2Qm08voRc9ySSQK+4EVdyRzXC
bH6uQfnayum5e+pwedVrTymYv5O+HmO956yOqLrl17K4p3OEMsYKN8Sr/jI8zgwN7VyEJYbw2ga2
Ms7IqcbArjxPXxvHQZqR7bzU53u20B7Zh12mN7gr3WiYo6gRbLgX+ZY4sPWd3/7eBhlhWNMsHnDB
FK59UwuWhtaO/ecsyZNO14m33rJCVrR/MLyhnZMs+PnUgS36RlgVGLft+nZTWtJPU973CRCdqjFX
5A8VJTUytpECIh3cyh2L+CHWreLwjHg/zbKM1g3rmUDqExSarr3Z9HtI8T+dupJpej4MBCzW2UmL
O3QJ8DcQp2Epy5BAFFmwKW8oorlAsy/zXYDnPkbY/Pc/Eyl/Iczc/v76W9b8NAGh842PonGsOR+N
HSnaKk5dZJ22lGcAS/eonA/F7bts7IcDaa18NJ33DPwsGkpsf75z+FRZj+yza6QC9xfTEs9j8R7Z
UIbtn7ZHFdiEf+JzftaqLrR0rrII222lVEWNhUgEXcX6jS81Vw0vii9W6d/z0GKQ8t5ERXHCEWRH
Nn8lyslAODD3N6cYLvLTDtgH+hs9LlmIhCe6TRja8/iEfhATFGHXW2a1KMe8rwC8s/aXu9DcCndh
muroQlS223ECL64G73t90DlF0KYe3qFeQNWjpyVBI7xrYSf55SeMvGXW6ZCrlF5BwD8YTrTCc4nP
83YMQYhxNFSVV8o7sLBDGCbZU49+Vxz3V+LasgPQq/wooa3aJAOv6ObxT3GaQM41t+UNaaZgZp2Z
jxdGsAsXqt40WyS1RloBZPESKOm+tvgQfLaGi8HrktwCacaXDX2LUPg2wBT8NAzUmTxN9drCsdGp
PrwB23rpp0UVw1I+O2haEDbk5qjwjhQpjm50ebkDaYSqgdfHU5OQ1zOlzqKYFPMUGfKwolMb4kau
8FfBPaFJJuOeKHItrP8cD3TZiTke+3W/3s2nGgfUtj5WnE+cO+UMv/jYoqsg8NlCxUaSNV5UWsDP
wh4ntf0fDwke6X8QGmVqHr+8iBctx/rECpkCTnidny/Op5/01WbcL1ZsPji36kIuaO87RYcFGAMi
KxxwDRX1ec8IoWeLTojlGq3WDnRjR2jusY19HAeiS66nfV3AxJbW4ZKrhuPTygv6/JamkeFMS994
70FcNQmkgvv65AtaKEqawqLvh7CLsgmExrmkdvjWIAhjTz8f47IM04ELaQQz/M+bgRfUhJsBSLAR
qFdv3iB8gJwSIRZxk8XRs48eMPHJXTNdVzjYUboeA3rwgPKhrI8+F2D9JaZERU7gpCtC4kaL1sgh
hjL7VPEkpL7OF2eMYpvmqbflPleDZI0wtXV6qIgPnuYpkUTdxPCQSKlIW0JkKdS9VnRlXZpGRklE
GJwoemPXMUpO4jRajswVN4WSPOntyWzj3KkeO0h41Gs1pCnUGZcnQIcRsXuS11EtysAY5vAo8ONx
jdOsTSL3Ft4cUSw/d22Jozv2nKMVXIv5Y4z8VpVq3cUsaMrDOqtTtnmFKLDgTAnOQNcdpJYp3vqT
XAZ12efzo9abgewsxkjJrM74c1wa3dOl6r3pMK1s0W4DckWm+XtWBEy5TgkmfpSiiTOGCwrQfWzF
VVJxc8KsRSGaGzt9+0JkjFRiPCFsO88jAAvOttOomFHFfzQrXgpkM+IxAMmFxZXpEbbLnsEIghSn
RqvuVhSInC5xY2ubtQt76ap5/MmDWsJzdswZiBEp8fQzCV3/JWFrpbojFdJkhNEByXylJG7jnWep
HiGxgOX/F5Fk7uB+SOgfaxhX0RFF2p3vSSuZhHnrN1fspmgwD9i5TUxplf9yLLDnI+g65tZu0KHa
4tJKeSFuhfmd5uvyj4GOVBlAVSdeIsnqS5BKhrnrQjR8EThieQ19ub/cAqXnLYoHNlIY3JsoovGz
9B4s7BaaukSCC2R0tyIJLphk88UXwqYFtmXa+rn8WB06DkvW5Az/s3fXiNRZLqfg4b7aPUpI5FVf
0vXZav6sXJPpufj54uHhWA2cQ3OCDGthVZPhyIBgLywV66/VqWuty4wdqOAK5L1SkRpbgdg2z1oN
omCSz2d3i/lb4KsDMlZsWJJ72FBF3Q2mDFGy2AuYkLDdK3+iJZTYpGbGbUuOMIz1/870YVRTepHU
D/m2eYwtGwApzLeZdar1fDpfk5THe3ZRUHzY62fuxd3QY+G0FQcKaqH6dp7zkrQu4DcnnlrDUQOS
Fgaeuf1pXAFTcOvyQeCv8mqP+ajsB1q3r7DpEpQ2uQ1TMmogf1+beQbqKaNPZ7eeLd5BlyDNLy0Q
Xke44o3MC6RG9qagEMXooTEUiF5Gr/bXtikt7c0LAq9cL19sRNhPjv6Z0TEw0zmOOZjIy6R/hxko
I5hED3BmoGFvkawsve2FRMYmsQDfqYPzOWSH+DTnuEYQSkNBRq/rsXplmvxLNxeCC7XNlOCDZUYA
bBzWKRn7ec1LXI3GtIgGjigXN8hxg5UtBj9tmUZb7JjaduF/UTcyXEFWn9MBS8P0aMaUO30NaS5L
yJEOrHB7pqMX6ABthcSkWvhRNf5MXrtKx2A9HmcevbUEgIu2+nbr2+WXn/rySnc2BDYipGVnaYAe
v7z0KKKNq+CTYUxZcbXhtOyA+lPukC9VEKYC5jwdgRewqcMhY4gO/Z/84k6bnjVyoT3ABSJ3RS/3
8Nc+bmyfoDNVazwwdJTg7YfzyOFV29hKoZ1yN9TTsU+jj+NJKMfXmgAzW79Z1D7TB4dnJfPPgFLo
dYvCNx1NJ/e10GCyhTkdQ7t8gppbHx9pSzjhEWBO4R0bb89PBJT4AvG7Bqf0+wkkHWR1SV6Uq6gO
G/wfmhEcRqlJ8dDJTjLAe1JDovlZqeFX8hYJmbQmF9ELe3aMw3H00e0fDYuZ6lmt7UPvF+VbW31Z
kEeERLJuxJBF26u9RVEJVF6fsC3pL/XNwsmUkLwUGdrY/s9d9xTw+iZHCdIj8TKYWIekVoZPOQft
kTio50kIBUJ+qnBjgjHywbSJ5yrJ2OLoIaBKwfkll12bAGw8FgYn/5cwcEk8Lr4N9x98k+UJc9V5
KpG5xMYnL1wbWmqcYom+l79xx0N8CspcBppO75PduAlSekqiAlvFayuIbyJJAn7UMvLNs552k5mb
EhodGXUYPiCYORTTuP0RbQuq91mdp9MJHWVEk7oqFo0etaOW6vqcNJS/AqHOI+BT/NchzRIe4XFS
s/I0VB6zBLUxoyKV+caIN5JxFX+uyYALQyEOypOiO6MC89EGYUl9hcfnQ2x3IJvclJuTWrRxrq1Z
CpDd/qY1MixQtl9Wr1Xla7dC204XiVCr4pMf6EtEA5/ZlO3b5KSjpv/rNbxzUJuapCvJxhO5XwqP
ji+PQCAc8t35bK3FRH0luTQKSdsiIPsvGydompTXOVWL08w/0PwfIdy+mjlG/DBxrzGvS9fXTUhf
UZ00+Sb2ImFcvaBxvqRY68PgbxU/JRcDa2mzvFU7WnVmsb2uvELy6samyqo8mU0ObzXfPvpyHAOE
/khqHeApPfJfRPmCUqa/J1H6f2pgKxY0Rdic9kVxs3uBwRunAMxMmkIda96rBBj7HLzk5kfqU6Eo
N+G+zdTy533zGkZmhkx2CTWNiC+/MVhGioUZhuCULSRiu9VyPuIisZ6S29UMuyCU26GBR+QaqB6f
E/PuD+7ByGqNzb4fvHuvUGoCeeoHkTWeEUlVNqzgaa4FPg+VbIWlYL/3EafCdrC1YgUlKMIdnHh/
IVTPVdpPczp/2EByxCWaHbg/5/capZXE+WnKEnlXEtue+sTyMI73K99z3I9Fi1e+n2WJ8yuXxuQ6
V/hQrZR3m+Bdwz44c9dvac5YMpVnEykV9vlAVUdiLRFghgxcO2rltWcpAQc87wvh/DjcmaFDIgSW
LFonZDfIv/BtekC3FOacgFWu1qNsTY3wjASl5Cb2J1S9SzSVZhOkgpK/iGJI0PmEF13XsGC9lcxT
75jjp0sWa/F9YVvvh78xoMgWVE3PRStFVJjVH14bSUvw6Z+KVNPHSENOcKU53tAewTyMlNm2aCLZ
3fT0+IAWwirQTw/zWrKWYLSVrzY/ukK+BtzCAUUvyGgKW4l+l1S6qB3z6OoDqTY760flzW1YtI2b
WqN96ulKxLCWD/dOxzaZxeC5Wv99nFQ/I0vBiC06ESO6QVHn7/D1NQ1LWoX9G1venU6XSFGgQcLK
7kOcAFykF7yhSa+4SA5eDTBGV2fXBrrMywmMt7phiX/E4L3HUQBegQDUOVyMjnbB1VwZUI9vdIci
+K0ALkhHdXiAmHI2xEQV27c9mLvqM9ENLPmWC7dSUFUFpNY2ul37PceuCXlL2hsX+bnqk5v7kyi/
mSkXNhyqarj3O8lrQktP0Hq44/FSEHyNnPEm7NPzjm6EDubXQjKfBrxMJC3qd4VNKHiupyZZ+r0V
sQT4kzIPLw92CqZN6YpdyauwzpkmnJfNnxsp+sjhS4DLsjtQHYLEufSTZ8Ea2IV/otWvMBQOu1v2
BTj6wgL3haJva1+trZAKwU2xcAvkoblPU/PT115n3AHcaSchIPAUjrNkec18Ydh3y2xIE3xu2pk2
XPoCe99cbj4xec8sgI45aMWxaeXM4Mpbvmi86seFjNgIFJ7EYmkcaZeypAHk12g1B3Fg+xDTRffh
5H1jA815Ni0Fsk4j2G1jOKcTmH5bbgYxFql0Ulj8dDaGSSzs/VegVSSEwzNXpnCsc0FKK0vxHvUa
MotTZF7T08ZugbBxVIhWgJlZZTpB2xxoOUyIJCJjbjFcbRLW75nx84O56+keULZ93WeFwro20nYM
FdSrigWvz1rxJqFec3QVFepRiSuep04p2bStXABHSmMtUfQiyYKQQOPd3EjJXtWnVroOUoKK5nv3
kXj1yyFWXhKrwueyprZaPRf17gCmPwqCsAIcz6VvrlQGANPQ217vqSACBidZoSVl7mrxx37k3XXs
m3IjgePyQuNZ6r3QC6/aZ8r0ruTg35iMdfOdg5115xn1N0+afNEvZKgA6F89iF+SH0hkljMW6UXE
00RKWCEHtazJBGoGYaNMhrFk6dOiQEvGp1A/lWqO9Dlb30/3EN5X4hqdHqKtEulVn6LaJgaBHLtj
1ja9es452suk+0sBC1IePGzc5uqPzsjpTuso5qnO/Ad+63B0AJ74oxLd/mkmkAQhY+fdEeXwKh/K
tJ442BoS8rfHgclHcNeepjapeuA5Ak9Z9OUFKUWHhGEWrQvkLna/Ur87oDuifN1ZKUcy7/OQQWwv
rN2MbDFa7XeNNstNsY3wT0vZy+A7OUqX0NdHOJh9oV/UF00thBdgE2TyUlpGvFo18STRSsyrliAA
kz04RuH8eSPhJflmmIGRsdI3dsjQ4aDiM6wNXZLHsuA6CAwCTGlGiFluxAnOelAQSmIEId7HZ/gD
aappwskUalSMpeInGWU+yPTGkZS1PlY7DBjOeOvTgvHlFC2Z4RVuqB2ehIS4vbznNQZIru9scHSi
+gRoVeXSCQBjOEhdrW1eaIaCZPkKHd3YDwo/V8iFtyontwEjCaWKAeLDloB5xc4qVcQBqDlmhoUZ
N4razZZHprYLksn4iA0o8DaI5Y80zTaYgrZAiVtCDhG7L59fcLddjuJg3V+cVmyo7mqx+4te2EeR
GwLK+TWD5pQoXruNQFZpMY1EihcMUGqVPXmatkfwghxGSLvmA8StDgt8i+O9ino2h/ZfnE90MJ/n
3VNarYYUi2OVmMhmODXTSDgzpKNuFITUY4osdIGscQf1Ww9ynjS7KzgoZZ3h4VYPt9iclmi4KGpW
9uKe6b35u+jJ62s9YE7luEZO1aUStjjB720jCV8sCSqCiWsyIe7lcavKavHTP+YHXQM3zwM74OWV
WXmQifcMwM9GN0bkbLvSj7jNqBfNMI95L8UDxJ9XtZvl2xi/3bLAnt0Y4UsBCQHU29+8fHlE3IId
ougqiuHWEpEtwOzG8nCw8xSdQmu1X2RcDP1eu/6AUoY3VJV80wpFauBcAYbeyGzOyIyD4u3O7jXZ
gS7Zs7IVu2l7vVTX6d3AMiyPpHU3oO8SsxFk9NeheeZKZag/qG11qFZmGCfPk69j1C0yFRJvvRqh
dN7/Q0L7kLmB0N4LAPDJC0QXyyjoXJ5Idr7MLiJ2K5Chet1HErYei1jUq302LuG37x+wPXWyCD0e
v2b+NsXOfAIgfzpdYnwWGe0ImD6+3S8MunbubKFeurkVtBZTPsTUJ4ODpp04LZLr2HDkhfEP3vKx
T1Nzi2CwjiTt0+wE5SmXLLpaTHRm+4Rt19xTj99FP9W0jZTunnk+rYvVGzyv0J28hTDFXQs2VMXM
0KdeaXciKitLWy2QEunixC92HBqXOAIGIjEje0eCLk9mFHuej860vOl1KSlG70aq5PvOyZJXGUK1
Aqj5jJPUjvi8uKZxQMEnpEB3MtRQzZ7DSTqtXbqPKngPYcY5xKN4t2Z1Q77L+t5TCxU1o9pL9JNM
OOvaFu3wDhJn1ikg/lGUVVCGcF03wFkAPUx4LEzTv7/fXoo1aa+giBxwPijCttAMRtcooIy29lEh
+e5dF1I3skqLKV3y5KsjR9H5NGv36CabYNJfNw7Vb6RPX7BxTsaTQOi9ocMW+XCkwsbVjXJn1MC1
f8PaDSAlrVo8qfNHiVJ80zI2jGd2pRzcMj1IshZiNTcEhUj0t9Zkir4xMLo050bsPrSFWXQZp7Va
CdQp1dhozNwbnjCrPzIIcbIv4tnFDrme9h11nxcvluHr4kcyRCQa2vh26I9ILN4F+yFZHcRX58UK
Q3wUKzBD1aK6nbwW52TBY7t0mJYtM9ZRs6+Otu/yzETHEkJ5AQGB5VBQArOFIr9SuT8J3d9sH7mS
+4tMIOoZa9Ay4i3hI1ZFRe84yeOhAnSzksLBL575dwbkX44GWFWcO+PHPiAxM4HuRRPKKbZSjQPA
Idi+FSU1aDkPUcajPXG68grRHsBD2HFQ5GNOakYbA12OPHjh/9RxkO7j+cPYQyV2593ClR9WWuVT
OY5d0dDeWrTZTWbt3Xap70lP2Xk7p10XhHY3LSB5qbtyNLpbvFc3HAsOdrPYLzj8jCOuzXvJXC0a
45NczZSCVpvPON7+SAJ+K/l/FEPvLSf2CIMUZuFCPI+ARRo0WV+yBd3cyTaHPIw5phVPBJHCbfXj
wXxD3gr2CHKuoz3W9WCRbOp7qlfVFt6Wsgy+z63BgUJ8WgRAf6R+F0SyiUomPiuNiYjZv0rMyhHf
Kz8/xDHQ4uFf5GpLDWBRoyhh1akULKG9Axpepipcs6Rp2Cx6ef5vu2Qy/D7O49xpAj2L9/LvDnAl
WEyzTCNeCF5TUyxgijIS3GRBNSJ5o1O4iNDNSkEXXo7Xo1Tn+oKf3A7NzNyCoKT+E4qXnuLoodEv
ayivZKgeFUQ5D6tbSCF46WiLtU4zt6ReTcyzhnEDvsknCQiJpz/oalDMXnoDK1dESz7kZv03M/Xr
hvenXZTGSfPl6YienPwFeeP8sAtI/TZaaIJ08YTQtKV9jb+cpEeZAPnXtLHLSXU9zorSlaORmdGb
ToLapDwcPhjvbx5Bw6zceDc/kSwYFHycEMEn9QOztjF4/FEPpNZlCY+JOl7aFmEzSNHP/s5AmKka
uWSuzSMG1mCJuTN4+pscKESzvb3TT6dpOOC+XUp/2Sfu9Vt2t/mR2JYM4OmZakU8QVjm4gOpKTF/
wjg1GBSwUJW7ALpUNC2gbF0M4hnBjQ+EYPpgqCj5GoigIlFfBUVzem09xk5VN4o8FTtjlvJy/se3
eeDOuEG0uhKdVMbYoJ6s12YxLOkYbuMHQATjklpGtLIRU6WiauI/HVKJA1vszMozeAPM1y9aPQpE
3RNzzY/rYVPWaY/zfH82uMGKdi1k1O/Y6x8vUfLdTRIxyT04BocyV57Xla9kvzabh5ifkeuKlKsr
4Mtr68WsOXV/qesw566pSNmlv4L4fLXPK9VaQkPVtzQ0rLyK7Dse4wZR9JlM3WXh/zbO5QTlGWd/
DHbMIudYwNAuhJC8/G0HAVPJapvWBpsPFCaA9m8oZq32WBmFRG8qWCzq7nf1LJ4+SXBhoVK4TDE/
CB+P1cViCZ5uQhBpsP5yv6aN4a3iiqWgEB/AwoeN8RebQHxRfB0cw2VVoTvzhoV34D4SKw/QYX//
KUOOc1DIXxn4TjQW/HRbMMZNoxFK4COQio9esBHU2PqzqtcmfffqRSn92L9sA5y2wB9TdWzHqIqk
YEcIa6a+09hakZ0jP0+xyt7VwQ+CQR9dlKi+nrvymFBG0hMDaG7aTx0N6gxCAYFVvEKFqs+EYXbf
tD5oD4MjyapAKbP49k/sLt5a+NCbQ8lyv00cTwSL5yfQWClIPb4fTtDzqcOtpii7rARrIrNvuCIo
WWOFLmSUZ2ONDMg6c6SFFNDDkR5TOnqHNT6GSZuw/V/IVV14IbkL7xymHmAp2Yh1FD3UETflAV+p
mcSH1L9sLExUQPz+SF0p1BHqWjUrlbvQWar60U5Fg67hZJEWF49/hFT7Rr1fmPaJaHKYaTdkgYm1
3oIEPpfH+h7nD3D16LCeJguNspgbyv7VYpYwm/zWJU0oz2qNBeh3geghqhMd7Kjo7VThZktiR7YH
rbSN1nnJka+Z+HQ3w+aMuLfsFNIMt2WuuIladrDfF1+/6N0De4yEsejCuK5aaE9aSV68TfXVZe3c
TZ8IyeGo0kzyhSvXlYb5ox17rWdzilJLNxGkeXPtd6xqPQlrkON96H0DZyd5wTgChdXveVPw7G0+
lAY9LczYHsu8M87NCEKtrMhKlXmtVBE9SGpMTCFNe8k0mrSwuENdHlseYQX01xIQ9Zfnjed+cYal
IcGWlaA/KjeD93q4qefIvAILyf3YmCi4wJY+MMwN38wqKjflwHCEo7V3NxfUyjLkQ07cFIwWufji
02BZEPO6zVp03pjaajDO/zcO+sJDRGBw8QkRp2LwTxTkKbPReKhFeEn4hShclSztsNGQRy9fzEpJ
gDideeP3MjpadyGc0phfOF8clSDOCzci76rBbk0lksj3H//HinycDiaKwmdCYc1hjJofxo0UEFhO
cxLGwqkDnJeltzJZjIFWK7VCgbYFbV50VOosFNEbmZIWxmylgVzhQ48uGPXaVfhSXhEMBaOhQSSu
H/2yqDehtJ1TVMIrgu5ndzvrv3i2N7hCh7nnPEpU0QjSqzgNJwzu7qlgIRG87GX55C23lBDB69NS
A6X6iHJbbzt819+aq5EFD6frdRUD5UG4UrffWTKN5DeQ8JkYs8Y1mNwj1mLzX3f+cQdC47jdsFF/
VPRGQCoRXBDWvO4jStpr0bEci5X5yvAES1nDWclO/QKuaE3BqgN39hvwmjwCORAJa/Jb7rF3EnkT
/kbcd9s1188OKTkB5NjwwaD+50N1uHFQNB/x7q3D0tfWI95CaSCsCXqz8kTb/uQIGv9GaRIj0lQH
UC9355ZtWWBH3A+vXa9my+h9km8f6w44lHpEuh8/4fNz+Ms+gCUFpvQbflJHxVCgHw8j+YCAftyl
oIo5zHBMw+0rZitwJLnuOlkH+iLqOOuS7QU+2cvrhNyoA2K6rj2DNZLK6Hqv/xwTxNm9tdDXoBJo
aI2chs9jZVq5XkK7mF7KnmUAVNtAmRGjFTqCCv98d6WoiAFp7FnFomF9+WOXx4LjWMqGIbfKbNxv
R4xpjafiVOK3MpOer6w5xba5i1NI4mgoDn4kcgSRaBg+rftrBw82AsKJPw+3x2I15tzj+RHW1sIR
XV38T5WfErIcOnisSEHIw+2rd1dh+Lc9hFMuvV+T9IIcREyzlVYTb8HIPDuyTAxymagrJurbOKPq
lf9ONjJCELxwBbHN7ch+xsf3jlMakCfPLap/4KgfEZtrnMoTUvka9NLKwlMpK/69ht0mSyx3vTHg
4OUVrxpiZ48DwiIGzSFq0HPijEb5/NRrRxMWh+ROge546n6784QiGZ6pXN71q58oERAfIXdawALk
lcY6YCeVaRmxfgGz3raTgZhiwliTxy8wV1g8AAZPgsJBS1KwgisnjpZowghHxMA4BGJrI2rl4eyI
jzJrpx4tmJBCteCn5p7HZDBWUN9I2p9Ps+cPhvL4jbuGcp3bkovashFMMkS6G2hM9Cz/XYWR+YMU
rKXzIRg7A/jdUX7v9akKgjwVejf0U4P/8fYNNXTWekY1kb+BBM8voZ5xmQ42YwGIPKuuAPjXZIJ+
fV9j5PdGgz1JbWDIx3clTH4sNpluAVPWyIlbfElNvA8rBHc08cdcsQVPDTY2ik4hxyNnQK7+WbIN
F3ajnXWlFo7/6CknG/KFCLuzECmVwx0bgwpa6BSwDznIEBlGTDpdx2iqIsbJZkfHBIvogLEudEcX
XFa4ycYK9Fr5QgQkbBc3a8Wnt4mTHR2G+sK0gwp4b5bkO7+F6c+GVpeJEl+wew9RW17o5fOpx5kv
tpIn8J9gmEN3N8ByFoWhnCo9YU0xtuuIAG9PiIZlWcHk/UjD7V22fx1wIENLwlnG6B2cq3+Vomhk
hg6eViyeBv7Mo2jFHQ0XcxhCgO0SzBfw4NSe33u1CZL31uAakfFJlQUdX+/5xrg9YB5Aosdbr/wv
jIR501kna1Ezl70vjIFy4JV71nxe1U/HMy+ZXsK+y1gz+i406j/7l787SPAYEPlNZipIaOSLzs+B
yxFbjDYAoC+zNxAdUj/aRUs6G1X0XH/6xSa7ARD89F1VWlajfct3Htdk2b+LWLWWEP2/lNWi/H9T
fn69nu3kKs2THIohJM51PmDXbFdyAaKff/EGdYTCjPdoqcNE92dRH4XdUaobn7vPyN6kfaEbFaD8
jnCof2alq9XAb5agghguz+oBRjsbrGkauGzE9eBESs87Q3rQpasvVe/ka0kuRDxG8VwBFBtqugHn
llqMf0+AhxyKDn1t2GvyrUnTR4YndmisxRmQxnTP7B0NQyALD6/WboCmkn8HIpAoGaUDD1Yp/OJj
5zYiE5yEsFfEhwtjclfuwb/ltnGct8nd/g7OBjgtMipXgKu/7GN4UA9A5Kzz1mZSgJDQcp0cze3D
U/CgCvmfS0ARQ0J0vbRqAB9H5Q59cuXVyWFBNGQRQVTNFZlp6Efxfjpg74u22koTkxi1tD0G/hK9
B4JcmWbwkF84/o/4F+v6B5fPJ7flKMpVywQjCsmWkVLeid9iwEoY7tjIZiKeernpf+qwPmj8FWmx
En+MSLckjk2JSHSscK7QYfYbPZ0YdwMYmYRo+qsVq7kAIL8R9tADNBFHOKmLMR5h7rW1IDUG/mZB
N+MSfqEJDJZYFlLxgK9IRVfUgX2Ye7wzRaox+TLIUYv4TU/6WhbLAP8bP3mNpbG9/V29iQgOVLGm
0dZFyFXOVq6q9ucTWEc32mlt3X6l4uOclVnSjYUISEuPBB1jmPmJzMrEdmDVQ3/HRISaiYtbsDHu
NhgvGyd9bIFnP2GvAjXLdLj1TaW9W8yijH5ORUh7t7FSdrypa6A0Wo33CjkzbjspQcYxid6ZwX/X
D/DONpLWtzQ9DEe0Homr5i7R3mnR1TzWkRTMqnCcbda4c747XGgkr0mJXk3ysn36JcTvgP5li3iu
mEOeXAH1JCTAS7QuIGRJN4+l8/VL85GK9tzbd2Ys0lq5Xkl/JwKXsJcBbEIESxF/NxF8AJVWjhqw
X/B6R/Y5FK8BAS9Ixmk5MeK9SrAPMIpIEk8w7cy2oMT36nUVFYwOBqV9W9i/cg+/TV84awVMqYKU
TS2X3kzSPpLeekDiSN1GREjsvlM/jXmGv3v2GClaAe18zOuQjC9AIG5GTfZe+5TtObGhk5bhV9HB
sa7xjQ/a9a/izxaapAh0jXDTclTPdzHxcStRIsTRwjPJkLC6pOZybHfPqrn3pXJrrrhwdiL/Sg6E
oqTD3HAF3yjVO1F3vqyqvAOUJOsdx2J3LWgt5scJC8QSFmmStkMaMZpdXlqPDErD20TAOdZZ4cef
305uwDznRjEffty58m0qrwkvGSAQIyqXPfKe6ZWADD7kVuh+kV9ZRMdGAEuIf7hs+zSBfpFOvNna
F+G3LPKZ5Q/JJBUo1JTys1Ym4+yeXCyt2XZb0trZ4EoMXfoeZSloqLFHJI8F5SETeXTMX6KGa1FK
IqLugMh9EIeU0TMMKEIjJBnkPeYNhes9oCASA2KD2AShxXeZDBy0J4S9wpSCPw6/ICJvQpTQuqiC
FI2odl1Z9G6rsc0IMcZIlKbc36RQ9UZpN5QC4e8p5YrAJXhkoPguiSpMtEVyZ3lCuxM3bo8kSVRx
HNdC0lNB7CLvesz+NfIw5dOcSXShoSpIUTYWaFl2XBXMbWZVQE6rKvFfGw7dmxQxvoPcQ792QI0U
9Ja3Qnc4KFUKarqpjO2SD2i/rNy9Vg0+KtqH4u4rSdW33SgxEoHrR4wqW8bsVc8GltL1wVsYGXEX
JsTpY0+M5djUbjrNWordPmzvv3N2wbEsw3TTsbtWojCIEskAPnuCAX2Ifltehh3vhxmrtsiX1I7E
6YT6+Xl2d3ExwWIo2lTU40E9PZhzmsBAJSCps+6LoXkcOKla19v39JM+9pQSdOA+hV7P2j1Vzmya
wQYPx0samsEssZOFh1TIA1ljT8kGTRr+c1UDeTGauSA2a861APblBZZmd2wJpAbYHQV3rPQO1IpG
YxnHvaZqgQQFuH/Y3bd2a58NeXEpzcol8jbwQ3a6itjOHzkWy8SKyrdBHOg/M7dsyTMYiroHpECn
Ulaw7TWnzt1MzvwxuTBHW8Kb5wa1zFVYqQVW6dXV6rw2qgW94PhkrS98V/bs4k8sUaKzMKvfOYe9
mfKVwSpDmZS963BEPbeDO2kpwY8DS4CTS1JMWvkI97F5CQpnrBr0bvNYkkQMK1Ih7Ib7CVzwd+/G
L4AyKH2sAIwzxJNY5DzaVd9KOBQgpW9BV3AUkLxd8ArL2KaPdHw/R7bqLpqheAcqtWQdWQCy7SDc
ikqHYzP2kn0foj+vqPUOYupdcXzG0tRsWdVgN2Zvax2euMXjtMn0CKkyJOWLU1fTyXONb2Z+m8EX
p9cirg3J9qjHr/bv73uCcS0/VevUQ/OUM3son/K7FldDlvnAtNIVDfduztrRUGGLPbad764eLibj
1p1ikrPNl7bClyrtUMpIAeDcSc/LpaX8B2YPzTSTQU4ktyv0DghcJHg2Aro/CD8KCCuSrTbdo0Y4
ihSSkTQXjEshUYBCyFa9BbDqud4+l3FHe9YUWNlBJteYxAPTLw4KYvUzgN9HjgX7aU88M5u4Ct5W
+82LOlrse1Q9qo/txA3R+SZRHc2MzpW6UHP/TDb8gIze+CS0j0/ppU3BXN3kIN7YlQA86V+i83GD
UwBVb1Bb6bwJbyKF5fnz4dS7MfHYTYCdNyD4buTnZ56U/N8kS/z8L3c7PJnJK8cZ+nJjGjVjJc1a
jIzUGn2wTNPTjyhzYsBMlJxeyhZy18VjAZ7lhL39KjREUsG8Wr0sHhNDJL/HUAjyAx6QrpECfvFm
CjoqEpWlOeSW1zE+iatTneZHxSGQzX0KG40i33qh0SPDcJA1CR2t59TEvn8MdB9VCoJsu/+YivNL
wzDpsbjuWkpfa+jlXu7bxn2ueOSnJvyBI9yS8DeqTCdgnVJzb01M1dh0NSWf1EFEGIghwX6kuj7L
EYMJSOPt1vLUAgrqJ9uH2uyt8d3E32LZLx+fsGGv5q5YMDieIkOz/8AdteWeTck3uOT77Z+o89ZL
Gl6i9mCheTIG6C73LVvnylh6uEd+P2zu3XguTiUlE/5+eXCjiTcx0jLNmkeoiQ/obu5EEEwPRjxJ
tDWzhUu/6zbZ5xqcixTEwdSWMbc4tfrmvuWBYpJnFVTD7eIwzgCYaJORj9r1GYH63uL6IsfAEfbx
ronQt0or+16XtbeLjQYE7UdCCTcn4EaIyGuao1Qkt6KCsV2fN7PkLwiu2VOe6tMHC/0N0kLol3gF
0U0mZnfSH2BGB+L/eWETxZQzmqZFag73g5y9fSu2WXvaEq0rigvYEEB6VDufyZZbNHuLw2+4Z6H/
90cLKQk9Wz+BKo9Wmpaeofo2wwfwdHcOFm/z75afpdv8B3f4RInRPSd9inGM3BBh66y/O8e77aoq
rm/xbRJ0+2MTUmgI/P2uqG//7CSHzgZm74p9qM96iKVIcOFyNz2xvh4SHU9TU71p5ZWa5NEnFl5G
pB6dXqKSFjGrvGemPuzl10THRMRzoG7BS2odH5tTJhj9P4GcCczt6DS16Eb9SOb6FiK2qzQbECtw
d7Y0biMwZdnHtufKC5ZfghI2PxTbBnqBmPakK/KUXaTuWCkEsoq5jLsBk7eiKV8x2U9jzyd+LrQA
LwsfRQOO2yIf96VXEqvE+fEMhXjXaWW4fYc2d91YH9SDTxp7qCvAYVfV8pqD7VKxgT45j4oLebOk
MGKo28rWfxtwvrsVKL2Qut34uHbtJrUXJ9XeVW9TJO0yj4RNyTcv4g4RNznkyU0xgIzJh1Bs52Q/
KtVPfbIkQYMNbFuTOHinWR673fbHQmBOv7nJTtluX/VNJhGupjGMqo1ZznVE7MUmqChkXXozGi3l
1URPAjUXJEGN1WjV2lI9KRgt0FHz3z5ntva26aYPcgMZc8YiNc7kRq+ylGxNHdi+Ifuprh/3kwcY
p9NXP6N2r6Bx+UzUYGRJYAMlmEV+OL333OK1PA3Fa+hI0iYba2Eumnv4oVhgO1T5kBb+I6gyrXMo
eLcTC1EukoGFOnCCNNCF5XizoIMuYCN+0Pq/E5BfHkiTaExsRKBMlz511F0W9tPGJ0RvT9CUeJcK
XAzkQDPLizGFfRQ3tJ31tmqaLrmscrLoLDBWtMBA0KuqxxPncAzx01aWa/8CAvqGJqDOxK+R1ou5
3iqgND/7kJ6s49kRsqYem0Ew1YOANixzqxAt7m+FCwT4RWkcw67XlE/xBQvmZYo++l8xLufld6p1
tGkWs4Jva3Ulcf47jwX5KOEqz1rJdaR4dpMjQRPwEq/7GY3OhcASt/1X8O1kHrTg/ino5XLjLIxK
WE2udYij2chojUC3UsfWVT2spVt8zqo+55eCF/wrqGoCf5pcEDalxL5zFT+c9fq+llrazV5J3ZgZ
BChnnK4WE9cNX1GYs3Zn54Rehgiwabti7myN8YCyf54KjFC5PG1RKQbGQzA+7I76JJWyz8Wxl4Eh
Wy/3EKuK93ZboDm58VeIcOkQwJ1cRE4VXSdHzkN4t4iPn6b/n0QAOP42te9yLArEbbuuyl9j+5Ui
GyDSSNjEQEaadG8+TzczWVAsiyFGqqqdLme4aTsfr/cG2+ylpbDy+T+207Rc1j519aX+boy9oTo7
jbKSp3W96X0P266Fd0JYi/CV8BN7jEpbLZ0eODDow4Blk6OVYUg9OfuUbKaTk7XhaG00Wd2EbFE5
GH58Cep8ijzCoDqIKgSe7uOI6/YTJtVIpSIdKsPrt12EoSWaMJiaxUjBCkJhDHEidiPB2YxQMlTx
7IPtv3QdX+qVZi3AoT+s9LE3eHxdue0bm33Swlw/1vooRBDIKrraF7+V70Sx4l/Ir6xL4TOthp58
bbN2KTO9DevneWu43va447OvLHDUAJkwxv8ZGDOpyTn5yB2rwZ1UFVlThfGWLl83GxEaW8HlAhHx
3qhDv5enoohs6fCi2xQv29zenZ/HOO854Re56GuNuIwbMH47LnYyzN+8zlcqhtuc8cv1elqjDCyC
rGdJubIsslnXLXb0EviK5dNUMWZn3I2HcL4BN1Ovq1JO3FP5TuGQTwhqItf5C1E3jadXUz31Hpuu
BwcJoU5G8aYcCprz3dfboGsy+0nggSnaS3gIJAKRIzG19mFS54zojZ2XHlxgKbO+fVvTlxi0Pvkz
mJ5mvNchuGzISv+CcZoANmbvhQgidPWQb3+EDCRQsKk3tt/mBbw+NQ5ZpSkjoezhE+SocHuScdw0
kEzMl6s9rg4kvG0mxfiZvSyokI8BEfsKpMMZrVhjfuWrjRYBi2pmtu9IOx5jb3qXHENlJXHGBxPp
HzFAvLcbapHggP9aL/OcMMWndueXxntT8Mo3fZoOaInML9r+k+1l6S1XEcLZ8wUOq71+HEXSCtYt
VOK4s6Lr/t2KIp4Ain4koZdTALBiQdo/SPC8/iGdqd8E4rB9e3wz7HlkA0Byljmv3Ad3hZevvAXS
0HwZroeIRfsa0dn24G+1gkoJgEexGwmVUqycJMYp6WINrgIxWmHxztiWR7qJj+GK11gHDUru2iAl
qJzP+55Uy4Htn8q7DjkZik0jdgMr+4klC+aydpJRX9NfykaA+8ABodUbsjG7whfwHFNYX8OeCAZM
s/n2LJXe2aZDAeABeLWkkYxTbYtv/Sx94lCxunk8i/N3LnJMOw98dWgF1YSbP9qLbzQ3ZMmou03q
l5dDFP2ieVp4ApKHui9drqXcBNo2SXRcGGF+6n0O6K9co35aILQkKPwOqMSi6v9eA5lCH2o35E18
Pnj3ZsIVMyjAVjpLTYVH4OjfQCjCpGW/i1lSfkFgwKeX3jytdzG7RMwA9Nh7fv/aVs10y59c3/8n
AttB4ZKC2gfLBPaHqef0bm8jfM1gzAf/l7/LlUFx2UoM7iyn1LInHsUKt9fMet3ZiWU1jc4DJtzx
tZJNrsQ4DZcn7wthxayJ+3ipmFT5awbI90cJuBnrHII49SWeLIhQVRIrUJ3gljk5bMKry4ht+7jz
EFdEBYhZVm4m9ZenEdsdF6nsvL3l+p+3Ku13Rsp74c7HTP82gkyRjLC8YW1mAWJfMShegAoYwlQW
uBuZHtzptpHJXfU0AzVTRVcGFYBiui/vKABa9zrXKJE4n3L087Xyhp7qVl7dDg4sPOp54hl2L8bQ
tTcUwB9OT/jj+SvwlfZlWrMSF9BFUOF2EQ7UKleCjHNEFh6eIY7aX5CFqpFSOyymtJxLfnrHDbcA
6mHyvXi9DW6YU9T0q3AvA52s1M4bopldzHLWFL+6Jwf9E47yUm5J2zeiV1Ub/5Yp1mboO52QD56E
6l6hcHMZihhh+77w/FSjKIn8i/UxChMKlX4yzyTbLdrzTtmw56IJ+LRQabLyk8fV0+PBCIBRmJU9
5zl1xJfomLtoVqxmtWjHkQj7UAVMxdWE4VtmQLy5AE5MxEuYcpmBQb0tUnC8yUbhcw4FOc6W7rJh
s2/+6ZLlirt0Z6s/Sc/aNU32NyCGLT9GUTX32A9x32ehulfTNZR56Su9HCk1ilWnX8NCUQCDmivY
cduPDiN8n0AZ/x/cbX0EsN/zynamFC83xb5Hd8t5I0UXuJbgDGMzpA10/SXK6jM9SsLW/8ajOpjK
39XmwjwRJqKlFxa8RycpXGS/g6SHbdayI8TohY2pj0ePc3NYmBAONI9f7/4Oq/m1e0VrR5VjIhlh
IhFNMmMzqKkrznvN6q/Zjqb0JLDenx+Y2Idse22oAYJdlwd7F3WT0o2X+bAVr6iBHHV1PTAt+cKU
5nA7967JZJogL6CrbmKRX+buS9BMdPEjLi6taG+v3JzrInNaGUHX6stW2bk/PmTQaiB7FfC6641S
wvUOvpGKsWXkmCW0pOFPjBnulWjXA/vDLF4Z75YZeKTW4ew8UcfSy1stfvHAloZCF1l8RGJePAZ5
0E3HAIA8iDX7mDLy5PHBEJKoUN7NZ6b7TsV3fyKwMKqdKq9FioWbRTKM7UBa/cPr5+7nNqFIHZ7l
MPmI1HdJSJgt+LX81TaKQTNVXhYTFIzEYOA8pRiKGUsKVyOIIKrWrDGSvLU1yFnR+HWfdNfKfTDl
Efj1jmSWH00Kfe2W4Q0HtP9t58iLolzJW8iAM8oW/Vzstyxd5r1cq0gyeoCT+Qr1uSmoZw2t3Nnd
nCVeESkEYJn3qT4dZgfXOvvQV3KirkwXSBwF9rAL+Yd2DFBBdeKQZl6UrTn+CktTD2UIyJVUdmNW
sI/v//xDIOZ074Ccw3pmZz5l+tUbsuO7DsoLUvteHvksp/97326UyNyzVz4KgZPoMBeSycA+TEYk
CMd6ayJqinHiGXB6FKev6EL+yMc1lxBtfTtEyKk5IT14AdrX6xB68XWOaWm1mJdz8RXpW66sSH4D
9MAZkcaHitAtIRLS9ydG1WI6d1QBpjlr0DVeeDneF15+4sBMKlnzJtQU+36HU/oTxj5Rn+CzmV7k
pJ3xo9ayRWtGkuKfiKVQJ4CSnnHWYs/fwMoL5hbDRlTxWB+Vf3MNkf52ppE+43urpna6hAq3hT48
3Fhm4vO1dvYeq2UBup4B8CPWxV/XetGvTVb4F0hIUW3IQWJuDrmVTyM9jHvt2dubT2Jg318gMj5P
cvhd8wms+IYXf4AnM8cTAhGB9VoKzzFUTWBsSZ9Lks56etlVf4fq/0hZPee+QKhuPf5tIOwf4yOl
Wa+UNO89dfKci57tVzTRemYPu1jxKDWZAvSLOqmvhYcVuaI0/qU2RCH1r4D0edez4FXYScVwlOto
HxcwGxR/UJJGS8IpOM1kODJcSPuUb88aNg+0ZTeJki8yzoTbFDazo7LHRpb83ji9yYyBTghIiSVG
Kd5QYt28ZGE95twj3+lxUsTtO4UU041uQXxp1d0I+KIwhRdYl4b3AvNmID1k7xJzCperAdwtA9KE
Fvct186XNzZtTQ1d0x/r4mIsQGv4LS+9BLcRKZedKR+w7Ajrnet984ZKl1YT77V1t0ie0Z+xrMDu
U+1qFt3fZD0dUjlOJDbvB5rBVRhvHKg6pXlLWl2ZlZ+DJchMTjtCBaHOahu9hl6Us5vVT0W+4FL0
wRq7ut3CD+vp8n9uKpmYzQZ3hnEcCkiPkZ2x/XPKJwbWw4Q2sFSiI5BKgpCW27ZXKd2LZ2J49YQb
WsMMzb3iHZru/rJuZj1aaGR7J2TnZOMLEMSbYbMu3uCm8GDCMWUlXOMcpHP0O5Zuwim2a7kyrDXG
lVHf1g0fRAcH4Yf290edfflKheb8p3QlQmgfXjdkiRouksk+z3jvm0IKV5q77r7z3Y0srMAspb4n
ywzjwRYg5HnB6tViH4dblOPnuxlXDjtP3e491YlOqdFY4vknBSVGHaowHyQcAUMDggAl6GaJUUH7
akaYsXv7mXoRc/s+2pJPTChZalv3TEEs+QTnoiIUJsXi4nI0uyQDMTs7brjL40w6GNU7Mq87o5s8
bwHPWhLLYhZB6jatdpq06YHjBOxs33CauApRqacOzIwC+Cm7o/e26iaD5QSgkX/qAM0cQxH9nrWY
TVR3nO7b6dNUN4x2hmh6Nyjalvy7nyvmezeCdSxKkF6zRmg3mK0qUg9fw5tpsxy7yClapSRoHaHJ
qd68IxJL9GvqcwvJMhkpOzLByjZBE2oSxki8aAoozCUFyxPTCtd4a+FfnaIH4TBPMghXg+p7y4Ie
gHpdzSrc/2YCIfYONLA+xz6QQZMwBFqDyplMcucLiu501vhycwnBqCCN/qDgW072/jYRnsh50JRR
4cAghUOiF6CFHAALDGWm51D6j/KDDazpMQsMuWSbzfdI39mu58m7E72wkjuw5unj6XRRiPNnqQzx
jzURUhfSOhFpFb2VuGYTl1PnrMYjd5j6xupocsub5kAx7OjpQjbZhXTb2e5M4iiNQph/gl3dx794
n5kvK7F1QavHVHRYBjq8A1zdGN7WpZiJxecMt9KO3Vwrw1wdkAEkZc/j7iByj5d9/0B6lttKY8EC
ZP7lyJJUdeh3cYFZGsVsNxHBX3ZD22oy+VGeGq/yd6wTd/9jVc1Eeu5QMKS+xlrQ8dKLb00wsr8m
3z7WQ9P6JN8TSpEpTwr3F1uj/S6iY3VQ2CYkoJDW6m4+O/4PDOIcCEn90ydufUgOIwQek+6dkS8I
GZCowj9ofQ0K4F9rJLEmNzMIoYakmMQxOF8TfbLALtVvvTGvedNbsGvdpwhEbdLw4xuUm2jDgg6+
OxRJywAaBnrcOZj/C+GNPvdgnx7LdhmFuoRcagSzKz8L+nTHI1O5uLR00tetNGvgLrC5l1F+kO8l
qrx78l664XYdYcSNWmxWvi/GX0v9B0DWBj6sHgTMi+zoSkPd6FdxLIFnD1UJKQowlRDYOWm4wyOu
SYtlA+iS973pRJrt+uXIdvEa9e60cIxyp9Mm1pZZ2rhJ7oWyHru8cov0wWSj9q7qyk8Etg+EdWED
q/HaCLLZIdyNACfxzH5IWiHZJgtpT8DpneY6KxKx9CdAWMCazULgnDF50DWfQoeSJAUz2/kUnha9
QInzX4BNWNtg2ult6pfEH0cnAN62f2Z+dL9Uv5mwG1+SDlGAFc7BkaJbb4CZq6IJFPDzJ7yJhlxc
3uzKauSVVnsh/Vw4HZkp/d/sR6WZby8FdzKbfB1JL+qfHgHH3B2E5LJ/JWFTrVGV8n6+hzzAEvkS
DSBG/f2bT8YlDs7yAU5ShutVgPOkO1nIQ/OicBWlSYTXuRtePWGFh0pegc19dnWCAglB21mQwjL+
krjFNXeF6g1MarL0gDz9KxB/uzIa4Mx/w2sxK6LMZ8CTSxBX8iGYfQTnTAKEvVVs70bMey8ZmXuB
6LGPVp1BkCFoCSOZwI/w1QshXwgmENnoOIkdXOoyncxwwvEaYL7MbmXJW4x6ftCG1hSnKIckuX/Z
aL4koLcJZCE3DbuPa/H3UIkDTxjapIasx0cHa2dWDEvoFKl8Y94udVwim2Pxr4fpkWENUeTEav7s
Xg7fF3i0hPp64V3WyLBKsYC+aKq5b1GorNmqOpaTJ+iUm/g3zyqJ34NUwFtUg5bkvdpYeE/Sy7rk
EjHye6fF+Sby2HkR19Wjm8Uh8EABs8GgOeqOjhALK6eJki/I9qBN9VIBrtDa3S8/VHgUuy1g2VNr
NWaEFWGy6zn71qMJEcEfz1/Tiqz2OMi/ZJ2GJW//wL6aDaNuFnOv4AnC4ZPH763sJB3Og2nA9R6J
2kIC09wo8jaaCCbDwNgqhZgmgzBvrTppC6NOq17+lS04DkVobJrEje7obGpjtk1OSEGiPPvv/mKW
VSdCcF4KzHDShYrEqFud3XdV/GaIY8XB5VMWBv2x6SOLl4a5B/wf/LSGhIsckUg7OI3Vq266ZV9M
vmFBHWeu12sN9K29MJREbPLhB6K3JzPlFyxbAo+KBvVXsdHG3KIEgNAhG5Xh1J7Z4D8JMBmCyJyh
vBMwXPiC42dkcNTOhiGWqsh7afYUQSc5etrzAej1333zuMCaW1ivHaBIdzmshMMps2FTGWzXAp3R
FbyARzDKVotU0cSIVGjWNBGqoTTglp/GCfb+dkfNxhpI9jqUSTzu93FPH7LhwVZsBLfLkbm1Tg47
o3i0AG7IVBpTiS/F1mucf05lVrrjYaY6u/r87es6G69I5NQhE97wDo8zRo/888pF8Xe03yn6jUXr
I0C5P2AkbGFCqsg/3Fbdlr/SmljZr8mgSeMSKox2zsknTCH3F2l0vnDSI58E4BRTdw2+P9FHPOBL
yVrXyPS4KSf/X8PtvMFv0MmtmbHY2BDwLU8E8YMXNE7OXC08dlJsiHKEsvBbWvOhxlO3LWki8cKU
E7mL/3A5ntsR450zrGyH/Yvx+jMdnJqXR6vm8H3wlGUTe2mO7cRu3Rxlbn1wpqg/GMivPtnSelgs
jA5ivqNGGRoxv3m4NCj23pXiahUp40q3wIboassqeKw3N3PIcnNgRt0CGIQm7l0m6LsvJWSmNNIQ
eP3L5VjS9vd9Z1kuerGUhTU2424cxzVJ2H1IrToEfW2UWJqF4lIjTLznumd8dLBatCE16b4Uu2FA
0JlbrZ7TGWw3v3HVSIGm6atw6EbJ41TnwzymXXlXxcmG94VAHXiIcVhna4qBLOp2wkyirXT0BkgP
Odp2ygz5riH70Pwx9Km6paYA+GJdMnaqBOA42bP2uRegOvmAA3cmZcIIQupFgw/JwPS9LddNmP/Z
JukAEFldH+iiy9zVifaGs8qA2D931tc1lBkVOkBZ1jo+c54wkbW7UaC0Lq6yyAzNwlRSZ1RXX5Hg
bjtorXp5irQScrV7W1noKdkx/psAvvWw+XYbgVkZ+leRH0PejFFvqS68IcBK4b/CMO5i/IcmWhvL
ucaKGBv5tFXEbVtgXKSuEuB/inBZwhtwe6uteGAR7sHIizZY7BoCnH5wt4+yGvpPPPQ5f7ISA3jG
MuxFUIDwVUSDHinRdHLg4w+lrDqCDZWGDrLNW1M5TQTDZPzcs4vTgIFiQoim/IzHqNoxJI1cB7DO
nalRNERI5B2V/oMhse39QVKsgE/JX175OqVa9Dbk8U+7m1QwEUJZSlbnF3xtzL5V3yL2CDurOVlx
rrgqq2cw7zPEbhVkkcq02E3ZZheGGxz9czZcw3MV2+95SKq705BTiMDI9/LYHX5C9SLmFqOB64Ad
pjcSrXyU+k++/2D9aaWoKrtVqznyNJBDPp7ULeqM/yqOM+ADaCMdR2km+QmYAMQHCnocteW7UkKR
d4jYIP3Zx9kF8hgcGMWONaBDTfqdP7yNDTY81q7DgRTwBuO5nkPdJ+zvoC/WpEoi7vu79c4zDJcv
9XiyxyfxWbvTQeDTAkRnfdQvRpKcTxTkyRvjW/Mlcmu3uehy6D75yXdvdr3HQqjOLTW+KlmElRLt
eYZjxg5fMGxYvVzBieiA93jrUEhyOy/O6TEVQUDUlAIUhpGQ2rJktl2jAhjj3ZxRZ6tLdDJKpEMW
qoVMRRz+ZOiRxLHLEKw0gfVACPjhn6/KmMSL2ydwekdf+QGCtQdF/lDApiAcxE5H72Jvza/yEZix
AjLV0Mp3gK+DaSrO/6RBVRrxt7Vylv38Q1lK6Ph0OlIk1hjJ9bmu1gESjzACSbSDFd7c7stDKVjE
LKfKowQOgpiEzn/zVBiJURsnmlAAltk1BzTmvLSO8HKrBT4q8BkUjQC71kjQFYU4RrlVSt2uC+3H
WpAiE6qb6RXTXsZ+/eTW5ToVcKiCLQrUcu7+WXPkRh4wcqP4H6Lujw9EJLikXt+s4aC7S/WZiGWA
caGUrr7DGiSoEi6X96p5h92mY6hGqGzvhTQVqUBivOp6JZMQNZ2Spd6ywEPMlsb8XOzewIUgduss
+w7n3CZNkpdYqb8/NQEqfqy93+ViBD2kavKgndu9aPYOyPebWjv67zfe8VDstWlArlREz8uwHjFB
+uS6blvZCMynesU+P78rVt/p9houVER9RHHHNC+Ljk8WOWfP/1RCt09tWx/3zoN7aOxN5p0C5NXS
KazXOi9q4NtGv0HmUVHD6Y+etNSg92+VGxo+sxK8QANmarbBvUyGu2V/S2pzt3djTPo44K7YKgKE
PcUgb5xw0ihcqr21Fpb7d7NztAZYOWZgjHFYU25tiTUS3CLw3I7PTDTpm1jH4H+k/NyVENnMuNWj
RlOTWJRJk2wyEx1zQhc3oVo4pc+FayMadcm8s0J3AQ0BxY7aY3zrCB8gdKVtvKK1wfAFjHIB9MnO
wMm23tBDONht6X8epiQi4P3Qf1KnoPXoHf3v3j4Ot42IlYMH+yG0JKdDT3msLiaG7sEgMSMAK3Yg
bkE9fs5wJGWV1Hd8bUcj4tlgy0U4kPZtKGDQarLUEz+64hbsp67ftcimONDkL/xM6kVSsxi5TFO/
Q+OBZiqPdesn2u7s0xQhNySduOINtcrTEehRsfUoorlql80OqR95zB09svI9DLhhL4n1o2D+vulm
Lru0l16pQJLWUk4kzAMtqnHeJDZf/6raYVkqFIBzm8O3aruI1tDZ64lkFeD6YA/nZcu6UW2zrhdP
pebj5wr/e1+TBCkbkUzjs6NCCqxixrmLMouJUsb0Fn4xKiHHZ1S5eg9CsG0IJMOazzS0xLLC4Ymn
KrDDrwNFZs9JHrLUGRo6TgVBB20MPw0sXbg3378Xl8VHYQ9eXoaFARFSyRUfJE708hIc5C3yKizj
2V2vRu8jxyy/Ndo0kSZlau77kffhvNanS+K6S0JnrVBOdik9SOShwPXz40MyR9gD3rvj96wU7Tzw
8W1Z2d1qPJjSzIn1fZF4x9O+01BPMHuz+PuIZUbW3SqDKjxjqfZx3INSQZzfYDuHR3W+9TydELCk
q9aEokp9TN+FYCtb3/vn18bMdDigt81Cx4rQAlYGuql37qjOrho8vy+WSR7a6effJeL0hTg7U0n5
z0Jogq+hksP9gNKhjokZY98kgYyxEdr8o5rHhXKHsIGpuhenUB4rx3NOIOe3sevgrBgnkwWMMMr8
M/lv1DMgwmTQ/uVDgrX3kimrO6zkUvgU0/CDF2ku7TSXBLFA93yOu2E+2SaTnVbgPOSMBnQcJ83P
ng6kddp5bsCWk7mcxWX+jU6bA3rJXEk+L0gkTGYF7RZcphACJgxwRlVyJr+2LRaqzYRTN1A1ZA14
Emknugy6ff8+91yojzTRaMMG7I7bw2ctIFdPM/dCN8Yez/rwbvrhSY8biiiMTvkZdVDYtRChaNwz
RH7Nf9SfuH6KOl5Lx2cXiu/ezxDtYcSFLItQfVnDec/Qs46y9pLiBjcm3VrZz2VGcok1TcY2Q8OM
f1mE1IjghUvt5FqPZVJOczUzsPvSheIjCwVz7rIv0HQXGDxAAcplF7/st0HcSmKch1KMVMP8uD2e
6uhBGakNf3WP3HLIyhTwuyLiyj3mx7vtwkqB6C50mglp+ZTSv0DyPoxdcLZH2H76W+qqT5LDgvV2
MB6+lbq8LCJy7b4eN4zUZsKcsS0l5Yyxj5oOIywIsIiP6mVFnPmkXqwIOg3ROJU9Vj6q9ZcBwrvQ
l3X2FWev63YzveirLpw9Up7hShI8q5L5VbIQNtdbUXMlQyPb6hZrdFIBP2a8CnS3+iuIQpQJEHkU
I046EuJPjv4LRw//4gg0h/+2EHyCj9hb5LPdzZhbDkjd3c3UBmb2nf9a9LDyUIRevSahiCcWR6hQ
mFKOV3csK+c/ZPzvxr7XMY7uB1KPL7zsx9Tf4CtTnSJlAAD8AEZZEBEXF4MR8mQxUbhb1iEt8vnx
MaRCkknWWfb/DSV2TY5ScSs0bcF+VuopbUsrAJ+LJDBQs/l02ZIk0TpJDbi4Vm+y6bq8WsSpgdeY
XTUDLXkcXu1KU2CTuVX6YkeLZBoNm58p63tNmy2rBymEYd1oMB3iyn5BlPZ7syXqE2fRGliK3B+4
iixnc9TPtHYjjoCmOEvsD40iqQLInhM+2uUJyyiTtsvD5iW8DPjkQ8tG5+hxkqiK8kHVB5kk5Kq8
8+k0991+RM99aicUfD8hVEjczZl3P2YGVFcpERSffU16gmD8A2zHqhFbHcBcvACFAxUH/TW+ryJ6
/IuHgRji8q/UuIwt+MG9OXknfiEhqYZM0VEHXZi2O9CRrwk8UgKG6CHVLit3ypcUJGwLtvx93bGo
YkquDOwkuPlqAv/djAE/sBY+fox0ygjSSszCXA0KyrQs+0+UGmwzWoPMih2qJNURgOh4oVqVH2h6
9iSsMRT4qRYBLDAFfc7EN/AioDJR3CAik8DBqGB6V5ZzEAdMQ1X91lM97KHrJ38g5PdJhunBuVDB
V8vdLCdAyuI5rgev47wFbf3DkV0Jgy9KPyuIpDM66+1PgTFf2O2J2lNjJmxwX+VDtuHfk66K9lUV
NWHmnBmqh1xGVzclMIrItXmexfo+KGS2lq8m1Jbxwhm4s8WJB80uupW4k/uurNAQDBFZHA/cBHpr
DPBZ3UNSbfjYnJhYHJn4TJWN8Q8Tjj4QXKXfmPEVFjSz/QX/UIsnqUJL5rKe5KNVWvavoaz2pmH9
R/lBMzVGR0yKLbqjdqte4nh9gAvj05RCmIqL+BFzcolrKEhgOqOdRDxgqiQBVeFoXxo7jM8iHzFj
NnYSiNnKsvfQfiz2/6yakBKySc0KIe1nQeMnEzUhT322rfXu6G3RJoO1MDs4/37KOSUHJjIVqGk3
H2vE3UW617gEBy+bllcNaCgTBp/P6LmASUJmjTmJhNFgtjrLM/blUJk52aHYPmGKY93PPeZsJDGh
9LyGipwPKZgm5XW/zfkQyd2BlXUnGUIOJuQPr5CueNwzqwN2jlbFTAzaYAXCTFRBKqs50braiXOP
Gb/zlFGntc4DW2+W/nPnUseQIZYKVVZw8sVYcilkAKa7JnOLRQb9ENSALY6PGpZe4y/ojiVG5Sq6
baysy5gLGPmiMW8r+7pXIfEvjdTePsoliLAS9XlLmd5EaRLlKe5lQQ1LrBAOxttbjat056zJOdSC
T6NZljYFZ4A9U/ab796gkc2wW5jN1NFOaCr0vMVzFqmTfwt09x1KAo9EkBKCHGCcwKye+azQ3nUS
mb29+5IbPfvBsKBJcLI+ercO6ppNq2q8o1Rt5NosQegbnMH7MdJblW/0BQPFwbD9LM8VfpzbEVpI
/Efo31lYk3q0l40CrZPGwrq3yRmMUlVTMWXq9NPskC4ow7L8nAeeZQBjBV8AeZ/z8xCBAMOapFtN
7Z96lLTHLoJXglAcQvg55GsJI/8s7CE+dhnFoLUKGl5/U8Bpy6jKvkRPrEjFcDXOmsFVYT29w95q
TU0UEi16w41OoJrVBEg+lcQtEeMc2wE+BIEKLPw47chiB8tahDaB04zJnW2HSSRMXmOVPGcay4IV
jF/0B/R+gtk1I5z/XiOzOUxwXRuYXpIkwS1GrTFJdyiHZCbAeQ1gFwIX29xA5ddpfMf+b/QRxTH+
hOX+sueZvyJgyB7gDK6n/QypDPvwvk7uE3xT6aYGoWadCglztTES8WPj3uhbrAdf/WpDPf3JTQRd
51kITqc3p/cPvMuHqW0ofxrRVJqTaiwQtc4rDW+y8Vy7GE8GRuqvieYvvbZnZMX+W51To3IY+q1C
2Twz3rr6KSQbfNALMbeMv0lZw/YGi2tZVSg9naYKYWc8oFMjm1J4x/OY7jWW16fC8QUwtJoiHDmx
f7f7k6IOu+ZePiYUm8mQYVCbhU9c75BxqOV6s4Qw387zNT95ld9FVqH1xYQTfNLcJPvvd9J/iV7r
ihMfEffwq972Dq5PLWCWsBboZ0KoDoCXbUQs4EdEy9bSyckvHhlXCmL7L+hK3zCgrWueFs7z/b28
0O10BeV0TdXausG3aQGRlaFKvsB52UDdxD9sjYJJgB1hrU1IrQ4+irThgYj2p8sxilv2WmubYax8
HnrcZpQw3yD70Cu7udPfLSy9l9AnVkV6N1QWODnC4xYAxZiauDNgVNCK8Y5wdEABhIJk05BU6Qk/
xUxKacDssPi4oa6ZNFGUUPMtBy4XFJ+1aMo7JyNiBqUV7xd72UT/nN96IPj+HC0uwayXYMVZOgfO
F1QaYl5Qkkfv6kx2WLEJjOr77JzvZ5EIg41J3scaVajWuAnYOfMkuB2BlzGXpQljVwbH6pUvg077
LR2sCdFbyCkPQAvrsNdbjIaT5DgCPbp8V8cGz4tPHFkySh7fOcIvkNssNjFe0QUNN+2Vh6wX4x/C
+WCySF+0usjuTGUaGG2sVEEz8yxINV+ezKRuSgL4r7blhiNjQFj1EFrYTbZfSKG97k00PcDuHUTh
PFdhf/ssVHpYNqceTbYBHvySJEesUskJBae0BLKrO3vmeR9sWSmwdKXAxCrJ+P0fjlpG/aqnaij/
pAV16jYN/dY8h1UrUcincTW0q2IYtRcAq7zzG+9kmvVMDXmy/CY9kA7QC64KDySliIboDqtgPKrE
vUMHnLz25oyPy1MOOasA6yXh+KgH9Urn6E4L/KnU4DJfV9nWssK3W1z7RJTysieWDSJhltu9BIld
vulA6CrIOaM5OVgZ0LEjGV2rPoi/lTGU3Y3pIJdKxoXTwXj6La0UwhVGgoELoBpI3rAPP7Tsd/KU
f3AUZiHOq4mMyz5/ZLt0AgntMi53DoZ5p4R58ls5Pd5/DGEXJ4NsnrJvFl1/ct02EDeH8NDSGf70
pHwvEZqJHpMVpfTnheGIml2MtDArogDkRVWe2MCDcuyOzt41RyaWXJ94qsADnHlxwk0ffGdTQPls
cn3wGXGjQyN1TS/vEY/GT11ma22WK+Hty4SFtI9m2hSJhDVI77yBT5KzxqxmUYZ4ABTJfEWcd3jc
Sli7GrCf3dHCJn8sBHkuKswqonZrO+i4N4q6kRqiBoh2gCO0WB88qyh0zx2+F2EZL+yr+qRQKkwO
e5GoRpsQg2qAVuOZP4WfuY2vy2i+XhIGeY53xvAejj10FYKm6Mu8EduPZpeTgdvJo2E6j1hf+lOY
lrSVCwTssAC+in3q/UBHWZV2i8DLsVaEyIIiCgIUL0YkbXkp+2/4wE1p6WxTd7275bcrPqBlyWO9
WX2ySvLTL8iMVSjDF+SZlRMecohVPqeMovch9Sc5G3xMvwCbtnUXQOwanHHJTw2a0rRltp72i6ao
Wirl5X3L630TRsEpgEozKGhooOs70S8iOPf2a4tGr7xIOcQ2nsY2jEDaFMp6Qn53n1Ee41L9tFX6
ehZFUeAxqkKjQeVvsP3GP6grDZJL9etsyIveI1SYdHeKQOynZ7ec2w9u+4A19WDMby4S0qV8J++H
iguIfEK0tied2Jp71E++iocW50tx6DNi//SNfumg25WLrThHsLsseTZBrfbRbs/li+OspWMTeOlS
7zNt/IBTw25tp6hS/sLunK4Cb/CaTxko4xOS/EfPY2eNZrrl/tUYGt2I94EacBcdt4BF9WtxXN+L
re/9ZKsWXjTV0SsvCSWKRBRJgUqAwu4jQXRm+DQ7RLv+SOFBc5GWpICtSr4CNBYR+tGmsQuaeTAk
g6tfB95yrLdz+icj7njJZebSJ7jDaDfkR3H/VaXTeAkcZIUZZDFnvZv6B9F5zFU5qUnsY3YvDA+P
Cd25RiK8Kf9xBHPkpUtxV+wK4jCmo9dG6QNwiACYWKUDWgo70n1cY+EvvbzXJ2zjMknEw7pJUzED
2n/TpInM9FC+F6ZxkMxSDJG4XG0GHSvBCg9SIFJM3MSoWEjkJqwuq0eW/PoYcCa/HyWlXeP7UjOt
8sUq0mrOPnDBmDLGG8Dw93iXGyVR0p+Q5UpQv9BEU4SNFbtDVFMUIoeg1Cr38gV1QtB9aQkgMYze
DZG7Xq44I0nVeYM0m5EA1jst1p++j8Af72L6kiSLo3bZ8/FSkACrX82B8mXJmBt27uAKzksLmKh6
x6ARTptbypW5E5Dl7eDC7w9acR7DtRcly/MZG51/Y8aqYBTjoWCi/4+EYV2vESfMsF54Zcs+KCx6
KoRCOUS0XzvgUwAGPKKDsRk8rSLcuwz/rWdrazRRmvQSqmQYz9z5SmivGM10Svz1lETWC29DoFuU
v3fW59kGStfdxZkI4+4XGryS3RSllR0nFJMOM4I5JAAqDfubLbwaDCeJL4BZi9re6BlocJLmH1TC
n65WvyvQsUGJRPxpDAPH5CbXIMdKuggnx0mGkjaxoCYKMtyZ4BJR4JSy64cWWslSwebICC5GStsB
kQrtpH7Tm0q3/x9AX/1f62u6Tw5hZqkppYk8jOfX9+hgalEXr5+B7k4OZ7uhCJtVKscrv1Yg/XvC
NnQih1rcfZ9q03mQ7O8sprgQY5lseGMgAfe5kEm7dqSM0ZFbVb0pIBYTjUq2klLog4tUdp1hHLqB
afRHQJrqnnvkNkUwNvoXohEQHrKwT+KmRBCly1Mnl7sslYi1JjZTAHC8NyNSsJ1KLbhVviNo4uBF
xzgtIvd6m58pT3v3SEyWCSMxhPt53/0hFXi458bvfb7gT8ZK0Aw0y5+j6TidBYEiVoBm9AGaTq9B
Fl3ju53On0bxzp4uGcjrCDHEr7QLK7AL4DaQIJgIKWqEiHWIDJ9DL6Q+9UX8Z59Nh+pyu2Y9kS6Y
gR6JMz330hheyt+iS+UOfpLUHqHsuTy81xOc8uMvem40bZnz2vliU9yx0Um3mjDVLmzTzY3jlY5/
bqnEZQruR6weCoFVXde9rgsn0+pCemPQCHGp1K/zicYM+4j8OPPZGxgW7+2NNwaIJtpm3WLrW3u+
EFB6f+D7hA7rndoVbLVbUBXzBgptYvCs7QiIqprRgk3fgyhqRGIxJ9bntiXxIAIUoRzYuStkhj8A
LuS5sEsy4vbyVyNTLNAYGi6bzanBnBcvOsHa2FIwmC0kcY8EmkgD+IF0ecJQRnwI1Y8WVZz+v7nv
KST015rcebvtYN53LwAsn859ImVrxFZdfGlygyLlaEI3E9a9Y8OWAO1pnHd7lFR0rFCBizWYWpd5
+milL3QQEaWzeTXch+HIyeVbBzM2VmsZ0cGDZFS9tZjNnhlX68XZRbSeZ7hubMWO9eiQTKcr7PN/
zhcyKEUuidmeV3F7jqbj2Ep2J+liSTUPsqhLmVYBsGEB1M/IfmhahJWPNwYAvoebomGnJHGKkp6G
X+83b0BubaV8+5IsfvOf03bxj+ucpCy7USHfIEFqSp5GdbtsvQwaYTa6HzOaPMoF4tNgJhM4+vU1
jhsQUTXDBTfXhIOA3n4LDZif3Dgy2b/dazsWKzTIIHJxObqehQT6kprsKQKfD5NL3dH58LQuXm0H
D/47v1Fv8EcI1rYeXIzpOEz8W94XWOaGzih6htuhzRJlJeNHoyKleDHfZvjSV5PBjNc9e+vu/4F5
ot3GwMfzogcT5+Cnfc1X7b7VntxizZZIFQBKQioC6NizMUaT2+zB1823hbNhLU7narlfv957+S5+
5Rin7OPrOJYhDfnITdAf5o6ex3Q/2JeXzYYKtvD0OfkFkTw62WtrvT2sxgMmnM5FQ+3STIhCUOd3
CPSlD/rZb69Ezl+R5VCTGRGb15lPraekeWXaNC1cijgW7MXiJF+KdKJ1Ka9z9tCTemDgPrBeIxo4
fQ9mV4ZJP5QCzvwMA5FuYRVN6qYATIrBPei8hXoCsNmi/C/J5UvJM7rfwLb/jAjOfds/DU4/dDV1
Z957IkfE01PBST0kuLwQGQ8Q5J01bfwWw5H9Cyfy47yXXcHJJN7nsgFTno1ACtQf0Y2MWeAm8wMH
ORCRRz9M8gWPJGJ1xY90upb6WQ4WvpjLHDbXqaZCV3wcdipAri0ZBCBizxJuTgMIfLC2iyeVLRgE
MO3u6GLRoL5pn3xfjSJQ++tHlZAfTFl5ItUoXfmIpDvQQtwE5KUSnyIKVlnhHiMkuDzqyYdq3rkp
43TPXN7q6/tDTj+9mn9Vt3Kjv9JiFjqo8LZoFg7zdX8RhGc/LkJDpSvHMgWI0ueFQRN6o9RumgBo
2fIlRvGJU1KI62BjzDfVEr9EsFhwe3RSTlzFTbxj3CRvtcMDChGHAELOekPUseh3+q4VuNHrlvZ6
aAJgXbhwOcyT6W0M9rCz2opJqkW49VMPid5cNIP+FEscm3IfSvbOMOZbJgyBoOfk/m03N73ICzRP
bvhgq2a9Q4sQlsAIkSpEcA8dsqdvkt9o5UWdX97TetgRteRggwMUyIxgfKHIBA3IsBlakYMROjIA
FZfO7L5EResJtD+89yQW1lXAbrekQBcgZp0p+9AlHzwWDWL3x4j8KUubjerPy5qF9yXGm1VfLNoB
1uMgueheFRg3ro2z3wxHQ5d0UU70SxDlTbW60+D+XSePWzGSFsKLL0m6WifswpLaUoSiXi2WtJxb
ynu4nuxsOWqqRfUHZ5j7wGId6udgENO9tJ9YB8+1dkcpo27p462uHigyuRVbyGnXbHLsmYBsVJIJ
UfYyQvn/beUwyi8FR7DAoGuxMvE8dsSrD1N/WAK6hV7SQKMc7yWXKgG2KMdJe3Nri974sYPfR9uO
R7DcIuH/h5WCTqO9HKEda9jiMTuVMiugApbH8KWZWwohdHrXREWJRbXT8NL79I/Of0L5pZsEDFkf
2b7bdW3D3itPpy/sYkrXFAqV57UA8iHoWldbae3EWF9RM3XSHExMg9/Ou/a1y1iH1uECZfw9vHqL
DuU+bc7l2T1SwTUZ0N2Z4R+b5sDCzH1nmy391Sypg7Y5smy5eTAMdkV4Rj60lyVBjWZogBbZx3QN
YKm+MbYf+A/HWTqfszFFNHbMcSE7ium9p8uN6LLKJXppm+9FJz18FhEGsGgi2vDEuOEm4o0Xlngb
8aRC7AfVndtNRY9SWtUI1qMgWTiZFLcc0K1eaPeHiPGW3CH9fwG6p5nmhWOTAAo1nT2/N+9nQIPf
hullEL7Rz5YwJMR7Ns4/T107HNP2W6f6kj8NMu6pWKgUUeFkCsL4n8+R44leJ+uWGpIK6fbwon6U
+9ixiAfmUzTQW1reZMwfGDWlB3YThVJMAEMVRliogJZLVWXgrw+UFWZtfBQORN3Igo87Bt60Dalc
Tpn50nLNZgC/26TWSZAImgKtzG5AUUAmWdS4PVMKEYeU9djYtg93/151GRbAFSqjlHBMiJ7zJUOf
cfjaFmwWfmlx7vpDuTGeluo7JWU9iVFYzdjr88beyahiQwYcK67KFO/9ZBkNJ3GT/tsICfreN+gM
45XAXe5VlmnRkqDMaSq3Tzno824m4V82MdXWkovcdW5+PQI/afHqnoLezSI9efj8VYBZZ06lpoOD
vsyLPHizQOpFTd9oQiCdxuomLgF7ZE0AZZdTcU0KwdcdFp33Gbit8aVKHAaO9wlA0Envo7vPdKYu
OVjYEXGc4VyE/aKsMhI3EcKSLbP1L7Xjnz5hT2HrWCDJsj+wzRl9vXRookxvG0Qwkbro4gVtKWq1
tcmnFJ+Hz7YFn8zixBrct4ohJ8v6gIUTAa9zbRfMOC6JxkZLGrb98y0+BhdkNFCwMzSB9aRv5ND8
JudCiyrmbk7K7dKGSPV+yq3YlNW+EuHsHWToiA3Q4CE+F9EfIX3osfmdeqkKSDJAHNJiUDU7OhfH
MChXZoCpo0ei4frpyI84BbNwhIopz84ccPiycZ6rYgxfVaOGF8ySehlipt6vLTH/66PVNwy1bhRn
yszFfxlyGxopZdEA+pS7/ijPiPQegBrXy9Yol5a803u0LqTL6QK61sovXRqv8eDrWUwXwZZ5AW20
t6dY8uXdxMlf5B3SuEBMhDYjf1eEdkR9jCPS+2sdohR1Sv1aStzpcKlQPlrYeiVlBhcrH/KBEJUU
W8LDHVNcxlPmChb4K1CKKXvSx4lvBgFAMXg89/Jxnbg63zL+p5j44SvmH89B/9EfaxgHwOPYaQhL
wa6pqboE4iLBiljTcDpHrG7YuuT5xdqB/sb33/830lHYB7G8/1JZrA3X2E7yxYoWmqc5osKgp4uX
lwisU+IS+055tZNL9x2tiO6IeZ6qH2TRs3E41Hiv/NBHxAwn7P2qTWBwddLhL0ZZtTFriBdweLo7
3q2XPD7+YCYR86P4/iBfhqBnF/W/Mcj5C02fqednngmE7SCFiDFY4nYKTopwE1d7vNuC+qRfT7ck
aJrAqlPpd195ZYxpPO9/B3MGWYevqvxiy19UQ7FeEVk/RDQ0TKaYuysG4/pX9d/Ak2q7kRR5o8X6
BqUs9bNXYM/23WqjKzvUQwcQWMy7nRmhT5m57YQwf6KcH+oT5mmYECaWa/g5EkPgeMF0l6CD0vhr
wj0uu9UI0uy6jifyJU9h+PKJ3HopVJFvehCgTIdG0F8MhxU57AmYnM18v5Aht9cMgVKbjowvq6UJ
KLiQqij3a+ItbAGjuECmFJUMR1OkvVwNuiH9BQuew7Y5GzQB3rObyblTKTvgpm0CS3uOJFx/+GgM
C9mmCaV5MxsKx9m89jEGQjA0Kqt8bxixjcMzM1oqA3DqNtKizE/utsrEIXC1aaMbSiYQ36trIakO
++vncMVH3wJQsf4U5wb5TrOnYPh60CJWn7jCYcawqJ+7iJPSjC9qKZNnnTdutyhfrRnRChIb7dmW
IeStBR42mUAFWLKmVsWZeRhKb3qV+bbwrKVQ6KgutaaJi65p+PbkMU/0QeRpYcnpnTe7ebPXTR+E
1qH5awv1ZQTB7E7NsOYe38fvsvOU12X8uMyJc+PKzpCbp7qPHWfAir/KXrfj7RBCCd7zd+mXC9eV
1CyXmhxz0L3AgjPul/0UR+eQpkKpCJD+x5NfJTrVCIgpLHpQnpv1BDeIh+TVHYvWqpBJJQU1dnSY
mLS7RVst4WLzsmq+EbNiCEjCF6A2M5syCKnqf0QWymu6mS0UYAhrbjAGI39zHfG3wkxO3NmcKJ60
62LKs7X3MFKHM2BJlfV31KQTN051nf6Ek5M0ztjDurmLdOex6VB8XVS+9mVpdurCW+anm1MBXaSJ
XNGMssA3qQV+bM0BPCYllMnzpPuR94DTWLWJWXwmO6joaA8s1f9ZXEXAVuioJE2Bd8hPVnN8G248
ESGeLhCK1p46eAhOnBQPyzeTeARPt8K9W6RkLAP6EyIjRf02mC6s5INrRjLdFDrSggZhG+9nno/1
CePCcTw5m6NQl6+QGcKoWloC+Vu8p7GMZ1PAN9qADgF6Vo8KZznnuZkbSF60d/elR6utbRNfs38g
toHZiE6vDwwR/bQoectfmsstmFfaW77jBy5XyEfVL2m7l7dGMIUtC1vjqgHpf4/R+4LVbXFQbDys
a4KIzHtENAMzNLDwHlVNGbSkUmO5AU4qNGSgBtRJ96fCbdroFo/sifnqqeeWFYTH56wD0HPV6n4C
HTkAGcxwVBROLyxbNSX4bV+JozBxEsBSiifXR61kyJA7YooHjKtixhQuhvGEhjcU2e5Rte+wRSmL
JY3pjUicbaMgRIMyNO34SsclxxkEyKGqICxo5UrAJSdCqNC0zyuVkCcbehXeWaAlsAiNhCN1ZXtw
YQeeOOR0BHpXnmlA/HpdGPVwin87oGVruBd5LOX6P44AJw3Ytv/c595CcAvVH50YILBGYtUEKt+V
6m8vkabwdPoQfccv5o3GoiKTtH8ByeeHsCzCj1o+wDpsrGl6AzSjnOS2lsVDqcyeBzoml0Vxmv6w
2KsIcR84lNoHt6CQ9KZZfJwpPUkIh7JJXkJfQifjYSnJaagXoyx/dPkgF3v42AOjxc8lHyFL0iA5
w+Ib4nlrTKIuq10CsMo/0H+yc0wfbjdp7DFxfax71FMGDcI4cLyVc/Q7tSLmrb7yatwcdSSM8i3q
wUNLie8Tgb9udlUWWDJ/Xc37nW/Jx3lBWwyMD9D6k1Itei71MDT45AbqMAtVxryFysO9thmLaemf
TivFZlyyEwCGYIT/Wj1ZqdLDdsEk7itdvNjdXO0BzUReUFYGdk0M5IuBL26tMssyA4p14OIFG9iL
FV/fHSylQGlWuKsjEl9WcZb47KjuFIxSBEJfmLgmbTgg6VLRXhfj0/CXQWsR4I3eITq9hCUonPsU
pUOU+EepaOfBNJMKV8hEPaOOSnVx02JHcJE2lkEIL5CwY4lbjySHA/MFGQ+rkkkKA7eNBFIr3Jk/
zcD/2rfOuhyYzzuOFb2nc97NCzt+4UBv4mTB5iFP20uOYdvfRfGTCKmX0vPDORRBEq+aEFZDqw4M
LqdOQMgCrZnvikw47TkoybntAU/LucGtEV4E21jmP1dLt1NpNhRu5wX2Ak/r56hhR1xjPGYZAJCP
330tHWvimYriWKhjSBNIX+yKr9Q77+bvm0YnQ4XSgUjTOCRXayolY9WEfyKhsqBrc8gyBIO6IdpM
FOk3nJpqOfVN30kQlL0iFK9m8jHiXorwwGL01LBv7fAd/KFPTNo59QOIAUguLiNlsgfXjfz5FYmA
s/i/F7bGvzBFmeexqbSPrRs+Xz4DKE+Io1BYSt7fD0cflkJ3s4igqeKoew7AqNHWgwp5Hi0v6XB4
TafA6No4pk5buPLZStblsho6NqCshrxNaUYo4LpDC1fjLX88UAsMHfG+tFWskonk6dLTAloKrBnc
FBB33ciGnzySMSL7gJ6HtnvqB/0sFkOGY7sWxRTAuSA7NOt3V1IpAeaI5UH5EesqwOfC4PAocBKb
pc/RBZ9TTtd33600n3jhFrQnDgKq1F508cGgQHBTl8csFLZ3Rh8pCpP2JM8ej9oLVODRxQtRBAij
kweqP2TgvKDXVwGigp/vRxA5gCBqGWILzqO1ZFw1ntaKHhJiAwq4pjBRE2IXW4j2WPYNcjlQCJa/
HyOWt8jDeI1+FFC99M27p9QwAw40/NOoPUUGROgQheJYGK3xM2BfSSWGcFzzs3gncRM1IbTf5nMF
05sPkUZVVYtTZoK8G0ulKWRD73X1o8boeOk6i9zth8jpDWGd48POd5xM83urVpDwQyHUv3+RxTLA
BOpbqBEw8CrzwH+GUXXmAIDBILezymQ98rC+8ynS/TIbdD86uSK+pBgukiNoCV7O66R/KkHHyPz+
ic6PepgwB+7y6SuIHqqXOeTUndoKN0a1QZAOr7qSIv8MD/oApwolEErAhdvObtxqTU6CRxEShl8N
UqodO19BIyIwBk84d2ZiLdJKV4Lw8rTfpH4sEiaZ10a+29Cxc8liLpSXgswHmLu435R3oXY6XjmF
RSdLCvR6EfWHHqc++zlXAs5YWv0HmdDkmQIcZUXul8QPNTwxWVueJxUw0Hm2kfs3c3u6bb7jz1db
O2OG1QXdBV/sZlJmxQh8KGe3meNd8Me/2a0I74q8HdyT+Luoup/x2SLqwkkYIsZYULpChGQ1CMTi
pCaddkbbawo0aIN99qRgwUVef/w2iUBKlrH3ZBA1cJjEntPM7fIJ1M37nmfRn13m7VeJZIAzJqCN
kkBAV6kZtunRoAZcU6zE+M7roR3Q+MqKrvXtLb/AuLPGm8Zen0gHRP4fnzawtikmNOJgVp2paeAW
1zimb4xPzk4+rpUEvj+evWBw7V4onwDM14rNgjUNVuzey6tr/Mw7MXgFelkd/XuOL/XsuYs/0S0/
mHZT2GSISxp5djcPJfCdy3pFL0C94/LVzCTY1dFUk882We2m2bNZM6AjsIWllXDoKWzMblgEPU01
Y6OM+PJzQWEDpL0yMtUJGJJGl0Ymm9jVEQvwjYqIYAWLw/PNPzbF6IwLUnw9/r6fbzthFAZu5PZh
1S/GvlQB0MoP3T98RTRNA5wzL5wT0lAK1jAuxwppvaU3B5KVoSXVj7sIwg6TDve9SSB5ooXiYN5f
stSEJysAJscEkzLmfRh9cnqLMn05VHuKXOUanPrsqotvOtgiZ1GZ3vE29v936DYUwXKxt0DGahQU
KmEOt+ItQqKYQIKV9J0TQDiU8LssJ5vyYn6rcpWj8Qgk5DPvhg8udzk32uGj7DmiPtmBoTG+b5GY
OKbGyYdod8JOZkunkRLoY9dvke36YHholy629A5EJznRkUNANBj9weXorkVolQ94/wCBx7ZyxPiK
ywRX4Nl7lAuHclSaI15PhYxlgRN+TVOMkONIgq/G/YSBoY2v5Wn6M7y9ydWfFCdoSH/xhVHgW9Kx
LFxL4dYgu1DCfNvtkttN1c7wgJaGVFMXXxN/y5eND1AyNhJ/ZI2makkxH5et8BhyOBh+vxTcnBkD
7JuKaC6yZCQLAWoSAjSX9egTkspGiPIanRdRxlUl6lrlY5Vb7m44pzoqG3CeOASooRwKZE6LZngp
3OQnp73s1TRcX7EnM+WaU+NhyMb0zPxiCktSz1ZYFsSLDvVQB7+tFwD4fNN5nLcklJjGPI9Aonzf
gF/cPxrUKP5XSFKB9kw0Rdk0Tny0ournppsF7dohh87W06jYnuUd9w8hBYVR/2HcE8GTdNDFgbSg
0cd/gQbPJOlrmgiXAr/qJMpEy00BCHXZ/+e8GSR1ald3HNGAsXR5Gk6F+juTMXvlvH4P94p/rG7z
FNuAgjPyRlFiYKDS3TZLjYRLusuroMNsqrY5kEYnmcmnIrKFga0ufimsYskszCmewd+113hA1wfc
gppPLkOoBFnUG+vSoF11JMhc+ebEHlyXkyZq1U3vYJN5QJZwi41GcVJshGOfGCQmXOxsXJyoqoZb
RvXeW1io+pMDNuJNluy1olFBP6Mqe0P2Vxr3CPU57v28m6KX2SVYUwg5iRuwiOAQ21TNUKxwmzih
J9lm1wo61qhTgJajN/JJiE3Q9666tj3d/9STnY4R7fcfosflwnAl7ZEDWF1ETPAaoel9QBsnU9RE
JlJkTJ3Qlbsin58g6kFAzK/J4SzIeHT8PMU8kI2Vgw/J5JOQTkvYiSFFi2+ClzdYt+Yih0MuPH+S
gClMqQmFeC4cgBUCZIRzhjjVpWFParC4m7LunV0nm2EY43cRhOnbKavEz4TrCN1/eQnQ8Pz6HDjT
XLbzvRo+SI97zCltJW29/BzcfZGDk4BbdOR559N2krstvrNG0EbVaJiSeE3PxYKV4O7MWCQA5F9K
/YsF+BYDyZG9+3kWa6KcxT8BtK8LwC/U6as0Bt7wdTjKX2baeRzlMkke6k1OgjfJOSZL7pYFTn/u
+jZr0I+iqnyfFybq+28V7/sYF+Y8KhuuH91swDMWnq6jSHX8awyq8MD5qjhtEQXl5JnbA6IMf39s
dIyG+OwDSAs08qSRZmW2rhTTsFoxGtFeQlgV9a+qd2fay8xYzJGsrSMMmvg0dUKWQxeDlAnveQyt
OsstfVwrVpoUuHYuT9q/hxWeN5gSkBDwaUCSv8yBC7ZNyD2xelY1vLz2rD84qRra33OzVm2iAHM1
xM2ujnfyPvyolP926cS/JQvDgdrgj6oyJwCYDZ0C4UlKqFVAb53OckS38shLTMgDFw/LGb2kdK4J
i0oXa6qF7gR13YqV+5+Y7c1UObqSPI/4DmkvFlrwRPfUfF2Cqn7jUyqafqfOeqq0FXbBWdfuiZNm
B+eXOgN+nSqsqcSPwQNrHhN68V5Sg83IuIigiyZ3nyR1ye2Jt9qixs0sxdkv4OZfE7BW+vB6ajPo
pCo+8hG3kpa0xMvJVrakDDXjjewAdUF722S1cByZWheSFS9qotDQUnSpzwmUBQrA4LSawNR9Ridj
BOBb4JwJxUkM16CJs5FSo0pkRPjkgr9PYbrjgXh4+wSP/fiPYVRHcOq8dhw7m6wPZb1/Q/370GRr
UWNX2Iwhvqs6cJ9GZ2XOrwJqL3j60mnPqOr1uN/p6YuME4L0XU1UEWG7EY4Jr7gsXoxmGBU+FgVa
BsaDW9XlvJe2SGT3h1p7/04VjuKQhuIa25jWXI1673b4kYtoFfsRNfBOeaQOwTtsgICxhBryPBAZ
UuJYdQ062LCDzI7goy8lpLXVm2L+UJx0xBFiSlVane6jiD6Y3CXfviUehQkqsIxJ4uHVgyTsAQIf
ZhBhXEbMz4dVSo4AOuIml44QyMxoUFBtgDSLQLER1jUgNQpJ9xvKKpnlft9Z7oI/bkkgCDLDzo8u
NWdO6UgLAn4JSfqBq/BEUU4FKVrnRAaK+t1CyVxXCgjtBIbrlhGsoOswphvWUteV3WdxWXF7cHCz
ZtWyedLFYuqRg3TaxTn9RLfva+EeWQJ/Fq3UMFmPZ010Xv4WSno4F1JvKoohIB6rjeQ491FmxDj8
f5QaBvpTSDWgtl64lSeu8xllZ1F+p9cJ6yy8HO47NTNO0N/F0koqnEnmMa1DTCmxB4oLwX/K3m5G
GJ8I3ZXjo2YdZsh6TSm/EvpFU6xvFTNNzioGEfxnPZwEIuHVE/6S6uaVETS5YMZmcW0S/0a9LPcN
jLo2f6lL2WCX5Xvqaqi8skcr401aUIFab2jX5kAAFx766+xFoWESARfDVOWqL3qfzBAT5VyByQ60
VoEjH6XPI6k///swH5vesdP8xu3SWg9VcFfUi88YDiei0CKGF9C/9W/nVZRk8rHyEHNL+2ruT5YA
Qu15MmMXtghyW+uuLRzJHDr+RecChpdX4/hb2LZh4Qss5gVHlkCp9S7qSfMA9dL1Wh7FqdlKa45H
eN78ozxM2nc0ioNk/O7nkh+GXTq0vyHpPG7nK3f8MmK9c2tYRLkPZ8BrGRZAkFFO6MtC7kfDdh4r
i2b5yLHIbpFolnw4tmrZAMhUxY+ly13MI9dgrlxlUtzpkWCCvT0Ha/dv+ENnpzXbfHjw0b8UJf1f
qvcapY45KFdWtj3FynOQJCStHLntdp9DDwAiT9p1+pMlLRYqScv9q37taRtXEt3YCfA/a2Zs6P8y
8HQ1jeSH9dcj/VNtVtBTSGBkV9GS9Du64rEEwA219K5kSri+aZ8puFUeP+JpgL/qTS6CNvHgrlcJ
rJSW2nSYBntVYr2LVn84MQ2IuV/AQD/mUpn1usIQ1mBLpeKDLBk1o7AOJ/LabfS5aAH7VLDemoro
wVocObOSFobmFV8Jop/G/lucNX9+cibm4Ol4FfYGUAfzMT1gVV0iL/9Fm40qbYeJ/hV4IT0Omq4Q
Y2BWjC0TlcVpXkgeQO2mNX3V3MEpwieDDuxFr7Bffu5O0GXKDmKiclDiGQ2+7B2O1cxL8wAl1Vr5
0VvsJUvFHrthRwMgRWASv0aH+lRO71Kj1aMMJF8zQfs6KW8oCVVhhh1Vk3Ok2fjvOFepTVDoLaD6
b9Uyv29m0J8uJCho34hmuISyJV4uWFNw11snDg+VimtC38G4zEb0BIVy8JfjxBTzndVdi3pPPrTL
IpIGChx8SciZxuK1M6P7rDBd3vYsSgzH5bQ6tWDnBiMZbbDUx8o9Y5kokFS35Spuyf4yelhDu41Z
Z4S+rTJx1tde83NEdCNLSUUetR2gr9/Lq7ikm0X7liZp5eIZA6mDZ8g2v1nKZ//7tlSgfSjlO2lp
dCYJWhPUXQNfFVQbM7B6dzAa8LyZA52vWS1bQ0yW134Mr1kuQv3fINBOQC632NBZPCtfR1rNU7rW
+iG0Zpyekl6XXvcuTyzZAaBOMg+jarTlBvX43ovvWD0u7WRnNvUe9+ao7YI2VelRBREJ0Q8HxHY0
JjWCh/dL+UxJ9qSOVYkNAJT+LAmuT8tXrBCY2feQPWXrLCRkkeWQpdgbTcbpP/XPQClKphRPMCAE
DMipsUixT5CuJovOaCAJFa0aG6KqkP/mUAg5UmhOgy4oeFgjfp6Sr7T3VM4/mTY9kDGcjYwF1tcY
GfFR6ZotGmNnDu5WMbuVXrYen9SoK6ywFI7YU6Rc+LlExXKUWlU/Sh9i0F77Qzx0XS425971QPZX
fUpW1whXkNkucadIXp4SzDNArLrKMFdMMXH1teETvkZQgVwonowfrNZhSs/XcmEE0QdVZOZjzueL
GEfUbqNSVipzAygQUr6BcGe9JFKKcQ9/zpDogB+L/0EoDY65n6znTsm9TlPjc7mcu66pPla7Eosi
aqwqwjSqaqw2Gwli1YMwyMEJDamydXsbaMZUULmwmPJV4jh1arGDFdlroD3SxLSVv+bU1YzTX8rW
YbItxVap/ss4+0Tl9x5oTN9UBbDK1TWOoSRsso4rtXDKhWoewLbGjc0Lbl0byzfV92+kZzxHm6B2
sbiCVThYAdIvpndgXFlPErC1raD//U7lHw6Wnm+taX57nQITqIpMtvK5EES/5JT5Zi+olrYvZYsN
aGXqKPA7tL0ljgVwZav2MbNqNHI0IG35Uirm3oVyvrHLWZiBwokVp6Xb2BLFpMgiawA2Wo3VS/YU
Qzrq1Kiv4MQu8csSJiJ5thW6HD7zFEGn2L9WUfguKYXKcWdvzGvQM9EP0kwTxW7OXAFsyQbnwLH7
Ebni56TbGaqAon1xmjMX5iz/K4OFZA3s1LUGd5CRWxkwY6a5xJNdrg1yLCAic2R7W0c8OzbNqqV+
Xr8wiJyqkj6SXp87NFPMzh6ncC2CnVtJwg0bUDub/EPDeyqhqnKjS2gF//rNlvBtzOCGlzNqME6O
bOWuzV+JUbHqwhZfqQaMNuhKFrsTFl7ZcVpNmju04/LOoNt4aMPUZ9U/5rgQ373owKHxio05AuK6
2lbJu3uvzqteoiocrVgHj1ijLMbmZLJE5SqSh1tYPpwRk5LJ7rWgb7pKAn9xXbWJcoHqr9VgakOm
a+cIjZ565ycn4KbPRKKxFhagebTM0KwKsMbnzOqkTx0ku9F3HLXPetMh0LQhyA0sH7SW+VpuTmeV
rBsKbB9KBskStzu0+2jO+gKtRV6zdlNEdHeNGXj+/aZXaxX3AIbxnUCen/TbV83lKUMCX2asiKTD
EuUOwi+Eej/Wruf8O9yj5Xy1kxRW2n2Al/ENWJAWmUtIrKy6ZLAMjYRhViW+zBMeCefEF+PWwZNP
CZvN3DHvIfTHLNLhXxPchx2mLUhk/nCBg7dubU3k32KM1OtAi3KcOhxrn2ufA6TZ808mGWmlV4UY
etC8Qo/mQzoxBbyV9ZrfG8AkmwUXnol8pxI+6AlST3R1tCznAUR2oYiw6uACRdYhgroOyGV/Prex
V6f8KztT55C8F5LVIJPj7fTWGyxHyTEF5JUeaWUvnFp4DEeFddeFl3K2tZccomiguNPPwDO23P5a
4AvWW6Vd30BCO22uADxeh3Ajd25lQBhwjtZOi3G3B/+PKxA1hV7JrC/Ok62JS3LMCtzPKAaohBPB
OX26iX22AXKQAyk08+OpEjHnXI5LgBgXei17Ad16n8l+R0hZvs74eRQUPeMhcK9ZhPLV6P5VoKhf
aXotX+3YmEcWaasn7AO5uY3nNU31RRKWjA9cqJX3kCbnrWVoIC38Q1c4kvjuidzbGQ7w2nfHy9bZ
uRAHFW20rjZhw+Bfdcvz94+Yrea690Jjz8sBnPrUBlha+szStTRNpaG6uKTqZUlIdUKj60ckWd9G
iAj8qV7Jd5vKffUO+rwTybX1ys/kGavG7TTnwWdcN71RmUZoOpvkyafIAKE8oD0SAatdU2kpugs3
p5Tz/yxR/EdtFGhA/8TBhVRauOpNx89K6FeJweKJlilmYjRIB4HvuMFT8K3QvhUAYl/7zSbyQ5nV
v0Pucc+I7Rhslq+BkS5vuyk+B3h2Wml7Xd70lB8QTfajr1Iwu5RghtQ7DU90Oslia12pH+j+Mtlb
8GDOfcWHI4Iwe61lHAmZ8OWVaPZqxIOpCjbB/0qDo0bCUah/x02C6yNMP6+6OXTMVD9V9W4UdVXH
ZxEbvwZh3bBZhtv/16IwJzHINIGF95/LHJB4iGlQN6WSBB4sS6x2qkwPQmyKwfaG2mzE3Oj7Z792
gqH7wd5sDRSN/tFaRB4aSf0H4Fruxzz4DLqkxVfrQrlyEjO/DD5+qxb6M7a1kDvVOcHfe/uqqvIW
V+YFe+I0h4FIszOhrxT28WpmGg8FgKyStx49CbQBdriwj/syCuMabk2q/GdK8IPnhCiWZrFLOJlq
qVrw+El9uxux/6XpgOhPhgE6tM7MhrEAcrjSCvEoTfIuZWiCxLY7zqqzkFwWVN17L1JxCvHEdZMQ
PHgxpDRHGrPHFOKnz5s1iniMct/8PhlYB82QBPgedOhNX4wAdCeU14kxBVAeqW3y7jcm7BbtEIJg
ZRTjBocs1ptFOQLXPVc3HRB4Yh+6llkqKxafl4/q+E+seEMRZ2LAc1POM7YKr23KX6UsPdtvzROr
Z2iLYXWvY9AECXukw2mnrDLqoMaXi/bCH675eDhU1EJAlbgUSX9kwfAmDgknt0cnfTfYjRc/YsXq
njdzLWPyPdFcEGmONL+maxdcxuy78ndQINpMFDoQ4rz5Xr1BgjmVDqJ5FWR5BsDnhAHAIGpVUuav
pf60+A96Dvp6A/iEKXpfO0o6i5SxNxeCPCtT71dcG0eW9VzZPnZu7Ncuq982oOfnJFSDoBYlQ0Jr
5oFNuM3RtFeOj3PKOVM8S7IQD203piJ7t6QrfZHnnQV/EfCe1T6X9aDvMRI8rM7NeV75vKRsFDfq
hvdJEAO7nvtj2syh4laBlsCN/3/eLSNI2qf/9JsphChs4wiE7ouZva0kETVsw1MZck6i9k1JPG/t
Wv75ZfEGZUEA8qoE4S5rM3+7yUPPXnoVqLT7L3UH9Ibn2kP38BNJkiiM/amLQgMsUNPeDMdKuCaj
sr8YpuQU1MNw+yvK5KkNOjDkqEWXVt8kSflKxPT0buG4jbwwCmNrrb5ukE2goej8exnPC8fSMl2n
oP5kID9FwRVbhVZf+kGo8EZ4TIifzENWKhoR16cqDeMD4caWS7WNR0zaUNX2tnT6ZEP/+eJHImc7
KB+SPjlc9K22Zsloo64wOXfLs/o5AN9Htj6XvrDow11D99Hx57rWNKZUbkEMhEw8AFmYSYPku049
NkkcsK1KQs1e3tEiP6zTp2LxPlwQ2KDzs2kS0SjHtGJzwxNkZz79/XOFOrAhkGwEKjmi5DIgZ/Sr
YhmAFzDzzK3hv2ZchGAvNE5iYWa/XmSMzqbv30MU/QqaSSDwIwwEESFE+EIhUbeuUuevifANwmo4
6PRjlvozHU1SJq5GpfSdJKSiP4Un+zUnoKCFFpQXIRe3P72aivwuPU0rA+/RzmWQqLkE2+saKYAw
qYSPl1IkMGVnlCR+xiv8kZKxoMbKxVBQbwlO0bkj0kiAFchxXu9xw/kbbNAt2QKaqrCpkNU2L2mI
DkI1nytM+chIgJp6bLz+HARw7lq7blAHuE3stIU+QJvYLuAEKsBcvsMp4b5+GcjG1/xq62ymdKG3
cMh+h60ohdkr9/OIDNtzmLbjRnR5PHTK8nl0+pJsB+sxs2tdNxqMUgqPN2OY5KJ+oUA1vK7NDHqd
gP333kQ1npi0/1BxNUEwUYKuHXYWbBq7P5EzR3u9RLAnSYD1s+5am2ly3px86Mbx5KAKZ8tceCHt
zW6QXKvRs7zfFzJrwImTAHn1l4Pq3+1DjoeweDSBnM6nE+axij2c6imGBZmlpj35VD7Q8xNnofFu
3nN7QyeuSuK9jnAoe5bShmRP1qEcB76Kj79z8wSzHaRUkIak715VNrf4DniQMMaNPxX72FHLvCnx
0SmREqoGckW3woJY3SAFrluVQk0SKza0V7obOtGFRbdJg9br4E95G061Msbk1pd7g14Ay1JQj+mN
Skkd7aGkC2UmvQUsm8ZPpkHeqmev/NM0lT/xXVY9Hknd3V7Nn0Nsr6NS7SqH332vuA6hq4249RZe
XRF30ZGxwuXQB2wdz5UyifMagB4ht+fcLvGxCjxcaM3qI4ENE+KTifSuQxjIRN2APaLYdAwO8V6D
Wr6oaFZXdSj4KYzF8Kz76RlAgZbmpOqaF3fWQuXs4pVNSXq+M8wApqa4c8EYNBC+e4nwUoNkP5N1
eYTdJwcqV4xdb6yIE1OhJZwGWxIADT1LzgQJ9ogAmxpINtezql3YPMH7sYN4zm7eTyjOq5dl9tMH
VnQTqgMQK5Oht3NiSXer0c/ChPYGPrB5Q1LGbxfOu3elPvOUY8z4E69dADKH3miszpyWgO4+aDv1
K8f03VguC0Sf8DE2ynlvEeJZtHTrQVhbcpXn7xqVtuN64CK8c24NWcwS3ljZ7prSwpiWP/KXsqS2
diFuawRPa6LFaKObhTKkIT1KP2KeH+yHFpwQNVukqWkQL0oMruVgC+ToM9vWj3LNsi8KvwqdWa+4
/HmNXyNCpSRyJ3gUdgRPHohBaYDvw59tygNuZk592wwZBnM8/vPYQXdMtkv4ywt1D+sbfofV5nj0
fjtNMJ+0IWNzuC4JFXcPNmbxHw6XiHKNq21XJvzflc3ocvqFA/d7mA/bXa1dy50dRFvyBUmUjz12
0+43LoYINRrkO2BXzI0swEqsTlLF4cgetJExLwVD+S35WkRX+T030fBY0Ans1g7Phbc2AwFYBTuC
r/peeh2bsx53U6Oyr6xokcqXp9EN57UJwkd5mjJ7JHApX2j1uDmWiqb8e7Og2YT/4P9jOBIEksMa
FRF2iR1bz4c6GFQ7vbJOowiOgnFRT5l9b6cMJdIQ/UOqAgDEQVB2ZNTcHrXVZJUsN64XbaL45G3B
5fJdncrLrUG/O8pjNW1CqLTeLOQ9A2jPHSY+o6lUC9cRDshxju3/hh1DKN0hR2RSA7hdsXBmJn48
uRlRA6f2fkfGiIqMg4Ibw7Gs2zQ9LIShcaz0/6Gj6aq6V5RSJKMYdv5ZA1BkC4NBuikpUgkGaXn9
WGq7Kja/j3tdm9pnxEmKMIhzClL2jsvD6wM7T/JHEHVrY5IoIJGxeky20sI5OQaM86PDQf30U1u4
p593z4Gb38rOT+mNet/QsO6pL8wUyCQzSV2SZ9RALHRgWJfYUZNfLV78csdLGqqSAB8h2g3zzf6/
37H5+OGsQ3mKahzSBBP/KGmnJJ1XAeOloCnCCSZnH+MZSBTEfxFiWtl3BN+r3RSrg9Czq3xTXLhi
V8LW8JoOnWTZ3cdmwzEB+UKpZVWyH8iVucxyqhZw/t3fusxkkzeHSArWfw/vbiX9TvGO5f60/nC8
rCYgOI3kyaEy85Gq62mG3Tj6dCTINxSLE7g0lTar9pmeK/kP8W2n28honBFn3Nkc2EH3+g0C5a9T
f3SUygicuUTlWMIT6AISPrt2XNtVRm6lDIXILr2YoooZfDesVOC5Nyz9oOs3R3K7dkZrnOFQAe6B
yNSQdGhJrGJffLTrBKAotUClbk1K2QpxLDgW0JHVKUNxO8RRhP/tqLrOqSl5Rm5zuBUKfkZSY6Tz
6HeXV+l1VSvJNIx+heqzDXNTSNnkWDLvRUgurEfG3Ith29TVM002St8ac5DOL/7ql1ahHI2zlvje
sPb5lArUnCo6EIPPSY0EqCPskfOIdFwmdZAhhHg9eCXTwtr/WOE+gurQB21HCMttkOsI0j/BXHco
VpZu06cgSoLIlw4OUITBKu9F5LGk6wIGLiy26ycpxMtYRVzBvgBAdYZ0Kjb8u+bgurMVQCHsATAA
9psg6bR3wcEM7dezDQFbOf4P4SpgcFhY5coS4MgWlwRyd1L87jh9UGI7OkP6UAE4gTs+kuwJEljz
M4SozT71o8zqPeZUHcyPHaK/YthZ3VcZr7ZDtthLCi7NFy/XiFPcF6b5TqxMA5nsqKpe0+QKcmtn
nzjLb7dzhiskHAuO9Dyr9n4j1NMn/DZVnhfrCQ2NfgII/zvjOdUvqviOufe9itzVZLuFp48uz415
/UuelqIbBQe95SF9nvMvFSLYkq2D3FNrzv21VP4+f79SCgxvIVvbSY7CZPN2IUSyn4hHi5Ve6oOx
xcxWP7c9Qh0XN7XhdomydRnvfLTii8c4hADvcPcSUD7aVOU99zrrveh7UwK2nXNyYKpM2eFEVjVX
pXmPgfZiWMId+XoVUvENnm/7/hBLDRbvQR8p+lG3BPtn3gx8+4oIjR8TAhH/K4POioao4lv6pCtf
9/2rFHk3ZlSgWmr4FowUjH2PLUFkhHq6qlnfOACNSlxNqP+ITdET7HqTrFm/NXu5wErpgkkRPC1R
/3EQ68O7Q43oMQdPK/8bemcpM2wlmpWssC0kurJVjdOa6Vkp3PBWeM9i6rKbbf9SnRo/MMpZvS96
RAP1Ilonr7D6OoeAb2pRF2wl4plVZt81YB2U9Bxrt9yooNwGiFxrXzR/oLq4186mvpyQ/WyTpJVg
lMtgPrmQlGAKoAFiFk+xmlVL9smzGd61NiG1hkpriO5Xp4jupZNYbWNbjaCmo5Ff0je74K7D2UY7
rVvydrf4tGOKirclxa/aAfPWwdJSTN5VqgS5/mF1VGK211G47SxlcfsPk6vNImwFpKdruwvuCChr
JV0i7FLS/DEJaDU8F9zi+ekA3/45UnqwcKRr13hGufY7DTSa8YlqwE6DDs4wf0TJyyu7BUyHv4Ug
hqI7K5akkWIBacYzHQEf6kcmy6rUz4S+WvI6K250RnGhUjJuA6+fq89ru8Y5zL816NlgZMid7ZNJ
0RF772nfGPAzlNPfRn4bP9Ff/hCazeGEs8yBsen7aFcW/WbuduGn5ZmdkEZeHeTBSt8wCMRAOGan
tlPfDLhWhn5QaFrfTi2LtmxKqzjiHeQnKYXtm/wPNXaYkSwLbXIhu3P8QyUVR2jyjkpa5xOlEeW5
4MzI9VzZpe9FIPR1YymANQcFS0Gs6y3ZT6Bpvdgp2CPXTc+2MugVXxt7JibNysFWcfRm+7AHqyBr
o6H9ZmG5xYTo1JegcjuwHLT4+3UxHgMuljH3wMHphJXKjXZmtQDBW1x96RYyO3WjOjmmoD6c2fKP
Rn0K+S6vEGPMEHq1n3hMiiZTrbNUETDnYhM5Myllz5RDRVMdgz/eZrfITS4DVbgPvQdmmj9OjlKr
ZG/O+zClRN4MWjv6r/v0CjE11TqKKvwoiIwIAihCo+0zLAeSzITqTH6lZyx/kPnIuuR3NBkEPnCK
tKYCOY5i9UY4iwcYvYgryFlhSRMNsDXwR0I50JE5a1FTWuM3dS+rw0DhgkQLlUUMk+LPLURc4ejQ
kds4yrWfN80rFkcsIjR1M3tiyBBrY3QltfAFW7InY0roh1a5sj3NpNUqd0mLJU8k9WP58+37sA2S
qvZem21qWKddIbFE/qAtBXRwhK0Yl1I4Uos3itbkyDt7oz2QOC5hKXoccZYfQk1M6RovkTWJc+BR
/S9iwXSR2CedVA8kE+XsOEDjTsyV338xyjrWw3d0Oeo0gKPcLRhAXS5CvVDyRLTtwmiWT4YiBgCU
Q+DN0M9Nw4LmnJAYesQutoiKrEkfnCI3qcI3UBrteuHDE+n9+8yl1rCJfX3orGDo3BSe0lFTzxtF
l53vF8IuIIzmSjusvNBmWSauFv9IwgPyjgqOx6pDoOfcwZ2L52ewCvYMiEyxnkwcj268+scy0Cv4
PegBRrPJO9ZQvsFFkl9KW1xVGmZ4XBIun0PRuAL9tJwGzOClT5wLXANQo4+fEDEiTQJrB4WD+UHs
bcbap9NjIhYeHmjjXm3ExB20A2pht0AlsAuQgMv2zuZeplmPCNMr001KyYsLJjAKyDKFe/zz0pPf
3kanLX9aA0Hi31ly2tOv5wSEWLIq/+XVr8xp6vTPlXdzvHyjD19G/FFZ2LM3JQDKpMgzjjXciLFW
BpmLfvl9ZOpc0P9ksRpk7nuBmwPW9E4d2QuaWBw8TykQp3Ilm4NMMquB8ct0zZCiMzEfTh3bdBLu
y8HfU9kBGUknluzgtXGQqfIXkZEUAuTo4DtpHrgtr4SSawrFjkJvEYZ7oS9oz+AFOQR9bBljEUdE
k+U/WO2UeUAp14LbaelNeWRPATWKU4mgx13fRfc/sQIsaJz2NxjgamT9zkFHQ/MZ/ILEKNiLD1vK
rW1UoYSKlGxPio/e79tjzzF2bvR9KX8lzxxqTgr81ra19PnZMUAsXZRIoHMdUXSsdMm69S2z16BB
5tHSK9vApAQ6yVf5dF8f8geUyCmNER/piPIYqt4e15liqf9BB+G4814QNRqBEd5lMnUoeNPkc9pM
aE132qBm2zW+E5EwFujWZUBqVYZ8cbxooJfGC1lKLIGZ9qC6kMInidMJ+g1oiEzzZldvt4//HYdp
HJynBMQbO/LHrrb0QyVMrrRqk5xAz7ttpUQimodKESxjoumMqsd+X2lSdzKMMRSaOnXYPOQGqwIF
lcqGo18iG1c2no5RbLyvAIQOuztTP7C7yE4tadgv5fRBdiqi+00hfPunMeLPpbjqEFDkziie1mPe
jvS8HGZt+gHVE+ClGMjfk/3VBqN1EnIsbzt4QwaT3rXNGu5LaeD5nA6W61nCeZsXBr/wy5y4G3a6
jIIoT7K4yOUeXKFtMlZkhnlAS+cT3pAhjn5pSg4WAaokE44wlShN+ROLHCWOaU4ZK9PAUdnA7Fs6
sJ7m8kdgs1iDn4OKGiZW6DbdhHav7hApMjKmhO9nGVZpQlIdt4o6iOKUoJ9RUU1cjIX8wGNMZsrJ
TaOgrDdIOGxyMAN/jc8zBuhQ8sK1LgeeLbQnOTn7U39cpFRa5uVTJKWGbh9v6fPRGUpquL8uG+pf
FmfoDzmcDPdKqCti8QEViuGMZrtam7zIqGGkKax4krdIOE6vgLQPvSzZhdmte1YGEKflicz/g7wA
U9Y9A1/ITZOvV6R+RiMcTU2LU8k/aztV5Ipn+WPsg/iOI4zW9+r7YEBUikUMdiMuS1H/Alic7Xzn
4cmvKmP7z1Lvk4NpNBOYy+6vIen7k3IfFyouqZLMq9yQuZ75QUUb1vElwnzgu/EaY571erQHaVIc
oPUywmNuECgrR5WJjkqXlFls1X27A0JwGW+khFTTDiRpevLuJ++Ikv1SUHXPDVuq9LG4dNXuxScu
vkP4iIyDe7EBzHUVF5JvynivSBlHeOSB1wkXc2LA25ruhVgM21Iyt++49GsxKo1Q/ett1nGtK10Q
iMdnCC3P67Lfx9fiCT1Inp3/sy2bYdR2B/baOWyoqzTohyGUSJGLA2oaEZ2KJDWCqr8uVfbs2L3y
2H9D6ZJpuY33CaYgyLyyrUf6FX4RWFeMVXFWi36KfJutFyMbO2p8Z6hLmo+HKa4x4XgVGpHT7Wdm
JC3g3GMs6ANAmhBI7U4df42FgvX9oYaVQyEcI8NLBUQFdYrEk6iyxGMsEz+dGxIz+I63sM1bm9L6
AgCrgpLiKLT2S2TAvDSbMelw0R0gtZLpjsZVQ6eSR+XeEg7gqJc1WmwrCeIJuyi1/WkmPdhOhd2j
FrV26jyzQ3RxRwAn/U1oQ9Q9QvejpfUKZPVeu5YTPr5J+SE1JJVFQUZlP4frqAkzA29D7znlRaIG
IHi9W8yCqCrdnnwmkIk80CqUoPle9BfsuZAK8r3Yd24i5lpdjtXckQgINyqXbO2R+efkKWHBnjal
e0PmmAw1sMhNhzyuv90ubN/U6bU/cO9DFhJMqwiZztd0Ww//y1OKtgaAvZEIsvjuWCjrrtp3MUjT
zbooAHs4UxS87VhYggPzNGsnPqqLxPWWYG/liCUlSLzcB+NZ8vyHA1JdD4bQL/iDMC9g5TVIaD6j
xUnBO8BedLk6GbZ4XkN29TlwqtkgtxLIGOS28bl7P2eW4FM9Nlk+T7uoq2YW29M2+ysbxpVJ1kD1
KCp53pPE2Qm+3jwIUpSDhrkbCZXk0bWJfQfdjceb3CvUSPjlka5cycXEIVYy7tpMXlRjs8Ya8lkM
gIsVHUdRM9iPpXPUjRtQsOrPPtDlwV5tMokgmz/0W8n1hvqVtqY4C/8hGnkxpwgFLzT6aIaWAb4i
d9/E6DxmnVzKYCvN0qT8EC81tu/PQXJoYLkXaROE8dywVv1aD8HpUzcpWTNHOUv/4KRWVm/cDLDT
vlCJLCvju7YNvYrlbuNmpYWIi0FAwJDKegYhKdW/x2NCLaGU8GKSuau+gwBL+a1lQF/IBABuLOeV
NseAY0OzzFaWajKpnaV2KJbBmkJwXB7ztx/VgQ9taeTsRZZwwqoon4oxbmNMH+FyBzvMByXTlKL6
tq/a9piVkzDMnpJ5HI/c5F1GU4knyPkGiCkCM7tvLIHNxbckoKrXNLcSlxGSJ9bqd9OJNfmxwvPs
2rYD11OuVfOK0LhKeYG2pTKvZm9u6M+Cr5QNG0SF48WRlw+5uwa4KT0qYlBohPGwzljl8WLUHbPd
i8VNxA2DB1q/TZFhRoKB7R/QsvFmgYPp8ZeKGfJsLXGO9xyRofO7keyufj1afQZ1LgV1DAFt3qJs
ch5194vueBSaNBrmU8CKu4ZgWCcky+XbZ9YswA8xoF0P5nT+aOwSBGpbiUrp+p4GwCEPfPZ3t/Eu
d5mTVn61RKYjOH3bPi+Dvh3zk6iqROlqUAUuJ/u4s+2ERX1kXjNRYEaCy1mqrehOGYTUGM+bDWhl
xIRcME96m7Zd2E8FHaGb641kCghnSx00+tSav/X5ooC+ahqegy+UgDyIycbdyKdRR1vHNydcWrVg
GJrCqj+Z2xu9gZwHN1mZ+qdMh4Pf5bl/IFLLNBIf3Mjgm+fdpy43Rj4WLFFU4xFoBRgv80gdyBdi
sj4D7HrGu9TRfVdrvKl2ZU2CG5ZP8Jkn1WR7YPtAdBCYWjeVr73xNeamd9CV5z8AbZmxJWX3UiHy
BvMYsCpb9Z12fMAe4EP1y/ryaOYAFkzbvGdpN02LzdngpRcwEwMqXjM4iK018XWmMSTOYT7as2GK
B6WGT4NnU6czyLuKbHy18heIrChK7NHLOA9+mEbM5zBM1z86/3wpCAB76Pwk9kwyK9ZJivHrBUvR
SlB2O5D/hNMdCRyWkyA++FfGh/cLyOkxUf+PwPJcRwcYYzi3oxV/i7uZhJCSzgBM9qxjEiwRmriH
Ei6fw82EzH9GX99wgX0/imEAUF1ItW2M4o1OOhwzex3W8PaqffwAbA/XJlrCyOluZhwu9X5TbR7H
BLoJSPv4hdXv+3YxMfWKPS+S6f+eNV9wnvJ8tDIQxnQS5sZI5L6FRnQNjPjbn3SxbSu8QOv86xoD
zvWMpKLduGoUrMinAAsrv4aG65dbSNx5wLXZ3FLi2h2I0w/ojddwwKjN7buZs/WSCI/+NJDkEhkE
yEqVr7T8rPonxOtKSyIKCwNdEwIIFCzUKW+7vY0dIRTtlBa7NvtaOxkvv6lnbQs5kZ625c52K3Eu
5PUTb96Zd6xk/Iq1YVUJOxNw8Y23l8vwDC+WaAKpqhPx5d4k8OGA8r+8GqctJXFOVkHX9NxD5VtZ
Jco1QSHrU8Z6n3U8fu/oipYsWnZUerlFPoa4j2dVzSjq3fjFC0YbBEOcdXxO9Vq3yt5sz9PVjDz2
hvSpY70Tzj7bf70AfyoaZe15pqAvMdVSms/0qv3/wNQVnq25f+ACnUJhUalFDAtNeb7uxc5zGmS9
MZlVjpsGktRujCxFNy8G/jRSPLjYAIfFC/ZuwLzhoctxwkaiIm5ShNMtiVaWXmTAcVTK9FlhgzeP
ijaTbI5rHOkh1uoYe4VjicZydkq5iLIWsAsvl2j8e/Bylrza6+lJ4QzZS5LrP0DFmGHBv2Ybfhvi
kY5ifrMlHQnA0uuo4T8rd8t2orYdUv/qTr5mEjqOP83mWHPoGgGPVQ7AUjdGcYK9GmG8uo2dHch8
9utM4vJeoYWTMgsbMtVUMd9Sy/zm3a25HSjd368tmpAo6XcVoxqrh7XxO/h0kjk3i60sKP+gyMMG
zpPjXPmfMrr/YY2mAb0HGlCKVnAxj0pkZPf7mSObOg7jdfBVlpiMjws5rfYmzvGIkcwa82wswR7j
MAEwG7AxegQTjqflSImC+ldzZ78nvK1K2FPpQKb5FZxuLtCzYwOcKcGUS8jhv+J6qa3fHCK1bA2P
MLhH21vtdWhYzEzzLlUOMZ37PBjW9gI3TY5MDFvKWMLevDWpSp4+9lFm26COemdCQoTWqNOe45UQ
OPfVe85iTlSGx+3/cvVBGNnWLRW+wJOCOa4HEy0LMoLsalMe8ptRDj2tsGEb8NW+FIqttnx6dBiG
lBGfLFS6O6OkJQS/4u1GTb57y0zdLW4YoxNiMELE0UJD08RtSHU595K1u+7bOSOFf+TnE+WjzZqZ
Nb4bMYbwXeLalt1zhOjFUqLD2Aa95kwCKSA1nCCX9rBz2wQMWxBSYQ2SaMUsMAWYCJjU5HS4vOqo
irSIHIEmgKOw2LWLz4z4rNUvL/YVd9sX9CGDhg5FpeW201q6WO9vbg85EmeiEHNqaEcIWFLHOMwz
0pf2PA/2nfsEYSQ/4fr4W+FPdJxH4Ffbln78SbSB3O/+k/l+HT4nP33oennyYCKTD6iVZsHq4luG
/O8tI6D/2HWf3HkKtfLJKfeNUMbRFExXDHJuAULhobN/31HVgFHlJ8DBPjzw5u9WPViGKRrAozht
/S3DTNYtNifDt8NuIPqKPqD0hxeY1MMSrQjoWKSTrKlng1QxbN1ulBR9mrJLIgJ+XeU2d6mN70DW
a6Xbfm6IzSmt/2hffMiWSu/d0bx6hHKDNGsO9Up7LnXqWLleLTvxAiomIChH12/TBm6ybbCCLPUT
U73EO9UWRpZqToiaM8+3OBGXsV3nf4UAeQmWIwYbTN89+lpeUIqPFqvA9JXgrDNK6Q6bVGw1NEzR
0og7099GRrAWNapKpHjKBLWnh0UPo0QmPeEXvAaGGORmwuB6KIDk0lHf4uMWpTVwCzA2yayIavIH
/AINWk5WQKgYcyvnxwg0+kjEE3UweEdhIGNRzZ1t8QtZd2qRPvOccXmgGfbkp9glaf/WKu61dwKo
F1n4b8vqrnsxvIhFeZTCTXRzJAISHD0jMu14bpPzmGV0OaB+Gekr3mG+qoNzHnFrEOXA5+gWmkwN
DVmLFapQtSN2fbLOWmQE6wsHHzH87YpTBs+32yo/tY09ImWPNURLepvepZT+kS7KAL6LG7EFAtJ1
hZ0e1JSOwBbdFJH/U1ZX8vyiRGXyxJAUFKl4XC3xmeZ/6oLB0R1x04GAectKh6Gnnpw0092JJm03
FresNdzzhtPpv/KYbUFnMy9+cVE/5ryf4CPgltkCjzMlNqaek6H7iuk5gLYrZwft2VkxT2hgEI2W
dN/RMZPwvTlvRgry2wWZb/TiLCiUdZWMWEnAv/EvpIEiWa9i64hTu48Y05tKNpt8qFwdz4zc6kof
InEVVOCoP++S2c+H0ALQZdQDzwtGq4D/3H2+PlgMN8JD2/YC381MYvTnMbelh/mBvhtEdwl8zWlS
xLRzsrjMg0nxrNQN4XkZLLuf1dS7mBklSR4MEm7Bs6wjjGwsSYIkN7pmMwF3M0ui15ffoxrLaRgL
4vx+f5xEPHZQlp/tXagHDCgQr7ovUXT+tFMDQ2TfUmHlgDDQbHnHdOdhcwzdEb0AtBfMQDIzkVIw
3pLOV0pXq8wgnHjQDxEhSrUJRI52Ctwb3BTuPDmPbOTfIHJY/6j+op3xCv0Z36bZoTChnKnCnhLm
qcjjLXU4r3vGAGHJ0u1xNiCSsAyuymx8rGsL1Y/+IDPI81osWCGNBtOUCCUsw6QhrIpBjh5jtJcp
+p34/Ph+u6kB/0q/Rl28DsaflP0DlgAtIIw3NJgLAmphiKzyGzeImXja5bk3VJeLSbZD+H8f05vT
AfygPVgSYdcm97AIhhylv79l0sZ+ZIYbgvKyDMWVe774VIwy7wf+RN0Yr4iMYwhb6S3qRX4ivyEX
k5hhJSaZAqoRnS0i8avHrR7UyZlNvEX9pxv9cYBU2/FSxy+ogQ+bW0yrHNUKqW3Iy13g11qb0ct1
anGq08yXsk5qgtELbG0d5v+fXMakQJeAxiZir5fUbEuOYTI+qkeLhctFTnGUCVOKbBMRu4h3xojI
UkGLsthnCw42tF6TS/Z+CTJu9PsrRSFJOdQ1HYgOdUWTlR0iSj4jDXSTnBm0X/2liRRIX+qgrR2s
t9cs532FlcHfmOBXNRrsTwBIEgwGJi2QsTHXLxntSE33pxFfdynv/OoWo8XbjzjwoAPkhS8mtMBg
kxkeA7FwRwYQDDOxdFlMfcx5zdPYS4eT9HeCbHeJjNGv1F35XBGj/rRfDqBuht+ZR4pgWfxD8g6I
VO4WzXNd+QxNUhvmdLIFAjKqE7wtVMlbTivuQAcfQsCKrq9MV4TTH9M9IUsjHYXi+xus3y3LIr+j
mQRy171GEFFrbcjsmE30V55WutB92u4R6+HFJg/XzcRFszSOwo7p+YEMM6mA1H5CuEJNqvUHvP8p
xibqaYxsFv2wu2DpRxVQQq9WQ8V4Q2NlLSFE84CLfEE/ScsncD0g78w+YWiRKtinE888yM/dnMOG
zDxHHDDzgSdqVEYfflMh7dMpKFNG0nG+drhTndOM29Lbw/YuiranralYuoEtiybjqO/+mH/2vqBa
aizVL+uVelzsVIRodANTUULOrnXmQIDsdFWgX06Db7PxktLCTWfjUrgQacjwk7HDAjQkIHcdjdEu
MePk08ucROqGXHcCYrCaWrT+QJaUDKAQKppX6C8pGVDtPIG0Cucne/K7BtG7BXBtJPysWxeR6Zf6
aDxu420WSs1GPV27slfSw9OKF4A8WsT+7UG2PSKzpvYjtZTNMOf8p3gBtg4dHMwMJqYYao072JDh
akOPCj9buWT22SuvQEjtLNk2eq03CVq/eC5IPMGCMzmdxfanLtabBiD0VmF6FI55mV8BA7Qa1sU5
uDrX0ITtNBsS8iMfolb3WDWzS4KHTx/4LJvi5hXoNmLcNVTLTsAr0IdL2Wfn7zRiE9+0kr2arIfj
IYG9y1RCZ1B6g5X0r0r+68Ifsxru/4BXUcPm+gqO7Idi+ziSrpgBxLiqb4cr2KNKnC53qHasv+km
vM9cdpXCeF/kV5xjHzMXPp+Yu9kSqrio9ZaB7d769Mf7TCpsy7r1oFxjerlOqgRrZz+lD/lY80jm
oibj0BO5U1LFTqnTWSroqDep33cv/m1dyT6sPEpoBxFTEoNhE9/ysX1WIbu+9GCjZTeW6tuM/P10
pl5fqEoU/YZEVzR/IwnzRVrSRoOHB6lV/YTYyBYuI0njExtJhLNhY/xrcC3CPuTpUGRHWM+41Tq6
2D4bBkzu6g3vNEIapm6BkOoBxQn0RtsB65ICZqRfuF4Kznn/xRp0rHNMuR23IL8PlJdHgd8llQs6
0Gz2g4qXXprhJJpVeyYL4j7iPb7psr2Lstq9ODfdO1cAbK3EXIGImOen7u8zvmKH23GSkQG3pMQl
EM1iAEdHDQRQREXcjMRI/SplRthFR260LtqSuec3yE+UQI70tYHY2T+1AiJnixNXpt+3cE5RXihx
FfMg4dymK94eMJadPwKm5GAyGtXEn3lvuUsIeL4eh8IkjyxJu12PiAZzeOZyvfWzRElNW//TJXE9
R64sXk7mfcMW7gtIuDqWCPY/OBUlGfGsxsKAjpFeIQHIctRyDy+V3w05fKF3DvK9uhXFyAXhNc5d
SiJpEwgA+q4G6EO0VycM63i7Tzd1OpXHKMuyG7EkCyAf4mLXxQQMVdQM0Is/GYxXzQSiwuwNtV1A
LIDcSRKaRZvGApGeeCsw0R8Ba4VpW308ogGzLiJSPI4AXAwjKznEYcduEYekuOWfhE6QILK+/i6u
c/pcX/iRU8HJmyB/Sadi74xHZW/J+b+mEsnBy1sizsSJ0YbAqJ21g6+ou/YQEjQnLzP0499lD7wi
zoRLvUVuCTT4wCky5KOimfbuVjimMVjkmMW7WFLVWp/gjElXn4g0G5EIAi1ZqBlpcctcMTPauPxs
EC92kcx8VSmCXBsUGX4G6Mdy1OER14Dcq1IpG5Yl9fAgzwZwCtqM72jA2jNLWCtpNDvm9leWZLr2
m0Op6gwBb3eam9JxCj5u2C3VXaBa7cTM/qqwQS7Ro+e25e1H3HqLJIQfJaWzMFxKN50pYhJwtJRX
kNiLhP6gqXf4i2rHHfWEM78ZQM2aPdVHM56ySIiOi9LV9Oznn0bp0Js0BKa9MlTnWu9xP3mScUps
s9oKi2Bs919g3iQ0GvVvTqBXvhMN7vXFXe5ZbKg/HD7kb8TYWRyV5yK+s60tKJOXNR/Pj0Si0SzG
vA7i8ZkdVsDeT82HozquIVTF1DzwAkCzVXr+/f2DQ99iDbv07Ui6G8Uidp8Ah1mMKJ9ASpshTJcU
ZxRVEzk3YgQ7T+lSc+H42IWpDcaNNbUSh6KZ+9ObOItGjc5W/aJkqjvvw+AgSwB0wmWyVBOYsfJd
zoavYh9TZN5LQnltcjg11IaL3i45XoatFfs0yQ2tLPPoHAc/2BPMVeGvTWOHMLc+sYtD6/O3skV7
pBx/lqxRNE5O2th1+X8MEugza9rMqQ1q/i0D1MD4/TVF3MBoZchZs90fv8NzW91u3hftquM78Y66
GqkU2hAyR+V1dMe21WuYfwViUyPth3qVOeAuxQ0BQNAh+lZU3S29Rek9ymRI7VMMUU+VsWdfkt16
yZBKU3xEv1SogsgFDiEWd0sLdNhZKgSrFzEHqIAR6z7YStl4JW1w4lUahL41b2PZbb1PBBiLdOPh
wp0Q9JEIZDM0xdkSWnPdKgsopgjc+N0zP5w8BAsbJr0JzqBAKpP4bkbt6j9EOt0mBklAaJf4vPWU
dDhA0oI4mT+CMFqCgbwFvCkaWXifx/amQNry/7uRTMIK4v9EJVe8cC5fWIvYbFRgo7/VCbSn6dpf
PxFgdDUd2DRxHyMYu/0JOJeewwMRCLfj0vjZjzqsxq90JonwNNphMldOQ24VqzDhqbtqYy2vrQnv
hiME7iCY4EWYcv0dKrwwkwaKF39vLqWjIlBZgKMSHbLAJCSNrvFB7aJ23yz+pQ6FrP//DOWWIF6V
yS3HdGs7Q86Lb4nZUAY4RrvQTkE5kvaWhF7dVgTIyRMLUyRIqwO6E6vsqicLSsg7luCg8gJGVWJX
vab8/l/d8fv2xbh0tuqRo7bwm9fNyTzMlOlpZxl4Z6ORuw0lkzgQmvj0IQfXS662usbyREaD9EJb
bYpOJpsWHZ1lOgw9N19Qw/og3fbwtcKkwfTz8FZIzYdJSA4XrauPWLu2ZdjBYbdhw49D1SuVMd4k
RlHN/ykZfZIqbd6heqym0YKzasjHkFps1r/c0fe8O/ozq5L0q05dYZVchNaybR5N6Qsr2+DrbQgW
iPAsQHgFuP8RgQ60kt3tHRoGSVNMNPN8g3Wv7kVuAUr3quvt1G7ujTCkODd0M9YK2TLqVb63MrKn
AbCa+cW3wRUhdQ105vDpeKrMUbE6OnikrfC1Ed62dz8vhOwNZv1fp7anpPxrhZ90gS+ksZDLO6W1
HkMXj5lMDXTM49HmCmMaV2m6Uy6nmLlfZmtFIlmvidM3rYS1JrpOok0MqqZxGBPR8jVk2G/ntitY
BqNVO/08zMM7+QMmdf6aahqII069Rg4qaZnzcPgoxXza521rxPX5C+45HwbSMo0SBHg1E72DEilt
uGx5Hr5IRxAy/lUVLRkPtgsxHt0Fw1v2djukhrP68k6JHruvX4QSmZW+/Fwl9kA+/TtcU8FjEz2N
7tZahmuN8Vf68QXn6SCTTuO8JQJsKjMo4dvuD7i3UlBXwgjeDaVjAlPClaQty5IgGffA0YR+Fc8U
pCJXHOv196aoGRqe4bS+6omwzedtfQhyBrp19bctQXkq7oedq0Spe/aqltvUUjKTe2T2dWzArCzH
j5LocDK0vFLko1QhGVGZ+dpufNbwvda/6R6ZMM9+RU3qwCXBIuJHkYI8RPJ62X3ibDjGmCnWc2FC
j9DbBuzlNeWJCsiH6RvPUXv6L+Ac7ENBvya019zC/5Lr0J3wXck4p9aBdIaPSe4rHYUFwofvcAQs
g1pPfgj8sVN/cfhqpt+RbW8dft6Xgmip1kkzgFWpglWiwuiY/c896qZ1SQQOQbVQfBqZMXkuZqTE
/ODpH+xf+tdhaEzu+2Fy3Bujivb79ZMAe4rZ4vmG3TJWV69dHD2NEfZtkntllUTJcywTa1wPhC6O
PMSOsx69FpFEUus1QlTfbyyWs1pMD8J4eT3w3uUoA7CCsanqqlldaCFsnLSlYp7CaGkD+472A0EM
aNYITuaUDX/JftpFRNEbqn6FjicTf/uhM1RTsddkOx2cJC5igVEM5Knnfmlm30/iOSrC6SpKfTT6
VaM9a+NYitO7eitipejx6MhHvsOKVEQSV1RBGrLkKWV2Xk+eSdPGU4fzi9PyYPTDPBdo5yuCvRx0
9oKLXSq4luzojwJNzI77k3DaceP6uOfA/nVMSQ6fdCo5ZA7yNQNhvpPoXKLgqwfXPJqDZkK3KpGE
19ruwe5yyG3HS2E/UcclkM0NqZX2QNk5ZP4MYln3ciRKiNWm1JJ9FMm2+QT2qACv9eOLss7uAB7Y
5pGWHP4tGu4Bp7O2yC7K1mdz+6+tc5/LsEJRJPjzht0Ga5QD9bkmcA0MqmwQ2Zu9SgYIeB8xJii0
Fc+F1O9vGCD6ZG8oXP1J/Tj8GbUHM8X+nZVi1GB7liATZNHVuzHKJ8/yn8eq4O0+wwAkExB/ldpc
edPPCT3ErfS8oR9oB4EMr8R7/IBiWm0mcrLXz3PNAfxD4a0tgSOOdpflOGgJJU2JxWFFtzuzCPq6
b+wuoci5DuWErsqZZXA8rTU5edHWdHuUFAnwCaAJQ9z9/TFayx4MySpVdcPQhWytfwliDgxPdsEw
rChbjsHviZe5Hgt3CzcGNkeveYPqgfZXr+qBYyiKn0XUp9d095u8avhsrHhWimKEuWk8sEVjeE+Z
7JcWuCz104EuBPoBlCPsDeMK15EXOlDydqZFXGnzPKCRfTONibGXAa5FKvMvuRC40tzF0e3k0uMG
Ss0XB39E/dvNlwnOjOQ9y8mLz76dK1wjvxextG69GqrUrc+5VmGPQ52Zl5c/fIAqg3GNHEF046yZ
IeZMpxFehj9OKhO7N4l7gKWHFoznKnJAaxBOUjXmpC+LmmoDXdDqaHvDOZBD2RRd2AMvVhyKi/xV
iBULVCaxXzq0iBf9KU1QNoVrj5UExIiXwWE+6GMrTQeYGbqI8cWEQveYjTZy5AFFOwhAZBSPLDAu
rkX0xn3Pz1UErj1MwEFm23R2frLIRo+aLL0CRBjJYTwzrRJr+effwl6Fxx4TTb8tixrGvVF0RM4V
w2Iaj56V3crS3m7yrzKzNOp8sA2SI96xGBP2LMVZsAxntCNgRyXqvRvKvzeVXop7Chtsq4NgHPFY
kviY04uVJHbs1WUGzm4aokbTNEaMcJfC776Mzpeq/R+1ioZRDr5UOtvhZwHbyT5mtpV5T6byBYI1
mIEm9gLvsR+dBCg9t/P0UkLCG9BDSPPYmL7PpNfL8uDJYOvDppt48XgZqtjC1rX4vViON4qes9mt
1QBblFVkY9iLRJovkVm5COYzJ43FrS7P4btlzCFdWt1JYa6BWV/4x6SntfaCnK54Jb+iBjmRV5kU
qA+2Y4ZbMbNla9F0ciZKl2jfxm9r8xFu/QUql0ewvsnyCivsk3M8JtNqZpY7PM/DlTLEl0BElFr3
3jAUH47wAAf1A5/Og1sYZZ3pTQO56YFUWEYR+zouiLYc0ok/quh02/ylgLEHNf5OqwMqNO5nqmx/
YBC+OUvaxcOc2glLPLNiFfqZgf533GBkd83MqYVOx60Ju+84JUYk0YZmx71qZYrhhG3r21SniuHq
mPtlDISIGmndu+BOztvHBzCI1lH7HrDdVhmkIqWeNj4h0vMlEwJuyCoB7XS3Bnmz//0/Yh7+TB71
58v7Xd6TYFpPyk4rH9e49Mq6HxbqSvdLzIZYbhV/iaZKSSJfD74jlkAaE2SQuj2bGSUzZLy88oQL
JTZRdLlQSv9qfvLqVB02wgNAYsfYmLdYfQ9GUAW2GPO04mSyWEH5iL5N+nd4KxJqqgFe6JKXRcWf
zMuwmgIGSsnwLBmRnXIXQ/UZ1+/Y8JG+pJsZoPUCOrdowSvYVOhVefvnRkk/ORSgyJ5H6UkQjQXB
LHr1JHFdmJhKNv0vBI6caTZdYOtHyewe8BntZ48/Hlwy7r76D7G2szHbWdSyT9mApB4Vn4W4xiZ4
M6JZhTHvA0ZdnPmizCHJXCUQgEPFefJWRGMAPS2PgHRkWBirwd/DzkLOY/tFqiaOUDmAcgOQoEAk
yelVmrezwgRnJePg6Og/NYyWfJXP2vkWsHcmaN353L4K4piDWv1A27Brlf2xLtjfGu7QNqlmYg3O
ySFpdBw1vrywH8Rk74HjSlPg4cVhGn244holuDUiyPg2mbusf3QQmyP11XAPLvnZf4kkXpmri9Md
11nV6Sx56NNClQ3JbxBu8UlpECCAEwMepes095GKcE9ZwNJB/LAeElIMNm97Nn6GhXR9Jp4OUNfm
VjBODpCYx9sNqTrKTp6gwjil83Ev2hBDwgOQCtHuzkq5mIOb1K3Yk39L/wY1g8k1JBsuTKkEDtAw
KIMAvPMm0rLlTo4eitAHOiXtm+L87KbRm32O2vC3i0XpUL0vUAw9jL1PbOWkveHCjydD+tn1Y6aG
WA5gDFC3KKGgbccBITF4NFK/UDuDj0z93btQa28Gdwn8OygxNSX4/adVDupfrTmAEeiTv2r7GS/r
yp3IRxjquaJ5/iXEQHp3NP+IHwwn9bPHpEhngsYD/9GdBw8LREaqtZbIkYjFD6MDjmOJIfUk2EUf
C2Zb/Pw+qHLRwUJtVHJIwbwvmteTVMqIvG/dJfaJ0O7qNKW4Ekd9G84lxRS/AilZdPVUaKKW6vK4
AAJCqXckMyrwkXFxh9zOFFAfjlQ/3kELOPNhfPnmENVbWCIvGP0UrKMoR9E1KcZ0TRwwPT2uWQA2
urJtf9ZTOoS0cnTwtCWvyqu1CmKaw3BZ/tilui1345j7hATNXZ2eQbGpzUbwqcYelba5Y2JgBPjZ
Gtw/oVc/1MsEGcFf2Ac+Dth4LsYs9sBnOvfKtDgde86PM+b1x8XnFFMUQkx/MgDFCBoVYT8abyXg
H4iyCG59oxiy+Tr6Ke290LjP5ByHodNr5w7Fkqbt8JNY/VpXQI0gyNrWiAefaPtdGjkIJuiJqPjk
i4CCPR4NsrVxnIMxepOqz9Wl/iIl9/ftyg6KQFj8kOby2SiwuBIW4Q3PrgdAYk7wu6ChDfotwK8b
ZvH2dpCKVr59DzNXwLgYD8Q6LG3ZlkK3kLDEJMj/j262nYJ53gQERKrn3irZOJyZl5AjR5qyERBQ
t37t7GmUmNU1NfcRM6IG8P5/GaJL8d0vd5AR3rMuMoeh/r8vmuN8qB6MJtNyw954ikyCyM2u9Cs5
4X6FDWKK9VJl1hqGFGtztgtuMOTVMBF/BFgH7X4pKds21OkEhhtvPL1CqgRw6h0kz0h/Bp1Ec+4T
ka3jN78mGsO7UfqFmdx/IXBJcFsqpVGIsoGP6s5XoPcddSTvlVF5xgHPRN4Ek3M+QMDQNew92Yad
8KxstbVcKRWn1dOQ+ldP2Y5jUkBAoIF42y2CO5pPXh7OzvtDHq5sVuitm6JJuV3MKp62Ud+5SEuO
KmuEbGBk7PaA45eTgcBjxIT9/0enCUJ7IxxbbMlSo9E+cV7paFayel/7uBUvN1Cj5Gr5O1SqnfXx
545ahv9UoHe5nUB5eZWmf59nhc/zvfNH9BKCVf5T+jsM1mDT8lVxy/k8mDcgLRPfxh7PNSUJw8UN
vRxIKcRXZCmIpwwIh6cap/qZtuUhvJdE71xn6I/OJjhnyDFAEK6qiB7d+1CCiAGI78kKBkRG3FDg
j3GkCGVJmo9Vc06HHVCoTujRo9JvaKhrYPw9xGVw99nBvC8Z6UQO250Im4zIk6BS/vIkUPtjzJVQ
k8nWMTtszBKeGlmvqUP96QWEfCSRm6vw79gLPRqyxO5NKeeij/U4RMQOIhKuWDhE4oMgDy/cO0KZ
A/Xz+E4wQCNKi8oLf1C30ZKMD83yuJOaCb5oV2VP19b8nfS0yr1dm81jJKvJr4xRbh5IFPnHKE6J
cnr6wlnx4jb3JMFisIs0m/ACGFTGtoQGC9OXng/+cATFZJ39A+1hFX0fuVeW22RuyCSfI/hBQ8GH
XdqfkVzjsuWz+ctMQ6Cjj5loR7ZVh8TG5gH79NCVl2mqx+by4ccwOfXSOomh7wUwQmfsAW2iBcpR
iUYN1Z/m+HU6PcMywd+c5V5eVFLXAkHTxWeAVcyEt6Ts8K78rFlmyYei1tQZ1c7ykfwYTHKLpxqN
Mol4viPg+YwGNeEl9QLGOXvombhCggyQnHQBjYsliz7hR3UP48CSwCEEa6+XiSUnzfZDbRKBruNm
5sGHi6wsvqFVowzVUw6fbqA4JSpUZ/9yAjRXbeaAd5d0Xx+ZwdW+0FALGkNDqxYRrE+xCGj8u9SK
W7LK3K7PJlSx/lhipCby2jqu+O6lJ5OKdiHAa+N+bf8LWB0cWGgMxdKuyZZBOH5mgm3nZcLHaDj+
sOMj3ynnQMhEYCb4YFidvFSzntqqdzIeM6NkM+kXjLbTmmHT/CSFyud/3bRLaLbwEJSavHWV0fzZ
2s4d+mGoem/iH0fK4793oItOSQFwJ5T3OdddKKSBbEaUryd2/1Uvlkpdec6N+WjzsWgBTKAK68Er
mpAZf+PkfVIftyD4h5Qh8Q0GeuxCVTN05AB+A/OdkHnLv056aAUFWLCnU35o3EvTKnnpm5Xb3CUy
sNGqQT1+m9bush+MtxwU4TYu3fEXRBbJwq6o3fTZXPDDvKD0C1+z3m1CIv5cXLYYtchX4mUClE3s
sdUVeQFQGnihuN6y0rypnsxLzgEQuQDARoW1ar3xYBee4zjeR/WAxk4TTMPIZ+FtkPASHqOWSNgN
7mk1NuiCy/M52mfaCveFa5T/ZbuQJf/Gluhc0l1KxAE+EpKaL/nwXoxIW7aF9kFeLGQSLpJxI9YG
5+Y4tkGm6x5FRd4wNohH/ezuUqzlds+rot5XTWBtcA5YYGK6EPt0sTLtZYo6aysfuzH0O5DKABaZ
2rny+7T1Q09x+AXkTRE25UOrUh5AybV7+mbwUZA8tk2DduLox0muuXCz6B/1oi+7r0ELbJ8VuwYN
glCwa4weDAT9AjOvx0TbT/QnTCUfTImX6aCmilkD6g947zg5pFTjFd+tKHvn4BSlMuk6SuUGUNTL
dRTi+CbpJRs0d7XuJNYyUESVKS3cwtMBPA+4AqH3S4SomVQyJjAdshGJfnbn5uZwiL4v3FpdreEO
5kr/Y0GCGVVIRj0xXEW50122/eMh7phOdwFTZUV9geuKgnNsaCgLl7BTyP5ZCADbzJZkXEZLETNY
ejTWBzYB1uwCj4+9Mr1UXfMdm7O+DMGMr0whkpas8Cp1uCS0mzfpvl0y+LXvaQefdfVXIKO5MNWM
Wa9qAizyxzKVCHCBIvhWQnlHXmMdIrL7bqxWadH+spWXvVdcKfxRK+sjUBvR8fOq6ZSZLoOLr5X/
BNTrnJDtrHib30tfQbTZsDNDLhyJxDI8R+Ass7ZhG4SUAHgJVgn75C+qtqnmGkR3LVe/98/Vw8Ur
4mwGsvwug3rcq3vAlw1nSmvBxLTCV/z+YUJS+gFEmBTjqt/hOVAoxbXMzjSY07snTzyE/3mzDcfH
95y3J7gzfqbRyRfojhJVG3llqWFOXcwTyVTedja2POb5xZvUvFklSTGlfrlNaRVXLk35RoVn/0kr
rrRNS1jWfvzwxu8Z+V285xlUex+HzMl0InQmeQIdUIk9O3UmT46mlam44rznI2MAmRs7/LT6vlXY
/rNuwG+9gaEElJXC+rtZvVH8XQjiKYZnFPfCnYg6Nn96i0rcqIBY+GsgcHLv4WC2vxT0je/SpVDn
6KctBIpTrZkljed+WmJKPMu1k0uUCr1ZzqFBFtebib8SXa46tbsFKkTYL3Y5M3P95mjYuUyYdfwZ
5d3yEzhwg9uIpzYxxNF++ANrDM4dKGOWT/3TRWtitVZPbSAfD88+k2c7N45Y//GSb26AJ/8k43hv
/YD5sh3XSG4k3itfWTtzhV6Ez6DPa0So9Pv7kIbIHFNMWKDp+Dw5HBbVGxdOgEzJ+BkKvRSWPKmX
LjfrU55e2+m+cqfIJTNKy57SCfbkqV4s67IO1iR4DjBOk9F+35rdv3eMSdY+7EvR2FzKayA8AqkR
yzOGecEQqVGfzHYAuUaG0RZTt2Qw6X2jtA4CXTaY9/WOBOWt3vbbg7FBF5NS6MhZRwF/oNkRXKGW
VuyB7P2gT1Vu9v9B1JXBDuNeSTdZVM8FVyrAzTc8csqzdpOa3ZIsEYtoG548+NxlmVDB9l4JirEW
s1HpZGeTqKN7C0m/balshWgzcOWETC+v1vvf1freDxhKpVVYKaiIN5GKP8uebJ+uK6dhpRl2Xs9j
2sFJLLJP15vMx94Z+T3Lc3oKF1GfNDUe7rCV3PCSjt/ko62QtajbTPl4yhwnsq4SXMe96V6tLK36
K5Mc9ZHOysK9n+doH88rac05oS9sUwhb8t1AjpbOx6FSIZKl8AKnNJwWoBw0tKn2sVI7Ce1q+ybK
O4OJjC+TuG4DpdDXMCUUSgtQtvfZdKtRyZ2lBY4ut+eZxUY3ZDn//xyrFobDn0OVGawS3JWttPdL
5OXRJz3PtGBn8omXo+6LdtqZxQFDaJg+5+yHZf327xc5ilUhMWqITol3sgLl2nJ1vOae3qfLUY+G
uT17S3GEzCyEon6mdGfU5H0KowXwf+N9kAbWWCS32XbEoI1cGWxSEAJbC1/SKgT19kIwktwoAIQc
up6yxVqc+w4BYTCqnFMt2xgxBore3x6NP5QqINFfcCzs5sNBWID41VMSPPbQXnzul2rGuPwbmMbZ
snwAa0rPXmY9fW2bn8L39dWNic3IzFENIEmG4AkQLVFvMpiozbt17M8+PlsMA5ayBXTTw1v/qKGo
+QTU4j1TzTXzYHW94YWL2XpMFMXyWnb0Mzvf2PNnI/Zz+B9gs4uiYgFf6vdVaiEehffgBrJmiESA
ya9BRFLLWTW3IiBkAgseMZA8gQ9srSgUe1yDeUA3vk9r3cRcKecRmNyaHobCjTjpTyzA3MQNJr9i
TVdgp2Galm5H6SrRQ3J8uZ3LVsfzskbFPV9qpOuQnXYV7XpXDrb3BR9v7PkFzp2blcfg/kqaQTEl
pMdrjVOmxn9GUy/gqBqzB6x5Z+4bCix3XrY5TJQaGvY+KIq43+RaKjmzA2QJbjWMMyWASTX1GRP7
ziO/uRwlifrvr9S0ahn2pqXiLQfUAF59Nj7vR1THnXCN2n1YCvra2Uzv6EQJOUn639D2IZfO6opa
5L/5zsJYaR7gFU3t4+iFfv4Zn7GrY3gISd4rLcACEdKM9EfZFwvU8VkatMiSpcCZhQjsUkCZ2sp1
FKYATxBx3pbIwpyeIhRlB56zIdTUv7KFO9WCVg7vRmfmwbPJFHSx5Z0ivmfFmIfyf9HBi6bi0CaM
uauU8McHMpHlwIOkLLoqDRYfjR6j5o9ZggCLl7sxEZ83/IJ9H7guv4U+59EBcE1lZ0x60MFgRc2Q
6viv8nWJz7M1o+0mSl8Zelkuc1naSEcjDedfp32I4LW56R0Ix5601X3WaaocrHHq4/JGXBWgX6L/
EIFJbv0s1e/Z4jtc+k4/1GySCDgkSfG2R+70lQjiXgUd1x9/klI+NQ6KbHMkgZmLA8Q5oToe+h5L
Bi/gWsfxSUKveVQMA57TzFUQ+YOmYqfjwElNbVkwFKYSLwQtcs7pp+M+73+FM2jOZ0UR191Ykjqs
ia5TLDMX+qAfdATAvLGX0EYNzj9ZVzUATBZDNxaGjSOVhHqZ1MTZ+V/Cg9vOy/eNuT06Ek5osLCh
K2Agpn6GIcMU0hSCI01lfFLVTO/C65V1p2G0ce+a4Bf79Y+KjSPhYH3SiqNDuKrSpxXb+JBXODtZ
YLBJAoCuKHxw9C3JAZjak/+4p33Tov5MTeo7/mtteTmHVS5NrpAqSKS12A5Bbli8NWHvsN3r9lC9
xXDah6uFBQM6uMXuZ4qSTBmDF+Tw2WIAPHhc/CYj5tFq7QotZH8HoR0V+xL2/gqjCtZL3Hcy+GdW
1wVzF5oenZmaLVgZpCl4rQXfLZinH12NnikkyQDAtSWKB6hVgDUsVP3mrl3DHXMqzKG3X7XgDuyy
1JjoSFQ4vSGIlwuwglrWD5A5/uRsgRvEyBfPrAv5bZ8i5dnD60Vnv9b5LBCWxE6AiWalzYbBQQfZ
EwQeKmooEbK/iJw00JYoflveMrRkA8oOcDIA5QthbsR8EbV1nnaaTQr47cuEoR5TfLnPlHRxoHyD
DMNPzU83zadF1bXLJnKl+ZWRzddql5NYKf2ImsQuFBlOQjoLrSEydNK/sxOaVjWIBLaPkcx5oq+8
UlD4d3Z9r7Gd4ebFrbAyyw4EaTO1wSYV80fDS6ZhBgYPgh+nvCyqH2XZ/M1A/7RsWRfXyawwHnWm
QmwZoBnSvrxvRRr0xU9YcX6Fd941rIZyFC/LHboRs9DZQFZ6W41ry63mnTJu2mAEpDYRJWIGOeG+
MmyUBg6ir6Iop8czx30C1/yuu7cJw/VMLrrPnysSppGrqAuWwx6p/0FXHAdJl8W7vVlyaYrb3DCf
WH99xDwTNcufzWXSqYoDnqFRMsBad6H8h4gFteIoaxEQKWG5hwKp3EdA0wZk9Ff1lXz3d/6m2oq+
bCyY5nyVjda5nlx8npZEj+O3GI1piU8P66nK1FdgnoD7mSF5PcL4N7gKqiHAAx2vdNKYEmP4GYa6
prhtioj6h9hdYPlvVGZ9mkCU4POrishdZ/7EuOYIrfTXVsUjILV7vUE9itguxeE4jOWNfZagXGwb
VRtn4Cye9bND9PVxRCcSDE8HlI99gVdPvK7jFAs8zx1hHd+bbebOtLLva6f/xD5AkmqU7Wch23wK
vB5ydJcIGkt0znuBi8+w/dO7LsY9MMq3BOtNeYFN3cIEFX2X75sGpjZl48FzOpeqnH/xNcU1cGNc
Po55bP+M95EqN3/yiTcDlsfiC4IBygJF9FgXI8J9YBZUBwqJL/g1r3NuUPxrgUNeSrzQwr8OyaAC
NYI56qM5O0vx2qhwfA1sFOTJ4tZDGBaDm2XzYamKbVuEyxYLCWINaQWZrT54HoQjjmwEFAMsrjop
d0oR0WJVTsW1tOI/zUmtWEHzLxQgpVpiSZ/if5UlItr5QiuKVqhs9pH+h+DN2XDZLlb5PqOH+p5t
WOnqzkaXVVmixaw1sY42HHBm/Np07rLqOXqn9VzVsQGAkXxDh/R/8mTSecb7ygl1BYHcK5sIq5R2
AfE2LDbpUQEX8gZFEBng163Zx8qSVtwYFjZWUSwb++TRjIrfXJvze0VligNOYbmfvRY9jlFN72M1
54LD7BSyAyu1YWJoCfkSnzOfo4ja0ngCJUtj4cj7/tjxV9wZSYIHZU8YKGkzhwqw196pM49CqBAN
teU2tbyJ7Ne2Mm2JqBYFj+Z6R6zfL43HJd7mc1OAaC0Nt7Uh8ePxzqfv31TCedqIuQBNbJKVlIQV
t4UhafzVKq2tyyfwNn6k2ba2rhUUk2OP0KTPlMwRIKRuBJWtkSA+kmDX5UuAcFybaIfXTBQ6lJg9
L6YoIyyEC0Q13EslSdkdpqLZze5pY/C5UqI0PU6zIIf20TbhyK6rG1pYKVS38aTg7q7sxrS3KYkN
+ItpqGkGXmfsVt7VnyoINyx6k+2o4PjhZPQiQBILVip7CEE4rdssZz4Ub0PPvTFxpbFMAx45SHXI
DhWzvbpn3JYJhzabR4X9NGPWurGot5AM1Qx/dvTLE7PunTWMfqxISb9BdDQkWyyKna5TIgBq/JG+
CfHXqL00qLV1aCqNw1LlZd2e4gQ8hYR4qf7fIuNUT5qOWPQv7H+zThr2VYi7rKrdt3dLZYZmPl0H
IggqMh9EsMISikSjeX81OK2oSddCd4ufAxmc79DBIr7Ww8FXkwU5sKnbjfKHtjNfUP0fRvkfgAFY
J4TN/jTz1slzim8gQE2MKoGCu8x60LL49dRUp3ocAF3wEXMtq2aq8prV8rqnRbj3Z6Mt4z+37+rJ
KEyUuQTvpFZGCbIlmYvPUvZGF2xBVL+Xzb+CRPVeBnldx56pQWiwUlqZjVUEGZxCrp6uYLFdekqj
i6nBTJsetcHOdZy+OcnmHjb3jugJVNBdsYy/iK7v3aWS6TCPze/hPNKT+999exvU5yPgKtTQbHRN
koiWCthfdDU9HnDPqVMzqZ7oRYfGuJXgKvlFIKPKbBFCXCFSisZVmXzrAkTgZFtEu1SJV/rmdwU6
gENBR3F2dgPIyvU5yp0jeB/x1lNVdHTalqJG6CcTMEU7aVw3CCZY7m/K+FYGxRV3eutf+gdm31Pj
RNXZwzIrP+Tu/3hJL8YVKCt6CJIQRYK3zIbUbQvvraTCWkBB/EnCRG694fRpQSN8Z50skRcRvUYm
PQ/JIyMtgpH5BdN/Ws0pO3RMA/p+qgpZqvWUQRE2TpAMAQP6IcERUoLjL3ecCKDh0vEPY7zkpsI8
miFamkeHkayNE1XWFXtKD8Y9kH8WRE7GSddGIUnTyLuLWd7udClxFfmyY6cy9qtcXyO6HI1PCFqh
fKkq85JJOgcqkhoI71Bujq+JjzqFbhihE/6gXZwvtZDqXFzOyciGuQ/7lXPVSK4N4tYfXZnP/vor
2FWOy6RXA7KXuIKhUQa/D9dMrFmwspBYZKBxlZCzuKsf8INuYRY5b6a2SffmMG3HWEale39QFD5x
p0KrolvA0bbv0lXgqk1YyZphEFEKroHnUXsHpFK1wLNRqyaCqhWkQ0vpHIoInbvVAIxfSYhF8eG+
5dXlMgl4uQBx7c8hYaTXK28DrmZYK5OmADhWQUKXs2Z+T3TAa1CJkF8Q274Ax+XLUDovYy6YIy1j
rJ0c4eiR0o3778FkTbE51WZcFU7QZNq7xXzaZwngIrF7yxP7UD7IbOlZSlDTh/R6FwGOM7mFcbIU
E5nr0MUmkxSJFttd51aYzKmmZfcyQONW/5QMdabyOeFgcE8r3yAyttDsvt4IbUcdS34CdDFG+EGs
UQGq5cQ9B9QYsk0h7yblzgB5+Bjbi+eNZzZnFUU4sDa+0i0gnqCA4JyN1+ea2ukjhT8EU5bgXCbC
B08ULV8/yzsHpnO+9q4AEz5nVo18Zs0xE1yVn9XLQ4lhTg8CWNfii+7ZtP4UeKJcOFdUgltK2BbG
rXbf7CnY/LeMlFXIyfw2XmCrd+5oJz4DgzH/AA0nnABmk8iS+I02bIxYhBFPDtxBgLqyu4wA/zrB
gF7/VxYfqihrmkcJ5d09MBfK4F0kbCMh9cET8gkkbkKc2gJMwOLkTlwBIjyMv4Q9+cnuZ7WXPix3
/P7WTqV1m74EYpie4uix1YsZPjVoYxdY4ES0C++1uvXwknAe8/QCUeWelVYsk7fmIAbz3kB+Ae1z
P2oxxDD9GOD/I3/6UG5cQUGGv7Za1o7Eqxxk7m1qxcbY72MkcZzyz6+gsxjw9DOSdRPg8eTjv627
2jM2ctqc1kBylPTUtDh7hNylLb6aqbeDaIxvzW+JjJoHgP65kBYs6uVtXsFezIfIQhbSSz/rmUK7
QM9OSwT4wryRAX9aRSLrnqsXc/VOVJ3A9fr4Ljeli45Kh3h96/r8WBPemN+HzDxgLUk2+ljprH2p
FKK/gRLkkGmH0tJaqDHNGJ5R20vkgAxIbNWhfLDoTTiU8W6zvjcbzefUpppVpllAITSxXijDlAHe
fFBjJlwGmxasXhdnYls78/HNYreEyLOyJX5xincJQ65JHh2mEszpDERfej7+/6j1+xK/MiKAl8KW
HEZIYfrur48bGJdEOofNKZlR3f3M1kmzePbmg9khzmaQ76z4TKUj1TjPpyrfO/IQGyRBxGXA8Aba
OqtbXRZRwX9F7a4lEeMENx8suELXbtMMgr1v3USG0p/8pldogmFf5nlPPvC5V9Y88W/GxqnUuvJK
I11KHMPeNKEYyYLr2p4ih7aKVHgZ6jq/c/4+wqEYRWS6SsMhop+aNNuV0kjD8WtYan3HbB+JXRiE
2M3cJ7mr3913T3NfrjglgY1QIIXiYFp+NHKNSRJW5GA9IORa/Iq2hSi8cnnQfjn8Rtyspq30CAk8
y5WLLBKCgtsisnQNVejiW7+AfKN6Urce4pK2nh03CrWK2+iO+EY5XqkCiTsRy7w1HHn+N/dXKBfh
mlTbw40dIMWRjdXsdqytLCjyVB6qQw8ilfx2DDaG+Ica7NeVmXYAR16p9FxcPQnSlDiAxeUXaHwS
DpjIYUI3ruZC3pLiwU/VL6tlNNWLErX/Oz3CJYOu7CpiaIJEj2eQYCP2R6H6HZWjSy2p6wAIPcnu
Oh8MNnx5Q+oDH22dAsFBcHO0I1vwAeQ+/fm1yurDGz4IFebg/Kd+0jmk/TbXymeiNrQYinTdwxCa
CFtrKpQk/qlFMFq7RkVCSByfqY3ysVXmU52MO9A3ELgIE0eScDDfSCu8lA29DneLInW8hTIxfFKh
PWsKSBQg0LncZaoy33J3gnz6I4mxv27jm/mN9koNvnupaZUaOZ9nNEs01k+9WGszRPTYz9VADGRm
0iwJlGCQavsD11s1f2JyRiEtHgQNywbzk9eu9lD1qcBI37V9ny+iZ8SxhKqKEw0sExhJjdikTI2Q
jAt5XCIWcNtlUvySmigMz5JqawVvnRxT9m4W0M5UvFk0RPK9dw6E1ee5ACN86OrY0UN7lqrPfDvj
risSFjcEgLPiCQUCRfLILdQWm/ZXUoNNw6aHnYvwgcGnDPahQiYHiRyJlfJX6/J2F4ilozQHKGDE
8AnqrKBzsjEfR99gIRmeHgnPqiaxbb2UN/o4YDRAlrkRjJjZRsoVGJjF3Q204eeS6avHLQTF3SJa
nEvRnqI7NGSGnz/nJsNIT/cO/bDIpv1nawHhB9PUa29Pju+g8aNvNiaRrxVOlrt+g4KAArtGWp6y
oEaQES4JgQyNSdHsqbkwlubRW8uAQWp6msk/USxzScSU5iS9gMWW9J+ifdCObXTnoTDIcWYkJPVa
QG1wFqu80JmaBB6Dhyxqo4xBGyx1Eu2Ygew6II8Vo3TMAirkGmnUbLGT4ONP18vlLxaQnRmx9c0q
S5wfAsjGx7XXj4KgDRy2lL5jvgxaljE9ZTRZSF2ryAzkq0ZVT3zyIbCagWbrISO11hG1eyPh8+Rp
1MagwSufw2OMopo68jaSsRxOrJeJyHSBVYhRedBcXYBDrYMFrLqtZnpYQjPFyE9+AlfPQLQle8Yl
mqAgV4t/5q9gbzwHCN4ITCJ1oqmUCzqSC1wE6/xRguupafmUUBVkmqOGAvu1P+l4MFkT8B+ahPKa
uuUYpFcJuwy+tzjY9T9cOxjH7HpijFzFAub1U49v1iltPs/CwpCgd9KAHECoos+fCxy4yco0jaLR
qlOL5EBkkHirdSsEvcFeFmpsXVyNKCd+8lGmIrpobBGVGtcPU3wVU+3rGj545ON5uo0zzGfi7vzD
YrSE/knOl1jmlljD/dmkFwUYd3Jb7rO0xr4n35JfjOBQq0ZSBroLq65gkHb2+M6v/OwU9J7M/xPQ
bHv14GxmQBN+1hjapuxx8req7oSh/gZgS9VaKnDLo9vG8a2e1lfko1sK0EwBtgfz0ORaUNBnLPm7
ODMtOualk6FNn/O3+eNmwVmdP7f41j1OBtAf9+wsZKvnjUZE2awYoPi+qFCDgPDzlSY05VJv2M6z
VtHi9BQnBHMwKe6KhCLiSiVl18rQnjokiDIVztfkP7tJk07KlsUcZAiSPKJ+lnylO1d30Ji3iU/k
Pn6T5XRPHyacSLFXFev/+UUXEfZDx0vs3lGKRfyp34DPic+2Lo6+YtfawWHhY3iDxbWjZ6txtfbz
x9Af+eHfgTxER7grvWqxbin0eGmabRIcorJAHtkeWWvMJS5JNwdrco6soQrcaHfkXyhqcR/hjZTr
hYa1DAjaxgZjNSLUcr8VuzAxW+aaKmBpSIiK366dPkexV/3gGLrgQzh6H1JWSrZq6gzCviLdbXR2
XAGEYqnlhsMQKbHqWntx3MQs/Fc3sPBUctj8xiqyCXDG6PThgXbzkvv3hPzHD2hVsff1TwbtNTMY
Zc4lW2ouVXyRb4223xJR363ea1Q/6hMgW+FPOw36ci5MAhfVzXdwHW64P6go91JWVXrNyeK0XieP
/fdxIJOrhDfJKRVekG5R5qRiKbbMHzeMsRwUnAIm1Sgg91eY6L51Xt6c6KqNMGk6YVHLda1SLvCL
y09dYNbZSgm2D/kt9evxyTkHziYyoBe+/qFcuCzx3WVD4go+FSwEOBxSKH57uubuT0Y8j/hUSYgX
IWF6C+cBK2MBF78c2RoagvRhlkAy5y73gyZ7zqxAfUVXQWbJ1kpBjE1DmQwKfCNMpcOh6NVYmWR2
SlqYbhZW3OWdfO9hj8d/yL51aPJosuIkiO3rNDGwyPwOrDb6eKWQNgmrKrIp7Chpa32k4NiS7jx/
E0LDGwUDUjZKSw9NDbdCL8q2NNqy0bsTVlSxZgAjyLD9aypsXHCfrwgYCWqfZ9iHVsSA8dZ13xor
xUXGprqGOSta2xBon3cDHf7ERDHBv0e8FuZO3SLXh0atXNKn4Kpcn9VUL0A9ulQ0lh+BNApXFbo2
2+Itg5178ioCfyAm+Mh1CDLB/W98O5OBVqMl4EjiGCRNeGTRLNI50TvxQCNeUPBZLquktEYdrGko
SfXiryJePGvVSqWS3ooqWss7yZ3qhWysCFfWjAm7ZiuUujM0FUd2HFGNwGU43D9yykU19+J2spdb
CFww8NSyNgFwOoMNDKaYfJzp/4EXvyqlEU4xQtmftKNuOFbZoLByE0Q3QLaWzELRmqdtX+GZN4PV
8x/D7hQxt6ATAFKjZzo657EbQOpbqove/GFweDIF4QXmZGYfkl9NolWLSpUqHoXpvJzeWb2cs+2d
FRlhpkQCcLNeOqLQbQ6HmY/EzWqR/eZ4W+1eKh8ICSd+Uhwakv4pRoiGz8wn1vyVD98MKqBbNBa2
l1RLPYWWJDROUBpVKw3vxhSg7hE647ZyU1yFKTwq9E9PMNMVHwMfghGOVhyX0KdrEGnjI43K8s5j
kapAkWknGmgvZUeD0BT1dVM/WlVZIKAFJkNciRrbdaAZ89Qrw641X6pxodnjs5WEQsVmvZgWB136
n4kAwD8BfmthF8BKpcOsXpV4a2BmcKjin9MYJmEuoBc990vqLMiKCubcQ3qHeveXV20Ftk3TwkV4
VofzFN+9wuuBmiTJQ0ATcr/4lDjwmgJ/vhbBnDWMVKsBvH1xIoi2aKXVf+UtelVTGLBgmTPRqW2B
jNTp3NjLlCKLzEYU88IlxnC9Va6EG0AMjPh6T5jVJypr+Hh1KuvKk6kYAGbs7V7olDkrB0iOrEQk
36T1wzmuzVuhKeFQeb2D2TYWB06azQl19/yeMJbxycbC3hES+P3WjMC2skY6LjFq6keg3826fp4N
vCOdk7rho+XzrmzPJpV0WHwbuMcCvbxKSYtE5hUgBrRiJ/GIy2Mty1jG8d+G8JsvB3hBje8pFLk0
jXiZaqXhDRq6jXaiKsyqVMl2QNKxKua5BohX9SHI4edd3i6pnRHgo0AoHsiUOLlLRmgwDzVv05Fh
t5mi5j/aCjwgOaCUNuAvujUFU2NA9orjOunv7Owjj3rLh2uIPTjn4zHntviUCBQK6rzFgDaV57KH
wcGkZyJfLf6eiwzBOdXnat2Q8ROVv18HXUvgvzlhQD58Fc6eneVO/e9AtAp6kmTZqJN4sHXhbTx9
ehzQbvcL1CJe7WLbH1ayFgqvptLikJhdwzzFE61iWPMUy+LzfkrP65KnSN4a5qt7GuS+orO/G0vz
/e/SHIBbjo71BBe6qN9UrthVnIrrl3WQDSeelM4kfWfNo2upORPcgA6kDsN46pCcS2MwzsFnRDJ5
DQExu0IRy0WJQlQoUF2+egz68nqnUu7gqgTYDu0n+rGL3jnSzwDvXazbAMDSd69WoyQqAwv4eOPD
ESKfohRjucwNFJqZIoPVOiqSw30SHTNiEsWlRDbZE64Fwx5MQ08VmBZ034T9DoD8yz5dwiaScMrU
lapWo86i10Uiiwwlo7KfOfxjyftgwduz9OXQjy0flgx5tB5mY7NowkcfaUPMvJSqtHQEZJ8FoFcP
sTMHTGwAku8D9KY6NL+rVQxHpfscWaCWbCZ9o07D2qjaBqbX5Jaqnu2L91egxQl9CxSlfUSaYwLw
xKFMlp25aTP82N3oQpWFnSNOZPBWhvzm876j6NwP7GJvzDvCB7d9Fa2WTw5jcunUpcW13KFtNcCO
PrCawkAoOCH3WRsDlmfrLMeSfLJ3mUNalUMC26zjD/tevEqHi7zn9eKHelOkLPASNePwiAkNXuWR
mNcp9d2pGz0ZvmkVgSbarzMUEtZGppezstSDI7xY3hq9fD34u/tVf5+oLdBCw52bZWCrVyUequpV
eN519e45S6dOaP5IHoUKQXiYde3Xv7zn+nMFpaCP+J72IK897q5W/JIe4MYL1+MIos7oMvr6PPO9
jADUj4i4tj7RrBpcL0dR+TMINNScwcKyagUQ0WURAiu8q0AWqWMXawnRb811Hab8gM73wG47xv9Q
5+6anzuJG74sKsvcCzVPftXRZbBa8USyIFB7XOZzk920cq7wHG6G/RJsKQMlgdObh4O4IWRSJckI
XoKLqeXXB8SdxFplLWDci5EyGPmbYlqWjF/wT5qlRcZN47ZdOBBFFdP5QlMDEzJdzcm9Phm2uEGH
fO/tzyBZ3CFwhwEsH+qGpHn76c4bQJUhQjOoop6ujtYQDJS37Y/10xib6UD2IxMU9H8k9uCJA8bb
C0eYYWIJbZo9rDKfXFsLlL3IxSdjBMPYI/21/+/hDy6k314x14CH9ViMRwVU2zyHmlVuaF1VM5Ow
MzL0x+Ve6u/W4Cv2guw7Vm4u4LMyKRFY+KdbwWPmc0lkrH5CBIQLtGdOM1g/DPbmwuoTGXihfaHL
qV1v7ISUdqAfgFFxEwt3IcZ3GKgSKfVi2lcS3RYIv02WL7/xIBx/NC78jRdN1EJVnw3ZoDvMOBf5
+jalybaQGTwnidp5TVpGUgC/nHtjQX4WZlA/LTI8X2GisITMuHbBIU18/90l/mk4AsZ2AdnlpjwB
cJV5QW4DIk6cWntFIwLTS/iy6g4Egx1Ee2xk/4RsKn5hXKt50xvKnP4IYBwk3mnmOuOkwMxm5WN/
j3vXJqsMxUy1HKcIWmWhhhX1euBIve4KGQinVcySxcfW0/VjvShHkb5qrazIKT/bBoePLEUiYrEd
+iJCZ/AxysmSCz9R8awQU9UT+uupCOmdAJxUnosQYjU80DKJBwPlS88hklrn6IE8vUrNF6frrGKt
laJ8gPab5UsTIWlFlRi/X9IZrJqR2MvCdrlyiGgaJTMVxotbosaSj04Z8kTxSogAUrhZvQHy/MpB
rwyakTd+f1AOJFtECsLi3An4RiB0k4zkoVwlCyvrmUeiGQ6uq9TtnjDMSY1dOCYAl5pCgszCCaIQ
tAZXO+FWnBlIMYikEpFtqR2eAG42aCBZ8iuNNaVs23O4uaJPi5A+fq2h5NgjrUV2RcE6fY+Vw1cm
HcBMXVDdeVvB1IPcR1x0XVC9uu8yk+n4DqCOX6dqAMGCESzCvTIOB1wIlNYy1z4IvS/sDbe3aJbC
Re0f1bBXYClu3zQFG77CZItkvO7GDIq9e+3BVVVwOtEAf/TTRlXs1Gi5ofPXE3Hc97s3d1cjWLiL
pxm9cEW68vq/MeO8aWdbxXa4FAGIMfCepv/XjsNoin4HumVJYQ4/Biu0uNHEj8mBcHcO037hPrC/
K8icRS58Auo+k6LVA4GFDSwj6421PdsVABo4BVKXPs4Grb4fS+4fbohYQ+7UYRzVO19QEi71DXqv
4lDS+OqhND3GykLhIyL4yWAlNDBLqB9E4xOsTOTww7ENENYlinXxl8hAcUv5YlHqnSFFY8VI0pGj
2kIxRrwWubi5uoNpAR/BTyLkvo96NatsgxUsw/X0hzeD7WxNAbgOJsziSWpQ4UCh1Cd07nla2q0w
s2QcvxcMTRs74kyB9MkWGRbVWQeL0DhOGbdlOyTb99FUcu7MzkcDb0BmVh+C3LqDVsaazaBpajKb
XUWHI6UXOsATA4egOetHhpAynQELdzBE6m4qSVgKLQJNfglTv8NvNOYycCIvG7sxFS2oHor8PB9Q
EFi6dTksZRBFhK6eMWraY01QjZTXb+EEItAKmzaH8hmrbC1Mh6SYoh4fYf2KhAARAzWcEf6Z6BkU
UjOMQ0Z0LjbrAY0jZN2jhFUKu5ynEYhcEC3VdVmJsMzXQumsXDnRun0YUHF355+pFIU8UBGCbupU
HbxqnpmICZinKKhHDPH+KTw0ufC/B1kfIJRPRRJ6qreiuxCXPsfov7WR6U/Awez8XwB8rjRoMutW
BekMthR0tY9yqVttaSZ8GGHVgJv+wQyHOBh3NDsAQjZPbAzBKPIN0S8c3PGckSB78xF20upnoqqn
TRAlin5IACc5QpsktZ6jElUQRTH2lugxIsGOqbU5NmVCbW0OO9MYDPeI8blU4xKcciBmiu2rFBDn
TmenYkL+PZyJq9OMLEdgwKqMzpBXtoRSdikxy6HwkU/xFyhzPKqh3kz9dsqVtNXGrmSKeoKV1a23
U9pgwyI0qmiIm0meb6cZFEbLmgVdOkglqSZ/W0tGK6p+mN4Rhct+TUAjdzIrzgfuRGOM1GMnj4zf
t8n1z+pwh52gz4I+0qBPhSnOv97vqzOswxiW0hiyGHkihKiRL0MQomxL3TnYb2SIxr4TPstxE1WS
29ULwGqNG8uGrjpHWaT5vw7oTLpt2QDZA/JAoemkRQheUL/4ETbez/SMLAfmg3Uu09GRwkBmRhIT
rxgTWDhYvvVJgHZTyTqRIG4kSKj5PuNz9uiWoMdFHG6j2zx8YUpQHo6pgM4xDbfjF0nb+rqzuA30
NHXf/BPAx/KFGWW7kJiK8LgpR0ip1CpIhpVtv+JutmUhcoJy+PXsVZbyKvrNvnHM+QHk5WyPJ05W
nSfCnYtYetU4sybqsiRsXL8/xcs2UT5nsJOoC/Njs/NhUu8fBh/UmsE820hK67BAUDCIAeohT1wP
2ffW3ay71KeOuhBlZlEJbu93iYA+BQyWQSPk19Dk5exd5NE547gJaf7wIy0pZGfO4ilyg9tlQRbr
EoWSe1nSkgGLohh/TD+r+vazD6uv/h2WVClLQj8IQzBeBVeEgR928tkL5CAXF+qX5F1i7R2sVnuO
LkJjq0jS+Zbs4SWypupVjePo7k6PEQRBxDPse9XQbUi0UDNvsWOI+xkRlMc6klOD5ZhW7tJl0TFO
2G/PjgFwOqImo/fX2vtZLt9TSkc31xpsCp94uV+EZoza5BHXhkvItzxwh9JwpYEatltgqNfox9UZ
lFiA+0KMug4hM9Xx19zu/zSkqpT9ERwrJeRDYdWRh04Meke0Ifjnr5fs1UUy+uykp9L7pV/y6GyX
MPKkPZvEX99jhb/WDhV3/OAMugfO5dmOnFPYyFF5+zgOz11/vlnPt7v4gjxs+2MlrIIwkSbW1+6Z
Zxbj8Kmv/iybAAlTcpB7CCc0fNd2rtBa//PYSF+G2ue18y2RYo1gu5tx5LpmqUFfIfJJov6Mmohq
JQ1Z2amaW9NLOjJa0oXULMdvpsD80XZknw2n+ARoIqSeLnHMELq6IuyLSxbX5qA3jE9ovH8zpN+x
6jmXt49WSPdEZu6fBk6vN8MfKkPLwhwToaMq/e0qV+Ggt0KAggbLLJ7BtbJBp+5p676Gfckw8C3/
cBspcqP/0TeNsgY4sU7Nm/dlv3ASHaDJpX+I94Yi5kWqcfAyZfLnLNlrD2/GDDyDK4fyXAipLpG4
VJdB2NJjDv5gN9RnozLutVOGVcA3DuSM8VCkFIEcBPWqI6ywd2fsiix0NYcQ50KaH4ufXkyUZF5h
Gy+JZrTTjTR8zoL8vsFrjhkxYY+geX0C5WxBOcrqRQEr8IrCkm5IYA4GlBhNmTW7b2U1x2EgGi8S
cxyPONaFK/WdzftVpo5hou4eaYUQ8/c6yAiWr/qIIu70S4fyKk2qqkUSJ3zUsM0q8SCi8kCBlsRK
PqOpufZMmEIx8MGiAPuqfbsmA/LNQkPxBrYyrjGXlbBIUtLP3RyhCAjAQXM0aO+xZZearsltKSVK
F2gLyQeBpv86KSZNVd86uK9KMINh/rN7KpkRPIXEBef7N87hCIdNOT1nkJdpGhDSf4Qy88y6ahXJ
m0DsWW9rDwakByBlXlzPyI4/HvLCE47FhlzbELhIdFiVaIKYq7xtbM+Llc2OEMOTJtiTgufvQ2Fa
lRc33cPXmXw9Njl39NAVLaSBMAwTCJQHDvCOMoecuJA9qYSbJkDGywAcVzkJoaiUIhz+wyZO36XR
5jBvTXWCVZ4wgZEblqGEt4S6MOmrwGSg/SSOdsocPq4hi+0krsKYLGr9UP4TKSl9Y0NlcsBQFfqU
GHGBRjQyHLYpxzTQfy8d3MSHBcCcBwHo4RffiN5a0EMr+OgVN4HebkrKMj6XFcSotSCHzYrVwezC
6jFNsbuei9wS6a67SDyVjJNzsh7DPPY5aMzL9gvA5b7bMJfTsZFYPmR4bB+d9bVskpnh6EXlXSwI
KXWvhHQhja7Dw6nWEhBXWOMRs2dKbCj4MDMYDQxahgohAhzH197MWQ1/uPAo8PWs9D4WiW0VKiUE
aTsq+C14cTv8uEqwOpOUxmoZC4W8f9LQ9FgHBP2cKg4cF1OCQELzbqHX8SbR5D/K0mhoQr0MC1rd
7B3gcQktOOHf8miEKljcy5TtHrL6PkPEpJeLe8HARXffRGzR6G5eYR2d5t7+2uSWKLxRLW03fXp5
iTf8Ll2TsUw263m9YY5B4Ef7/k8HGRKJkKS6B5l7udkx1zbGc5wPX71CtBc34SdzuJxCWz73BvX7
ZYcOHiQwqnbXeVO6sYaRsOJRu95YPrCjjtdYxvYF8Ech6RoM7WW1pmovFtuWlhGR9nfzZ5Cbpnnb
pYDV68ThTvhlm2I1p0MpuiosK/8xcR0MpCU6DaAVZUqPvTfVmxln5uIimeQ9I/V3W/4GQsm3izWV
X6zCKN3b8/EQxP7Z9Uuu3KyIZt7EjG56uWZUpv44/R3PFKCeGZ+keKZ83hxy4ZXWmAhMwMWsgXMj
YSlTmPanBxyVsYE/VHexVvZcFd111OBJg3AW/HHBWhcUQ6I0aZCMx6JqFVjgexulH83j9fJNM2sb
dOf10y/MAIZQ4t5EMbuy/k7RY4KwylD35T1z+mLHPZWKXssjPFHUN7gYAogvhEOV5xsELlXlO9+N
yYzNajCVPMmdC8hA/nXF0XAzUhvqL66tARX4tVU9SG+/k0E6QtRbU0CKweZNte/ZA5kYuzczRzyp
6iCjpZTHVqGWBM+9kZ6VOtKz8L58ZOD03TxA5ABTFp5MHajxCjCD4ulP99WtNvf95f3P+mmzjC3+
LO5lgHpKPQo9xx8oSshMNiA4NVaZItLP3XkZ+av0d/rZ6RcXYlZNEzv2fKZ0TbJznLi3foVDV32c
upxGNQlwgMRg3gxylykYEgRgmW2jJMOZMavXQYinfAoFcrSKPXkHWOYNQWXRV3VUIy6wp/Tckwie
4SHO/RG7uxZ+eZEDAq5itxunaLZTDIcxbDu66UCY5Ji8hycj0+pTQj4G7J6694d1kjD0gfHOHKdR
1EIlW/yWtY5nJkPvKJt+5U1uz8XafMyywoOXFZXq08s44XKoQi0+GeKgv4Qo+xBOhjSwyY+OmX/j
sQx/z+iJ43RIqTAUzLMSFhRfGjVi8cd32uVMnxAxNpxRTA7sz8uyqykuiA1w+peAGhpyH040TWMQ
x0movv9+gbkmzKrtGFN5NlsWaQTeuCp0518O+i7Eiz8rLKWy63sWbK4YPlk2wF1sSV0aaEPNZY3W
euG4+tYLs3wOHt1Y98YnV5fOHi76cZ7wbF++z7j1kyaOwrey39lM79lA3BFtZ/9zbLlpG5PHmbY1
ESv0bFIrcjAEEsshiZM2sx98gV+Um/wzKDcQcvcsKYl5NxvqZ2PnqXYoS8P5AiTSsR6RR0djZqRL
v4OrnkxZlyGnflUzV7wxtK0c9OIN3b7LLOsP+3D5updjEasxe+nKLzGnicfETjj9u7cHKQoDrdJ5
gfNwqyFvU/JAYm9XvyHY4Hd5Lq/7Y6vaOx480d+ZKdMYip0QBBNjqnkhNaSRqW6zixkEtXdZlVhq
5tCULxtxeBr9X40b8kX/onjQUxf9avuVj3oxz3XcD07m+lLQUALXoZLt/00KW04848aLfRaM8Fdr
8YnFMrSnqv9AEBaOF7wQc0zC4fDcScx1TiGeOJUvULpLxhzYKeqmkX7ckIUBJyox9ZqNxq+jT2LS
BIALJzo3m+UVfa3Jh/EFcrKrcGbGny+1ZHBbP6axQVEpvAuq+LCrkaRKAS14S6vB13UqLwSnB+sl
eaVrvmpn5w5ZCuyXmADOZbeoR7Y2NXx8uTq7wVxQRpUVhJJ/5qTKLyF+pPPAatzZYkCHKuWoJydT
nOcw75t2aSG5pGIKxG2QqT8zWN+n0uq2J5uPZht35BZDR50x2dPI8Ogvvf4/Np9KEbq0O45AWU1+
J6vasKTC9KJPo9rHSSEAtkVKuko4FZaQt60A/BidiPfaNRVoJkGrIUIJZhwtiRyxHNNt13Lqx0Hc
PaqSvk7tbUih+1P82B8vibnjcfZbeu7DDHjeCGP2gGgavBcIPS8VShmTIZy/M/nOeArDoyJugyRl
TFzs7DGmGT/DGGO9sfxDIJe+IxnyZkXKZgcW0+xhP+TR9XSMMOddsp5U1DRfdOeejyacfiykbEpT
ENMu/Cl3Ff78jmab184VqhTLf3e8iyry/bfk8TMoJNnfA7UNLQOio3aMOOaaEhHxR9BUJk6ybtmr
yicU9aErl+EVYY2nHD+1vqociyLcPK+BH1iWazfOLHs+1yGVP6ExKgdiKmS5XwezSVdK2F1cSA7B
V3uQ3kF0rZyK+UHtx5LSDG3RtPd412Wd7F1zycFSgUjRK/zxqJO4POyTy3IKlRfzd/HAW6mr3Znw
mEy64TCHrsCNy/2Sdq+eCUxWyGK7nLYWBAJ/wp02k4Edo9Ba5jLA/VMv6oa/MbH5AsnPUEaW4yfn
dYaMxkqzY3UdARIN0xtl5Nlar4ne37y788AWExN0hpEvcLMOdl4A6/Ys8rRBNKlHW+oCDoWwGweJ
cYI0IreAp28EgecrwvZRmHg+I4b9/7JafpY975sqfDhvipvC29nIl/U8T+8xtoK9dStu2RgKbxkL
Cex8t703jzoYcaj3IarbbxTTolfQwl5ygLBEE7KjUOiakYWtWvLfhg+Y3YQsAnnASoWUxMIC7muy
jsHxdeNMEOig6pHTwieOi3ljTJID7ZZaE2OAhZgYtVas8Wa9VNiMY19EOsgTHimNaiNbhh/noQYE
FsE6w5+Az78FDo638VU72IvlURgopT2lvGRO5FarWkDUCC26+kPzTmOQqfYd/xBKisMfJ0t4/eYe
CydbIgvN1tlspHgUjvIlz2se5v4rKGL6sJQmizmV9TcU7R4f6cdfCvQ+rf6RDSgRm9Looqftt/sX
Ys0Sj8b5DIDAKVox6Nrt6bzSdV++Cbs0ZyKqzT92m159A6oQRKmuI5Q4epid0i1TKHfCq/ZvL8Me
rhUEpbRaETVyixQ3PJyH226P7Jpc0dv4T0Yjq9txPXgHVngYLk1ZBCRyqO3GWes3Y4/Q2DRD7I4p
0oULRRnwT5yjGeK6hq239BtasXQL1ZamMjcEjKN8vX5oj4EVivqPKCUA6PWiemjUnlvv/yBudQVH
kCg+q+Ir9uQiiH4zNj2sbgsWYZ8USv8eFhD7dyxGbaFc0RVci8pE8FcZCW9kEHC2EA+Jl0LU8m07
o9lAVkdoxX1Ej6a6pJ0FGNplv8LDGKY6GfY/4hVA+u1sbsvfkbyLZ9fL4aDhdVimlLOTpOo7/h7n
CvSoHLgu6zRfxaap09aeJEwrbIoDv/2Al/v1yA70tizz2uTXu3R+sREouOwKS+Dqb7PzKwxJut+T
vfO/Iysen4XX46oxcG0tQjE5OxTZHWLeamygzxot1gU6T3b0FGtInZIGddS6mMmnsCF6htHzw5Oj
fOdFqn/IyeMzF93jG0EWjWR/h3xJXzcf8FrQfykGjrLih21YWeilsztVWcoFodEPijNVXkoqn+ul
yS38XBldZ2n5evd6eKMrwqBFsuMrL5UWTkd0nqSIpclGRLt2bDRHuhvZ/eI52Tc77YNeIlpbGoi0
/ng+wZW+V0Rf0FIEM/FjZotfZXf4mhZMtkWVJjKNJ4mmuxnzqTnrXt8lBsZ7BE6DDcVu9DsyZHvi
nsP+h54q5eIU741I0tB+drbGzTawjTtbgwvuXoDwYwek/i9wqUCEP2gJ5nWXumlpGcnIS++7Y7W4
6MXE9hNI42H1M7Bz6AaJyeA0f9el1uWX6jFL1cmL9sfCF6Uak8l225c7mJ3JktSTS8wwqdBpVu9X
SvaMJVGrIMh8Rs54UPfEQ2ezCQefaMgH8UaQ/BiXrBIzkXru/OmDvkZYxcJS2qKiipfBx493nOkW
88dC+qL+wJbFHhGid+jLwBQPELebtP0kKdjvc153effQ6nv4Plzx58BhZYmk2ZVgfsCd+rb4J60V
6T5e6F8z3DJPJtGtdarUrYfOq3qBih8m7WL2vnhfCVeYHrGUl1cp5pnfYFC46EaTum/IWsDBic5l
BirDI3MfLKuSahFTbbJhdAaEnr0o/uWfaN59zCfLT7my6KKCjF+uOcYJhAeewiEedkJRFfKJJ/tg
bgTCsH131t0yJ5l26EqALcANGLDIzBWJyOKE/75dRencUY97txO/NQf6+upSSuQ63ITFINR2fEt8
ehvCU8P42LINt3GGRK00wAl8uYGn9HROIQFltaxnpV4Syy5x61Ix/SuK3+/STfl9k4Q/Ly47K6cO
R3egzzHPCQ/yYdllmWhu0C6WkE2oqp5b68whRsiagJd5MGrkOw8PwsauCXPIZUOaUAKGRTmJti4R
axY9HN6l8aMje9FKncrdwlP6MwPDFk6GfmKrvvaU4ROWfsn7r1quYrcPvDvA35FANHKflYfQI4tt
h/jDB5aDXUDGWqmaO9brvJxwnaEyvBDb7NmL+6p3Loohjhgg1YIVhoO4O/yZ8o0U1DCDiFyskIAK
RV6Pc5DT5bMQTpdr2NIvqt9gmo4zT3u5HgDnRQVa4N8NVkeEE3NyieZeeN+dhbdaRn5QkQQ3jjVR
Fg2+nzhjY7OlolrO1P0JWOuQYPupAVDyNrJg6hvNgwo3oxXACSjJDRzniH2EMKgxElO6IbtJ8bqj
iooAUx62m/mv3ErTuT+l3jLrmR2X0whL7C2AR4bEqaKUeII/XKbeI4X781BgUJj8OMKuC27N9zbE
s4eEYxclhIgLNbAKu/BVZNxdGkDZw3d/hd3qeit+pHQwJJHXg+Du6lBL8lls3E2r6FqS44zpT9Yg
KLqyc5nxjiBQWlEALHe7UEM+jb1n+GZY2xSxREY/dASgpX+29PWM1GOGgM73CL/57ZJe581J7zWH
Uaf+qpjH7hVz+rhAzE0h0cpAntNDrsGZkjCom3dnYDJgQPs5VmtfoGfTEAevJn0Gh8XeFui3rEvx
M3Pwx/DTpTCUngE1Z/IFnfu61gmbAwOjLzzGjcsUYaP99tmDaQ1I7TrbxwV33huMp2kqRGi7xif5
Eucgt81MZe4dF6fJggj/jPFXn27xBL+gm7cFBWa3LzS7o/YCjzQZJIDn2K8XSYWvZGSxzNqrfF35
OnMgNwYLBRl2T5ebrf9hiv0fVo0a+JtM7t4UQJ35SdLYZHBlWv2ztRg1a2PH9w8RzrryLCO0dwy2
eo42NeYPc/e1VyYMKJUgNPSjo830dkChGXlge4PY5/FP2s5K9vJNYdAUvBzUud58eYVYBwcZCB9N
meXhXVDcx7HpLc51zb8kmkWQdZ6ZR/7S5SUZVCkRByuTKAM3Vx6S+dSQf6v8CrHb2zP3h2uOeCEk
omEz9KZ9H41x2//J7iXdnfX97Q1kvNzgvSN2QW5aqvqq92rD2Q/Mj2+AUYLP8j8v4/+adsnMATXq
4WXsKXPako656FtKoXNprUAHooE8g3/boYpTmFzEaJxx5JuXkVmGE+y2jVQpdHsBOYa+XWJTDFwb
lV8ibKqg2Rc3SsLCvzySzkz7Wdchw7UFjeFGE4ZlmXIRxvslFZ2S65EqF0lL+lBmze3yneIfDEJV
ZhzCHHjQPgjkn7tL0zQsWOt8c/520kUJDMtBr8jK1BJ02zeNn5jsSGgYnTmzxqJIg/uJg8O8rReK
2tXgRXjBpFVtj8f8Ty3lOIt56moxogQsnCsTPSYCszJK4aLJXGGiDKX7NVN4d6l8bGpSjVJ1KgIr
x8hGgVhEQFf275r7op008mETdFtqIhFXm7tZDNMl5XSYUwB9E42G2NPVmuYWY3DnyOjpy6wwm9mo
W6PXopHsA1YYk8sIllHqHNdfP3iUdMwSzUoeMwPsI46cBnYSQPErfPLjdD05T6akELY77nnY53Mw
FzwmSGOYN4IOAkghJXINyIbrVnP6vGfrJ4qjp4SyHf+YxF6LUrKFrPP8RerBYHh+NVeJYiu98HWi
ZBNIElpNNtzREJ9P5QRn/JCdjmueA/+AKixq+uOdrOO3wS74LrYkv4hcYDx7g+hq8TTBZ2+vNFaC
L2iYnFcxhov1Hviq+gevUd8AROoYZYr45bbK/rc9mf4cg67l7GIFctdEuQ8sKHooUW/bR1ZA4OWF
cqK5teyIUnDLiSXs5nEwo+oajFjS9/F0WTuwmtiziC6ZUvIcnhSvFmcB+tsxDXY3gPfW0PbRfJZV
miEhrte/mksLWkVBX5iymzYj+uKZ9xJaIPIU4FsK7ElDwOQbS6wNseIWie54PSjElH4tqEcSLrQ7
Ng8YYo1mIyzNg0ZHoR0bpAsy3b0l79148fMPubLaPc3P7OjKrfSs8t4o//6Qt3zFfLwECZHIiTKH
gi3BiW8cL/kEy+6hAswfsiRPJRJ2kfj0/MKo/ewnO22OMon5g/RoxW5A1CdUHn+9S8AylQMuexAO
ZJsxAh8hJT6Wzwh0WVl2ZdjzsxYGq20lMT2JM1ZPf0iUTONqUhNzJMIjvKCDYaKsc79FMeHIZ8F0
84n/MRmWZ4pTuH/7lZKKAA1sFdpX7GqQ4L1EXbyGaJsXx5sPw7eY2h5ZRpNvvUUo6BclO7e0cUwp
LUk0TxMAb7A8Cni0rpPqqDWBXfRN2MUXRwPCz9auAYPS84pbDwFpqHv2wo53vU36rwFa6A9Fagja
iV6NGXFOFgOzjGn3qsaLVfNlE/65oyvilw/uJjtcKM7F7VsyAgbR6j+etaLh32k1oh5gY41KvDSz
K65Uup7EVent0koT28YUG/flYayKyhfTnPeZYV6kgmGthpJkFyfmSPoaf+6eeKcrBtSoKBJN6KOt
oXl7HKxX13C+1JmG3kXU4ZdSZJwWmICFnMwl+mwdTCS6QBWeXAOO6rnWrK60m7lJkSBOoIo9BcsV
I/alx81fdAdj/Jp/EX0E1MyGgtu2Z+HJj0xoVkqGzORa9oVDuexOMuqxb5ODA/hR+yQWK7O+rvrq
FCNO9TTDJionpeYlsXYsvEAGMwfH+W9xC+GtiSkvvleuoK2yzI9FMLBlgtj7aZyZHc+O+eV4MxUu
GH+bs3ZfdPPft6EHPK4qU+J0fW1+lN0SERFZX1PbHw7BF2+loTFKRKyOqNdkfbZFooSnWozfzFSd
aAFsIhM6ktH0aJa5PwencvGpByzTwJOiED2gniGNCtda09gzmEncYv6G/cU35zrIfrcvW1deE4CB
3xe7PObT8KXxJ0Ng6o4WXIzU3Te9ZSzsckM5WDKldiJkV3Kw9jFfSB7FaWjueIkzzr9ynWv6D0Aw
88ihCFNEpl7nWuAigxuHWcaRUCvsu260Gwie9stURmr88B1UYlytsd7A4VCYrR13qYIKHtnZ7G+j
zUGMXg7dJhmN3G/liZyVzcwQw9AcClX+d4Bg6/4EMa/y5W6hh20iAJspUqCTI7ldm4uPhHB0bQN7
scG34lG/nhMTFQ/Cr7OpDQkwqDLe7JvvEbEkO66aAiCqfrpK5CSMe919ey3VN8uO1pJDBL1cidrD
ZrHw0apShNdCnmYqK+kMN4CzHRI+R6jhHnNMQTV2iwL9IbYCDI93wbO0/bJkgPDqk6Bv0p1ZOcCi
dELq3Ja0D+ofrAqIW70ffOBEbIgMij7UZEgm7L7KS4rWq/zWfOiU98N1S/DcvjTEFCxZA2hEu4+4
wUeAPFD4S9NMdkKrOmR30SvNIYdy7O8oBz8kDOl6FHFS//caHOejgKOjE1ILR2/WQov5HlWra45Y
CF8ysppn4Al0M/7OK7ZT4v8ODO9geuG/FxLhVuTn/+Oe5gUnG7QVAVDIJ2flamQlfAKOMSXpnbsa
VGgSzz9nVuOXxA0kGIkYHWrr76tO4+RvHViPfwg8CCCAjiqqIsAGtowE3RawtpyKS5/xSMGQPt1g
fzvBP/+Osgk9KOQ0Be0Ny20JZ9J3GZbnANmU5UxJ1opnuBpDLlbPaSValg8CuIhXxqEcBPd+qLGm
p0iXMqzikdbnXG9vrNAeW5ROg67+cqcIdwvUXjnpxFW+4YXZCsPBjGd4m/5RD2niO5QRCbUzoNzK
tfyIQZGnSO3mD59NQpbboqa5vc3Z/mXz083tfyGFsHMZGdPvwqGEtNFnP5UmMKFvT898EkYaA8rm
kFwMNV9Aw5mYyiJeIMXdInET61cpiU86fU+wuk7PtbyKo14476yS1CNCTkAxRbp4IBtdBeoxlxM8
7ohJh/UIfDG8nd+avM4dUagVqPClK8glP5Q4WU/T1bpJ/XyN08fCcntVTcQ5ixlHHzWdgEMneP9L
0r7HvMWDxnJyROlGOWswewxQcpLEBjnyNCOAfIrDL6qy/FYYBBXI5Xpjg7V383E2j/WgRhzTM4DO
Po910GlQyYAB/OvCELCW8+Jr35vx+opO2VIHVUQhCt1clxV3Dec1sfCt++f154RIm+E0YXqH5c27
2Nikj05jKW28kHlbdn8e4cMCTsc4+1wE12msUh8RT0OE0Ntz7HnP7m3JsXb8BkDgc2EUS2dxmsqE
QMQ++PooAjOY0bT4N/qVh7EZj6FaDUZJe0+EqDJsk6UrJgI5lhZ2IqLTnLmbN2npCMxrKk3O/sVR
L3l88pSyR0YVlEery4fwtnGRgUpv7K00tlBfGvNJgmxLKL1Wk2Iz7kroyy0rIasVkdeeIQogt6LY
9FDiyqn/XRrxWVho2AUdbQO18/r2G8XxQP/RzYG/feQjmIg7ujRWcpT+YscFV0ehgLT6+qCfRHhb
U+SL1zpdGqXnuJiwrm4RmF2Rmv5rcqb5ds8QDhWC0HS3RwmPzF/qE/tsd8+zGYiHbj4XpeuStr/H
j/RgMyvXomh7fbF+e/CGojpqat8rsYH+aYtdguS41UwQL7W/3KbvVHA5Fi9gIej5rlipUMFluQJd
tiTFveBGBltShw6wBkCXJTeuPVcroaADaa1nY6miVgyZXHujhd9wNHJE9uWqp85hHUb50sOXQaqT
3xT6q+OeSMl0SWZ9kP35ZZC+OrU7jW2xsga1wpQUeknFX6FSwkTK7f0HCDxxlYA3svWVZmn5Fe9q
5qFybnDZuMIRIUNCd/4QiQYOSGUZQVVeN9vbfi6Ybqh39zYekIg3/X1q2CAVn6L8dwQr3ulSMN/c
xJsOkdV4J8z1HQDeBuhtYWECe+9s1jalbuFDsfS5KDFeT0OSgrTxExz4B2jvzzu3+OFgY/UWqjU8
C/H8LxffOMko+WEYAW/CyIdCG823L6H0xzYZbMPLjLYFk0+NhkVAMmhI3/IZWXZp3alNqdlURIVr
HwZdHhcKfrsPdAdFwgDET+mKZPqmUwpRPmugr+asIpNjo4oG4oPUVyLNWLx3ttlGUpLcdQSy5SWq
SiZYycAyxuUMwW4WNOI85o7WL6gOy9/JCZ3MjcdA/WEW0H9oIJy6RXvpz5RtgdV2VfMbN/DSgojD
6lT2WdqVf2FJkG9lfGe4q7CG2UWw5DiYCxmoMlcdkqsu6wVtUtprTLAwhjkVJlCMER8gVDMVISiq
7ARP/HWctGUZqu76HuXkXiDzq87t4pIpcHjStA0RgAkFwF7s9hFZ3wqBZpZgRORDrMXMisSxADXz
ZWjI1OHOfR5rBySenMSnDrmqHI5t+Yv83LB6TewdzfXTwsBObsuJYiThGe86wDrJ2EY+qHbZCtzk
Q4x7WOaow/xSCPVEtJbPQHTxXxPp2I+nauVzFwzRwgRrUx7VOaz8Jd9qnhhRVmuUkN2woVPA0rru
MywUTQmyD4P3+sUc9n2l2SL6ot5uW37nb7hE2wjZSliajI/42/TGtx94NI+EYymRUGjnJfgfNwDJ
vmhTd7Pg1O9XlpL8Ol11lMsyPFE9RKKw0z5b5xKuKf8d7ZZv8Uo2e8QfnulphN/0Rn+nTyJ42BMl
3SFirkcIRTQ2kENbb7EPRGM9dZ/2kPNg3u7VxAj64UQErFi/5SEQJxWQrD3DVK9xjXmqls0j5FQ6
YyBlDYPPn3PjJLYr6p1Vylb3x5rAuv/Kk4QTNEg5dg0XWRgG3OPUcugyL+nER3ryrz/LCL83rbhj
KWLXNNkBDiRVX6A2Z042HyuUSN/wLGeszXstXpehkklXg/osGxguNabGHenWLfBtWsx8zblHDZ/B
TIjyOQzo9S6YUA+M3bAO8s2w1KaTmFvao/vwUOdVhcAn3Lmi/UXHTyKhMdKIbqL1Jt4k7leIm39p
PZZbrwvp/uhKjrhiw1ANMbbFDKTd7dacsnWx7YOXnqOd+k8e8YoFHYu8ht24ZMwjohq3w/J9N/Xh
b3OGHdloletVO5sVnl778L58AaOdGxe3a+JtcXNMJp8O89WTK4+jlseAR8cRA02l0uFmcS+tTP5e
z3a7/ydhS6iSM9bZhvFAGvsa/WjNcHyPSMfILFx2OEPp/yWq8mE3qYn2949QVCcHoRBzYZmAEpTS
6iEigpwN8tIPe85gbJZz/YAl0c9MjTNGKE90ts8qn13RT+qRJ2wsCKNTme0jhvYeK9TacNI+5XCQ
1yo431p6w8zj7e05KXjkbY9GeZh5HLh1OGQntM5oBVkZdz66mHFInilybBXc4tW/m8wLLpwt67D2
QbFWofHFleh0JaXRjcPfVXl2W6sNh37Ok/hQUtwV6tXzosAnlubgHa5l8Rq42AubrFGs51usfScc
oSh8mMJlgdH2qWwj+ebszrt13Yv7tZ6/WubkgPkaBNsHo88E0aHcL+s04SBKiG7zjHIul+XVBBTY
4CzXXwXffOAywIlPW2XHQAO6z7/Nghla5mWX9zJyYw0dAo/YC6m5kTrnmw98QjEdJcafL/mXFTnF
Me+lR2ReFPFpupdWq2jS6fvidVCJ7j66HGZiQ2pJxXFIGgcZm+cy0wHyEUJNcchN2fBoRT1P72NP
xpu4hxSGMi9QbZ1QaIm/5yHiFxDqmySw0aVbxwe/LRVQuIHfwDCdzpY00Fe5h9O2HAgIrwhYeCE/
3iqp7uZWRhOC/ubOIHJkwsI+QIVrF9l0luu0D0JP/rZnRfRjVIidsPTN8PuPDNp7f7d+myMWNyQa
6toiOKJkCRuPcWzQTdrhSf/Oqt+BWCLav6hagma9hfoLAdYS0jNvt7L8m0h9adlm7hUarRsyY3fZ
Sv6LqS1r+b/psjJa9AR/djkoPrTWCgzFH02G3y3Ps8QYLcQln7pJSD5AtojwFZZWUAiww6oekodw
jnO0Klm1eKD31UpVI6cwKbFHddtlujdI5BTPDbES9IbJWPxoAprGeSgnhF3cnnmDX5pq5uiBfjRu
7KHmXq1TGmItKSrO0Jvsos3PzlQhw6ErJlNKBaMYf41vBe6aETjDBTGBFIwV7IUCqKXMRfzqkYZx
2fcj3dWJjktVbZqgG0blwk1XXg5NGBOzLRJEo8uRpVcvVKBCJdtuVVaocf18EPM9aTeoRk///1sm
y/guO+Zcs4UYU7GdPl5QHTVvOBABFMr/ZIT2OVc9ld7mYbuk5IjmfiSiEhJgxDr00ds8JHHKoSsc
tiVen9UWWLXq93SmjrTCkQtuzVMCKYGkiZZwPfXKrLlIFINWrOuyNQQfe9UnnQ7rZZ6M/ysJqkCR
c+f+so3BkpN2Jhtp2u22GYM3gmEnpN//rc0O4Sh7cNCyJdCizKDy+4TRrcOpcaSkW9RgIHx07Oyl
NChrMedPMtBReEct2ZAfmq6RMfqbultSNhAFzl1hTD6NvKL5XnGBCg/UOtPjmn5QwfpsXt4xcyVi
I6iMbl3vXzvO6wBZ4OMDlUDzDI6cC5FuJkR3dQYGdrcAFRgplDPbvZvhLOno3qu4eDFqn2anm/y3
RTaum1zrdkge0HBYlkPtv8tGLxc2DB/tERZ/J6AmPqQeFgBWnqTz18dMTC3hjtk4cc4Bzn5wzU7e
isNLRG+Zmt+CEZIaXCqkL1m6Dnkfdj+HM/56hQT3ayvWp6a47svErCDtxH/UY55sdt0Zp4v8dDRq
fieQhEk1nQz7Qu7fFIbzJ3h/iJhUhPr3KYMzrIkfXLK6edvJFsL7TJDHwI5I5wX9KPvNY7Y8kYCu
lE7g4Z0gOGaRlOwNx3zo4WI7tRIsqI12nJsw+d3IcFNBh/vMERQ/KuNYTj9lbeJDH5JqwULqUo1V
9AhkBoEc42X4/Owq7HiAjb4pIZRICQ9pw2HJSjbIQ0mkJyopJIYitzhjvmnwEsR9h7HEml2pfRxO
YDejJE9G6k21pl/YHaFSbLYeyV2ujv5VmqGd04nBkfOn2D9SNedONtI8FTRMRqridUQFj4WyE6dn
xCvK3Kw9VWw/Bw4Zq1RNK+12KmrzIlr3hqhWNVS5SSvDPnJPma7x4gTQtYRTXoIC+5JuroEi/7Uo
pjvAFaoKM9xpJpVPvmrsqLDIZHVRcPjbxcNatuvACzUS5JmK/IVCQFRDr9QBI+ioJL+nAUehGhnp
1zyMweklGctKstb7AkgmkHVN9cRp8S8NGtM2tCVljYkGXfvZOTNAb/u2ZvApoaTHxTGwzHK7APS6
GM2N8i6KtrV6AxjZ8bKRbhm9kAuGh2XYEB38Vqywr93aqEgsvIqcGFK1LGlFOgd7WZ2Fua0EkDs3
duHRmOkx7ekhnXVv1kW2vHdLiJYh7JT02KoERffoQcJrRJfPOM2tX+iSdXS93YWGM+ZzFNPGUa8x
IZnxhNeUODuPZ2t6XGlXW/0JeVi9Oyc1hxoth2/huRT0HJzRExWyZLWuboT4RhX83FQ1zTHC9q8n
Epvf0A2Vhy9mVvsco4l+Z/xpOn6m7Sc1UireczTbp+bJpQLe1Fw8lMDH89XTY0w3jKsJs0W6P0jh
CdXc+cAI0RJcQehM32HAkmCthY25bnjEYd+k6ikDfe+aLv+V/2I6207daAWS2BbGDcXjz3ho1YrD
VosTdjlcVlA1gfv8GOmeV3jPK4JLdqZr9lJ+jlGQaKNuO6k5nlj/9a7sk9AX8BHQntAMRi6IgsJ/
L5/YRvnKbpGIn+fzv6sof+ryyqRvzUCvI6csui7yqh+Sp65qUTmzxTPHTiBObVDSvwHnNu2meKll
EbtSj4z4iWju9Cb66fyV4bHaMz7AYBmPI1SGLAK3FFtm8DH8Nfxpddsr4mLyzhEJQJBLeYMJkCeq
34Tn4jiEha4gWh7pBlc2F8r0pdiJ6EYcMwhoaO2Lc8ZXDlBwg6BWKjwPaCkuC5UUkNAQinimUYa4
OLpQ31C09zs4LjZ6RKvCozu4wseIFVu5LVagStPh2uUEMkdXCyZYWm8A9ImLyWsLeWP8Gs+hNkfq
ufX2haQbWrKz9ZjWkBJsPqjF91GDmvmmlPJD7J24xpEEIpQv05epUdyvveIM/V5XHDWFQNq3LDxW
VHyx/ztBItG+KqRZwduYZPO6Ckb4Wc/EPFGgDb7fLyisPKSQi9bv0fQSK+qbQJXQHbV2jyrskHSH
MqUMN/13/seOMqoW2cU1TU/usQo626jkjYNj8jnyY68UugcrNfuhtVPjMlK2axzGkROT3l2BKkRM
PMv9GnAPiWjF0bUPBQzm8TUD6H9SI468uPWvhtgAX6G5euzoFBgHuGovdztPXLIBRixJ4s7CkpUk
SHJRG+qgtLX31ACeAOaAYCcCEm+T5+WyxjXvEdYVsTn/JqZLh+I3y8dBNjhnXTSJat81281a9zJE
ea6fKUhpJUjKNCbzl0Y3c4tHbEf+UaKaFuZoV/xtrEVdFH3lOqDuEKCqYklh3eGOSLMw8ZkKzibf
GSEH9fGeFq6oWIZZCc//mhYBR7sLNUHhNZceofcwyMadTvDw38K3MrfooIPlU1WPbERI1Jsmyfk+
KPSwx4iQDccXqglFFY+5LyDvkZ0BOSBeez6vVMXXo1OO9NyhQljUXYiIfoz8WemAxxJBHk+ya6dq
LGgGnYSwYNaU4hWKfSuDLbZY1qLl32Gy0VNeUzwspn2q43FJmToILGqT9lHS3PN9uIfpTfKZaUfe
cy3VP1uTLzwkMg0C7XwkLr7WbUr6wvqchSstGbr/6k1frbBARZSMid/ZoWxytzTJoa1sTxKRzbmp
zANh33NCQo/rEl6PFz3x9P1bEdXrdib1jaosQGoRk1Ak2RJL9e9hYumOmRPqQ6nOvSc4YcfXKOa0
zGgLIerdPSz4GrMjuAD8C0aMlPRzGwpxhRbuAybWje+/PorPH8KTd6trAa3zXfR7UlzRmrijhgGA
LLPLsyDGtg8vuuzEZ4YVlE4KEaDIK3NSxSMOd33Fn0Xipc3uH+sOJNHigtcb+1kmUGd6Zvqqh+uk
AjIU3WSqY28Fqsm9UEYLlXWJM2EDGEJInLlwxRA1BFG47Ds84uDxfRPpHIUEzHVVnXNNqYtC2Bw1
M3IOoWsE9c5pz6k/asfZzkdUn9GvACfzAR3HPphbKiR67mS9N+7HF1LTr4qTJll1hy+0iAtxbJn0
xP3oCLHetj5w7fOGIb2wb/ChfiZfwBFTl78vntI+i6/YQv54YEnCES9SmdX52Jog/bBd0lI2kqTZ
tq/QQ3UDcL5fIhkueaZyrd/KTKc9pOIa1MfF/VVyZoVyz/YRhPZeqeFJKCHMCyL8+C2plqQdqYga
h1x6WfwxPisimY/1+wB+Ke4RqcW4kZpUHh0sFPTEuqvfEYDjN0KayagAvxFA+GAtSPH0a8o8tMBc
hItyQOMQYfi4CiZLIZAF4K7BW/7NsGWcpIVTOtHh0oB6rzQlVHGn8uY0sk9iVGTA3wrREDkneJkV
GJlFPlhv1owN2DyIWoFQzPn0+q8KygDBYWZmynqkxJUSAJzffubDiGFegvGWyFzzYPvnBJfTahsk
q1RrdBRiL+zbQObpG9P6j84YxF5hfPl/lYlJ7xNT8js8MRkXy3mmklk2uhTdyLSYJOWWYz1oVdvw
PlJcIcAC2FngrAoXP2p8AVfJOxP4HbpRhS+3OKbMW3HPaVL0Tus004UQQXv7bUDAdim86uGjQFUe
zDaFO+qACTDStSjg/9X2uXkzHARR6gmZMqUVmDZ3um/rhZbyaSarAzIuAqRG8P8BxDJSToWcNE+n
cNWYXdvrRd/fWXxZKKz/xp/xCVl1J3d0a+fvzLsufh1HHbjK0LFoLL4VHUMMSu3moBMF0/CcDo79
bVU7R8cXZ4lgYhAJJ9N70Hp+X4DfYEIF0ttxZ+KmOv+HVEqNJfkS1G/Mkc+W8fLTU1qZfI/yhqXk
iYg9NJ6jTPkB4MyOcWda5o2RhynU0GIXrqmDpnFM/V6NyvCBQEPKgQezXnSwdBCkk0acmbOUDrni
wvBMplXVRE5zQWyEef0qlb6gNl34+DlDxd6c3K0dg5EIO3Fg3xdijx+mAibKppwOa9jG3uL7VN9L
ooBGPg5c8siHY6l8fbuy+zINoPJAl+KFghjxkKA/tCoaOocNqsOuPeEL2q/Tm4rrU63wutElYysE
LBrEHee1E5f/dlX/eAeVh6xOkRlBxDI4loCocSyzkRYFc7nN9CUMp8fx8TSLHCSu0X9CMlZCNVqF
weEB/BGJwJMU9XGCmd1rjtrzsSMsVBBwMOBUL+TUme+QGGUFN50FXJo+vO5I+YwWWVcfGs+Prgfk
g1rYbDKwaMB7dij+nghu5me5ER4Bs4tCVP3bLTIcX6YEdYQcuFslLpzlqzOjXJzYlmvZ49Cq5OAM
vKbwkdDltJBFbmPptzdsn0dibuqkY1CLwfT3TrbDHOVv2KUbpyikCl6Tb5dYcJwHH3NWBF/G9pEX
xYBSdR5Otlh80XhpYjvJvpUlqtmtPVRilbo+nHanMdT+LdI7I9HXb08RHQjtjscU+9cwaPhD1nzF
hL/ExvuEZu1h+btov03DeKT0aQHruTFQ+jSok6TuwEZ+kDvWalkwt87Fcj3OATytR79twym633Mb
0Zd+sXcE092RQ5eZmNSTeoJZ4wsnzGpC6Vr25DD7P60rprZLKQt9gXux+FqiOeG0sw2LYnrwNDae
f7+2R6uBVqyXPI0p+thUpbz8c8UGfZuLi6tdBbmRQGNZaETeq3dKZ22QhvSq5APpAc4nmoae8DgH
9UM7VPr4AzI46Z95nyuyOP0LvYTZytTgkNVCMZP5ueTV+gwVBknPW5afiNclLD+hUfxBj9XRROa6
eL5bZ1ucsvLEYS4iRA5/qij+UdkJlY2xqTMP24thNIW9Xfqx7VavHLAI7ZRqV1LeaGzaz/IkDPh6
/fg0oz3IY4FonsP1ZgMNOwigeQR++P0onRIClWEDSu9aKPVlkPYPDkYqY50xj+BbP94wBscbZdrk
IYJs7URDpQ8MK7MbAPyQapJ5ROVVM6DKu858XUcOBBH+xwM/3feEkmD12ceNzP4fi/7ROaL9fAua
EtVWj/Yb6qBZfuOyG+RJZtkJvA5rEm0hm0+ij5VRqfIUCIf9OfGD1mR2TzKHDi+ZtnCVwKQodUFD
Il39q5vOoaaY88ejudRpVKxWayjyCHrzzij3qYQeSn/1oU5pwrOppItYJChmtVQDQU1O60AQeX4j
sIGc+Smtv9J5Y1fMfg44uA8di7egEZ+oK9mp4+KkzetpPek8hN357YWBpVnTV40rPt5G+4ZU0Pez
wvLBZvb9ihiiLM7LZofiQC0ZzHKBEvmF2YBqMbZVCp5I4YwMSfXL3le3jV3eDNkPeyBY96jtf1Yj
Sd18qRjGl3qGWRBM0Gqx1CPyfZVXggZc9k72ghqzAQiQ3AGUC9irzDMuA/PHj6WIT1mUDnZfVDP7
Cj6r4ijJ2aM8ou4tPidpbmi+memfcpWmhD3AN/tIF6H/pBg3iEdAoOHmRfeR4yWC82iXUQAA4FEN
MEBfB4Jr26T8ZBGfU7WgrsTsauPmm1Y2YTIEamr6h7Oqa/WwFdh2mA8g5QLJ7aiRq6pRBOWGQ/w6
b0GNjqizAjRkTyRzBAD4vQPiTfQl9i/nrVilT8Ax2H4Tnz4h5NqWDhXER6WtOtfEIyIXcwyIacEx
aUQJZUmcyRRWNKtT6nXyq4+9J7rxOzR3mcx5twzoSZTukdbG9sAMFAid5XrY+h4UIZGQxdzV6Lqa
TwsjvkOmiTAxSh5vRLha2CKav7GlZVxe4G5u27hDiLCU81rCCaNtJkExtJPhBb55PumPgLsFShn8
sd0zaDDnaXFVUO5UR3ckzPcLOO9xr/grguuzxEYgN0nFGthzjC7uXEv2ll55u/2J8WLieXA7gyiV
5OyUnwiMa1po2F205ok2fjvpyVFGoNeLfKbQZ9yh54qHoZ9JAMJFYFG2FwXzP985dNGDmIQ3SxZf
mSzNdaOo5khvw1L5FqMKIWkIb6EP2DvtEdmYn4Pf8m97yUR1IlhN2ZgFqImyz1zC65B3u3bTG2Ne
O6r0+Ee0abiLSUcmj9zjSyGtS/UCn7xH+1jDEWhuXa31v+09jriXxl3R30GeYOivT58MGRjloC/M
zwvqm5Up3uqK4NI4vAJFKK1AhOllXIVkOFjfOTa9Lx3at4UQxAa4De1l/Q5gODo80qDI9jy/4qmx
BciRwJ0ZV5Jg0dIJTq+B73NNcpWOdoCFUlGyLcixA5U3qNJWvRIe8vWu02oIjnCX2CBzr2vAm3Ly
hwreUo7+AeHNoiWYxkngmgYg/dpjenLaa/3FEq4e1dR8ipOHmgcZ+P1ShkVzJBcatPWuJux4kaVP
NrMLJLNyGJVnRE0hBi2/nf1YC85sfYRyv9ND4xmx+3UNTET/twINrkR9HXwSGQwXyt0d7N38AFz0
VBdCkAWG3VoZvpfMHC5S6r2i9u6Kz0flD075YFOQ0nGYNLEVYM2LuPUFqjeRJnC4vTZU+wEP5np+
hw6ySrKNMZVoh95AeTii0+PSHpmjuxLtUbZ+tedYcNtcuxIqnufHT/OqgPK3GDl1aUPFkYFX8+k8
kAY8+9BZDxU9Mut/Mr7+J3I2B6ZYOKwudSwaY61rcYh80XWYaB5v8WEa1BR6aWAOZzpYmCAbwxFC
Zt3aLFFdlZsGns06N7aw+xrZaOMw7kgwqkCIjySiFtefVSbVfK/qEANpik17mbt4HEzE+Rj6VhbF
8pYqvpPRkWj5Oyl+CnRjweD7HUAPVC4d9FjcFbWaYIVpYI48OEVnB8QNAPJSDGifNdgtTK0Dx361
JZ0H2QsfkiynPtYLgRERJQb5clZz5zrRA1rQDouwcYQi3rmgsh+OHuelpIYrRQxiFbWYekpSMAeK
86uSxP0SLHH/nO0+uSsbOFe0wmvmq89AScmu2JaQf32HsVhnons/Wz0nvmMrL2RBrjNUW1iV4N+T
+Zo92HRPNHD5SwvH5HW4244at5ZQBrAL1lid3ufNaL2AtFzM/FBIcsMupevCn6xwMU6KySk6wm8Z
txSy3yirfF0yULxcxGFQDYaOGCyziX6a7QMCjgucfP/CXC0L9pXL8uAdTMhsWYTw5RwYiAgHJ+dI
ZLv6ZrYRyeamLnI0KJZoVqvJPk3pjxnL76n4zOIJ4LQm6JcGrDTucWM9Y4b5wdWUpMVsii6Vz7Ig
O4xZ9f7gphZhEpYFIkDCFPBb+/9gSA7cMUbOJI1RTgd9yTiaCCe8xoP67eLqYKZHPrG+ANryJ+KC
zWcGy9/M/vBLWnYCDzNCelWYsM+yl0CRgkbBk6gY5DnjNU7DAE5WNzxfceIJ9I6QluZHHEU1VQpO
nVLM+ieIwcY32+bLOFfgBdwVpQSny5zq9Bo1NZc2tNIsF4yQjwAoHoqSJUnUTF/NnKWm158Oz7Eq
wPsKxx1GMpugx3cRnpOV+nqQlHi4ai9h9et/vzrZy83MKaXM5p3HxL5DRExuY4ulyxqJobuugTfM
APIM5G5QiksZNuutMw+GxfaSngdaGBEr2grVRnNVUwr/LrapHl1Me9b4DdiCGfgYYv3kwT8FTI8d
AjK588Pb9uIcOrDxU4e2vUWTQ6k4M3lQc0qSAwnp+jJ/xxyWiRamEASQ2diOHA0leHY2Nv9KLnej
s5oFAG6pIv77ReFDSotTrpfSUjqp3n1IUU0jtZ0GJbSz1HhBypNhRsrA4HyCAaTph5aadHTc53x0
qNJuTCmE7+q6oXBBerQFjvABzGeTcPzuUQp7n3vTGo6JdyMhjiLR8le1WV1M/se8C+HFOla8GAev
dWdINKo5r8kaTMpY4v2QuotOJDVpVTS5Ck+1jv0s6MO5BQp/H/DLpHGXyErxueD5f4cWMK5L1GLa
svJ8XDfA1B77Zk2kt2gCQdcvpxUbb8CPTYT9FOTD2q75Wnw3LbuEUUmUw00k4zsklKRwUBFaL86r
YQZTDIwp63hoFFvgTNW7eGSt2S7TlXsCxcee8PLh2TtpfC8hGuaWm4LlrzEWYf8FZRatsle+wxWB
l29zaCPAZhRH0pZKyE3eKR5s3/hCJpk95gXMimtLa1ZcdAMWZn5CJD4tLjBImqul1D9hf6HbSn19
TdV9xevJLxEJjuF9GXiMitbcWmjTBQpEfLttDpcWV5MwHK6nx7r7IdhUtsF2lboknjK7SoLnmmof
KwN3ZPN4qLsC+qdw/hiG42ofytSyft7e9U5mZyMBWJt+WGitXGXkwhROUrDuU9vKtithWZ1ZQaZU
Zt40wJ/LWseEugxT2dURw1wZiz2LLAmmSlsSxyw1xXOTDfYX3Q/4AfmaBDS0WkkTk/dx8DZQ0qFq
YcPgb3HCkNPIpHnp59BCSG6v18S22DZwKP6Qn0Jygumql0JUsquW8LIzyVCDec5FWJdypyQ7HnP8
REIxz9LOCxD+YkayHxmGgPwFTM8o/XJzinIeJOEwvzQntmA13WMGEzBuCrWy0KGk8MNtU+4ZNJl7
Rw+YfA0+m9vO+OctLE9O8HTcEnHBfdvt8V7djA/4GQdrkX7vdcJND0FCFqKN6TV+K9JfbGblInNU
BnI+72/QzOtNLAxeU044c44+8U8YNnTe/VpArFJHVE+6Dp+z0U5jxQXNPCJwO3s8ppmxIgPxMRCp
UM/THOwip0EyV7uqUiAMQJguG5sk7CTTT+AypNtBoLKLiM5pmJrsRL+gzBAU0ZWlRhbkiH0gX6zW
xC3DVX0OqYNMNJiijc9HXNh/57crQkrYCM33WfVL0YfnjhsD0D4vsPuLJj/BmGGNa27P+eFoi6hv
aFMVV+gP8MvVNDiDJJmdCT4rKrXhiuZLBZJitUm5/kojwPQopYFQicf8NMJOsYsmEDJR9+xP4n7I
LnLsN43vOEGL0P7xlia16MGLbQjXnSDVUb0ns+lHI/gK66/a2dgb5HL1raDsDQPRqWKxz/8rTYMl
KO6TLbWu9PQuYQh6K5nviB5A1zmXEomZ+txLqMqHjCMI/cQivFShD5CaZ48IUtCyt8KpzKi+LoBc
AD52fMOK9CShxn2K0MdkTYOlsf4wo+V6LFm65j7UOMawwg3rodnOpHqj83pKIAPIzvGAnMp+3kU2
eeyGooq51ZgbjuJcKNNU+pS/+/TPmAaGTWUmsK2leE9cBIXv0B9NvVrz4nvuaYKiD66fblnfEvAl
SC0stZ9ZbvMjimdnJAPVUIecXZ6qXKKB9ziKm5AL4p4v9NL4fXKNoz5Rsr6eLh9bv41cz/yGNGM6
HYMBoKkJGooWT+1KNhiWg9oUz3qOaaxWoOEzRfDzvThAnH6fO2lgdb+XEQSvAmCdoPGYfx2uXzAJ
2r9h2Tg2GWPijAQYzpvPR+bcaq60LJdIfobhkJ1EDY4GqvYB9fZllncmxuCuVIQ+JlzZ6MisnPvm
RLBK1R5tl4QLu7LfFWu4DCX6Qi9Hiv3663NtUHvDJelNHIxun1ZQN6h6TfnwjfR9eUAE0U+KFiwd
XAVz+HFCx4eCmE2uRSyBRWVGwN/6CB9Cq3AYonM6Vp7gXYmnuiqZUI8ctZclQnxnCNwoljBFmsKg
G1iXWdtENJ4uNyPU5m9H3bevfiGDM000KIBlRVGELOgQFuwDjm/lSZ1U5SocUN9m/2FA1PCu16rA
31EaoG07AB3EcYbDsOaW931flmd5M9yjaWeb8qFqdyubkgLbXCiOF3ALM8AHr0gKlViT9ST9brDz
rdzmMKDTieM1nkHGRj9PLF+IhE+QU9MY2DcmWO87s1Gum4E8XmwKREUZLrqDOEmhlhQa080xWuJ0
UhLJNsTnGULHEBBiCwGYlWIIx8tHfQHpRU0xb9mULRXwdrM6tsO6BkCECoU7pcYKo+qV2JSo6D2k
cC0IrW0/zsYnvXGJ7fezrG3bQZck0btYHk1N6jaZhpaS0Eyl8rWQgq9ISnwBTMVZomXE+ikr0dEo
mmi2T3INR7b83pF/iJsBP52szVnLEyGZ+vf+fzzIWpAo+qHH9cmAOlzvYWAYej2sl/w480SOeUmW
YT7Zm1WJC/Cv32k5Hh4HUJZRppQ+J59uZ0nWLST6Q6S1JiZKEVAcMeojvUBw0HA00obtxevZ1rT4
0sZ9/lCLOlVb+wriiam8VsHGs6DwIbY4eEe/pM2C+S1byREipru48HN3ZPNRQ7xKvW/N/BtsAowz
SurVscBAMoN7vMkxuLBdPVuQxWpr+jQfjOkGjYFmwNLF8XLyz990bVcVE+1boZrQFqK9zmqb1KOw
zDb9uD0v4P0C0V1gIWAbwVxbGQ6ajuOgGS75lgZ/mKoI4IctzruvW/cmMBnfEniralgRuk/bI3Ye
cEJNYesUKjmnxRIEteA2l0ZLe8L/eBF56GCuB9efVBtlIW9/Jtpa/AZXA3MxPkGJxvyRjAdIqmZO
Xt0DSlt6Kb+k2qOKoNWOlVYxXcwolksd0SPUV7Z0brVmnTG/0U7uY2iG3Iq5cdEHZE95Ovsqst+t
zMdXGjQ/FV4s9oT64bbRPRvaHNdX2fpuStcXPMie4NElTdz8UPi5dgqkcTTya/e4cEijdgZxntXM
hLv97WCs0tso79lDOdd5JCq4K+3D6/AFmRLKsb/iUK5qx2bxvo/pQH/3AAbRu6mVLbuXtJ4kQJCp
3GQ/PP3SVNbfLD3kK+qKcADdrQIAh0ZJwucQUMBGIgKhQSsKuMevRwxjmu9ErgZPXzuMikPrMi6O
MeMo1u60CF5pBOsjVh/Ah2UKLEN+2AwsdM4mbfgdvVWvWRQpxEnyIWc6+btjK7SmsaBhbtRCtY27
+CpznWsIAlVa/Ile4RR+EuOchpIjgDpEx9d5XX6SG/EoPVBNWgPK2pLY2gDOpcNj07DxUdzEm1ql
IgUGIovPPrE4yIskqKbGHzjB4RCCz4Q3C/ABgPbPcgJVbUKm2bIcrLkw4xCuayIB30t/MWdqWKVU
7IMU18virQG5vBsgFfyvNCY0mcqnGNy5LBGEGhpAinoc1kYqCklmTAfs069B+eRHvnj+p/0PUXQI
EAu420J5MCLDvMbIMgPHy0DYTDti/KKatbdEDh/jh6HqOVzs/GBuLKd+A9xojHKvPqOggEmZ6IW2
F+baq7tku2wzzeAbjTwpwzkXxIzLO/zQWXj5EHoo6kdHpPY/BVaFmOhcln6NiVJvVaac1KUUO0A/
lrFFNNoOE9j2rt8bv+r4MIiOXf4Xfqq3X/Xsshx503uH7UKQhNjceIWqtgEW2TcUkpTdvRB63cWU
vq2ksN5qVJ7bWMu+tCHrHHxdzoG5b4A13j5TrmfSFW789V5nxJ7bWIXuOvf8pwoYKdHsbstZB3JU
WVt0yzfdxs2ht2hpsBHDGk7qMSkHfbjkOc603y7Rkt/8X9/NoxY7wIY82pUb/jR1MBTGpwYRyiP0
mrVoWw+Jqd/UOuWhlx3uWLQlEEz7HCVS5a+ni8+uoorNT805pRgwzq3biO3oXQKVJNs6SbgWAYHu
yiKeXO/wQOHZcUc9kVrvakviVt3puDlS/ZTklVdFlXHVH8bcM2Y2Q2rauUEqFa3xFki0aJWuH4kU
qL12kStpbiCMZU8KoqhFiGq1XJ8ya6v5vcKQzoGuC3axaIxHqtvoOxDuNVcASKOXBGNoU0dDYtQo
Uxh+PwZaGgufno1YKogpSU3RNkhfXojV8iBOALkdPyDCCg6Krf++zRz9aaKfYXYiFDR6ojzEwo8T
AAxU9z8SCMBUXa8LWbukt+pY85YO8Ts2Zekj7UTM+Qkif2RLLfQJAtDM1utN/n0tnJibgtOgEVBI
R3KwX793chnfbXP7Rpql84XpkMlIigd8vrZS+er+d9YZgzPXB08q6QRtimRUmkswqqpOvKD4cZoO
tEJzmfCsnfYwokR4HySnx5FCuCyNYfntIGP8iI7CtZj1YVOJtLPew2QNFv9lpJWkKJpwsuf38ZFf
FeoOqw6mOCLJ5SdeG48Qdxi26x+I27iEIbOwWUvzKokZ5ZZrvbL+pf1QVra+H9uTF/v0vxgS4haC
Jqlv9oP/qjX2LN0t0NdDLewR9wwnCMgHB8/sP91bAILe2OQ//jFIxxpAOxQ+sqjmnIp9CV6fb9oP
xJgeS7is32cyQi7fefK2rsjdfYA95UMcea6GIWI7485MKSYeIaBsJj/AQLzgOYn7bsllJ0fzgmn7
5Dck1bZtc6cZm9MAr3+JmzsKWqg4dJv6Dzo+SnmJ6jN2ADQeZo/LnUeqol6laEHpTQ8pm9ZtzhFG
QRJAKdFUJw+WcY9OqlAXKyRLeKsK+LU2Tsun9VVf9odCazSvJ7G6jf8vtGab/hLBNU4jqgUirNUn
3B8iSwhn5ZeW/38I9/Ay8coQwe2TbEJQcMyEXf6eVeDL7mf3vx5YjL7sTAtWYVGiFmrAQq/XjMe9
xzxZpOaGgRSq2oLTVnlwnV9Ua3jDmRY4LH+q2nlM/jCBK/y99MxDIwsmOdmVyM0boHSDql1a0bgT
tCmvfmdajco/7wG/sdL/AZFiRWP2bpkdu0C7XZrpc1NVqhO+54hLjAVPL29gsSAPR55X+cG0f9v+
fQgQsbhgspzD5AYVk7UoYUHiFQjpCdmCEI/19o+h49AJSvB9pTAODbTQI1Q3xH12JLbFNjiPEIIe
nzqjQt+JKdrjKfnQo1Qmh3x002uRByKHVwMOLO8P2KIdJYpfov38zLj1s9pNewbz7GxkU1d4wAyF
sjrWbi2A9OWgywQplOuOUpjIRkWrQFCM17G2e2LLi/a0dkMLMzCo1eYQYnC8XDYXkUmB6Wq40Lxn
E/BzNB3LtxYNtnoH9DvRXfD0MJ7mWYP61ppRGDCk+H+RoB1cYk3Z4Uj0JMZMunBKB8JZF4kHMKfr
zpoicLsr2eh78Tlbk66p6Ntd+1yxpUjbnR3T4CCGUxC7StCp7hvmlSLHB1FoWHvyWc7W3WsezinV
3HWuqSeAse1Vfo3nGl3X+5vnTP1UuwJM5d+Aup2BtaiHi7abegvnLk69i99q8pEh/MnvrxEOUaVP
FNOiMgpXBakXTFnfrX3JNc8vZL11QHmvfKVJAb7M3M1YFderXQ/d78j0/q4F5Z+56y53+6Yavhqf
GKCKeC3tBZrNk5BsZdzP64ki8tNlkj456f3OOO2F+BOp0XSS8MjgM7Y1+nzs6h8eEm9m2l5K0U4A
61k0run9vQnfa+n+Np24ks1P/9awaSMJVe6Jo0jqF30+BvCsvssYDF+jpqrCHG5wpj95vB8k2H8V
IOn9sD/GUVd5ZE0+Fr6BTXbh90SKMnHQl9b9UO4zSDzw58OYzg0HoopSdE0BfhdfofSfGgOPFtjB
LaGGbAcv+nBWz3eKC3nNGtGiZh9h7N/LlB/2GOf/RsBO389GICRJITXcaesuw/vmA0rSkJqsksdM
WKnzQTSV4ay96T7c4fe+LaYwyfwlR/+sJQApNeWViRnf6I0xtK9l7/GAMm7oqcvh0b+YKIaQAXlk
QHOrQ7MezTc4b96AcoMmVKH/Df1t8lu59Vh4TOQckHiUVeGqEVE9UyB+qsW6aqDEL8k0QGy7+9aR
G1DqLCh+fBceEm1ONPdEUjbksb7a0bxFAqQoFk/AjDGUCone+LapEW0ZzkXZRZurrddeFtDI8ju/
C4AvBV90rc4LWPsqJFc8GoTbAhayaXa0wSQ2iteDrpSm2wOc5bsDEGKr2i3hyfyRScPD528fo1UQ
M3odU1USQD1ENdcWKYjdt5JmnyHZR29ZLAFU4CqUFT0QOg/ioWS1Cjz7B/RfDd11VON6svzFhFRI
Cs/EjTO+A1AgB53vROjusj4OkPqe83X2z9OTAOw5z7E5Av3PE5Ubcx02pRcrbmyAzE2PVrdAuw+C
XP7yDjfZTTorZ4R7WMHiN6apzwib5QWgd8ZVxPJigj8Ou0I9zt48sPwhD6OlBEzToQlAA3TQu1Ol
qOek7r1N4nGdUx7rkcG6BclmgFkd3mR9sBPOr884cd2Tz0FRbd/lkuDpqkaN7AVNVm01DXP5boRc
37Sdjm2JYAFZAgl1Hkr0I7AalOF8vXWJzrXW9EAnUwxgMDREJtgt8lWV2KER4WBcw1LNkDR2MURn
A/V4Q1HYWoDcIyUwGW4YtJAV1IjtZWfc1rImwqY6J+X0+Ve7/SU9Pw6hbI5/DV0LixO5Uja8XkDZ
cE9rzAQA6X+38pAvxbH6R8cetTCXzZnEtKauuN4eOqWrnEfmWJ4PA0xpVSZJbDgineSH6TH07c2n
6j3ZYf/dlV6kcxz2xxcqeSzjEy+tMX1WDkVUWCzy8RTbYCL93ZVuPUZKqITvwYUM81Jer5Y5VyZa
g7MXI1Tar/yk23kpt2w5z2q83wwlFL8ppIa2eSQMLgUA4MMvgW4FFW1RyT1BoY8OP36YhLTJGycL
+fQyCiYP00uZAJF03MPm8SPO+JXQIEiAbuWG+yYfbS7vLzbbywXC+71cuRmnycXv6cXgfCvlLPO8
l8UyUmZjtgre599TZEFDitiT5m/SZq1+VuaoAHYuZRtU7f1g7dFgHX9ihRNK/Ost9446RfbIrn4K
Bp/KAKq2Ao0M3l4rACC+wNPOaPZlCShqrHcdKfNyZKTCPWYor2dDHqL8RmJy/wxqnEpkGuYhlP00
6YPUqVH4vHBEMzhzx05BzXtCHzIF/hKMoE2xMKHhQGt5uTzeuEeKGVqmJhRLk1JUVJVJRR/F0niI
HQ/9l/Bkweh+04XAaOF0HrR+KGbDeZQnEySbaM/HLMu4NSwiTPMFR9VbnXfFiXuwP+n9oM5uBW0Y
UpWDDGGb+sxp897EPxX251MKklClK2KwEtIAZu4MpaBgbhqJSlGdH/TbKm3rmN2b5eyPzHMMTc4S
IBuU8wcMshvpII1TaENPYgzaMp9VD+6atUKOf5zVTt3UNzUvOmgWPShpEz1owCku6ls5Et5LEZVw
8ZeA5x6c19Vw8hdOyduFO5m9g7hP+MfgeI6Ox1BN2ywMH+xMGTxaDj+7PL67+T6KzcStICrxyggB
WKDXDWC9h2vgkk4Nzcn7SKFLbsKSXKPXz/W1635QAw3Z9gqMq8pGYYsJgV8pq1MMCO1bjMcsuUBn
OUXRdVG0u3265k254sNoy0OPEiOwDjmZQhT6khgv0T5GU21eBN5a0OafMbDIA45LlWvMImsPoKa+
BIWguoJni2deE2Tjr6Q6clHmOuOa4sl89qSHgRlsyaEDWK8fhZaQUONpskFJ76mk2X50QUE953T2
8S5IwVExoPiXv0OiYSPTZWV7goXuIuhC1fYxX7vOJDs0Vz1CMGUksEgE3zGnC0WJs1RRv0fbuXNL
w2mwBgp0jCejssqlGzq5iYhbzMoINEc4VqHAnglITaRW912b702/1GaSHhdgr8rPUEXwPlRGA8o/
UxTHdIwOnhVNWBLkQbVNA5vJvbMXMeivOguLYKa+NBisjaO6Y9xWAZkzflpM5qapgQpk6DnQTk2X
73QAPDDzXE7YrpSC6Ukw/mOLp2YwzUCBWtFZZW3eZOW9sCq4cdD1GNM/KVVufTfJ9AFU7LYnBHea
sCY6C+3YOSQvDDvIPjA6Cx48lh6QyHPSftiBo8VoxNSEYpMjL82fn2XaQ51n3/rutcl5Ki9PEjyo
KEQSA7U4ZXmA1nAB7+gkHLIgFcuvMKpt2Mjdo2/5BtSL0FI45dw4xPfPO7s2Fi7KxF9Cnkt6stc5
c0/k0fvbHqi0zazejF5uVLR7nyfmspZ3hq2PAN1/OJm/VJC5GyWxVBEmFagQ72MrsKQzI/LW28aS
mj0tmn3/aQPxDjZcjULFAmdviyQNy0upGiT+aocJaWVC2AeUHpci/xHOB0LA1AwKVTbAAG+8Jyud
xi9X3VJYiUdW7i2sguJa/epizalH3qBOYCSfmeWBGtlthv8FjyhHp03S7ew2ZZ0rt3AH91sNuhWg
2waNypz7NzMxUz6e/ZZhCcfIt8HyM+U+LP/sl5eeEZ4/K8urskimdb15MwGa8Pov/eEvAJXHRqqK
nAHUW/76f8aGoRR/FphY/Rz0GrHbyl0f1DrQeA4WfDFh+IxxT6c5M8yo6IqxRz9smHI4o1vMqdWO
35sv6iIvJU1w+SRU1icMz4BmJJLfAXZQ1vfwk89wxer75gzC4gklCw/ObjX0yJBWdluVmeAP2LOY
x5S2+Fhf/J96JqUIlUSFhTu6LmLEbWBTuPmUPwsxCP720Rr7kQp2lfOR+2QK2iQQZYwdJRw5nXOD
UYd4mwZJlbyiXnZ9OE8FTlyNUqjIqf0DK7P//5lOJ6zTUGmiEJCMgbI4mYveACEf8IdxM4DIDVRG
HbO+V7PGS+/9c7co6VtyKC5bTCqX7Go2P4zcILVsB5zXBTJxzjcbXSeLMIrGkWQNY4r1x1e1xQUU
adAJx6+hBBKIujEm6eeyjt2dV5y2+dUBwHpNp2Q/ZW7lftCt824oTnw2JvnOUzZvfSKlju+5qvLt
n9wS2hxpEuJMcAAFfm6CEHyXSNws4UtpRjN/qO8Ej5IOMytNP8H1/4OKbFE0l7ghU0kGMAJzqUdN
5nXTmA5faNC/QP9EcD2aNcXASz7f9C3Mnljnh1afVEVUDXcI1w5Cq6oJeqhjakXS7bdoJhKBQZVQ
aUwgTESteNV5zrNog45D9EFq8WGQZlrWPg/EDMPQZgQpTEh/rlYmYBtkuzub8gTBbbe7lXpRlRlT
cI7N2PwJGGorRrPZhty9E7ooEeWsu4Uyznh5vS/PbQ1V7PWL7Zj56PXbwhQjO6R5NhMeJ1/PAJsu
85Lx0dWY/aNnlrnmnwHZRFDmtdCtrS3rgpi058mRCsPuHlw6JeN8+STETxYwxEq1T8JFF1gSaiEN
gtb3YNzy43yX3aDP2ejRf2Xo+LsSGfZP/3UYz/hvobF2AeFn0yTvbOXPBR2OA7Z6up/Jl2ZSRc1t
7ME0Y24l/7N8YkqEwSWMX4f7xhqJ/VZ0xEzPoTUhDLQ0/RBpnjW0fRl0jfd8uBcfwFDCpacDsyKB
jXIxProvFO2KqEpmFC37I/lQCs6dAfXoBhZfhIeINbJTd6F7gOKMjc+7Zn/MMFSiUMbnawwr6fmO
x+wV6VUH8BX749kV1oKiPUFB53ToXnitIvx6onLctr81COwC07wrSIuW2enIKCm9cTu+o6TmRo2k
9gfWR9ZGq2ejUwKjWCOxnQruWQ4Pbr66IhJnkxjdnTJJ0mUqoegdc2aAo2WIPkO9d+Rh5NzrJlkI
pcARehbO61hPRASTN31nZpJGmISHPevW354Kh9NGsBAPP3m9hK/r18QFsCqCH4X+bHo1RKSJIGpu
yiQdz1AK/xWVpbcQUIp/S4Wk1+N0MqebNPrPWW46ac6pwgchpEv7Exiy+BwLdGnPoAnMvsrMxrem
tbGDP/VpqXFxoVxEqpQANoU/wMm6T8kPRbz6qF9+h3PP9FLtjBAqLIEwcBDZj1YehDJiJUh9ncQ7
Yu7T4IsvAxOkcyzj00MNGSl1+jJTP+qUtHid/pmMK+AAsXfQxfWT12Jn5EIFr251xy0Ks3Z/W0jr
jVIIHXUIXoLT/vzdWReGfwig3UJr4IXfTiwNbKjdMbRGkEG56WHjUmsamlrrci+37sJ6FGnxm7Im
MtHclFBwLpZ4gbys59gupaTZCafhDNhrzVfWXiVZxd0gZ8ngXzsjHpNHijd4lLFFGj3WUlAks59e
0OP9fpPzx8YTZhX+u6q5edcHwrohLzdYgHGrlixf8MeLy+RkAHYK2ECD/EHSiXHFw8t40WUuAgff
Q9UzH6Qh/6iz0w5pXYJI5KGwdVG+520r89PM9A29wf+fR+zVKwLZ6FojtphanzsQK6CtAJWypUzv
1yez06hGjm1ntfIIFAPFepUGil0xy+gvzAnpok119SqHQ4Huvt9DJYsaCA1SH2f8jysI3aesj4MG
H7W6mmysF4wEKWqygDEp/A1HttmeQjR4HGykLNp1lhJgt1/c8tXscf9RBGDYn3kji360DEkhzIy4
0R3KftM1Gj10KeN69KB72GMSRJrf+p8tOK34ggWEkSRqB1eMjQi+Fs/LLBruFZBVKH/vDTmMhoWk
miz5ngYEOMsPANIg1uu3X3m3cEVS5vikN/k/AUdMgHfCz3BvPQK0X746Vovkv2SL47GciH2RjsxR
vdA+ViF3yzLXf+ZQHgq7+/zuWIfJ1oIE4b3lX1FaLc1/8ubwGJ80xNH1IEfy6Fl1xB6tNSCx6Gx2
VEM0OUNYoyu8DEhuaxMTj+bey0ZEo8udYHYTyD7xAklTbe1G2Nn94qNU3TMJzqVzB3f08n799nkY
Jh8QYyTdm3N4KPqUECruXBAA+T8vUGeLa8NGAJl1FzFNdO2EpRS8OVBvXTYaxakwoybKINEEe1al
Ef90+uhvLjWFeymfgfUx9RlGZDlh5qThSUimRutHyuBN1EXvdhF5JWlqYDVzJRRLbybWpUDNiFnR
Jz3Snyq+JCKwrexPudepFk0GY7cbH2QrTtOlB/TVW6oA00UIImW/E0vzV6jYG4l17AtyQ08CyYPx
3QD+HjUYlFkPXmUJvEzOjhxoQTV+5ZbM/egvjvGQlMVl/X6IhuwDyt8qtutym3dtrXBZiruAnkJi
IzfvqkHmNOX423lqXRmzs7YNb9p4/MH4QZQ6rEcDFOLLJCDJZlyEGhA69rxQ3DZHpoCFu6EIyi0P
+0lUUYk0T5pyF+RQdNb2nYxF8rOb/NUL0CCjeqte3Pq5PAmSaIUJduGa+lKy7seZPUuy2WL6w40t
Zd+mdFyM0hajuKhFePkZ5g7nXIVDgegnGxAKOXNmHvFFb/PomLPxDyPPkUIe3Rl4CnNk0H7Nsa+s
QkEL+qCkmunr1De7IuNxzKG+9Sjf7iTobJJiaEduA4tfPlfjGF7zJOFyNmxU4AubI07qIp7s8bGp
VWkY+uOlNd9iMdoFXxCqUxQqt9aS8ND17P+Wysm1iTb/j64TrthvwtaHZ0SqVZHGd4i3Pm1GW267
fVNtVbHdW1299jAA4tT2fgz7vUarogIk1CBtk+XY189XtVraYtNIWfu4XxbSffwSUW1iUcNaCTjh
p+uW4l5vmQPO2E0ww3JXM8n/BpL7gqvj75vDTjG3PbUjyh1uymID7ePk9PL70i2J73pPZSfIkw62
exUYIpYZh86lP9ZkaJkfKlfo+AmD3b01UHK7PQ3kx4BBSuBxfnPTWDCYBf5lNWgJSx55/jH9zGB8
uWDpWhS8QBkk2bdeNwMvJzhnayox0xehvaYQhNywEFmY8084Olylk6dTpKpCuHVlWQ6rBTG0sdHH
KypfUqYX2LS0B0rNOaK7O2YGhMiJEvLp+J5MjUpv5zD0kGmYvNJEbeqakfeksn+kKBCqijaDrvcx
ecIyW62Z1taTN7U48xwU+aSeYCgNjMOkFafemudmRyHcY0G03kC6u+/89ZdTtcykPrmvw1RmBTew
tZVMnqODoxch9HiP7a94oqXQB5VTvLvZ1XKnfOAwsYCZ88ltHUOQ0PUFj9IteNQywWriov20TM4L
prdRV+Z0rtWxJLg4+8X6uOtjz81rcFNOBP0MoVcxd+jnKA97gihKs17Vsv5uv7I7iexCGU/f4ywH
yw09bmd1x9+BfRpH4fZWeBcx6Ak1do9CzEWkmHFrTcESDQUx7EcQ6vdgV4D2uhfrhngPP3Gm4tEa
sCaX4hNt8xJ56RqGIHLgq4oZI6Qf2bSTgQTtTODFXTu0Lm/0jBksn1qb5kKq3D3uGQ0AeZA0UyY8
+YowxHhgnyF8x1hrkDDObF6vG2exklVpvepi1QDtMZTmA7Hmhxgg9Fn8dn/r2XfQFMpRiXY5we7V
u9IKaytDIat5wj/r2740RusRSdS2sAq3DDNBlxbdCqZottlgKJ0FITePaOwpBNBxG4/LM5B85CjE
ZMVDcX9TIBxEYGgiLp/aOhchMgscHiaBgYlB96/56K54Ejwfhms9TnCfm57XCg8/PzDG2szsLRx2
M5LPHPjoFTXpZyOar5Gb7q53MyLmOTaMynQ49mZA/S+JzIbR8LwHLUw3R4wsvUn78fZnBbYkpHW3
/fqoc40cmO/9G5Jx6X0WMAWPNnSUSqmhofgyiyOfogjLCg6KOnyx0cTa2AbFS2J8/U6liim+ToA6
vofkxim/x2Z1kwokxc3YmzRJf+par93vS2N0gIvMUZhY6MrNiyWDPy3eVqyCqQPNmIHUaidBBMhV
2vXv2QH2zUdXY4+0OXTpS8tZrtlTwP4bMgyujSJQFaVbdWITlwCdI1wOQ+PRS2iBYG4mYnGiaSYh
5cTpAkaTIrn2VPTLU/EjLgEvXxeMo1G7StKvcyC0a6BM/2t/+hqMC5FtGRrPpfmvbwPOhEX6EdQv
YUu0c7ld/PAysfWCsre8d3WT7qvNQtd0pvbj9Z/l+5BTcvBmbTBCwlwPsadxQueyg7AG5qQ31bUF
91ANImlF1kR3mBR0UcSn+LNNTcd43F28Q2M2dzJQdMTvPFtmxRaqzPXvO2yD7Zw1O8S+bxKMQq+n
QHK3MvkZ+NwoXO0mZSjHZJbCikDKpguV9f4DmlbsCQZb28u/IO+Z4NOx1Bda+LGRap4ciI6r8sVe
M3+Ml4+p//5AoUXjv4wlUMuQQh5F3zgOuZH0OceCHNnq1JDdbwiC13RK2D0NaxkcdSNRgYkPBgvR
Ai7B5+Cx9yOCyrS1dI37wtuKndnPco1YjZXts0rNvUKH63JsTH30quU97k+Qx5uJyd5G39x+U00W
yn8b2V/sWDxq71dr8QYDHICyhND3VsOyutJO/elKEwUf62HA1Q7EB8KGC2fszThH9HAwOcOckg0R
yBAbEVqUMo4SxQ9Nrq/j9ufHFdsVyODFH6fyFDWGOXDs8XqIkGVUN0D9vFptjrVOPP9IR3VDFL1C
uIx+R/yqGZg9ms3LO43qlkLM6MZZscpXigrs4X5t9/0zFiatnLcQEmXluiPZwOaTxzXn1ykYNJwt
hLURiQddkDWXPeRXHJoGjPaFtZNK1D189aAQAhWg6Jo9AuvImQkBK5PSm4UZzC5xd80uKWUGPloF
Nc9wQAV3CwhnsY3yUkaEHwFAbvhuTSO0L72Lu/9rzohSlxStgCKAedWUv5wC+cAW40jbIW2KXq+i
TGHeDXSucMGqZAyUA/4Fhs1+JjzUEgpiDx3BpFCWpayqtavVeicsAFpQIhq0AsqSqshPT0Lnzksl
0XmBslEIH7zv6njbrBa+SjVcTOTkSrbGs0WZmxoXFWNzRa3Vt3tQEpvko+GKV5znWcu8NMjpU/sh
SRK6JRH6rN/0C5HtKi7Q5XktdYpdI1brAnNSWkhAraZ/ZDBM9ZZAWPZx7HLbM2YPvChh2BpjW5zN
z18FVYiKfV44WeSRRJ+6dtEsmeHCcgv8++PIbZ/Apa3509rKJRWFSsR3Cr27wOYt4YGblyuOd70N
dZY6UTiH2jI2qAMsgm+J8xtJ8jGh2RV3VCY5zXh/BkS39HJAorR9MomuJN28VPKV5in8L628/Bgn
ynSEv6C2/DNUt36ddWWGM6TE2HiLKSc/vi3GaR2isJWQhWNbRnw4FdLMesHCNguz+qYAtuq1vz1u
rT7I1VHQ9+37Z8PLXZb5X+Cixvto13IwaycuATY17+awtNrAicQxUcyPH9oI1YCCxC7qnCkuw0/J
AQz8yGWIWMmNsjb9Rsz/J6QwaYOSzXo6F5plw6LVQu5pOkRZEbYJZmacsaOZ6H+iXVqJq+HiSRzL
nLjqisDFm/Qy1P/EjkPwHJ7dZoua5rt6M1lH8zh5EiLhcHycWGO6bMmunltZYEpa8cqe9Gcs6cKL
SrfXCtcoXCdXrJI5HMOKjNFEOxUkVswgbMw0BOf76bl8fNEIo8f5QlxE6TSWUboiXFcKKXbW1t0x
1KBdvcNoj47nEK9eb02AyzIHZep0cxaLyHAgWB6tYGDBSwiC4bMlkddL1tNAq4o/ydv+M1YzhEU1
Mamc7YuD8U4C9bNwW/IRtg3e8JLlvl/TyO1P4ReW+EwHLxnn4As3l7pbpbxzldCC4ACcHFXa5CXg
3gmPPaWg51KTbpgEVjXsGWEJPqztAGQvoM+4DoOdmi0Km5QS6QniKSvkGwoHyDVEhpIw4BxKElmi
nTcGq7JwQWdbAlyuQHtj2rq6LHea3YwF2pgpYMOWEhbaUcHxoFkVhEgLH3LFx8T6s7t/yKJ7hap3
7KzKAw6spxUKzOR9sEsif5ohjpPnMfv9a+X7PPR6Y9oVE+ovxMkoqOXb7w1ZBJAZ7jn9g2biLU7M
4rFK5JhavTsd6Ky8eRo5lrOJrM+Pko9mTuMj/fgfDVpVNUTklhT8tLIyUkhXlwM/VDeRzrAn1a0u
n5NqM8BlEOqkpzuH2nt4BfQWs7T+G/MJjSHu6PZflTl2NUFxrIlFY/EZI36X74K5q879SkTLL1XY
bGUxa0i0kXJAvFLlNigWP4tLoK374XOik2rna0mEAZEvgAZZVQARMdDzrmeVmwM6n3mUmcKG4nSs
Ei/IfNfui9Wo/L0J9xNB1vFnp2RD19b9IfyRn7h7lWNCU3rptPs/0JV1+joYWN/cBHgXcCCZS4FI
C0b2Ew/2GrnOJ4fSqwa9AOYogseNKstbGIUqhLQd7/UzICRbXabYinCe2R3qbXw1lGFJc5FCf/7z
B8OOW4/T4tBsn5MNFLUEuPKW8XIP4aILHKOYwbIx86mg3WuIZjuirsj4StKb1LM1V6aBh5Jl7J3j
Mrj0zY8v6FIhshKfAjh9d9VA++WiApYaxo7Oib4Mt6JvRv9FYxEEClF5pZDlVxAEoAmF1i/t/N9P
b2vV6kmtp5Pm/kEIAKEoFauJ5qEnk2P3K+LqX6Wn65bWRRJjUUgE3JjY2tN/Upu6LdNCBU9Uee4U
uK9uXNmtejE85r1e2Q8YU5/TsI2t390iqhsS5UXWCPnZ8WpVdHTJ7rDZz8vhqryz2Ut5WBhaQKPd
EmzGQiy9sZ47bSSBCBHpkaPWPtrfwIpZTmA81I9xrTF24033Tc5W0lnkxtDxmtq6apuf7mlvFFbI
+t4FoRGKDubPpLigA7e783otZdK6TfN0VxIZIpcj5SI5PxktxolKDQLVipH5Ga60nFJR5UqHAvk3
9HS+NofUnx18Khd4BMa+slB5OtTKEtuJwhCdxbCIprVazAUhB76V3TkGXnc7b9Q67SDLdmjibCme
U0BU3TCz46U4ymE8L9q7ENutBJFxJ5XuqkAnwM3jchRcxF4EsUdeu9HwPuqgk8CuG1YOkKxEOTvu
4BEKJnKDJDQGhnD+qtKFgMa8f6cJJj4M5ioHPSByPfKKajSIzlOon+2XU5VXKX0dScXHD/d5LkGz
2Xpa/NTIfljXmQrwbtvfsMSYWyvMfyG1Pg1SC9tVSUSyGs8yZkigJ9ivDfgoNErnslbZ75bp0J9o
i3e/GfQIEJw0INf8pIdz+opKlOq7DcKwNza/rfImjhahJ3PYZwctuXWS/wXJig+IhvVmN1y3boX+
3qm+74QNL+ktuwsp+SUGOxA7j4GhbbxLTLfqsdRRIihFgc0fveWmssfLIeGnAwRtduY0UtKUZo7I
5coRxJXDOy/HGiGAXK6T245uRVeJuHcagGPnuF+dx+zJ4UeQCsnEln6jtDIaOdngBwLxCZLeWhel
PeNvRifE2/me5uKi3J/cdw41qGGu/sNzCULRJOrWRyPhh7U/C8RV/5i/72O9+ywV6g9hCiWJWtKB
3jB5QzbqU6fO6MJDhEZWEKrqTli6RMu9bncaBV12pdU8Z48F0T0SBfOEDlrr7Bqt75Ol86xjwE8J
eH0p2lmoNjdCBC3sEWF3Osi3I/ZLr+rCQ8+MtySk11UjGf2u3j4ePFg0VjJXt1NK/0/6wKdLEPMS
6SOiFX4/FBAQ9NqixazHTMAsXjBdSS4bg8HHcAZ32ju3BBKfXuPgPzD9zXjUuIcqAiD4z89tBN2M
SxVE4NRD/FUe4YctZhQI+zXutWkBkPV9x84pHzmtidKpnVD40QMYzJIBfSe3gACieumnPkc3ClKm
TgRM0j5zzdfnoM0VyyPxqXmIjHVKg6htfsOBYacal+iv8WrtaINML7pmwXzwcDJAIabzyUDfEJbp
4XM0LSPwsbQbpJirA2ogT+y/tpiVmjyT2Vq1qJNasiMa7UzqMpzzrcrsJb1TbMKXIFQpNta11YPq
3gUVJZU3bA5Pl931f7QJzNnS1B2e0j6DAEIMocfaneU6zyRIUAmPeouMJ5SuaV/VVSzzBnZ8Br6b
kok57GgU1RpmrnEyCn5bXAfW90w9UHt55pTv170qjSJYGBn5FjGHnFEEAxLCvSgnvSJXM2rfAiOm
UVY2TeTbfOW1pYZtu4joG55U9ChEGS2r6hh71v3Wc/yqXUGEzPOzQdLSbxqtaIRcNbfPC+sAY3IK
wQ5DECiFykbMnN3b/fpdm6aJ8baWSb0UawW/yDkDA3Mr/C6zTxGN2tqtqXtrO6zZCpSXGb1Mp/CD
AHVDutQHlDCEwlb6IfyYAZOdVIdffS850mwbJ2raEIeH0RBRO2CaZi1k9vUFQg+kYy42sJEY3ZIP
aemYa/9PNoiWdoqJ+Cl+9FwNCls/oBFybNrCLshRZsanWSinBddwxjXoBOfHtVB6m1tVUXqEbbWt
lcVVML7QB8aVts8F4L+eLTLwTGsqk/bk6sPoTDZdjwn1tDKwqu0miCxYJ+Fef59KtINUyN8Wq90C
XsrzTktpW7XcJMWYS8mJRiDC4nDrmx3tCK1qKOAXOJjKh3m2uuiPnDJbHECmlr+WqsGY2kDny4hH
Eva8iWpCk1sH7yiBypwMnW5RnAiWUOVeDMyYlnvbkHwZEEHQ8ZDyBQAD/CSvG6V6u+BSV7GpEcfB
tb7i+IQ/a4EjCWJVb4pUjD3BSNo+lgt4jdx2gd5LV7msdwqrJNISzGHBnOOo5JfypK0R6DM7489/
m7UizDqbSY9Ek9mwlI0lSesyVqvTCqBnNRTOUQOCtA/DNyHkSkY8vzNOdkA+nI0RH9PBTBXBcfq/
PAraqfqbJT6pGcPgEVlsSxN/qtLcJ+zpWKE/XA4gy9QmxhIJkeH9X4b87pVVm5bRZklBe5ma46H8
pRpBv7EQz9wNQ42afklMymdguDKVwRP2LQh3Y7W5GN7vVZd7DjYFVXd1DlV4Gg4S/W+454WPOoVe
1BElasqLZcvUO2MoYCVikhwxU92lWBh1Z4Xn+r4MFI3FXltn8UIJyoF1UxA96aYxKCnQr9fJxlqS
MW9I/Fv0LleXJqnOarVDk5t0k5cX2PLlbs+2HCHYTdR7nEgGYmHvOtn8kp+n7dDBMAT1Cn9yXdcq
+0AQtfGnP/qSto4J6+aKaI5pzJBoYD0HUdmxnOyWj++XKasg00fQ5tjQvq7vV4kl6dESN1zSp+j8
CEV2KOXU22Ubmg9ylMdZW6Ku5pQ1fQCT2GD9X9GRinUy78bdZJRzyhbqtPWk064V/V/GAuj7hmwR
e1usFxPukEFUNGe2JaT4G+D7fzUkztE8d2YG1TfeJiHjMoQceEV4r5gkChUiyjwt3yC2/rQVZqhT
IvHo1NcdqbKjLRgIvbZxfF12UAY8OqUoQia1OGmNuYgx2qEX3M5MwcedIdWZO5HwoVXsjcaH1RsL
Ueum1+FtfH9t0Pdc5xSu9nBMkYsgAlvBdrHHpmhj0YONQEK7VOSRGVX1Dg4LdbsFHCvWJ4S/DHnK
zzkWf5FuOC+vOujP2i65LvwTagh5h2L6dOvq6Q0beKY1I4SnybmYUJP1fLsQPZFPWwrabBY7qhaM
sGCgXNrU5D23YmH/9ajF6w4atGHodGl8jAkQVWkoW0r313MgyZ9eDGdmFixeA0ivTNPTtDa/g8fS
WbSN7SFa1+2IiG2jvNo2gPVIhAj/QEmNWYwTnBo+Rz8JdpPuRSy7jZIXWbdmNNwy/GuvMNzPjLvH
Iz5KxHtKsOcZ8/bp0zFIwtb1JwIwHX3SbMR98srRARxjwXms6eOZprQVhFQi8CQchvWNId9V1weF
jGQYuoAWHxI1YzWzUqUlfZMDsF78icFdVgCdhICeZu9l+4WzTPPGivrUPqeZT8HRbuwPtsxs6Mdg
sG9Eqx2yCq7PfpaQDn2Zcw3viIamUUFE9+HqBAHkBKZDGFKwosrK0FNBuKU+HYH5wvjUW1D0WgiO
ZKdj/4oBZ3CZE4zKfDE4GeI36qgURO0wE7Rmqthw5fFp8Zxle9F6++IFWmwt6HsM21jdORLtvTIb
gNTuerUfJelXXliNAQWlvfG3idSeUeSkdKYV8N6TM3AkeF47S9wtwHrMuQvExMFnDii0FDU982N1
q/o9CDPAHfLDz2pmjeBK45JyaJqRVYI33stHQjcZHfWXN0NSuiLY21pmtEqLffwxlPVEWwUqLSC1
2mnCRQIFeocXVguO8DRPI//A12hZa/CP5qZcnNKLHCoEee3iNcXf+/MqGKYo5Ktfv62ZGQDbnJ2C
Uhv2KbK+Rc2koFKr4EejnSbtiKDZrmcgqUDhLuaJmXN5Ef/nrKN0tYFJIOvFgeD5/t9i/ggj1pS9
IHjTte2mMvSamt+WlTVku5OO5uKdVs1hd3SAkZzw4fr7trNUF2VPbL1dRy/hSgXg83/1i48pPCCu
X4X/viS4UBDQcfgLSk9AteaJ6Ic4oubsDJ9LjjLKN95Gn8S46PRAwdRKfzUkNqKUzfoNMwm8V83W
P+ZlxDgnzcoHdDx91qfrB4m978hxW9a2Td0PS/llD+YS0kmZbYcfx3grg6RU11+rtgmdmPT6ObhC
HNUj/LBk2T17l0SfVyLnb9jP4ltgTAhyldSylkN6J6XuU7kiPKJxTlqzSbssxqeaZf0TVKfD7Qoa
U1tSgsmi/xXAqooJH9Qb8Oet9WcgSaQZrSQ8L2U+M7h8YQ0VhZtpmpjP/y12cFt7FBHOwtpR4l0j
3eomz8zpsNqYvndbkWbc7jVajoFRD6WYCxy416S7Bb0tnUsCYi6JK0ZuXRY3QIc3go4/UEL16UZQ
GR+yq1qAmedCcDRWRhyPbqkZrhwcAbDmvuCyeUiSnIwPS5G/KplCJr/YiHHKxoYcKplQgF03FDru
ZRjNw8sTreWv3mz5KETn0PgnoG6oYV5qHlWGYFRPkXR69UmrAsqOZRuKxuP/bOBvIzOP1WX6tfIb
+GnFg3fXsmZfH6LBJaepc1Qjx6VrtXtFkpu1D1TM/mXy7oFsp2NrVqo3NHrHHSrNPzY1s4NBfJ12
LjbzUQ7rzno3dBUt2hWqL3ZHBtwjtQWRRmR4jwQ/imCgWMxJKO+0pSvlnGEyb5x6KkHe1MuYjWbU
PNXW9rD7ic1RtMiw4QANJEALGyDE/OeUfcPXsgcRnSOwiOdzBUVkOptIY/ep+q9qF6BRYlPw6Ns9
sRMd9xuKIoGsrKHEbS4T/HD5C12rhr6M5QBoPTynw7v0g5WD3e9+5vrB6nDZe0QpwsgkHbVtEEHp
2S2SNByf4uce8x/UeWuskBPGsY4Y+py+haUMRRDA7xZGhm0Bl3ibU2H1pCNjt3OLNb7fO5+ZMrMw
QIAUOd0gmiA8nFUSqEA7Hx56Ic7DzZU9gIYh4eT9AXkEvW1Vb8FZnm0hlq+i+5hjcKbcD7ziqAyX
1d0nKOKA9k3PVgwr5q8BVOBgWUOHx4tAHgKg0hLdad6FisEaGEemYt0ik4CTB+ag9PdqsYU+7iqI
bdtAFTNWgFiosa7gD9thwPqbimvqkbRVP1gW/vLqpuUTRc3ZVlFmRipCNNbDuhtUCbcknqHh3e+p
o7b2j1EgQl2nAIA6vu8bMx2OlBKWYsCpzpZ0qqtGrFXkzdZPmDOfCgy5e9XYTHL+nLOG4ZNBGvCf
WnDr8mftaTj0PgG0fkDN6BHsFxcJFpU6F0m3iUK2Ath1SdgZtMlYO/odeofq9Uwnvz1J0CBTcyCt
pquTFbng9VFPRhkePuiiy7c5GnRi1Bxem50aefok+ohyo9sD5GI5Vy5z4PxgI0T7+7NG67cVi4MK
TiFMsxApmUEehAJvpaUqY5AjXxJiP2BD+kcuFhz0FnUcf80XhQfHz2D9qjJK4HDP/Kjbk5PNK+FU
EGTMI0ukMRXikJgMONMZytYxwOnEDaLE6DSsbMfEE9H0MmaH0fktZcDcAtIMOFc9SEA3OrlKt76s
IUE57e5dFlZ5WsDDtRnXTFcWxmbkU6btJ2MGG8jAhWH92cWHcftgs/kvRbZe5A0llpsUCzGKTOAA
Lx9q6M1zum/9IxHu1uNPmGa1LtgxD/4bJbYmcjJQU/GkHUX1wV1oMA6QR5E+zVo6+aVxyqFunKnf
y1UlrBC8jVV2s62YGaRc1DEoos9JIPBKMCRRS5ZqlFfLZDCYp1x5CdcCzpYO3RlXcQ2irgLmAuq5
G8MGIoFShB0vMeonq56YEkXiftFGb/8qTVHeLpwZSzruf0i9qbyYccsVz1ITxEthetFTGWLEdEyf
gIwZ5MlzFz4kX/L7r0t0hBWZ1XNBa3rGfQPaZQg7wtWg4hnSyRSL0HV1EI3D8zXArXIpAqjAbwLA
f7ElqUVsa1dF2iRakaCHi61599/UaiXZoiPuDF+BvPLd6ZwnCcqW39N8OQ2qVNSLQ5/wETCNdY1O
DBQaRGSIng2doTZr1pnbH5zg21QWGJzmYyACQ4Wct8SrhUmqGpXkUygnGBD3hw3PRcjKpf6E6Gh8
JzYu9aSlF6fsScWJIp/KeEfG44aTiDLyfuwO5iKLrjVPbH05LZGKjXvAvE0e4qeGRIESTov68ivH
nG72fbb5wF+IffRyLSh5y5gUtNsLlslfBrgF61UjfEEoaOeCyM9FyEa/E1zd4nK4ZNpIMSDtymtM
9dlTKOEz9ABUTF5/9WjC7LHqNsF2bl2yRTI4CtDjh7o2AkXQzCu8rjgmjUKwyecXVoCtvqaQUvoB
enDyyPBLeUJ1N6MI4Qua+1tVChQt9/ETEjGbgE36YzafvpNdoxK7kvcP5x8f8pbY+0lHqMrGcyn+
OhFz0/PL1VeGEA0taR/mnhGzn2g+GxoY03xO/7JrF4id//1F6IdkWk1cj4IaF81OOpRaiPGjgDNE
s2py1THj4cCPtosh1dY6zAvUf97wkLJlUjkrIu2SXES5ThuznlNyA4B5YdZYHeMy+sK7eoSIJKoz
9yIHma+mZrjAJjq+nNOr0wAVV/rkg+t1YA9nrBL5+w0oKpNdDlaFBIsh12QjtZS0NYTSOiWHVFAn
yMevSbjqjX8JSeXTI7TKCwE9hyI+SaFQDLJMr6Tvbsxk15Ld++gdBct34YmUvK2dmOXAJNhHvzqV
9w+SkBXmHFD9N5iwAyUyQHj/GEoZDQ6IN7rPoWDtMy16iOIvkrqPwZC10V4bcN1O9RD5C56PaAOb
HAn+6aTyAiep12ovi8rKErTMepfdWD2eWcP9s9cwUpLMhKJ6UeD+E/+8/n8EgpHhCtwIZjuznlv1
gQn5AaPKTq0FRu2ii8DBLIPBupj/oCgm5Q7IUqv7TxYy4ANTE6PYpZR4xNLvUuQZrtIBo9/m1bvq
/1r/xvQ6ShZnDR+NFSwQh3f62l1j5o5R42orfmDWf2CxqZ02qiWDs1X8OFrxEEfbz5E5+dAh1yrC
RDGeWkqTthS+k6DoHgZD3beCHu7e9WiDmgKCtiSrDXnRQrAjojHyiP7zzB16zvv8WnwUy3OPvk0l
+cODLvRw65aYQmnZMvtM8CdK3pYaWXaNdhMIe5X/w4MripWAcomIuZp+bk9h7I/SKsxTUL3Em+SX
txO3HJUhCJWGaL/ObPSQfEryJDrxBKic/OWTY2dkAIQsw1Ga8WEFxMDeqwpccQfdBuB+cq3h/Vxd
Ox+pFpmxiEmXj5urpRvP89g82j3mPFtZhkpi3EAmvWWsWK9pg4RwSGUSvgrwqzy4fxKc5+/W1VLH
S3ZQxEXRrnDnAbYDy51z0RGYnYwiHmNwurLGAjNtGXGbrep8pNIdXduUdl796khEm/X0C5Ov1eWe
+Q6wwyCg6aiCp6oNQ/ae8Y3GOyoC5XU9pSyW6cVOUFPDZ5M74iE+seB35z0Yb7fH+B1aDtAFgGDL
Kf3YcrSngKexOUAcsgJpfhQTlUofeWT5qtOL4F5A5V6QxG9lc57L/LqUwT5P5HDd3E7iUtgCN9b6
g8btc7OeVdVOn+IaLZRE8WTfK6ewbrOUSXHUZ4FdjkrQrMG5pbSY+cXajz2+Dqc9d5pv3iW/D7AE
INXFjf+IVK+rpM4wjHLzx0/l4ISVKaA11/Z5C9ebPQ/iAMNFoi1xavE4JWfGQNpAPUsU8dQqkARH
Wb13SYrlLnlwNQGIILAWVqirOMNtrbdbbFLlDmxXYbo5I+8FOhGuucJrgRn0ZO3/CGpuLTFJmhEW
YiJiCDd9VX8xcf5796IGLIsB/KUOZlEXl3Uc6weGbK3hjk2k7JQhCBP4Csdy9lsVCTPdR99WNKyW
qkrytAUYnfirgLv32eXRrES6/1sdX+tjBB31Uuj4bdXbOQgzaUiDggMFWn/27Sq+T/x3zVJfMU+N
gsUDFVaZPSWi+ucrMcj0R+qFWXw8WBiGx8AWflJpmdvvoTOR1tgulw5lQPJMddV9iKNnsliK1L39
i+bUGHle0jXr1XThdV9U8KSVmIL0VfXtbyKj/7+Lqwh2aIKpSWB35y74j/3aF/MiFVNSqGcnkdOV
y+hIKAXm2rLxUHsfJLmkiNZeAX8uw21g/MCtlRU/YkRe7k5ppBb2wRKrXQaWtyFAiSsnphJSCp9c
MZiM27+wTM9A2J6wj5lK8+vkkJWyWKNea9pFISuYWyyt+cSy/RLBuWlAaD5gOZ1R/O6kEb4iEvt+
fP3aNcpPHUqAm2jQhWUhsDhns66ECWFYZ+w4KnhjliApfORrmaU6kdBH8jFJ0CBw2kwaCClEXKwh
BlGpLINLkkzKIGtAgFhz/Uczucfl2qJiiKrjINmh5EwHnAZzzHqb5cry7O3WjOCiv9H3oc3RLHca
ry8EDxzXD49U0Lm03EfZtcZTexfoltPjkY/8PazuPvmL9zUgECjjyuzOIDOfrGeNiYleGhkw5vMU
NwUW+8yHOrVEvCHJMjsf8EJoG6T52s70aM8q2PQvxU2hY/FXVp4JA/uM5wbodIDCA9h5LObeWU9p
N4SXJARM/m5OT+Pi+Y2Pe2QS0/xJCr4Y4xGLM2m4gArAu0PQuGmfIPjBaEhgnm4viXYvIda8XhRd
w7N09BcjOjBW//mUCuLv+b9b5/q+RBGmpoXKOQsxYBuc6XYDyt3GQ+9JKA/5FoL2jJ2XH3iYg/IR
ikizoS++78iaa2FqCdLrV7IcI9C7BDqbZsllFZ4d6wG0jNFXoO2K4vICDnEJT40hwlxtspUYKk/+
ED/dWQ5Q38+zdBJzDuh6s2+9+jbYdKkopHNfWs8qKBEgrJsxrM6c6T9/C1EMr2sGyQQk9TbYZW+x
4U9S8w9KsrA3qC7gb1sFYK0Cv9OxWsVI7uvzILo11sKWi3PbMUSKZmx6rvAPa4sNMTGkCCThOyVh
Wk+l/Uhz5mJGLIPqVacQom79rHTYdMi3rzoTnr//IPYujfGp4ni9cQjeozqrPWQU3rJ6Hu9Iycmi
eX3LJtB1TV/uz6gl8kjipdLQVjHTgnvx6WVHKg5lfNUFJclap3T++90FnDwTsSzHq+mo3J4pNNKj
MKI4B0CAUGvqYfSRTQhyMmqx3/NGh/ph9wD7bhoLjnQqlUbeyuK2UPwAtBI6UxtRR29XrNPUEZIG
UeEZ0NydX9pfXm2DVf9w6i1RQ1XtvOSDJtP5Gcvz7CabyL+6QSyoGKBRLvv7718rTAibQasahzSa
OM9uZrEvpn9pjULjeeEs99j7VklAx9tCpCLTk2CaWU+HC+0hYGqr9Zr1rE9+8D5GHHwitaTPyXoq
mg29H7DCaRANmmdn5rX9xyeb/UY++a0oYDnOL+vP3kV9pLkr74KVFQjrrx+Sjb8k+bWfvlPyrp2U
kPfNFzD/cLbSrlhl5sQLalewcuJTW5LYDQncU6HK3jdlpAKCQph96sUGdLGqTfTNItPNJJ5WD/tw
SFVXZTZLEorl0CpBbDTKNW8Vwd4ZpcMDcHuUQj7Eci2qnI04Ull7RTr6Pjav/ldCJJBE2zgXdwAg
yHimiohYulAKcDezrxtqRRQ/bbeyqwj8BqL9RN3iXWxWv/L5K0uTS9C7zdrCTvTKSahbxp3lspu/
FvU7EUT77et8un/5jpVdEqT4yS/mz2GGjrJAQP0dR7m9Qgx0tGeI4C6zacrHbf0UzAjWDGYhkp6j
3HwgcknIS3TU3v0xVqdM18Sq74NZrNwrRwDSAmT1rm34FBRrqIeW4pPcGs5kLGvjBgLuq814RF+H
CpOJCrArR+hXrOS1FpkeVeL6pgBf9Ij9dpEKdNuXaa4r1a190ag2VT2BHIrggpb3SiQiEWKMXV5q
y7KnVMcM4VxKXF5GDWEdc+39V7i3xSzQlC8C2x+QRZ3XMs7YXHBKHLsxhcAg4Jk5hNLBtlv1Zv3J
ozML08ciRXn1HWwCnG/QPdMXvqIuDMa7hAZZvXrXM5LzHxUTlTJaGQCZG6Qh5qlF2aP1l8X2nUCg
P2sPM1+WxKekto2kWmBIWrujojWxG8KhQnIvzTeIPLCYG1i85nJlU6F+29khNNko36jJ6UXdgYiG
ZjYNbrihuWv/kvm6i8SmpT5inlS9YlmKZKbuNR7/NvWRF3qke4Y7b9MeOTlvWj+zRt/YOaSWZlno
hAUEi5HE8EhObxU4vroS/3YzmlkV6Oq9vEcWtXcmJ82BoPrqdeYC76l7QO7NSRkBLTCTZDz4BeCN
+hML0NLCuLVp3pUKs53o3FABey0b4lQs72OUhp/uVaOqCZpS6Vb+X8TBkL9TxNfEvXoZ9NdXBbbp
VwxneHNLvN92kaq+fkt+hjNgJQjYL+cUQXdrFhq5WBCijIjwl9X2PytQI8vKTsoMjVVXFl0ZK4Iw
zN86YdL5OB4m/UySKNAYmGLBpiFftFGTCAhc7dMpwQ3HgzVCPKpFHh5eLUe7zktsouNsF6O0fD8b
IPKD0hznZsEAGamowN9jzU0s3a/naqAKGeizMO6zTfcd6HypMKH6cBRPm11attltHlGPJ3WM+pT0
yFbYMwGjdk0Sn4UDbxuRN6NU4xSt2vogZt0fDacs4qRGIEVMElak6mL1kTrz6PwLNIgq+jQnGFiN
UuepJ09u9V1fLr5sbcOIHzDCW4royK2eU957yeeGPlQoMK0aEB3Qk8UAHKlCgcO/ch6t21Gf43st
nJ2HvBJtoaPYHwbaeZoBrFG0r5OPoIaq4o3UqggLoRfYYOobsHojN+2w5YwStPL6CD7rmue6fnug
E43SYDnkt2zkK80AnDzM68MVNOsaDvU4F7HNwZdDM7+d5i8WU4BRqaN66HlEvCnXBmr6VlZEdoU+
ixkdrFToUhgctjrjRnBMy9ww4KKSdVEc2YgO7r7/cJImeu0Nwa//rYFEeZIjAjc9D8XqBh+rUB5t
Z3fOE14BWXXNMFtJgVWNRbgmFJu94jlshJmDUBnGvAycFNulHXQkGe5QfZg+fbFBIgktppy29QEe
+OH8M92tqLZzDvYe+faZQg7kWQVJSjZ7+sHATY58SoV4KzaB2We8WWTvpjwNSYdG8E6+SPhEvEuv
EnhQxWXfRNGoA7WCNU8QIaDZ9cA3JTwB6YhG5bBUc9MICrUE1ekZ4lfQ7QAoopRHzN9QEbpfKb3H
wgbhFCgClO7nI0iDnRgur+Gpx4Kl0pnelrQQz5q6hBbx8wAhE9RF3MITEzaT4pfieyKLTxSAUqO1
lSShDgZnjIL8XTxqrUmK+cabn9JyUt96Jz+O2sJRsvqHdKko+Wsx4WtobcDMbKBWdAwWXY/52PYS
RkkVOxfPm2h1JkGeQT4S/9CPk2haeyejYvEANi50VIAg6OO4vz25WcDERUbK5aMDpodimc/yMSEd
fmSStSx9RHnpFwGpJXlR2NHr/9pouQBdD3YEgmMlrYDA/EK7QiP4Yyt69e66GO6yyGcqGp+tDtVk
ApOagF/D86k3dF1tM5Bzt/08w8xQjQJPBQ1qmItdojO/FIICfu/ep+bWHzRQn2ASKSYQUzYHODm9
SufkO/4yUbGSJ2YU3vT2QU1fPzay/nxMyYT+DCCWMY8TzMJ7sAZIJ/h1ygY798Qfv8O5nRKfNrzF
9AfO/W8SMczwzS2sNwQdDVoq9DqzBY2cFrqphiek8O0WAJGAHzPQYaMUUcJPgcosvr609CbFUbCh
8v8R4uv5KPKzd2nNkBVko/dm5K43v5pKcZ4hAg42lig+hi8gxizgrGiu6ONVxOdAjrYBt6A1cX+E
HIFICdlx715mR5ymZV2iwST2TT4q2zF2mybmmM4j3YbUOopRjPEctdh2zRzka56b40i45J0O+fv+
UJTWCqHyYgoCb3yAcWDlWJ3QGLRkwa6AP/MRnhWrQBZ0MKUgZftJw0t1b9MQuJLQfq3tFMSkuG7+
OYG8U6xnIayp7GPBjSqD7MAo3NRhZda+HsXue/jQBwzc6RdWvYqwwESCxT+tY4KKj2GnGE+dwhzx
EYt1O70c3x987MRRATR7L8+eoWqZzFB+bwV12lOShj0q0JbzSf7G9bpzp3sjQvPSaQZL0sI/Q/ok
/KhByXo+RW8JuJ/nudBuHHz9nAU4kcM+Hdg60qKRrVtAEIRhdYXU6wRLSDqCyn4x3J7D9QNVGNyN
DcY6NK2jF+vQ6dWjhcfBSOslsLKzmajSn9Wjr3mFhFhrZ4ydYYwqUfrKzWR/DP0CFJzeUtrkwioF
sPo9ZRTDqgsI+nEV+j05GWC5l67t5i9lnBUjHSO7ktvYwMzEBGFu9kchkA1R+eLFPMtbg11eSkW8
G3GthcA/1ixrIJXEh+Rr84ZjIQOt1NxCcJfIQ7J/zCiZfmR5hmbmElQEjfaFWoElVgVLrHnxuGnw
b3YB8f9E/0C/meTLR3Hlni1xvmDKUltDB6nBpNbkr7wuslEyG5XWZAEppEPTMdNgNQU+ul+dfSOU
FhrRPF7M0gIxBXAjbfGxTFpfcKRqPrHFTnD43f1dhsFtlbuxZ8hcVETWNIaTugw624vxl43r/Vx9
un4bxtkAO3PAowKLMJ65Z6ABPZg+S36hz+axp1jbBsy+hpGj1hOqTAkgyVI999VeOW9APMYVSSQl
M6/zDQ3Cauv4auD8ZX4s013TNOy2KO+60/QgJVNogQgPJQi3qFJFrXH18WraGsMTomMmf4UYJWXs
VwQopADl4srZhH1pYsHXmZqwSpj1+/L0DtRHWeIdDsvN/S+2GQ2YtbSx08WEBaxcTTSkrC1IHYc/
xAQ09uQEQk5j82zKjnIEKu2z1czbbRicF8Pv2Iar2lRcECIH/DpY97hkXa+ANwigp6O0X9g4gJAU
PVsr7RVui+KTGihkMHucOwBCEsXMZMgH+V/bfyiebiZPtqoGsMpqHrtkE9OElrwKxffgTl5e4ueq
urqkhgow6V878CRyYK5dFf6Q6hzN5oHewsGSDWLY+/KslSPrGeAX6Pojkz96mzrauIa7gjnb8pUq
vw7C6rIsfuIYntWiTOOcz5EMnEmrJYsEa/OfZjVpp3L4I0T/avWZpvT6D0JCbBltlt2P2S30hKEw
lraUkMXvstp8AgFd4FHTWcISQGH6JdQVd8pZNhvYlHT4Z9LBZbsQ3kjFK+WqVZ8Cd4CvVQNd7Yfb
tuaVl9R5KVf3VxdN/ajVMGlPJgA5AS0Hrb7ZxC7Z3II/EI1ZE2eGRA4DV+0h+6yDuwppLvduOGKS
piJ1xCN7b1RNero4FQjCojHDW8UVny8Tla2o9ixg9wsaiPrXJgNWcbKsquIVe9L61gd54If9i3yl
7jias0GowVSo9nkFpPLOa8/a6B+VNRYaLFZkP5udvHhT4LgXpJbgvDiDkyhGMf3le0bXYRm9K5nZ
7rE+KfFZ7R75WkK5eEDH0NguPHoHKvx4FtWjOLbxw+hEYEvBH020Y8Y6RYDMDRhpACu8809GTykc
8+VlMgeGLh20RAh67x061F8EmeLZXr/azeZX4thkJglUwZWESrt0YMyg+fHFtukETR4Aw5Q6x1TH
s9W4IvGMezhBQVJjCavoVF6lwjczu6LLYGso4kLzu/EFVAGP4bWkVq3IckR35C1tkoatRxnQsvAB
rGIKHAJuLM44YP9lMmk2e4tu3DLywAh0yQUKZqCFWnjOUHAUrK/o2k108VvzwsRuPV76ZvEYEbOL
+0oPZ/nAdnlDOsvfPsCAS9Bxd7FqbmBsp9ZE9A6Ih7lWKD9Xa7ym/RialtkxqOMHK5uaxjmBsxfu
bT3TS4M7zElc96mZast9BpAFSmdllmwmQzkbff2vAEzEaodpJX+xMA9rwztpiPq6i4+qgYahsSFO
UkJZ+RANF7dv3uJumTDoUtdH9pHgVghvFfessfThr8zP+OdyWSadbYAGskBc0byhvoUKMBHvywZS
WZfPNp4jWM2kcH4URHKdD/+6Q9XU/A6HHZDooUjRPVrCdZhKU753PFvIMjFcbR75+tcnEFGm/NQ8
nKA+cwZ6R/O5R0FMSw3r0sAXtQ2bw5uPDDk1UEZ11e65tJFEHTMag8vPkx3Fv2ZC4ygy95FnN6wU
Sxdqq3Nvsi+sXEMXNchOYbK/oWsbUyc7KnaaBnT4Xtf8Sn68l166xmIyMznhFgh3AJbLYxyBhxW3
iRVVEMV1dlMbEk6VR+sc2VJ6nBNuJR4V7ZOgvZSWE/kHyEeZ8eO0ldPuD+8iU2hSCfocwkXJvxVU
YTy1W8wn3WemRX3HzDsz8A3XnG5m82cnacLjVfmCW35fNxzZ3QxcaZuJADUQSqCS0Fnoa0aagPwA
M0mpGK2dNo03kgkkuROHgOIgtKHF9o2VHSLsUmy5gUwKL2bdKhy30ZFdKxdT8WrK12CQgRj2aUHf
xNSKLTd+/OXccRLoPbrPsWuAaXduGG9Fq+OZOeNbB6uQOHmMxsupQfx3yF2b3uqZSwNGJibs6+8f
u1m16pQjLZIyXh/LTvTgwSYFZqB5qAmLTWoc7z7YNRyXxseh2YTPcYtzgd6H7es+PMSJAr9bjwzL
E9hcmhGWSZgaN07RJzRvYM+buF+qaiXl3CIWAeHIv+DNfUADLue1YX35I2giwij1KBDDRszSQkOV
05+tgn13x7EyWg9Ok000aOsLBGwxkqwNG1ozAhLMAdUHJwb21himuMlO3KU59ObDEjuiewNurW0b
vWKQoS+jB8XVz7dwZlWiu0TVMZn9eWXwgeU+gc6jekmmMW+JEA7JUAYX+jVqo3eRZgVLyy0n73Il
q9n9uO/wDSbjC7rYRXh9E4On6MBjqOPfIyvjZQwXLeJP6hCucoIpRisw56quPFhNAxEaxRraHfNg
zVfvSr4+YVVvUhSjqIdBBahYszgXJj3NEE2LECumdcAWPxlJwcVQNq7oCVUwb5BOcVwMT9GcX1F7
XmQNyRF85bRvz7L4wGABNolE6PUMdmcD0KP5SYXyT47nv1x/IOy1pI9n6+XeFY3xesh+iPHfrEsB
dTbcZsjkO6XumY7JSlYUhWAspIGGXaOnKPLbxyXygru/tbn5zE5nilyamV72leh1DhUmWPYYpZJ+
3l9NEpU0OMkgQ5I7GNn39rgAs816TVVNDRk0/S7Mbdw7ERKF8g2eKDlwh1vEDSdT2dSe5L3W8j8p
pncR8aH+ObwT3twMqqoukmfmqUkiMSACeJFlpvxZ88NfIEB0JsngkNuAjG8e0i6JAcid9645wTBy
+U2TA0ZWZ7BiN5XbkuErE24FuUgCxcyHUT0xbbhm3AGW9CR3ApwWPGC8J43zngy0ILRQrha88S6N
qGKCK0PYLo/aBWD/JrnrT4LHGVGLUB7lr2cf5lx33iKsC3BewmgHylJV2Is99sVae/05TS67M7lA
b6w3uwwvPe63nGvn/aMBaAA27v6AfapITkB+0W1M+eS09pTB9pSWWreNFky29mncOqKnU0RRSsDH
el9a6yIvJNNgjAdIIJUzelcG0TcCxKPbUyKw4G3965JxVlynoNO/42BUtVfPZIVHlLWPMbclgNCG
co1sI41qwczI9aj1x3VYRtoaTYiMIYIHX5BUM/SgNsoRIZgKIQv/50rUMsgr0X/wl+FDQn+Z+MN/
Q0B/quex2IC5/mN/mJyY9yqRKLeH/lHw/A429x31vfaGJBCkAfFAjTbD9Eenwple1jfrOaei5lY3
83Z7xE4f0CAe3Ax8/TmnMpjhnQsubmQ/xW4zI8SrPoxDWUaMHXDOJmtunkPs7GU4a7bBg33ZD+CN
HCu8dYdp9eDIb6SlfyzFJ40qMrgypQf1AaUrWRuYid34nHrWvU2oF5agieJCoMCSngLJhXl4DFI/
WgSBVp23YXxVUfAV2vGz9gIo6KwpyltaGtoLz5cxmZdPFrGmAYZ5LHYHVAbFr8GgW5irTymAXodn
90WHG/ZnjKsT/AOjHGdTIWD+IkQz7vTBel1Dd8KwECAWLO0KXRpbcNSI0UYwVfmim0HxqxNORNDK
Qps7jbteXCiVTfukch5dHLOJaRViB8VV4awvrbC2ZLsWysB5Z8+P6YrZJktKDzGG2K4ccAvwQB+s
z+CFP54/G4MYJxf+SHBDzTxNzGAhDGo/oLeZqg8fXskVjRYxy0Qweqt7nw5PAeJGkLTKIgg7Vqvz
qYEm4CpDIm2ycVlntQqOut7cgEvvwTcI+qkDH9qe7Ec50vpnMEtn5adXzuONHD0PSDgc8XXr3Rrp
VFG7am79+zlHzN/WkDLHyHomDzziVNN1deVJwKGH2FyK2dDrso6Sr3seNGqXf5oskfB4BjL7ouzF
+4TbGwQ/EFS394Qk1J6qaW+ayNwzB+1SIxi9EEo1Uxb5RBUqLLtMWkQdscnQCtA8L3qyKYg6cwWD
VdzIX86uZy3wUOqkNO+PrfLlg9+r3lEOjElr88XC+F/aK3O8uEGizYoRbeGnPIypjY8rKk2yi8IT
QkeAwJ8xRlgCnN9wXnqPF/7uOXrNQUZpJAf7av1BAGN3ndiEaVHH3XrsQVna4mbArQgACBGzfb92
5nYTtQfgi99v1nkCmjo1YTQsW1P+QZVDPQBWpjuDycr3AsD7V3bYHflPcbCLfOIfW6hP9Pw+Sv2o
WxCFvY4E2ECRHTSK7NSaP4YqCPBZ8LkY/3rBST7+ZSX5LBnRKvQZ0juSQZ0O38DLM2q+F5XHhdgR
0fN2Y4NFL9wcqpWy2l49zRDUnax3Gn452bNAx+7NJntNSyQL+wxt1yR2Ek42IAEHJ2nTcDQz0904
hNG0C9GRqlvTVf2fNsfyLzqwpUYlM6I+bAvr8JnyFq7Q89uN3ZrfPnvzPs7ImMpXw1q9kxNGn/EB
z+oCIFDFmncZhuKhErvLoDyowDGZUaWueMjTFPjCm62zXV/E5BYJs/vXOxiCQvM6xzoR4CX0soYL
ZxdIusSV0gLQklTbZ1FHGgisr/tR5lplQr7oTVrjvC9wtKDA9WuLY86yMcIPTEjb5ZV0xec3iNef
TjtoY4/2D54iq0mdceWVzwMlvqxF+rVPRBIqwJwv1WJ7dUBikMCLmSHpsFCZidgNdRzlERDEK7F2
4zQcHhpOkOdFAyqNP3Kmb+mZIVXMfmcahgmhls/aKL7m0LZ6wxrttIrb7mIBQjfIeJds6IjX80Hj
WWmzENZGEzmOEegDzYX/GwhwY8tJh5+8LDG/RrPMPVTNFsGdCXWpXQDzEq0PK/CT5MdDdfi/LByY
M8H47IdWxfmrWKQY9SKGQDo+wQujGa42glgq7vWBTgSUG9YTHSgPxfd8L2F09VP95crCzeN2xeD0
7Btq+2ncaZ35VE2zSgsI7bz6UcfSJ9/yiQ8gb4DgxV1DBBV5iAxAvWQ08JLDovVGDwbAXqlX7J0M
9cHhh1QEaauPn5Hl+ZsQr2X9Q09HmPJlUG1XB3uSPuAkTiX8KEjYz1jwtKUngGVN0HQ9kxpumu+N
U6dA4sBRe4bJ8U7oUPIac6U5+emL3ZerFzgKKa54ooWfbE2DBHAsfbfXOx+yyRUWzDwMLvVRRsg+
krdafZyUpi/IAO7NoOBkOSNvIQ5ktOJSDiskoUSJOcISdQK1EkHjY7sFFqA2NEI8FGqHi1gV3n2h
xmeeq0/g0fghDXzxMhzGsnzHW1U9UznSzM4vwkKtebknEmkUcI2piI4ytEBVDgUUA+/lQrjsmJVw
pzPFBfgdZlppYWYjJH6GVKknXfGprOtabfETxQAp9QCyOgekuPXDEj8OCERSwyZVsx7GzHTGTahZ
GMeRtLajWRBybFwkcxntrAjUqxhStAcDLVBHhwa/ogOm+UBxONzGImzIeP2Hi5FeW5O/6HDQHwuh
WG02/SmhmIADpXozdKHavm8N6Xt3fynMl5Fa/Lvv8E7Gmpw41/EWMzuG9PwdP0/a6SPMbuu0exuh
VeYLF++vW25BlDjCWZEZfNXEKsbwaFbrxcXJ1eUUqYq90ri1fcVE/fGsH6kgxRQq62+YJsS0O3fQ
4Cz3kYmNBxENH2bURWFyhgMMZtSHs9pXhQfGz665V14B9dXsVx60N1IWm7EQ+fZhsZr7NCdNkAWK
5nf8wv5W+Zq3x+2uOhnd2CGxtxTbvj+eVpEO1clnYCmSLvCDgSqE6ZwdR9bEh57Ka0JOeo2af8sX
/cE5/Yjzm380PpVuzWaFIdCW4Gk8i7983SIB+l418ngTzkb6iuDNBXiclZHIzGudk7eQUxfj9Ihg
X4/3l7PtuDZc6I4KtHfCYKqFxRFtI4ITb08JbYrKbOBO6qas70LuHQ9wf07sYxczXadbY5h4wfY8
HY0tjUlyQ96ZEwK9J1BSwvbz1w2QlHmEPlR+RUXJt/B50iUNtRRWKpS+aq+kcFI/2WDAe9HPazi9
V7dyqLmd+fovTmQdLfM4TN0Los5uF9fILHShwevXpXSDlM2Ney8SbZiWGlonNmhHDu9gneljXtWA
9Wqh6hTiA0FjMGNy6wNidDNgRncaHuh9qekbMp8YyiRj/Pz27LPQBzo6SVPAWWL6ylF/7RhQSzDR
iMZEJ+2Elr4huRi6GEV9bosmnI3pwlwtMx3GV7yAu17i3aHINqjktZx9XhC+y/fUUZ/0zfgkyL3M
VTa3Aa7a8upDbxRhIdhEMoPgYSSEDsDMhfN399eKI0b4CsgsGjyV3l2fPlx935Dr1o2/t3nVQhZH
rYoQx13FQYv0ef579hHbUhzyykgt3WRBiZAEQAaMU0pr5g1CgshApKKhaQFvW6k1feNTCcoLhw0p
Ea9Lai/nsBCpDYvfjcwRcrp92xOyIbE1h/teFhhRA3BknZ9KIyTIanLm24673+1nwhGTeWQSpJmW
xpCOIDsoQyBOMoUgNBPOeE74QfbN+NkC5WqWjQJ8WAPG8mYo04I0cU6r7OwRzpB/+nb+jrqr/XyD
xAF6YNldJkgZUu/GOeOyk0XsUGFljds68bthCAugLlUP2Rp1H0d3BHVjakWzzaCbPBYbZ96ysSIA
1lK4fJAxKrOHVbQkM5zFpi0XTOKA9xfkwXfVpzxVM/pm0UHDdzwZ2Qe66M+jJx854JMbwDWDYulA
XhvlKld2/aAsE6iTh5LO9Rn+xtAw26QMEuTtx9lmgx5GX0c3BlWaMdXsuWJ2FS9virxEF4otwuPf
uC3SS/FG9h1adMVr8ZlmX4XM7rT1WZyZQsUID4t40GiSldJSTjiD5Ksx+hAKcuYIhtQsoTRkn9Bi
Kc2zGMKBXocY/o1bfqqzYBv0juijiCLyhr6tHBbkr/kf7UsbKOEelL/dHlVSiHIKabB8ozV3F2jt
L/bA3YThzxzL0Bze/JJKFdNqyo+J4zeIE9vLucIe2zXL+ZGboNb6OP6eJls1Og1EOLAL03nR6/Jb
DPRYO935s6aB+Eetas0CaTUwPM0yPZPAvTWTX2w+ODDl2ROlGVpjN5O0CklVnm3Gldo7l7uzwYev
WPzB3o5fT15py0uUKKU3SERYrdJhlqBl5eI6HIyZzJLEPztinA3q+AJVBBQ3E1aHU3QPvNHmJCuJ
kbmD5mTa3URt4aCbI4zYDB86iSIAB2G9toUvMTLwIKD7yQoGqqo+/pTC7kCZuYIWvWT7zRQjojzl
Ya7+OrqQTOz43BwmIGqmpnjQUItfJofOx5OB+eDrmUFqz+egkZsHVFwxNHSt+kYOtnXoHIx/DW2N
ViElumaF+Egdr/ppOwKzmUJADLnNAfvlciKRLCA9kV90jgGhYJ73ZrOfuaIludTWXh+f0ev+SAvB
GuQ+ZWsthXBIA763v8Nq8P/pofOvlxonRWrt0N0Ov5HqAt4dR1QcWL3r3a4B1Vd8sLfklvy9816U
YzoZdzRjKepAgSjLRYjaA4h1oJpE1XdjkclPtTk/uze/Azxv6Y9dLkMI/gw0SxKaLQKqpUDZDUwx
uXmk4/WVL4CBh7zqPqwlNJFw2l7MpUt+VgCBFp1B0mM/WXolbGR9mIStrl4vW1qL85EL2yjLuzBd
y6sTlZ6kUKgbNtqud9TSuGUAApTfjQC7jK9TU/fz5L+eIIdEFcCezIxLTbVFISssYNutlsB73uMT
HdokH1fsN8VubDu+CH6sDNdnFlnwufNvvdWVe592dfiPbCjk01unXbpNniqhIa7WUyEoYQAeTy6S
2SOgnhW3f5oT5Y50HC+SyxWNPj4cfduZFlIGaUYkWdNTvZWKWVkYdiyZ48DJ8GX8ldNZjPQLGe3p
1sYROCMsPpGY+a280bGoucsr3cXWHxvFjeIcmpwogTJzyVHGUPoR8OrRfW02zDumXB8pxRXzI9BF
bINjC9OO+Vok/FwBf7vt2+Q2nIp+gSD3yJZW7Qw0FslN3+e27oUAniXXJwjJfI81TObKVIp4JPPV
Rp2w36Z4wFmuJvi2FaXqrgRjcaedwo2kfLZSoM/d6Ty3AFGhATingkd8FJnf7CCmOauN0iTK0UAt
/5i6utRAgVYtvXOk3NwYYbW+nB5xlGE9knekOa1ghbD51NK8JP6JnkRo25ZUxGesIP3f9sHijhm0
APXJT1ZFGEHjaFwloZQ3CGjiIvLTSXq+3xM83/bMnjFFLE28sM1ARmGfhd8H04Vx+SGa0vfnXLfo
eG55eckhkA20easG+DFM/oJyngCGcMcDC+s4/dlNPCD1hJLfZt3VMddnXsdiSAOrJ1rZB/xdD9pH
jBUMcDtQxE6BS31P3EfQeO2gFyVicqMUgQUk5dm4i3e0EV4y1xNvmWsZkpxSsYn8Mx/9gq09EGc4
1S1R1mSLDgAowLIX/IqsfRUzjqDU1pOpwj01FnTyblrX8Si8EOBzWvXNlQOLu1PZQWk5ouDspOv6
dTw0IbupELIHil1AfeHnTIbXtHeAoX3MwofXYpbUf6EKoyrhUEZ60k/vd5g5MgtodvxaEJDFHv9H
btyFtnXY9Phf3iHGTEAfuG70lVUYZ6nr+YLSFWpxUxmo5Ne+4YDce0008HQx6MtCBbFyq5Y9zIk2
mRiDxOYTT5xDlB/WVKxFe0psvaoUW18FvEUqhSXr64Crp596Jnt/H1h1NPPxIsLUDq2UXycT6IHl
1/ZF/yqKcr7EBxZ5+RiG9kpZeO7M+MalEqj28b+6m15EMsSfKZ10CmTy7q5ooRPOwRaRFQBjbYvB
lA1GNeGifsWwBnzqJyJ/tXjUKon4D/sfF+LGo2guBkk95fHjRPTvBrXu3N5lNE6tE828bHwT/emO
coEr8iswpCvSpswWIVYUyvTpuvVVUMBhznMo78mR71Ul/Ql2Nf31UAPzDMT7eULOchoUbASt3u+1
tk8B3MjbmJils92G/LzZYu0t+ULnoSTiX4GYw+OS1KXrw1ny8nEe359fFY5Ub4FtFTgez0Biw3O1
IInmvlF89q6agUkDnnyDvMe+u1lB6NUc58UTluN06eanv1OtYD2/Sg4ZYjctkRqjLi354+d3c3If
vq62kocVNJcEU/QFG/Sl7hqQXhOS93A7xr8ARFdAUcXWDCfNWRMQEUe96WJunJ0wpTykUeMCEgbc
9/xpfMnqh507MMKer/4AV8liBXXXUM965AA2Gpv+Za1+A82c2NXhi3G12ykpWhMZ8bJRkpjf9/iP
fdP5usbpKQv/l+GOl8oGWuvZ2pMzN1ndfBR93pTk9pUnWQZzd6W7atwR7x4Jkj/32hX1kKy9O7xv
KdkwIgSL43rHO6kuBV0Yn9+eBqQtQp0wSU/oDj2NZSQM3SPQwckyVwL4wh6vWCJK9RyLM1uC9f2v
/3G52EuEakeFgW4YDdBErCNorp2fhzbxWlhqGHrbH6pt4AS/D2WdHNpYk8odTayDuYEQWZvLID34
crBjh17AlkwRwwHu/kfSX9HJgJ44VGjVEbFyWQDYJzpjKIOsyxRYrFv8YhvAn00rArheCowEdjzR
+ISYmZk+VAxfbiz6G+fAMp0JpVPH48zk2Lh/xWCwxk0cq6M1MVqqL3aLWI0Mfp37pY6jUgE//TJI
ohUUD4WnUHo8w8yEU0zQdO8t+yCTH84TU8NkBfMcW5KtavreCYCiJ7xlHzYqDllxafcUlMQgOIWU
2QHHkFiijAzS//CXW8OClSyy7+CbQ0KaB9KBlgTcpgdpEuK6C7GKoqP7n4P1gvSGH0NwcW2neccX
X+A4e1HaTCAcwGMeISKaLpw/nUA9ugewzsdhzMLNHHlwf2IuFz89asf7NZhwg4P9NXU9uGeLAQJE
AbxBd4iMdOx4yj6Y6YCDre1nyTBVc58uxpYu4gmQj048HkjzFKZUGWxxLpYt64hvONe8dZtoWCEP
Ln9gsFskyyxu8itxcwkli9VIVDQwnfZ2YJ2Q6TxhFqVIWTSNX8zcriIucTVjTWJ0RwRG+W6AEHGZ
Hwxfgj/nXLNRhD2Poq5vdCtj1u/oNBzTPvlsL4eRfRqvJE0urcnLhCxB7F1mSfIzvIa44/wWRFAc
yGfzaZjseIo4XjQoN2jljyRKaoOTYBku77DTEcyOJ6r4MYMEt6JhscpiQZz10mCKV9nOR2t2rjHO
/jRTSXsw8P4v5vv5aIH2k65lk1ln9743qNo3K6fav9HiKGwQ+BfoLtSFA+I0sN5MPMSF2sT+a1hZ
6pgEEPHiLqAQhNwQEHE3CIwD5VvqJ+KYT/KPQgN1M3ptcikh2qQEpPhQAcnPOIQZ3oZ1bHViYrph
bOioOaZJGiyORXXkU84aD43lmT6lXrQeHJqHhf6587XpbKfdrTFpgJvaG8hddHKm2wBco6NxyhKu
ICuxYL1j7lzvQ3lE4S652Ow1lxVDDHtmz2en/JeWj34uNd5QTKOU5Vuxa6XrinqS675iZxuXOuQ4
qkxlKBcvhEHBXrXoB61Du9qkbGPBYtU4o2bQGJOs4zAD4wHeldp4DQbzezPgG/I9VK8WAWgc9dvP
yM/hRy5eBKdnGtlWZe8L+iEOosyueDYj43IGTFncPK4UyCImPyWgQbNfRq60WGsEJ+Htti7l2Tu4
9H3kcOxmDLKdypqYBhS3WkNiwwoXjQ1sTU2FWw0o4e2juiUWkF1pLq8OI6ImfMdeWGUaSwaXJjkG
GqYO96zLW/zSb1XBJUENpx3xqtZZtOhkzRs5XSvS7izmf7Q82MK6CgmMxFwmyuozwX54bh5hPVdf
xQGIq8cZij+BML2ENh65VUAgXQp/SIrcP8mclxnNFIcZYO6WiGto4SHHdimhcEWK6gIpcP5Y/tYX
aVcTzdKFQwKRAtOuC6QNV4ZQeBsAI69lZ7N8YlFPu7L+2RgiwnOFht8aib/bkYLewPYqbdgj2Np9
dtz2kUbW8MHb6zA83uLYYtjHk/DWqOjfLeGxVeVnKaGzawridXuQ+fA9o9vUsMKONg1PeKPMqUEj
qPtU+u4oPwFnJZJHJIlsUMFOZbCdCAxEE/N2Bnolihw2uCeE7cNaD1GNyz857KcI7mFn+aAZlgqv
cGojFny2BgKawcVkVF8YcRYlNFm7F4zMN9J8WTCDinh+/gsJnMov6hVM+8l9MFS5uznF13VnkWb/
K3zryh31clXmRvpYD0fezIHroE02E++79BuXiG4Ro1ys5GZFOrK9nNA26qTtYhsyKKHO5oOQffGc
kQscbn2emZmkDiPTtoji2rWmYZmNQ3Ztk3oK7+xwbzqMea5wNJtk8y0sE0NChqFHxTreED4Ds4th
V5uwwK2CM/ttKhjk/9SrVoznxLQcp9IBQ4Bqe3Ng1qRVG3GSZj616V23w69fwljY9ynqZGV9Ulty
5nU7T3WSVV+e0sYqPAuiPY/xOZP2Oy+rj+8XOLvsORlJCl80GG93/8g8zSPq1lZzhK5lhttzOlLQ
kWn4ETrjNKely03AafH2qGYtRb2NpkV1u3Clp3FYm1uw8xxGZJzy+nmv3AeXNp5s5PpTPCfA1hl5
dVPGdmAOtmKe3gISV891MjVIufqOkSE5c1zCOjjK0AKXKX5euqMaPLRe9f18gfxKDDUUX3qVJEvZ
WM7w1dGfYrC3sg8OM6qdFa51g9213dkkBckAFqcCjLrVqfkZZdOp4savnAdS2MUQ9gyCBeCSTSuo
3UuAYJseASH3nKFZbmaIG8X137zS6j2s4XhG64tyFrkNnj8+kUm2QQYXBKDzS348OP8dJrnOlXF4
B5C/QLvSnebyOEaiNYQf5MbBclxiYB9nHpQKeM1OyfMb1vQTyzEJI9WuDui3q4RL5oFu+uP1tAyC
tjE8ChReo3V8splWW+dPwtQ6V3TkXLvlDr5Uu4ZCYHc3K8svStw2xci7OEJXYeHnu/7i9AdsCnIa
q1vHNY8cWKY8dYzzabf6Ex9Vwuab1sPSTSKojzoAFIweP4mZcf2nBMmIT0An6DuKc2GdOBkOo95F
cDqEM5YC0e/PZOpYS5ejuhIPFTZgXJFjBF14azKe9kl0E5I05/nF8SQc+e8zReb/dfKQ4SldMd/u
KjFb1vsfkZgo38VSv8s3PJgs7SUxQHVsw93/wuQBoN4geDoVkpiKpQeZmQe6w6aHbkGor2buvujt
WnfmGoU+icheidJoWIl7qporLD+LemRzMtuCOz2hivgdinQfdHly2v+7wUFkS4YwHa8YHpXPFuNi
Nj3ZBSwzIJyTP3wULVXdptoTlTJAT+7dCIShk5Oi58lL2IotaP8vma27rAc+7PgGZsqFF4qYiK6y
6c629qPia5jZz2KN8Kk6EiQdteFSHAX67YctlqDWHHPAQ5qzjEtI8/7rD4tw0X4tdDhNB/gQoqOu
y/FRy9bON3DUnVyC96jfN2/NCrz16spxEIwHGL3+KcFhTeiOddhmNqaN2QK0AqSsunE2D6jFSxdB
7f+2KsDGb/hD5dQ+P2FaegFyN80getbzeCbzrjwxfHHtTOGjAknDYWVYH4UQZKvEWD+WFi7C4Hi2
ykxUbWsmc1s0u1HgHKcuK1Kz2KUW4H8w2rBglHHSyWyaaagSNjTQd9nol4xNuE1KeHTa26jcFLbI
yNMrqVVAP1+FCqnqgKeNcxKcq4XzK3p4EBXd9Db9edyMKmlR44lMVuhNcIlIK80B5Zbhtr8S8kzP
gOFNVyEpVnjgVKTE14VdSb9q9taMe9Yni2vlbQCtP67oXjL+b2syXWH9PgMN714QJ7+5Q2J47YCA
m/U8mtjQZ1e35+0KzDcysnXh2CRBP55FHtk9p7A5MUZcjoJWQh1eNdqv6s57L8JgWuo69j7Y3hrT
3hIQo4gRdKRsPZLwNu7wWWbX5kbZwNhVZ3mCPxf6G7lwXT52kC0bCVb4RMjUhnwheBsCy3fNHU2a
gvHSPWNVhPhiepL05dwSOS0YGy4xZqrLNlWDUMGNQGxHAW5/h09tRU83cDs+NL9YhHN5Gx3KLXcC
GK4B6FUayHAzOWHl47vNdUTCv8P/CSWeIZGYymWiK+asMKLPTRtlKGaUXS6asm94FuQwxV8HLmd2
vIjiAv/6jZmOdh0F7rEt99vJ4f5R9C7fdheWacEVeUHPVkBPZpwemAiGN3mI4ejjPbTSGl1j0IIT
zRUM6PS/ytoEjNtIdANlUDoCSr010A52PcIDJeeAZw9UBluDej9Gx8b+tE+j1jVd2mlRnN672bER
CC5KUxqgE4RsSTL3fOKkClDlV519wJ9pI6okFX9dUecJBDB1IzPiC7tfp+hQiGcNicq4Rf85jshv
bNz0jaV2jKlOeIIz1qsDmKVXLggVuNkUkAtxFhdCCctHuFw91L9/IL6WpbAOw6Dmw8dqMhisQ5vX
p0tURq7avpQhpahgz+5rE3yoBt87MKpEw0xtMdrjv9mvjPPuXVoO97D2+4znOUu8k1NbXqcB7H36
5dU28rNid6qKv+M517Llflf04glqTBAUhU7wpcIFR+4LMZHRlOB4cSv53pGEjB4a8XY0cxvVEacE
gadhoJtDeQTiSyRWhORNKDBPwU/LZoMue1f3qVEEkFnnmrWD++vfDL3oyRVKmfs8Iom8dGz53bu+
Bllypl0LRmxNQ8Iuc4WOTEv56HmEicpPPlzO5T4cCgbAseygnZbsZMPG1OwnsK1zBXubf+wH79gb
k/9rV78SG/jj1AdFSJB4xTwwYjrnDcEnH7/rb6X5HJZ/W00iTV+10cO1sRCO73Pbd13jPCtM9h7R
QHbJ9xhFudxkRcyrK+KP/TU+ovAkiGeMQM6cQEreb5yxF0mV4puscVBUWGEU97/PLRt/4rThzUYL
hofbAtYD9P2PYg5T4Xrn3kBCFb40BPQMb9S9IO+csZ2UDwYpkrHzxYul6n4AHWHqC7e3oAPb4dFY
JjkuYjL/aG1d0vsqIE6QMskGGsh4tvjINpGQ0nvr2pB4I/wN8Lor7wHvzEBFnmxOOiIa/J8tOM6v
owM23rH9eaqgAinIPJD9J3gLLyrjGueJQcMlDJBHPghGvXWrvNXvIfzeSqEm6EiEtCztxTDtsMZT
i8uzvbAX9qJFOLk/rAXViz93tX2SxCQEPrMBcKQwRMDE36GRhvchguhQbwFJMpb27VRfr+MqmuvP
xVHRUO+QWL1i6u77AC0lbR6xtK/rmVRLx9za2f4tDVrgvq+S4M7apEs8vOwXfd3bp6eR5L0t7bqL
CVIYglr05r1UpvMRJbPcCW1/vq3vCb+o7PDuJaCozSeSekHeGGcWdgqfOlHPWJkOkUYcYGjMARnE
v3jXsAZZFecbxBct8hvY9zY4v3+pf+ogTZ3yharomGHEqS/x/bpy4hIc+baHVZwEAVKIGCYMzurO
cSXicCLrBHmmQz9ca0hXjKU5Z+Glm7Sho/N3750J1KKiDUXkO4R1Qbb68/YP4sh0a+H3CKp0H9qh
yvrn6okSzFfV0GTk6xC1YrXuHCf2aflP20MsX/2DgWVeAHNewR8fOCzTdV0X9Nnmzvd/BVsjJkON
M/1GY+cOZdXD+sHMyhRcfCHvcqj9w03fDkPNxegTxIaL5CaHmzR/NM/PbuZgHSA0RHn5iwOqfiuJ
dZpsobog5NsXG57e3HcRwcJSF4FGvWSEwhcPPJLIz/KWtKDgpEbyItfTkdTMGKGFim7l7e5iKifz
j2xWv7thy7yE/IeEZdu+X20Hmvbk1VPqP212WK56r4DJUXhmyqrYI7J2V7TDs8BmoLGviODA1fSh
GP5zDtFrOnro+ar5YJ1a1luxjfzrDBwBv3dlyT+yolC2IKuqm9G8zF8Xve0+BopsNvgbrkrHRv4O
u+PiCFO0Qtl8gdChoqfPzY/gWC4jEaSqtuZLL/Y4luOdbj7T85ufcHP2W67PeaMZYs2tmwDgHQ+V
swo4xn+aH7UDhabW7YfL7FLX149ZLokMto0hEtJc6EAJErrfZ8emW4eUw6gv8A8WYk+PpyFOBzm7
agfnK9SUBY49opfL72UTyyWXblImQ7sNsd9taPIfnDplb0pHFn05+vVdy7SRpskW2JU7H1DE6ws9
/TuANQ8TgV0wvnflsyJHLLffB83mqUId/30h7JZpIevvDzfLVeHSXMvHXkvCTbFokui4wSbh9ZTH
xBEES1EcsNjCI18H15gVRbdhfV3bNBILe7cCu93bXxLVhMqUjju/xTER3Kj4zfddv9ZFQGFbiuD/
yKARnMvE7LqVWbIYFhX8kfmxgpM4NCZFCb0oZ2GfpLTapqnEsVzjSi/v36ZKBow451dVatPQRNOZ
JPTZjO9XiuYDAUSmF4noWPxeVnkh1UxexEWTLTdTDq4AKET+pE5S8akZ9Fie4On7fz2oix8zptTf
yPv4NpEz7iuQDI0cM0WGi2UyOo08LmeuXBzn4TdVhaBlQ5F54SKQF9SO+AJcgMlmS8W3TLzdvcRu
mXzphMziIqoTQIFh1jWKN2lhAy04EgHkNMbj7PNycBWcvz8hE9BzLa397ACAVyJ6lLDP6VHnW7dF
R2qiMCbNg5L04LlD77uor5UTnAZjQAAmtV0djqDO1InF15k5qNuWgXKLTfW0kdN8tZ5yXnyw75MV
UE6f+FyqReuuGbZBAOzrKYOhcw/RGyRQhi1qo8IH+StncGNZEc8dOme5inb1sxyNgo0VL7YMjGmC
0G2MIB0QUG9js1YtivLoMe4msBjoewZH0WYMiwsE05f6voM0UuZbtn2ymDvK3mBMy0P2CVld0Vuz
SPLAHj+3auyRah3d1KB1vfaUUF+iezsC3cY07iJOSW5WebdGGmHidXpy14cXUait6wEIDtbFiX1D
CqaEhbTd9mTdR9fL7a14dssyQNnWzAnh+ktn4YkmRNc+7t0kVh9bRqJ5Azu2CfISjsetKZcTp3Us
nrZargALfxRH2Pof3dHqDBt1+pgO+vizSHa4eeaj/JDq0Bc0W1/Ohs6e848XKozq5H9rmLHlci/H
zpS8hu91BLihnUvxQL5Nezghpc8XZnhBV3mGFuQjnklPOByCuU4L0GaziMHW0PZg/jj9J4yn3D2o
gZImmLc0F5cEuquzORAygTJd2fhmLMkEg5v3myBSq6y4IToUxmEwcfgeGlvep3QiVgl8cu1QXvU5
fXoUE3KvCjL5WJ+vYl90Nbc94wBmmjA3GpsQCzrhETlDt2dyY/cfOpr0YmrcfA9f8rFc8WDiEnYx
3Z3k2ztMwnGcmKefmSTlKp1wnryBtE8VC0ywSpaJJbFc7Qcz0fEX7RJqfHRv6F4zBoDCtXFlKlLQ
KcpaGOfPM1ulDxbkKHOmSDi5De27iYN7mJX+DZmZk999ZiPDFPnOswgrmPnEYIE9/ILpQ6bGk+PI
gKjFA+6EnhRDUxZKlHHqOQyS8EoB+ZFlIFDbWsUdJaYa4Yit1S3rOkt0T3tgNskDRBzCTr0W6iyC
dYgk8fTQNBLcge6LaDcevkv0yF4jVEYIgoymltfPfdHoTDegwUqC5kqNWeSz1V9W0Hk8yEmHUILL
i5Xg8yxM5GwWxElV4NdqsMhLhU9A1r0l0mFyj8wz9LpU9OpC9lEJEmkHRKHksSMJw+v+Y3HPKROP
H5bJEMxdIr3R0xM4M4cFgZvk0lCX8HfR/xjiAHOf6/5Z9DAbrJdPrgSFLs+KZyn7R0noRENZgofp
8TxFjcwX/XvcIKWnCUPLZdIca+4A9v4nxEOHpRKSakBdP4p1ZAUDBCejI/kI9Mhko4oivadZnh1r
1oNKCPdUKdgjvlp30P+ubi6ibDdyHwmDpf3D7KetKbHNiYfUk7mP3CFzClAPdUTxCHlHb0Z3MHgN
YMWSc9Y7sVI8M3N8a6/CxchnBAEhrITeNpa/V9jtX5a1ovxZm+FkXmYyzNoKOVisSLB31Z1T9eBr
RhDJLKTW7LNcic6KyJqKu/5hiSiS5HvMt+vPcY1isTaV4ntlnGFWitDv6gWI8igzeB9oRCD6iMSp
grl/o7fPRUF/XtEnMVA4In8GsCL3lExARwJGtQKCo+9nr/LcoDuaYcj/NnCivONatFPnpQa5QJrE
7/yIc8Ga4gYk4NOCZaka9JqDKTq3rsMA4F0rkilRJyDacyeKVvEZIUC2moy8H9TkkcpTwJxgbmZM
T62LLBM2jkwCp2m4bBMHUVQrgfm8pyH4RSi/WJr/ac/cXgYL7hePtjoAbyaHjeukdMhXNBdlaSGO
F5SciyLNLiEde6CQYiVbpGAk4tS1yXbVJqNM6cnvJDgtFshvDT3nkfSXs8NkKv1z0Ay14c0f/7Qk
5ZYyE/fbLEGQl9YD74vSzVsc1aDwExH6drlERhOwiNt1sPQdFt2osXcssHp8jnUycPcf9qnFrcrj
EGVvH31HYVlMrDDYoStbDwUIocUz9aYMX0S62Gh5qjeGfjsWOdI3caQvGLlUDo9vDM0y0kerRyLw
VXJwJsis9yMxfCf2D33eE1EudvfbVzVfOJmJJ/pLrduKkg2fA9sDJnwJ+hqlwAt+qQkKqgfwOmE/
JLL0FbX1YS2RpOj0CNh4YEja6BnAIDxxF1v/jy+lzRitKUCnhlGnE5fcGQG8hbtZyzCGNa+K+r8J
pBG0p8Hdt9t7xAFOS/LOeuFJaz0r5JTeK+LQaMRPGlWBM7Agm2vU7VRJH5OrJRJeb5OtmSE9LCRa
WBp8C0RHlUu8/QcbqizrpXPKsffjIJi7Y4K3xAMxZg6pNW8Mku83AjRFoU1CtP68M4bRQH2rlurl
Tf4s3zjun7BqNVP3QWUgqcWaf6Ke64mxD9m8R8nnrl8xmecfjkY2fxyaKk9H3oM6ojf8Ob2C3OJq
2BhBpvdlrWPFMcbx7PbBoK2U7ZDh4/dVmv9V6+iah2aigMSt5ec5nTuYd315QiogenB5zOC3zR3t
k1oLjYb7e7w9Sp8zBPZJKWEggReoiW+7wQqhaKaAvyvXCkjSnMrBNM+JNhJ5xnfLMrU4+e4mYWiA
qFaFyAAFyjoO2411+rKaRs2h6ZbP8QpaqhsaiIho9iEKH+PxW7U/V/9OeEMYopUCAPdt+9CCBwMr
Ef5wIITmIguVNr8QFJePZlUqjqbzVeKO2FRkRsTK3KcKXw4Ea7SnPNWUBL0BKldd2wD/BtknDGMO
gvwP5Wz3NQ281/rW9/BjV9E1P9lyfgfTBBrZs/ewIm+ClwAyrC7HR9VaehJXQ5H9HvcbTsxdcBPE
i4Gro63qhNLuf96qfxnayBWNaJf7Brez25NNlbMS6qN7Rb1eoUtrgeu1qAldQET66ZwWacYmbkhV
dt1fCSWYAy9+kyHhA2KHEqQ6neP8JSrVAbnQDsMfqvzwiR4rrqKt+64Rk5C6U9Otv5sHImzZdv4E
ijtZLerBHRF1+XDh62LH33i/E0q8ti2+tMP3xQucT5knXA/NwaCmTqVEEs18q8lQE5XPQQCnEyVv
pBgyYr/lN5j1BVAWPOgEh6aTGGazH559hnk86W/6i8mLI5Yoje2YISY+4mAHdGeyo8BBN/AVwvZy
LAOO6NSkaoMdEJzDsbyWi/27xsjvJsnjPxw6fOPeDiqD/Czf0Oz5vZ1FGt5KTZiI1LcE+dcwM/gX
GdsiGaZtLcL57xsmMq+dJBlSjXf3J5ljDp8FZZlvAJB5Lg93w34Kbm6eHF+YJH9y21yEuIHZHipu
aAaiAPNrjY9/O+XQ7LTH7uP/1UfRVr/sWIo4HZI2JooQLlw1gPTdmEqPXsCGj11Z5ixMcnmI/RZJ
cftH0+0M99UUttWDsASy4wYISUex8ww9pvaj1246wkeTnywkeeLAKk4fSmTFqiqOta7wHwlDu33O
MlzOVUUWmY2lko2ldHjxpsyBR5ADuvFXYJPeex0R0K2h/IBrZVHpUaxSAGCY135x2mEmSDaIvbUj
27H9QpTwBn7ByLj008onVKgvEQQ93p+i02AgQdrTKkDMeq3fFZDlBYFNemJ9F344Flc6xAyoLwuU
ZXiilYZHoxyKVpqFRRUuLpxd+ADz/oU4u2MViFfs9ZGgyXHQ6R8Qin2Hjh66gFIBdXCI4NhgloSC
35EWAdgOcvBdqrY1zbOUnMZbCw4Q4dGj/2oXvbJHXjDAyqu5bjI83u/p3zx8U0uW9rGHOyZBA2wU
svoQv0pzHmVAKFQjnb6j6SrVvsupscDLMMpFwf7AbE7lyMFiJidgjQRNRdGFFvEPceVDLlGuvOMm
eImtIY44mln5CUB+7fEQp4ltyft8Bw4W3RGINJhvRhn2SJbX6y3YPfY8Sy51sIpXTqs0phQ3S71t
Ksx0qySPZe9ZUvfpVscMgMNd+XBwWX1PEpsVzDh9FfF9lGnayG3FUsmPNt8gKnBveWNCU/LQIQqn
aW/iztOozZzVcmntatnzXZwxW8E19vdBVF5n8vg7cZQ5YiNnAfIdQjpDk/287djd7u9EjO7kTqGR
Fgmg8c8WmYf1smLoJHRGf/AAZCWKYMfyfTbCjD0QpCauAQcp5gs4RjAtll5SKlqGCugDLPCj+pZM
yST8l2wlIUEVdb8Z4KQa8tq+to23B1vKGUZaqIGVZMBcddQXHAz6g1ObW5ulbm9LE9cmRVp6liXc
BrLz1moxbvp0oy0O3gYBfxbqYU8xHVjiUB0hERKL4LGtvUayfOYfCcDP0kO8uLda+QdsUn1/7NVK
fAJiXtHWMNVaG6fOomZ2IKrnsVLiirfj65giw5kuQdwMoYVIJMimU4hCdGx4XBgO0Ggtn53epQrI
wrr9RcTPrmYp702086zE7DCvlScBZFr6jgkNfI7sSYI0veGnsZwEbOGNf+W70VcC8+St4qCsc8/w
A7h+kqf1PpOjV7HHoKN8ZWM3HGXfolHLDEBrQzr2mVN+zeKBJMDOeDldpiVMXx8byJXzQ2PeDR1Q
UOnd53sZRbpCNp1Xjk71uap7jPITIpAG5qjfKWufPQUzSbamhooTO5Yk6jyFMhXEBDs8cAwiHYVa
3pMKYUmBlesUM/+NYlM646tr7lrFlNIFDcazlf5CEp9yuk+Q62Q2+m5yfeaoANHxamZE19JGYXZM
mC/OJAPNEglEQSQJo8zHrQXb6I1jHzIKaQyEorxHscFjiJyQj6kcRI68OiY80oyAU4XF0dfcLuDC
i7LhK0HGqMF7pR56HFkyT9pdEd/TXxuexU20auQetrVz4D25t6nv5f9Zb2Zu4Ibed0wXqyWpiuv+
NCPA7PSHpes/nXCbWtMx9irAP7/UGAlA4cfuQ5r4x/N/m2mSVVjwU10Y5YOZfB1oUP+q4/7paRni
EmVDukyiyra4mgoPpo1I8w5N2NMZ8rK69/rMT1G1+gD/0f1bYyxMpQL3/zojnTv4qjEBbMEfIoji
vmlIXZD2Ul+JEjVlwIk+jH71vHzFnGPjz6M1V1Fx1ZPI6bBpL7/CBUEEZxPNoqDFqHCngqWP56hy
PRuA37+QG5BpjEJjgSwDfS6Vf1J3Iuhgexehmx4wCCAmc7lFiuXNWh+9tmI7GukLgJCA9GrqVeMq
u/cHx1Tg+wyD3B9r42kIlNi7zz5dDWQ81xvjSOXltOFAy9qufrMTHdiHhh1nQhMEXMD8MGsA68z2
oc0yW+VTCllKjPHHmSpf/7Z9t6wNDrX2hOFrXWBqpda6/w+1clO9Btp6lBGuGyhymAP4Ewww4sNi
4N6LeGlu+X6MAtbmO5QULqrdyR2m6Z634KcEOhLRBvukGdRp+PfCmbX6MsOb1IbQJ15BPgArLVE0
SxhNu26l7IFAqow7FL96JCC4rhlvhztuFme2by9nYLXirir4PcgByU8UlAfe1W2iNTzkwB5UEGfe
oKiTuB35Z9piheGetRqPHs515/vqxJqqnUsbc+XUyeTEScA63ADuR8QlmzV4ywavwvrA1p7X/yiC
nv+tN3ZTVuv5mkqy/LbsM2hCeJQmJq7uN/jXZpFyBs1SLQfZvHlne7DzD9bgPX6ygrxLGVvSpqGb
2uRlbnxs1wROwuHVC4Y2K7dcrQ+nEBBpXUDcmFhZeO5dKAnsMfQX4HgHEIgno7loYFPeHBTm/2sq
72z/K0sHYcBsKk2li5z4iAYzd6KlqfIqOG//18Mv1BAn6s7Yw0A4egxBssLKi7XMznyLG2oViz99
8jAGaB3fiSgiMUgv/tcPPlCqi8FNoLRMs0b+YE8E78KVpgj8nrc8Q7DxWKc8fBRKK2QlECmA1hwQ
8wzn8YbJm4e61ZxoEF1nOaCugteYKIMYFZ4P0ijL3PUjN2pGGLaFpFaQphJYlt4U0XjZLnhH8zlZ
FUM+hFmCLu1OGpCjlu9U0qV0Mwn+bH4vVcGSO8DueMyl/zl6Wq1YaPrkehu1jaCib1Y9GEEBA+//
YayqtynP20SdFZx/DS2vFSEzZE1QvJeKz1+8IhjEAM4PFRm1hpuoGYIh/OKhN9jqawOAyqKsk2kK
Y96B5cgwIhmpWNcKyl+cihlZnYDkw6b/eEEt+zxdRDHQSRgvtQqvpQZ8CFfdcMeYyrNhNsx9FoMN
7aBzv5ubZPsJtMfwqJymniLZzWkFUI7gzR92xJVp1XXSlzaRxYq4UzErHDaQqvx46OHYWqsao80L
a9V5lg+66HP3x05YW2TdHtsl1Uht/rgOb43rsbMEsJL8BcIMPFih81o6o8cpRiJPKxA1iVhd08ZX
wP8cHDjr5A903ZoDRpRSyG4r/C6AWUJvVhnV4WfeKTMpxgWpKFzCBdMvpCN5fLeq7wgvGFAmfv+G
+/YgKYyNYdMlbmckHlcQT8d0HZisvHI4xWpblpLYPdU5Rbuv/xUrM/eoRZqOeq6yj1iP+9BZNMvo
Y0G37g3D25OQ46nrtB207f/hs9t7Uy7rqq8rR4S8e9b3d+ItoH2EVlqtryXRxr4q3qTlN+x5ooaQ
MiH4ce/8SrmRXhxqCpBa8Vklhlou2Xvr6Wt/Ggx5UWfdgLbm5DEyb/10esTSPST/TOLBCuSOn/vT
FpKj5ZhZt1R5NgtQS/RTJ/RE3O0FaRS7YhDPHrvis3YKFtw+1fDw0fqgJKaUaeenaiSHyQb/DJUO
LJEH6YqrOP5rsmZV23VpoTBsNFn7A92JkDufJbej8/XW11Vz7YEv8mtZmQbtxwokHs4NklSZAB2F
aR6xsgDcUJBk6cnWAb48gWwGSE1jzxb6ScadyXY/nu19BBAXbVatU8yZmTcl5Qy1zQhGgbYby66v
rzRWYdRQGsietvPMn6WuKcDuV3QHTjexde7H4dB+b1qS2vhDs4FVK3WGeexGgFzpfwhE2SzzcyaG
h9+Lf3b8DbaiQG4uYGpbZdznCdZu7LIIV2ro+b01+8SzTm97EcpwaiWlc5FhyVr7xMYL6dX3wV6H
qeUf1Y6W7ox6ES+2BKQaUAYLHCuDS9JGl/1LsyvlpPrE+2V1AX6e/CTMZcvqJaXq9wVixJSQYQR/
kv5N/d6hB01lvUopJiVlpOCv1Mc0yqSS6qU52RutH4By2i7LD6v3byGJa16ivwz0qFVvDEqwr0C2
5PCEEpJ/FJMcQb7TAD66cHoGNOJfsIoZHrubQo0lcHP4ArHDsXxNj4otMBT9vhfb6gDR0Ke/ZQKl
Zl4wPE6rXukEDTmn0jiUyQXqKnmGXwl/OhylchDgl7wkmd24OSWjrDbBg7ktPjt0Xqk+iZaUvYju
xtYkuGO8nMYuLxtH/F0ZHnD7SfH4wVeHE1U32Gi7k6eAbEGgGs6GgqOLmbhNoRzNA9qXKiR/zYgr
nC2ub6IKScVNts2WzltjQM4ucF/pWEUFq3nizFSBqDhcZIiZBrP4Xqqz9f/T0zDytHryHNjcLfT7
RM4Ej+FoyapCM89h4GlhKPJk4/U83FgSypOTVDx4ToEqs9H6KptdOxZxlynkrQyntTAR47ehG7iM
h+BrUAdizocQ8TGp/DhG3W/Zvrb1UJEQbXc5ML1NzC3tkfdHw1vnBpV9N/E8TXVNHM2uJ/QtCkcI
7wnsWFRQR95HCo+N94EcYwY98wier5MoHJ9Pmy/stKfMmsS6Ps8bmqR4d3ut3CNVSePPKY1kxgsX
Gg84FVH2I6Z0MGRPe2sYK/WBzmsbkxERbgNsmWPwib8qC3IMyrvDf8Rn0CyAQNCiydmjA5dCkn8u
ula/BBHbbG9mbFDkb5fWUQF31KCpgjfHkV3v4zx13Fhjkg8nl1ImmR4hdSW18nv1rmRe68GPkatQ
EoUwBdV57G47dumMjAX5g61+DRMNG9KkO//I4/MQ5OpRE3Bb3axHdM7W/MMNmBOhSJPSu/uS+uxr
2IYA78DD5sEZ1+ocCb6WYBltxUIFEo7GEAQ4iF9nddUcOZAYO4TVniniEigeBCrx7tsZAmEx3TUD
JzWEV1ypN4FAhL7B+hD6pvST7zjLNf4h/bQR8z+h6EUNMAesMkjoB+XfGW9JH7T/L6fEYIUWjZzC
DqDNJWRNSmOU/vNz1dAUUC06u7aGqXuTxt2Y4xjqkQJ8f0PD2bPkBbLnAn3wFWGpMdxDEIaC3har
0DCbhd1ZlSRIdoZFK+VIAKMuAgQHmz2h6bq51rJPrN4Qsg2M3H8zWPdwBhLGUYzaIcjY9fZuCPi3
02fmbPmpPv1LfRjwB8jdiLsXv2KZU5VQrmb760pDZzO0a4VEqfS/trJwKwfqXQmhhDUj8TDMI9Aj
XwQsN8HTi6axgETUwfaEGxekUVawZrqGiAye7STmLUxZjYH1ewFTi5s+cHC0uX/DXYvoNwaAeq+z
zJqWfzazTIYw2qR1mSqF5/aTnz18R8P7djOZ3LAEt2HManW3InRhEWC7pBl8sK8HHxbSu3+NMiyh
YaonAzHgOFkgX/gimIVXE8k+c2pVRpBtJw6PrZaZhnPgBv9sLLEyZxnP6BSMCRgZzPkZNUr6u762
g3amfj7RwWt4l6RokYCuNPrpxpoy9iM2PhkBKoaNNIWhPFMx3/VUY8ukkv+77KFvbfFvx9OAnSEC
hLyMS+00qwHLgko6BzHU5uNa9rahjd1Ky4FCSR82K901qAERFr7JUgqBjn1fjLz7rZngQj5RIWRP
LC91vJs/n6wYrYq4/2bOa6YW3UF1zBMJRchgJZKNEmiM9YkD5fpy+Ckk2annJmn9TaBt+ZkDj7z4
ZHvI0aH5gaEut1dpeYDVQUAKE15rY+NAcpE6eFEJy2ZK/eIze7+riOqxjLOHC9aqxfzRAc6MTlNi
ZIo+CIxbN+dBId/2hHbBFR/06x4Ign1p5kLwHt4+F/adK7FWcTV/xiIwu6MQXeNM0zlmXSTRVz1g
vCyQF0f8Q9L6ORLQigosJa+nCNfS4nx+AECxAZeZ8RdM+R0EtjBBE7jmxvUfKDTTvKk7P+7tvJCM
B2ABXGFNCZADi3RDDMsGQ6rQY5Xb8cBrEIju9uUwrbawJdKCMEeFqMFWg5kPzFbsR8MwQSlDXwsj
t97isbzWEPrMifQSMuhKdWiy6fm8O5wVw3BHk5L7BcnweY/lNIQKZk12B51brbpsL2oFEXSpJdSN
T93h0fE67BZ0j9TAdzD4jtS11629TAl9GUrWq/fQRYECSxLK4vh4P9pR3/8tbxgXEvyik9Fecc+J
nxweHXiSooPGy+DhIMmfHlybd1u47nE9jcAAZvSWwN6PgAG3yAMq27wjRwehLNvY/RL0Xs2X5SJ8
favWLmSfFrit1QV6pu1ElwD50PgnrllTOIHIaaQ47MIzxGiYy8/nIfF5i6oPtLte1vF93sVdcqjv
cxEPSXOy497B33/SugstzP0aJfpP7Gww0o84FTzTFD2uY+clHyELhlxwnHxskU0yfn8hZqatE1EU
TLFWpr9mArXC318+jHyMG8gV6npr3Mq7n/10qRAGOBsSPtXwdLE9zqFsKI/hV2b6tzO2XDZgYirl
tEOjYPTUeFIrUiaGPIjxg8O+STUkoFGNeX7FIz4X4wqPpKkilJqF+uuuACC3qvVgVT4+2nY4BSbY
z8Y6xiFUH3JBQQlv3UW0odDz2TSWDkYzLLFpnKF5KPHMnp13P/slLR7Q9Ng+L80M8ZnPGN8tbtvv
VfV1Sg2q1tbPYDKJQTvvteTrgmhyIdbmRNPrPbiSoKVd0rtUSzs0Am+HpM4lpuyl1DUncLryHuYo
meWAN3RcnDjaKEa6U/TAIjA8OPX8Z/qfHldC34Nkd7Jyw/RSB6VwZuGkycgFXGLIbSNLb8DiLYCy
txviwHT9b/lbQvvexBhJXsuCPn3FH6TWL4ztNV6msZ+sy9VbkA+988u2udZMWlAxRgyvwJfP7cwq
6jqPmufv1zvxwj8YgB2u6vAffRb4ntdKPV9W2vtB3CbmLs1StwOsIh2G9EwIDvxlJmO9hGpuZWN6
0A7SuWqA8D6N661X1c0y2bBUDAxzIeEd155/YWefuMyNOxci6c29LxHpB1e/wLau+DTDpY1Ss+xS
RbiazP89MuxlM6Rf8eaBY8GLz6vD0iVb5VBgIwKioS0B26TIFy2z1V5DxHlRXHFECAgjAcrZPcnL
rV+OxgRqQSW3VIZDvKMOoZfJQhbPSKGrpNdWEIy9hoxNDOzsLnWYScD3lOwcXWKp1VfZQzNNEy5y
wCYczEWdVFUfHYkTuxVrmhLkzZkcQCnGwgDj3qajLNLcRDgBWpAUfVIuiibK/+ak39jjpkmYLDEk
mFa/YqBvXKKLI+ZE8AYLGUekzqa/P5OpPOLsXgNbmbut7bIi+KRdi35T3Hu+bNx28NcAPb6IvZ0N
E8mLygCWWUNBU+lLaQqyPcugb/qKSI/gZBMu2q9IeA84EFWWxlxQlz5W/yqcjzWRiVo2qS1UrEiC
bC1ua214PfizP6z2Kqh0ePRmbhY6XbnqMqX8aLVv8lwN0sHZ5HTWsy5HL/kBHnXHNmBw6sIHBMhL
+awAvfn8tBKaeQA5HAMnUyo0mQeW/Bm6Au6iqqGr0ltP6mZYxqzygm9Q9krX62QIq1mjNUySL8uy
u8p9XXJla7K4LZEhmswgGDk8+AA5kmdvTvbWzmF4Tb80eiJwE2/CEHAk9l3SMz6btX9NHGi+udA2
bJlrVoRiGdBe36kiN7RZwFjRmdZElSOXyZRcYLFXuKyxgtntGbOSD+LS2wwdfo2rmlnlgVePfMTc
VrTB2Y7ZUaRFLFCpbuyJ84N9PU+vfP7ULyP8aH4dE5KGw2Q0W/lghKNBjDnsIYIEJTWIPIGTozbX
LLC2xRFICik/bqCk/FesSy2w1SIHp9oYrh098b34nk1CGWGR4TwMN7K+6arz/R6pvfkt6d6seLFF
oycvFVmvVp1Ib/WnhinfQGXC20IKym35UDLcS4F+DrS8MLwo+dk+YFg46shzFQZvdkt1UgndPSiD
JG6pTg0pGuDfizMNWvdnFeCwFA0cLixl277h+patmPbR/l3W36qllI2/UcTAlX1RVo606Cldsjl5
HQwQeUhrwqafnAOnYGPvXyxU6u+gCx6cDnZHsThinczyJO+htZwM1vT6I0+iy9+c8jMPkcml9747
8pm7bwNf8DggmYYKnTiFiPl/rcGXjeJDUue7wnJR/DEo1WGH+D3Bb6zHvUcaQr8ahLUp9FaVv829
DKCXi4R7i/eT0vQ2kBzEN/9RbV7EuUXIXYnfLAkFf4FvkvjR/6BajdhNSOqXug+d+ubYh/JQHyRC
+mhwtYzF2CzPQFK3FuOzgYztZ9HlO2dA7sy9F0NrIBKITnEB9TRRILgxbe6eH2SMf6zfJWmLfGDp
NTcS0Ng6DL4UUeyoiNLtZaBZJuBF4l/VgGzaDDQ3J7qLmiVf2ixlev+W1pMRl6FkerU0DpRd2CVR
XiL5816nGTNRAPzjps4uD3tL+mIJ/W/fmUzYmQUnTBPRwVHndHDWtSjaKnvWJQ96xgKK7CJvcrY6
z9ChetJQrB2F6mZ6K7fp4SR38AcJnLciV+Hn2+/OoCq1uygu3Y+k9o7UzJxGpYDroxEYvtVJ+fSS
NxBOH4PbCFzcAsIy8viZXBRbm5JBdyOsZONNkqhHW29hdV6lWhw1D8/FuDvgwT5b1f/I2bJFMO2m
JWFIfPhGp7iCnIon+OEVzQBjlwD+Vn7p6zsr3663PRo8iZPMJwr6dORiVbViG6I4Ow5T+J+zyUZX
oOtQNj5J5MU+JtHMydOjldLXycgv/NrGl5FenMtMvafSf72rsyxnnPfnsLIIP5yRhAHB+1z4EI7f
tDOKjA3Yd88pzRuxdRgJnuuFrHij0RQHZkbSqtIIUtSc4wi1nXx2vQ1wEqR4CjoH6VeYqEZKMibI
BMlb+kxK4VzRIoik5APpYvytNlEM1ndB/p3TXshH1hoeJ1JZjRSnm6SrMglPXxXdabMiJHungbrQ
4Rskwp+eRloddeMyrB+rVPcIUTF2VpQII/XOZiOtlj5+Y+hndhsdgcnw7aJZJ+KfYJSzQudqb6W0
jwQCCnqTGX1VIARm0i68jGi+kuyYwto2xHtyHiOfc/mRycIJc354BZSl8tCBMRRcDHsjYAJn/hqZ
XwCQFNrAH/h7Jxylg8Xv6r93wMvoK4ZgoTvdHz6OfRyVUoE36rqSH+WMHgdnfBFm4uRR/vMVv/k8
VMnlfPxEs1W2xhfZxtUSZUaLR/yFDtXbERSSC0F4ymN0MLnilU3v53LzZ0Zaxtd3vsHhb9w9KkiK
EZbM5E319Y5M0m3kHnGdPAnE+cUegsspMCW1QjNRM/9S7CpLMLKC1jSqlnyN1gqBddtGiAdmwXmr
FOPFQhTGsJAgijyS8VKbtSpx3aOeMJKQxA9T0OYlhgyub3HLyRbxGRp4m+Gs71eUuopxPtqIG6BP
BcLhJ/Dacp+MioDzRGc7jtTM6rtDBAuJxancUWav0DQB5gP0hIMKwbRx5b79ktm3uHu8sds8LZSJ
Euetuyfaj2dhz+qQIT1PHp5bTnZeZ8RcjyiV+zPckxuchxV9Fl7O8OgsieZoJHAVG4Q0hmQ193vl
ITbDHTj++o+fJyBfLSLmhEiuFkDpOQ783Zks3SXL6eeGh9KWI1xG/CIKgzGMYwg3Tr8cc1LUt56s
gFfect5MIUFf2fekUrUFqQU2Y/pdy0LzJrlTqPUBT4Lajpw31dWoBQJw47h+u41xeCInFkDJKJgZ
0SrTX8XykV/LrhuIw82rUvR6sddbAng+ChyLsI+UgHuGwr90cYcHD6tMNBO2XDMVmSSMGz6VBEqx
yOPluS+BSxuqYBkRWsToeoLNEnM5Fw/n7wARqruDJRSv3zXkbqGtTXhgXWVZmnj4USIejaCnpsKe
ySFeLup9U25rAuLDo+oYtgYyGZUG0sEF1QsX7U9pYYcz2hx2KBLxhZCT1cJaajb+wJFxCGgpno4u
ZAWOh42i/gaikbUBo+QCPkFsM6CmgMAI3IWTpVTsTohLHHC+sRb+ro9U1oTpqBEenLMlyFx++Ayq
gyq8wmSyDuuKsHb/ZBZUqRGBxHtXF3rwfrsD1I4S6PGv97/J7e+ISct+6Im6m2fQgvwGzIn8I+7w
lVrfa2VqgX474bc/YCPUY34rRFDMIotK8TXGXr/Hdfklg8N72fV6TrlFhtrBv2u53iH7ruE3Pm+z
tEepUeMR17V3e4+YiTQJtq0Wcka2qxrPcMdB6BiPvisbkeLAMj6VEvRq0A9db+m31WFLs+JJFePT
sAE+u8nN5mAWV0NOp7jILlYuA+v3HOd6RGEIcyEDxyJ3pnz1yBZjCCOaOIvIne/RaGvaXfe2IsS6
bFYj6rMvTrZY4QUdirgJKqkkNxQbJXfItEvmk6qT+k+U9hl5rVKSvYBlsFR5hUOgZkrvs2mNl8d2
4OzzWbgxBJzDhd9uY3tiJtQ8jiCbGm5QgcR/8GrUYTikVpHJsHXtopEUOxm3cwzeh4X6otXX6dEh
IBTgQ/Q1ZtMqaal52dMVU97nbuu7GnZTicNiUmoCieuSsXS0RaGuqlZdgmFMfzIWM8pJuRZ09PZ8
JJkuMD3S0wwelIf5FiqYW12KA8jpLEZl4wW48BeAXVprDalTX21BMdsQQyCVfjsWXYEh2zcML7dw
NMwej/Aj0lxC7lfG1ioGcpuqME2Re/eYyo6q03bCgk+ItpWYawiSJdgn3hPFDalTSrR44DZWtqzy
tZvxbjX+EKFs0Mn9nbE3n5zbf5x+cJriQjaeLFVJ0WEwkQEBo53aezgeh7roiy++qLGcCQg8AZOV
riUYW3W8WORtYO2E8gbwHlNelHObru2yc6IoJ5t/b+g9ZhAv9K5KdKLPHdjYNUMyajZOQeVKkHD5
YcrloBvl/XiqNTdjfCUSCEaXQZgcQOrG44sOqC992F10pYt/Dcl3acJsjW/8+TYrTqcRLq4xMvl1
ixnqepq0NaSpvqokr0vViNvB0wgr1Zfyn7WvQsqW+zR+QhnGzq4o3xvLfgt/w81Y9efqLj11WHDc
CKZMVC1Amr0+4TIWd5omcApZNUZ3exzGK/4AvfM7jUty+0oDilYY+2p7scRBS5HBa0xPQTCJYMFU
S+bpEVbsdrVSnhJM/WmcmY7PZU+W09S5yHI5m6LFW1OpwxBTtDFAEBeuOEdrzYx5Drk4cNN45hY7
sGucqBnnfttSqXIcW+ETMWUJP12Tb870sv5dok/50d6JWTK8f1H/60Xr2YP9OgfaRroInqLymi2Q
aXrq6DOE+xhdFZilol9kfDqfvkQrw5mdigEmXMw3i/UGZYDsJO84iwfiSk+HMye/mJZ0vnaL2z4p
eelRjBZmcyWkhWe4YDiDviRAj5e2e17va3zVGAbPpjCdzZ9/xr24bVCQqkYL0T5ozz909wtl181b
EWbnlPT7J1LR8HGvZ6KT1mrcBZor0cw4kw7ml1Xa92djP/+pnYGjqcIN1UOQQ4YaRHd5cipzoA8o
zECIrdDtErkmsRdy0PeGCK/iK1I47PQC+pK0aE7mHYo+mXYVa9O+WSLcdVWgjYxgOy7INaxviRI0
S8TzXCgDg1U3MakNZ6DBfHrdfiBFfaZK+kiCl5Z3EPCznRMzhRmsuaf2pu9yakhiU++z1VOtVv0m
3KE7JPUxg0nCp6NWJYMaTmQFmw0SLZ/RL5ux+9as7exxinu72/5qMN6wAJMwRDWItiIoHo0rr3mk
v2UH3F6N3h/MRY0SX5S5Qe6BQUtJkq37WWCAgTH3RCbcajJC2o8ZiEqsguYZk7zASFfdwQstWYqc
cVSKXf99M7JSRwEViSRSPuYSQV+xvi61wUtyLv0+HbMnLOyldradt4PXFTzRog82JkpMN1bk48kR
P3zqTcm9z0c/d+XEX/Xe2TaKY1pUnXwL1I6VLClKT2VMZDQTSP320i6wMtgW8rXDreSiKn3kHA5Z
zSO1D8MFmt2+CukYpyF7z++XsI5pba1HLQIrn0itrHerFnaFj9/c9WpfG3c5NYkM+nYIMTWDCW5m
C01iHX/hx2W0nu6Vi3st6+125Mc5C8PaWla5MqZnrrH3sXbU4pHzkIHE21VNOk7tDndkUG83EZ69
HzCJpnzr059Jpky7INhpdhHjk5XHJR6znREJk0DJGSbVZEOZ7kXudDIL/nzGaDusEaotLCESUs+L
sG3y9IMp9v/8QYn9sZ7oQHHgUFP+lQabUedl8UadRZyBPdFxkVE6RgtY7g2zkD68W/oSzvk5ZG4J
qfGGZkgQPyczupsZOaTv8ROGJT7vwMkD1ySR24S6cidss3yn0+wDcViUuy99Asu4WOfUFiBNbPsp
LHNSfGgh7d6dAHEDha2SB/Po7RL+u4xpUU9xntXSvZRrvGjuOiZK06hbudcaNNAKwG+gULzVXLLv
vOS1ofxPcq6Y2jdiHRM8vqadOZhI3wQC9TGXySA15hS6SOnfsiWxWQmRslAUwt7xmyAVd50M2wyU
Otwq3WvW7BI1h8x15W+c3bF6xz8vE/iYS5F7ETnOUBUxnPzBnRUHTo47O58iPQOVJ+pyKDOwOVvP
XeFmKqzBQd+UFMaLc9jWJJpH2a/P486C6lrWV5+yZ6L3Li09FL4HQ/4jWceW/r+rm+YqtjybWu95
j9U1TKtUtXUPyQN36HZQa0xTIMm1iiM7duVswInk9OXImHsb7doizlKputNa6/Rv/YaipY6MtAcL
sToIR9TeknFiCVZob9X2/zpxc4EiSFuqA4gcwExm0CNUjNcdXro1+giFZeIQ9u159pDH+zsoW7/U
VKCgg4FjSSuYymdu668wFuTj7U1SfN3ETN87COSOp6NxekbAzkTYLl9tm4RljIf90E0C9TN704CW
eag1V65Khf9ZmtR5Z7YAlPWXafMYY0SZemL0l44zIenXq7hGR2ileL1Gn0H0wHpCkPjQQCZaBIkA
SCBICVDj6zvLu03wiLvbkmKSd6lV25i3Sz2+WagZS5rlbSZQ8q4E20mEydhopJ/9yEYFeo/kQGun
+RTcF9T1nW/bO3+RuwykJRY0sfvT3RWF0+usm+V+81Vw4MjOYxWPq3+co/1NiYICW2AiT7+V9X6b
6JusDBG3OqlsKgQhLDItM8aBshXzXTOStRAJ10J5GEfUVr2UoHk0sB804QpwEmxpQz1uSzeaQ7db
9LeWTbSgZ86jbeBhDKqxuXFgyepQYfP8rK+h7aMQltSE4tD2gon8CisvsVClxkUvEcyAE65Tsflk
KktPdHeqEAR8Vas9I8/0fRcN+3ZbjwKNT6g9CbTa9P68+KPSA7G4JpVmJXCeyvCP2uJRE0i9DUFb
/g/jaecWz/W7QYmdDWuiI+8YdmLkiz3Su3PjEilenfZUdh6fwip++u3SNNFLicu0kKzeEzF3ZBcz
gnm4Bv2H3RO/vjTkjq0ufClqGfd476f7h69ThIpo+Cm/crIlNz5ycqCMnoitTXWBsVlAvy5/rDfi
qyV7Y156Mf4S4WUckbmU1UkWkJ/Q2gvIl/jGvtyyWvRJ2KPbGGScfANGhVwnxA3DqfZc9qspuR+k
ZPh5Euw92zkA7XipiAlKU24J2M+OyaYZhyEyQ7cp/NEHbM7dVP+P9FGdrgUqChDZ/NCaO4gOhbzC
3SusRaGfp8h/JS/UyC167KRG3uZ+6rkPArXek+ahzdlIAJrp2qezGXztjiinqMvt6NogZvQafajM
kcEOfRjB2lAp1Tt3r3ArTVbF86FO8m4K12tZQO56SoC+Dnz5r8PWfWyPfrTKGVvPHaen2eM162OV
eKeHQnGZwXroZQa0/pI5To6A8gB1WwCGP2Wiudsoa6M3maPc7Hfeq3cRx/b57hjeohiS9zBqlh6J
+L7DlZvEqOnljEAoztuKTEyIu7fdufhl1TjSBstIMuc7Mw6byEs9OwncWfDfWgnTURLB24BFeYFc
VSg6sbt0/7AryBgVwxSQdd8L2o2PS3aZDlQjAAHmM9e0ErjPG1yNYTmrPm1z/uomQnLh+usSs81J
Zu68qh5PqmdoBXtP6GivtcxD50MYhrnqz4+UJ0rZIIbBLVilxpWb/yq7ycHRg6SB7xwTbBMcIFoO
/lF47T9m9WYV/1Q5AqL3No4zl0+RJ7gAOgsA4kS7KuIaOli/FVKi44KdIfaJF0I9bPeu/yZe/Uof
5MOd7a2E9Lh0WMvfGNv1MWnwmwPfkLWmN3yl8LEYEBUzzW+F7BMzToTujZGW31M1CalHgZy3yL5W
2BrIeHjm7Nnbse495eqx8Ws6NMYmAZKjUChZeA/QRMY6f0frW+QpCsDht8gWbD1NnLvIs8MB77in
uaPouSco/ScRcU1f8Oy3sp23PA36M14OEe+jT5fal/t5EDj9XrnMQQ1So8/Z+LpN37BT3xUKXOqN
ACjBFUpwE1/A47cxSpTQBfzafpXV0P+tSXY7nGybFgSzF5/UURwufAbabi+dcNG9mvXL+oUlHLE8
7TRttF18eAuSVG8bovf8F5dzBz+8wnutlD04I0OikmJguRfEzBj6jS/tyN+m9iw4q06Kj2XdSqvA
VfTE+/jFUhjvCLKMgEH89oXiEHVL1sCU4Gn/BD/8qe4nbmHK782cEJFkJxlAmpf8h8V1olOTSR67
YYbW+znG0QkjDbz1+iMwVH09py2vsW65jRwN3JLp4SRhaGvdUeE7HVry4ESIPePuoJvaPKYr1h2n
IlRfzOxC437DvbmZiNu+962Ii4FoE61U8W38anacjzKLoXd+agI0dzbm0ng+yA0jZ0mj0vfiDvZl
doXmJkhoEv6bR3qBpsdtBECyuND8Zc7G+2afUZfQQ9/ntzv/3Zq5cld9gVktgpIhLJDTvGw3jT5Y
qDM1BnMlIUD79etaQgxk0KQI0IoLHV3j2fdmX/9SWbdPdQ2lXqUEgHMlFJJus6+5BKI9H+IMLMsd
5HEwB5+es8dSlxnqAUnej/aB7FBD4Hk1kKhnf6FV2bcLqvg0h97KBXA+GsWL62+/MhF2+ImuNr8h
cUib8YKfGnmOUC3EbL4GC6Gn6lSTAlAi1CBOhfNKB/HzFlx9flBkWKKrxyTXk22yHT8c3Qvk51NU
KqFUlmin6eq6qbX8AWebXLnDuj3hMEh8dRJQbL84BVksRvf/1PMfWt5pdGTrmmEZIs6yHjDBTcRy
5NnhN/6b4QReyF9udcoI7+MS5qixQp6d2hBqJUcuqfQdmbeoUBaOBgioGVQYZBIPyB0ICFLhhulF
AdIZDJWLjPtOyUbXzivcxXpugJlP5bEOz5RnzBsKpy1oGQWgyjKw7mVJY2WVY36TLgJ5W4sl+JfP
Sev9AK4iRtR4DsUqbG+mglFTorxr9+YVCjtX3H0209pVOZbfpfDRA50klA4mgUZSChX5Wlpw4RNo
9b35LacH7AFsjqHGx9Q+cSJptalBVIRykX09wZdJLnBuYtpfPiAWev+JQ5fu8bSd9sTitDF4nT07
7dJ3jxXMw079we4ZM/g7iCk7A91JYU0JUnwIGFf4R+x12+K8DSjLKQBVIIshHxSDmg7mw4MD1gDF
VmnVbHHAQ9diVuYAN1LxVBY9qPsXfHSvJKAJ6UQZ7yVlIQRQIM2ItN/h9kHI4ze89nrOm3VVLA0d
5O+YTjR6WDW2M6y27AVdcvtQ8NZSKLekNfo2I/T6HjS6BDqFKd2A+IvFkyd7QT0dkk3loatgaDWg
YNKxQSvyvW/z7pVpfebOGvhWIH+y1UNnpv1yQxsTZTnqfhkrZCOUazr1vfPypvMpT9X6T6AzCNXy
0fCnLxiwVAgNFGJpzd/l/dW9lVQs6wpAZISjhPotaq8j63avCEu13x2lR27vDJXEtJgf+V4pfBrY
gO6o08zVDFuIRVM+eLVbhztAuZsR0uW5s3IbRxIK+45fRrZ8lcl3Ejz3y9kvsvd332lj6IC2u4XA
d3Oz+d8/V2RZYMFNH6yStpG8KSafYqcWEn8FdwxltlMI8ZaIqMFZMQzPa8ANrgSEkwAlDIZXuAL9
jBEWGZbjQlpa6SJ2+LO0dt2P6mkpApfKofmTVa6YQoJ+GM1ySsqPKd/M7wWvNZ8XmpBqENjUS27C
w1wloh20InXD48BmKIx/uX4RbgwRGjPefdRvpvMK5Otl9xbV9zj1iQ8BPokg7MREtQJc0fCSws5Z
O5dCJ8RfaQhgM9D+oN7kd4E+7i+mcWPjl4yaS5BELjVfRStmjt4n+Bg0xqW0xDGCTUm+SJ2/uk2v
ExVWFRLZ5WvDB7eVWJhT3U1wLx3tK6rRNNPxYjsCyVR1a98fMg0V543AF3oKzCCsqG/N9S7hUSvk
Mq2UtdYNPF1jOcUcVh3gGk7z3heUSKjsOM2iuETBhrbnYhqTawB/rmbtfRKNF9Xds2e37EXXBGYU
EX9/9PNJAII/I/ZwxY7wOX8fATJAdC3QVio4rP/l9+ClYTksWPmM/qVXyt1/CAm9GbqxD8x9a5mo
3ubkiOz2zojXwWp4kdgujWdaUKI7Ge0ovT+/FcHnA9fgLV6JpXJjLZ97GBDDUNcxXYn1IWrzt5p+
cZPBp82o+0QlZJvWIa7Xf8BrdTgdfsKFr67JgLatAzW+/y/eGD0G1c9MmeG5SnGyM87b0reSZxeG
7k0HMzXjvIwdpsl2/HQ+tPbJyHR45PYkYA/YtyCvPQkj24YA0fhuRYZPrpUaE9Tc/WQ2U0s3WZJu
Yi9gFyhOg90O45wNF6arwLJSNpQfEoawv0iIwpsYJ5EKzdcTQ1Qa/gXhGeZeQ7A20mjj985WYJVh
F6lJbTWW7QGlutRw8xbTf02zowgVilXaezzo52dtm1VUudXJiNhU5n3sGjStNZ1pMBC/3Ceg5Ewy
CkxtoIwOqHdPuLvmKurMEOfOyig39FPmXxYWPXpFfxYR4a1p0LrNNPsxMeuCfMbHhXThwp85ZAMV
FhqGMuqp/4K3ERPTf5gt2AHEbRk7EclhqRcQU5aonuizeUG5BbYtkjc6X9mf005L7wMBP7lO0VT6
Qnz2uLkASEYRNIFkM4mkh95+Q4o+iMWte30TPvTZZnJmQRb803RtY4sKPYeSyKWPKADsqmcHn3xo
hPJe3GWeFezXYQo91in3wn9HvwJmjuv2jnLG4QP/bleF6l0sVo0gVxcHWAQOubu6GyHHAxL81zm3
+arb5bF5Fl8An1/MfwoDTkniF3XzwuSuwzX+lzKmxdysfgnYOcWwuGkL5oFIwvgvEwJtD6+bWhbt
yjjGJj0oFQq+gc51SfxSoi2zmLyE1uxtQBLiAj2LISba6Zl88j69jYpozWdicHv3KpB7X3yQW5jJ
pn/ybNIo+6EPmVksgbERvuxxvP5PMIh+DiGJEUGsTldUvLIMZvHni4vdA6tdhy21cSilO655AL2Q
qQ1Hk7YQSMHv2bXZQSZHjBrF0GRN2fDRtwEo6LyMDFtAjUbYrRUyHyGdLr9wTK6BXV+Q+xyJFhKJ
74IR621tl8NjlCwKGI2ti7YAXLSJ4OUQERizPuVZRr/a3ZRPhSa1J55HKlG0F0iiE6nxmlbYbJQT
QbEcSTeX5TiR1Cmt/Nh9x3cuflm5wiuaXNJ2318GcNdpjcVpXLAvLNquwae3LtBC0XvcKW0n5/AZ
EsE9o44JI1xCIQIn6mS8IRMLTEZFcLhWDlVgEZuBW43x/HLVIV+S1NCWlMknw9WdZWHKmQViH030
ZmtmxZtA3cNltcHcPMlYlStoAB99ob7y2bnIi/hM+MfoI5p5UHhuGKDtxhIUMlN4Oh45wqO0IKCI
ky7N6CAcGGNPNDtHFA+IcFeR4NrWgryc3kRVIdfheX27oNwEByRkfwYT/Y1GDtQZEIdzOBUZ/kGU
psoLQx5v9vm+61aTNtjcB4JuScdXUG/6+YUvcD5bPX/G+EKK38LSLtROXDVEcdSQEJ58vZ/QLEZn
bE2Rj+xIYU7Td+o/xH3lgstnB3xeITdFlGYGn/0PRgwx/ErIlzih23pQp3MqWLZuPSn1JNyhk5iE
1LmYgGhowQofAjH5R2FeihVMHZQsSWT5SkH9adGxovSePpCMEJXxwpuJ2QZX2zCHg7trx0wQvQWR
9v56JzBxOOyDdi1y9oOGVjWhbt4qRYi6VOay0+8gfI/3+fgBl0a+xZUWOf8uowJ7jHyw6G+MZ/il
hfEa8/5DoH5aZ8Q1ySiKqt691hpz031fOF36q//YvJzUut9DE5xrzGU6AjR5xeK681+0vrJYZsJL
YuNm/oE59CIAsi6UZCPMqHo1NjktbKEhgYZiWHAdHRHS2kHUzGs9XeO0ERDUQfwc9ThuQquMto6w
ds+pJEp5/hJmhdU9zbnum0oCpG+e6Y3poN4zMQE84gyn8emM1tYpgY6hhNiwXr5GQfcy+uexZyCo
aQAdx1U4MK6xKa//srkilWLF7CAMOBGXhbx4kg4SUWb9LL2I2IMLFt2yYtWKUIF3IT16ZzjqO3C1
qi07wZ6e611s0fVJV4r8jw/cjReh/E3yLZj28dJ5OP8zcp2Uc+eKEtnIO87ewP1yruSRBXYClfiz
MfLSefnFb4VItcRWlNzhnMBk8I1+0IF4mYa3lyduWLoopZYk21zyAq++mZ58yTjXDoi3iHYnfU21
vB7rrLBFt/iEofoMITaHvhsVckEPaYUFD1vIwg13sY45MAy0J9/22x63I+k/PMJwtq/bJiflb2M8
ikwX8iSAkwwI3HIY9YQhyG4JMpJsmmLOArYS566hzP0o7Ti3Ptjz7sR3s2MEbIv+LUBEkn4ffQIQ
+wbA7uRezlF4kBBkI8rfizB+1U6u/+Z16Pp7HL9ox4JZR75iOlTfSKWcsv/ATTg0JNEqDXEKwdD8
8b/9SHJZcA+bICIWpVCYCK8JLX/BhhvcjMHv+S4gtsJD7A6IpyBg9JQQVkGbIOrqfm+cWoxwAScJ
GgNuTL0F4eGcpV7qT6QlUKms7VmmF/A/wWydLVZelgw77MZDuuowiAEAkgcFAeFa7nGph0yuKOlY
EBinYDl/YiyGQqcJg94w03VGJ6w251ZEQON6P4K3/Cgy0wTxgDQpJVAqd6Yrsn4oTi1x28IND2Zc
AC1jtJ0J2Fp6ANG9ndNu1CWiO5VlCnJWMrBwH+6LMx6tgzNZ3M5GQv/9SErWxoAUurG+8aypjI/a
jefW6GYhQTAi9D9sK5cd1FUab98VnTGfBqmwJ5DNjDnoqqUz0TLKULfRmfjp94MhIU069kzu3Hlu
FinSMxg8U9DJLF/W7325c5X1yVGxCZGiE1E2eIP5OoVJmrFMcvSJQgIZcah38YHQSuX4V9GjBgDC
MODgUXTGVYMJAaL4/zCF0Cynlhn1D/9OCwF4+Nd6GL9ZP3jQoX5AiaRonakZDVDxme9GzL4PaIFH
VNzaZodXAIuNV8svBqo4W44SMbsN2+oHaG7TIeuVh5sI3FNsjNR4eus3DhSM7uu8hoxmKQQ8Ig2m
vZZPIskR9fMH+f5A73h3p4zUYcDqN8UHcRQvmfrnvaL/Fbi+aDChympW78jam/w/SQhKUKdX0sYQ
2BU4Zo9PvlRpw4/g1b43itkFeyOSmmcx3kbbqH0u+tchvzLz5BYV963MrkFCvU/Gm0LKBQlIVhUD
lJ80qBtQrd2bTnIUkXG407QzboujsiOpRDxAWZy9kJWHyiwKStSCmnKZSTkxOJMVOCgQiXomCoux
dNdMToCLvAhTjxzF/m1Sv4Mlgzpr88an6rbRH9ViVNwBiwed/yvcGkH43fHheCBjNk6+KNRmLzWz
O+nr9YzQj2sk48NlnhCqUe4X2E5MSYiBYaV1+AIz2G5OJfYrpGSphiBU+LjG9pigwbqm+Vq+6bWJ
k8XoceESVBCbX1YpUfJWqfnQYKgMItFbnG+0h6dXSDF6Tv/vJqC3icSQ0D4A0KD9QTH4jmtP+Cr/
gh4zMmSkCqxK2EiH+Y9KzC1XiHFH1MTzG/fFeKQpuoIzeo83XcIskGNSzwKqV82fmIPJEqJET9oB
tsl/L07jJMOP2jx75CytSZFK/MqsR5vTHOUJyjnabXK047HLHcVE6NIqTziWplJZuHn4ys0uXSER
AQe5N2nVU9liBzBmy37oueyL9GUIpV0y26QIBnkjQ+qrJ1FryQR8fzrVIif9NcEac3CC5OLN598r
YA+3oHh4/e0MmP8rWXsvaPQhGQs6YIA+wykpBLgBbCzoSUqWDi91p5hObtI0YJpVjCPKBB4IwKvv
ryt1S/KswRCGTstsyqMK+xACJRd2toPKZuDnFTeFgPeuO4XVamdj2tFQPBsBm/MGT37WhyXgMlBR
AGIBqdBj8Ofnx8UH3eg24B1x5+kmCt/7CyTG44Y5qXXe3DaMAV05ml3+YddQw9kvZOiIDi+GuZvd
Ag0nrElQQ1re15bld/OAl2mChFm/yGNfolMjleV5yoGQ7F6HWhiLdb6bJsFx0XZkWK7ysLc5jkvX
IxkX7SLjpjWTq9TnU+d4YoFkAtNGUfZ2G5G8vM/9GHfd51nPWaEV6Wt5D9Qof9KZqDQh3RG7tDDv
6NkXGHIfkf/h2DL6M60dl6v4ubtq3sUjqF6kjXnCro1tvh95seqpqRp0L3i9ajBD6vu/2nzaN47/
7N2/cOGsNrNP/e5eGLgqKe6dxaF9zR05MP8vroPgORvT+Ve5Ih49pY40KabrNiXvZVJO4OOetl6X
rBnmH9y159r7t/v4BGIWd9ef0uZgfvoFQDIZFzt/BwnRbowC0bqE2yWsY2e6W5hR/d2sDIFS8jpQ
e3a3xCRBFpCES6oy65WWyO1t3iRBJdsRJ3UUsAcRC5Ye6TkF6DzH0dYpJiNQl49LWtyJoAycjiFj
G6Pv+YPhPMxSiDhxVCs0S0ULJhHV1aaeyTCvOx0B9/7R1FjSOJxbQhAhCea62MVwO+bfKjaUg1zv
7KIPbYtXSB4FnUOdk58x6nxrBHbUmqy4KEPdIEUCUBgH5XAQj07QfBLjF9aQO78Asl938wA53kn9
OEZNl8wWrLDk0Rjk+nM56loMqkGzqX1yCmwPIx171PkjMXdLJsOr22LS0t9GHn6MdWsyavg4g8SD
s2ihGcUbDgJWT9XGbe+OWyUsKrCfc+d+ZW/bxQc9gYrnCzd8NETUptL0SODWiKQpr67TeNj3XWjp
7QCMM8he6fvmYrr1O4NGEvVCf2kX+Pght6Q6bLmSUxClx83yeetzkPCR2sE2iGTresFgXG0qlYTW
avi9D5jAFnQ+cs0UGAh55hEEmAiYkkok3tskzzzceXa5cXHALJFJATU37YTxBFX4J5gjzfzrF1RM
Vi6OoJXaBBu4ou10gEt5mMx2mCypAJfeTWsU3v3Tkd6jDMcFquj2g16ymuSzwsOlP4O7boobufIL
PY++yi1q4XQ9fX5dPw9A8Zfy/2U6L+Tmr3So8hf1YWQ8NAZkjAPvozmw+9JvnxcMesWhqxSW5tQw
SmIy9Ulp84nBvhxYwoo7btWEE+hVfpaemsQ58M2OmHh+I4drYW8QMMpjfG4HhQXjOxQwBkwRdFxu
lwoPPBQhybhHVYXOuiqbmzEF/wJMMQ7MzjJA33RSgWuq8oF+KDf7pBY245Zx9REiu7Kkq+jChL8d
uBDVqt7bpXbpHGFyUZg3nW0lcsoNIBzRvnxowDBdwN2QhTAipWP/IYmuxEO+F1mHEz4bftN3HbyC
yT5hEV7nfn5SElE/vcTMzd4i5Bs7GHKmMeVsn5isKnwfCTvDyaUP7Vtb3aFQHVJxnwMvO4cP0Tyi
xRQ9zxEbrlor1dXq7XGjPZ4FLruR1SOURrDH5Fxydp0WJlxEnPisGwf0QQAIfwqVdBL5wXmydoXL
rUc88uA8uTeMwF6WICSVVROSe8+rdCxdFDcy8XyzwnvLoR6Lii55K6Wo2ncTpRnqV+9uY/OD4daw
lMNd8yRs8FaguISK7gSGMdPWevoIJtTRRWxZEfAWBAHRV+8lYDvCtxV7bIttd5AwXiSkjloW4Pb4
8dVsOv3niKf+VFWwi4w8OBdjRuscdL/qSorjgrE/rtTPI4cKEgpr9Ys+qbw1EDHliuWQ4hawop4w
mfwF0opHZo+dmMgz0/6rtbW6qUtCYCOEI2IIpyu4ptKXogQTRD5auYla/wfeX3CK7D1vRbjwwT5e
PYBXCsHnWcHW+MOSDSQ8+wRO5xm/Bj0KcSZpAn1GbjW5eN/FBYG6uXr1jDgfdKnsEQZLyOAM4Bpd
IglwpnEvXEagTxrm0DWyPsVVkO7c3SN+UBQDrVm/6HBG9bCvvSV6Z+mUeVxmf9n/Yf88C8SAC92g
a/rzwCBAGMfGp/7NsSzNG7P5/H1F4Od9fPJb+F/TxMd/zRjzqIuP6//NJ2HeMjKJ3o2nBixDBHCR
lElxZZU/PuMEoUhTDTapeEUk5KBOEAI1MiIAWdlEXcK67bfcPXGDhgaCNEsMkfp4ULqzPc7TplRK
5MKRXQwTavWNJNeQb5QWvl+FgV2PrgljKzpoMjrd9xH4XhsGoGee6Q+1fP7dwtBElvZfwPTKOZ0s
6HxCj5iCcKqiHp8rT8OhALuvixESG3FNi58OhiDnFVjGJREskp3NtVuZcYJaatDk5QKK0E3b8fW2
SMsFlcJXvSc/mDOqJNEw0xFdeCdfFpO0H/e5vfugAQY20YvfsLOU973cBvgduuFcYKmQHfIJ/tZV
xgt+T+jM5HWKqa3SMNetgYPx3mg8aAvI6n0Zo/rg8ChxYv9eUgosUo+yrzZVs38CD8y6vnbjqEkt
oacHHUP20aVeUZiFhKPfTSF96G4RW+A6Ra9XRxW1h9Ryw1lR2B/Zcln09qjMXZlkoZtvCWHewQd3
r8/PLdFwBkbNaxAmosyzhhwsNDThi6IDRARDcDz86AxJG3V8o4Ll1+9WjHXTQpOCex/2PoQVSLib
jVVPU5Ob98MeMKmdhwu/wfYd4H1tQ0dHrJo5Gvwp/UCwyHLm4Q98hitmj3w/hMe2QUlKicnYgP9V
HJ3r8I/3IIPsBWsnmSD0J4gx2mFtRFvikni8ahb1wFNIt9xj1wQ7L+8YOvkWfhCwA8qAvFEWyXt+
1SvKTqWF1gy5clf72r1E3qpbkDeFm9ibkHk3DCvNFEsBuFvtTP54ZzDPRUU40V+2PnagR2b511g3
rtacqiSgmjY5FYdBATfYV3eaUAtZ6wUFsFdyi2jLSvfyPg9YYn3ZH3l/sHlYGnZareYzGgFa/fQc
sF0cS36v+w77PpCCCg5tf/WMD/CjcFOdyfq8DecS5xQmFaKg/7+JHxS7CuLjN8Pce8zaghcvv2Mn
MDAxd9v7l1TwJDx1n0RsD1yXI54OJWfqspqdFP4ZFNi7MYpYSqlqrhXfyHF7HK/AemW+oZ80pT+b
mNDspEryd2MI30FAnVR3egkT7K3TDqylgr8WAE7L2ksb6kEOkGpJ0+NRFkQ2LEXoFFLVI9AFHpIB
KhwdOVVL4BCblOYIfS26BWc9h3ZFkb5iFRoeZuM7nXzqlk1BXjASy2bus++JXKNK4lGm3nD0sde+
K3bLwHHGn/QAjG5DrSRt9d396m3fFsXb0+6U4UNp4nAj5rK6wzLktR7NvvaIpUOkmchp/Nu5fdAh
y26D38SAnxSa5Q5SeWkJZ83NY4tw14FYOULjpPgP4VtLyURHAof5ySR5T75lnXa+Qkn1CUsOs6aG
RgoF0YgC3cY4TraJeH/78VU8Czv2DysSP7GhgWgIv7KqDQZ5nNq+6EZp7Vz2wlJRmOUZfVTNXDnw
Vx5k+effaNpM6lSQdgcKL0OtxJBmZgEvh+2kxQ+dgensfNOBEjIiei8rcH7c3O0VlYtPzXxi2WAq
1g1nWHXh1xp0cJt92FbEwvUAV1RNX6ovbDVziANz5u66caRLy8WEuKYwgqhGA/YZTy9orVzYweEC
/dFZnuGk8EYhQI5RgEuYQxAISKhx84BFFey6L2eWQyFiOA/HpNKwbdYKHnywXydkV1W8GLiubsSO
oEZPQrSZcsP6CXdmmTWbYerpUKNosAhhPUfPLMHUtkT8Fi/CElv5QIzU7iMAhbJGnhTzAgY1eXD4
OoZpAbEFVGW4XNwClLNAzaSJjSJFITiQprlQmz8h5SG33ZiW9nkeKaBLN/QKwwAhnhJNbWQaZ5Qf
+E5ym64iyO4g7X/lJnuVQ9zY96FO1ozOvAX/axydnfsjLbLRRgk4ABCJnCN72nl2+RVcd+QjhuPJ
PBmFoeiShK/U1fHN4n+NeNqcd8+9eFLxm034DS1YyGSjjAYyYxPnHc2iPiMUrszxX6E8XtRxHs8R
ri3DZPnWmgZqtTSVmL5m4zFc6fU5OPRbHWZoNyWhxk2uTS4wFXCycmO0wKfunutvrEOHXEZrrTzD
fZskdnRL5yz7Zw8UQXs+wifljq9E+R17SsmF0EFr83SypgZrKgNG2GTurAr6vhSNdXemC1EyZTp/
jmT7ybZd5f9BJ+3IAx6j0Do0GPYXNquHTJwLfQ0DRjM05154v6qMrFGwvwopjjCI8SAE9iA7l37H
x+m8VMdBnBRFvL5MCf4PGXYDzcS7FU8EMuCPetmvZxYhJtWs66MwPfVH7SCnzbL0p4PhD93Otoz6
okzxqOin+HkHlboUjKxKUaoNbHgUb6Otk88gHoVUJ3OuyyjJTTdV0JAI4WUr9RsmvHFP26jnWeRu
1llMzIw1eq7JNgvFZriLYFDd5wmu/LJ9H+EWo4R6RhM5K8rUDhtWk5CtDomnU5ZW5CposY7Feq/t
9Q07UBZ9Gl+4CU5YBgpxwKcz/DhjIrIkETvLxZ+Ge/UY34l0N1VOeQGHYwpqg5Ma+KRi5prUPx2u
mSpKki+7L8D5T3a7POb0wpaCFWkqfcK9ylcBuAfYE+l7s8WB3MvSUXpOutB+MiTT59hVaIGEX3x6
27Jr3nKLiD1/Lvp26v47+IZYLu+0FeFaYog//Q7vIqMDd4VAkH/qUFCLbseN6Q4HI5Lwhtw8Nx1n
HegtegkjUtnwmsY8sg670AqslHc2Yh1OGDzmnzyrtuYvtA00SbHllrGLG0oEohLHA8CDr1v9XdZc
9b/qLYluwrhZypQ1VHnFl4ckf6FVAXI8syxOlTjM3s7kJzVy+c8ici6o4SUyd2xA34f+9M6YtcVh
6i05rwzpKMH1XgT4jNq+Q8KcjpevrJlvUh9v0h8bQSGf6aUXgRk01dueVXFLPLH948Y+26aThdRC
cdGITlOLiMoTOArymb7nVOycELXy0kdZFA6cIcxsoEEEJMcZBJvXS3F09vy7wU3j107R3lywnNNT
Pf+SGnhVad5ZgDRvRFvLqH7fAVH62CC2C9f+rHe7sOajNUCF3JkyXB20DMJqegMAbVJK2Bn/+snq
qd8vEBIjGl/l3Ucm1VZ814p+e3NCOMLJ2kXZZOzsPPM77mmzP28cXd117PQ6CgmYraug/C1juvKH
54PNWlsIWFf14mNIB1+iyvxhU+pqawUzjV5nDm/cruSWduF2LvluX4y12BZjYUjZgyJjXJU+TGTz
1pKQYUYM/emyR4rzA0asrqo0nYKldbrkpcTsjVafiyhlkiZ2bifiJwt322aura1qbHuJQQ+EsdTq
xULXMvG0+UzEQ/Fkzy2app9xYAb2419ZJ1ztGCvgeH3rBSEnn1A1QpY2hEXgkiNRwOjLGhM4Ot2s
DDGH8SgMzFvA8Mz8uKI0/TrwJK8f+F0zuyVwpv8mJ5urUdlK+/8txA2zEwuFJHfO4YgwHqqPyb5a
uqf/9ZqaZ3Ar8UJFrvymkLUurJEvcLQMwm6TijC2F66ZmitPg8B1y4u7RF9zDuF+jnzaofD3tftM
hzugeU25b71iZ33bKgSJdiwQtIru08jLGkh2rrD6Lkueme9uE3/EVS8Zu32XOlgKrIja6iUPtWHs
Q9wX1rSYGsZ3Wz7Wv4WnpZ12bgFJPdJZi86ZX7jkSBU+VgVcbbL4p9RRIakBePU/8P0OpE6Ig/oQ
xq9aImrGtd84lJCdEueNBJsqXXG5wXBBq8pQyjqB979YVQldApSDbRBeKBKjgqgP9Wp65nFXpxF2
TaamkrBh2eiv31le9mlApqEcGOeRo4wEfzFNx3elPC3N5xfakxUqIv9IyR2kf9mpJqyrjDow0O6U
kCzBDVa5+BAPtXI7T4s9xr/4WTpMiOXRs+RPaQpSCMqRtFCAuIbWWDqID9pXKkO90ATqfxeLW+dp
FG7VPg5PQaCHY1OR5ylG5+TipqgK2nwwM1eP00y5g2lh2HhGWpmUo6hvY6mFMnbQrb6PqSqJ8Es4
EHgjoUafu5C9DfVtj1fkvt6o/pOUS0IgsApvFjRQBxKY/5Q4E4ibnNIgTBKQdbXlHXlW/7kwPjTd
m8RcUCasqZiv6AQyRA9ukzVVKAYQFasR1iAeoWRrC+67hKUux6sXHRtuFQVtLX4/P+pI3LuylgvQ
y6+54g5S9AUb4NBhwKutgnOizeRgEh1/kJk0ab+RKVNgB+1qNYoJymQu5putkn8/707rCJ3Qdswm
ztngGO+3AL76Dili2PVx3BJS1JgWPDo2VDc65XAVo9VsZP8VAk+jGvDuzZPzL6VRzp3UB8o7MsYW
ui47pmfSJBodZaBid0YChF7qoArmlM3SqxyGQJR8+WX+y6pT1xQAtxLnw/m96xQKBgZaAi+kJn+R
Zz/WzZKMwM+Q5pVKWeeMcL+LVcABRVk5U8B+COQo1+A5jyUAaSodaIn0bAZ5MpYnuvOVH+KkSCLf
SICaCjOQ51nPZ44Q50nSgZTOR7SlMBzuyB9/CRm5p9okvcGx87qNp/laT/AyMvVbUwma9DYL/l/e
loMFAdwbnh0aj/HZx6jUXss+EAAW4adtGrsoo/txemGid1SlUBk0S6sdUL3ugwBIaY91vbrSeTEf
x5R81jUM/lqt1Akbrtd0iE9jVqLI7hXfDHR3lMju14rlyYDZjS3SIzF2A6QiHPCGaX5bu8touh0z
jSWRsCekBxWJxEOqbJdrzusblqOJBHqli2EdepvHlSW2eHNvumebI2CsOl9Xtq5Yw39K2OFqrKYf
p188xzhNHLc0B1PtzUfrxK2iUST20mIERMxADUR8dOTOB2/itbAda7QCm1vduH4xNvhNSzfJ7K1p
aXFQ3/ez+pV36T6ZtKSYnQiiKtuKei0Ii7BS+um+hHw1YrnzKGwLgEyP+A8HwTeksOJ50nGTgMu2
piOR50miUvnswnvB8Sv5MA4cfh+FJVOg6rIRh+KF1feheAFXuxUWHBkdTU93qOWiP3PFe0ZmiL+7
wUVzQHPOvBLn2wE3JmKKK5s5cmDIjY2WAfFoHCSHfj05tMC7ewRJDcRDhWUfJQLrzQOBZNFrNeQ6
4QVjmw232El1vT8+KhUnPQnzmCKYtF7871mNycDOAspQOv5tRor8ssQIrAHN4dMXgeOYszC5wB/i
mjJzqEohShE/iSwFNJejotYk5jxXXgpTgcs0mkcFMxt+qQhEu5uwvXdDRYK+GPURMb40xR08VJMq
EAdalbDid8/c/EBeajW+6KbZrF1jnUjrO1DBzExRXPyscOa40fd8eZBBN0tNqNmvECJWPPdUrcnQ
AVpA+2wCALnUfO4slv+kPaJjqzkoxmlWU9U4vREPh0tZB13nIpe/ah5V3zhzvs8B/fKChr5b3vOW
ot0Le1FySYFskNf0naxvHCXZ0DAqT2cel5KhUws/N9ArKO4PCqyIKhv3vZb6+GuM4MbwylmU5KpF
okByTDp8zVOUO/XQHQHddVTbaLx4f8d0PHxJZUhLIaZOVMm4y3ql9rYfVkm7esytqujjpoHU9EAI
6+Ugrlh97i/fpWcrWwjHWHK36ijSX8nMTeP+7e6GohaBd6TdUGDg6Vfh2AEO+i/wsjq9dshn1SLH
4+VcAWr+K7/6tAv7wLKmCBmUrL6Z1jwinTVviwpMlStzU7kiTtoirvKDCkZFPlBi+nf/45+B9ora
lkbiYLHwz73tXVoOr2Ok2H2yFP/FuRo7GPIF+Nzf8LRmLFanWo751VfQVNUb4dA7uRWygqk6rq7U
eHuXagaNzFJRrWu56scZksoYWaXHUHzKvYPdoAyZs/0egd8crib25/Rt2UsBAUbcNAx8cDsQODfO
lz9I80vHDlRYwWSVK0jJD1Bv6Okui3NsRdsY1MOvIu0/wM8PHoAJunpwWeWtS9+3ktW2B0eyEEuP
gVtT1ea+DCAPXRzpDXi8DTIKLo2nM1722e4Mf6mi7VYi6O5gOke3fqau7L47VEu8EuDEoeJ9U1aq
cs8nYcAm7Y7cyA5w3F73I+M7bbaJpBOLean1x4o8N6hSCTz7bIFcCOhy3j4mZQsDP5CLtIjEIEPS
90yrfa0XlRvoxa/59mtoSHYhDxYe6PNyY2jBVJigQ9+oXwdem+f3kuKYgDxTPhTiAByOI/GJJPVl
NBo7rOLkDBlYfj1fCC6IsST8Iyh4JOlxIf+NE5zCJ/srGKu9jKndmI6Rq+B0Kq31a+AHY0GapHzD
d+5RMUZVmV7a0rKxxy/stOQVRr5fHCX0nqunrxvsr3v+6EKDC/qCsDiSXC3H+Ub+NaA8qRhYjZvA
fql2FcGnN0LFRXT1QGLda7wIOgPu0XQJViXVkJP9g6Ogg7H8d21vOIvqyzeiKdLxz6CikXNs+S1T
1ugxgq0PSGf/EVJDHlcJPsR1QQzhYzpPaVQyeHV8oZ1U5XdTyr8NQkkrpgi+EdfuMW1RFAKXw+fn
5EUTESaRLlNFEhtypGESS7ZpeV1a+QFpRXA385BMrP3jNeXYzDEvh0wPZFXuqO2qZSOSAv6g2uqU
TcQltplU6A7zZewz+kJdK+Bk7iHbWzMwexDt1kE4iw6TDLKlCDwOHk5IPB0TPIByM0xIUWLiDnKz
6v5xUgbo+errVtQeln8LLl1Gl+4STEbRLAcbWf8nWJ8LpzreCEx19Ah7Se0zdGkk0FMDFsvk6hVS
ypjj1ytIbhIw2UqHF7Z5HJrKzpYsCLNom0N0DJruF+ks3Gsazo3hLdwIAK/EeaVzQCU28YII0qsY
Fvc4MtEm9K1vRlqtf2AXeuzZE3N7YudlUgtU/U8Gihd4nFP7gq+wFxshK0l0Xv7EYGmjlUKMtK6L
awMQMXtdi2dyF6yqwK5k1hnBlfD/szRGUZqAs9UfarS9W7iLKGrgAfvje8N0MvAWt6z/CMdD7nVT
BVo8mgYiRhUYvCcfjW63C0fQw7lOdwmv6qYZUxB6AKgdPIu9rLuFcwZc5CoZaiHKsDQN0Yq+g0jA
ZuC+hACC7lM7g4bzAeqYCKLh7YLELC+x+CMcYbb0dNS56Vsw/dL1WvHxZaVw/avrm7GJgOhbrm6q
A1nzTpsoEtOmb/kq3kHGlamGiHu/V9kiUtmhrmTDfYeEdZBoh7REgXOAMEupKTR2Q8BhYSYBFntu
vw8igeFWHFNfXQRHe9jrTtmJUYQOOJYC9NcmipkmcRDDQpfDcFfTVpZvfW9PMm7xQLJ9lDlueNJL
G/YmC/TJAS+j8lRP7wgVaTvohURHvN7idAY7m6JyFqCTTK1GwlgwNScYBfJH1SnBE3BryWLBxwpG
4kysRd5B6zxvjFNwE/IXmopJD4Jfy8SGId95Orv9CO1I+654ihpdBZHHNz/qYa97dAfYaBQM/Q26
7qVpdP34/Yqt5hc9ZpgcWKpeujErYTL/DtdTEpM8YDDNknle+UtZqwO0B5ROa3zzk3+uxp40JVkw
zcrxeJxmRDHZGqBLYL6rmMw/6YJzRz0IuYsw8suQkmk0OCh6hfI3rjY38yrUBNll+gfJovVIWjOH
os6hhhJmVOcQAgzlgo/o7rK/vxia8zcVmboxF/gCKNU/Lkbi8FQI6zugq2V25oh1gpkOxShG1DzI
v3UGxLZfoSzxwrFW6wCs/SAzFNsDtYEacayIT5rGB3nPAiEKMjhmJ/zuFHXPI8HiasiHEoqaBsq2
63ou/IwZxW3F/Kv/hmqPGU5qzDpmk9zlUAP3RKYoC6djSZ/0rw0SILrYJ2u9SS4o4roiCU8Kpw16
m4HbBR67Vi5DbpHsJv7D96d8QGWv7phDbBUmGMURdKUGZmQ8RRE+jqyoo8Llj1iDlW4uAK9P1rhi
bVtqdKVLOyC09xW/H/KHHUpMfuDSd4c51sYYcYr020DknREzVZAg+TafMRSclvVOkXHlz1oIBWgQ
dsG7J+PWkA5KxsgwiynWZ2GYwb5LTTx1EzKnFizHKIWDJVN4n/9ahX2fyJSIiFLVp1bPWcjejXAI
ZSCzwUaBMqngt4G0jj06e8dxX/YVG0uFc5yF1pWEzMndO8PcEah2rDH/q8Qn6ZWKSgDVwoKnQ9Wh
LwEy2MaaO+FXM/6gjTYJuoLNejJtMSb5CWQWvY7fJ43VIcu2qNX24MczqeUpfLzCxBE9nJ4YXwAc
u0J1GwBozjiyEjzipBPNyf01a7bAi/8vXEvrRfWbJaLwTgOwAAaEDVUmGhSvmIPJUhGD/6cWcBj9
FMu+i/knSTGhV2Y/t+27M/6zgdIKFWUJVPKKgUu1dCHxbEYwPY98JiWUv6hfpZ9+vmL6AUZVPR4Y
RxaP+iHoKV7gS/bvIy6F7UcsKYerEKoLPlXJug/nrgOgLaPD2I41R7Y42Mjd0cQaLT24iHKNJioU
kV3IFSlZaAfSaWw4LAqEACgwcDrrJsY63HfzmZ+iaWfH3gyJS1kDtluShRkk4JxQBYik5V1+w4rZ
4SHpdrywmvAWLnUokfcvd6RyOwCaLXN6pF2lHX1hAvyfKRfIOty+g84dTn5d/AG0rOszq0y/v4XB
38adfrqxztx7bCHK+FQ9ymiv+Xs9f5YFI3MSA9bBhwqSnmV3F9LjrqT6YzwLj/wSyuOyvzzKt1Yn
ao4jX9+VnKLzbE2qL1uWRy4IenL8hfE8mC3TvOkbULvsLnxNDrUfyoWpXZq9AY5IG3l0HzFVUjVb
W1uOsQ0KCeGl3DXnsHiweFxIAma5anUpxbWUeu89lGVeJak2P4kVh5BjB2i9qZZeTRbq655OzyTF
LYGL2DnSjErfvDRyzUukAETS5YxI0IWEm6p9timupyu28pm9p1rPL7Het7ZmF5WK5watHriJvheo
O2WA/p/UvB8a4C5T2bhbGipMkc3ckPIb85Gj7jAkwrTHbdR4LFywo/nR4Y7kQnQivnF9dJTSXxBb
FLKlQsmcTJuhHwScNiZ2a5/axOMkh3wjCesvNJDDXRF2IIWB44PlFRjP8troQF97am27k1g6F6l6
vtJQjGc4yGKD5mtpeFi1NzAT9FwqkE9+CcOcU+8Qm+CbEwMmU1Ux8GEKjknAdukJ3cn9IZoQ/df7
m02DgS58fV3Rt8oi9WJn1n82MNKsl69TKkyN0L/uEqpljV/7f/ro0YZwAH56Xw6AzbJeL/DCfK7i
SPet0JnRcClm1uea70VEJFH0CLOu1iQsIwwmeVXkvcpGPnSLPtef00GPm7K9QktfTGn2zj1rwst5
Vq1AwSK9NZq9H5/K/vRzCQK/rJrtNzVtCywbM45Dk3jqi8z5QgX1jOWRKmMZnOxTXq5Y643we3YR
hTusJSunj11xoCwqjLOPLrzBzVoGNT4fK3KsHppMjyet2zCG1bN9AQYOxkR66AH1bNEAPuIrAb0P
o3aydi4EYQ3p0YZl0sWIbQb8MFCEhQHN2qLwvOwsqpXcLorBLPyPueb/50XRkm0Zi9fpwc8p/A0A
0QJUwBoisQiJfPC1Bfuv0kW9ehWjlL2L4ji+5AgqplUJP3IHl1cVrJMMAA4H2cxcfHtKqBN0Z4DV
1NFxKI5TsN1z73RuNm0g7D4sDWnoCD0F1uHzgWim2Y5zs+idtRCtlAJ7XkdYV75Bunpoi8sEkwpg
+wSKG1pqGOgqQAEzT9kcS8JpHXEM88/6yL9niAgSLo/tRQpDtDCKNzMk8DrueFUnphbT5x8+9EuY
N3r80pUgAEEPEYCLMSt5qqL8AwmtFgPdYBfJs4f8A96t1gbQjgP6GGEunnLE51w606ugZSIKBApm
Vrwtq5ppBY5tisHVPld+KU4nlvKbt9KwyVcqgOc2rGkH8vpwZLzbsKN8XxIxl4JVcPgL2dxmnbUI
O5cK5u/3W5Xv8VoBDkdtnPoBeLVT+Pcbcan58TqTyWZboCrQmKYx+ee4SjEQpHE6d3MT+alvNRb3
FHFPAImmMXYc71YeeWcgqEEMDQ/0VNe/lmZFDHDuL1dnbLaL3BFVtVKkQTGmfl0j/prO4qk5DPBO
S7iZ4dmNE4xXqwTWII4jIYPKND4nPdZbP2Xn9HnUdazZYFWMvY6QYupPCbZfToP5tMx0wVlC+TCv
EN3xo5CK//oOvvFGIEefR+OqMyGxZZIPJcztn7nyotxLOHanVR2c3U8UcefOY+SjCj6EaXBv390r
nv4zWvRtkxG7dwluY0m+ktb3KW3Q4ux02IdLxCN0DA4eZraGK35UyNlQVdHHEB7HbOYSPtPhCVjm
Ml0rkoRxvbFF2jgeGmIHmaF8u5sW4+cwfAempT5bVE0h8hXQdQHt6yC9WPdntS4JKxQ3VNvaWrGZ
lhcOW95pPw13G+nda2J7a2GL9cB/le9oGCxjY+QsLFiDQcYq50GPZ+GhVQdoJdh2WfyKlZTUcA/7
HEIxYfi+hlsiKH2ys07eFK1sZdd81CfVd5tZbb3dXXW9tHzcio6+O96X8dzck4kxuLBXU4Bf+uaC
Et9fYn0tA/DhDuEVXxPRHK8yzmXgJg4AssBRiTG8q0Z5Psuqc6MjDdm6OPSSu0c6ZdT0L+va+6UX
yeWPSaP1sosu1Hv2IOPuI74Yjvy87aae72Sf8jopF9O/3bNd9pOSEAny0yKMqLpjmFW0eNqL8CcD
BJ7nuG7ruUP6nqQBudf+dTcsh9X7v/YG3pUEyNJ4697bLi7U/tqRWfb87RyBjVADReRYEGjbqYKp
kLDz6WpCl913i8LnCL5kivyRxvOlLKa8yx37LLsE3QzWgQ3n/CVaCTH1bs78rvonopesjtrYfuzf
bIyzTjgLjJaBIozJBPqI6EOcJqRf6EsNjf9usW7Pqwsesxb4U2njlx5rsQy1uoFAhAc1ZXrJM4c4
whKZItKdWzGWb10dSnryTom9ql7WbjONUrDMzNkNL8GZgSlES7EzQZSIEEBp7Orj+kA08Q56xxUl
FzKaTU2ARFvfaGwROnivca8UOxCmCS3bY6cLyqpI39++wKXRc7EVb/RhPgh8PMcXtI3s8stnehXn
B4gifJlKDqYwJp/019upHEIzQcaqdxsyUbnhSTGAvZd6NEfCAd6jBdQ+7c8ZXjj9JTNc+15pi+4y
gXqh0sb+0bSI6VsPQ2TziEvV/QrFBbECqHXe14ydNu7whtLRRGk8nQi5o/nUijTbEpc/CAIP0KZq
2WFg9CyeIIrLDeSbztxfMr3UFHXdsuvxGooJrez5OZJsiWO1WzXMZRwhzZvPbGZBTdj/0KRNlM2Z
KRWZRkJLSTrYdEojr2xMUVQlpwEuqt7BbdF0i95FQSRsP5VVJOyVaWFtucWGG9YYlcVcGHoCV1wM
B1liSa1Pao3mc6qn2YWkMNk1ND3Kr1dfvrlquexTzEVmdHhmE9Yok4r6m1dPTH8kcvHG44efLTdO
F993B8Nvp+rXkeZNFeBYyQbYjqMImqyIj7m+DFKppSuzcdM8X7wl7RV2UnR59cAldETjFkgsVeMD
JacIlvUiAfQ4mPZv2iZDF7H0IHrbIgjkHeRTN5xZUdyePxuZwCeo7wPnlKIrdQBbvdNrQfqFF83W
Wt09R43Vkt4c9pym58OX68aWgkxA7eAnc51AWdifooUufP6KlL9TO0oUl/jUk5Ll9+qOqEi/HLyQ
a4hXxzi/w5bAvW57MgUXXNaINTXhTSdwYKmQxTHzieWWPcSsmb+BBwrKNb9wJUIeigNTvkbQc/xj
nyoDGxAZo/uunx/5dWLx08POlmxFRc0Ep2B5HV6rSzq+sm3xDw1Mg++FzJJA/WJUvBTV5zj9Tr2z
JnjwTNbLCYq673/bjtaJRpwBZTOpev5P30TtPnbHDWQ7TvMHGggDk3TLAAzmjcVGDaUNJSUml95d
L05LmIFyJ4x1nteZYaMBaGZUFsPuQ3EAu9CsZDP3xNFTOIOf/QCk/FqCsj3+p4rkB+FZbWxKYiD0
0yjpnbthr7C9A+o0Jr2hDNtNRM5+6IwY/ToyYm85Bp3gvY+4Zl41DIRZYuY2SToMsUj6LUpZeYVi
L7w1d5kYNrlCPnjIepXPfRiz4YPBxmgZDDkjINPrO9KJQhAnjUGP5u/7EZIaLORjFobosmGVVBBx
faypm69icIK7JO00/kn4r48pGirp/1Mj2pZaQpYjHyY6x7ZyEbaIJ8o/RRlZg21CZk4bHw6NGNvL
PxuAw+20YtRg3OnA2kLLDZArwwY1H32Ke5EdeMxRb12WGQjOliXnobQg8qhChYNqAG5R2y9PQIn3
dwLi3oopI5tE5BF7S/g8qon1k9x2gzi4ZHc3IEgijfSJmj7Ogav8FzqM1gGweaF8e2c7kp3TEIpy
j3hnAHryLRJPp8nlbUGO5z4dP27Yn3Rs70w03C6L7cCmM1CAIdhhNn6Fgs1ofST3W5MKaBXBYXYe
XON3RAdulp60lHXYBRr9nUXJjmQcJH0VSee+aKllcyPF1nk3EditAik98gdcKr+8E4JI+vHdKkND
mL4QenPjV6mKrj/S7omZm9eDGe3o1ZK9dyObiHsWOnL9hUgAcpmcyKNgjJPuML2/jworXM8o8s79
CbJuLc1ja26On405DkV2aAi1I9l4tosgyN2RNHolXxcNjVhbsyKR6/46cZbdQmlCzqp9Vhk7OmnK
Pgi/w/5Jyo7E+ErqSLuIuU342V17Vn6lR45xMCLq9tuZgRo4UhA2Mueb4qE8VAq+AHsPXhGQ9lhx
zh/DcAsP25VeVilR3Ax+attGG6v+GOG4PPsSXjYpt2DXngQb/XFl4ywIKivXUk8AcPAdj3kNvBEI
svHmda8DghWLh01TOU209VHmF9cC99HQGMfD4wmrZKh7IqeDCrome0VfAFddRSbnnPX473p7m6rD
Ik4Zt5co7loHltTrdEQjpLTLE3ylZrerujUrW13bx9yZRnSrtvzPsZziDUX5rKSBp7TmyYMtsXe+
iL3kKom8sHVfkNS6gqytctiOD8owPacvp/BLuHqtpHjz+fAtEl4xCNQdkOvTje0rmC2sobVbLHFr
5QsE6KG8Q81gc+hMP1hzEAVzvtvnOuWnNbVmfhOHKK7eX0O3mBop2KzeRcw+Lbcsenm1cTu356ZF
I8eDF/p+OBy3B4zSUTJoBNzvZKl7og46DpQA+MYJCQq80bXRhjpaGlmRc4sg4ZSeaHE/lU6Zmf/m
5H5EmZbNOC3rezOfIRGNyf5wEPpniJ2EngEOl8maUIQnPbSL1xXvIzBM6OK1WtvOlAZuDxO/KwUz
3LHmeO8mEvlu0AmHtwakvXyEUocDJWFJf2S7dO6hLqUiKi/8QXX11EFTq0LZXYzVInfTE8SbudqU
OB9hlZlnmnuWU/spKu8j7zoMQn5w7p784Yowc20alR7AsuoIVLV14XJ93czYkZji0QrVpTOaWp4D
9b8M7cEje4F4AIu5shYlI2Ds0Ga9kflSQdWk7BoaHoRW606u+312/A3AGqJFkvjiUcgJN3cZtQgD
rMt8CKFsfL34fWnwAvWlmPfnWuQrr69k5jW/PyBIYF5glz9jwr25+uMpOsPHZYIK1eX53dRTRlVh
x5aiCMx52ho/OcT/zC0zPVgEtuQZN4Ij7LM8sM4bnEKcmlKcj328O4+xWXdngpkyAIPcEnydQ0va
KHgN2e1AXAmxr+MD74HpcdiGbfi869kz5P+hFE3nrlpA4aVofJm8GVvRqgtbilQZSJhp6KDYVzF0
x1/x1BAYWVCTCPUEnUCnQ6A8eMeVOx1w8W66QC7+3nd0LonSbGc6pC2nFxIH1ahrjmncBDA1M7Ds
iIrsuogex+jJsOQQyIF9nqxDlBba6yj0/FtJLpf4O+8VWXhQ1YHA0PAUgHCATOmTn+vSojhRdz7F
p7EGPpCqIT/QueAorFKtL8+Pq62gBcoIXVbP7qLSkcBxB2gWiBhKnBWCORlCVLqm3jdsUiiQJiYY
flzawFhVqiY/zyBoJNtgiqlxNaTL5mFB1oe0X832ZBjdxCzY+Pb5UFhM8KGwRrg25hqVCTnsCo0G
r/C3mZMinq6R+jz3MJ3iSKYegpMgVCTHDPeOcsN8UwsEeZOaYoVz/x8SAZ578hmiHo0gggscy17F
ysSXG7dMatJJ87M/vBr0g9eqmFvRymeXLkG+NC6T26n0W8FRb8mobsQPfAqgp2MsUxQSphCOpOxU
PXqZP0ANSLQXeN3D8kg2ujQN+zjbFq2nd1LW4+u6+pVM4DdKSIx5V37yw7GsBBeJkQVmLXLLy2p/
OhpRZlxRx3eTzoGytSxJ9c7+i/ECaxbY0vq/UUzr3xndZbYN3h+1UKwsW+zYNEdJLravEvwclnNh
rum6w2MseVhBe9TMeb+9zsW8n3PvTromZFdrskgmuCoV79RVU3xF06i5gYwN3fp0zNY5/DJgEPwt
Pfts57JiwdV83YgY/UMMMaJkf+OJ76OHGT4X3jYpPO4FD0lZ99tgef29V3E57+Fb8f6kNtL6H4Dh
fmrdh3bagWzrFN7iXPr+Yw4tO+9tJTq9NZx0pGtUqsepAjWjXB/Au1xtQil/F79kYoGmHYAviVMm
OdnBMi05t17axG5YwBNEP05IvDivndAd0wRRM8kFZkLxZKGbLWf2oA44UIgHL3cHYQ17ooidUpeR
I8ttgg74WPuGp9OP1dUIVCE4vNG9AGac35340hOjYL0oy+XKJtzLZ2uCnvUsD50b8Kp3VP+qakHN
ReMi/Hctl++giTMHnyToTwiGx76cnBde1DiS2ubRXT3RVqOuR/v6rWu8mzxLDAoAjSqKUR4R2u9Q
WQv0fbe8bQN49rA3Q1o88sroD0GpOwz3jWPaqTI0Ry/0AG6SpwAyuoueVWQjbl29NTNSy/vz4STH
M52kxpuCUYKQpZuqu7oQq86rfI4cCeKGRvNOepj3f7Ggxp2/lDe+TThnJa7syO0IYVyXCEiR1Hwj
1/hz6SgcBuxIwT0qMCwJQraQYN666H4bCfUttlSTuLsEu2EUk/xTfC15Q21VwHyQcxZ/dUrgFaAv
Kc14ChFar7w/tRj0h0Telw+4k1Vhg0GWBBxoeWUstPfN8tPQ+9M3Iv8+NnmhQyXQPiMcS1Oj0qxW
EYRRfAOVQ2sP+WVbgEAjRbHWKSKJDB5P8uCVjJP4dqYxhsDdOnY/ApyZKXB8Z6uHns6+QdG4HaEU
JbEjFUTHw23tB+tjU2U62hX6Kh/zc4MgURsLLBhOScA7BXGBEwwZItjoiR6E5THTvuUpU5oSLydV
8aa7CgCJITdURZIQDjC069FTbgRz9YMcCw5Pzl3sW2Ol5naCRgvN67L/DHqx68k0Xg/CWaN5mr5W
/UOSJDb1GIMIuxI0qfYql388f1RxXo3xeDUz2xUdjsDmCvvGM5x0y7+ryLFEzpWlxwUFsGV+mwd9
/KO/H+wwLflG5Ezmokq3kDncBmTHje/2DoLam21HERr1tjugE2C+mNlC4c8LwmmZO2wM4Mc+rdQA
9V1qrtPYLlZ0pFRzKqHotOkSfgAVxvkjQy3hdhrwHd1Y+/ouSB7u7sov3kC0MFNjCEMmdFBGh7XY
kmUA+93qxKY5iPMjtwbBBm1jq8dq19pUGnwjH8tE24OcTgy2mk+xuS7boolFROS/Eor/G5JrMp9W
6cluC7GQDOosaXvft1kRKtFmmXRRBN07f13P2A0xL9xeKYKOIaKkuPmfe+q2SxysKpHbJcbTExY+
JQbi9owK+M/BCDiJf3JmQOe7U8EOBCpvRYXmF2CxZyU3mmHNrgo3BPyWIoTZKm2hpQKtddK69ohb
b9FLUW/MBgUsyGOW6Vdlm7Vrrf94CDYneazHqMf6dIu4mmDxsd3cSsWTJnN2EFq+ZgfJ0Rf4BN6+
o6BHko1Urg6Jg8qbkmQnBLL1FZ0lkj+ewbvHIbbAXpumIdD+l4PDCpFJaA1b9pJTGVHUh9208ykd
5WYuNW+OxS65qNmn3laqz7IllzS2jRFKHeEBES2mkjzIpuv0IUr8T4hMbDzjv2djbxk2yIxW6rdE
35z+xM2pjB2NjwkVJ17+b410m71/GC7pZDFBVqhjhaIf+Wl7EIPPq3Eew+PlnTkkmBP5h/LWAM3K
TG5DvDLPyWmJlBcFa/xiPrI8x5B1yc0AuT4aRPn7h43X4WLha26F7erpAtH4MexKXs0jkbVM8PRM
zTEP6cuSZOgsCS1cCxaG6GZOoAcKShY6z4VmItzWy+GY0MFzj7g9p44LEE7tmFgEu8IQFb7mJkSa
+Fd1apDvWQ0MIeQnwhPdvL9bcgCRRVtcAVs2QcvLgQNt5kt/m+8MO6Ig4qv2EOxjbORo2zbHGAG3
dQsfrj0M1goLWYO0Qz8UpMPuzvjCYOCaVS7PfMDhZQz5CUeuuHsGG+lzryx/FNW6YI6oRbGl7GnC
KY8G65Uzv9/lUC9tV/Jtqajga5rX+B3gZ8JecnPPrsA+OABfJv5dgHsz1tpSAIDMl7XQP+xrork4
wrSPqAhAtlHItYJ+DIxmM5RERMS8gR2qkrFJAwcjZoNHmJJZNjcs/3nx0inG8mjOevRljVDyqb/P
gEf2W4m5aE0SCq6dWxnDiEBk+Rci04EM1aiGPNnaKPKyEn0LE4h9nocFWjzkIK7A6VeNI0RSmyw0
YlHbw0ly6WRy/j/luUI0ghVOdc9/20GDGI4qdg4MpFFKylN2XiUNyI1LxASaHpbUTUeWCoXu7D8O
x2PwfD98+/+an+c6A/PvS62fR9W8BBeL/sWvW5ZXKdieBWs4a3+Q2jTFb64ibm6Ay/aMsROSU9s+
1YQ3ZIF5n/vOc/18/6nph3Ut4AKxM9/Waw52dD13k+9Bm/bEJ23eom+TgCXlL0+tvP/zkx6ppCko
8Bj80pi6QXeNrsOjbU0aR9lS0aGEfxxAPVUAq7pQ4Qsh8OuSL83Ai5IcZQA6F+ugyh+pkjve7QGN
UwcJeybJzMTBW3PXxQ9KcZBw+QwoTsajRDz6cSwGdwUVhnoVgIHRnZkPpaNM52VcO7aGVGGqG726
uOnSUYLWUftZObGaQ7TxOVecZPPL6JITuRA7bU1zl0unlhUDvQ+IMdjkCmsiZK/LQf0pdT3CwNhY
H+rpBaMDBsx7wPonVo+I8mg2oWbYIs/ls5boMmFSp1dNu5SFILsEMYgdN9xY9YO2UpZxJzwddRG6
EuOWe0urdoj7jaMugMQlEJOuCsxcibitVhDwN81ASbp08CmqJDVAxstpt2KlK83BVwHfg16dFoAA
w/Kv7N/5mzbFHrgr8zwCvBcToK/uOWDeb4gPUsT8q/UcsFSuwCJ3mU6HoQZbBbj8pUdCUItwi6qy
SFPcZ2kfi19j/pvW6m6MD5g5Ap6npNeExL6kP+X0uZpY5q0+r+/GzNeAju7BaQSvxXBCY3JJTg1W
LjfAYnb3jqsfUgAno5AovkRkl9B0wphwAJuPy6hGd2hRvUp1lokevKL/zTh//TzJAy5XXxlRXsZe
8TQTliCvr3qec+68YoMZjUiILbWbM0YEmKAEGZ9+WXZMv6d7GE3iNZbd7mrcVt8V8ExsMQ5bZZEl
tFRSRG2tyoxDkF3YB1L0btyPI+wHm+ZqtiOg+G5n/kzAAFNo/yPuvCTiF64OFA9IOnhGNmeyS77/
ruQaOzn4M8nu/B6E0uDKJ5bFdB/+YWp1yeaXNud/24BmukeDVpmVjYDje2AgyanWRS6IavAdQprH
DCQ9/Y5X8VMLYej8LVEUziC7SXglXjYtjBYWG9WCMuWYuCtKXvFFhJ40xW5xzyEKXya8TGM7Flol
nTFUYJXXyNt3mO5y/4eqNG4aU3rRMvCAipyn96+yggYuOyewVFhIBuoJGUaHScDnRzjKRK816tXV
N9fry3IrBka+JuHhYlrtHAisO+T6sCEz1xRDDZG+rEkFxhCmuD8qL169JIdiq+FG/JNPNGoy6xr6
6y3T3Y3GUfMx7/QvQfEzWW7knsWZ12vOUN7+1z+c/n6v+Pqz5ZoMA/0cysS5ynjxzHfDcNDpg4xq
xv59IjNasADobeH/FA8SH6nOOXMvIFY/wKhBi4ZXUU6y8Xc2OYiVzII/yAT7jeCwG7g8jyaMHTDq
p9jDh/QLlfK/QKjTOjSo5k96J6NfzZ/5Rff4M5/0Pm8rf+MPNRuCiXmb4kIObeaPJJR2zhgMGmHs
hSSF19vNeLiQSPRljDqhnjoWER290X+xyfFTpMtYWcvAchmp8jWb1m+lrs8zJXxnTCGoonKcqHsv
XNNoJU3hQagLRK6lfWVEh78ujqtgu5ZclgShOXrbxziSkrfI+4f9J4jxjKYkaP2B/e0ETSZmGcUu
1tmyAWfwk9qtQJzC26NPA4GBkhRyN119wteSi/zForcGbD2d8gs2vncQEJiUBB49oc9ox6kjLNBe
h7vScEQNRLhZpFgdCrQ2n3Dm6YgiA2laH5Z2Q2Mc0BXd5+oAPL84xNUqEuIAj/4kXTL/KDSqiwvW
57Nskj2nauLYyX/UOV6TNeeQOOaihsHiBnrCLAnyjgSrw3JaNCcDVGXkGMBjwmTn2l+/dBKqCuYF
bB++nkiy0f4LmjhrXoWPe6dT4mWJRd/p9YFkt47qKJ93Lvp87juCUGaLoOH7oDRBjeYrAo+2Mo14
eu/yGWnwAazCWK3YIw1OB+UiuY05OdFH+u4hqYnf78kMsuEebUdvfYeY+u5VU2HXv51GintWL1WQ
RNifSVcosOQPe+QCCKUqG4w8Hfs8pnZndcML2XD7eRUIDqnKhg1CVDMdlJ+xUkuzSVdaY4uA+XSQ
RvjRBh9nXixpRmGlcvTDy4o4K6dRK3b1PgnWjJivK2Zp3UgtMl7TmXKc2lDgZDqrxRTyKHMH1sRP
oIJxg1pJk6NdXHiYv9BTvZXOLxrWijBA5x7N0bmAniOeIOkFRMbS1NB8xzGMwXeK48l0kUTSuyaj
x9kfaOef6E7oLM+7U9roqNbCTdJiWvLwHAJjSKtT/pVBWF1wm5SOO2YqY6u0sy5wd50+F3zONsn0
NoScHmgU5aeWxVJ2J4cRsV7l7+KhORnSlttHloEu05thBqmS49kX2HTtoEOdUFPz11KJ4awoNPwu
yIhAMfKVI4KSCDV/YNDBdPAuO1TtCRSBFJHFulF428NpTI991mB82zU/9lw/AVsBcNRD/SBNMsrg
IebvHkb9O2lz8gO7JlIqBF8RG59Ml8MUNjSCEH6yzQSmh7eZADazrlZ5woUL+82qWwLdSQumzqin
eaXkXl8+BV7mJrRnysHL0uOIRhWuhBlHkHLJY0jnQLsgKaPEalJpQZPKheX1wcPGqoBifnDE1Zif
JugR5sTQ7kL43eseq3/kuKHKhrrlpVKkaRAGfk2Jdl96QpBZ1l55IzsGAQx3nFt2Ieew+h5UI0eo
E+adwQ+Gfjpxq+/5JrPDgSP8cGPj2dZ7DOwy/6x/Tfu6uN3uE3cUP7Caw9wAglRu0jNNUGssUT5J
qaBl80iVjV9DJIUVWz7bKcpqrWqI0oE193RJ4WeF5M+7dVWIaASWbi37Ei/nN1jyCD2x+AEeZtnY
byfL/JEXzwoqoVjtahIYknshcAoS/2MV0uwbZv2929AcBNiHVIR1vFqjN1MW949z+gdr+BgcPj/N
rxjySUHyYoGNQR80LgJ+NzOuB4tU0bbRXqO4xLj1IIwYYbCQ8ET3Ox1U68rPNdqfntLGOSqP5rtk
bDYO1KveSxW7EASAaPXI3Y86kACRI1Bmgvs05ETAoPFlVGC18DgKbwK+4XPyLD+Vnu3SXhfvZYP8
5AVVflyr442YNCvaZNJ0j4r1OPESG4ymmg1Y7MBEjUkYjLQuqxi4CHK7KLaFEKOMkaDmrYJMv4JS
GtH/j2nmGaHsPmXpTu0VzZtBauGbJTZz0zX8I6FFs/DwrPUZcwWkoGnSTfrRF4HcfSMpSF3qzQS0
JBDr6Kk9f0TNWBdEeFoeM47b2bNV0RyvgTo8UoS8nJuPKYWTVtQdLekJMHszqCuAv5yyBBXpTKSh
cT/vVCi8LWB4Ei68x6K2Jo0//ERJrNPuDiXPVNwEaJtbFcYP/DEanRbGG2T7iR0A0r0jPFbiTulD
wMEVH7YbNVu1XuzP5SmtAcJz6dVx7Gf4zcgp/uNr/TEzOOHI8G6bsmPAe0py5Fc4GUt7VZB8jyUI
Kp8DmxLLL0r7uhyqpruAZmr8ZynDZe0P92qDDvUB7C5y5XR39ssCtpEHUM6yvxDIQWfQMoz7r7jx
ScB4R8fSKAiNk/GjWggGQVJXYj64b50URQ6SDh6h1wQXH/3jA7RyG1Zk3WsGA98XFjdySILslDFA
I3U48XA0kDY8w3g4a61FfRAwB5Xe78T+dcrH9Q1+stjUh8KyNsOVHuSvk/4QP2w+0cidQQwDQQhk
LDUSJFjzsfpTVmBYYezIgeGqloAiMLXY1SAiiu34ppHp0EgoAZ96twxrECVza2hqMQqrtwz14XFB
ggNWSDk1RbfNjly0waKnCtHSZ3ymVG+ivQXs7mWv8YZ/uOqnNhtSKBktAR4N9mARcxsB8GNxPpo1
sHqC1bm2m0GDgHjL2XV2zkIF0fm+rkbRRibcMVz6oSbFrBK6bWQ4Na/UwufyrSOReI+Ef197m8sF
TcP3hsz5XXUdZvzi1y31cwGc2Rm070zbCt5HWZuVxxAloBgr9TRH3aJjqL/CgR/XddthBgDDxKUH
P7ksHRJY3nMvB4cLD22Q/Z9p6/dMnL9y8z8dugpbjKCje/Y6P29MhLwZHaT8p6b0nYT0vZfFwYVp
M6Wu1uqz4U9210XZEIEEWTLrXILgzVX3+GQkR+GVUxFVv9hkw5bEg2bdF+pTA7hFxw/b7Fwy+Mhm
BhYTlXA4+nooW+wnNKgFctP9EuD7j1++zy/Jw/wwWXdSyXL6faH8zTQoRpqjRw2yjgJaDDprh0Vu
EX/+HjIQlIvLkMqLAFwwwVoB3Vr/UrV+Lvt/nyfHgBE2mCleqX6MkQ6WIdsnaddQxzkNbfbxI6Ea
M/JEpta0OkR12c5Dhkn+SIh3iyRxoMApy5j3hdaqxENeIFiLB6zEcOMQ7QHx5VxHvxyd9/AmDXhP
aNJwnwBAy/1FLM9AnRraL1yFCpImZhnp6/hs6duZNWQDPQK1+175M2Qw6Xc1xvUWlfXgyVYfZInR
bydtYceDqjvP0zO3OP/Io4wwnhGzITlin8MbXdzIo1mboRJQUMFVrDvYqj1ih6ml9XT8ALwJc5WT
27AyNR3kDRkazBPFDDSw5S6N+nAAEWwP3VlCTIqONdnp1qpAsIKdRKBWm58LPZuEuKYSWXdMYPCC
/F2yewhm5aXOtmd/1pm9QDL8zyeNAI13zTMXgHWHQ+3pe0JBb9aMniY2eGejLWxeYYwXzx4T/X0F
i6eEGu8kHVJN3fpN9vVrsHnBK26ebjdPD+gh8EwgrE2nEKOjkog4CaN4HYQykAIDWaiJyP0epBsw
0IqiAetcaOHqudRhFwbqhVZUl9l0GL10Yk1+Yr3xyorUyPxn/FHKg2Uund06AFILyFVeyI5kQ304
v5FNP5KBPqY2zZiLuu2CBZsTypObZqJdAqy2vV78t6ZKbeUgmXm8dp4TcLumS6SCkhSsEoO2+8nZ
+SPPDtC3AFKqgWB549PcfWn9LWGrxRsErLjhTYTcdv9IJoAHqfCupfw4BzdmCPo2Rhj8lcsUcooo
1olsjnRnMjw5Aq5E/2xOjA97zFXX5jYSNrxisFaRPUJuOu7wVcmVoW90LszvzRtN7jHFXEIh07pB
RVzyiFE8BId7TIJcgNOP9IaP5jvwq6GijVd1q5g9xXUMIKxfvoi1jf48jJu1Z4RVdea7EdiIPHh/
Lkosfh1Dx8ROVj0qP6+8C62tVbftL2ZwTRk7vPNMDjz2APtUvxIjqjj1CNfMLLaSnnULetONq9eB
UIxYkpsH3icVONyDFaZEGgHrMRzDHvINtitRSHZ7nDdoxDhMHfhor1iC07YgBqDdI0ga+0CNh5V4
Vh/ds9ThBCwPDr1ucveliWwMqbujsf7Rfai2XUvcKm1pAXbMc1/xVslX+zao5CEQEYPZVGn8/5mr
BLxMTMgK4SSihivofNu1XO3o+TqrUeCs0XUFbGTtMS/MrgjOGuAH2VsxJ7vh3Mqv4ysewX7hlDPl
fG6uxX6SYXJiQuRK8jJtBMlkbs84njNqX/Bs8U0lWgVJYm89NuqPdR12/Fo0MWznRbNgzRR4b7Gm
+lvTYFpjxSgv/KRRcbOLz66u8XelHg7krxYj0V7MOj5cgkaMvMoELhMx40nb/KKQ4BUkxi+5lLzB
99VICGTprPGHPxILz2x7x2JBG2qjN1WCN7zhAOBk2UMwSD8HRMbp0d1MHzopB1uwrzhkB/xl9a5T
A7EFgKBzulKG8F28gVN242/DmH9Xd5i6zvU5TWzUQRXhaDfrp/gvamdQqjigTF6wviqkXny3yjPS
h7rvWxwBo8uPHOQiwDvChLtysACmOplg9hew2dJjC40GItTJ2itsj6q8Nrw/z5tbqJqtryw5o3YX
OxKxgCtMlNOXkbfrtXsia9BZv8CBNto3X5VfzmOwgCxTREQLHsDsdQIbGNWqAJJX4/D1Fe2VaPEX
sDtifZ8Ut6OOI6oWCCf1qXQVEGg/3JYhKKDe8d7FNsN1AH0xEx18RAL2/emQIhahWdBC1/bHPVMm
4AL42MarJJTOKjneXk5D4l538wkGUjpLH7yiEFd/j7Uipy3S65WrF4vW6+PRrp3AlLU/IWCXkD3y
teTC8pL42KUD4TwnztYTp3aaAORoQQM8MYuWwrRciMI6l6wCdqER7GmwpV6H3zrry1H576xIH85J
t3MtlIyQNT9LaeAa5AOctortU2DlBUoBP+dqdvcginerj0Md87Z8mhvFK6GVhxe+81HRipUmZOt4
o8n6mtbe/PeUoqjD0i9/+unIe6PRk+8DUbIfYYf6gKrHXKWtjKr2AN/E8Dzv0nNFn9RrNCTHZSvD
1jrVUnn0PtwX+PjgTlkePfS09sCQrzGjfP3jxltTvcUZoLVrxIWumIytxM6LzLxpe2NfLd0H284P
Jl1BfPorNA1J4KH85xR1X4DD1WyzNtLHBNWJk7Muvu2iN0DK8UnIyBhZV4EpCwGzX/YIqlFQPOi1
nOVOnuj3VF7CxcPXe54iw1Gay86VRdoycss6lpl6xikiuSzcJFHCOd0O68GF/asedWTVTIkDyOS8
gtOIc7D04ZX1mxRyPZQSNuzetU4AlcgtR3JuYNBgoYv9QJWtWQMmIzTFvlRBOmyLIxNgCIF/LYo7
6N3Y9GQ/9pQRBy6lZrpLk7Q42I4NPQhUctH3EzAgMmyLySX5uc5CDh05ODkelZ0PnRqilAwKFP5k
/IZgpUwf5m3a3vHlAZV5zaEMTctvJpWSyqExPzYUt1tW5FyVwvgkLIm4Sgp7/pAyuUcPoBxx/aM+
Idda3YxsoxLXHdqnMwXmtYR935jjgDjAgvlbRW6HrtVdYwrHdwRg3btso//hhz7Mm0GmtjZcOKxG
vaK4BQ4hp9n45yWE0gnmsmUGCISEGbkmAdlfhfhKmrSAkbbc52qRTs1n/vlzJx6RlvVrQf/rEZ5P
Q27bQYZVEI4GVxHRMrRB4AAF+JwNM1ujT14o7JoZnABN8oW9RlQJvUFf+K37CPvbo6CynPNKPSjw
cSx9LPNF/LBxg5VUxrhb1W7sUOnMNzwiJgRjCVjfzKePcfnbuu6Z2d5V/MW02x3fTTyaTnhMbwoN
1saDXp9bGgNm9GWmw+OSUd1IADS/wCHtdFZtVOPvCMLORBwDrDJjjPZW3hDcAlPaI0bNz0iEF0J6
+5HRYKKZcu96Oh1lUrPgx2rA5gqUuY+TiLXjQQ6K4TZ2Gsx7tTbr96uLy5tbUMf+Y7pZuTkOlHBo
6A25oLoqBLJInTtASKiWg1Rnvxf56lSCl1IyG/ob8p8C9mEZUEZstiUQio6cqMo2w2/7FaltdIXW
WjaTyWtrRFStwxhpx0f7g8QAVJuc3OFZAQxb7zTS1kJrHcOthZirDUV6lkyfFGR7LHvgLodRYhuI
UHJ6WYbLsDkVBDCHLRwcZDIyQ9oW37Whk9QSK4A+VMcRmvnbqKnIYjykOBDzx91kL36uYAoOuoAK
Q3z4j/GFv4sDtj4z9VFeD79DtFne9Lm9KGPAjBNSO0+XRHpwFuP9UqBzBwFGLVpZnQJvKt/MG43T
th/HQoIN7DmBv9rIV0hCvmXpddT3WuDrSPb10+onX1N+mcBfcpBYZwLBT4D7xwjS8FI5nNVhBn6N
My/wM5HDsuRJ9AJ5+TGvVyMGz6S3d+F/EY7OPQvEBqsMVZuc4jdI4ZyjNv5Gl5pS1iFUCXat3udy
ozPFP6C3HN7hAY6MhcFOVBPMrbixlRUo+sEWyazoHa3H+R3UnE3hE1ILH7gT2us5ZAobFNp5ybm9
MPNldaMDRNzw6YPiV5BsetixR9R0+kDpxs176SJ2vGNYwOHDyqKDSGZ0WDakmA6o+VkYqqaCOEf7
xM9ozMExT6iD1zWXdqb4yFzMyk6cMldVAzOFAufeP48IFVQV/t2yMOZcZAsuXPYY/ZD/cQ9cjtyg
Yo2Qu51PhIR/PdwxwxkxRmKP4JWXp/P08kmYf0FoGMGwIRM92BztkPSd3246j3s3Jaj29NfSxMWl
d4vRTG8p95DEcoYkN7p5m9mGcEgw2YUGQOmFdPHJxcb46WLb7x7k9NbOCsgPGkbbvCkgAOsnkM17
Huxhl5Cn5aSoNAN5U3WkO+pykaC1ajk4oerE9MxUn5surEO1XZ6+yig5Tx0L5ujkPPSM4uKi6jXg
XaW6W9ZYXrDfQUTsJ3q3JeOVhhVWldj8I/CX+WXstk7EWYKoyxTa++gLH2Ccy/rmr2bJpPLvcROe
1gVKRm9UCEJV1aHEhEEMZajxVX9iJ7bfDKfVnd4Oa0FeAtjElX9ucvbuXuWL3OXMvK6HEAGgi/6/
WWtyg82tk/nw0TNg1CTMPIolEtf5XwjC9bKG025wkfvhk8iuhmaRDAFJ+iVCS2LlajH3uTQ+nmE3
i/7tdC1cF5T6brCm8fTxcQCmlrigf/YX4OBop0RGBhKWnnq2kpz9UBdL8odVLU81FQd5qfBO9xCW
RABmSW8S799g3/MuNWSb/YSZQP9Em2C+rZ3JfevaUy3OH1sXxFdfPfSU4mGauEqeRKgudvj//LBD
HtipVtRTVB6KKVox/vOLgYEu/RNqTqwAkMlRw8NKVhT0zvtK6VBb1TrQDaZ90Dh7laf7H9wV7jdY
hM7BD40i0J+gNVwg4hFvF0B1ceHxDBBju5D1RBU6uZsGXkzTzSnqNU6EhHFVTUulstzRKckN7PTn
QNwONd6BGw5xU32dPnS90rhw4IDbP7pM+6NWdxdYvhUEW9DqD3lM3P11zqnDLE+rkJo5YQPgBGlc
pTT0qcqehmgBOgLVwXpf8aoYBZUnzGKJT1UxeE5b0olvS0YCf9sY0Nv17h9obJrxRMw1bAGDyw7z
yjpZiQ1nvY5VppZWjVAAv66D5duwc+LvQ3RNrCNvr6KaSCNQVEE/WIdxUJp2pjSyxOW53uubp5+O
HEEwUfojxnGpKenNDbfTS15nRwr/lZlFmggatX96bm4IwRVVixKO5Sdr6gtGC/xX5I5GghzR67N4
+Gox83s/mMZJs7ol4aptHfDT2wO4uFQ2mbsJAnxdxjLb1YU5pSd0GZkCHdz+HaTweqIxu2Q0OUQ2
Cs+xLSlOzEFFdZzoHbPrNHjF3httfCk/1vAJ5CpTpGqphyxrZ6it42p4zgmbAzoBfSdTdWhCnUG9
eHTiHf9einOysZTAWkNAivltGTRGVHJzCkmPxYGHuVnLOvDT1E1m0xpH1OF2OecobD5v63Da+SX2
zotK6laTybuUPHKWq8c5ikZkIRiE2GvNIHGEqbCTS8cadf9GFs89In37WTy7SnkxO6UJuNPYy0j4
UcC4alzhq5x+CiehjaaWGG98G4vV52UjekJblGCXgUq9vuDA+CaWp4TW0RzojZ5HIsuc6XzROk3O
wQR9Y4USsz3pi+GE4iRQ8uZOuE6VKflsvY+ZVdlMtlo1hz7wVgEk+b734jXLyH8Ipy16m9M/wr3e
IvF2FnXUVbNANwBz2B3Fza/cB+v9nYJApnUGxzU2b8u/jiSYilJrKXG44AZqIebFGtuSq3YYBzIR
aN8qEWlxm1ZzjiHh2PSrgWzTOihiJURq2JSZ/zicZNnjm+X8KDQG8uOx7J6bnXd4LkCs4ZaKsDjW
8RGyELFYUBbxINa2FiB/EVy7L6pAEOMqvQ8GZrPXIE8pX4NEF6bPQvZ583riLlaC0lntiJ9A6qnt
8CHjN1uOtdz5h9fdEXd32pP3AUw6Jgem0KkqSKL5cKmpDNSVIYz46cVvzXjyaUg3RJYwv5sGNDnI
x1sk5nSJitg0/0lz+xKW7/OAOW+4ZIljE9BGAvuyFX9fdjXx1OAZ2glPiGP9/wqh1F2tMUpf7blI
HWhs3jvZ6NPs7XshjB9rKEukedLLd47rvOEwtYsYYfp/ku56iCSgTpL5Ra/ij4HDao1y+4XFRk8h
p4iUlhPnfCi8m9ODTqLo7blX6bQAAnw7REo4dLUHi6lcmlTVO4HNG7wsvQ9T2XTHSsli5mad890D
8Q+sUMcIxQOmfN4BO6Gj2258URQmYiP8rpx4LGoytaCVdhXufVC+IDGQJz5jJBjOixZvN09bo19U
tsuN+Rk1N7yoVNbN1c1SVc5EMCEfFzhsHvSX4imrkcqKVKM89zjl2XsR+xe5wFFrxiHQS7voUpcx
x6VnfA2lOCkLJUllaXlNk+Ws13hFjlKu6jFpr3OdJJ//d5hhih1Helu3Gk0NwnzkqOQHCK6WYh3j
FtdxQ3HZioIc5Qvd4hcI2wUjM/NZU5ZmgzEMHXSZ8EU7pZhaTqwh5OQYtOWoCdKipc5x/8IClCLD
oAoQekQJuysja/sJjlaW0hNHxsZLtAsbNpYg1LaRKQCmQ17NmtAonjqioZ6GGsJx4ZkFMYUnNao3
YXZR0cDBMQxYvbFK20QYEXlOceVf4QzTm3R2OkBdCEffAAXfsSSt+LMHzicziJnHU7v7njFO7E2D
gJw3zIk2ONyOqsFR0tK32VNOi29XdKeLliI7FRx7MGHMXXbavjmlTDLzhulinjRwMCf7W773/YHS
CY+CH6D+RfkQGGq6Ac49/CZi+/bVNNFv+K1PNgrHkYN4qaEBT/E2a0qx+CS8UmuUmFOLEENrb5Wg
t3yGhGt4IgkYvydSPF5sYghQ69Cz050uCOHSaugcT9MqkqthzGj1AIVPubKDqJyXDghg7vZzCU44
yHWjAFd9zDwGKH7k2hdGGfMwhkWEZvm0m/vlbuVcECADtHT/aWVGaXgiGtA0GJ3sw7qEvRpZ+K/u
4uJalLn0IJTEXh6wDYTEU6dzk0kurQO6LttcHM6OjTZSio+jFefbngk5YwADAVaU1q9dUClrxMj/
bp98hm40KJjiUzyyoqqvyji0z54eBcysrxPOiyq0wY8M5Y0NQ5+FmLyC4KFF/smF5bUheaXPqzYn
RK4dpy62W9ZpIOM6sZD2yHszOKztGN+apvXaVLTL2suATnH8Bv7te0gjHQGfQwnfnBnjHxbgDSb4
Ic9+gIif3Cse6J4qxw69HgTcjs/UADbAARnZEw1CNGoEXoam2/C1gO4iu47IAElsR9a2EM+/cxc3
VErPywv+W3MpQf5pXZ1o3xgtORPqWbNOWuPWEwV4957YE3mpjOBzogANhHBZxPKUXpDwkWbv1Is4
ZcrPWXEw5jvzw3xpxdsshp++wwu6iyiYUUvGBHUl+7XVSsSZrMNn9BMwepz/H66HkRxi4xeNeEuc
0RAmrDgu3hfynWhUA9xJlV/YNfolbV8JrUlI4uxBY45W5VOOSIAGjLiF0vF2bp/VQHDYa01ssy9J
PRZAtClZ0vxLOEJaZjOR0V/qJ+HYwtCMZu65EYwb29Id9Ev6oDDha6QYJb7QWswsywe2TgJlNqhH
H6AY2lwFdBsD2Sd9QGjDO1BplqJTJwg4kMRmZoDVSm5FZtCX7556KmDRZxxTIZ+FL3/xsOxvcLQQ
w2YMPKk8hLxS0MtLTeTtjxMM7BzNoD/U6qYoExfFQ1VMvPgUS2J2qybutRj8HP0Yivy3Ix3KMLJx
fJc0uDEFV5vBcEdDoVeEDZeUjpgQi3iQPTlRmsJQNdWCkUdYFZsPQmW+6htGnoNIxDGF99qrL6Um
uWKF4A+4UiCweak7whvEQonPKCzqKqP8Lz56wsR2bMcB/wBb2tbTp8q3g2hjUSsxulnxK4PDkwVD
Q27agFi+8Pg2RWvoTC4yKqwDUsFWOcXPJrbDW5m3YPCFAxere7LcT31r9d/Qd+oV/5W8ke1g4T0A
yys64yt/kEPWdP36ZI1Jfu0fUQOkn+OdtosMqmq4F/Y74SJBP5KLd0vFEapaGpbb+zN1TOAqJL1v
T65NRbaMl99+uyZ4l8d5zhBxe+wfRSP7pdXWTmnX4AK+pJ+x3ELZAwF7SLtfMy15F2D5B8yapj71
96+vYeqz+3jQBXdbzvG6Qeo9AninvOcPSH9jLCxaN3Ne7H0wyEB9DdW/ShGYQZWWqGwsMh8Uhedj
Ov5sllbjtipHk2ESoWcATlF3EgJuufSdOBWAW0tpCV6N/HJY8v3albDWMckhtrcoxZVW/Q746tT7
Qb73VGD4H2MYn1368elxVifeiWJShWTF5j6gUnDFeWoiJ8RISVMJluIg/KZWQB/jGOFkHaQBf4bo
LE6mVoXCnE/lJeiyio2dCa8pR7ylOT7rwPMxG04yp4bVBCHAASWzTZOGXyF5sk/jNbrAM1G8elwO
06yQYr06TOpO5odwiXvbB9xW2GVeBIuhsqz0bhBvii/JghRTrMTA9Bfx94QonF6w0BaEOSTCXhyh
FxUYYjqLUvN3NtcHLSdq3sHLfxcFZ0RSNjVtPCAlIc7UGB/LgxfCOyoZ083OcwoXFjDHZqcYaM2X
a88jYdy3M4GU1MCM5cl+U15VCAgUo/iw2qW7cNpY3pwdGzI5KSvwoHc9CNwzEHsTOLAcUAALYtyf
YM6Cnz9qmnwa4VmtVT5kuPCuyqiUY7Sp1D6eaQaMpJgFNEJ88Y8kbk0z2MArsPUA4FqtoVV6jrbk
6GDC5uHF5CX9U+kyB21IXhTLDYan/tN0bG8HLgwcart1qakWrmznpa1mM7EtnUmrVGLPzuwsSA1z
xmmPez1pd3/PaWDmeYy05ju9SPfVC2TMzdHSa4ziT/YvYJde4dOvQvbS01qL/s9/o45SRxwFL9O7
6Fg/5oem1eqzNIOtUccJtJYWRqVkhRcOJXJjV4hUTGd/mNWFABOpoGmC5I4TdvjIiTvxvKhzsUWc
6u99rPCzkJmivgGjZCQkPBa0S2HVl7MHjdM/JvRNSN7hfEVuownGRFjRcVMPTi0DG8S3eo7kWTR5
pdTaxHK7Pi2yIsOYYCMivwiybW49cMZZqQWFYBv8XIPRN2xQCWIqufpV+hOfiQa9V7y8DHGCEjUY
iIqSFzIM8aB0GhbWQ08ydbOGpsdoFP8vzjS9czZgRcBLmdC5CWDQbzjCfCVgXjFcA0Bie1a3kjkY
Cw6+Z6YYObTePJNWOL5QXOibaHh43pDPtPQVOSG/POffMA87HmOIjtrlxN9nUj8ztUSuMIz0l6Re
mUf7j2uCKHn4n032DdwRt/Y4dPMmd3mb9/gV+r4IeZYWVXSRQr8/qIpNmeq2lI+SZaYKSoA64/eo
7ROqsvTozS3eNRRT0YOBCKUNKVeXofIhDa+JrWp4iIOzHnTCCjUIa1ysfrk4fIGucEs8I/18zv6p
oh1TmunMXyItJuIHT/y/8Mzehk9AZq3yO+EyCiev5NvbwCL7f1V/F/1CD2wHgVL+tGxpzId3labL
E+d4IerwiYrJqPAr5hUB9IKeV5E04pFy5W1p6iL9k8li9e5SSfUhiRRTxlAnGawRY8Z/kX+GoE4E
4W2Yi8y5WvRojzTvGeXCgGJj37O+Bdr9zVD2sVSgGofQUXXEIFubI8nAZFi72YTcoxrM69mZ6o9f
6ju6e1LOoLF8AUoVSls42CJV8pS9jg4pAGyg8X8hDoWExGY8N5NprQC7XWukw1bTjiLhYdTGfLDk
NtuY2gyR+divyaKvvitq9yL44DbJIUxCrvNyWr5lJOIZd9G+XDvVM1yTgYv2TA6M+k8nE1zh9oU3
63Qsg07iaaQP20rgbUzxypME0pgR9vVvhM9CeH7HXXve7uHk/nzCMXbo3wrvfVDpA7sUinu4FOuZ
DaR2dHnrwRahqjb6KWXVHGsnuG/2zND29swumVXtTt3CThThCbF9Sdq829k7lvwT2qX9vjwKoBaE
mRWavdgl1UwuAds9uxzcqqL1r1Pa7lBSec6dM3YRGzYblMFHzXR06U0Fms8t3++6dhmPmtYcHS7i
5kKd6A9BdsYoS9m42YO2hvrbP3C0AVBE9/bMjIIe4kde4rOlBY3ecnW2yZQJXzJ/TRjZenR5KU19
ISh67orYYtHMlwH89FXUIwfMhosB4TUkzKp/eB7HJ6QsEOeWGzKdjNh4wDnUNF9Amll1bQ9BGbGL
FnRCcL4zdbgWJrbML8qHe09mpBfBzwmKtZY05q2fZAYPdRcLISfNspYUNKGHuUsSLXRqtaZLK7Mt
MiEqF1B5vU4+SLGjg+D4D9shzdTfwGrvzAdTz5noxaRN71CI9H/3t4JePVsPMkNvfpjgxLXvylTx
ZLrvpFIMG8zQ7+Ohng0sUoZbbeWrZrB5lmyBbrZ9PUsPDHez+9l9oG6M1tQllGQ6n4w70sI7N27R
aHmcvTT5B4vpQOgwTTpm0vjv+9biFnDDiWOpf8Fl8BrsQ5pZAXuHTFw/RohyviNh2Q5j94rBOlqd
wL3DmoVbK9BgJ0oRU+w/vDL9dlQeskHrwWuQTkI4d8nrt/B92fi/YReVBnTmwIJn97eV141NSOFf
aJMe2Wps9T01VqVUVRDBrGH1fmBK8cSGMl7kAVegOEaAvHsRp3LfOwNfB+qDtYBSOO6//BN8Fe6Z
/AR3ybVj8s4QgMOIEEqjgsNx9Wzdr8HsKnFzEucgumXaZGwUfv8xhfyECTLmsqDnDFdW+/M4zbIA
fx/jcO6u3oaoUsa/m0gNE+oUJkOuCsu+ysNVzM1kjpLSqIN84n1WzBUYRgawOkMmAbmbU2KWWoyQ
LfSs1r6V5ch6a9CItpEWmbh+8kDz2sGj1Hp9YA6UNco48mxWM0AoY7GFk5MOGLcSOvBNFynkZB9f
XU9coIAw01JZXkH2Pl4XpdaKk64Qyvvv1NO4VE9Wn/6kIhZdM+yUFM8zop+cf07gsvRE/Qcs1Kqa
MWg7RRHjErIBruLZkpxLdn6V4IR+ithT6XyXsqpBiqtJS5FvR1WEbxmPBhmHkadEsx7WAMHSKrr9
k9aWl723i5SpojRDVAz5IKsxKIZJZDVjOUZbDBHULwIZUAzp9YrRZzFjkMPl/+0k8uLFQnunwpBY
fA/RzWfWSTgv3FBWrsKDjcmNkwonbyhaMdq8yoKFvpjr7Pfo8zaa/GH/ms8o4/TeRzPEt01zYZIE
gDQDOpq0LgdTGJjlDGviqnfN3o3EEo40HBJn56Ecr5H+t5eu5wIzFYje2N1F/n2H8uOP5xlpDQ6w
lSDStuICnak25PtSPrNOaYNGfqitukp9QM3yHU86I1rwspp9efx9Zc3CRfoYBwYQp/XtXVhl1rms
zgS51uHxMVfxRflyCtbVecUJS7S0nKz26bAm0jkO2nRmuNF0E+zM/uXk5w3//+GLuwzPq2lo/1Pl
YkpP8xUQ4L1rGJtkIY4Lu3YPWSUkNMnFcLx3e4SIE4sKofOQFgBuP/1vCdSlugl5Yj4I0XAW8cQG
y6DhLsetIugFAQq/KPTae97fH8/wG6Gx+1WzMEBd1Jpij3AP0opR7gRBU3iYoGIW7EGG1g8ky9zn
gvFB7v5iNP8QlkZ8gun/lcUdegRVhxB2ySFFYwoX/10q7ObWA+6QZrOCXwWdzEeVIVH08RMUJVBA
mivJqcQHhFRigcHo8ESPH3gnDRXedjjsibDavOAxlF4J2B2k+8GPbsvbWY5xVGdZVK3b3UFfCkAY
nDVYzz9vKMKsdEXb3/uHKWocp6DlFljszXcGFA9O9ZFyIhdn7sY6eNNySpPETIBuOJ4/l3mFTiZF
NUGIXMVvmS5GG4Vc7B+CSyiZduK3jeJqN2azYubUdAqcU8LySUMDhVm3ZYpdLzOJtksOgZ8lHtuj
qdOCnxKRyNCImfHnj5ev9x4m67+0PLoEzKubVsiIYZ7zMlhiiX1+xtlPnV2e6Q/xjfPJi25Lv2hk
xHLza1+dMxYRLY2QkmX5LwX8++KVPCcismR/0NY5/ZB/wTvgPou/S0Bi5qyBMI4YiTI4PNQIs78L
4m117Suc6n7CDYjbsoe1q08/Kfe/Yw9DNhKK2R2DGzLVDr8dWI0eeqklJZPSm7MdfBPJJMXBzSZW
3dkSaiPtFnygkUJXCpuNOvCYCMe1fWil8KqajD7cXj4XdfOzpffhcFGxjb7AGT7a0eFTdcypxhCg
dxtj0PyeYSsmIj0eIv5JDxRWf8wALcFEJe4TM299C2wJhdV0VzRlyJIqOzug4GCrU9X9hc91sJEb
H6HSM3At+v1KRb5NDhHd4HJQAQRCLXgmE5Ww8mweTd5qG1CTs7hGDpuqqtWQHsJALyslkxBZjKW4
+z/dKwykU5SmcYdEcNFQKitHLeR/1sKjTualOdzYPXM//wkvrqu268Cmn7GS1OLw7ka3K7WpkzMs
4f84cLD4njhuArAnQwuFVUOOtm/7aBWFaRfmSRO1ua6JLSKnUPvc/n/ivTDQBVZ1xAmy6Nyqk/iE
FZD7dhol+lqzuORAj5VqNr4YoreDBizYh3jyxMsoWzRFp295AsIWcjUNPfRu7myRPoftpHF9S0u8
xt5A7Q7PnCTGRb2l6dTGAevHJLnNeBx1MhBhX9BU9LqoIYghYVu9/oWrW14IT1qYNzjXwq5yl/3q
oelPkWdWW7YmW+LelF1xy7H/DaVk7hHmg9n8dKRFMxgNvFhGnNJvLRvyyq4eldXJBdYnM4lmtQM7
Zc9dIEHGQQvxnl+DFe71gDsjrVSxiyLIGvSJxyb7PR2pR8X2PLtiam6WNYfHmWz/don926cFr92l
i70gJyoPTRU9tosT9iK0IpVv7TBnBZmnOsqGtS3s/5GDqK7S8sXDREqcB+mKxFtmeDoHkLWDzwQJ
9iOrIRuiLEeh1vSiTtHfbGRxu7cSSc+FxYRe4LsdXOHbyMRutsOFGpwQesXoRXKsU50zwdob42Dg
q63tBGdd/QcZENGQqCITAIv+91KSKbpa2eTvUiruHpcpufqgapSJVNkqRGRYR+5y9i5P3moZFtK+
LnwSHeKSvkt1HFyU8118s6Jlpafb6CFkRoBHtHwVhU9/5fKWWyhFMU1jXwKMIQmj5EQ1bHo7A3SZ
Cb7pG3d1WFpX2rxXV1K/r8LvtlwNTghmdtUJbGwqpVgWJ2ObShcVHhaNYpfp0Y27hCAvelhxy67B
VqJDJ25qsc76xq5ky0scqkrP/bdg0Bd2DGnm8nuNPgRChfLDwT48mMTh7tlziO/EN0Fnl3AZYyh9
26V68hmQ1OgpETScebArrBCKgHU2oUgiD/hFf5vQGHGm/yRGFEPtUUDRgzD7bvvFeu1dGGxX9kx3
7QMIknkCmBXyiqvkwG1xTYG4Pp9Zm+dN0pln6/CbljZIpZiO0wJ65pvCmznIf1Ka+MzqzJP8ksKo
e1/Y+Xo51q8WLknCvJai/AGYXi9RLGSHjR3d33yhmOTH/kAAsYNwommhsxtXCg4xjiohYNwxlE6O
yApGjUFeHl4bNTknFlseam9XOCMzhyzUfkGi7QCP3GS8QbHQRqtbmR/1wfoHvc9gOj/ebmjqpSLK
amnl9a3O2Zc6M8OBmLZvi8rWyfHPTvV87OIxtUK/X78kO7zFomXQ4k2O7oWw+ePE72MOWb1vxAD/
WX8lKn9GU7EQ9dcsZ2Jk4lXT1zztnZBKY/i/p95Hbkqj7GGpZyqs6bPSFxKwqcfy6wgBzdg/Y9Ds
TpqQAR6309+MMndYNPisJYhHhIg7ex68PeD9+GtAohkeOgS13A+4kwrgnCl1A8wshRFEdgvLiA3a
b0hYAFlBjqn0IwU3GICjHr2C0yWm2NzgrMhK28iDV0fGefFiJpiVR/FsMpHKdBUFppMd225Zt7yt
SKZwCDy5uIr9WP5OJnFcaODWD5sW3LHXPob+D+BWbaJdLX5/Iq8ftif5Mzv0MHKmWgbfYWMyDVBN
AfZPPQuagEtCcnliI0gZ+2M5PLgXd3C7JsH63DiHq6flcXmk1hOEL2fWzUIGkj9jf6LJBglSvTP5
UE5xOcJSpstHlL/o1mDEM5EbOdiIjCc4qBMFpo/9I0H5Bi+TvV2QQwK4vYucrvVZ62Egsm0Clvuo
Y6sbbHXh2huinIsXL0phVN5UWGLxwq4xor1MwRuECzXUiPCtr0ErDxK8Q9Pi3LzQgNXAxEE6Japb
Yxde1W34ZszVzGQSkyT/yAL9k/H6KqoiJQ/K66XVJujmVkbv2Fwn93kYZ2gRDlc1ciHSrhMf6WoW
lq7pdZgINjRnotvhS1uSOgNhETNO4gmmJ9mYghaIbPctdVmPMsaEh7rjGJXv/fNavHaaV53HCgSY
4TAEVztdmDQGw8iTDJAV7QrP2C9nyqr+5PF392jDHlWnrxfS8/H3Y6KJ0B81Fh7lqWS+Ien8kktb
lpewUAcEebVYA+Qsddu6EOR4+mbgjMtgIxr03YZSAoRpTnqirR/RJQ3fThXwgeXLF1pv8KjEjTvP
ksfblz5BxT+c6IgBsOrMtJ/mpVLxlNgWOUuUmNXj0dSkcLMOG+kdgMpsQN0yKU4Z554ZjjJFXqk+
qkHG1xsN3JHS7XjjeerodBMdp3iCnInMnZJvFTUrWUttuXMKY7tGyuwuVc/P18K/4Kv/FeAyQic5
KqM0hQsb4syCjIHipJHKnvagtiD0hW1afmIae0TJNmVbG43fGCFUwsUnPcuPW4JdfG7BTBYSIWQ2
6tvloauvVM3InIss47DrDzVFIAyJG5zFH7/mv9jwP4wQrKLIbhXjctgFNkG6wYT3dY/ocqw+2cIB
/z3gtH28Cm3JlHUSFu+sq7r8rpfUTL921px7L73tF8LeDnMZz6SFI9/ZsDxMD1PoT+JL0XGUfhvg
g3kTzX5nScByccd7Id8l541ZZIWlr57uPD2BXoSf7zkEytrZHvoLzQCX1at3pxHWQhsSJWtXWAcb
jeiJOUGs0lb+p51zghKPE3BC+KuHzJA69O+J7x/Vhce2ny8pu0I8b2RZPwh5I/eha/znzM1JHxsx
3oaNJQ92EXZVdSpO+xSqAqhw9fEbqa7mmXK4Ni9/HK6NOZA5vQfxdBZ2rhwo2elgXQjtE4fW2YDI
yY45unsyrZspwbEoZLrfT0GP/QiyZtXnBn4HXNUFkrYEfaPX8I/KL9WWo8XTiinejJVAVs9jB3qQ
dDK7bKUvi3AoGFxU+3GMIKog/5fMIYHB6GcuyzW1VKeDpsIXIIJgScfUjnMLawAKrKIVidnHowgM
GoWtHzP5KgG3VkuydvGLbNwQmpD50fcHSTnsJrtEMrN8ZICodHP/9tX4yZEbtJXGEsfZzEkABtHS
3peNd6qbr1c8Ubq2scVI/wfkezgge5MgM7l4weeffjB9TgfmmhPYKFs0XjKqKrI7jwqnPquDI+2T
A2qZPHVFw80CwJi5rTCzVwUgb8ny9cmYkCajG7cL3er3TRLrwXHgPhvOVLWUbSQYGHPtebKkDshT
HuFktyQb2P0W5NSO2MPqBw04sgu2Gl8Rgpmg8OLEK5T7APZ5O/fnMAndq3iTyh9y/tmHPrM+eV8m
2L5Gq87Vt0Aq8efnUtjxbVBQNrvSQJ+imnIzVuhaj0mcbgPfwQUVDeza3cb/KP6s/kqJfJCNv2KL
/GCFQXI25oa0Tij6gdaLeN0Icu5K1OpQUProgJDrgfIUYKEZo4HkCL5aIxSlgLuxoOSpHXjvR+Dk
+fN2NKhWhubzF7ZJoAo22kmTnJcCUeuFycVovB1+AFGnsiD8yYyGAgwetHAN79gnTVdzEiLy7Qte
GR5mONQRfeleq5GlHVUiKJQ+EQVdhGtz/ailTdUzGoZj91Wk01+qaCR/1/WSMWHjiPCogJrE+0u6
9xFqNwhTLmfSZHZNLYRosXEeCJxcOO6YygXd7lLlxAjRjpPypRv+KXkqBj6ND6iCRO9dATL2as85
gOATNTUx6yQwTHuwCZ6h1g+ZJCvSJWLeVaKLNgR6KeKR8uavsCNR4THy1xh2yc6EGirpOQxi+S0M
FcAnnAyI1Z6hLcF0bH+8k5KdOrcnNVgmkwbtunS32zg4plJajiAfdzV9awQosEphgnV+kYoi3i6l
msqomBYfJBoaA2ZYh1LIwgiEiJr8F7HB4kUD/AHwbOUiVvvMa/IRSPiLa/h6CYESHnN4AR+xpY9K
CjZ8Ew/NHQRYhXiWtgnHW6ElQukoxWULx7Runwmromm9XAtXvz7aaIQ95k6S2HcA1Wd874yObJwf
Cpj6z7Wuj6J5Q+utKn7Z/SFxk6QWFKErvIZcqqnfhPouEXgYh+yqI76jCRiD3gT7xgApfp6RXVGh
q8q10udVTXHJTirnFAwhBkkFnElg8NE9EtrA7hX+osG7WubFVBcaq7tiM1qig/AfnLeOQOJR8ekH
fBgdjrYZSSXtqsgPMVMqxzkQmBuIaGz6pcdL3P8+PcYegOJasPWI7PCRR/j4HRe/vMRN0OnQ5g3q
hMDUf4TF6whH7AkVFPIvIfdyZu2wTfQUE+6OREGEFta0VtfUdHpn2dYp0sqCkXWyUhLa+hC3Vc7y
wCH5087GTukwQ9bA6/Erh+6LBvV7BZ/q6LhkDibUDEW1L+JAOrRsds1RGkWheUKtbQWF5LfQmntv
MH/aCgkrG77TzNAaRBGvrKWtTs9fNnwhSsJbxlP6g6XVvSZVtTvUAcyEEOCpJ6FYA2brQuyGnlNE
kFBEa0R1hktIc9DOnFm5O6Br46NSWbmJc0dEuHUeO47jZdgS11LZjCX0y7gUWZaj7cZL7dErh4iN
f+TUnJ2zTq0bPB5Z+leQZtGI12pXg4N9hXRFozKw6wdDmq3Z65Pf2GaSrCXDfmLKMuTuVWL0seQF
NtINKG+t8WlZWjI8aIKn4+UyfYU4SmaFCVqBUxXGcbCOdsPNj3BNHL+FiCsZkRLu88uHwF70l+WA
w5XbFbJp5BnAHoAcB2T4mU1Ye0LjVMMahIuQjOLQ6pt0YcitcGZPs4TMce928YZR5/0BOXUA1o7F
rLFryLwGk9IL62WGkjYxc6zZnFyUf47jYd5D4BxFauXUc651EHr9yHl486Jwk4Wck4b9M2Gy4vPS
LLXXPqKj0gYQSjmIEJZzVYl/2mV02HYi9qjDqhHU5VOCkbBgQzkB+SMyDX6BLdkzOloRobLl0svW
4oubAqzfSD+/H0TzBhluBL3tCIm30ZJXEv+lv3wSE2rMgsVhaZffAYSs/ClmhzCyRdpf6BrH9vjd
tPBty+DRAYBuyUMbVUutbS1MeFWmOx+52oEsnIz6W+HJ242glQ9q1go44Hzev2hJTvTs8Fp+F1Xw
1yYvlG1FowVKsE13CgXaEi5EocKIUIiGiMS4sZVKpMhTPQgPcooWUe+RKpNr4yIU2Klaajn/yuBd
Rp1Em89lHOGriMEDxKmIyhqcw/6bD/KPZ2Uw+AprgF2vkdUME3wL6biEkQtXpT7kr/TyPfG3Fz0j
Y9QsnGUKBJjVijSwOaKbvmVyz42+6ErtLhf6ag681gqWn9neMxxSq84wlhLkwbk9FxmzTTfotCNG
rCKRUaK5Dx55GG0lPhDqzwApmKKQUwEg0fEZQUWfwLl4p87IQp6eilNP36mk3V7SJ+YXiL/zIY+0
UnIqFJiJiA8rhBeFMyje5Xh/TtT8BzKIRTCnGLhsJC/NFsDyE10dO87Sm5iZ7+TcyJA+7lAOMx6U
H37P0BcOhAhAxm/FHLH7QaMo5PS0v4BnPK7x/SemZe3W0W2EkZlPM2omQJ+E3+jx99qpXVZs+nyL
EvzYK17908G62GV1QNTUp8ArWdLT/bp6gXP8lOyIhELjjbVTGEa+N7R6kpLJy2qZkI7g7+mv8UdE
TZTaHlmD/K3fS1vPJniUdA3bb0qqd3h16dgIjtJdlU0EcFv5qI9FLZtxlOk/bv5rnoOKHeCk86c7
xkve4PDTgkssAdWYK+VQQJfd0FNmp7K3NbemKVXxcTS4IC49ytCStNh2uhzGj/sakYyI5jiP0p8Z
5ILGOW4edp78tEdx6JW3ni3bLAS1vHu3OVJUAAwOUVz8m2QOjXfCn20ecrPvoO1tLqNNMFAjM2gP
mMcdfE86D9EgkD5Bn5fALjGJZ+maZb2jbkyBmEtOeKj53X9zqGBUmbYaQIBt7C2kYBnnsjVAuGUT
C+MJSj0rKUt43FdBb8a9UE25C00Q+LC2fkVd0icmluqj1CHNQYLdYvPDFMydbJxnJe/IbyQACDI6
ueLweUbMr2ZCHv4Eiv6MBDwsc+OF0S4FQhwT/jyZVXvID5I5bUXuOSn8xDeAWLhkzjKHpkj7BJer
L0pvovY+XNuN0pa6FIa/vwmWCaRJr3WWj24Txg5NZ/1KWdqOSozxzBQKU5LyXEYF6ZO0O74u5qf3
NYmR7QPVJWZxQf2rbQL/UY9rGYT/e8n699IVGrBLUZhvVnPyhc+PFm5RQQtw7/ynnYypgPs76ZLD
8xTXbYMpL3jtUGGnPmp8njHBy8wWuuZpFdhDcgcZtPxFsE5qr1WwIf+g+jdiKd7BjL18Bso+4Cl4
1LgDZrxfEZw9YuCSEFH+Pdu8+zmZbfClJUzKkv/kISBH/P7vU3/+oust82TNkdR7xiLR+piqemUY
QkXT9BU7JdkoCeVEfjOWC8NI2l/Lk6PxKl7DtnYgeDz9WJEfWU2fmI+SI1TtITOpC9j2vKI8pl4m
fReoFqZPzvkoTficvxxD/A3FZdNGIF+RUGQqL6qkutaqjobsPU0eunQwiIS2puBIhs8dhnTjf2+I
eAsESjH3OdTmDE1EusnfKMuHwNPOpWvdnYjtPj2fz7xSSt5wu8jfzkfBW0BaiE3F7XwfRz59KVSV
mPrPV4qbkMoCTwFjew1qp1cHJla+oJT00urhzdtD3TV8+fqewxVWguCWaYgzgZT02cwcUSxPj1+n
rSG3gdrXtBPGecFFbOfzhUegVG+lz8LnT0FnL0vqmkyQlL8CoHFXY1Xae+TAiQ8UoTH9KzBULTtS
RE2J55KkCUMMd3jcxqUO+/1AacfteECUA8iL21IgZN52LsWS2C/yM1C5gCMLErL0VzEVk4QuCoR6
Ec+EYTEOBeZ43CvST1p+V7GsLzGY82cc1TqzGA+yjpTSkdRaltTICOO+wIVjPHBHEBWKXHOzs/Ti
pkJWgR3DVzlFhLWTXzw+OiOmP43cPtLUI1dR1TvM76MAIXgG3sMhwDxuNfoqD+0Z/fiEfjGHX/ML
NtpQ6IcSgeY6EazPIiNNQ73C4dyknnhCB5kqdvZaE2k/szH/Zb7CWcMP4XwvDFlvmUbv2Z2vK8Vb
YrZ7/FU72JfAogK0Y5eDVJ9SNbaApHx9R1Lx2jDdm59e7GAXgXEu6sHPPSTN9KCELKhHEzsEglpL
EbzAYXF+hwPHJ1+vxWr3rbSLJjbdY1/D0QLR4uR2kn24ByfQivac9D8Zuz0+tgANMqdHeH+gldgk
3W85d76GJjrVYvqT/XkrdAgL+OUR7FNzOPSOwedMzJBF3TVJWzcP4fg2ksX5TszDsw6ZX6QEey/0
oSl/gcGN6jKILRorhFlY0DfdfzosMjrkgmTB08NZv4NMoSRsghWGKEuh7mWCxPHNuJVsy216FtfQ
u5/WPrUkqPq5XQsHvslISXgpg8iaqp5NwGvePpIXeL+rGm1FSeh4JN0N+eQRDtwNS93K3JlRgMiG
/CVwfw+T7tueSsbpIFZW+3fcviKgrkF7ToecZpT5oxEAyPTzqisLjfjdZdJxBixwVvfi3GNaYIlw
N1IX+ZqX8KaXt8P2jRAT94eTk+ltePNDUaOSDtBEiJTiBVB/Fqkbc2TA2RuSNPTSZUwQmu+toxku
iFXWdU+CVXq1XdpNQMiWSLB8FN+x6bQKH4WO4Y0erCduZmaXAra7iiixxV5yPV8LP7JJe9AHRwTr
ule05svL28EimWY3g8NO2Koo3mNR4pWpubm04qoV2XL7EFj1q2fBwFLi7s2HuzKC96TtxqcJyHRh
F//84eZDAIRxjU6UrtSR51+2paG84HXO+GwciuCIDPHxbXjOMa5RkzGW57o6RoVkOHbr4VvqeNrg
NzB7g4KkC4paDayz4JnHCMPGijggJxNyiuhgYWImXBDj93zPkA92gG5rvXMXg0qITFjMFVL0vu76
6uLnj9RVHMjAQJJ1RqExZzFMwJPftIUGqaaPnUj5U23Yv547DdCQ7zT6OT+4ua1EO7OqYVuHhLug
CQwj8K8FHO9NieEg72X05MB/lLuWL3ipfrPKczmOzGzFd+j3qGUZUFhPCzi8IsNKjBl3zjaOCgV/
rmI6kIOgksqQPwsiInR7puDRsBOMvb3Iq8zxm6ZVuxGVzx99B+l4We+nSJzlqN7OvTHtRBXvRhMV
0ogvsx12n6aSSeCpLQ/SdoJSXMDRDdQPTybjVWSogLWILsiXk/faPD+bT51EOYhhwkWVEKucucUz
/+B7AHHy844jdHDfm4bOg4VpL3eetGUfEGEuqntkE0HUmG9l93VzL5xpIQGit0U36gOzpDwd+kj4
IJKSMMRUbC7RQ3c/OwuYN5ctGhCcCt0Phgmwu9xNep2BgVERhhB4yfgzRS09XcD/s+h0VYdWD3Vu
JKCNyO7zuoMJ4PwphPibhXBKATdPkUwsIMpAS2br1QZBwWJS5OxPN7q/KgPLOvoUwvIl0KDUqYY8
cGwqXQ6oJtrt4fPHukA7m9ELV2J568zeCLqQ7832t30Z4ZmKb1M3iXE3EbS8NYbyt54deEA6F6JK
qpP3VLpVR2InDpj6EtH7KK6u1O0uAPRmjJhbyeZJvvSiW9Cjv+vFWpe4XzRuRkgwQTybcVC7pNIk
UhrPsiAowVSKUuXdfszdI/adpsXk23P/xn2R242znitYyWMEt6yeBXJmre3J42sWUTPQtPmXc0cJ
4lOdJNVnrPCe6S01f7VWrprVO0sCJe17X0LD89jVkuapCgJcAn+Y0M24ZF0sONJvQ5wzpfbBdo8K
12bwOBjXv3NBnTRwlc43Gkwr97cID+/dxKKne7xdq9smwVLP+tb2UTs4+XAcEPkV/bCRarPX6Eqr
1gkhNGymXLIgIl9h7G9wuYfq/mp9FViMmzjO5C26mzFyn7nd2p5KIFbcx0BUkTLv77hetXraO9Bg
Wqx/VsTTpvDLG+GgC3usZhLrmqcLjriL41AjwPN+HrVNpF4Z8Gw2v4rthDrWSw6doCwAcT4wqM2w
QF/rl/Tua2rcLG10E+NO1s2rzzB3YzBQ1s8X02Mu9gPoCAAAeIUbnRFg7TjTnGbu9RSbTFfUSSsM
NhmGXp2GAU2tBfvdSBRLGvObPJzhzHp8ehcyZOLMe7SDuhxh2KPeW6IAWsNILqg3d6QkHVmzB8KT
KcesYv9KCBKnBfTZ3A9gh6IcA9sQrrXMObe8Fl8WpvovKSBgdn2iT9W9116QspZXBHNdKnSxJ9+z
uZZbgUssMA1AS9d/Fm8WXxsLHtmVLDQVrd+DJ0fF/aWG4upNBAf+NtKXfqFezxgl8ocvjfyVmuI5
/Cw4q9y2/qQxgkvHoo9ROyGdurX5/gIkga7x/yfYB48ZNB3q/bBLDzQmt3G2Y1VpMUbVYbuhbz+Q
SJIv7huqG7VoaRlZPq/eh33+n4UqGbNIWD0nFSjj5pUtlecgOFm1MQIoQbiXX2Rp36UwVxBOojko
rPC8nBDGVga4pLpTws+dv7Kfluaq8YJKuE8nQFlUma+E/7On5A5RmRsGrDsjv1tXfTAvAgDVwkIv
uJeiGjQ9wYFsy2+sOK34rkCi6IYKpG/+hLvl52+gQDCa8agc2af/zZL+nATOkY5kYrrmX7Lwxcsa
WbSoiu2g7/zZWkcILkia/Jh/dT0PBWKQzakIOgv3UY19XFKCc7gc1DX8W1PVJgou9xyhorDWbbB0
KqxNHxgPg4BXrhGTl9/sVb1TdU4F2c4B6d9X7fAFFMY0OZFbRWd/QBVpAsqn1kCxo/NYqY00uAmk
0an8kIJMhVWe/y9J7ofYdE4NTOsVkNzbDPgaDQD7ZArFiA7RoZMQfzGffRNisL+pWc3JSTvAGPXU
qW3O8JINylWLW3V1kFao6YNCAOvPlhFjlKObPQ75bQ5251W7mdfIJ+TG7cyfRfGqTquKXcn8DOg0
kVvWwJW/JAcq4/76tYxM69j3XUCU0nU3CABJdCUqq4e0yHI82n/eWhPKFpF5klfOAekbEaOyR7EK
J+zbfz0dsAYYeUUIMFQqfw/K1wnupTWtQSE/ulKH1qyfGEAmECWFhOxhj3Yi+hUQJ8D+FiZsNqyU
zMAjRloMRXgidQ0oki8nbgi5u3XHfwg7jfMCahrXfgX2e14zeBn7W0/bQfE+80S3SGHB+E5L5L43
kMOUTajseLGsM+/H9ah4j5dYJFTOcQ2hGLYnK4LVnZh5JOQoAPO1Tjj/yhtTem5rnXI0Gp2UAusI
WDgu0EaE5tC/56Mn+UpHkQ7odsK3SPWo9Z5uL2P0JJgD5FlKLHjzJj9U9iQXV7A3NBOILXvWNTnB
I77faYw9a8bE94BTJc5dbP8uIiYQwMshHIhL3eAvgvAsEo+nA6OM/J0IN35KGHQt2x4cLe5LQnNy
aGGnr8if42ymf+ngvYjnpATtjt2Pe8LpxA2dv2ZSmkxAO0/Xti3kMAtsyMGGC9aMAiDA9/0lxpxG
WYS1Uc9iTETOf2KxlMZBMJOznBnN/lH0B8SHEPu/mfMaGgZrJgAgTnnWK5tVrDYY68nTT9is+4hd
MuXT0GPZtJW8o8Pv0I5/ANp7OgktVpf0j2y+G7x6qDFh+/XKRIGwIXKYzxc92cefNtYex2oDWeDV
iRp0IO5/QToNCrgUXYtlSJ+e1yiQiRK6BoiU8zpcP/RHy5PbBvME0phTpv1MD6RGszcRe28K1qef
91wjUQzklvO7ZVxvitrH7VgeVL/cIPgZfOeHCVcBfLoZAnfyyj2ai3nksNbRhgjqEGg6w66Vn1zm
3IDStpLysm+I7rWqf8RXHf30d4bnLLvsPoDxNDOra91xXdt+pCJ4U8SiiPqD12WYjq2S9tkUuLhz
l04sdPXU0k4sbSL20vlMBskk3Cxlfw4zQBuN8GwR1/eAW9fJ31N87RzGbBOQlBI5IYUyqtHjBjQP
5+UpXLOvezbKVosWXCobEAm9xQNd2+yGN6peK0zrQ45Xlo+pBw4kwdK7+ErIBeyv64cJfLYT+hrb
v2K/8c8PIBOxSxj2fEfz0RULGZceyx1cfJu8xy/6fQFnZCFLaCFEFOGuIM50VF8TmK1j0r0mvMjf
ddaHY6Cdh0xc3C9u7HJPUYYJLCUk53oGecOwcqSgXo2BF/0GR6rc46uXKCPHxIEjldQQNTLPYkWq
4j/liOecFIk1r/qMl03tQ07lx0zfOD2GwijWOcAMsstzNs5MIyHLHjqr0FN6GyJ0rInPFJST32LT
YY85QyOh75oMR2U/NrkWaCoO53v6B9ufV6zNvvwqmnsVc1OsCHlvUinYSjZ1++z1zc7ispAEneKG
k+LpZuk+g7i2Dnjbhfi2lhGHcHVFMWPfETx9Pt4bEYHxsihBmShsmzVonY8PKBAlFsv/yUhina/b
sTgdXQUjj2Pm8D3qxfzgJ+f42W5zCoqAnZ7357ohJ2zoEqZAEm7fIvAVR1SXyBlWN+oSanzO1rHy
K0HHmkX3HNOTwcaZ0nA6jAbs7Ne+OiQC7powBK63qXCJoeuGWsIRrLKAVLmPumGAHgcnvl1UduAX
QUUPF5Ud5TPYWWHSDhKAI2N9rVRAKm10EJg2+qIMAiYY2mY8+1lnxh9YBS0UUGDVy6DdZr9Kn8NZ
3KpzDUQAj+BWIXgL5pz+2SbqTsjnLdQzyLQuJxaAVAadsXmmZjB1EQ/q/czPxQaR8UCjqLXe7qlq
w0lr27DjQWpp4zdfJ4+tc9FEON+uCCUVVOZaLf1Sbi2kuhFzqieKZaNBvbMch8YZHAqupxquqhV/
H1BY1so8Ssev9W/My76mYUWh7jkOeVOa8kiUnJOE+lgnzwOv9LKJso4/VQMQH4nZim5wgxHsOQaA
KAL+N7oBu40OXViX0PjzXBgh1dpGY/XY9dPom/jVyRoku9AEpx03pHaE0KROwtZ0xs2SD9bZeYzv
iULtXla+XCiYjwA2wuzWh2V9mEXAAJvHDQMZXTikHqbw9KU71tp/4uTH3okhNeqC1mc4/VX5aAg9
2Y7oZfAE+iQltkrtJTqh3nmNxM+hX0iC7rAAt/vTzvEekAi+S9f5DugdSLCwjwV5aIKOo3YYhsm7
+Q9Gqq9X3IRbtkfjMauOXbzv0ZE9C8kLb4C2JArpQv2JhGJiZ87DC6n85fu/Wu+HAf757/xxJgZf
6tpJU0OnmrWhOioAIDKMsi20dd7hDHqCm5Y8lxvlpyRph6sSjT4SmW6RqWM07wmAKtw09WY7rt+M
Gck8Hk/AGTUGZRX4Dwx7XpqVt7Ww5Bfh9u+WpkrH426UdwkmhT7NlEzgn74wUhI9lS9AhZYANMi2
JONFtgmKVJY8akGg8o4UwLpL4Awbc4nrKpDYrIYsqxZFKcqPHACBbhbjK3zwY9Bi652Y8huB7UTE
85ISzXmQzVcIlGkQAZhKa+oQKTaUTjgWirIQO6r2SRzL4yhAq/SB56Sob+zd4VHLYQH+4fgYJ+Eh
ixE2ELruJ6jtSD5TpSp5IlTjaBRnuYaBEP+rozYAehWN8n4yl9KjJtGf3RB8o/ke3Bv+I4nEDQ9G
ujVaw+KosxVrJICLSSPTEypAQK9Jhe/IhNgzwAD/YO8NrZr/yI/yG82l6pzfFno2S8Z+9bCUuVQA
icSMLzOQB/uLNHLiGMCb711bAcMG9FIQwNSDyrIJzg0L8hEpppu0NlfOEgcxvdRiMzTTcFpfWTWI
HROp8C35ZHPzCNlFTKkQ44nUElHWUIoRUyKALUk9+8GWAMDubHdFe8a/vI+1yywQ4+8PNzOzGKMN
h16mjlJCvPvSXos3krclTo06eRzFdEDwR3MGdXNBxon9WnmozKGY602vT+xfqRIe0gfa1uWkANXD
tPbChGLqePa4O4G0NGL6pEJBBKUR8QHUuT5y31J6wHjJfRGJfGu0GRg9knSp9WvZqVjBoEF2PZOZ
tmwWP7NE3sfPUdToDV8XObQongfme9KG7WJFBFETAnw/7Bg+R4KelVqYi7smqfeJpKI27GzVibS8
RQqZHGNU/SBQRoPB1Gy82Rq8sFrpiDGpNEHuNDab82p5IMgsNKnuw63lHhYXT0plZzz28hiEMeVy
xoA/qOBeXLeZ61/R1SQFC+2Pyq/ifEUB2f/dVJfuQeosWMKG166pAZwY+SxBVuInLg+ennMLqI/0
umkMtGPPT2JgCCDaHdoPdpUR/EqjB9UITq0vIZw1CY9Yb9BtEgNlHr+TWnEKz/FaSCn+mAxNe3Eb
KBfBkn2uvNQR/ckvhn6kDlNDeUeNuboEegdvwG+xil3F1lPIX5uW71Z7YekqMCLJQLvRfZmj8pDU
+T5hWBnAsOdp0VoqmNmScKVJLg59op7+RmU+oaOeJ20sVuGnUlD1h0NRpqIKiNNCQpWueJDwX6BH
cOwzm0op9OgKWPxPD/P1WPNoOR7FHS18LvJm4gScmX8DC+NvddUm27akatHdXdbI27clOSivaMOJ
QjmZeNTsANG3h/K68lDtjRm03emTa/2yJSKb2JAROpl+2y7ENiScL0v0srvBDC0Fv8NCJFGZItZR
KNZbDyiEQRg9YwldNVg5i/h8MMDIsTK+rOh9Dm5JJutSKRHDTiic1mO6+itbEN60S8zxaHDTTLqG
4kXcX+LI/pbv5bUMEI37/2CCg1QsGKCylBLJtAGnQyAcb9QRkNao7xrgfgiANUQ0bGn+hnx1ySrI
8aaWzCuv194byGFFAcZTbmx+Ru0ynfflb2Boovyg5nfPzYW4pEdlk4Q93Jj9DjfpRdrg+AvYeaWb
5F8aee32G7BTHblgTIsWOzcjF9owQtq8u/hOe8re3gl7QnKBZ1hzl1B2ReiGDen7QvbdaS+w1BzQ
NnuEWqspy8BhxULkN0a6M6M7cCNEbXnKoM7zyLJHdI0qotvX6RigfEFBvy8wMYw3NO6Ca+ETFlWj
+F4Djf6R/jynvETNi0Cv59hkVDRAzi6cdBLzwrOofSgsD9RDESrm7GSqK1StGq0QEfflfjMXi50o
FjHYRV2N/zYc7ERUa9/X9zdAxobZRB43TMYSSvDngr4mrzTBtAWo74I+ld/+mHSlUzwzYP2vpJc6
a7iT3Gnw7DW2e+d/xztstKmiWR1AwdTDaV5+LRsS7bxLDh+7iZDFdzQDPsMiDuT3V69AHFW3e127
eCx7YvrKQhi5oM3OewTyuVs2jdxEkMOofP6manZX4iowNV6sDfJXkP6UHeqYUSaARYPCRVOCiW+f
ekrPD8toB7I6CfeS5fPOhdxpeEPiHVTQlaIqCOmZDKlz2SA+jC7LN9kId4WU16GIKBkEwBEExFpi
BHy7zR+JRKzanIO5hMUBdSDVoDd8Sg9q8mqfrPHXA/I9I9482t+uVrzRc3jzyRWP62G8rIAUOZiv
cBf68ajV5/OOLT2kKL7JJNX/wnwV68FST8vLWOHUZUptRcpjrV1Jau7kYC34KE0vwtyhbaa9e5ck
4NqJZ7uKiUj20cZR7Nq3qGjzWUZxlf8pWlohZVGFp2sY732Kp92RkZ21k6fyhafl9RSH30Rz4G2+
V/MLo0/FOUPHFUw5z1hXaOJwndBLHbozPYxsNUMKiAYHoo3J9lynVgpiN7IezKVI1QmcEcarw2+N
SS49NN8Onyj1Sn9Ff5o2q3XVCxNJYDlb7rBQefl0rJsNGJSmF2/LLgH9hoGmDVJc7nq6tzjnYFbN
vUf1V0o6bk93exNXaXWOT7Y3Dn7DfSP17SlDRkJ8EvHiQJyYqCFYz/H87N2Ed9KPPtoAgoz4/ire
mAt7EQIPSH7tL4ItFfc9y8UxYf431T6epRIjHAmtbzANe0h609Ain3rly6pz+TQNwusIe+cn5qtS
sNy5AQQxOm4V/GrfCqJ8+Y7yLmJu2LtU1IIhn7UpoAIqT/ukw8ucL6QmTUtsV2NqFFL6iZu9JAhR
73plW7l1dLQe4hJskVAjfUiiMQPQ2tV6Xtq6vLUfXGbKeuTnsqgxsPtzS92dK9cd4dIsk0SHjl9e
N9mXl9Lv2QWjkDt8M3Bth/+VoXH++aVthixXr/JlnkxZlc+F32NmdpxGha/bwk3UBpfwMD6snJe1
UWcM1wuK+HP8BYXwB2Y2rrAiGdzH981Vq+rtuPLCE4a4DBymzhHhofKrkz/3eaMN5nQO787Y0sox
Z37aRlSsYx1FzkNRe34w3PlutA5uxlhQR8UqRLnhqKXT2iq7lDYRDRco+IsJpoX7deo0+1x2EG2m
XS5XbG4gJQFkdCOlbIVnGI341m3aJhMhV365J6PyX57Km/IAmhnWDWNWqFvJ51uO/k4cuXiHw4Q0
fRaM+bGsxeb12yeYQBBh5IVkkzUP9R8K8+gAXecKmdYokgxzq6xhMlGYSrCFnvokzXKTC1Talw4D
j7oF05mYWvXa4ccPxI11D2M37JtPhUqW9iHTflwHSjmEhmItKTaISpAOwnbQNuZp7avQC7XeO7us
TSu1173SeNgQs/q6y/XEILKs5kumwwLHwwbulSmW9G/p/UN1tpviZVAyyjfGEK3g3+iC6mwcsuXF
qjZdjd2zE13r56cpBYbtLaK5GTgC/g+jZ4cYa3sQrIo5vuuYbRIXmjJ2difIln/tk8xDtbsocoEn
vRv4uJ0U/zmDvCpfeXxb5xaIocDOnaOhJD8M/0bLwfuX48tYc/e4g+9xwtpsY679vbv1i+xWTPhJ
6DSLRc6G5vFd2CAFueMIRd6CooZZz45rzCjePxNROnv9Qas6JxL5kYOv7I8sJek7jC3cccufSgXH
OS38axpskh4J2EwpGfCRpTGWVd9s1CsqJ0DhB8v+8cjpXvIgvd3AC4cTFvi0EZsPixVk0bSx8fNw
1gg5Cm5Uk73qZvmDefzj1gL1qQRLHn6mEDJTF+Skwen5REzAqSa0vlanCvo6TM8dg/NnI9PnAPjA
wTxi3ImTDgKUgJSq2eNyIlEOFOv4edNOBezK4UpHxsD4VbVYzEK0EAGtftqQQvHVuZ6kGzkzPa2O
IIaRicFl0m98/31YojzVoeqwo8A5AVPIZQOxq+heNymn2GQyGdyE1RMwX5LKYuxGHGFAkVPLq031
9HagMovFMzcFEAsKKO6RDFE7A3xf4/JBJXZGLDU74XBP/snCtduHH86L4vyMhjsDBQMmIg+aqmEQ
N+m5Ro2sGyW+dy0WMy1vES6yUiyQFOY94qRC/XGR03aEeAvNVGM4LgYpI3KnfIBK3Zjg5iw/B7xp
71F9Gg26hDzgc2viXcFgskrCtf6jak7QOq9Egs+kN8zbbCX/rssZ77+nmvtOmBmALG3yx3kyjqAM
MDFioiYLCDZMD5+fZAsJF+yVaJW6XLl+4B8jWRbWKkYSlnCdvmE+iTEBy4QV2EhIrBFPc4BuC1Ij
5ipiQhHX7Nstl9HkLt21bBOg8PNejhntLFE/mbRLKHRrbs1Ralo3gvcQJT7isM8XjA/uVVXZiZWa
w5Dq5RUC7R6/I4/QWz0TCd0SJOqOwFMDZgU7jnjX+pBr5SSuJUlh0GJJGacRUF9Cx2Q1ENVz6DjC
xXJtz/ZETYC3mWSqPNuL9MpCsSZpuzqmkzoi3kGyDShtQ/9cm4PCD4Q3XlEVelPKSLcyoKszoLP3
TXnn8vYiGwGEArst4A5/XrjuImrSMBE/FuF0Y992VZKv87h9cXrTUV2hJk5dL3vAo7wjUc1x2dpg
0abSXLjTSOhPWt3MPAxE8mdRVT1IHucjVFAsoh5BVU2xH8/51S0bND01Y6GBgB7J1TU62I4begju
Fe9Wm3fRuS1r+vBsxKJKAfYsgiEqmSATmRz3TVBPry4+iSnlEllwU6c2Q63/7MyLNAJUwWEFntnx
Ir/zIb3BqybRGB0U/mi9sqQx3Q4xoNpgQwaqX0QFaCP42n/WnvM6TpNBtn4YxHd5HskP4IthRSdK
vhsKxjU/dOCr9W6KXGItILnqm22tLRZYT22WZKZe0+0N3VF96CgbUmDmjfXfNuyfAaWbYPfkcOV7
aW0chbOVCG9jRFdheTDVoh3LTOoDFlaE6ULCT0XNPyBWinqBKe01tU3o2zDC/w5Pdx3UeMDIsIkF
H21lxLMPpgA+cicypohdsQTdgr/6pLIm15/bX59VNmPFHxDxV9nO5Qa4AGL+ymRzJIAnCvRJ/dFE
1RyDPAhmdubRowO3zmh6E4K7/NCTKmw7j1LZDOfzBc5pWEHlI2MCs1o9X0Hliok9qt1VQc6wsWKS
aQpuM4loIL0DABRnl9w4ePTq2/ZfwRd1E/qdwHHvNrGFCP++5kqPMY7m+pm6KyFeELAG9p46Q6hi
wg/zhuZOCCXPlLrp0rAkrM4C+hvxPJBdnnvCUvNnaeHhqffzNf7C0h7d6q9pWUuFW6jhw05Q9gXT
4ulS58tyTMcRJkcBQ2nXDOaZVu+mHfWj+BS3kyvGk3g3m5FkCDoE2K+5OpblFkA0LyCdTf/EeZsA
k8mE3/juRWLAu63R0LvODZY7njkGTQOwY/ziveA9v9gURnL7r3pe3qW93QXv7gG8a+k8MahPzWbK
HYX/IzaCswetaZvpXrZhewqhZUb/P+YMcEcsMUMNuDtpOmY4tkUG4bWUZ41MFuWr9aog8WxaL3be
ebXMEQaqWyR8YQzm4/Hsu4hGNWUjeYbi9r6oVv1uCPQxJnNKUZr3RSLxIV/9JJ9B5Hfn+J/TQ/xL
CRbZM+xL3FZl8F04zuUt6xNmrvVd1uI80XR0O/PSuEc2YdW8MvuSXAGTO3t90rHr4t43bdlS9LBf
gAeZXlN7xc6dPlCE4xucK9n0rwn/NY0CCG29wCr+pLz7SIuUGoAnzg0zb30SXTr6wJYBSbo4JumV
QY46c0zbzIxm+SqXGnxEO+GpCf24bL1AiCnbUhpeLcVe4JjeCBPACvnhEVi4QMCotD/OeShbRXuK
0gaGehJ7oQ59bD+F7tfJY4bIdGDDh7vzpkQ+P+R3sLs7yBPYdXjG4hOB4LotWsNdbgdH/dVPTDrJ
jFNwl6q1ILHUxswASVzPFnydEAtQkPQTLDCe5ouL9GXK3NMfOl2Wm7RHUcJ6nRIDejj4v/sWi1Qn
fa8jdwF4xbb+d9TfVScZ1lNsS02Gdqqi6Y/zlQzJp9kij+M5/Ckg7vBR2ypX+XZpj9okJ/0JYEbH
qwIAOQTqdYI1c3yR+AZlJ5AH6Wtje4X0HV/JC3+QWaw8VmfT2VxfJl1UHuCEBiEdmqXNvTvBuR6n
NOXMxBuEGZzVZ1OhZqmbo+iT9RhVYuGiqxRMid55XXJ33Kbyx95mj1PsW0E1UpdoRY/uBmAIh8dO
H32Gyy4qbKySO8L+ci0fSKQy2uVQ6QWhUtaSEzB27Hsspxl7t474OlSh1tk7sB+i2wD7JQmgkPGd
d/GmaeOjWa2b70PxLrby2Bd5FjNroIZAoki/uqzsMDDNmJdVNiQgYYzX5YqcVoxDUJx1On/u7hr5
Pu2gns1JB5kaZnbYE0gM3INRDirauIE/n05E5wvJ7EqMBRf8aR4/2V5EP6zc/wWJ8c7+3fzIy0mZ
phkK6tS3htsELogYpLffq2gBikqne3emTRVIinBC7exsDMWob9DLYZKmfXfWhhxd8F+aqwwjYwam
WhcTQtklWRRuRt2l5Xf6gBlCqp3yKfxhQeG3qdSruMUHfP0TA3T6uY6pdiNQurazBPDIWGG24NZD
ErgJvXSoNTS28ZYP5lVPnItkDkFjWE0wFSBpLvin01Fki88QFkbp74IRTnFjSG2za66Hq1RpG1nH
OqUzgWJ0wIcwqGjtEbcnFKvOZ0jrlw8LRPpG63z+SOKTHblIqoxdKNdEOhE0HHbh8NaUlCho+dsc
HzlcDwLOy403OhbXXfAhHGxOtEz/bNq4UBTqO/TzWqWE29pDoQGWDVpHQBv9SrhDBDeYtVJfHkVf
Ysyu/mIdUa6NGqamu+wZy35MyyYh5VZP0jcc9BCANFg+mD1HfZo1XOUHIAs/Losw0chk/AaXH2MG
OWHEAu1bNbf94djYVLN3xsIa6SToPAbSvsLMuz7ErN+vanIlO2iNbSZoa4LNybHZIYrMghfd41s8
P8/f9T9kzYz+Bn6Hrii/v+el6b5UOrTSu73q8Eir3hEcrzCIwL9wT8qQjReE/Pvn0+SjX5jNETmi
Xx2VGqSUpHrfwpe6nnk0m5Qw0V+jAjeoA4yHFONZV/FX58nRhaggDxmkSbyE4CAsi52di91jgGZB
iIFdjg/Hnq97YJsx5gkU49q9uioywC97FsMLgI093Vj6x/lrc8PKUKzEsCifYei4S97hRTZePIty
+CCwuyo4ZUrgAjr6XqeJ5adRCVnwrikQbL6hWZ9S63O0rpnUX7+tyXFTmMjokmue6LWn8M3Y+cgd
ynls3WUoyLwbpHMVn1Seu6r1UPw3byFqWhZIDnMxBo8gmy+A3eLxj2+9dTSdpHW5OzbW+IIQUiiY
4YXmRqUZdIOvZKbaIXGaIZwLSIPCEq9Wu/wRy49o9WfnHa5YDyi1YGRRwpoTbb+cmvQkhqbOqd6x
qY/OL183oJiQ98oJivx3YN1QHpG6hn4byt8iZVD6APXE+rlLfEAG8hKfOzBbqsyuPb1VDmM9h3gv
aYjrYxJdzkMJhzwsrsdQZGCZ3+3lM8tIbBa9K1LRd6rKKP+srcBOioLn812QpPMDucgyGXi4OuWt
jshluifPnyqVQfX4nzkjSFI5pmE2cXlHXNSrd03p6EACRAD6uigIoEN4JFVTu0tl8agWvtQ2nBkR
UOmufOtKk7EE2E6oM3myh2B2FtvtJ5xnXWs0z/Z70s79aqFJ/p8yybSojdbrcFr5k+GXV0IyY3gZ
giUDqrrJZlvGtYTqiLl0MYq7anLYSOV8cA7T0ixMEqfdMvSKlWf0S7vFFthN/J6Q87DQZU4+gGr2
dgAU1r8EncxAnasAuI8oKFvhMuo6wla3z+6zDtWw0U40NSyhrYYkgtJMrUm0As6YG5+MRliEI0bk
40RpTlIpQ6RWGvLegJwCaqNBi8Dy8QmGccyE6xzZd33t4pdmBYxDlKgB/Vkt/10wSzR0uoD66ml4
4I/31wS74XiCGRruHVz4/tWuBoxAX5p7FZuQH+z6d0XH4+uuJYrrKFDGPXmeZCel809AEYwahwDr
bb3GIEkz9tqjbSfazrFUm3NTGhpohiyqyDFqBI9aXKf6Hn0bYQz58N8R2nKVrYFrwIjOFOdrBLMW
/+0pQg0eLVtY2XoXMdiqXVVM7tG79Sv4l5Jg2Yla7ti9x6QC7e7apuTu1w8ivvDAuFDbzNMsBils
CTaE/ueeawVE4AVfZ+A+G8m7fJ3II+Ya6qu1DTG3+qpf3jEjlW7EdwMMcnh/tNCL3Zw0dW6MX8V/
zcufwUcNWRXbovaL7L29RaeOwj5HChUVLZFd2sB/12jNqXX4exh5F/5n8kHnE5pRuWuC3ZSX2i7t
TwUUL2A1a906GhKUW09I8HEnanYR4rDjBqwqeISnbXcDPZiy8xweHXns6HevpADb0fp4gYQn/m8b
Oqc+VYE/YJX/cNQd3557drIIIkIBP08EmqqaE9u04CgeOlIso7aYSHGZs7Ztb00tvFjJyeKXPr1C
PnPsfCJqHTvyaTgSDUSWggB8PSnri6ujaB9I04HgAETs1GmWuoI9BjAtuRcFJjqyroYQee/lQ5+z
5seN+irbpihp/Ow5eRzGcvbrxgG3SXq1uR9LcNzg8lvHGtD2+QU423sKVYfi1Odid4QkRc73cuHS
HPPD9kfts7Caqx6gxqyqj0BRHM7DYXRSTYKjc91ToZy/y9rxelYXWhkvy+zo+mGVOPEvdADQuH1J
6C5k4GfIIInTxFN1Lu5ZU1P85iGSle0RWgmy5rmQKeq6MrITRsGNgT1cGRQ6kH7+hrQuv1woIjgs
RDohYuGrnFjlqrYUpwtXGuxeF1vX0GcFEc4TGr4zAW077bTU3gSM0M7NoUwh7qRIxrG47tjEsxpQ
gqEvfQs7BKnmKgwfhdASx9CWVdRleHnyee+4zTlBdZ6F/tDLhxjppGxherovHT4jIAZojqLTiUFi
kmWql9q1uXBQFp+ovdPUUDbNr45EDVq3fVb1UEWs41xUYqui3P74QsN3p+c6tXht60xygbXuiOAz
vdJmxeS0/oa1zdBDzs7ykH9YTHs5Q9PsYzNB9Tcbj/k1yYGQ5bpFxe9eRzWs8BBiyPC9FHIUStup
94hUF4U3ALV52rlLK8FBh8CHlHTSxzmAaQ/nTjH4n27nO4OV3+eWNzHXFK1PkyE5nlyhYSrGf7fE
iavlMMX8JOT9CmmkVssgabwMlUxYtKPT8UBXB8iAvFA6WFf4poYf0aeyjzAg/exZ7yYfiiFgwuVZ
r8jIE/tUY83BQiSzBG1ZYeyov5gqu+wnVb8Bwq6Rl+QBgr9fNEKLo6A0CAw4nBkVpjlVJP8vFdVw
ZaIVNUPBMH+OfRAdKjoIDhfJJC1D9YPb55GFtny+tlpL/5T5956pKjbWuePqQXemTiF2ZIkAG4mW
+fHTnxTXFP7NdP/8FmqXQZJmN69yTBLXhcgBqg7Y6bbwEZYuPg7NCk0SFPxVnk0zBh0GWNxSXQoc
alieOcacLIjdKkP+9T37ENvH13ebFWQflGuQeonAPxDtns6DNCFyMVIjgX6tUznUVJrpeo8XmEpf
H8uFTxPlXLgUMoe3BTu2pC8DfrnpCcJ5keYeVxVRzV6PI9cDh1qutZzkgP/3zeEkD15Tp880Co9H
rUNrVcTAVdgC9lVi1mqr8hiHwx5ewb5m/x/ISxitaVRPrFstEvryJdhuq9BuePNuklOaEEeJsxmp
3vYvRnh3mCvnoACc6DQLeVIaxRTGdne4UXpJDWgZz+53WjXwtHuTQ7OxH3ms8UvKifVAiyKtJdlS
AweufcRPxVOMKei6/Na0rYDE9hYlmV3ot7C0VzgBM/caUSvcMfqvloMr2CwXxOlYX77R5nNCFqK+
oivABlMhazGF7o3ezX71EIloVi7cpqTHOqrYfQW3NRWKBGyQAonJobPoCoFaGjXHsk7Xj78s1hrI
jy1izcxpysTobzDEUbjgtQ8oL0Yk+gQ7n9IMtNCtw2DBmTWJ0eSxGxhYJZu2HgFwj6mGtEzMlMe9
6fIqlKFkfnViJViWFl/yr21ahM/e9YDY3NPU6sQ3UeBBmN73ylXMOpUWxyoQ1QfCDMSQEFlpViZy
s8Vs1guC2dKxTX4zEldYchy6biimg//BUpMdZ4hLlAsjjAmKSWzr8buK5p76X3h681AceVASQ882
Zjyt7RMirIT5Re/7jCr8YoUTI4nZD3RoY2vWf8w4fBfr6nV0vqFEBuTwuUG4W1wzx21Ty7I3gn9l
X3s1ISeT1J6n7I43284x0d9QbKKobk4xO7ZliVKUEP06J+qUzEX7gOxSq/p4TV3t9Xwj5r5/8UsN
ETg282IdshuWV2YzkgkiCWpO3zP3Jo/KrlBSzVhDU1zG5g+A4K8sV3mpu6DBF/en2/RZj5nqW/Tr
u2OYsvuN3ljskdWWHP/9iX7xmiJsnH/GVMUZ1DWP4oJoDGAqs1Xj5Wxwp0pu5sd4eA0eYx83Pkzn
IGaqHkw/LBQAYr1/RxIHtHfeLcwC1MqgvdbVh6w6bj23Rmak0pxPhIldP6fhrT+LV0JZdom8moE9
ol3YYOXhkWKxeKt6OFU142CjWkFNcJI/0NxEx6fKLr8QnGKdAa1hFFexJFhw02hCoKJTHBundXL2
8JR6uToZCx+fMX3lGKAc4btUjAagZknPOPa4i7xPsDrluF9Wq/oIrnPZP0FUU9C6u7w0PS0xnsv0
wBp4vIClsFgGRo2mDM9NWQj5c4UqQu6dMJIzVj8IrUzbRqMkYlFOrQyWrzmDREwyMzgBhSK6ZWuF
x9FGUp7LguxYIz0akLOwPuaYAspEpm90majpADEBmNgKTSOVF0Lfd+Sc4gOeAj/dinkL2K50BUHN
ZfXKfmHNrahYljoXCnwz/LBKlQhupE0zPvEN/taVsCCyvPwk4Zkc/KypqzGhjxCk8t6mPdKKQOmS
zIUr/0sIy1qI4iwEDWXeJqvkkjVH4Umlu74vC8LD0pZRGuHgbrYj+W8TkXcW+M0Rua9LKVJ8qonA
2HKuoa2tgV3GYjQD/EbT0mxbarn7p/UlqwGVmNMQMP/UfQRS52z9dP3hbZBs8Q8Ko+XpzTrtXLAO
Eu83p9JKbBOc7lEyahDRj3vjLyXnyG9mr2PrE/ZoNrxsBVrUpD6fB+vfyhULp0U7z4KVTPp9blH0
1mtzrE/+gyJI9OHsk+gAJ3TV78sKG9/0mZyRTM/HL1pWeQhoniGB1NuvmAR+wEZ3pY6LD/5KnNHW
FjARI0rPBTImf8gKjF6GIiPaoRXwZUjHaWNFKgbuVY9VgIiq2kVyi8neo7RkYYgDQjf+01Xb28rl
DuR1v/f4rHsxtnFG0MTdMcPnvaG4K+37y410C/7DDfy3OgKdCKeANUcCJrbxAirI8p+WMYjYRgca
SNfJk4cdot/x4W4Ys3taFdAjMwvw+PgnX9O/QFPjn48p7+pxGA8iix9GGHsfbJYEFpLH1NOZcPkg
jskmRsOr5GnnKahBsNw2tPytB7nv44X1D+BRvqRRQlW154DQvbLAX+fn9BrKRp9SUXdcfZE2vkRw
IFk4KrNTjJ/RODZKyFZBEVDMFOvCAHG3IkGXiMZlnd8LqjFe+IHlv/XVcOKHU64pyt+lE9kO9mtV
z347KynyVxLV1WwxEQLYqncj5TlHi7DxnbxWJAqlecMV/XxnIRZeEOJjAA+hcma2oQk5yycDxBLa
vEyCfzT/Tq892no4FAL9nV1rLm0g5eC2ykgVGLDFRPKAyisVebfKqvMvpH3360vZAVgdP0+OAGmU
dczKOhbBbm77bkX802BacDF8vyYy+Xy9lyFCVvSIoOQJDGmJ0MnfyHq2zbclRJPesRY/0bMrjJD+
lbZUka5L3uoLFkp3phPANPUZuoffnOSoqgAeUeRF5nda6F9T4nY39TCBm0EKMu4jmUEvyJL2mYZI
6fKAAqCngFJVfwV5OjZ7HqnCBs9DdcQFI471D/vcdpvL8srUcNXQENUiq6cuH3zPxAn+o+Wrk10J
41/n1Cxiy+6lzHtMCcjlcOyMkNnvVj6Axdaa93zmq/p6qUfPh81QBoOMqlgR0ADHgQHdLX9S5FaV
rhoWL88FRXTpl4kGriwaW3h+ZOCRrRELcmBzKZMPyH48xYmlQ9Ozb21LdTzm40pLx38hKXXh+b4U
qyiA/pNdgBA9KwGGUa6iwOXiw1QOEazpqV/gwBMDWf/IOCFSCmeAu+T8TkGkXU+sk9tXuqUwvePg
6dTH87vvw4VCKK4wTAntOFBC5TFzYPGeOQKMghu/wRVfFDc9fUvjHf1qFNC9oJRNAgPy05El/HBY
NI4H3kQkNwK+g2Wm/Qz7tW97je5V2p+u1d6gZ55sSoFGKadO5V1NWfsoXb8Q/xVsollJFBEpS39b
E1v5JuGAuOvMwbUPFlDeY6FmQaahe+e91r8n+JdvhG9wrnqRFoxNrQR5wJlRqo6368bFK6UFAiDN
q83DDfTQDo+yXvivRtr2Ri/Hk18AWU1fFLfYD6zqU9FGu98S8SfjK/eoItuMQ56/BXXffeBLqmkO
KN1FmYgU9MT6/bNObaRBwHfzbZiRvdtaNOT6Dy+NQSe7bqAVzsfHh4uWGVuJWJa2x6Pucq1Vjb+D
t1nzpRg6q2gaHTv5ClTXTnam9BLYzcWbEY+Y13V1Z6GWAJ9+DgDFlCstGYI4YeeZw/i2jxQAUbC3
KC5bWWHj64AhF2wBUl5tNipATuqVmyFBUVIMx73ycd01okJ2ENjTt2OzoBRj3HYPJ9gW7GCFT1q0
pDgh1B794E0J+FRLdmsvK/3pdhVuGkc5iO3+K7uhx9/lMdc1mua1IAbCRJlHY6b+LUBmpJ9baJrh
WiEkcmfaGN+/QNHKFMnWXIGunjmBcqsR+q2k4COr7ADYSXipvKphTvIrlnzoaOHFzWjnmwy5CFib
UyLENqv8wBHJuRnhlnUQVIKQdBurc+CuESAiJhcOZj5VRaSj9CxhT95ADSEnY41VySBlo2L1e3by
B+QMqhroMV+SDbEJoBEkjhkU1WtxuUkbdZHKZrYWMq5gf/UYb6CUiTb4RPYO8ZjQCEir4xZ6ct2s
hON9S18y2HLjeKD3Jx9g1NtkqAqGz6wF9c74cyEDSe2AZv6CpDAey2K515mn53zdJtgUV1RKQXKa
FZynqZZt91+OrofciV+IL1ZYu+hVD0N7+X2///XczuMFGP61RMZy3ir/QjCcg2aDIVCx+m3b9znz
tAqoFfxwUB67CAGjweyS2P41qnsoGy7McI8gIjYX2ydcD3GOItkd6qKnvPGyyR8VIEQ3BGb4+Jgs
h+k0r/rdTLbvT4h0uO6W+Rx8yMspjCkRa7thi+4PoFFuCJWSxmSFwzaVqgN4CI9TD0wCwGgz3k2b
QOn7KvlWVLOgKWJHWzjcYYczQxC5go5U3wBraAZTk/o/DR8R8gDmMHw0xS95jz4BrgwrsQhtAgk+
LURZhFHnFZB8ohqmPo93EgvClA6A+gNNPPat6k2bG52epAGX7nptTd7I9XmLxeQFKSVekCXK5VV9
EhEoFPOao1H8DkFTqh80AMii78S818kiqRhHwTXuDyPO+6u5z8Pu190RBEGDl4oh8HLfQtKGO4yF
OxNcViMPoZkfwKE4VYpPUvitfXPCCRgzplqL+8/imIiEYHdklsfGi300UEkgmH0ifyv2vFSLwL+5
uygV5+xxVGq4JR6KBIuD+mZMNY5v8e9YYzu9BSCW0y7R6quqHVQ6yd7NPUsfXRhvImsycy1+jFR0
m0ThCn9Sp6Cbpue/4uIWHcofVAUljbwA6gMCuVwijTF58GQpt2snJPCGY5JGa0o8nQMQgTRK3x5w
NOBsaqXa96uiEcV+UO7coVZwVdrnVBAaf6UF93FnkM7XXtSkQXE5u+dVIQTbpj/mcnpLzvwnZfyh
i8AzIckl0QUVjQt3pRV1NK5hNuYmOajzWIAht43tTEP5e8evw4VAQL3u8JFIEO5CFzdoWhJ4MUSj
iKZyjWn59saqmsQaLSwPfGpzZhGe/mypw1ktXKxHiVxPtBcg1Tqg/fFspdMcaxQEMWXyemwtLWub
XzfK5rnyMzaGrUte9ywaqDDMmjGWOCmkxMnNLHezMsCqzSmqxz+7a9T7cV+I+iIort0NqNuK4L2O
pzR4w9umqAH0gEUaJXrhNUOeO9ISbiX5GGUbBTMzF34jC9Q+1ptXccLmDnvGZENfQ+4LcuxhQrsE
Xzwr7pOHC94XnjSdiSNMkkyoJVo4PVJ1DJX1t6PFZTWElRR6jXZCi9yQ8CtpPWSzNmv03EhaneL0
zcS+7FsA7Z4yQEBq5YtN4SZms9UrRC9YWuTdPUO0AlONJ9wx7MV3Wtx3ZpINV3COuck3I4QoVKy2
7tJKukAP38CHPCG1RhOQF2boQFoeyoR1v/7ZpOrWY3S8sm5W348cNA/ApS3cTTcsyPDcauY1Sj+Z
azTl9kNoK+hOfuVfmk5eW/ub7LcLESGCpXFb9jQKSdB2D5d51oYWad7x3vG1DVyYTr1SjrIf028J
Zp1PkRKe3ww22Gfvkw0fOW04y+O02tl9CQbQizUaSldnHff0B0pH4JnlHe2TzyMJ9nrL1oCTEBN1
M+sn64OnSZM9NQDgxqqHIbY7uAD/ZOtKQG3h3GXJcxVHLWtV02dB2NSLdXzYGwLtPCsLR9wAgqWU
bJnEG1EW4yFmTHASIPrXwsOEorXnk2gaMb1ZR28+y23PmxAq6jrbG293tM2XGNCGcw0zqhJOSrRK
kEQ0o2Yg1EU4QjOe609c319xZctGTFA5wKLOOQTk1BvYNDCe1DyhYgu02qinlExdF4evM1sd6NbU
f8nE2ySIPDCMEOdLY50Pryfps078GZ1k7TLvFDO/Bz3uJ9GpxuyCb/59K7dHFAQxu5MCroWLEPpS
PAKg9BcOtOSU7ZmyXIapBHt41Vy+F4nMc7V1V5Pl356nN0ga/Hg+xBKHplh7EIxyXtIGiuEOvC/G
KE55SL3w7MX3XbFDj8CH7jl5QOqYlcjfBzxcCEvxU6qseaYSnv09H2CaJtZEgI4GJYVepvs8H3nM
C+v3RoTb1v72Ut+mJiSMYAjg9qZ+GDJnCWwu5d1lWl2+VBFp37egMcSIBuNXGlUhT71hXt281cUA
vA4JJ03XBH6Xf7q/0x/+yrWOJQQG0mVllqcMjxvX2Q91HtEXLXwTbjnmyl4qjotX8sKJ67GqvbqH
pib+lEgwSfI8892m3Rb0M7LQnp+FfVZrHbCq0Yyn4ugeUNIkEhDs+KsAvrfd3hWsBL+hCJqtNtFv
E35k/QgWSC9EsGOdq69Mpm3FLsyW+5J3EjVM42f24quwvpeLKjBmcxSCfBPTFgF976QwSlDkpfRh
+4uV1neg1rn2CbcosENa4FbGMTVq7PXtLJRmqR1re0jBJnEuHxfJ/4W0PUHpvu7a5uFNheQa2ECG
qpcLipmr1/b63v7FDltgy+mvci8vOyrQY5SNw117CpkaxF8iXQoRh859kjzsgi9qQDBKosDN6goq
H7OFPWJM8pvhs1Uzsa0cAwLyn53jK5fRpPJojt0vLlUq7MQWcqREMx7Lnm/MjpGpsceh4G2bYWMX
neKmW6tJyZgzvpdxa1FUDAwPCgvIqExBJllwVikbT4eFbi30F20zKSKg3zlbd1zoQ4BprUXWm6zy
rUN0J5LUkyoueheAMmd66r0KCUpqoc2TEea6VaTkEEjbhmP6f8hRv6XIyGcS/22GJGLh13JT5bAh
tbhYqHrJdYNgHHC0i+CTRlIkKEyLMVQj9OY35TFfEutRLbyQhGqEHorPCm1uT75EvbG3wLDiUtVF
8nNmO6rRI9quCpyS6NVIq4YaTBvNLkz0orZg1PpL5y1Kw1PYGbhwjp3jj4KVIyyi3R+19V6zQNhk
hlf3mb7oSzMjO2jPc0SH3pEFiiKExWdaql+mXtxpBwJ/2Safda6Jyy8ziORGlZMWZOvgGdA32KDX
CeM1btZZ1kWbtYgyFQRcPsbTvjqgelHTgG3/WkW1kyuTdnzGKaeTHuNbII+TSZ3vZeU8UOIsKLL9
VB/yZ35UdLxuArTkNPL2xB5qZwd2FyAUP/x04rZ64M1+Mf0wGwWjmzQ0MKQ5DaaTnMOTb7JIS5Ik
ajwG+Xp3flyWwTOwWgCAboszezp2dlAhYh/SwMg9m8dX7buP3Khq2rHBVR8H5k6yss9ueWsYjz3I
QF2yLaFo5Phrjp+ZDTCWswvD0lcf3VHz7x8ws3zZP2nEeGXsFffubtIovN4jg+m3146fxeOF1Zve
/y91nk8LAp4SaBQSywitxjs8XCDq/E1JvrSBucavoBjKTlur6Ve1WbgGPuN9/fQnQOHvGqaOC8II
43YEJVWUhYB6vbUTsmnzhbu7ICz63VoDMxVkxFXRDc8HqM+C6IImxZ5TZv8nCaDxaAn3A61pNnL4
AKr37bPktkIkZKH1RBvpB29QKNm8c3snTl8cIX4YlvHW+4tnsSolcNR6CkJrldsQ7MBK0bXOxjBJ
jj9hGzo7J6wEmh8h3xAwGZD5I1jXin0K8R9ro4UG3djQkWpS5MAkVap1Z7srlY7aiw+/ptkqsUuJ
cM4DWRuVB7GfzrU3UeLgd5msM7V6XfeJrag6axH2AF8EpCqNLPg4guVjz58UFOo57827NBoPHqSi
9emlRV+SiWFq0xsGyHrV8Q818pmgf1iNZZiFY3F2EZPpWuZYOOS+LWBoNc55Zk0D+gVBTkwsKarF
0na8W7edtJ1MqyqZS538ucOhXAkvqVK+EZxa0EI57rfnyAtqMT0tnfZQwknVmGavLo8aTeJAmWN1
AA1Ap/+7AEnu06mJsyK2I/gMsradkdoJLzAsLnFmea5naug4t0Bpyn8Qix64c7HO8u++2/MJFGWJ
9wOpRqmFKSjvJ+jQr3O5BNfPfQT0C1wzwbqIYxLZpGRwUZ4eh4n0rgj6H694lGHeSvu12DdABBTX
mAVSGaWZc2iRqp6xiTkI0KG+YepiJbJ6WpZu6Vz5HHmaQCVQHtHBq7dS8Eji2a41ubqywZpajSqK
q/0krRfaYPQfcUmF9Ni2fP/XHcApHeBH4u3l/iiQGsPNMjBF24CW9XjnTt3NTD3dQr2u9g7iNy2a
J1TZ+HSIPkJX7QUN1oe1wP3IfpepJ97pk05NG9tx/uJ9P0Ymvq+Il/0becnM5vlHA2x6sVcbeUkI
E9lammZr9Dy6wCMVSicEqbqPIHTQf38gSoSqyFAa8INrmV/Te6KOI+9C2UZXdjQ0WxXlUxHEFvTn
ZAAVeAojqJ6ldCkjBE/XqPUgsXp6OVRIABW3XwVAqgXqUSeACAL28ItTB9E0RQl7LLsKFkA9Ta5V
7xbv+tv7iSD59jQiq/TkuW4/Mxmi3QJBJYuWiNXHEG7k1WI07fB6NkyMKZje4gx/3nKOj9+VegjJ
Mdgyo74b9lXXMUviOnqOqWCpuaqxlU7nPjhaV+IEqyHRgdn8MppmSs7RiphtfbDNWVQWh8hs3jLZ
p47VgLUbbjzkFbpKHDC+37oHJtqmgCdgfyLET5ifPcooR3Trezrub7UwifMN+1yeW4p6IaGrqa0H
lu/nlJ5CXfwKfHGddXhticAFEktasvAcyb9Uoopss0OS5xLa+/h4MVNPTjgyrV0nG6WN6BhBDwSg
7M0St9h1PvWicLKZ+DGXicZdaMv3q/glW54XNd9rHcCLB0/5NACtP9hLBTUlBNVEOQUBFZtyJkgk
f5ajJgGvpDmocMfv03oKLUDPW+qf1jnHEHTtXp5HWYbqzdLTaM0ozQh7X+P+V9TbpeWxbONcHEgZ
CMyhDgLyo38QIBQBSS9D6sbxOfr7hk+Q6Za6jq2lhCNKhsrGFJ6Jm9yD2SQWxuu/10x7Uy7RRR3g
xm6J3WVoWynu5m6pM1I2la3JPcxHE9HJGTB0T9wIFwFeZUCzNw204bEePqTIBAM7dZqWuku2mriL
QweJUCeWWPcgowNdm87TVOXxoiFsQrB06wmYWGXuhwpgVwgkEfTa24BjLfMbKsMRH4m9ilEHCB/8
RccLm5ZZKBoW47xfZAV9bLhc7YP6Gsm+VrXBbP1ofQqBEH57eqN94BJOmyF+LRxcSRogr89HiQd/
/NoAP5DnNmysHnH8H4l6TRmEuuEe05H6bFacUNctsL4s7O4WgiJR9zLoktSaeLtbs0IJsXVk6b+U
wC6lU82thlVAFfMgy73rcyiCoA0udazw8XBNi4NIOaw7R4Vxxfmud63qrkUxxbG14+5/wsmFHwts
8A8caM4Ah2pCZMTMaNoaJ4ETG/+3EE9hN4jNwyO4bvj8/O5KDN6jBLMl8P9l+DB4KKBxVZZqPcP0
uQyIqfkLLD/yCIVVxcq2CBWtSU7kBAQb/047XLbB/L1dAhh+MrzavBaEvXrGf74Z3SQ7NFTOFFgq
FSI2ytT4Vz33KuMnXpeHldfh6gP8iV/y/l0WkK/K461/pCCTXNzQxbyPhkQtRCJrzLZ7xJ4UEEsE
YL2OKmyScJvW8sFOZAWfHb6oGyYieup3X7WAhupWga8YvHfwiz+Ex56wpYxy6CmCZQREC5SRb7Fh
DVv6XXr30D7QidlIDurGUSVxkuW7gA2HfMRbyFNIYP+3NKdD3z5R1f4Rc/MyGSl8uxF068E2pgh4
NrRXMb9gpwZjcs9BhyCu9QnUNoW2dTv2OIGjfR0qKaosgkf5UjsqsX6M6UTMv5tO+dNrg1WedExP
dMJJMKIo/PyeSP1uo2hX2T4HOlf5GvwvaeKyQWNsQRBp8aS0chv830KTi35Dep/fDKH6gJWuXplV
bVJbocyE2EGCSGVPDlawf+tMI7mdiJ+RlUFuHDAC430arNBhAssSKQbBJqQhpsX/ZIR9G1amjrQr
10tSxRttkSoYYnT/O436cDwH6AuXhTURizBouxktOE3H1UY8Us/v/yxc+7ZqiVDABvSXXXZbX8Qm
nXOtrSlxdhCoog4E18advKAPl844LtR/R0WvuiYCikrqXuUSihk+QTuujqyRW44KugaoRY9303ye
RGPTI4rsQQW6mYqU1QG9uN5lol5M8tjQZ2X+9ZkPwKE2vZgx2Gc2RI4mnDmKcYHpkPJMiosEEBqA
TxmYucZPLuTLAKy7hFh22YKjoP5HhvspTklpl+HNJjbJ2rccPpwIY8w1+hl1T6fX2wXRnCB5VhOU
9luh4AIFQfLn3nwCEBITYFW9vSSElDikPqV3xHKM0yVRumaAXdkOp0o7TlWCcShqWrsbNdHp7xRJ
El/Nbpk0tCCQa8PwpgnmrP9NUl04Eq8I/wf27lo7r13ZZXz609fZafJD7fzzGjv3omBpsm/PxdPh
mElK88VbbH3WBJr54BQxchM7OY7XPJZQRdVv6XD8qyleIH3X6OAkBrR07Q/zRPjIMJNTSnSZQNuY
cfwmrMgjOFLXcZlLV9RIo+4k4nXN6ba1XOaoWaO4ACPLwZV/h+iqzzQRQvTeOP7XeWaWdH+00yWG
ap7EmuRW8/b7cZrt8Yp+S3/nTTapm6YbLjKRQSb20Ktb+SH1U/nS5DPYzJVMMv30D8pdPdmPggGp
aeVHLqRIzIwv+eb7NvtLSQzj2mTInJgaqb9smMETN41hFkDpfxus4ghbiDq0EUC9xJNDbjpR+3Ds
Y1qXX4ku/JauqkZ06LSlj7gBgRwG2kQ6WS1z8Jt/U09xnIsQj5gVBLGZvP9uf42QEjmg74Q8NI+a
WEn2jDf+VO8/pN6HuqgVPRwB3/r64W9x0RHlAmjpjA88Tz0vvDJylMJgLUon2OjYdJr+kfzwDGWS
kQ7ZRXE0r34lKP5ZhDqmKAZIuUbpdpJnoHL8RCCXtS2UEWuRbt5U5TFBTnFg+go3en0ESVux702R
cMXwR1EZQLQnu2wIYOVGPYkkaP4KMouFwM7qvZn7pzSwJ8XlfkmxasxabW65Yp3y957R00OdlJwM
mIHKMmSqWNgKmOYbPzslwMilZISOuF/X1DBdzGHkA54YLLOn2rjDW+W8QkPyX1XqQv6mkX5hOnWu
dc7Zn99eAny+eNpqMM9/WWnY0kfyBwccE9df9ZPKG8BYIS0WSWwJHop4dKQePgr865Im5W8EQcCd
d4xGevB6FXemLiJO4OJ2ZhHnvw4hiOcI/F3XG8bBFtTJZOL5JvDJpIu60mG2gb0rUApiJV/OWphl
VGgzZe6YLUQPSPvaQbXF9qlZpLzQuKJnihUad1n5e+7bs/URtpYiCSPN6sltIzFlOKA1gU0L0EhD
2q8IUP8jjNc8AN2TnrbDOeZaeGCS1q1QHQQvcXlfYp6OOyR2MS0w0wcK7Iy9sGZzENaIOsn7yWcd
tuxAI+hs2GjijXAyR+Gb6pQCNPsr/diLzT8HBBFcy8Es4PRIvrd0GsPhunIudYNrCaj3L8p+oBdr
5p7X8hC2BTu54yKhjbvioKwnnKC4uFpogMSfaSSikHRKDJk8v79eThtCUyPIUZfHcP/gAbUuQqUl
u/hyEB2gDFW3/38Vh4VtcDDo3uRfL0Uq3klWy2JBHq0lXCk/eMSkiUJ8dN24bO4wguhHzfw+e/XA
sc5rfkYfqhrMJtBSiA55K55QD2Ev56ByypfnK+IYPbHFKYnC2+hQl/rHvSjrlBvTWxNKKOPYHYVT
yz6iOjArC+TlCPK7UNJqssvVzLa0swdd6SATkdrYCJk3XRR5DHwwpbRWophgR7WE01giWFHsXtgu
ZLr8kFrfj1OKeDif+Jhb36OTEErJ0TfROF9pSgWQvt5lNAHve0sWKyRTi0PqDkz0flcPj7b77dyh
kSoSAA3nCV7ftB3zQvSRXs6JL+l13eCcqMC/pDzfc10lb9NnvL0cvNAwthpS05TtAPO/1zz3SkeB
sOQ+9Pwi3tO3LD58h35j1OUaPCA5+DYmmo4sW9GjxM/Z4BueT7EZjbTFjQblUKRJqxUFoX3VD7H+
qa78webu1x3cYgNlXTFPZIkR1YypsXa6tyAxQCUQRgTGZVyrfyr9rexDpOb6JBlx/bZKQfTbE+vO
X064UEZx1I5QOt9/DbvCPp9zqQ+0/+VlGqal5MOF1Lv/0WgjCnJ+Jgb7kZF2Fqq46hatQYPShZF6
fVH9TlU1hsdKoYCjB1otphNWeJmKJllBm4kX4JmpL7AUNAY3pZsQokAIcRMEdGEPC4auvRgztkkK
z/RuPJFfVvjeQ6v2DlyRWexb7tLtdn1rrovJ7zr5y/3EOYVN1ilpIk0KcFRC5R31zqdrIm4J36C2
g2zsd7Oh3ZVj+kYcm7h+TqGeGlKVeRWBtbcr4YarQlDGTekom7JX47T/tPhx8+BoiG88uhDbxgsc
yQQtLNF7JGqR8DxsHljAJsJdCMlpsHMIgs1q7y2AaUKDvglPnJLz75+vW7uc72QR1mjGeFVxN2jc
moRdApUFV2FRhAMUL4JcYGU+YRbN0mNzfHSQi1pT+JKGXvnQkeXy8TOvACG3SEm0uxCgo/7Ymxlw
H/O8uWW7wbACaCS3e85v53OF9zZxE1SiIhN95qx/c82LY9ahJUoQqNYVtlxrC1jZL0bcusAkUuXs
BjJ+UzgFuOoZXn/2FY6MYPlJpsgult2ey77H660ZvxDYwMPYYck/QDxoXH4kl8puXPRrXvnFYL5m
ZL2vx7ObejbDpHHGNDnIYCEDUSu2AaHS2ej9p1cMnya96JVJwAVHPC43dLUnGBNJGXM9AcYcEJK1
+d8N7f17TiudASKGB461m1XCFsCd0IvwpzrAObhtMhA0qwJMpf0dnda5bAzTlhKsKCWT4Z+jRiuX
55DnYxaJh7N1trll0jZCDZJUcSpO1ltvEGjte6EHP8jYMDrPhBVe7th0KxbSqlTeKzNQ7kMusN5O
9HomVDI1rj99YNwITY4y3GCHbPNB8Qrdt8livwmaiJWfsbks2thdxqoT/hEg8UHEuIQFV34yAUwF
Hjufzn07JHzieLySWGu7hN43l7vwLEOd/BU61rGJz3AF0SqhyS6bWq3nieu0/SBAppu89B+MItH2
7jzlSD//AmzNganWYnQpUkC5g6Um8B1kyg5MxIZPYLeO7wn4/DlaIb4X9o5Jop84xMcgbLtkB2bx
vppLV6A3j2u/lw+CU9some/wVD946qTiZ4ADmcRDDxh+D/Tloh6O5SftA2kZDXYctxt19dFITKly
UB3aWAI3+n1e7MOXbGXLPLijNI+I02UEYNIot9lcITBn3ArsythWc9Cp9APhPO9LBpOpFQOMkg8Z
zjqhy63Gjp9J7umI14xWEtmu4c/WWxRGE91VC26BghbBGWaJD0P2Jy3sBU/pmf9oUwpE1qQGrZgV
9CElbEhRN/iSvbairI4vmWkS92CtcueQO80OkniYzP9kvsOOJyhmfdRDvDV+rf0tit9qGp+DNA4c
ixqZ8e+Lltk+NcDF11jwXYbz0RcAvS5slpd9lBMPgxHr2mXig/wVgS6VwD68k5N3ClbY65Uok8LF
OEGPogutZbJ1Qeyi0ab6TPtcWxyinx2L2+WkTTncSMJUFgqYR5w5aTGzNnTUfKyCSeU8KaFwS3XH
W7XB+eMzbKslUObMqaFh/NFPiDnICxj+ZqUxyRA/kJVJBikB0DyEVP7QV6jAVehAHCJvnWANL7ye
75oizhECYAb9l46IAGxu+R9K5RRgUvWJhe3oeVGviCtasdlAH6izehGJ2gaAfU3+X7dD5ofUMcGM
p7ofB3NCpyp00fvleBUs7K4V9iVqhShT8EsNx8itg6mBHyNFqhNP1sf6VDAO58QtlKmBFvBVftcV
JhNS5VzhCt97JLTgZvEUNeWWsLqi9bm6XMlV8a2yxyOkTc6pGE80NghiDZPnS00N/N8vMYs86sQK
7HvB2S+dr+I9GbSjEXAnNz2FCYLSmZctGry9pVLeDU4BJHJXiDYC0HFwJ9xvXtHWCGldX7Xy6K0E
kG21t4jVxX5Gs9sYZ89kldcru5BvJ4EpE5p3eJMCVXeOFLM2x0VogSxVouB5htj6DNIwY3ulsFmA
pYBZX+YzTWYCxZhiRfU9aP3qlXPIiDTmAAwcHHbDj0WJ/k2UyvLFam8wnMBxsmbzmGsZ0rx6x6VH
HTC7iQF3344f7cez1tGn7XoTQQwZlQsTfQasXtUzNTqjm+4tg/EHaVHIseGF3br5yyunJbwPpmzl
HXel6DvyMMkvAcNVu1OPlsGrnjvmA8TIZH6rMK/wGagg75WgFTCdXz5t2PQrqgU/NBLJeXYmuKZZ
zQ8UJu03O79ppXUi1g5WVy2q78FWleTCPDN7Lfpf7AAutHFy9V8pegKDEjfENvEphq+TIF3AxUmi
+89R5QyqQrpPlckG703WtQKDuzDUDSitbZEiM+hgzOS9vHRkSo/MlI6OzNHpFNubq4p2C6J//hOF
l1zs2iEYN9BDlyLQxwuJQ5jQ7VVwz2ttN+zwsi6Gy1T0LZLGviEqlJEAMTj6bIC31HYTCJDRVO7M
Q4UK3fa+2WaFjZeXcOk8l2wI3mAlbiwowpaf3zdGxtUvop0yaLrv1cnOFy7lwwlNzbfj1kvIUoyU
m34/9EgcQR5HBQ7zohBQY/64Ok2vC4X8Z70FUndPCCZcdmLZIwHCWka9TnvjTEi9RzkkzV4eiMzC
HXs3uAjALunnEh8oGYiqdmQBH4ecNrRvp+Ao9nP301rJAfI0yZ3M3iJKfbVeDQJ+MzSflpI/F097
1FnzccfzaWGUOoMqe1CTSrAuT2CdkiNn+Qe/L7UBaLvgAs30ccb2XyqKDlVpjTajDB2igIkDhAmu
DSsxgmZizujxn7NRZYdBrdNchyr+sbx/aEqP/QqvbgWAv9U8SEXFvCnWnbfq5lG2vLtY+LMHp08p
1ePjRrc1rZ1a5sCiRA5DB1jTrH7Lq3x/nn8jYxamUEijUfAMBtvhmzg/MDi1AOXXh8Yqgiq6KCUD
8q2PU7G7DXbW1aJPoBJoPsLHjt73bIo8N+Yg0N9nNXovX+HKfgEkXST8iBrInjfr5yqeDjKSqWG9
1pXUOt+FvYqsC+iDlHZlxffCWaAXgkzfwadduqv/gmpTAuvMfISN3c/t1nr/Kxpw2l97NjWxotuM
bRMMSzAYJdVYwg0mjGzSqqOF1vDgiKStrUS8BvqcorYtayYAuZgxm/EPBOVkqiGk5qUjBdyVits1
Oe+B80Q9sw0f2WnW/IvwEAt1kPciQvVsFwc6/LvZsSf6lYWx7I0TK8gr7Ffhu/4mL4e4ki/k/Qoj
1rtou4veB727ybbwBu0z1xcxfFWhNyJlsyHF7J+wFe7XoGkzp3R+IqikeVsPeGZUU6XenyOMZpDY
zuVxBIE72wSp9a3leAHZH5W0WgTqmsqhL70yuB1aaV8gRsNS2Q0QM05Gl2wuLjbk2Prwxf274axo
JMPRHjbGmejIas+sSsk3r8KKzBxEcRIoUhMcnItqyI8245o+JwqEjoQFJxPbq+SBbLn1duWCSJTR
vZxrvIOreAPzSsQjTrY1lbU52jbsa3c36/TO2+iEDun39hZokDzVyQJZPdsHbmah7jwiYSesDwRx
WzOE5LXc0x+4NBMKJtl0W+yJ92JgBJm/luoDt1Dh4BKyYvzNtNPSBGg0JTeu6ryo8T8nJNoWe8Pa
vlkUPedts3hPvqU5OvrQSD14lDxQBgB1DmItB+Jz6EW1sCWknwceJYDujuDbOspPFgkfvYnoyTTt
AiuUIaf1i8mhOowIy9ed9G5YOvwQDDWIef+alvqhx8FvB9q0dRWEI8fSyznobTKrFt1HcPSWj0Kj
8sk0n7a/g9Tpt+ZSNcIvnxGNsD3GVU7Fw6OAlnbDZKoPMLPtyEk0Se5ilCKphIENJoMlG/ChlI4+
QBYOfu+b0qrIzCiPouZ1Tmla/Kq4HppHXVNYq9jFSl7nFVK+GjHfULmIQ6aehDppqHd8cMBV70uA
Ik8bd3oNcOWPoM+1/D4BCod4H31qk0hSirCSkszuBRCvk79MHPQjNMIexNfoKkFViLCoy9MWqWNm
U+/CsBtbKTT8eOoSU22tM/jxuuUa5QspCcNN5xf4JAcmlB5ysjhggkhc7V8IEJYed5+5RPSwtVJx
NWqo6VCI5dlugoRg8Tiol7AITHTsriXfHNAqSEJmH6ptbr4GJoY/SaxpWJI8BntzdS/X3QjPQrdz
AChVOOgMbKq4G3ih0ewg4h5XH4CibAs8VYjNOgBExjAH1Z/nHWemswv+KBnBOp7J3gWPi8TRPVoB
plTx/6a97oZ8RSwsg18hwaqUe5RHdGdLGX7HEPUzeUgX7HxfnNI77CEA55ToA2GevxhdufQDCVud
vGHiUofouifMEffPwZqmK7Iq9WG0r4xc/cTBZl9bY7mRk2MsO3LHlEleYO0UBwVBN25gtzr6IKHz
Khb/5mX1tiGZtV+/udIUAYq+Dg9WcDZDdfOhuwxr4u3b36jcWddxIu9ado0pVZXI6cpohZGQl5aU
xWxLO1kncjhHVo83LRuJlPHi65u+x1Ey+JaMz82Xpr8AegJzSonPXXn71FxxQWkxzhlYt1/BQpbb
S8YEJ4nYujsF22IlJ692a5DaQvFcxxWhL9GowXLgl6al2Mt2hl7nXgz3O4qKQnnuSvcOzWYRBhi8
gFs5+j24viBx1ec31U0K6OYbYb0Od05toc4tdKmmVFcFdXmhixtzvZMqsUAhZ99FulyvGcQQRKvl
fZi63FSuzdrtH92gdwkJpwJMvFZ1M5ntb/jEeke791S4r08YY2xUyljShrORU1C42epld+ObsOv0
jAkwSAQZl4ow/Vu+f5oxr0xFeaJQ2B9cz7I7Hz8Nes6ZXsFBz8FTAAI5yjHTM3GwxP0IxTMMWWFR
sLFskzRNq80dXuBKAo0nV8dJ+YS7EnJHjBfaTVIopP5oNToB67mQB9rxNoyu382f19FVvb2Un7BL
7V4S9F3pLI+r3lsoGeHZu3KLH90rsaU7S9XR677a3LkUouFe8TpnzPn0CwgUhIMmA2aIu0fDOG8o
Ko9p32Hfv/Lk1kQMpmd0EP8ZR98pV+u+rOeCdEjNlno88UYgF9VLpyqaNq5tOiibuTB0TA9IdvqM
2TA1Q2jsX9dd8p3GOHFrXeZOaRn+mJRM5xL8RHMfJ2dJBoYD87BcxLdM80MaPHXbFr8aXolcOQV1
/fo6M6zVEEUy8lCxkUltLHgUrgaOlC52pEfncRZkAn9BZ6iviROdt9cp0HI5xd7LoACLQhyFGSoS
iIPczRUJBveb7kQxV5ffB/9t9qlQarwo7XE5CjENJoOMQwJpubGPetghfUIx0xspS7BSraJzVudh
H/5cQNz+BpHXtGV6hz5FXMly7FfkCzakRoo+Vhvcr8iZp9XGCE4xNdIiRoEN9Dx00SNOjqgfoA8+
XrFfi7+D/K+HQePzWOglzRHYdq88GY1aUoqM+NGkzR7HP6JDFKy8L0o2bdaE3ugSPNyFyhmBtA6E
BlUO4bkRZWLdyCe+5rLZ9xzdC8eR73FAeatajki6M/ZmfwfTdV+vY8eREFVX4leYZwujeMW469uJ
6OdChxPtHLRFp6lsaJlBPJULH6PtIDzUBKa4JxABwtLQUyU5QpbncBS9kj/eUPC7WqCtU5DlgyfV
UmRiISohGx5TIEu0FZuPB1deEy4toOdVv/sy7owaJaUrvu1niviMsRV6d9SGeWe0QcgVda21XTMp
FxONZjn0wgSo4ekg76xA+6OaA4ZQ3/gixWqEeg8qb2zvFqiDB+zyJ7f/gg6kGpUHUvt98QUvI6jK
aMQftimlaFZR2EU4nL0p/fKrY+DmLX99CP8Daa5iTO9A3wimvZa1lE92Ky2NKmKEaNzfKM+gq2vY
7bntbUtDvGigV2bwNtGJPBu6USlnPplx3qdD9pVp45Uq1eyM2A65BUXku/shsdx7bFufN1M1tSf7
SdMolmch36GMvzjOzLYr7pVf2JbXVLrPFHksdjHGQGENt2xKUKQOrogldmT+MLunnr6g/to3APM8
1sFuCGwpiMu1FpJI3J74K/ojt4areYSVC2dyKmhEuQJCO105jdC1qLE+YuNjErPkA0nCkzw8mHI0
nyQrmnu/k5Fw2uhwxHvwNBQY0IGNRyAwvqBO4rS/J4yQYUtOIhWgWLLknhESn1B9nb/biVFP/Byo
D9sAnK4K7RkMp3/4KbyVWHRMCovecQJkd8sW0bPLPY1oiDZGHzLWMJM22o56SMYLHz4I/f+JkcXx
+o28r6puH+tT/OyS051t0CA6L3sD6WULZ7RqPAVD1e4F3QS8iH3h+gvOnCUeuFP0tnX0+hOnGVps
n7odpLNaUX0T6H0L85rpCTzJLwPXaY/3ipP87Hhm2NbhgOmG6a33P7NwgcImLef4pjJsSsF2hNx4
ikXFcBliwdSqpLj9SfhSphjb2FsEdsLxSULiSaDddwmeNxj2QfzI7jsGfr7s6wubi6osWMLzyejf
fKbGwZ7uH3idpD7xb+RbKt4v627i2nF8qW+d1p1uNWhuskcNkK1SEp8LdYKeeC5k3t/4iiUUTc9U
h30pHnD/rdqpvJaB3Z1YeAY4EcS65DOnO+jZNcqSKlpVdPm2ByYHFkjXssLpX2pu+FqzGy9IDI4+
uEHUvyOoFOB1NQFlF1/UuiCLJe5ku0bpqHEzFAzMdvaCenEdRVQR016kW03Nna1AqNC09AoMeHXP
LR7gimF8VBNWZeB85+sL91L6jRoifYiPT4fZPN0aAKTdinLB3GPhEUo+R3Sfy/FtFreQQEB4E6Yr
KcrYddfj3aX+ImLwT8zHoAJdRU3meXtBOLdVsOomogH1KD3I7mvPa12AFrmjRYg1ur3Us9ysQcJv
RatYrjrIRkb0hp0iUMXNDoI3lWTWlbBAb8yGREij6Xd21WwIU0f2+ty8Z5IH11Wr9VwXhkH446px
fmQr6/7nZ3Cu1l5dMsPrQ3ZsbTDJ+e9aA0cQwcLqHle27faoMtrUZYwcI/d7fTPLZhB5S0Xx8r8E
R140e7D4r3FnIm/ZGq8+TqntqxzJ6r+gF/NKC8kHDtIZFmLPvYWeg8T+qfgXApSBFfgjtgqq6zNx
GfBrlfAI6eElBmRAmYukMfNIXtVJ2quIqJN22IN5SQ12doyig9G1Pe08I0aLZEs0P8gbgJq7+kSs
icQkKuqebDjawCtxZfmbqceA1+ttNrBB5TGMXMRWiJA7n9ONWOOOo7bPaK+fs7T/tExmeIA9qF4Q
x4pV3DGZ6OfCsbwc6gfzZOwARe7JA7JNAW2EG9lmqcf7jgW34Iy3HPN3BieYnQad9lBcNqGFKQQc
1EDMKPPBg5IVWYUKE9f5HpX3u4Gv03CEw6JpvFF2ClVleSRbnOUv4n82HTnWv7OAEP+ruVsaQK09
RdL9og/5RXczXc4yzYfeLCkn5Do0vWhPuZqu9QEE4jDxBNo1f/HyvkkGMBsG7PBqImjgM+0BM/e5
OafKKCresMXRS1whrBDxjzHsuroCSDJZzuT50JGtqSD7gs4d2Lbr8XtwbzqDicFe4aD7a3xKgRN+
K/6n33pmQsFRRaRALJfIotDchyQjYe9LPEGvnoAsCG/kD+3wVaWhT79iA/3iMoqkwJtjor1An/Ez
/ATIaX8I2GHWisI81GRDUdaE1A9JhYGCg/M22aYRELMAoHbh2NO3XBzfAxvw/5E0ZRjDzmGjkdfN
J4zRa2XgpcolwJvWI8rnthJbDuRb1BDttwSulOenyCL/CcoGIEKnFf8kMdZwxvVAcVkpJ16y7ccL
oq40uriKmHQWYEamDzLAsSmutPwJmXQYqYweisE9FcWhOUx7mA49O7SiCjAFQaM3mOC/1hZH7utm
wwIe/cMKJjlkFnQIKUa+b2x1VbizOVGZhmuIfsYVO+yb/8O4A/1SkHZJh2S6ayvcUHvOY6/c9TXm
nqXVkCgm+bv4ED/6HQex5oCktzKNyS2LVcAvcQlC9CiDsSF36JZgwTnwC6g+f0lizC89yaZn5PTu
Q30SAurnNXi/V7dGQIOccmmMsEwyBaB3V8pbX4ZKsksWsOxPjNPOu7M/Q3MZHweEKNpnz9JlGJjp
3ujCmRV40oWnCM3blxwAoWulNWnvNyav20iC1zAp2nLwIEiwglD1OVfKrW7rhsSvG6kxgBp2HSZS
rP4syf6bZ3NNqljzA1nwrA2USsVOR/upfV5SjgEFXO99TKumhiOcmzK7ig6tFFj5PVS9fS14xvwv
mMZ22SkGuB/yirwXv6ijgrIic2pajjxvAPRPQjGn6IiMbid2LCbpFjNeZsDdNN0VecPo8YkBuNPp
eFhevcoeT/XODbm+sPqeTbr4u+EWthcyZE/ubQJNHBeq9Y/J27isWDkNwUgSooNVAQJr4qyNuXtJ
HjVXCUz2dYxmVu1nB0xCRAU1d421fSXTcS8AvIbIWoWHznB9T4sonfkaY0MxOtQe8w4Atomvm5rh
a77qLU/rTVGC98PrSqHudSj7/vNTIGRL8C0UT1e6gRfwsxjc2D9KOZGQIk4sEdnGmrvldJJpYbkS
gkyTCVNXNAMNr+rS5P5nhq049qiNM3VbPPL4sTxwlI32Biefm3ReVDccJdo7XrBNYlQhcgYVGJLu
W8yB3wq3lKXBSWgqNzGiuX4M+9xkSWCLPIoC0wG7M+ITTih3nZSqcV7C4QLya0uKRCXYs3QaiosI
NodM5TxozsFL5KEcQ5mCI/DMcd0fXyjpaHKrbaLS4RcA0ofyViJXGBmLJaRfivOEUov7mpostiKt
U5fztOiZCEgoJ7LpO4dSMBdSBg/e/uH1UzemxfjAOXbE6zQpSdaemNyGbHvefboPf0tOkJVt+gh1
p7wwBc8F6+S29zyfR/etA6P13fymwKo+GiShyW8M0WGFesQJNGVXfVPzrdfctzyccl4uzgfdvRqx
rWQ2KQTwXYzeqtZKqGwASWNfK6SXHtBqwKqwAyrLxOsgw22GEjY0XkV1+tmedGYadP7agTvhuYM4
Pv2ypqdHA9LpIwiUVHc/dKP6WLql1D9Lm1VLZYAXykxzil74++FR4UwON3QP2sokfBB6pDKRcfkS
EU8kPD4Mlq2BJM8RKvdbq9VuBFYx4mtHyLiKfW/teddOEsWrL5kLLGUv81cVhp9xB8dN1Lumly69
2ltf5gQbTnJaLMS6sLFLC1B10GJoKUe+WTiUmHbhhyJNfQpdomYS5GXGlH1aN47oXZ9Lhzzbg9FL
a7+NN9dP1N0A1bcM8BLzCtAzPTRnmkIS7uYlLFF2yuJ1+7kgOPdgIrfU1Pa0y6Xb88M7qEu7e/87
ekp4TCN8SdT47n59pcYfDU2QCgrOUbISKIJgei0lwc3Dl0zmku2kaJpwVd/+lvYad4WDXE1RkwDO
LGqhOQZATO1Q2o8Ht1y9fUcyB2Ktj4Uoyu26LZlM85JM+f9abROxfGHr3PpMOP5RyegCjzsXQciK
w1/E0rmQthRITeosmI80xcWrFZB74nOEsAyOYXXXhMhJERXKXadXw+QaRII+2j3oixWR3ISsvKHh
PAyng57mBKXCEoQVWFjrdVAbOgXA1rSAU5P24g+UMY0l2AoGPUZm63CNB+Ly7YXYhnwNMPXum75N
AfLHi/PNhNg0AoRrs4yo9MY92ycXTjTKF+PXZ9Av3IB7c3WoAQMmDfGf8a3PlYfRwNsd/R6js2gP
3cxe35YaW3YhuIXobfGNNVCpj9aMTsPywBSw/2CBLZnl/SWqXTlVWjt2nmTLi0Mjho+ftZbc3qr4
tViOqqOmJhPqp9aWNAVseV+5RHu9f6RnkUjdUWGXmx/afEHa9YMPObdgd/LbqwyJuF5+2IyNsfb+
W9aKmDyzsmT9xXsvNCl+BjPLSWquxDUxv3WGlJGZJ7856Ib9a4S63jZgZ5lpHHCuUvgYWTI6T2QZ
DnLTLXxgCFZTZ1r/vgTIdWz6kP7jUPtlWt3ph1qXEQxoE2egj5To/e1lcmE8tP4bH3vuP+A4w63T
OkZZS9dYBaXgDWt6SxC91J1w2Vy6MKY/pJzoY8xHh1cqDB0Pwb9BSevLD/KwhzohOdlaWvefmU3a
/iBY0rBB1txY9Hwi8IMGnLA+/FYsyw5taOJg+Y+9LkBqQKT3XLi9HPDj+TwzReSVsBWhTI78PI9w
2HS++8E8vrdBZ11AOY/DitEZVOeYrMUqdq+l3cKhqP2z5wxgDj6wYp941Sb+TovAfa7e/2GB5Yv/
Pq+M03Y9UAeYcnUNTx0Y1QL4THgPrfo54QyAFu2PCg4Hwx224WZ9huPDGO8NS7Wuqsu0uyr0zyDI
6B/NWoh+Vz6eromdumPtfr92BNXRAMyBtiAefjX7FUNE4WGm79eJBpQL79DobB6sE2qJIslU0ioa
GbaWg6U4en52jjIWfdoRsS89iOmrsnEdgdJtF+GbohSCpJN/bkh/RJ4TtcdCBa/b6pqHM+a98EHj
YFZUqBSgroafrTFRsU+yuqKAMRE8P+n6MdpT4GWHsXAZG/eBAkExbNvdV8ukFPBELdmYKqcFEiOp
dd5d7i9V7swNId6WYTNbXSCWzRCSCi184JSqTl2krhbVWPevT0siGhV8p9kvIGs4jT/ltnsrmgB3
r7K93Kx23IpN3dV6OAC7C7WzEL1IJGIVYN05FClXqEj8YdesPc5jLptaP/Ox2NWDK53ex2Ry8wFa
LdJsS1T+GzoPImeoltHf3ssPmjth6dhPof2OTFu73t7VtykrA/Ndih5ZNCi0A4vbK0cdwjM5/lVx
IzsO5pBJuV+3gGbWGwUcUNZrh4whEL490VUuzRmwWWSiN0Bn1lAYVlKlc9/T7WTAyesZ6V/z9tTB
/ijKx7X+MePKhSlArFCrFfjWsy+VBfdlkhHTkHKnlLqNGW+sw5Drrqs6fkifoSQXPBYRT/zr0BC0
HMJo6tzg9KQQw5W5yoiASp/RDW0QtN+PCfyz7dxvPOQ9sY6rICj1zcku+Nxqejj6/aAVXSMZb6jK
MHZSaEmv04+FyvPalfvCEjL7DprjSnZvCJpi2bWoNEDYJoi0+ABhlx2RACJFcJw5qXWx5HQYkcvt
yIJnJqFOY9vovFjA4VHocC1iUr9wyhUqeoREjMpHXobjs3pqXA80IqCYncB6lHEl77AFWH1Etw8J
hp4RaeqVMiArn/GYFyJboRgNNJxOpCmys34kQRmA99yWY2R9j0fEUqdMcekIBT6PG873V8c+DaOw
rnJhEhve7gYNNA0FehtuYI7Ao0hVg1GkttSpTGk3WjCEm4A1sO/6YkgPJzX1+CM8FUY6Fdl2HusC
Q18ipxBBArbp8aaFnnt6IXFeMvRQFat0uxCLkpz3337qzPqnCVfLQmAxrhiRRq8yNbC/BXHt1xfe
mypwVsGeJtAIDj5USilpvUUHm8gnaejVno/LBQhpT8dtYu7EuYwabiK1wBGoXkX5iX3RSR031I99
7MjsGb8y86SNUQQ1gpbeWFKBB3zX4LChfSWXuhG4gH+sbY5dcgEZ7Zp4yAkyUgGcHITVDelJ3JQM
KlbN6R+vjUbHejRaUfaNREjGlnGGs4+mVyQOCmqgFvRiW4zXAKe7MdEPKqhVsjCldUNxOwz+O8rv
hDcsy2aTn/KN1r5H04JFPP78pDrOpJ2dJO7kiWnasrnMn/oJoTMUEd48VHG4T8ItZVEvZHiRL9Pn
4ed3Qs2BrNH9yqT09ALCzNXDeOQ2nZr96K5Vep5uozALcRd7ZcjSASi1zCCrcaF4j0734Ob3Iii2
zuLXgm6GOX8avVQWZqIIPfJmvARZiw6MbruF7UTXBgU7V5OQdCEqnpuzlXv3/JJLSlmpawlePpiD
2NCciCnDWq9TH/wBPmwFPPc+6cyKPCnKL3Jk7mltO0Eez6AtJ3qJZotg+D3rkKU4/3+txtXYNSIy
2d9dUKjgtt9yKKXj/eJR+BQaHGcNSfuHAN8bLIfmAcLWPdlpY4u81W6q1p2tsDwY4v19x8IZtuYL
5k/5X2M4tBUGes8MFWKmK+8OeyhIjA3qEO7iqdH0XLHJpmeqid3Rqr+kU3WcVoASM5H5Priwm0hc
RiLni1B1pJBoBmzWakPPIqjEWtjl2fcTGma5d49Sm31X9imVE6viapMxqKWUqnNC8Upj/v83j3kD
/H5pQ1ODKz+tvBxLXnA/sEcRzjyKd/zFMiUJlZhNcG2mSK+r0s60gMPI2utWuLvglRgdKhgAKS9g
9Tm3RVHExbupLXRLRvAaUcSi3t0kGmfP8+LhXLYpn9r0LJelgVAR9aMoPabZElDCBaHVCN7m3Wxh
qEOJwaV30xCmSqgrY0UZOOQDNcNZs0k3iS9v/uBTyiBAXp5JgYyPsRHOYRQ61w2ffkyoM+2H+MLP
qOS4V4hkpVWlanlJeMMZ9sNXMBguKnk7G+7nQx17Q39QN7rm9amVLHSBMYiNwI4QXf5N1SAdnaqf
gyqmIb4jMbvAyCoLukYpNHjW0YlJaDW4teGVZSaqTU7RRjnbej/AIhoUHuRMu3G5sU/vMcx1ooKH
l4vKOEIpv40ja3BuYVyUyPcQ4G5WNbjr7YOL3Kw1dxx/zUSQWhb9hKnmPKOPsdeMtqHFKdmHbn8U
5oFg0tQrq80IKDKf5ci52AL4uEZC6SPu+mGNTeqk3t9FZsYcNuYgvlxZWEeqXf89nG0KRQh1TD1e
Z3ZaivpRVS6JxjzSZMYvSMZiw4J2ZzXf1mufHhgfBISRFYby7DNug6U4WdzN5M08DPfU8TZgG9Uo
uRBUXtZgDY7pM3UvRLDd10C7mWc5dXenkLjMIRcDeDOiske+AHB+DZ52NyjZYzcHFFe5LLrYbvjd
vuaqpcJyV/U0+bVKstxj/v9RcnwOzodc9+9uFcZg8RlfxffEMs3bb6WgXydJI9yGeh+Q75VUah3I
7r4hEKxQDk6e9+h29mWgv5EI145jQwJbOYr7qVoXXAYiIsuplycbINcLsfEdWhst76SXCU5GZk6X
w70YIpC5+JGmqpng5LvN+29Sh/D1lS0aDpxt5yXrpgPJYhWS6/YwXiTjvVTyk/TNaaXSsLUnCxlv
BoSV4cCXV1LYtVgV0qi/9PWiL76g/AZGt0YRzN111KSHBb4sQPY6gaH/tZTPo/H0O4lZcuRut3+2
RR4OZdn8C1IyKqTvzAwR6Gan3SyokWlOFfLlP94dQfa/kXy5eXHN5CvbiVrF+/eLiMMtV+B6QNju
BjRexLeyk51m3qr7lQGstoi4rGBOAcroj9IZFbXH+kHgdlQ4huuvAjfjpp+V2/Br95mAEa53LPDG
uwWqsSlFgIF3P/8Sht9o51E1Ap3uchhaBtFmXiFtOi9hAsBruF5PaezUi0YlsBJjWjCaSOtdHqsU
ouuxYGUoZEuefJ7G754YGMH8aVNE7+aNLJcXJ4etUZ6DaI3a8797zlf8iKQ9LK+m9FUDf2C/Nk7O
b5xxt4B8GZ6eYwUzHmuDY1N1zUGXDQq1/hAE4lpGs6TdBAQH88Za59tEiN7yQ5pxdEJoseAdWjpS
o9XE5Knsl6dZVcgfOrq3n9gqaWhtsRDpYwQamqlI9XJRNuJPBOQnji1Y+LRIkF/kDSOT7JgzD71q
6QkCJo++T7Z9bbkgVbFESoChQjBuLp8+Nuxwl5VjhpHlYSgJivj78em6xKz3Tfkh8CLjDAqSe7H9
Z6kwv52qXA76fc3BokPF95np74MiBarT5felIhJFT+RtrRAUhtXkOb/Zjztm4QZFWsI9qZuKzkfa
CtRUwLuGos808NKAbC32ti+KFdI0Q3b8r48YdvEwp4KPelHdgK7eucH/AAWf1go94xSxF+8hMKvz
bQC42EaPLRdddh4dh3LQb/EnMzGxiFKVU+ps/XaZmXkb/cIydgxMlilkIxTvY3UM49JIoPE8w/jQ
6gT6PCoDC9CaXvRTfdSWONi9e/d8YBVZGYUdSFvznvCo0bFUsck09ya6S1Ng2BBK8uTMxkfIhI2c
Uvcy4MG35DRkGCneDwzwqW/jMVv3skId1o5OkcainYN1Z3oM5nDN1h0opeKHVSqVxlHH7sYhRj61
9W3601e6dOW/dnHPKaAPVd3pE1KhRpCx05rds9vKo7YQ5DeBRe85gVhJAkPCvhxY9nmW9W6iUVE/
LIItsEhNVHurQD7vDRkgI/LFm2THVSbk6PwIdAWRd/mZ/MRvulh1BN0S4TDpANQdfFm8JLhcza9Z
MdpypoZQygKC0lzBphrhuviYkjJ3bC5/xaI6254ejZnjiLssNArhLLRspKfx1grGgnrCiv4X4lhb
6XQBQJ7FFOvjwyQ6G8PvTziO6oQYZhIs6O90XZN1UiUruQ//TsrPEb6iavTT31I8SUcW+U2KkNW2
sTRjv9K+ZAxtRHE977ZQME8gS5yZCB1CFptdyF8o6ivcOchtQLUYw+TeKwRY1OuYT8TriUyjrnCF
slt/vcssep7CUVhm7xHabWrMYyxKZS1/F1RQqUy2S0jyHruYOcBfhk5uxRGhbe1KAwOTXvmQmmrD
d1DvTY7VfL2zkd36R2iNjQb+uWVmGO5wdZo1BALluPDYmLzZ+ZwVBqCe/nH0sXEkcMznNFPXUc/T
OERjzABPRg91qMLcRW32+isA6d7CNFP9WtduCeHp0M8idDICfAQN5brMb73Yt5DzSICHZtQpJ1PK
JCwzBPlqcch52OkFFPF+SuZr++zNQNxG5zrWz37WZjcgVeKM8n9kFEBQeMpDYjVxjQHDE/fIJGb/
uDPn4iopqqmzEzPFZZ7rltLvV2VM9rON2Nj90LpmzYt+geiYz885xA0ricFo7gKeyqRF2RTG9DpJ
UARukoO5fxlzB+KIK4D4+43tHbQMt8Vt0rorTX39+3BSS7OIRv1w/cE/oUEuO5cKX34assQNBLDo
SJ76e6sPZSW/ECp1Rw+eC+HxyaLNVjouYImNjShgUBrP/DF27Yzk4U2oYxmbuWySy2wYd3x/MwKF
6qgTNuR0KeHT0wwv0+YzqKu/k6sew6gVxacIVcCqCeStJj9n/jpdIWR2u3JKRhKcNqTFXlPbzI3z
LRAsgku+u19+Gm7XC966ozg3Oo3FHJyA12eHtgVdaL4Zni5Y39LJCbavjvJIxuYKa+GdS0aCIKTu
iHlCxOTW9/wgpbFQg0oulqj8Ju7DdjpgZFn530Q0y94av5rNpuSkUqAN7oGd3lric5I+2EhNaFjx
GcEI135FE3n5kZvyDS3vzHVlNiztC4kLS0Z1TNPb+ehYF0v0iWt5h3Rp+Z0elfnx3fBKjGZXpIN9
r+dIibZGi8Dhvcj1WxcKI46ZvVTITVhpW3rkt+fiy/898rrsz9oGbw/fBv4r5E6wBs2y7H+qiucp
xz5BvNTC2k/4yvjIk/j1wFYU4WGsVekvIqtW7+SEB4p7KNxhgnVL7BZNeeFnFuoRKmWB+4eyyVrV
cwbXbsZWlfv9Ci6z6EuVnt1JA9823TU06BGdZ2/R/tRAumZX6XfOe6aQLkdr/Vy+RwuEyn+A/XLX
N8ph8IiC2qfi99sgrjinIt9uQvDkH5Q0dXUuOdbvNmKeqGeVI5/OizMKpwAKFqq00fQ8mO/p1bLc
0HTATn80gAkmebKrMJImX0b6x4IUvTY+6RkDq0v11SjYvriMWBMSqwymJl1W4SwUPiVqCZUMWu+M
V4rDMu0kSTR2QREdaw/ZnaPL/qHq5o5GywEy74g+Th8d3wcdctka9v1dsJx2zzYz+m2jMLktMwFn
u2pvGNUjPRgg8l1s4ihIyQQ4a4bLejCm/3SXzhK+083tWbAE7bW85Gn6hp/GpKGVx95kf3T/AfsF
1JGQqe7XFgx9UkRG3jKZHe8uiLY4hmxHi1H7ukBBDEfMC5N8se16/Q95kxiOEd/m5iEt918VnWxR
vZlgPi+nbtdSpUKbZWE0c6tA3Ktivl85QZjVpm4TvpkrZdzRlTFfDelT/NkFA8ZNDkdifyPflniT
gVjU9iSNfIFLB62wcmjgdn2NsfjxtIpnkFovF62Xx7CKJur5j7JdHaYcFbNJPH7NS/2mrocv5Mrw
AAkOru2LQGhTkkl9AlQB/8XS147P0qXB4Hu/lKfdRa+p7Y0rTlJvGpTYhGoLmaPRtTSINb6nAEiA
E3fJq8/qWbCTguARtuitku1ciVUzYIaDPLnXfAh/N32e4wIPq5G+0D2KN8aIO2m1RO3ebx9PY9Gv
y6zgYqE42IkoG/fGqiIwkID0nAVMddPAeKBC5KXD8ft2Qli3H7Z30blY+H+ZcnzptCqlYYsjPF2O
IF6tSR6KLcz06KupcwV4m5RAcjSwG1iUgB0S+5PJA8Ybs2ohqk4odsyGosfEQKb1W0K60SFsHWZ8
s5zBGVzElAWLHEuNbCkAxBftZ4EdFsQWCvAe77mGv4X5zOZYs8FCzw0GR0EUvPQPBrRewMX5YZx/
FII40MukU0ZFpG791Gy1tyAAgYwQRdsXxT705zhSM0+ojizXVvY/mluuWieMnGTtJ7zkUcQS/AE+
DpWyHw7iZgq1bA8JOAFlYo2t4CnVUcF1JCgHSb2THfLxe/zze1TrUTpuyCWyO5mO7rlSzX3LOqOh
9vmLb+sduii+na4HJxoLRD9rNoJCsMYZqsEPBbr+i5cbxBoQPQiTU1E+ViCDN16rglHChVjHkj3t
LtqHaIzNHhRFoOSjkhwTJtgu8Sq2NaivNEm5U87KBlfq5XwpL4Odt8ddPoN3kolmBL2KwhSUuipi
/fjTHwCzM+aqckm5tam9+ADtcYmc7xNAHUsze6kSayXaD2Aw1G52QVZ2PDksCxIr/FgA046EaqEg
2Rj0VJqdKuVBWYPMFpT8B/HzufnXMwMq8j05wkyPFME2vaLWSBMzJilApW9/cIQKwZwhUyQCwDeW
AyFTQefm5G5OM8IFTwVhdE2KWjGwawjaZA69TRpvuBS4UFeHA5Gx0y1Y75J8t+yGVE4c5wvNKsUK
Zz5HnO2VdhdZpmhfq7VufgaDfdxo3KSHxke0aaGpN9PpDwM6knHEsP8Q0jLsWkyEXnP6t80OVEBR
Il0Yb1AZ8CPeekq8Ct+b/htCOaup9RqgZ8KAT6qUvrr6dHEF+BPeGiMQ6KpBdu33BdZpGvqB1qEq
IwszPQnpuV+V+WvB6MzQLszmQ4e7VbajGiuW1dMEjdBJDjT4b6pfck4JCWcC2pMQNjZmxJcN4vjx
w89szMBGtnFPm3nJzI4jlFLlD4jIdjuvpDUkZcBGn3YQNp3fLa9BWz6nszXMuzqR55DBO9a34SE3
Azy7B6pEQH6faKh0gh+mREK/wySIe09tIy+/bcKaBI1k+8t/E1t9yFyBNnnGhpIrMr03lISH33HT
eKqXFpKUcB25CVxo+YVzn5PDyMYXtATpTep2wzjcOSgXOfpz6EDaAHDeHWbtkHpbmQbHpMw32qyt
uy855oUSyzuM+G9r6K6XLXbnUDgkajWGGd7i/lYCYmv9lS53QPNHjStq7goJTNmfi+Aha+Au7IJw
eJ+EyVKtyNm60N8gHz+tk6WbrMZB13rxHv/lo1Q+hGVbLH0wlME43DufZsqMvpE7r1E/fEtkQWbn
UuxvP3n2tlpQ5iky4tvHfZbvi4cZvPqSHivBKj4Dw39ffCmB2iVNqjabl7dKPljAPvyZeaypERLm
+VxAUzqG4GSynvUKSiILIc429kZLRfTwc5/jkP26HcjYu3XJLdKOqUt9aGik8Jd+xS1DOOnig4vX
NfFm9eXWWggn4Cr10d8EDge9EylUhj/P+2YIqsq6win+f6FDw4MgM0F+Q0ZeNlDp5GdKjf5El1GL
TLiJj4vsKH2GLlbpfSLvGCbqXUVCA74bjwzbLgZJHNqJ7GQbkiOth1dmhWnBgMWutl/vjFi8+d9Z
z548wq1Je6nSpAQAQpoN+fJXy1t5z7cXGGU2EaHMz2+lPgjm87s1QGuXRaY2RKVpH08wiecb9gdK
Kq7FSkU/1dFjImBkMC/aLCerqkcNRgpsB9pAXU5IYXIKBalbGEgy1mozPdlSrzyO8FKf22TDdU/k
7+N4afwAy0EERihWvRHox0wdjjCk1+rXo7fG5EyjkySSmYPJaP5GZ31cKO3CTDne6sOJ7HtRZQv2
3AX3wLNffs8Cp/uK6dsr1wbgInsuFA608SYF+cC5PmU3iGQS3Aowlmb+gjxlq5BLhyed6DnbpLAz
L9weUWOLwwZO0zeGQAKoURJIDGXp7twdhaSDEy65gEeWY/sJHYR6ARs/Y5bq8mbLY3PKUgZFMS6t
3/haOhM9FFsj5rwsqAWV9eMyZNsSLv+MT/BfB2mY/JzNSTG4MLmggQxmrFgeOf30Hbr6VoTXbKoD
YjHFwPH+tNk7abk2IB4BF2jY4STbjfDBdu4od06V5P0kAaJ60I4z9Dac5Z5r19chJn9tzGN9PvFf
/KUzuUnvihApR19VyRd5JEfEt1bzWqHCDo6LdMJdbuvpMJmogP7cXvrJa0JZLYj9vkMDrKd2Mf61
RhTnDAOk2GWo3FUkZn4hkT1WDiQDI8hDP4CIJFfouDXsT4tRyf1LUAYCF4XFy+LGyKkDfLNKRYuj
/HDg31lBXytMNHdqTIqeL1P8ay66XTaglDv/SHnrp55ynZUssfcW8/67NBYtGc6MVGdOm+g0XHJO
RxAEljn8TbLsZVsbj5C0VL0WEoAzPYGVB0oCrL7b2HzCnnRDBEAkX0jJY6FCsJKTTPYr4Nv4CdiO
+HJMhSPLxPa4aqlGrJSH6eAnmn9qrpv3BKkzmwiVp6Yfo+8B/AfUqHKRROIomZnxla4Z7v0X6mUO
1ib7MAa26XfamSfiBWW56NrC3zo4SWh7VUuI0QtJgzdgjl/0n6jmZdNA0L6UCey1NV3WI2bNNpuJ
VNxgut/HhR/opUsgRWZOCcZQGIKGKmdGX8pQwZVat9A+4mcbVn2BRAfLCMDGt5B9dWQIABpc8dP/
ChxATkilfSsgcxQ5tLGA94NMsX96eZ8kbhXNWqsg6zAyBrL1taEF0YgK8U5CKv4ODrGQbnQp7OKc
dd5IjLTvI6uRGM3s0gLqmqGax+Ar+IVUd6t8RXxBMGaMPwep2RmbCWCGUsEOqQCDFNOX3tRYp0Wi
IbW/lGKeHb+o3/J/Bby0f0UfsMxBVPWU7bw0qT1f6fQjWFgwqGAiaL9eRIwamjGk5twE5o9TUS5z
Zx59EdbmuFvo6RhQhPHfpBiRstAXh6y6LLH4tbz9xvO6w0EnTmreZYkdEf0IltHlKw5fKrz79O5+
AGvfTLZYGs3mAMWp9iVaVY3eIMaiqriXhrevTVUr0NPh8BCP/MdOQN0v/ilmmyEmg9T0o5F9yYdc
yh+2KWX/PzwPekSs78/N4BSKHmnPei0eSnGwGYi6ZNAB6v0Ku8CJKSNO9nh/U5b98JSoLW02edqZ
8TfRqDFsvgYgnuT+ZXAZk1ISxtgnGcqhgFnPSPXt/euZ8DB8n6OI0wZ1sfLF4u5sMWlaWohwNlKA
L5Zt1dPQm3HNGjKsm8dXz0Lf7A8LeFaM4xifJaT2YQ2F0l6kD7qXI8vMPy7Yf6W3cWRQ18kg3BnO
PAMw8pG+TFoDuOnfMQYU7+Pis9Azg5+DXbFgHZtkh6bm5ATxv/3jEZpg1pBjw4v4PuPS/xxaJz4I
r/kT1vUsjUiqTD92Wvz3blf4bVxpFAN0VZGWHNI6a7OAAfvVJy0kUlRoTnHwhRfHZ4whGeZkaS08
QpOBUvzRZTB/m0p+c8mm0nqtoYry2fADpgUUQlo1uR/kG0DfwWo5cwBhcuXJVV7wPY+zJl3q9Uo4
d4Bid2KQPjIr0VqKl9Ps8Ivmh5ACaUImGVFW0W+K9iFoRlCU6StBLrL+1QlfIb+Bvav1rqTxRBVe
bolXy85l1HslIw2/lXk7kS4mSOJ16oQvLsTc3YkiTrUMQeinWYZr4W1V3asd/fQ8SvRF4b/zmOzX
UGf8upAvnHL6gCSe3RZPiOyPpLbwr8r+Cc+cU7BSzRxA1EB9kEbOxtyuYBisCNY3OYSkvNrqyJ0n
8pEVfjqnehM8aWdOZHaIxZqZsdXA5tObTDVu3d3OJUSQOt3YTJhx7ANLtGdmijJOznz3Jcpf5nWS
Hlwf54roAggfBeQ7qzbStE5rEXhjahaYl0RwLCuyC8UxOG5QhtNR2NzEK9rxP36SDNJCNos9awwP
IZ4aWrXksiYCQFdmeRsopaj06eX9g5RfkiySsgk4UmD7U6IRU9pgz3GdpwXxIHOnNTYS6QpJaYLV
xZ3bDFpOZ/83aAsZtwn0I6NxmG5TrvA3puGDcFt2UGKDufHUSzqqld8qde85CWphUtkPSffE11j3
AldDfoYoC0oJDbkSImsDye/5jxWZdO3NeKkWxS8noHhzY+6ezgiH8sieuAmrE9d+O/WxJ6meZF7v
3UUmTDVncaFdryOQ7oqtrgjolSWmgDyDotmXEUmBqOkb5g7nxpSXUEM6fa+KNpBIUm726SVF2zh6
/XZ1dhqiwr12Pg1lELvcihHYJrwCG5/WBn5XcxQxgVsKz8l3DZqBEhYnryJ2nPAVXowg9mfjMG6N
kVKjsvZTXLIOIOSaqbPvX98rpqoY2Nsaf7fFYPuBfE7KK6UE3UQYF1umQ1RBYo1pnjhVLf4acPC2
+BGLOMbpwfefbfyw6azJdZfFTWP/B87fg3NhoOTC7QuG2tIR7f9/EoD9HetWCCKe1bONvE+RXhM0
q6YMDJSOiizkDVfc9MZOmw7DN1sPb3der4B7XN4lny2IAfPKmUi5aL/9xl15rZ5dBorPWDH5jMcO
DLa9n/yrtwt39Zp1d25s9kr+dMJ48yPCxkvVImuc3Rob/ct71Vky1FtuVipQ/f+/dafCkj7zNq4o
xgPtA4qGbG9QH7TFSqYK0Mx0zNeWwXE8tXDy4KO1vGy9HAmiTc+Mle8gD+deiWNNgwFJLc1B11iF
vTw2HYyP1jOD8HlXEiGhMgpkPdtKrBsrsaIBrVa92o7MEZBliNYW2IC3FFYvbzdMLRDyE5ZG/ADP
yh/Mz9Qq+06BTVR7o6hEo0pf1/Oq93yjRauE5L2qK+udzw+8c5an4XRNn8vN2Rxuv10lCMYRGd5E
LADzSFcYVNE8vuwHeDypopNv4w0aAwfm/d8sV1RZ/uzUa5L1OMOFiUomFxZmfIXz2e7me1KByKwU
nke/2Ut7JAkv1xWQaMLSSDgKZZJwHjMambgzSc2XbgSI2xa9wyK4Sg0dfBQhYRjMaK8M3e6RWhDn
m18CorJVEK92Jh9v1iI5FM9nmJDcFBnr4msQ5mRf3tcmMgrvSU34VJZvmBvSmYMG3Fepqrpb25Jz
Fm1j01rR69LjdQ/gt5S+bZZGkkwsRAsomhM+vWbFJE+7I0ekotfc3vCz9htVQ7r+/XRl+8P1eSS0
MtWCLSDiuZSK0aSjP6f2YGXahk9m05bqf5n+w2pcAPJIF4UTDPYj7F+4is04Bsq8ssuHnpdEROWw
4bGPpIFeBnO2douGvD0Nnp/HoW+2PGcGnqcY4ZADgZnrJpwerhFA3vNdePiaRHXawPqCtT+4ltjJ
zBGp5p1l/nyzT4KeCGUMOm1sN954eubUTJrt2jdx5Fc+MRothK2ZVsBt9GtewkiP00RaGtRvyvqL
cWD7piJzFqw58n3PtRU8zfeAhFFD/j77sjDwdkuak4aJ+N9ZPiv/PBGpa6YSpvIudinMkwjQ3kAQ
05gw9Ihu/3M7TjpA8q9zXLuSxLfLcpTXDcHpQrXwSkwZ5J5FE7yiQ/mcWmkOzHRtOJnNRptvmF3K
fpKwk8+JlIPI/8Mjp5vRMoZxWMRjug8eb/eALFmTsUQ0W1ZPUxQXpEpWreRZ/w3zr49Q18HIQez6
LWBwhTACnUCPDuezaPsPOt7fsYvEllZW6yL5VU+X/eQjAwqlbVZGreCcSzPjSevIOdsJNmy6Xpyb
GUGLTXzgHxfMVqe9Yto+i9cXHlrD0lcMq0wDyiqbZr6HlILw7q3HPjPg4iMJbLIphrEagZRNrZ/D
XpqqxN9rz9zo+uT2NLMbQOZ78AkKsGJpZWUK3J6axs9KFYxY/ef9iMp41ZIvETANcoSen8Hp7KVy
2WNuN2aEfAh+z5/d+yMDeKMufkUAtt8lFs7kM4eGtijCytd9H9SjJXhnlhG+NbwTwVRxfL0f7PUS
2RUkFDXFt3q5Y+w7ewzWTPFvURlr7lkcScP07WCZISy5Thw=
`protect end_protected

