

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AEDf93kkZknTAYDLPy4q67UmP9O18ta3jK/RtCkxR3ZqpY2KlRt7rza1H96MUf+qsK6643W9A0n0
TP4few4v7A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
erRjv8zI0elbdGyufePGLqKRctW7EMRy4ag4V3lsqysjcz2IbkoY32VNXZB9TkYq6LxuID3xgPR/
/dbN8HKNlVJr4fTV1LqzlQYnx177n3iaEwIdtrjwP76G8DtyrbDzV/JISwzd650MMmyKJtHnC2yw
alWuAIIBdbSW+HbA0I4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gdHY5LRWuJLwhBPcRYPMx1NPD/GuGCtHF8ywmbYLyoAM0rjTxb8zBoSHfJbS/2vKpgG8RCdZOknj
FMJ+fOkJbpOMFaFsosZ9XfIryZEhroI0pt0zugw4Ha2XsmQGqxGDd3IyGRBNvDMKRw2cnjSZz2Oy
H3SrajtWuLhpP/vuSzlhtnqryvgbp0USaL81fja6LLlPm2jXTcuqgEPsJwwUUhxjUSQyRtABTEvs
3Vjc63pIVZUYkpkoaKpA4243dOoRhazlhTF1c2Dp3uyCrdGZU4fWhJHW7m3Cq9Aw1murzYGrPLS4
eQrf4MTXbiMtIPpNK49OUBbEpUuLfnDwfATFaA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fCQs5S/zt//IgxsFc+FuMl79LHVh3Px9B+S0yADLC6MfIDCRddIdSKbTMZ5DlFrngWDJwpd1JzqP
cRXcul8iGoVMrVmrEStKWXi/mhtK5UkWTAd7hoyj5zcI+N7wWWxU1eBAeKZQ7uML2SLN8mYzQYLY
98ufqGLyMQeFAWp64iY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rLzkYB2xv7C/3jKaA9rJ0Hz1NLTW5YORm+QksBhLo7WkyUXUd0Olk6yTtcSIC82lRfBo8f3njqY3
dhmWfikGbTNV7gixnGfPYVUvZg+xsJ7adfqwnApC/cK5eBJGeWXZ3Z5gEbLOhuRw/04o37fRIoCo
Rt8ZH/C+LE5As0rIpYw6uzjL55RYR91wP1R/rUwMQTNJ8XwXPkAbkuyw7FWG3uW7vEvZ/CGu+T1f
VDCUznG/Mry2818W/OOR+t5yQ5fYiXNh34gzkO30FRWgtIR7ZfOn/fgLqv2Iaq5XPzTdULGOHjv5
Pl+0fdEaYyo+sJ1yt8Il53T+ZdgLTjEgv9cjPg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 30320)
`protect data_block
foFSF2cUxo0FD5CO6hLhcJIULXLcp+PJI9tGA0kVaQfxF4ekLtRzHdPP3vVezYfybQuw7lff1X0A
LguqI8L6ySRGqHGGSC5mCTNFR8hTZst/q74LJYJZ51PjWkL/t2vBtmw9KlqTdri5/iRSbCRNFM6A
sx8m+sBXhGH4x2o+XzcFFS3O/jhDSSd6XrZxkd7tF3DVIpeQ800lIV2MjSz1uNGrNBDEK3FcySyg
UQeUThQrxQ76PV/hEEOBP0JmFB1ibCS5jW6OyIVH48pbJpUwSCzboLNcnZazehdifGVlLG6pUbGy
CfLA1dzjbcfhJz/xCeTOcqx1OgBMq8lYdTiCZrXHjUKV3TMnyca33phGO9nBT9UfHx8pyb0fS4GR
qyBcD/CiHm6hvrKOdszMjlki6Mh+k2V7AEqD6HeECVHandbs/4U7e2UGCw6/EeVn23XPZuSMr30S
0JPFWAMSEEtlCyeIyYP/MdjnhW7sDhsZ2eox+t6A7Zhad+uiREs1DaukuEvLCHuREJZ0JXLSZvfb
19H6vjwI5HK3YifLaODOMx3MDfE8aphfrEqt16flI99+dnJrfIInBjmtfA6xRJZKBVo20R6bTWc8
teWf5JSdFuhJrb/okoyesj0oYSngndbvTTNkCZ8pcr0AMgt6BOSd7owIDv/8zfmgrIUjx5GW4/Rg
3DWDCxkS6LU6r8Bqdy3vDO3AjjLPIy8NOxHXvSn95dsXEi/1S2QhdcE0eSBDTirsrs1HWcIxZ1ve
qznauRa6auGigA/Dcmf9Uw3PIYbIESoE0SjooKr4cfzaGirXTEr9t2s/Yu4P2HjJWZdjL/L8acFG
a74s9U1oMgdRWWtNjHnHx5yt1vhkuM6qGCWzTxemCWtSfjsRQz3pk2AKneYXDa76JunlnS+le2DS
Sjd++k4P1Y/nd6P0LMA+L46Ot7iMCISef+8BNegQworPjZO5HOYHTUNEeC50B74A9o1YCrP3vhM+
x7TbWocf0YfmcwX56H/curm8ipMltkrvoc4c8Qbt+PcJX/MDCIxR96eswrOXZu4He027q9XXuMll
cGOKuup0ae1djcGhcKrm0ZyYPFoEkKt6HuHlghsXTV89z44JO1rI6AClM18w+t2ixWCH7U9/2vys
/U5zImCunXHdehKDwm1D7kjCDZR0M8im+l4s9rCbSoWwwm3UMWkeBag4OrQTuGgJcLTYdPnPEe7U
Tq9pIlZ7gLrSwg55LPbfFy6PI3OYnGwNMyDPYAbM9dQsHfVAu9XRsZUxed4C3dqMzUWpdjbIjhE2
fLEB9V8e+YBUXOqPdBecC97+pQpDWQ8ba1hDfO2iQzWp3zM/a2UenOty2Fr8e8HqRNe7rIbP/7mM
TLgaDHflkRJnTddzy8QnAgfGjxJ1a1oTH7bvTTXxp3zWYohleClXJ2/qBlglrNGXzcJlJyyMw/ON
tCitG4wj98CO3RAKq0Zo3QO/h2ItNk7kV3ByxKhRnUqLPM6u7rvAgXiNz8Q9Mdp1QjSFW7Pl/sXS
Cy0LHKDQRl+reOELFDIZq48dJKJ7mQrTFDeYw5tfUE0xMoz8OdN+oQ/03OxgRyLYwhnEVDlHc+ei
SW3Ns5S9pFZNT1KsaJwQnuTu9UlZy+UG5ApPtrwUEJXXh3+chf9HYrUvAOHEzwBrzMBvGdIbjNQh
HXPm/UUcFd44ryprqcKynDz5fSL2q016GV+ml2EgEkxLIptGnKqzKz1BbdTPqt2Wuq9Gk9L6UCPZ
K23zhV8kFnGppRxdp7nUSacunJnaKbgQHpYxFgj9d520gyijxHo62oMLYlWMsnbAY6BOg7aWKf+s
DgBZm8oDl43vGZStS97qb+/toy8SakyZslLcnOuMAsKEQ38fFKzFeVk/F9gl4RQm53X9Ysz8dCna
010PdiZOko6rG6hT70kjxxuF8THznE+x0Cv7M8eSMxOt0X2OEiTwWL8xvPnWicF9LTzwoH8BNp6y
Tz10k2SCnQBpPTxK0rDguoYSBGOHlMC9HuO+aN64ZH4cOiH7PXCyV4e01HtwiaYAkOiBKPCoIKoc
ilI8OMIkEjh9W5kjOncCuBVQanq0uVLDvt0xGCi85TTH4ULK7W8lcT7RotWPNcxTEct2p6dA16Sp
Aqwvf/Rtg2Yyv4M0+Bo8zm53uR37B7ipwNO8EMPn3U0FmSId1twXuYaYZUE7Sx96O5DuA4Ow5kHu
hsCJhoLa5zfIS7ZeTML8wDH1Ll0Rmh80T+DNGsja53mqprEx9VkmBtkuzdLmuCWbf0zju/RWS5aT
WKyIkmJ9E4gzGcx7UVOFc88y+9KL8noxMyxSWvUfwBhxHxrPHGOs36+s9VqfpqBZjCexKa/O9kVH
NNl3COYEZHGUn6BzZrQOemoxsMV92ElEfhR/5Y4Au92hPzd46YuEL8zZETcPsYBDzgt+o5CHKXCx
kMVLtqLJT9OmfCcyYk4Qo3R3bheyeannnQ0hH6R0Ju1TMGlTgrtXocA4y7XN+NyXjVh5ris5tEO6
VPPFq8uv+fOqo+P0t1dMDGgUZk+A5QVHUvm6E+dsc6znrdsTYf3XsaDyav7ilm7F946O40QDf374
6TvfpH7bSeDZ4tkirsgiG0AUXM/jlwzWsS4ZDVay5qmXj8iG2LW9Hnv5hUKphD7WTDpwFX7U4wye
l6QcOQaFUZb9uP88t0tFgW7JUdxUSC7+ezaHGzLrPqX1SOipPFde7JCz5SjfZxdW8m4xh5MoxabA
niESnUuy5Twz4ONitmJ2qaQvJ3ZNI9fKUqSRllPZ4eUsVNTXhg5GYUhKQZxk83MY6PUH962RFzvI
fFrcsdYJfe947xbLn/o+1Q3CtF+qoUewWGIcCEzYqOnCa4jAf6gIXsUhp7TpF3wEERvaohLzwRoO
alC4UXPNMWnG95ranDlXcB5ww+qKNl3Uq5PlaecLBES6GaTi/YU6GMkf7H3U7H0Y2WW8dEnja9QV
0l/RwHqukCbhgc5GjCngUQnGkbSKfKcpCUZc6QCPny+q3w5KBYFgZBRt5enwwQ9P/m/FyAEnhb+T
gIIl4RZrqlGOZ1DGOiu+0ke+8iqYUHV/XnJ8rSU9xcWf54zQ2sb+5ialI5nhRv3VTe1XW6jVombO
LperR+mfosR2JX3iotcfgOIuqlE/p6hkEmE3rI0o49rqqRA9L4PwVdvMeKaUzMHBpMpm3E12iOVw
ncbViTh+y71ATxQ0U3SoxGXFxxUWCKCgqSDOMSKUJcIhqWcYJZZFAoS6xmk/2a7LJEc1yaehQcY3
lOtBGokYehgrR16PFc82lYTvvCuFELrW9+Uvg3J4aplWHUyA1sK+FV6b16P0wjgx3jZ5P3z8Grs9
3IKVvXRY94GaMwGbcy4vFxjqdglO+kauRe21TLxQKUG9wkzIaAIXgNJP/FdR00BOBbdSQlNZ+2Ha
hGKApf5rVVlTpzpfxAOrQpDxviV+OBfWsDL/tqFhlTNCqGAtd9rgt4KB0h6wcqImWn/BPCinRQSO
U0D/3SWmjCNpbzhKd8Y8rSP7m24NRviyr2vlagGcV46cv1GCzyRiMGSqlSQD/Ni+flE6y1xQL1BJ
kA9YqyNS+rLY511YyUKdYACx7HeM3ui0NlpevzxBfkwngt0DfuBlPffDNR6fzXgih/VURisu5yiB
q1iUW8YZwGV4RU51JLM4pH5518zY9NHP7svsVZBqVHeXIBTXXG0Q4HjSg1U9iPGyZ9YGHeiXUFJ+
aEKkWA79yeY42XSTET7oF315KThzk0bFuphW5v0FjIBuTk3MQJS/v/C6WdkTJIMry9qwKvtHHQhw
xwlvQwIOVvF8hll0Expe+e2n7oZ9AJg35VXcYtQxpbQTIypc7Tc7koEAp2qVvrUYhAVJ53v8Pw7I
bTugBkyDlK/aH9yu+kQVwBgtDBktjLbOybfvkEWmAHnkGY2HOGIO87yPYj/E3tBR1CD7C9HGQep1
wwjrySr8drzhgJRjx6q72Bt3b038/cbiziKYRoAu7EGAevu+l6SSsJIRIJaRrOFQrTxNSWAXbKej
yL7ZVZZywU47YiKGD7mER0kkjdAgwRz1UohVRM3d+xy/SDNGSrtvu6ZM4OQ5G25098ZB28hZrtqh
6+LJGhLKHeqslIDrkKoiNtAQTPDihI/vpT26QtDPMRnV2OlDfWRhCEI7BZ+0C9tZjH3fCQNAGBp9
/GVzS1p/zEFlEyqcmEZXC4tTadXCHZkTZPnE1MFcuub0rdFntiUM9zBf62zboqexVRkKl9CR0z9o
QeAGO9M2eQ52STpD74Fx4ZAm16NuuyrNQvS5FVpDpI2SoOpG4PdEEo7kYQ8jNd6MkOSZ4ur5urLK
4nUWBUpDov0kGrjYF6VoJdh5pbv496SDCDj6vxPVdAEn6OpBxqVLTW/2hDDff58uNd628X2rilHz
3/xuNEvBzsWG+xfjAcnjuVj0G8pkllAq8HrkM5kuuDfa7ny+4iFcoctrdLf+CuxoI7riQSctzDby
NN5ZVetmQP6vu3BCWwYYoWwAdZ68xmCqj4R/DIIcxA0XmRYnFOftlexjG/OwWJDDOgAZcTVHgX3J
Q3afZhBG1FOb0RSoIvxsF8zs5mavBzcwSwNmKE4yPs/S4x52Q7UmEo9BjY70TkOd/BXMxg5pHXoU
+O0oiL26KZ0j7r5Oz7Iu8dfJZC5Wsrgroqivf3LtO5FToYzrUmepHOmBcpEUbeleY4ZD9drhyUzY
z2J7C8PCDnXKlb2rYVdHGzOv0jO4CW/eX+uZREMOuRpZJYUQpyxioC45zB9WBN/jZKqSwdIzuidp
P+9AOoeOmqDBD3TsUcD/d9v3LkcIUx4u8E0SYqcIpOGrecn9r83ZcYTh0bONiO4KW7w4rl2+Mzgk
n4HN/LC9kXqPpnm+VxnXIE8Qgc1+DsDjL0z0BNBBxP1z0kQPVRQiKEy+SyJrjOMQyXPz8kclGD6U
bBMEXDjoEZAYoJagCOgbNKLn2Sa6Eo+wSt5p7UVrsTZETXZ02liRr5YpTFff804mkakRlGMwqeTp
zKHZmhlFnCWc7U5/imhrPveBMZe/aWk0UlhYgxYXohzadQSxk03cqP/vqWiYIYg9pvmLg4v2LIUm
1RRTTR4AZqgtzWNEEUOhXHO4FgSrn2Js+f4rYlSHT/4jgp6/HV+WZZHDC3qHEkp/WYanHqgogCCz
4IZTjM1O/87htQOpaAIsKE2JN5kzO0/jBu5WCPrRK18691UTZiL/4mIQBA62gF0EoDS+Bg+fLl1J
f42TDKokVBBaaSVVzPCmjpV4InQAq2SIanhD7wupzWP63wTjptPO+tMu+xhpu0VtMxSzijPq6iTB
a/PS8zJCWa7/r/46jNl9kmGnub61yx+75hMzBxeH32ML7vzvVR8CiZNjIR+FQfjNNKLLy7vVEB1A
/gQoPi2rNR6l7zRbFVNKFheAq9k3U1l0CWH/I7iByd8A4JDnw2MHDp+bpC1/rzcjV6RNaZOwfrX+
8iRS6WGT4M/Bf3qlzFXD0Bldcfzile5NDTKD1sxz8e50ugakbSapT24D9WkXbjVX+bqywFUJ4f8G
gaOb9uA3XecHUWdrVPAy2WrDqW7gzJm9h/emzxl5/aX9lNnc22HdWnc+0lyEokPgQjlXvNaDYbXC
AMDjOUjhlQZhJlvvuTMLpLdHHGCLvVBrWtOM4YMUEfLl1yiHjNtHiLgyTGgtXxFuYSF3g1uVRUd6
WDJfg9+SveN+xiH15h7rR5PMSd8cL+qz0OtiYMh9JDhTf8Vl7ltWmK9elDS3mrd4ymBVn4v02ep+
f/YWbXM9Gw7EGY4UzVvcuspTw6KWCaPLYoP7cKR5p4y+5Rpnm6F8gEUl2Enyg9JSx0Fjz7Sc3v+G
bX9kkvMsTbB7/hMIruk08FiscAyFO4DjKOw4OD3yDSkIFczRCNHsj7gJ03ZLji9v95SJI5NQKC6R
LhNP+ffKTrNm6u+Cb4usNZBxyplDhVXa0/NUOVFpfVLTiEzhUpPzJ52satVfJAjv31a+SCGbIT7V
gNN5M6Trn5rM7YwaBXMIUPHn6Kq3paAR3fwhnq+ia09SGDJx0BLv4tO+rHryKpQXVBa7v3dePNx7
fZaDOTjNGEbqj+ebsswGrtvlnpntkXpNrgO0ZKbKbcAKMg0KsG5bbcl5huye8ifYA7rwqO3f4LTv
iGV5rASCIhR5LZuDoY0DG+UqZ8G3Ypi/XM08rz8kqYXYIdzo3VmwrNI01etDROwMt/IPMF7bVePH
Po8huXRjjFXqsLA5zESt/Qf2gzLYDnv7FeZ0Nqb6F7iCktx4Gl2WW+qTXyDlLMlWxI/pUSt4Bk9Z
k62tiZdfWCaF2PIsLklmJP2/BkKkYyJSaN376r5YTmw6qiRThhFUNFYqEOamJAxR2E7bwexnEZ4P
iNv9z6d2tQ5adFLkMIMLZ0X3Sbi1jwoGgqbuLOdf7tduJ5xX3j0/z/2fULHBfM6FUjuRsD7w+h+J
2XPy5TDiIScxb1sddlmiwymU9o1+2umyAwWzKiSzgpwprYBM7N9asxIit4Xb8SgK0eQyDWcF4uH2
Q7GCnyXeNs0Be3SViWesg0vP5mFURGYTdxRtUK6veu2SnAcU5H2wspoB6ugi143yghkzXjAr35X4
LmFHUNynU2raKbp9ZxO6xmpRbTk6fxR5ra5c89Gh+ZrO/4M8Ao0QsRg508OZ4OevkshELoVghUdz
IStn+uDuTaRfGbBHOrVKDF34S+kuhhs5eqt+j3jzXGdgVaSfmctOJyic7ppU5lLCvGS16OsS7T7X
hvdE7QXehi2UuJNp/fNXL4s5qGqNMet2DvXCd8y29DU/J27uuNW6+oSofl3ap1Nd/bYNMVuXW5ww
dd2ijiIx/Ul1YBzsdI9l5pEkP5yfnycLi2DbVTZ5Uk8DPkaR3MC+5dOftfWzAU6NmrrC4RbgkbSH
K6nnRylB41/1qHmByRNjVcCb+gGsKfR8UoiSbUShISUC65T96S6B3AzqEyYckamr5Eqcr2mYd7ld
Zj32QZeQ75jwutENNlL7FEB9jDbntUct0BaQ+v1gQBSxxHo8BAEQ3bGL3d7e6TK6GwGx435nl6PD
yn2jexcyI6OaROkTPb1yJHjrUCRRZxkXwDKalqBJYyXCpBYdvt3j3L8mGizH6/Lbd9IVrWtW9WPR
So0iZuCbdIRZ/HpUeahzRaVBntdl1fH2/8MNtIbFYMuT4JrhN5cE/WxhPQvd0VluG8FSqsUaV1OH
iEl8p8nyw2dhuEDaFu2rn00mHzSfG6kFpQHk/2Y3aLHNyKA7JCGRVqyH1CrF+leuyr60LLovXUgL
5kejEi/T2eiPZ0bqyBh/y++r+uxkZ1ZsEaDM4Q1L/mPbRAOpSeV4V9zFPTULcU8wwGafvJpZcT5r
DKHsDfMLyNbYmr41daIKQAUgeEDFiAEDBT6Xke1RIzDo126uQP9EIAc9KWUNWZco74qOJ/5bzdqh
nR4DCvJvkGYrtLr2gM45DzRIiZgd+VP62eqa9kjSoiLu9irn8DC44x+nHmSc7DFZ80H2agsejyKc
CkDsMreGNXnleyb7waz/WDDCkg793ylsF7TF5/0dRWEUjCOPQ6MZrKc4QOaOlO/PJSUuAHpQnabI
ok/P9sR4N6nUtwwWoVv8fXLVGC2Bn7EvpR3LU6zhcAFAjYdJCb0Zb7yXg7xQj+pGumDR5lbHDvvf
rDM1MIVPE7T8ppgNeXnxNVK/t+7So5So2t87mq2p8YwSXL2itX2tIr8yyjtg0AFw87BOIUW1Ibi/
ihC+MyjHXap2rCqdhBD5wLFc6JtrFz/ya+8dOMjxM3EDhSSbb3aqwRolqKr2cfEcPauRFmVDVTMa
vrhj/vXPaY5DWGDFvUSw2HQyTDtJ6il22EskgBXRJcuXN5VRYP2sOcH3I24PWDMffXJYHLxo9ezy
V6BUi4bRAHd90E3VZsiH3V9hasDBxWbPRt8IoyHeNIuabvEzzMxkIv4ECv9nAkm5D2BAGYXnePG1
1KBegowsmE7cBJYxD0ApR8k9QJ3ZKyH5YabywmSB4A+0yPd0mU4ni86Z+tr+B0DjBFUJXfbL7RLE
/ff9pcboymM3EX/9Vif36WsOs6519JtmJxyusnDWpIgH5U/D7viCZnpOoBBOcUKG7nrZTSkezMMK
+feBJM8nMzD6JFWTzwMQYIx1+AOviwHd2VTauVFm52nOOvRDT4tgbq47fkHcNc7OjOpKBriRslcV
wEFu7No/EZ0ABpsuBzVC3j3F8tZIdveGyhFvehBx5DRWTHvp7nLLfs0oKTnELIA1GvlZDY29xkvH
VxOBwBEB/qSaCU5jzS1oHcYpKV+ttHl6dd/BWAHctIhM3vOdZQ+GWpTE8WyyNq4WT1Vll9sJp10A
rpdSaU6hlKiiy+MP6TGVX7e7DYiyevjjSzFlz+ax2pBfD03DA8sWzUH29Q5FaCLXV99jmxajuYOH
oeR7xR5DIJbX/gthFNwsFExqxu8EhjSyFeWc/GxlCbVcAWdUMDKJ0/IhSlDcbXE53Ir/Db3jdzUo
LnDCd2je/8tSWY0G6YaIdEqXqmTW+H2RxMr4twzuT1LgwP2NGDSdEKobRLO+8Ui/nfOYv+i1Dhlu
/fzN+lzOY/ajc0RT9o4FIsWCdmpnVJ3Ff4XU4Yuo2Cx1V5OFeTS4wlyY3/3WtTUp+77FqqR/nIja
5TJ6Pjrung5myM3gQFwmO/Cv89ZUGAzppbPBFhEADNCz+13ZVfL2PAhSzHYjowYOqPTrwIoahJIt
9wjW1xyIvur96/oLuEV2mZ41FyEDWCfr4ricjzAICsiWWh+XbxJl6i1VjE5Q7EYOA27UJuzQVX41
iDOlDy8xJw1FDPClmhMPklQ4Nk59EgzVILL3EFjZJdfrGvW1jZXT97H0BNcYNCcqTzKJ4NOpYb6b
XBjEZoTtdalPdV55iOnhojBQVbXmnOYoTByk9ntyEG/jEzpSnBNNA5+zM8vnBAtUnnhtH92BEmSo
cMFiovhUxOCNb/LaKQfoeVjdQ4ZE1Gwhs33YpPj2p4fV3r8miRzHVPi9G8tJft03Na0bngFy4Gkr
GD5FrzJiqQsV00E+S7QB3Xt+Rh68TNEdUOxaiAMxYOYaYfmFnYdNsxrjqNf/wSiAYLnEqQg5ksNX
f6yxV3a9CSXFwOU9r1zftE5y6yc1Pqg5sAaoCRwy6T67e/NxWaBzsgXSrTJld9IQ17smAYdm7QBa
gHxPi2IcxRYMxmcfv6AephhHE+sP4LpY8jf3s0nOf1qagz2pihda8LnN/lbi2MtIgdZ+9dm6jaiA
XSjED1aotAg7pUiXd7it1ryfv3428fDRJKEZ792jIYt7CJTWu12j0AMPBaui2W32tjy5/VRDDwYJ
2itXrOQxbjOdDFDX7pmV4A5Li+1BeEQdF/W9lNbTBhz0hujPe1UgJ/OWz6oksLzsmBuFMiiZbPmd
JhyShOHw8SOGc4M8KADB/THKbG0L+vUISZz4uSYHyUdvim8j8PN+k9NEfPM/9Rxfjz6lsdR6puC0
Nxm34VMEGBOUzqeFTv6f4oU9AT+FCzjlw9T4dNbhK1Et/XZGr14tpJkH368QfFUTINIkLFut7m2k
dC1Adh9DvxPduHnDbVKTKQWdS9nRZdZcbNU2V0Mm2SUPBypowpitpvdVa9JUWnPleYrXZu+7B8VP
kWD/DyA88iXDqgpbzKwxRZH3SK55DhTel+DZ5fHntJf9fXAuSbMRv0IJjPkSXA4BXIfqr63IGMsV
7P0DNAA+8BUXxulYuQg+ahBR5K5TqRErMIcXvgQ6uls32W33CEHRvkEMO/nHdakEWkmP2ytPtCpn
pkRLohfzJomuJO7wWa0dbvXwCDBKVKBWYpEuqdLVYFVI7piyfcztwzZShlOfD/WiRwF9q0Ynrmnq
xZEilYrpblS8/WIpqk7WKydlqOAo8lhRWXNHbXHuFiJtmaYDkPQABLhycv/7i/t6M6S3eqapLRIx
ZYGLSwTF9kAZbe8L/5C96JPqVmjQZ7xM5seZ5clNP28580d+0qw47vWY2ma5G2kP4xLUtwOISilJ
E1TyviOOyIMK979IBsp+KE8C0WY6Fs9OYGM78ltancrdIBiQ2sw1RVJ98VhVv30gQ8lCChhIoVfs
dXp7aQtAwmfs5K1mzYtRTRT4oZh8h6hFrS9GYBog4FIN2A7BDBVXO38lVJL6ZlL5LjDFWxS4Lz/O
QJOxQGkeJQJd/IPWHvp4+FHcW0cAZPUpLQFnLDL8Iz+4nfxnvjNszgLKzScoM4bC0rH8gngsBR+q
AqX9uKtzIaV5Qn3nhdFnC3XRhZ4wOJfPGg4cBQu5E9mKux1OxKmV//7SyhlmAe5gnhFF80iU47fH
cqnm16v9mPfuzom2pAwwLXCYR9RAMsL0hVDLE9cS3dwqhvFE87r8MPJ7zshx5AXsePmNC3vJH/4m
BRb0QqAIOz6bZpLtLmflouzqWkqN2nTTzFWaQDCrJy3VITaoqUFgDVS+xzaAje2/esMD0/jz/m3k
AowL/+n8bCLO3GdbHnoWw8MhnSMYmHnEsOj6j0PO/0jZDE8pXGiNLnDD6qKgYre6t3VkRjIaVeBw
kxNYLe+NdTpp+K4+pPTLN4mHJ6zX0r7cW3FzAsvbBFxJ5BgQlSUI5JCz0dmsPe4B1GtLMx0cxHf4
sqDzentirPb7MraDPPns21JRgPyfEupkqQaIhoff4/X1BIS5ESvhhcBbetIEqHDUDtaSLSZBfK1N
85p0JJ6DQUPW/9MFxipBKVe+VMS8GhvyGji2bSO8aPrXXKR1EbUR02wKO1QHHyeN8csqRQXnG9z6
0RvJwpAhnvxUWR709wmWeH7AvklZ6htIMpCCgM/2bNK+KHV3b9VSdwyhWBpMr/OUfWwEEopzr4+C
pvQ3iX34+p7cE0pq5qvKJPyYXYRZZqPBg0lVnqMSY34KQACVaqblqPkGrtagrnx58Yv19KhHjVDK
OqBqQO0Zj3+ka00bI1vbF9U8SK55PggmKbjOqmruZraNAWA0Q7gSY3GERe48U5ueUTAFQ7quI5RN
On3eejHSld2IBubiVptryjazN+1N5jv+5u03DPtynTOU86WllBogbSPAlYnwG92xEQx/jDR1ZaXg
eM4rxzNoae2GFAcxNy1M6Tut0K4/g9c5slMu5GJLeGqQTsNzAglXj2ar/ZRhQ4ia2MuKtYHMC9km
N1KznAIjlnhIdfpouUpxGBf0UTaOeebpJNZTKu4GXWL+qAfwwTHG/QRrvTKs/5hwimG1p1bIsFVu
c9fzoLuFqWFIHpHdYthxCBg4LKY/FMibPUsop6N41IdQnpqVP1EVyZLtuTEll4u1PrwRx2wr7vyy
RjL+8e3+2ahcBYajoK05lDiWL5Bar0mBMI+ygP1HbRr3tK2yi46G87OSPHSHMsC1nMaqoBwhzcQW
qBRH4JM7XT9EaHnhxCv8U+Nu4NfAPMC9BTRK1LcTb3binVtLRdEuDUMSCNTOzKJJIzKPHvfJSb6d
r1fmB6X8Mckr9NRVwVZvSSNdCbVv3T6ZDn5fTsOnOFvcmmNEmX15p3EYpzt4E36JkLQluNdk6hhf
uosqS2xLdyFyprH62Vm/rYWCCQ9e26Dbq+EebnLubvO2d3zORNl7I5GO5gqPLsDhIvHYh6WgOLjE
5N/V1ajL5lQq/9IMC+11Mrp99Z7hD2+AQ6L5M/cSCFz7pPzre60TZrKUKduyiAmb8pZk1gUzJqTm
AST/LkA3b2aPLmMrX4YbKWFUr+yoiN1PYegvY3nNZ2Jwa/rwOfJKV8g7RdPBxLnLV2zKW+awil5E
WnKsEmRQPEtUQ0PwB7oXQDoEh7ZMWwT03uMm8JWO9x8gtjwy7aZB4cjkJi/1zdMhlt62VYhVPvMZ
rqwLERvhOCXg/g5N4QDVTM5WmcttM1Pb5FPR8EkqdjesyvTC+Thx7KxlhMuTNBgIvQobds15xDmm
Sw3hrJkrhZPtA/CZdj32ul+mV/wMc68sU1T0sD5jCzi/VN0JpzaLs3EIjiefD7So6dZl2XFj3VrR
hW3DyPe8Bn9lQRt1JIGdTDHlS5FzF1yvcBbXUQrdVC3/dTCIq1IdZ223wytBN3FX55sCAENmeaYy
ybAw9v305h2e8gHdgwVjya3coGdBxQ2zpmlEvXtL5+9U/SW8RzGNGA3yjwilcqLpuoiYDDWXGY7y
NRHy5Ks4n4JVU0W/bbYymlhw7bQnsDiTo7+WU1TODt+abqxjbL63eIKykBFBmRrYvBxOZaDU1pDr
l3J8qGEXaMwP9r805GwDmYlGOWj/YDcEezLQnR5INGnXorullTAPCaOQejZCBrtx1l9NkXAEf8jz
3dKVd7/9Q+TY1Fg6Z5iToAF5fd1FchUmLw4ZbUNj7Wpzrww13LiJP+y6akfnygl41yEzVSnjzcRY
c29klgBGXbH3MHR/mDbMmVaY2qcM8QZMOdVL6qnjS3peav0gtAXU/h1xr1+wBr6vAHLFfvSWEyZY
2NisYNd8SGcB02rVydQkUejO76yFprVrF4bqbuhkDkkyOOzLuUD1f7Hw3PoEKE78jKvnHjgPdJXC
tN+oCKGPZLNcn2tOWanMOiiLJ832iLvjUTjk4VY5pBu4pFkUNKo4h8EXhu1yt9pWb9yBLEsXTewq
lwWHc0Uoq6OWbq9IABUP8Wm6rxcA89R1r2t76fOHYVVwrfhFplQaWvJlTJ8Tjoinnl80UANdfsq4
4atFlG5J8SayIprEzY2LQrwC2ByKMsDTvOAXnw3mKzEw4i7FcFJxBz9+BcfewHFB/c+m8z5/m1Yv
k5TMEoHG/8qd/WGGiyPyKHt9ASeHqAmGOgs9Wd+9M79hfSTvKBVKk6EcXYqoDokqqWVo5iJA5HhL
MAZd4y+LRyNU+wngCztJ5xMIZcvMRzU8vFraLQY4sGWG/BK6qFmAoDYccOh/qfLqINK86tbI4qMb
zzri62elnUOBO8ITpJFELLvQDZ5liiwhRe+hfcdgKm4uEOZ4m2W8tBYTMP5+9Z4mOPCFXTZKbC1m
fKYbgNYHaYws+AA0DiZLa9zlF6nSka1mfXW5nhTk3PHBSBsB67Al/ZIt9m4gvrJ8L9ERntO0Dm9D
SssX5MC+8q1di27yU8sztD70uSK/nLkEP5C+0zp6B6N5E5+oVoerA0zendJjevxtrPNu3b+1bxXk
JlR08iYu1GZS4/f5iy2Plv6tB8u4PuT3tR/342eDxadNU0mGnF8dk7cDAlNfgQPzUgFGx2mNpnVL
1/x1w1NBBpM5PTJHAKEeKCeEEV/wanyvj/BHWrca80BH0+3rZV/slBrLUiyLG4IWdvV+kReoRlvR
oQtgh21BZgIHXbNaGEzU930zjNdUBrmnScRkVfLQEHU8du2TQ+VUXnRqS7TtmhDAQ2sphRbltKJf
oJto2/5QEpnUllCq4ObTxNn4rUo4x94sPOGnK65KguIDDD/FZdP7bXGq0fuGbKEhdzwnsjo3+iPs
zZQoLjDZX94kSSTuLpbV2vN1jbhvHNI61qsONsodoz0BlhPKkXesvwsB4nPUw9CvIXF8VHQZrJ5W
zoxs4DlddBzNvcoidWOs4Me4hG53gwUNLTEwoW3JnN9AG7FolLpCra1mt7C6SV0M2ljnwb3jvF4M
duflIwMrYOBYTcUfBv13WQ/jWLFd7Bqy6mY79l3gtrUBYpVUfbDJrT10SLpJpSkXcwIQoTnBlRM9
6u0iaggrbtyeJWad1sbr7AxTR7h80+L2zDxHqGGfHJ5sxNpn9JjqkAA0Hk3N6/SoLESoz0bfrLHT
XYXG2peYXPir19ZcKRny6ybt3Pa9iN/b7LhQ3dzoEPku94q+R6B6Xqlr3rl5R13EJyu7dJUX7B4z
MzevFfp0+yhoXKBfn/bmnGLOXwfBzD3Y1dwsov6ovJfPAA5tL7i/DMfz4CsuGcoa2pT6U/o6rmRy
G1RXMMNpj0SDuvnD1CCvWY58uP8y8V6/48iMgpRTp+g1rvAMETC3TwFjMDwFjtfQWQD9L6PQGyHz
jMYUWNMt8FyUJmdoEUPD6SewITQWmOthB6AU/7nM6XXhlQ9bpPGcrnEOfHGh68cQPw5M+/27lxpn
Q+wv2EJdkZ7ZUuR9493x7Z0S6LFa2zWVs1hVUKGWrD77gmeh0qn0ix3pyyijQKMJZ3H3dtHXzRJs
IMnJaGgybFRsx6qZUm2/xneLuZL/jNQdFJPhNfiHf3njegwsxtw8mgNRl7ziBwpIZ/81u6a/43gb
Hoa/EBMzMZH0qKmcKYcMkYWRLqkERG+48ofXbnUYWTQKiLtFdc0juEEV2Kl+VqsJd5GlSaIm04Rn
qa7PeixHeEx6eQtI7OZl4VMZQfZcdkwptmK5bFWaSZ6GuuotWH8BRX7WehzzD2mXVsoo7Z9CZW01
22L/esnZyMslEFH9xm0ZjuCWGbtsLTqXme6V6utWGwGGn4kVK/6mywCADOIyTXuahGYDnI9qrEh7
fDdqr/s5E5ZN69uVN0cpPLiYjmrC/vBWYv+xqJiTXy1/WFH9He8gQsyS57PTsnYkt3OrDNd7EB+o
AiSzOX96bmRthiN2FeJdu2mqPn80MNwqGFFE0k5ctjF1R6L59rX2VikUsiYkPdmUcjrV7unOgQEi
xvH+y1UUNUNLS3dHbARNOocET0PKvlUOabwhbJzX5OfiNmm3IPiB3XM81ZHCQijhiUpWlFTRbGlV
x6q56tevNHXle8Ye2i/W2ZuEOX2R6SmLGIV0Ikdy8qa5kP6d3Q7p/EAfpUEPKqrlOsXbQGhKgew7
Ex7SDjNxqKwG6sgiXajQk7jAYm17/aGWmoJ97hBK59adhASgUDb3GkSfdO1B41fAeJWaTAps7gq+
akIlQTZh2e5YzMiU5sz7PABC+arClxsOtywIyuc9rsF4ipFJNrC0HiVTQ3deE1UI4s1mL0H3i63G
9BDONJ0cCBVWQjC/E/Jxix8awHOVJhX/Sq309MxoGV05synhRg8OorlmgMMFAJ4AT6ENzhd0jWNv
wxWE0nGVmXgzLHz5DwadxtbGxiOJ/woaPLVOhdNeBiCltE9ugw8puBnsb6/Gg0asMn8KvHYZ/i7U
7kkxAyxX2zm1nmG4Bb8MOJg8EgGTGiysz8oNouUpoVuSH0iX3T85iBaj/jVIYAH89rKZeW37ssv6
W8VBLQI5pkdQSwtIoSPh5KHOyhfEWq5rPKCLntUsETwp0imP9RpN70r/1DFHYnXxsRs2GgP4VNg3
w/lET00sa1f+4MhL3AookJ4cQ5I7Zw0FYpVEZFcvxiTlEh/xCfWyd6Y4sTg+/bCIw2rNd2Bw4S9T
jkeGdbQOj2DbetuHrOnmk3J00v3Pt9n4lN/TCFteWU4xOVRhhQA6veW0UZBGkFJO08MLF97NWVRd
WBNI6QRWnNNrCo8XMCsBE44UdmKUdr27WOokMv58m31lXNNpq9s5abdi5Tu5ayj2mFou2TfU6Odu
WE+NzwbGeCopgbro4qczSs6m+nRYzxubNdRf9bfqunJshrrLae2zeeoZctihwywFMAiLjFqMmk3c
r3p9fVK08kIj6+r0NC7u76YI1p873hD7y9Hpxoks5O+PObuUyq/Dri/B/AGNKTTnRc5OeQSDxC5g
xdNNeO7XqMI2bmnjWDGOekjXJZ4O7NvAQbii2HcruWwrX3WwgiLkUgzmieBsUW+duShfFo5q0y+Q
uOLZ2LalTjprn4IZ7Hg+PuxMoySUFPJfZO9ZErqeOnG7+Y09QQyU3V/WHNbz2LwAVu9mJ6SNwEzR
H7+9UfHmIje46TCrT4YDIfvxZZTrYOp99IJhMj6ngWmLHivuzH1CfiZLYnpe+AGpfKapsm4PlJJ2
BQqheYIRHooSshcywrRqu/qtorHHdPYRt7ZKIIB6rkOt4i2PEfqR5bmoR01zjtZzL+6GqWT8dwwd
58/XXc5kp6oNR5toIPZ6rwIZ7SC9Bh2GVCYXfXaYpgiKPa/4jMIrUhx5PSUa+ekLR8jjhnvQekY8
OvDI0KX540Oi5h6+MVv0O7M4uyOMNOWyDYpoiTfC/LL89/Ofk5DjMHV9PjPWDe4X6cxc7PM22yMD
iEKeJFNDAtFG1WIizsGm9GPxcb98RU6nMrZRKtF6HtnfRejCG6UugiyHzP3d9304u6NrMNRgzLnX
oiRCNdi1yyUggIWUVUFQz1ttHrS2GhgirVHIGfOrrJWlUGkt1qbLkUSp5i7rLVpokMGI4BJ5t12Y
vuW3eg76mL0B3JZu34M+WUFq9cv+VdXuRrBupZGr1BiL9ZEtO5Hg7JmgwxhVkS0w4TEDwl00Wpbb
RF2FMsR78/se2LccC6k4Pvl8lOTK7mKWIC0A1t66hsr3ZlsGrd4INBRn+CpITtxnMOX0Qi7Z2A9J
Ed7PBMPW+klDT99kctJ/mh51T5M0Y4KcPjz0Kn1bWqcF5wiYucK0QYPNuwLFVavM5XJ4Jw+dOxB7
rYzl6746FVYnT3YQ/qGuZJ8swJPT3mXz4UzJZW2QJT60ZQqtlY8iQ0V89Oxo9KWIoIXwHo/18iAJ
zsSAQ8f6V8kZVqN1V0TSmb435piQm+Wv+KTEw0RfZVcmgF8whKbmQAy1SJJzw+QrscNohfbar5X6
G7U4oz0NV+HTm/+3VOb8MbYZePr9pyXrs45+aUajKIJrtr3Hr16gQTUET3N/kFtp/Vv6JVJMycdw
k/7ZJZBgvb+OruIwqoVUqJz2IPOZH0aM5T+0fUcNIOsNdcl0lSsvNiyZg2sbTNfAJYxDehU3ruyu
d5iwgED7Cka8eg2nR49IEatf3X+jqWeU+X8EfTO8CUUG2FbsBoSsQYsMCBX3PHYhl8/Z9m+5H2aY
t6/KVmaxKbNYMbjr5ejIUATCnLzUeUjXeSEI9zTB+ODcd4rzdwLX/rHNrRYKFRLsZ/H7poulnwFu
wYD9i1j9DW3DgOJu7f+vBIzci6dMAHbgFW8MimIFXz5fzGmdAjLllQQL2RMxvmkWpWVHlQHrUy+p
okg9H3xKFfqdCNwDFIkkuXO63CVhx7Y7xqzKYvYH/QjF0Y+6s+f6j/cTOJXOXAJV/GB5xk5MGItS
Ex/Tm46zUknpAUswWzikFAxZhqB2Sdn+E2ZXRuwZIPWgeVAsluRtZX83VWtZntQf3XaBEOcEf1eE
kh+aMiRinW28lnLh+vR2nLPFtHXdLtY08LC7UuQxTdfUXm68mUNXnWsNBC6uNZYt8D89yhAprQj1
cp009T9TmJh5QOVQ9TIJFj0T5Yn3cqkdiIS0dB1KE7SD39nY5G9braIew98Y/JybrQtzdA85Wp1l
Q6lWdqH+34d8HYULaSEB7EukbsO76+LZurl3XAZHBjttTupsrorpSzIKz1sKfJgohRt3G/vq2Xlc
dyGCmfXKWEslq53W3nqR+tFS+BehJzSNmxv9+laXjtlHp4kYBrbgHS4ltzAMl5c0suy42dQey96G
Bar8dMkhSBeUg69HOma1M8qtSct0R+7OLuARejAptYxby1S4BOYHOvB3UuUuJD4UstTBoGVGI+xC
5Sym+oUC7Dy72mu680HiS9DjwqAa1OB0Mhtn0DaOpmMBAjJpCVonX0iBIUvfwAp3XkQ2IhPEwZZN
HmGu09f2jKllt0HqkLx2RFmhOf3T1bZR3JamiVrfM5dwoXohgjgHBKPiaeN4/QsS97eC7mVh7fup
BIJ27EwxaondpBXE7XvEjZYjL7R5GsFPGDG5uf5qlViDwwwHxpp1BAQ7p9rkvcsszyFaZTqgJ3xD
eaKZqCe8LH8gqvGUzJiF8fICaLN9RZshAER2VTKewz8ulKgRFWdgmQsYEPPvNGrLTREWwDNwDLyw
OU5lTnIbpf7zcBj/th+1hFUN+NhlatO3ata2tTGaMtBZJwLLNcb1rg0v3hnx2KOpG+D0jZk4LtNZ
vc3/dFXXZOUQKmLEEtbsBHS6rTZ/ty2npuenhxDwSbAjpY4gOdBW2SLtg+81CATuqNNYeynqnH1/
Z46IIjm2khW6OATT7BZdU5fMOdy3gGbnz7XV9wBtFJJCuvJ/faQ+AI2zYFwMqj1qytFR3x2G6mId
4euSipqYKAikB7JH1eihuYXRhQ6alj5s2qUFNg7xDKUdqcd6Vd0i0So5ftVTx/9YkD6PhhF0EQTT
+Rr2+a/mFYou1ORqPXyfvVtE4FSyO3DgjlGUfEcJs+54qJVNnGIR+Dl4s0OSLdUMz5oSmCXUqIRE
q4eyeN4++KhkITKsMz0GuTSGw5kIhm3zy2Tm23YnDQq4UnuFkI3+67xMkRa/jZsNwkGSc0PZUz9Z
UdmXF7I86Th+S4tDCiUBhtHFsmk1s0ep0J5XCyviW+EOmpz51At8Y4q9p3Wa8mClZWg2wtkWCqH2
/NgxqNV7WtMA0eHhHY/Ly6GoTDo5hkgYnJtYA1gTcB+CKRZ6xXu468SQ5ldeWRQWthol4Qm+ewRX
5ItaOKpRyqi4ddlyWe6HIgRvFoD+pkBZ3MPA5E0G9npdry7WUQoubR/MNqpKvT3wZ1Q/L9UpPdGb
ZL4QrvKeHoM1qesjeM1BHkFPeeyciX7XJAsOrLDN8IRhwEubjz/KWJ9LVgkJRm327dDNULTL1Uo8
7Hi6T9YEM2d6U2ykiv0n6H19oZrDGRgF8veSvZ+uP5yLH3NtWJfPOykNlVTQM6tkJ/3uFOzA3i7z
C7OahLWXBHh5NZtV1LuaHfFqNjB0u8eKaMyWkRf/DXNrxYlisqvz4BFnqGrrqP4UMnIQNA6JgF7N
mcWhBWGy/ovt/RMLzjCpTHBAV3fWT7z2Un06SNfHTLgSkMHstmH0lWpL+H2F0CaKiA2DUIxbtEfF
7GstNmUgKHozspbaLeA55Jc6HH7Go3PbqLU53HdR9TXcn91TlGNX8hGE8iYf1wHOTKMpmFABBEco
JMk7qlmee/iglv/hgrFLrrEU8MqZe++YdFRGnlm7Wm0JDbfCJeyn02n9cB0OSl0Eh1TfJn4SIuy5
InPSSt7/yspP84brL3i5iJ0nWnHVY9SyuXhRhy8lZtYrVv+J6jZiLr4Xa+RJUQWmwvVH8PveO7e8
rXZYAw/+qWvvNRUNUX1Tm8bTvcLJdUiMH/gVT5vpyj7I1t3pPbmoRxHwrY3YpW9veDGwfSDcJPRo
0GuvdGTh0tFgKO14H7ZZGubQWortcUaeHSDdjalatxl103GRaZ+T0I68Diw+ygmhmleoud2hYy7/
bDRSkh4N92KxEZgi+inexqKKpeuXFnfPDxPyIfyNKqUwXKGWjbZGnUQzTv/z7X/lN775OeALDTuU
U4QpaTGuCw6EwnzlcDk9OcxJ3MF04I1pPHdInG4H/0gqe/qa6UUbPC2H+jcURwv0XB3Ow+CFbzKG
Xr2tAZOIxaYVqpdvbSyRrdO+nCowEDhXAlnvUTTIE9HZhJNJyQI5qNnbBFYtTKHjcxWJ7ybbqmCc
7GIYzsfeHsM5sl+0rc377vRYsUSpTMEqZqfXiACJfu1iJ0U53dL/T7Zj018Um9AYgGrPNMmsmek6
QlcH3Btp1ybCqFYp/nNdQGdGNRJcKmKoYdBeF/xZOEaWMvBtdVuQw4tWvO8fiRGEtdIrtQp9yX62
gP+jvPWhwTRJMY+1UaeyzJ9Y4EifjAkAg29aDRLmFlq0kvqS2DDXXolOsAibXbMVvuZilfIfCji8
QCqnwva9MVtB89Pk9iBoFg97bZLz0dPH51smK26dXszU/hat8p77n+OvxswYmViGSEhrHeVCs5G2
m74xlREmTcpFbNuYjmeVkgpbT7vtA6uau8sfpoPspUQ3SE2uFGeCJtJdZQrtrxX8hspBr2MPduaI
rWH+vbvk5EsYuBe6kLLpT97dewN2levV+EgDI6fWVikTqR0dCTqa4k0On9gtciqCSOhPetRqMmoz
B4rfYFBpZq83yBPKVRaXxLRg0filqlwsgxPZTMOkEB8E3pi4frLYTW/WGV5FfVYZQYfAWsl+COeo
vdDoOZIj3zOlILDZqSQqQ2IM8QSX+lc15ehHX8kuVdPfDgrr38Yo8J1a+QRCcVcYk9gwQf6M9LOU
ukRUtZNAWWAcrzEmJ+RsUOZR7i0frpbFwf3WB8nCVBdrJ56uO2bOJELD+Pm7/Q3r2xY0bIFljcaf
NXn+Y6G9SjnyIzxmDfFcq5l/zDnOrZB+trAaAG+IqD5nlZbVFbK0KLU7Oxt21DZJpbnGC+Oc9RI6
TPfTFp/IbJ//JpIbvoOxekFnt3fukvmkg/XzxKf6ZC2aqv8+Yzj4DF32m5zuOAarQvPzUXBdw2Uy
5HWHpWxSEK7uBvYzNomZNcLRGQ7kSnN4puJfwYnJBEfE3Sm7kwCbjNtVBujwqUjH9nzABmYrLplt
JucitYMCTsIaGwi2pIBIOyiNsGOve2RsXgHj4uoy9Qf3IC/KjgjqnnV4ml+4pj88cNTnLoleXUGS
bffRQO8wsCp5UiPsk34Ry3Ahq7MZYw4FAh2mbpaR2cusvmWNJT2aol4T/G54VGde7zOlk2A3jIYA
tkB1NXOBzXdiZ0qd0Os598D/SfjOEsaZ2mxlRwLmyHhf+/hGM5c7YUM69v9eymU4QU2Tm0Jqr+kB
o8chiZIYqOOt1ADR3ectGplqOeHv1LMOcZmxQhNphLP+07gyaHU2LthVyp02QsQ4KpYurYtWYIkC
UX4ytKwBA+IOyMrztrDyDBb5bJEoYJGN+GmmVfPsFALBAv1VjDhPXsdM1mPxCLbNgja020CaTC3G
rV5oy6k+saVpdqpmHEOtuh1d9Sfge6LSq4lZqqvwAcsgI2aec2AU72SKZzv4YMtAr2bOl1wlP3FP
YB83YMgYk7Re6OBDq2QQ8k/jsjujFJcgh3MdEgzwsTLlI0OWkrQtMXegPqz/oZyARotmByl/ZKsE
YCpu1sZIlwWfRSPUBXnIQp3vLzOFLsCbULnYziXyu8vzn65js8YfKlezcAFZ5DXUtxE8okkhrpK1
ms/MlGvnQ0vTkCbvW8nuhH/2oV5iOJ0RXfdbQcBUdM5eoCVBaF2Af4EXFXZTiMEnpPWSp9LJbnF1
i/aixO42kLwZU2uMa3CS7UN2saB7AztT6Mh6CwbTkyH7wXAa5lERd0ejg/GY1UcHzOW5qunYfTx0
J461NpTqIipGXObpmi7iTux6FBFYYwftvJ6totAY4QzkrqbsCWWrKjmHB6HGpkxWchGYxX6lhMQm
KecINYyneFc6ITLC8TNEq008jaVEPobLmQdq5BshVNm+zOyxAW5Cci15YPTcd+mCgUH0IJ/6LCp1
UAGKJnJFDHoXhsTXMhEV7d3EJbBL+liTeDc7Rq8yWn0OJ+kpIcghxX+hk5NJJLr1kQvvLm2FEbEN
f4oC2T9ut6knGtDhj/Oa4szaYrXfvriYYmJpI2m0Y+Hr21CgzLN4K7pTxsHNWmBiF3L+GYaJezY8
M8DJAWl77+Vz6LBoLDNwoWiKuIRkIRx8FAugnVae5XGPBe4GH3xl9bosh1Z9N0dT4LsSNfzF0Zl6
ME0p/oPqWqxspRXnIuWnoiwTXMVeRneVaxXZwUfdhaq/sKkVDQkT8df+30+hideXP5HjXSPRQmp2
ls00ONPYv0YeFEDphv5hY/b8bq0ol31EBW/zqCBZM1FZUrJYpcx6mTAnZxe0ixRTn+RDeJ8AiZ5k
bRMlqBTEyafSBISOm507R/l9O5qRZL3D2OROYuhX0xCVhE68G+D/VLdkAlqmStT0wRr39kGAxJH/
4qGJ7SP/YusMoZoM2RIV8UuWuodixPhquzSygYvW58yMTpAvaCzRJCZzSv1Q6TPT5j2ls/wSL4oj
6OUb5b49Ekq0jIUS516yarclpfiZAdlU7rfEfLQvocSSNwcgftDKapTpAzGxPFfR6PuJVIG6BfA7
QuJWlZ6JXc6gBU0Vtn4gObM3BEFkCSFv+gV1hIzvdHIOAaBvbxueorWoE9Bpl3+GgPBTWbaMxafF
I4wPstA8bOLrH9pIhViiAAkAJYRwp7GT6/P512aU73bMh1BdzRHNin+yVXZd1Dovk2luI/x8FAC2
/XQU5YQKPwKZFeBefPlypRf02cAzEgBhDmVyaqLViElP42AvPu5hMEeIdsjf2wMOUkc/1JiqFhOM
U3uPPhJ3eDzJOCoCZvj7OufSKSEqSTF8B2AMVnwKpJaQw0UnczJ9/eewbeQFAUE2mkNWeb0bVKjf
SGvu7m8yjs7wF/A3EnAr4GF4URMwffka4xwBBPpJ+ySOPOxcNn7EDkOrvkBpXH8lwFAvlGm/18Pu
PWEtOslG6vAFmRjNMvH6udDYfdZrGIZHlJ/e93RruRoTJbBZa4hG1qqVRlXL9ZmYlz2RAvulJ3fD
vUlY/M9tMmri9aT4LTF4a/w0IFTIrXCtrKdmmIXOS/g9GQEWbptDMshHBQ/QuiBsHu06JEKSnkK2
wAW7Tuq9K0GRaDG2TbPXKjoxoN335qffzBX6SVWrrVLdUt/VYu/r6tEnh3OHXM2mrQfhcU/z2HOd
tM2CfD+3CJ/eG9ZUSC7Rv9CeBCa2pdysFkUZt/ZrPtF0w6VciXU+D+hnzf/yNynTeaAHBm5kz3SY
jND9nKdQKrvPQNCb/jydD9WQdDgdMZV6O2DTf1u6EDDJ7tSOpRlQKL7NEBTr25p5ZgDX1+Olgban
K+NNS0HcynyodZuLnTGpek3MHT9kxiOYNQdfj6v4Rp/7fy2XLCSKONa8gv7M5M+7q1nMvLZXvEgj
kuihFb7im9hEoCjMtWTHnYMPPDYYLJKQpCHx+PN0Q/A7l+1RgMHuCgw89PqCwS+Qw8tNCdGJsAuh
nwf4IbeUACDSz/SLRHS4rAcAvUkkGmL+u1wLkwcML0e5LwWUUgleGTx4onXJ5jKjap7JbodM4eon
XjKuK5jRFey7v9UOtm54zNg6IsuGASexeGfbZUFWfPTlnVT+r1gQJpvth6Oz+cnzKD//13CppQHT
hcm2BjCnAdQ39pQwUffDBGgQQ2lPVmt8y1TRt+TIWLnrdeIZ8/lRf9I4jT4CAM78rlErrq8vxOJi
wktEk3mfqf6S7qu1AV8ZHm8tHMEVBhJBV4wKfb+sbczmOPbQOGPrkINYPbtPAP+BC+MFrofFAp17
eUDJ3crQw6m+8YkE77R0VMG5raTINe/IBJE8Nb38vdAC+d4JxRa8dDc3M8Y/yfxE8VXfPbATbUSv
dsehUMB/7kBZHI4ewFUUPcKyAIvpFBQjNtkBGkpaDApmPicEBzuji5eM1qwB1RsqBX1zUMIQpwjO
z/bmwbL78sKYtx6wY1BaZiqp2W6R6ZklS5J470JmKtGo5O47ZxPzvexYGjn/4PUBkVXlBfr46Tjn
jEVBaUcHlYLD1mv1FxQNXZfxqrR2gwdql98lHKGjFlzh7ke+/qg+R1IRMHhkwhHO+hlPHJ7BoQrs
0MKz83uuEx2kjWZ2LNHnQY1udH0b5T7OEo05tbCzIlVtJHrI/2sf0jSYq7ZWFcWZ5edrdsMm0Acx
JMlgYNOYOLgK+8ssCls2zlE4ykgq2NJqLJKNb5BFUYfK3a/AzV/9y62CKZBn1s230nTptZOi0QpC
h9PYbRdf7yo9aoyOobErkbYnE4bZxYCmNck8yUOfxOXMopq2F8G/dDsAY9hzSrwpqtg7K6uRlAzs
qAdrB07NniaORoC+2QT0LA1OxXDfatl4lH6fhHgt/NBdTscAkoiuzoL8MLhzwZR1T+XCl6gPCiBC
N/RIi2XEuhLo0+gdLHRkCh0A9CGE0jGhLpfaNn/pW9C25D9/fjmVM5zMZSZp1IrRj9yDqErN9Ovu
+U5LcKEF40Fq8T5cMNvhEdxvpnuoBCFuTkjr2PUrmPDtWBXjUfx4Mm4VDR+7LS68Eq1tU/STlYfo
O18EC6PYdecagOo/akQn3CwS0IZdjZbXJKcE7zyWfDO0JlR/6NBu4b0AnCyD1HsiVSoMay52Ce0T
azWFIUmVin9YDFREhCG9VBH3d4j+9RaaMvgd3OjxPrk2z3mwoeVg8C03JHr6gx/kvQYv1yVRfEFi
srmi0iTYVnC9kwoCyFRHip1Ufae7768oU8eVI1/hKmWh9UoWxqqAJ48GDpvitPAwrEbVyJlYFSb1
SpWjsOikn4zJ5B8yK8tZDzYaHC5XdYAH84IWc+yEeF8IoJCGa9AXe/9nuZ80/RlkC8CFg7UBV9dx
bj+tXsGHWwP1kuq2ilAEwNcY85KLk0AUJXa2xDC8q0ycZCzz524TmSRhHcJ/1FTOzcBU3D6yRbY+
SOV+8CpoboS79EckJiQslJ9+alDT9mmfLBFBq3CKAykHFFQVt26j99PFmjtDNAsKXSUUvr4cEyW5
qvO+v21swVwPth39hAK1jkIBntBX+1eiflEAADj7NyQN9n6ATImS1r7TC83Xj4J76Q4z1GrlZmZ5
G+9HlWKJdH2SKyDP6KkkVjs+GHp9TQK62CUTgSVWRw4u2X3t8p/nSEBFTVufY2mknaoojHqGSZc3
FbiSgN1x9vIJNg4qdGYL/k+D8Iltz+xqNHMfpTU+ZR6wxywDzimUESTGmfHrgHH4KFnY0qcQmy+o
jfO05EqTvS+syNGGmjeRgHHaTl48YF2xnYQKt1czuDy91e9zW9nzMiLU1NVWku1TFFhfEfPP/NY/
Ofe1KQRkjpcS2qGxrg0xtLuQA5rYVpxPXj4TbmokN+WuOm/EGhR5CveZ0ubiw+LBH+m28s8V64Ig
nfwBWdXgc7BbnpWINFYk06AVMMTiLOL6x0il+RIoYmi14ac9uHO20jskApkCOXGkSozSLsP8kh4H
Q5uLXI8jRgGxSIpSKK5h13rltrVM8PdkBQ/b8PYef+/OCJZ7KLZwsQXinvJvpQB2clfhpNsiryv3
7Tl5RPWDOnyGcAZ1iQTZJJfMUyR5hg+El9XTg+R3oYlxrRFE0UH5h1slmJA1Bcup6WR44ZpSt+0n
Y1lFgsRhl3oV+NSljzXmn7/WhceJNFwcdXHB5lWkvvULTcar81CzG7SGgWu2NMghjRTs+8Xk9ONL
OUB8nNkCupDQzaDxAv+EsRTW4TFhjnTx9WhaIrnYZST1LklHl0kg8UAtTZi3UmOH34qPmr5y0unM
Clw/kZ+y6GoUSIdRzYOKxBcX2dxvbhUBEjsy0+zulWnVPCnGtKTBLLDbExEEfprBrmJhfAzK/WNc
V+Ma7yXhJBiMBDEmXr0Xr6UrVzfl68OPE0yh9DjQmkV46+blITE0D9Of8Txn7iBj2UmLb/lsMTFs
zTNbe35mybkqBAZ6qlort7KlHTKAhJm8sMcsz2iYKKh/1sfvvSffwkkZyuYSvZKQf2gVtVbzUzMk
s2rFoOKxV+YgXNUpDEPFIMtEWBB47ofiEUtym7ID3XU5abs3mVP7obBzHRZPyo9zz+DcoXA8/8mh
4CZI0nZ4SRIYNH9eGA6K4PJXiXDoFSTc/kOPd5aYQH8fUBphdkj5WmVziqH0G/p0R5iHRPqdx3P8
BmiuPMIlI3l4oErdtS3e1IuD8b5C51RKr+QNKz+vs83ScSK1hfp8UZ5x6bwlGuTH1F7+iRDj6TwA
zyH0l1NvgVhTmCu6EUrbE/Qpbw2uUQw+cPw7IW1vTRJx00nVM61O7haK0+YufLy8oOSkWbwxBMDY
x6JmKLZUmI7Igu4tDVEGknpXSAuNwWAm/X3m2fZzNPYn5OvcXJWCiCnsLH7LWFiob4O4zJ65OcAe
ux0FhwG/MTt1vALJrPU0E9SKjJT4sBdJfwTpi8h2rqsIbmAMzbWl/m9Zd/LpNRRJYH9dX2h91+xx
/GDywmvHnChU+9qQmK5nrEBLkpC6aCgNeMjLfYAjoNt98jWSg9PJNn6otf3aTBTTox3r+2wbekIp
Wd8rEXx7QU7m/lsMNv9HfAKTv+z/YlTRo6MWkUfklRV7hIE1C/gjrGIsI4582XqVMs797Eipx7ps
eXyXPNNbjF3jdmKJDjCDm8xrLwgypqdYv8zuGr6+M86MC1uvxGgN1TzIRfk+LgyPojYQYZjYoHhm
2NELu+98QbiDZB/+HVYyhmjzXKfuLC4VylEr4P7wcqDQQ1VqXrWC4AesJcOiB49iJqAZv3GYn+i0
NRQtQ79nMUJ0ey9oSPSYxvDZ52P9PiBn4Wd+Z+W+LJob/EiFpKotSViYRkwi50R1HuzJQ5UrZ5HN
jiSB2X5+ugW3TC1fY3ClMWlOri+7Zp2YcaIjwvRGWiiOc6GcDeTEZ5nvoIiDCDcTi685johuN2wC
xwGQb3t8M/IHTMsl6fsms/jsSONL628J8nggloeqWvwSarX43xYGTRLdbmoDmotUaRv+BuS4ylBi
cIE1e0ZZybUHFScz86r5cV4TYg5RXvIal3oT0zN2MNbCLoBgp0T8KBTcjgef+GKUPJP96Xbx2+vK
j6MZEWmkltVne8vG9PvON2bx5z/zmxnFn4V5LwJO/vpZJAT04ryNiNhY04VMgrPG1eHRRMLXp93a
ZFB6IfWOPkC/87TCh7YQbcEfusBb2AclQD/hhYzhORn8RB9iICvf3GAyNfJLcJQqg4DFiGirU8zE
Rs5yUTwwJ/CFQJgUl0Bt/z4vY8uzjjkd3G2jNCTt1WCyqAZkJInR2Ot6Eea+8kDAZOVidD53/Rs9
qYRFRl4qqsLtmMZtuNPr9uiY0ASwkNTkHwEXo7/Y+YXloQhYDQrC1pZFw6WA3/OUkC8NsnGjR4rA
o13PB8tAxUnCCEvwVmgJgrb2uCaOvdzQHbvd+EoymKBZj04laCrWS91gTzkcx9x/HU895DZDWfsH
T5zMOeX9lSNykwQO4ZQGCWNlWY/5i7yRW+WPsWMVnD5rv7DeKKSHBZrZkrnlN2iCuhPj1V/3imyZ
CKiA/s0LMJfTBJBr8v2MPYQe1n7HkCctfEIfWm9UQwS2x62D4F5ZaY5f8bdwbV7PxKqM/EGldhd8
Z8ZzkFZ/eDBoQeSUr9IMRB47s3TsP/+wKstoDFPHFmplfIPETgA6pbjo+Ef8Vw83g0jO8aeAa8Gs
3X3yucyuDmviIMe9KeUs76JzAx3Rlby7xmxNAjlXxBR4CFMilZ00fyZm8bdBJPsrsOs4nC8i3QSM
07cJf4/RWWILSUmb+ecQWwWOgoJS/YyCDL9+c+39j+QAG6H4YXzXBam7L9k0v1myiT/Xykwz67II
DHA9uyPM2nSXASipT0atJ7/0ytKSFMSz+ru/oTF4yKNNRud834C5D0WJ+Xo/4SW7WuAGjC5fXOkv
M2G0HzZAcbuBwfAJpcUHYs1Uz3Bpx7wU6OmY50VVPGHGNAUoVuu3pOD/sFqr2la5IcqQSqLKyoCw
t0/vvNmFVObuYkaL1A1HnlEdmPjoDbjWzM4mfD0bYtw86CufRlogQrWFC/RQKvef6U21OEEAQHcB
aAKCKM7+ihyXIwtvi5l2qxWeBkyh82H4p6ONuAYBwgcssEAprwkkB68+ME2xrjLOFngJoQ9FKCAc
SMoWB4cJuh1Hz1a8AlTwWa3y5EfXa3k7sj1KnTwuyOFaAoYH866whu5rDUwk4mf2lsxsbQOfU3Q0
mBRTyURGssh8Yj+bRLgHQ6353lImuGX4VDgn5mkQN7HEAwPs/FJZRNhim9yfux2s3pkHpoBnuxON
WesuEd6kB9ztaOxOIVo7DY/6Fex4zdoRFYD4M6Y/7a4r5nrwiufJ6CPI+p1tdvpZMYWo5D60MrIz
Ej9H43QH1iKcu5WcSJ7XhDge3giVqztqnkENKhij8kONTnjIac8eZzuD1CpLYHFkmX5yX2kMPWv1
NXy97LkjXNnUjDvE9+c4RuMZ+vl6OTDWHdsYwmx4liOaeGKH6Muv8HPnCxQ3bJZDbhsnBejbTW6T
TWceBoTf/qRk4/tgtN3yPuBND1llo9ZQvGrIUX5Wj3XgqmzDtVawpWgRs6SuCl1c7jtPpy5jaOef
pTBGCrlq+wkvVzW4xRHTaAaJ1HEz4uROO1vyN1vl1z6HaTpttp9W9xSspMp5JpF4kwstfFmKcn8n
FvyBaqk99McudilSFuVe47Nx8mw/mPstw2po+MoNEP9CA5L0T0zto/hGufdxR+DYWUe2YVHzGQoK
sq+8N1E7QEg7QI/lUIet6noiCHf7oNAhLTDzt2n32AKsQyJO+R17dhdkM5geKNHCQg3sZxmse+gZ
ilyOX9YQq7t5Ji2Gbc1kJkDkOtTVGJVrH0y04pZI4JEgW2Mgn334jJDcSllQ6h5pvC4IgsfGNVna
EN8fqnbmFNUfKo/DnzzG0GwZkGYS8/O8ckCvKV2wh3jQN5hRALzVlwkWPSz8QSRp9VEIqVZpYYUA
w3w6H8s+9RQoDf0jOS26oxlRUvL5/H02lk2o4qgbXEnQOvoFb8CCsrXqhH4dB2ddb9LfjiVcwyCU
HS4HF66C7W/bPi/GMNpLVTKogMEaUlwZSwnkkeYOvny1JUVmz1OXXGfsiGj9KeK19dwww1b0F34u
m22V916HA8KtLp0HEC4Ixi65FF9cbvwggtVQJKTc4Wr0Coh5i5y2ukspv3DtJdupZiRxMbKIhO77
5R0NAiKkmyioZ1YbP9ic2Fn4w4mzBGPErQkIbvvf3Z7a5Uv4cR1YZmUL3KWy5iNLnGJhyYkHcji/
BDhe4Os+kRoU6uisdfxN5DZ+JRT6R5AJm8S+dMwXtiAPVBZVrOXFLjHWn25Anub+JDUMHZNSloCl
upPrgXPnL0fpjatrgR5tDkvcgXMnpBD9GCKUQLTuWylxzjNUZdyeYMPVG4Df/gm5JM1T+I+hnjBd
3GP9rdgv9cYRrUgihs0h5GYLlk/FkDSbEeV90P726Klf87w/9Hh1YY4f/lVc72RoVfOs7GVutoYd
YWoBBBL1KF6AwNoFsCpbj0I1hyrmntf3r0I84eIYnZ4FOkh6s2o2PBPb8VLF9NPH7bXtRGHCVyJF
fX9+b3UtcNtZ1sHhiQOaFToUrFhRzJih8Mb8ix+VF1oMU4GM80+ej8EQJmXNYowtZ0lmKWNxYrC9
z56ZM739AZLvo1XjnZjkxZNdiXhBNU2mFjeruy/DQ4QDyg2w2J0zGb9t6kFdamehWUOhMPSt6BrI
DhndlWsmsunjIe2Psw4Q43xT36e0PPaHJOjVM5NKPELdrTc33veZdJIpKfRwcswNbmovTNNZC7s2
5yw/d1gI5laNoOl3U9uxqiOGFjyYINfhWGzw8ssKGNkOgUlk0ri71G1Rkzn/S1mU6toUoVl8XW6y
ZZK0rWaGWrIqEQiCH6eCjV4Dt0uTuHt+aIRlMrJgB/3MaRCxRieiAZtcX0tOVgTSikwTozvVQ5qU
4zQ+mtr3BNtk2udELLCpwGdd+UcYQ8HgLBkpwCJ3l7q30927wOFpxD8P6oZK1nt2T5GXZlap/KYK
3Lm1/ORu22I6rRZ6nBumg3zB0ahqMKpkbKNfzUdm4xce/UnEcZVIp50CclLWX9n4D+fd8E+PFfDS
m80AIAkh8ZCHg/4OReTb1CA6sR3/7w/JRmmA5pG51yEAVewgO9cBT4FVqjnY8vGVV3gExdCYUbr0
LfD97ylw89JUIQUu+Qqw7nUNAeZ5Db4Q+5iZsBNQ3S2UhD0vbkT34WpsLKpMx+iW8kzps21mOqhN
tLuqffPUBM13F3EnHnrUrXSKV9EpYWtI4fNYvO6m90F0WMsZTk4UlDrJ+0UFJQ0P7EX/x0ruZPys
kqPJAfe4C/NLDHwXsMKQJ5pvR+6Kw4hOvAK62jhKWvZxjUzt9jbBLLfl76Nh9L3CeEWQ51LZ5OBg
/YS62AhCS/yZwgzsPKaERcUr9BFrOUET1BCc9rfaOAOHeM6A1lt+8qlonov5BFgJhdFAK0LqeKSZ
WW2Tjbb3bE020QvBrLS7Jq5I3A5Ne/fM0zE2XAr1ftxtr7NS0SXwrZb0GpvOfPT/7ppLO/nskazM
SpkwoCUNjbFVms0UBzM4YJs4Pk+4y0CY4ncDXM2wO+TNemmyO7EBOY9hWzdxm4I2X6rt4uABBhRi
AdLrC2no7Ih7ms4t03b4EzP32QHXAA01PC8wSBc9endcVSsbdm8cR2kiRjQ0MoejqdV1sgHHK3V6
tHwVo1zccH03LCDdvPaqbFvzjrg1aYWAouHB7fGy6ZPHvgo3evn5pvDJWktZEM2MPBn25Z4FGewD
y90YUlRi3ahZinRKySLHF61PLmTOptr7R0he2P1KDA/YXUW9/eQ3rw+rnTXCP7JjcQpHVAn9WhMQ
llVflHonXhsW01cyNqqFEuitgY33WKKZCQuqumesqM2pq2b+HXEK7EsUVZ59bVpb36hf9ciqNkLS
RAQolnoBKoN9CS58lE5PjU1Q0WiNIh2BNg/LEIPjlWXdNVjTrKH0rFt6uu+raXGepIWx+Tp6oyce
5Ufy9F5tdLPIpH9ocTcF62aphODlF7G6vu4d4Xh3NZ4PSNFCbUTULuIrAy1HR8De8MS/IBy+9TKG
A8Oow3+y38l/cUAeipWZCmDE2D9d4crIu8luGwdSqjyhgXChPiajWGKZ2kh3RUQ16mtlcvYAheMl
63chYNMRp+NJKiDBhXtPSuTP8KUKKlyB0JaR8/MLbNDqB+Cq5JXqU8o7gSQO1u1aUqMfeLgS6Zx+
yKMrwDN915gHgL9LBqKPQVVI6o4Ixv3suXzhdpRfjmI9OQFBX0oJqdxCFbyITICLspqxZDycg1+T
+1y/xZ5itfMNpwN2wL90pRBSRnxCkIZF0pByVna41PPyeqxMIk5706hLOx9+X7IMBZIn5bAnErCj
UWQkiW+YmKKBJwPfnNyC2TxeZP4jltfGQGiu9LmSOi25VsUuOjfzMeeShxh9ibEvN5YA7ILgypgE
yHMC3pup+zOW6BUuPPbLyQ/axACiMCmzItKOme34nNfAGA5rag2X/k7FoOZum+DMj1xG3NmXbL2E
ZiO6mJhn5a1qhQALaLrMYSjX/TgXPDkAXg4RlClzgRRvuxc+307x9DA3+AtkZcHstBKRmXaEgXO3
M3aiRNoqcX8Hjx20/nrHyak9GnPL7jwvDjLOZiwGWKE8P6oRe87DB/zbS9ra8vYKhynTXBnOgcCS
A56lmOb7catK90/PtWkMMRkXETsQykvpPrAtdv3PvRrEhgfn9ij3qkye1KNYiagRFq3k3w1Atxzs
S5CYP2Q861Zt9NI5dvjYlE8pZNExuuEhchcE+T9S33QDseqWZuQtoKB42B7LcTAsg5/Q0BNYxH9S
CYq6n5r1BFnmkA04j3RtOoHx+E+eC31npxQ9k2qcyHiI91fW1oOQtqoyMtq2wXcZomY/gckM9mJ3
+mKjwySKkzTyF9/hlzKugJkNr7KgTHr8SuSuIcUuqbx2CLjRGDUaz8YJzRbsKB4w955KmliXhKft
FwyT3Eh2YHCutsdlE8cXKG4u0Lqei/tqTiOhHoHVFSaUQ49Yrm1pii51nx1I5686mSu7wdMIT6OH
KRUfGfVpXAraba3u9cSdvwdWbfHWqew7tKyfPP6fcbkPfMo2mIj4w1/SKH/hy5HCevECWU99YrC3
JEXby6hJMw8Ev537ZZKiZ5SP8LDa4Uvt3zP4YcTW912mKH/+zz3CEW5ZCAR7JqvE2YS6odBucBh0
IR1m5W/f+vteBH9ClaVZaNO8XKBCGvFt+BoBmFHjmzroG+FkeXofNrBHkWlUjFbgdLcYtaUxMiGX
KQrGP9yFf8dtrspbPeRGgJbOBrbIIULbs1kx+6l4Mx+22tWLYNImtK/0nFxVadH1xJyAbBUgBr9E
XUonHfj35yjTe2DYPk28H/EtdFvbJ66TO2VV7JdwXEUeK/TJDLWjHa2h1qosxjrhtwPg4i1JIe78
VHYv+qQ27lhhYwrpRAbEq9fFUxb8m2pPNjk7dODMcOruR69k71+MYeLAwMUoSuPmHJyNVnHpX3uT
8mSONinecyEipS/90HFmrgOnf7+/Qv9e33UAKoYDg+vfvabk7fozd4w89J14ugzbMnkqfrgyToO5
S/qf4nzglTO/E9Yu6AsmgTkgMSHhjtZhMu+DC4QVKqbEwD3y/Xt2dT4MlgJcZ7Wr7v7IUfTivj+t
JeYcjDmedli17Ou1AxS4/8RvKj69UpBeUaDl5S42krKqKEvZO93sXZP+XsjD5C0btvF1RRYryi/v
By+fOrOMLMiKQU2M7Yz74h/Fto50xKnCyfhJp/9K4A4G4Yhk+Ed2kC12HIitoBaXWrJ1aYuAabix
IZWHxfmhoCfTKs35gxyGCkI4zuhj02R7F6/0SxB2oPn5Bk60iQt/9kf2eYNKbrCGRGMF0oe8+BVf
MxqNCMZsgt420SngP+iUwrMn2twSQK+c7DK9DD/ohIlUXbGe2tZa/E0lLMBmZBPhybTxAnILtkZx
cvlelq0ggZaKuM4R3W1borb/wLVUIYXsBZ4qCq8ne8HOgWCem7VCxJ5suTWrrVtvIMf/MaNvrc1v
xqkFfuciQzEZ1QIBfoZC8SYOz/Sp+H5UGsRRC/z0S9AziI7QvaLYt7qlegL10Sqt5JYu4LuIhMLF
RsO70NdMwZ4+H6qBQd0GsXwUUpmPh9XRNkYGep2LQQWNC6Ald7tT8lzmUDRyqr50JUgVJGUhbQXu
rPU9iw1p52lZVVj9gFqYCyIVvgGsrl+pz3GhcsZH4mXFO3tftY574uWSoJ3PO2wKp6Vg449FGmo1
n/Yvcp9P+tIIu7A/86hZn3UjtfK3JzB2tahDsCRj7fTLyTlu3R2ISUbfdKzX1oTK1ZTNN2sZkecy
ghABEf4Ix1ejmLZQqy3xNzvLejhRq6tfkYgxPZ/neJF3OZKp5LT79TVxSHwMFtbYU8weY+IoGzsB
pv27ZLxaodY9pULVwAg5upMJjxDs06Xg7S3ckDcmMuLhJKDAZh5Q/+e0vfmBSp7FaSsXMMsXERrr
aqomnrB6ppOyz9TmUizCceEakvYcpt/JLDECGDlWqDloAuP8+3LQC9dioapw5EKEjL5FalXPDy1n
33HJIgjirdwXJtZ7TFz441t7dMU5IzHL1CM389XMrcV8LK1AIGpehN/HKHHi/jGKdsZJF/8bVawN
Am9V3mi+IiMv7+VfXZMiXC/Xx61QbzHwdKpvtE1XD+N8iGt5Az/pWOlbLT9X6hOyTLf4p4Z77B5m
hibjDFYsN7/r/bK6nvNzirc02xs3wzAr1dU/4Ul8ppZ8OBo2YJR3FmqfbPJS4HSzF0RLFKBsl10a
Gn1HC24BFFEaDMYONc5phgTCvvCHfuJmulM0oCRjLVfRL96pk3LWpRKxdqx9t9P6a1skHGveepza
UHYHOATJMeOpp1xX2L5KZjnUUJVfUBgKnxR5c81lck6hgjWx3aV1BcG7peHMdKf4txHWb0nT5G1Z
H8Yn8Z1EL9N9+HkvWp9XZf9U2iS1qejgZGvyiYJXP4HjAXTj1igM1t4i+XrzGInJpgK0rl1UBlxm
/sWALUIlKjhP3992/zJF9nEmyEzxv3jMo9hS0p7lPQmx7I4zR4whBiMyEOmcWDWm9Zk8FmSHrlyr
guou2+wlJUTFe6cuLMM/8bl+3T4ElmeDRcUVlSh/OLUbvqQ2rui+/G7C18tehdjmkX5ev8WxaQ79
QJuByhJytDQiZCJzv4FullLIjCmKrzru3CGghoqW+7VXIvxQ2qwd65lqASxGuis1bIFqpyIWDwVS
I7ohZmG1QJafeNgwJqFT4vZqu5G5Z8NI0o+HWPTifEt8hL0Vvxv5NR8DcugwE1i3ruQ0jcn/BSAO
0DMuibQhHZ0X2U3ikNT+KF6+kxDeEHGQXAosnMC0k/7nIpzKsOYbDmBr35YRKbUiQ2GTNDInvAu8
Aes/e+uDwuTXexL8RyDPtW7N9aIjjn7q6fdspBJ1kbKxlJ0BEG3dAXPQ5ZKGCzEfioCbTxvdK7Vj
L3FVqFORacO5z3zLvG+wKZGV/NXnBnXBwOUDFcHt7ZWlpmxmtARsFKfoty/iVpNPGIZ39W7mTwaV
KnEWd0Q7FW7nXnk6mCj7ztOXmQtDac36wA/OanKfP7NIbcGPTAuOXmoNfoCxx1tomx8IKXjMGBBV
p7dJR7PaN0xHtxm2l0fdThigUUHZwToruaC2Tgn0n7cLoW195cEKckkVfknlvxZ40MWjl3YonYC3
0wuSQJjA5qQ+RBRblUxz8nsKNun+BRRzHcgsNDGv5WaiJ8vsvukBk5KPGBCHt+mwn7V6vYvN3mJo
gS13QiYIk1bMDx+ecijUgUfs2mwTuIGBbLwrrcE37I3oMK8ME79w1QUoPyX6AGhDYx5/EdvITk0Y
brevfrlPJqZRb8IM3OHhiJZQZi1rtpvp02Atro5lc/0mqg+SjkTpLSBpOENAALkPkoM5Gm0c3WM1
YoSmgsqw9TIZ74DIYQX5duqnwUy4GANi2Asc7PNuIye4FyR9a0qBnppM22OI8aFLrhl0Ecl3nv3u
qFlfH4iIEDvfKSkrrCCywBRuwjHZxIQzAYOpaBlDu2xsNDcYKMsHDhCGbNYLKGIr4eIL+7+l4guM
/xGZcmP7CdZAE9zGqG6QUiYKWx1uWRS3pLldEwFydi9gfCAm1KE/3h3fSwF6+QCC5jHnzXCUS+o3
du+05Foh5fuw3kAnntVV4ebIYMtQcemTIpNg+tGw4mxn/PLQh2Xj9d8+YSeeGdvgJJhtCoeor8IS
ArinVWhcSdTAAX00g+4adiYTJqp7+Y3C4SVkd1J7A/CLFHMTauNFqwvPVX/w+cL2X3W/uozV0EmH
sEoG/ooALYvSk0QVwg5NRbKU81Ta/eg5NP5yRp3awu9cQveR5rC+UAUzODZhHP1LnGb6HlsV0fOC
4odo8nVXKwD3k7rXvdwwYqyDFCC4hQMkFMe5h/TljmFr7SwzsvNR/74Ejhj/gCuPeoaVH/AptMUW
2DC8XPc6axofi8jVh5W2DxiI+dS8cDD31trZ8hbViuuLZ0FaDt8Quh3UtIsXygupCP0xBGfoIsak
4GI0y/6N4Ve0NA1MI5Y2OHE7jaiKM7eGnyUD8e77H2lB5Z4jJPj1rUNpqiJEBlwHCEKSAJgzK4bm
JJIdXkQwIf88iO/831YMMWQtpE3+2+cLCsuGnzK7oVP4KVzJ3xuBRgELpnHGoK1Upg9fYgI6WHVU
6t36IXnoA7LNG1aRAboH4riHuFw8KojkG4ssN/Zd+5deSexQXs9sm/gi/v8qn46KMLkPmorJk22P
70mkKm2MSoobwMGDNY1txDrR+P8/vGjVNOV0ZyJXMe+8wsCL6tspc6PVBz8sN7j3JsOvwhdBfO17
L9oOhSH7jNTFm8BiXNv7/J5v6FCoE+sSFvBHE26IyysOnG04kyyYDZ0e6B4s+pq7AxgzrlTqD/1I
mdJeHI3fUV/vRnxSlXNZjAzg9b09EXi9rsfsTLae0oi2KhnaHsdPkxa132UBUw46SoxUrH6ez8O9
DU4AQ7Z3k0gvU/sFM7TJ6/BvPeLRoG+Lqgv42retLZmlPSMPSfw9joMWv6r9ijJuNcSMgDqPCA8m
3Wcy9Cur7ra/br78jLlqllEnS1aukZtctfaJJmVkuhPaifp8J3duPuh4QUNbUdug7uuo0yI3tT6I
kEHFj7mIov1tUdGboe031VpVJ7PPWHL415e8UCS8yJP4iH1WIqEgLK2QSFxTTDMyVhNQE3PFqLL/
KFJP7IqFSXzwZbm7UP6eKdMO84i2iUJpDP2bbm9IIPzoNLOH5xSLhxv7AdeCZ2MUbgamsFircrJz
wLsYFKrYmA1YC2wigWHygsqgpaTT7DLsZs1bnpMe9Lm0yFDQ2+2SA7IDB3inAVzxbPioCvDFvPGn
1yahkwaC1dNv4p0idzk38htuRHHzplG5W0yNUyxoatK7YJogBjw/zTwvvySk30la8rXtT/CKkerA
O9CzHvS742umCuJcc4WjKneIMqKbjR/3ZNxfleR5t/hl54p8y3oYS+SMRIWa6i7aiSSIM/MCxunG
AW3csYOCVAypjxW+OvHIoePiGnLa8kGcd+Ov3ql1RPevlUGVyhEZSAIvvH0dJTomXE+yf5SzYlUB
HShgqVDDJVLwCoKI3NN/3VHnEwdbzbG/cjALnCm1I/+JQncNqB7NqLw85FbSu6F6/bnKLHbMAcg9
aED3w4qgVafv6EpHjyii0Owmr2xTJi5FIxHlO3ynF4KSuRH6SRzRnBrBS6iSRYwMUW+7pW7jtLti
wwbZJWq5sfjN1KODm05NLp94Pyc/OQFiw415Y0SMXHjrP2z9KpPdg74Zm2kdRflnfbv9sqUqq/Pg
ZUSL2TvXzIHD/WHp65POVwkG85ZbX/TxLG99Ev78TjvV0meDow2ipo8EkP7WL6OMDiWZsoX3FMez
Z9YHsHJji8iuMkcIq3T6LSEru3xMi+JbaaGZEW4wZfGXGIjW3Xe0lEzaLaqHbUgXAUN2eXUhglI/
qDgC1718CzMLk6jCoNTjxWsEctF1ZcVN2kDP8GwXdXp1G/9T5r9rrs8Bev7aw7bwEBtwyT/xPWJ2
jAq4s1kVEetbUQMrFoUGqkrPIO0D+PH6PDvLMI9s72Xz/8BQ9vhLbsmonfSnqSfATGbZYoz9pcDW
BNGMOZk9NsNIhJuAT3PSIbE/PkKWgWX2FQfmzD0XiU2yE1DWJ5WGvTw4tibZpcU0e7WcXlBfhxm+
KEToP1zsnqtGuTF5vrBiJZXdfoUMFlPZEQ8ddSC+0cXJCi1cmKpxnj5OnN2zZwV1FRQWziL1MYzn
O5YJMtMSYN32Fds+9UY0AiKd/Re2eWvPQTbyqDblQ1Aonyhae1wFojj/nNUdcAQIOS5xVOWUZEOG
IXUNEdVlO3FePX0VFq88ZLbHubvo7cLRuOHDr4t5JwIvISa9SsEuZV1xuPY988Hqhr9YtLfZTl54
uoTnenqXihnz2uU8Ydd6pCnkgo0EkZ5x8rwmVX+9yppd30wVodW5oaScFueHiRGmjx8QqChPcaOt
ASUaUwIbnfmua8G/Y6uRji3pC8UoDtteZzaFHvtqdmcRgNXG11awQG1xPEnGtMMH7dEi1U3EB2zq
L0jVbakk27rRnkOKKFJ6VH/jqrcHwjIBnOU/BoItUysnRLv33WDCYXjHUxl/bUMHbvLwF/oUmHr5
f7ky/IU/TBrz5S5AAojrhgahqBdEn5YnSmlp+jDRpMP0E7n7EvKYT2eY5JoeSw3lnVdKbBCv1HHn
XiA/i1myF4Cs0YpIb0k39Iz7wPeIrAqHp00SEp3C4PM5Od2hdZj5tZ1jSm+udZvUbsFUG1OSCa3e
cRwB6WBhShuDwlTiHNMKOKxdKXisrpridJ8r28hWue9N6ctBiFvPLygOViW2wKEbsnQ6lBiWb2Dj
NU7AcBp2U7BPQ8N+NKADb4x/awNLrI4vV9bm9Ch2uqGIFJV4xXxMXkyJlAs/mNx+XsZu3D302CZZ
J2Nftcx/9XDMJQh/PWvCCqduL/N5KdkwBxD0EGW1O6zBfgJTtTQTssB1vvNW2JkZNpAtlgMbLEtQ
ORGDD0pCgZRPkqu2PRdc+fyo+W+0D4ZF8mhQE5rJGdad6jOiBBOGblyIO1hTVHKqOmFi+PPWSavK
ndWKxWaLSQ5cHugK3fQ8dUy0DYqmHdC3ShfWb53nsL/ytWCBIB5iKOczJJY36C2wS87uLf4sft/X
7EfQPRgrBo9jUyXbk5cDPe3Q7FGB9xbN3ZwFUJwmWrOtY9NXOX8k/qov8n00wzcslMdV6OFzKZab
Cm1lg5lRE8svUdv2opq5uad5XH0Np5BJksGRshADiuL51UjsPIfNCludCGfHf5588xNd41ip0go/
eoUqsK7LSaWz/RdJEuNwYubNxsaJj/sjQiVFBI2SKC5o8bYoaX3KyQY6oSUphrz5TwdXyjGcyB2t
/PpA+fRSuhS1y5mjY+KpyKEyzoPOAHsu4daxQInGAd99aJ1bReFdSSVuQjGguCPO+zuhpzpnQ0oG
cB9cnTB6r+IdZE/VZP4PdocIGfFEACtHpK9tuoUy72jESbR0FtUHssFtbyBeuQu1efQEhRKyFBFW
ug6xwMf3zAcW86FTaTQi8r6ipJKRF1KE5z66nkYF7W5soTIkjnJoVB8AuBvDngvI4P6VMfZG2VgA
rlAGoGby5X6fzmMu4u9B/sx010dDWf7FEB+ihOzcQ5uDzNg8SsNYz1ofGhk23R/42jEVNkUC6EKx
5pwiMjLXoCw3+BJmZP54U2DJezTeiIvkrurS8zwHOC1zdm84/ymQjW0s09zJ2DBvSaMDuWzUxwol
H5qI3yPBYU9nPaNHLfKVyMIyABXb7a6zoNGieYlwB2p0UYdtfn5UX9G/+vDlwL8L7n4d/zauDB34
A34uVA4D0Btevi28uwm9cMg2mDmtV9kSwn7KurjiDj6eh7wPuAJPv+ibiZLC3m/odsj7zD8s0bay
8R8SSpG0iD85EtrFzDLqxQUcsLOQFEdTWVCa8BlGztJDSvARbvrooBkdA9MDDHlkNeWL+Dyry9tX
S1iU3p0fDVDNd/6XW8TJLsYaVq9TI8ny2SwOZnCk22boLAAg9HCefEWGpxGFsKqWj1bGvUAnCXjR
MeLJJvOd6/MKwSWWURlK1S7kBSrIv3cbwcyQaXPpkptAH++aTJdYzbz6ZhGBUXVgERgM+oA7pXEP
B5y0Qnv1eQJfwC02ty4JwGNRgh35EdVV3yIcrNaVCCZVAx/PkYHrVr6n9a1D8hWD4q/+ghqhHr1y
GSHdj04YvoF51X65prKuRpste5uQryHAp8y4guNz4gUkq+YnDSWXynWlmCoOkP5w69VgYAsj1rgM
piSf1vIH05WZsEJxMn94BQBLFytGRHy4MedcVkMco+qwd1Em0+EfVhaEFYWKTT98fjnCdXbAHxjz
E+YsEgEvCENF92xkZr/p4aC/nczALORU5b2UD6xOmQ6XF2tXLuw1sORIjP1SqTnbX5qKDKHspY/W
RafK/rjATokxr27Q2ujRZ5tuedbi6BUFSWFrvSJfg484b60F9+J82c5FFC1UXNfMC0GeWrUmpQsj
yQXEYPd4b3V3WT2i+Sjtqr5UO07zWrRBSZTbgvOIZ4913nml1R71IhmdjUI9Spz/72H6HAzAUADa
+1Jit/ykNTPPCIXBp6A8o+NqeiP4b2rW+GKA8EbL3dz/vNJ4Rl0sTRUpaUCBHl5EuPaCjrnrERnO
WzZvkeNAyRaQtRRTu3mfGHXYXEV+U/oWsOBJDalRNYt3FakqkyO7Kf+BJMxCenRSSxUEple4bbLR
GYxa36lRhAj2AtgrKM50pw2iU3REryPy0lLK1hDDxSOxTtBHOzg9SjpuNDyw45sdaDUnX1MzemA7
VIUUK0jn2s3nk1oXt1Ni1x50kRt/H9Wc5BvaFfU6icgZyemmfaaiUBlssOEZlz1vclzPu1uh0SP1
H279wPBwNoViMoboCJdHg3Xm1njzFz2bjANqYG+3LFWdL0Jw/G+f9dReBURDOyLVMEuMNAJsr2Zd
j6+j2+4S6guvAmIRNAxHo8b5KQI1AHMuU1wpea/gOIIH4MMT0XcMoIcydMQ0udo57YC6/2YJYsbY
oG6HrL7c+OQrA5eBBRIHTvTdi4Zu52cz1vFc6aqm6YnQ+xxzqRr7iW704xTr3x5HwRROlQcWHzi0
AbKRBeEFVM1TFuX3nFG6K5lys5gyTqaRYUOAv1CUzPfkIv7yc0l6tabty5rXa2jnRdd/TpCvrKUc
QLM1AcGy6vNJfx21P4fwmeRsrnAoBbgc8/SDeH97gA7SvfmD5VFAufLVQnCFJC65QpD1/SWHVPZY
M8GOIg2Uri607w0zkcq1hKEExxt/HO3RyipygAuuB07x6YyBQCIQXf9SQuuUn54g7A6Aevem0ZYy
IDlptPNZdPHmHMmgXsFOuyh00e3kmLdrf9yLVVNqW7ZSBT9SiBDKlf3NQVYLqo7KmL+FE+b8k48z
V1yAqKP+WS2BJcI9WxB6Hpjc30r72CEe3oV15Sf7UqzhFkC2MDUSNqNZIchL4oHVIAyIax/kHaoM
UnsYIB3wl1voitgNHs6Wh5jbpwCEHfrd8lm963xKHiqQGYt7+CILhYEIY8VfNvxM0okQ3ylnE9m8
sTMzkZxzO3hHNzZsvQ58OVT6Md7QBOg5gHME5rahMo9jWvXJZJYjuj0vvfZOKo/uPLTVa78I8wUm
J/TVw0i///GJDlNVUDN8jzdtderpZ83mBvxWxMYUOmE8Gq3YyctutaHekX6lWNXIul/M+2K7Qkxo
EjyQGi5rLxxliTZ4zAJUQZRcA0NYH0yzBlEVb2wMx70+oOKa555BYsaEWjwt3PPrTKJkcTR62sHr
V07qciZXiRkgLOao5nHilX/PkCGN7BdqPhiLXYe1LBNSdy57pKyAup+VcIAH7gzk5R30js8MHiUt
U38NSQLeQ4Aeytle3XPk4YR0cE/6mjNORRnbs7kmt3H3hgY+SI2cuMqdIaQRsnZF9MxiFlEUZeZf
gxJOIzzjJX4/BEyYks+s4IKJvg370wX0qpNCTGp75AXqwDn+aDjsZisoHFYY4C4wsHakNLY7+uR7
B4+mhTeD6qeOoA5Mz32cEaukYpmdSgdolDyBmS4ALr/ztFpL+tFUP5tBZ3Nf1hy3wTc03Dc=
`protect end_protected

