

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Zt+Kvzwu2Ua/vrjhNueC6ZHFBDEZvqw7CYHtLwQCcRpSvR8qcFedNcWPERpPju3eJt3nf1a3JFkv
PrBPNZe2dg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BgYona2Iv/0k72I3J2JPeYuzuEtaXjhj+ZWCoU9nVssKXxrxRKdrDHt5tFvberHeN9tDv53k+E0+
zSJEc8s7HUTXqNlaEROAMDRbOb7ChasXXdVxfl3WOvXTlUGfsx+NSKJ4/HfkR4Zaiz3A3zH3MCLl
LSzFeWSNT1Mt1+XG8HU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FzDw40mQxR9kpm1uxLfUoItwH6249dxMvWlSzzE19zJKjsyLJvf8oLgoShFkGPrtSiP79qKNxcUe
hzH0hyrZBcM+hC6bI6Mi60dC4BhdqclOgz1qMMvUNpZqrzZ5JB+kSMGHVFW8GUXvnFCCxYuu5mP/
ywkJGUeSDVEZY2th7ObJJlKEA7icdJ5tzO8g4W6w2f+MHJPOeHFy+SupHzB+1djuSlirLlm4nhaI
hraNZ0zRKoeVe6z0EIEqhB9JNsFNiC91BziwCnpzBdkOsKtsrb3RxMWbRRWbmc0XLssKg5Ki5yKr
zZaZTZk48RIng0NJRYTCGlINVIuaWueM3WuBUQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gVm/uXv2qQX1H4bUmXuUswxUb0GUskWeA1MPfdTQVCi9Xt+VdX6mOhlgO6EFKXSas+dhLpimNzTK
aBHFEULIiJVFga1QEdJchUQ/rBMO2ShyfVm62wP8vvP25+deZ0Ac63uVlMRNhE68fori8KTc3x2X
Z6Nr7gpu2y0w16PhA7E=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UyIHMrvI7wZyM6hLJ4gE4jKiSWW2iEuHADz2BcA+kHWTu+vXmBlODWfGdNNdgy52INFMV1nxlqnJ
XDvv73yssq80S34n064XoTXJBVIQ+OApIu1S7Z1OlLjdyiOtUW3Rq9q1U3A+hwbuiZ1x4LA5dZoj
5xr1PfS7YeIFNi86pALVL/xngSOmrya7h0pb27Yqn1ZWp+ZFU4zxAnMBdh6smb7IVFLN7MVgfSOU
BFsRwVHyMW6sC4c5q5LyBHJsVE7Cty+4Vqow0WWDEITa8OtbnNcM2JZrP1+VHJVzH4AYNHP/h5/v
rWvTg/dH3ZrlceYDFRqzQnHfQLNZHJkGerETEw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 42448)
`protect data_block
Ge+dgH8gto3o9DPWq7bd4+6Lib3bvZLMcH0fAEguFjHJ6KbYBxSVMWoi3cKT1708z6bktpfit+qt
doziRyiE5bG4r6d20qKfAoQngO5lGr0UmCT0tFxhzalW5dQXbunXbkfgUwbYwH7inYe+sPAjBN8x
/tAAjpWcSwsIFrPJ8BN+pZHLWIUe84gifM2bROWplmgBecGFbirEOy32w+FMqwk3iLmgGu+se318
39pAgUAg/LkOH4Qsf8Mei0cvzBDVqEHGfwUTLcNbdnUwleod0Ue9nmyZOPDcralK8kwv3T7oLIbg
RiMgKctKhcfQ2jCgw3drx1amqT7KmIjA2RE2NWQB++O0Gz7uforJwKPqBD8NyQk6QcWLHS64jqzA
sDAZ0YVMSWIWOetAhi/htYMwwHjTJ0hGHAc31eEv2MyZuhMuF/dehv9KaDxdYXtX6Pzk3gpmAL1r
ZAbyM2yCUn7vIix9665yVLWYa2A+BvwpATsskLO4hKLnZfVzmoWZ057bepI0qOpWKkVrfMjJ5gub
U/C2iJ8+FTh9YoKT3kRwOwT8GpHCA7fJQ7dSIBsgUwskMZDn2uVAOFU9w1MocatdlIoVPHugqBDn
+e0qHTwPuR8DxWNWkon14Ror246fWcA9tir+UrM13C8tGrvP0TJWldvxQssUHHthXO/x0q82VN86
ap0n6T2um2eKgc5u2VTih8DD/Dbe76aH1aH5khvoeOuNfhU6uRHb42APbWTQNDZZwprLfiWD4IAj
/baPjtn83fqxBpt8D8xCHi8/gIz+AnjTo3kMOxhO7f4UaH+fjMJl65yoCel3ZgITgPQOlYNOwZiP
sZ6k0mDefT1jYxq3VP6mVEPjLqpXPo5zN/9cOiUa55Cq4tMcx2FuXUpuRzFkpfxwTt7JOb0+RfUu
isBhiDoHdNj8Iu52r54Z4vBNYWfW+Y+plIoGZhrg3IDcS9arqkFbijVi0t8RX92UatQkjbVAKjpM
vpOk1PIwwnesJt7/CHbW6i/5p13GA2qrmhpOE2nK2kroLXbexKJFMPXwB9faubBUZlHQ0q3sq4OU
fOoIdUX5UD1zjOvswlEkzqgD+0McuNDXMcyBZzO7HDdn2vaE7u0ObrmF/0fCtpXgDmSrJ7WSCV+Q
mA/kFy/mYbh9T6U7u4Igd8G7xWka50W0zFyskFSUo+5TEIpszUtQrdqdvyhh+pUSClMgzNpwTePc
pafr4eQ6QYOS5BO/rhJPJGphYu8OycWEKeSc4x9Qr336yEwngckRPyTSkNBM42uESUQLGchOLamO
lA30BSGhip3qVUWkq1aSrU2naQHWGDangxs1V+94qkjQge6pFtayLwHfvv0LwU9BqXDcJdYOVF8/
pI10miX6+qk4W4nqm8Owjgp1qH6T9Q5wpfv66OLGxoyXBabanSNfbma3PA34oHDKj+FVA2TX1kGn
ZnSIlQdoLRwHe4OwO7K1utRenku6zK1rKJthOaE+13YGnK0iWIP91juluLSwqc7GarnOtjD3ge7y
scL+wK7WaD5virxBgNsv6Sqfi8ySCDp/Uu7BAaJkLEjdrEKJQhCZPf6dEqSS3vnXJM+lCzAUPj/L
QldlqAhK5og54UG1eoDgRrdLOIygyC50sQMng9oUm0ArgV/CeQfgZjqW/LMJNVcbKNmkdYUgUqJ7
Y+m7rfnMhFYWykSA/EPrPfj6wp3rlIOs/aTJV5yWHtfE60CPgUXDnPxrSn+ZMtqG3xO0VL8H6jox
2+Q5FE809KK1bWSkrgzH8c8I3h4WG6YWtxPR3AIDH1cJE9ljQ5OGO8niuMA1vxvYTF7AF2a0u15b
6mRb8bGuRVug76zkGqZIs/1Id8JkEXArVkVHWAmfRd/DfdIsOqw62n2d3+2EZ2jAw3E9hLXP4ErW
rTlpTP4ijjr5mCj7bX1ykYNc2l9TCIUszMZHgRgMkhOKWc5PhJ3neMgllrfeqnCSJyXBCKVPjmqt
0VqlX7f65et5KKGhSF6h3aM9Yqj8CVwm49ECMOqagU79gBLl/e9nTPN2EC6lAfMYsTkHdzSTzXiQ
I4hbAgLpSerOQ+B+IKBqMXIE3Q2JKVV7anJBCWvAmblw5YzImh7C/6Xb6DDFGx+Inf1BdA+jdfqK
p7LqNA+szr0loXygup2dGCpePSwGCzoR5TZty14Ja+uJfQBUfDWgm+sDgXxCTdoqhTun5zjLJh23
4gI7gPrdAtfh3MaYQkNh2dK9ZUCdyGi51fL8zkNUdHnji5FQl7UwLMMzeWjVh85WoNH/kb3p66rj
qul4RQd+2dYUQwrOLo8/K0m7zLIQiCQozA//YYdvZm+tEgTjAKW+pLANx7xxfT66c4RH1+wRN+3p
mqd+LZFSgY0Y2gO/d6KTC+pU7Gk0hZmxoWNOIGNQKQW/Ddw46DDtRctp+MZeqWKynyQmXR1rdc2Q
s9b3Ie9tFlbV/5wuh1BqErH1hN3zCLkOXRJG8Q1Oatdak7s9WiEb5SUq5dw4ZE/SxJ+dKWQYKW6T
mCldnQkCWfcHG7Z5Q23b/5hXQy8JchSApxpPOq96aYIJQSUWN+kpkeQLw2bJk5LyO8lSiRf3QR4Y
chpAzALlNC8WfraUWWS3NudG+Y/gp6sYLdjeOHHAoXWpHYMzUSvSRZDi1+8jXkoW0B3z8VlYL0lX
1edcpwtECDPS6USlg+DNFBm2qAxTUhoXj4x+5cuGq7VNRXW4E0eSgnk/TVP/vdnRC0Snop4Rr6D4
1Z1c88n0Qy4hTJrg3OP9xO2aJlAIjrfoa7ZhIUp+NwzApTi+e0AjlMJOqQjeOzhmDYICa5fxVk+h
J9PJumVKnOg4OIv7Ms9E9Qij58TrEtI59ATOz/nNu3DYqJ6vf4J4M0DRm13dzd9x1nbQQ6dvBijs
B59VSi8xB+u+DwruIHZcD8lzyhmCszhHweXV3zque/E6eKR7zthvrDCmBDOPlKlsmyscaag++hPH
Am7Br25r7jlW47sCf0gw71+E26Sp6DGNwVgLyZ1YpbxjjNurjxCbyPoH61qGncbOAFo2WYhfsfVT
QKA2eEExtVElzSfj/SZUrKhE1EKrT+Cd/qs3IXWfAVOEgA5u818jUp7ACQpqrC8/5AvqHXTLsd93
C+L+ab2emriWzZUkKSX+SluPtibzT/CXgeNqxgBsLa5ecJ4/hb6tzzBK8HTbqDgb7wult3zHVgNr
ZV4eKMmI5lvJnG+ZtRYgmesVBJeDLzxn//LGdydkcjo+pq19oQjId4Aix1WjRvNFMmbBBSzIj3Zm
5S/LdbuDJT3Kq7xPz5/XkSK30mYSFawstxY1g4WF1Y+pyOrALSpJ2FxJ8bpWpkOcT7fv6lxlZJap
IujBUJnYPLdcDuTuAhmy/jw/Cn1iWEFjBNYO/M9NveWjl7XWB5uSjdsmL2/OvLMQH+yWB8xAst97
DcU2KSACEGNS72qgsHhj7x/ex4Xjg7e+L6FOSU0uweDZlUzuIBwkIQZ/UHrdm9hKeHdlW/5L4tlR
MisT6axLSo0xYX9b1nqJ6b3tMB9sD1+Kj6l5ojfpPkpgLPk6C4iNs3Tpc3AyRQylc07fUAcSY5Ur
Vq2qQ1ecn3s8ZWfpSIHFT8+Bg96bLvimap3ymWdG/xvNGjnaRXt2HClI5jo9wiK7v0Rakx9/7FsE
fMky+GavuxD+WAFk9FzyX5ViFX1s1xRYR+4Z+CKSNaD2Zd7JTHYOV4JIUgAg+2Pw922Ej7GJ+0ua
u3ZdY2IDVPYZFgFRTFW39YRYf0gPF406ufKXFpj7SkSuXMzTujmYN66krDCELvsEpWHzgqW0+Sib
WMoSjOhhNk3uXYisqBdn6qK6ItzseCAZwdKJss0gE+V80Z+3pA1SfC84Mp4SC0v08cTRpV3+k2tp
TLna/YtKJyf4tDbNEszo0syoDOvXW1Lh2sjs4wvEI9sYn319eWTBEtvHxssOWUd9Tnvn5RCT/30V
AKaTh/ABkluswIGSMliS6Sl/kKcd62HG0AK3CXwady7hDw0nftpmp0jHfUZgZrdz/9xhW2mWK8lM
drkjka/bb6wJAQ72B6Co8XlMtlU6hpvR2joSczKP77CcIVnDbFFwXUyj8bXydpOwV1h7yHKIXoxI
ENIqDkVMZwlnVezrXl7RxtZ+srjpVIRxdczMpv0fhxu5DTVy0M/LZyOi52hFVV9/YLJkvWdTfvNZ
OvFSHwCD//NJmzAcN/S13KuI+KmP21EHcr5UqBCu8lwypFAe6PLljuVkU1gQKeu3f7+blLQ3EvsM
kfdezRV3nrqKhF57DB57i0dYawnjn8RzN0zZYgOvXWw/ti2cWMXy/J+Nallt85uHuJZgvE+kGKeF
AyQwFZ7DLeot/+RK6pAf+WeI4bLU5LkcqiFN2rsc4NktBfg25iITCnn1ImlNMdkKp2pfmmeAcank
+fSdIhLNglOA+pkIzA76y/XTShZ77AT5saiNtGVOa46eU1yXxUWQx1mZpRiBM9P78cpxP8xiG8lZ
B1FjKKVa5eTnOtR2eL3dWGPcwD+Qh7DD1v7OIRJJvSArn4c6v6nmxVKkcAGXl/AU2Br5h5gOxUeI
IKX61siaxiyo9za8IE3JPHUTsmLUTkHwXP30r+pgM8WkR9+J5iSt+6ouIvXdT8QG9vZRwenJ20Rx
04rlMYUBL/Vq51V46aQPZDLMHaahxf3j4S0JSpJ6miWKrLMVtZ3VW2InRKBejmGUAB5rZrh0LCLB
Wqs6VZYmDPMy9lKRBMSX/uqjLXgG+1lqPrOeUFLh81WVSvoDwojPJ+MrJ52DVBqSuIp9E645GPG2
JElWYs2zvQkiYA5Di3kEdqJ/lbPEuDakaipWu26Fies3erMyZU8+EmW1YezQN6Zd2YLmeB3ev8Jg
HpKcNJKmBB4Y+qlnaDyoT+cG4LUTg9wvQVCZ0ye2Djw4esTBaVpUkLZqXcSg3wnGE/ZTLSAuJP7D
Jty7lBLVATdJQs85RCYoS4yCBVtpJIggD9Z+P8sskDELhhPSB/S0BGTl5gvLzcPbGv88VLvEmabI
KGwuFrnvIXZ4B4uD7CklEF73ucuWdok9PUf2yaLBLoBu0TLpmzSvC6f/AQkEMNSP8IY6PBzdBNjv
TK9cj2ycel8rL70IrcwpxemyItxOT20JiBsxgB9r+76YIgWJun5Un3uiBBa8wEPA4qfbITunD1L7
lJo72L4np+139jilZvQucnFnbOrPbKuTrWyUuCvq1lQmLojaIW7Den5at5uX8eIsB4kaQCxZE3+P
60Cg4Y2h/WMIysq7oh+DBOXDg+h1q18sBdQwFudhPOyNaynFwBicT8+aqPoNlAgCSuRNbZTcCpR6
zRlTH0dzCUQFItuwtux0smTA5TmbCk2ppitcG5zrlCHo7Kaa2xqkRBYCJC0rU90vBBnMGCvqUgVI
ipSCxXri8MRTPAzPxpPN4bnAAqK2+17VJ7zg+EJtK063fYwQnM22bMwqpGZC77UMPhQiSaW78tyq
hz//5rI31GhoQE6CnQEMUbbNz7nHBheskZhpYhoFPdsWdec7ElE49WSP8HzzCwUpTSWzKus3aVGp
ApvTDtj1mdLajeMB7SGyQGFjWYuoXlv3735asr1qBmwSiKXMK2hrbj7vuPgF+Qwd93Yr6lWqXRNR
VoCTIObwsWHWDrik76x2+iJz+xmqFKWl0+yDZdANFddFG4NNy4WpejbFDIG1dEQl2cp6fcL3kuQd
nQXuqVepjw0dm9tiDZ/FlZJhm0K3KXUsahm9TRRg8A0TncamF8joSzaWToOcSGDrkbov9eyoETQw
kWLp2sNYbBJkvLCkZqyEoOFcpfndyYYYT3ibMeHUdMUcTMkZp6xhUFZWqx7IiQwI3pJipW1hHf0d
6n0I1WMFPFLqejOFklfnR3N2BfZY+FpaCTqNTBeOTc1ELP49rHyIlzQxyVYZziKGqeqEoXpKpvXI
D/EV7JpRNVi7A8a7yTBfbyQHLKJhIDOk0f19mwwctw1b69sSNhYa1DPQBt9VWK3wIY6tonnKMArK
mJaftcFqF5znflwuY9ZKBAJNJq6U1idpFjXtmyol4sUYRcF/Nf5vlV9rzIxy/cnN2XHIPTyFGHl8
5paeR0WnF3en63lcYuCxfGs0Qnxg4OPgaCgz49huqj3T6nPLYQKcbcCRr9d75aY3hmd8+FBkiEkO
sZWw1NhZ/zyWZwp0sR4ZukPpzPc9ZbP3spwlGS9UkGhNEgbyENAOzUyP5S94QRfTJfjADaOn1UHC
u7jUG6ELMAZ0VQr7HjXV/jyVB3xwuB6Ey/yPUiK8Of7aLv8k5t3mOWsF0tIbWfbBK+ZmEehpCVc/
lhIZd4F6Dga9dd758GgjR7cNXyoQ4Dim2utbyA79xcYs5BABtBkpxaa3PrLLhcz4nTikX/G4qag4
65JVLPLokRXEHYRGhmdL1PdE1K88qmzaXeBHbK66/Z8zcHQ8Z+lvYIKMl7QgdsCRPDmQ/QGbTODR
aOQPr2Hvcb6t15toC0EM3DnoOdOieEtvzxSjgVCqMEZBMu2o043gVaJMc82jiYENHrtbSpB+/xU9
RP+Xsn+k3VMRdbXlyvLXnvKRMdgP7xSc9bIbDhl4lgjk0qaEvrbDqzPL1Cls7gPIZg+HihCaUajo
dm9JjQ01fskN1gOzCNj5mDPFJn1P+HLGuw+fiUgghlJGdKZRaJien8CfA5hnUBd+fpPqRfXJKgR7
b3JfUEWqVt4MkV/P8zjaHaYv2X96RM4QuChKCrR3jUpj3aVSwJJ1eHn0/g64ngwyuAHBO/S3JJz5
aKAZ9zNtVLLYogSqxS9MVZHKFGZrvtoY0w5OEa98fOQu95d6jgqG2UkeOoLRx+x2KMPkpp2bcJDw
hShD8DL0t8pGfu9DGMHToIcp6ziCqrHVr3nLotsxR83tC4gtKlVjcFJKt7iiRqooCLBwpINqigVb
4SHebuzSC75svYTgQss30ZbZvtTeTk+ctaUR2PUGEZ2CidzCzPzOIKi7recRUZvw9j+/PMvITSpW
1EQ/xlumkHz9bTj/tyip9cIyzyQ7wGILlSYnGMcrQxjrdFRk2DsD9tUZL/N2o3TARALwSqrLTlLV
WXNo+2uHvWZkAbWAjSOnOFIdYMIaJr3ipQZaXYSFuGlmbcMNeCjaCpM/2T2WoSsIXPtAJafZ6u/a
0ETS5drkFcfLoV25IP/VRzqoMbmYlgEQy7rRmxMQW+jpNSWMm3TbR6cRuvW5WdyG81ZsezhRYLK2
ATuFOzvSP+PXZ0arg96JSTrIHY/PcDDgm+B58GeFFS/40hZO2Shu7PELtJM33kKCEO3DhH2l7Byh
mRdXdy1fciZcXCBYaT5ikFBiQBqO54WTwDErIVcWx7/Il87sqTL5mmdkGQdNomV2Ga8YczDGnCTd
RwKlRjFbG+Tc4yh0gmLwCmKCODuH+1oYo/WJguEcloBPPjgXUNtQrGrjXSvTBG+Y5o0RSclI4M47
fbtrez2wJ6VNnDa91hjTj6dgP+4GPmLRyKyEJHL6dcXNp9b43PDMvUDq+VZQvW9JlT/Yy2iZpeQq
jMwJo2BgjpuqZb7PgLqSPNofYGghJStJywaYvpxYkaOc4IM9uksjQHEwadNq+cGZZOjRPb+Mzy7/
e5GcJhxiq9Mw5hwCizglGOs1OhGKPsOPUZZMUBicV5eRzsgaJe2sYNBDNxotURDHoVRDQ+eAEp09
MLKzp6hirfR7B9cw2V2U2FjVlvAkcfx8K4IOw61D+AKjNZm8JIZu3wP+DJBR+RBGppaZUiHulg2T
Jy0rumWjEY/kPvpv/uyx9e5dh3oSm3k4qawKHhT84fhsoOHIrrFUlt7h5tvI6WSrab3RhpUpn9Nd
E+u7Wx9s2k17UXrObdn1v4XXAAsrY+Iju7+DrCxUqMKvn9qHGYWMU6Ktbz8G5WxThymOsj+kZg7s
KninzQeelXZ77yNV2Qbrj8NHsunbLz+s0xzrviJ1KnSjCsXmjqoLKCssMI66e4b2hiwzYgBgxN3P
qQdspBJ9Jsy3wD96wLWa67EBv+PiZNKKZoZJofebS2vdwT8ZX/ur6d58Q0OYX+4buH/FHSwAg7QN
vS57HgGY41DTUHD43ae5KGIzxm2cWwhoWGLYZyzxiujRHvQKSDf8Dh8iwp4UaY1n7m4KbOitaGf7
5Gye39SH1IaYZx4GrEV6lDCiJRixdY31A6cPr33Afxy+Thq5iFssWbSgHF32Ah08R0mdcOMlfgPc
TVuw/os2bUGLBd3IUwBm0sG7WaPl1MN6yRssQjXG/8ZQyDSOWBt4hhxaoNVyAMBDDOZfAwSzPxgF
OcXH0DU8CX75uiSVTNROse0QCSSkhj6ppn74KS1Bp59riV02i0w8oCM4wRQf5wspy23MzJGQDX4e
LTUhPPwADtLm+VKf63UT7PAOlzRM9wximTO05R9L1dsCzP64lvSgtiiOPOVWg+QWObn7baz/A5NC
1hQs7I66uU6d8DH6HnvB4LLDffm1AlMpne3v3x4ogxcbW816+MJ36sjo/GfzM4+4TwMQjR8zXgLm
XD2+DZ6Q7HPpYfROHahhwJRCrAwHaLgk0nN2RbRJ/t5O8kUpMySwYdbMypVo604iDuZkj/J6YQ5F
Ip/nd2XONEZGGoyFiZKZq8s4t4VFh8jstBAvkd58elKf43KLDZln6oZuWIBXtqJjC95YcatlUdsa
In9lGu6vogtaDnsYqJjJmk3kuBxQ9nk3Xm37zEZfLpwa6YjUtrItT+f+LUbmLbfRJ4qy6B4GaqGW
mwZPp4kHatlCOMkcVmvR1iTS1FOGbEIrBnv92D7gEMKysxeR6NVLkaP5xwSbNUli2mpwSFoOENiU
LKwPekcC+ydczUChubSFqLGYU4fv/jQPWSjYYzojbHj2j2Pi4yAsNycoIL9GHh1XZkYOzLgr7jzq
lzVklhGWeCfPez6g9gSm185MliBDNov546JUWHX1O+7Vu1QBq/kGvU1Y0rWzERyNrVBtBEImGhu+
3l8ZoCrG/JBhyOWESzV2U3caP0Ko3UPEDRWzMA6qOGKahbcWdOsUWLmhixGFAqGpbqouK8JVMUuQ
MiUmvveoVA2RqMyuXlx7XGJCJSmiFUXrZBX3T9mZ4eyfIdxax7IRTPq3QDIKNvIHvwDeN9Ju+LkJ
S2KCPsSHBZQD/5r7z7sfwZh+OdGFqNUKVkOR89jabZypn7KljXGmEXRORAQWakZjndct0BxT7Vf6
4rzsx/0kjcf0YK6bbiCxLn/tRw4ptvOQ1x0BdMeCvp8m0SrQrMtJRO4bP+wtwSRQf5Ymal9K+SMb
w4+sT7GljSrLNn3vOS3L9eg60kXPXAktvt0RpNdV+hOF2pZEUKiCHdXcm4TkPQyf4l4bRymQ7H81
jFk8UkAqD0KtincnBJXcFgnjJMFJRi2f7LlWeqiYYxmiHcZ8pQ9X78sLZ9IRrvz/IsJaEY7xVSrS
F6zopAnOQQEGuXv4l9JshrVKS38e+wbWUVEOKyBt1KsaPypdmqCH5iE2wvu4oYSOWBHNwubkDJXk
z3LvP0MXSFPL2NN6E6IneOTbLgyXdNbehAkMfR9e090pcDteCZx1nM82I4BEysHl2qCfdIaUWVP3
K8IREMA2tpfAF+3iH2T+cECamLJtPaKWRczDTdSgVF2ygeTtjejythaB2Mf0VlscGPUSLEKoHgz0
Kz1LE59+WnXhXWlS+MRDnVXg4iDqczztukvq0wh+As6SKEk4PFUG9ed1blIURNf9HGTNh4QYwx22
md41Ox7XRt+vE0Q4BZ3CL8YwggCs5vM0n7GRTk3v+Z5uJYcNOYZmqZU+bkTU+EnuipHaw7MHRGqu
NwirdIgm97+RTc/xOEAElhTJzSQHhpwcrfi3zIuAB4G6b0euPRj+WLGfXxsYulvB91H3Kqd2ZmwK
eMg+xY+TUayVvvjplRvCa2S05x0C7wlG9MXxXXclgbDDMkghspURFfTRN2xtMyACgw+AiGnsZIZN
MeG4N/rJ78eMopBXmHEoLXlisijh3SPoY8ZS23UsGd6FE5zZU5Yki18kDxZR4k+/Iad0pxXVxSXg
4/ktlyFviXIdstYWCsCnbjwRBsUzXLJDZJCzDkcOeXQpPCqGVRpb48Uf2WhetY0jPHfiyhIqk6U+
cIntF+Ii1PbR+LLAt4ugqLTzdKWHvQuv4adE5fz0rCO70Zw0TepH9eiCy6FIMb98JVv2KaBVa8bV
+2hIbMJCWGT9QACH6MM9IHGixvj+hb3hfkSsAsgEBlGI0cf27dAdUegeYnRI/rgrv/QZPzf6FkeJ
TkpgMvb3sGLTtPqJkNNAuoJfUAtaZ2t2/jigTYg+XU/3RbPW8hsfOOyn16wI7LL8T0Bs6gq+hiu3
CE+VfeHama7/BVfd9IL0Mj6zejfVaol46cJRu2xxpQzbGAYg3FvddJw7EIwOg4xrsdiy5638EApJ
YzwQwM88QGRiKG//ruD7bU96/D4YsjmW53lrJUoPDCIth5pGsHYzJth23jx4qXEl+dJIaIZWvAu5
H8L7uhXkE/0pvZR2h3YCA/CyjwN7BiEOqA3l20R8jSiVisC5dF6W56H0Fi7Q9Y+hYjnKiQQpqRnM
88c/mPi88+P2PBJVU62DD4pvaXEsT1pvfjJAa71UtisrpZWjRSluhocupLHhIE1001aVgyzFX4+1
pR1VYsXszPGYMxOQByoRrEYY06qz0vysy4czqEK47BBYZOe9BFgBLZONQAJ/k1DLKHtbqP8UVz4U
VQTBgVW3exXPpsKSpetlRimMUYb8aObMM18XKsyg/bAwa7htT7xfsO/WWAKnukQnUzO81HgEaEd5
UBGjfAC8HgnlaXuEWTmdGWrN6BXhnT39QHzr8VdP+m06hkSy5IW6LDAcz9CSjwqU//1ktzrFwb1C
AxuXF9PSizZLuRnQtLjdib0P1m4Yan/M/ZL2bEuQ7r4QJZNiGcAhV/hC9d2+ngQ3PXXetfBqGixy
oPnuui3kLyqFWnC+fx3UxzjEN8CjaSxvMCwfEePGQVYfGp6nxSwsDQfWXtCqRz1+k59/lET0FbBv
mTMDK7ss0ehpWksX3xjqKVPhU4M5Qz4FvTymHI2tkElA909MX7lhVm5e/vSAp0fCFi0NiNTHn9I0
wPwu3fXvH1aua7UAeZONzWXKnetAV3+DPZsEWreqIPvH1O+G0FDbRaSrgpBLwZFYQaLcWCx2iMld
b9JxZs5vRTXOSG9hgb/rfSkdUhtlgUvIr6qcKHfr1oYn4/iKLAdeAKg3CMdxITSiDt2fDnTmy/l1
ID6A1PVdiVA+VxnrFYEvGrwaHHKIvBuOmZkXzc8yfsB+9FbF96Srtst+umeiWGlwl45GfrrpsZsN
/W5rzrjM0N6A1JMig+tjxLwAiNq1/pE7aXvE7VMNgAFgnhjGrTBs3UC7i8K9TKua32vqk50awP/j
0qtLBSJLunO6+aHFFxMJlcoM6Mk4ZxnW5IQu2If8seB2YMoQCyCNUh5VmMam2kW6LBlUI+scsgwo
1IbRcPh3qWJaJtoyRCqQixq0h4jdNFIbuJ/nfsqRz0DOedL2rfdm/zts0621wjhqpBhFvHuJyZh0
sN5P8EeBMhwm0YNh51PIDUrLoc7zqCTu7su1wHEI2mTharuFPo1BgJ40nAGgcXgDBiliHoEB2Chv
8g2iW7rw46D5ir2PS5oP7r1HTZcjkp7iB1qNLbF/p6EfVp3VaAxUVO0VEuGccWeSgu67k6BjX9YM
DVgmwgmsnEyhwivsokWboVZm6T3BGx5fa6zYGd9uncmSk6pu4g+YqGOeVMaD+/gA+Nyus7zFUFTX
9xuugNPfMEN9+KkK7C51s1eSAKTccM3bRnQaZJttyKiqdHKUy5K5uiHkmGK/CP+oehkLyrKi/PPr
GfxJHg0gASngbOhDH78/4DkZF2B7876zZ2WGOTBnuj/AAjmFrx/09YSFIzGFxGZj2WQMDNXobfoQ
Ze4MKfCNS+ZGsWdQlceIW+WUkA/gsjFyVUKVjtdGFH4DUpPSWnuAMHDblvt5GQZnkZT5Owp+7Zq+
0VfyO0b5bH5p1Ycubz3x67bPAdhvczEH5Tl4kcNFf9YLtdxRpLRMRIYnjS+5/Ea6dFewG8kruL/e
43PltLtXK2EUfn4tmUBbYwd5eLNoesf+ykDGw2bQEMmmV6uCVeUGhbt2WVKKhT3MMudDOvTvW8Qe
yTw8LbUVeXE0KFuYs4Kh0HTAKcXpsp1q9G74ebD2tV3ZdgGLlmH4sDKraHHh9XUeBejnXspEjjI0
0qo0MkjDe1xHIfVntjj3+vXO9AV9iGselRH/UA0eYLNhn81+wIFBarSggk2hGqK0bCJr09nf9ZxM
IpFTjEjiq6Jmo/0NgCKnLWAtanDwEt2BEoep+01yDzGZTpR9b2snr6fZOY8MFGEsiHdTPUGu5O/q
i76EAv9OBtGU4wYcU8S8w+W+S5g5s0fcigzOiPpTyfSVQ+fXPRTkJ+ZpkDPAVAigqoiRMNTd5wO3
/iLjcDwMw//WTyj02c+YghdczWiogXXjnuek2+pHE8zNYM6rETfWJd3CGd0g05c+UzYRVx3VR3TI
QP9MMS5FKQqZw2AKVK62SXop+wWpmGO7zrK1/8DGj1PqjcJ7vR3NaSBTrcMNgTOT61yAqUI/RBB0
i9gZlGnnxpevaEGZ91ReSRnWVqdkja8Idl2FScGcvCbWysfkAWNzKr5YnVY1TnvwvlR6rRUz2abR
xExqQfLfGcj+NE7mA3dobrhh/0XbYAAIX3noZllbqkP153ta3un2f1w96VuFMkK+9OtwCW7Mtd1B
cYkWSzZV9wnMF4wtQjhBnXYGxmzXhaC1QVJNFTP3+ykZiIrKqKocRV/QsQJWzyVqfN+jDyaYkJMH
pT9MuJ9np5onDZDb6azMnvsJnSlsWcBnUAX/yclFkzxkP5WPlmq9ZVuWVAORRo3QJdP+Wsvzq6xE
qxJhoDXyjeoroZU1ik/lDSL7qq5k1J/3ZpaNy+xXsXRLqS0UCQoouxE4waW8RtG1/qSV80Ob90Vd
5ac96Uu+4lcAVoQyldOUyjunCqbBo+ph/Pn7s3h5u3Xu1eVGEfNZaHyyMBNZZZHmi0kFjNqQtwBk
LFPQZrbwhi4PshmtJ0c71jmrNnlpT9ix4EKIxrvSndDwPnLd9rGcQQ8br97psBv3i5kvibVOvL7n
tYhQx1Hm7R08l4HjqtUWu68e9F7ymi9/yXC1Uz29TXKcI1ceX+J76zdPxZt1RUQSrILLU9hV60xh
YMjQaqx9tII8Jnzx14LU22XR2pkytGrhqpyd50+xZlOItGrIXKDsl4lvuDO8IdzxL/rUj8OXJIGH
feXPWb04XkCyVXfggYATqFjlDSVlAQn48zGhTnKw5bzfuJBOcwTPLmHYjEzbajXJy54jqjRGhNId
cexYm4Bp9fhBNj3s71PD3VX3/sllmpfVGQVv14a78Y5i3lbmUfb0DgG2amL7fYwL9kJUfwy+gVjZ
8TgFDVZopt+R9Lb7kg/Odeh5OAvfoXxFZGZZMHgshghbOuH74n5VuIBCpMM2LMPpP0kUILw91wDz
vbgdsgkMA+tJ0AzdFOMv7Y5/3u6fOvmNOw91bkQZkBsJwsVdJopIwZawzeHMbKhGvDiJv016MuPx
2FVVDdZwxZLnjcC1wLwI19RJc4mcg2u7gQn6acHH6TD6GW/cP7WFJl6aKJd+3onBUcfxSOHYMqVn
NI9zX0G5U1YGBjvS3bxba6NFHtUVi7mWS4/jAIdGuuyPlzBGCx/XkMKmgM5DqKdSXnmdLOiF6bET
vAMbTpsT9YqljlynL++sc4yxZAvyWm/jmnguuFbGvbkWa0/SyQrht5/+Ji0Y86rhLVC+s5Lx304r
vhFKd5viSpuRru4l8Iy5z5qgO5OSYUNI2dhm6yzQXOHaRwkUN7REBBoYtA5g/K2/HzrihXvcuy61
h81y8JE9dUhfrTVDcXcB7rbnkY7wh0SoMJZYcUsGtDG56qZuTipF8JS4CeXrYJ+Eev86KXmjd5VU
KrHPnyunXBLcc2YfXs6bFqBnvrNu8NUDQhpoHvMfw9+iVZqtACK96FjV48+3BGFZdMepO/zi2R2l
XmHCxs1AZv1U2Au+U5CHWLJLlZAOHaPg4bdVSpvsa79rv4CWIB9mdNRSecr2aXdjfc4p9JXH7V5B
vdqun835UFj7pLKc39vOoHi6lhZcpcszCPL3Pg2aY4/YuTssdPB0CIO13VVeSDKeJoo+T5oWU8hG
lRJJ/RYzcT+CGfjcX7FSnYWK6RLUShud1O1XPweLvG0zHO892DEDy2eqJAPfF0CY0yd9kt5LX1AE
Ad7hScPDGE6wcJGV45OYVdXqubHpoVzXvyKH7qYZ3+r+V4iywByFyv5Cfy1PImnTO5yxImNJJnPc
ezWhhRaSvAxjXSO4BdVfsq0mMe2wXDbWIR7mCZxu+YlmUSCrvlOxn2R0+/IpB2jkKEPAOyl36R9z
N9P6h/3HGbgvpgQfbs84c3jA1yzyzkbdZouKqeSiMiHiB2Yda2BaFqzDGLLLLQ5ppDyCHQj7yTZv
G3N4J35Wl1oo+EUpzBeYUHlkSWAC5OYkybsf5ievUk3dXu9/sHTOP9Bwk8kdBeiO2Pcw0eSnNo1a
8/J1Q3FASL0a0LqK2YsMkEppUwa97BU7LANKImsFzymUoEnmZByzqthapaFrGM3nt4dBH6Zv5cCa
iteNqIbo5dktZH+QyO+fZtZDdzjFJfVqEzag1d529YVHCWMjgsZ6WxtZLbI2uPZAVzdbouFmotWL
/pSl82onQ9FR/OycJ7XaBhcsdXf/r9NgHDx9T3PMCYgBTeTuYDdyP2IOc3zfj7S/d3yPZUjOfNVu
yqpXt9aHO65qmWUp8rmAt9+/3pN7P7Ooo9TMNJo9ZsYWAUaCQzGS4csM4YK1n0twt/NwXvPCxp9s
H3Gl22sh6vJmEksQM3Wc8vI+FCZmuePD8wmPnze+1hJwClwTvMeGU/+/ADHpqUG9PWUmFQOP3cjR
tsEu3kBDEc1+DSeG6ZYnjJNF6FK6Y93PzUq3Oa1YNE6tKGk3qbpX2XL6HD17B7Atkh9aSdLmm1jU
9281NqdEyBTZW4VgjDE1ndAWleMACHEGGW5mc8qcvrFofKDjCBeVBasqDild92xftaN8KcFqZkb6
yH6xG2RUsCZJYNhzFWn8zvhsdBRtmL0bBz5QAedn/J0UKKaZSmnLkhbGHl68zn4vG1MmCeQCUCyy
jiSy+icXdkNljpiCtaaxjuSYqXnSd0o5ctFfK6EDMTzsooE7WAVwnZmYefnrRJr84xbcRYjrKfHX
baUqbtisPWUmjqDZ0XHG83lKfcQPnbOjKGLd20LLIEhvsZHYDCyUfA5Osyf1QFxScnSHnus1w/SW
6ve3nwBGRqNH9oOF/lM51zPN78u27gEP1/v0BzyTYtFP+r8ufcAGQBGnuP9uU64V+okk1kYSppTL
SM8UBveDCsVcGuZYdDLIciWk44oyz4ziZfv6+QOYps53+QM5Glftn9DYeaTsqxylzr+Mxa0lZnr2
4X5xQj5XHbenbt2Csp11uK2JQOqLqpbm46oEcBK/tXq3Ay8d61d969XG+pzMBwWH+k1Qa2qBRb3y
cF9WRvnnyMqBi7uG7jRYQHDbIADwPOnUGCHKVIabiCZbzwGdGVOd956E0twbFkgmRUdAkaGbb7oP
TglHt20eyCNtfFDkCDxtD1Fm5O0x7qYA8Y+ve+gNv86FPNAEWW/EnJiS49jKChBuLqfDk5r10Xpg
ToAftFjE5TzzOdxYZDg1OwKzscAW76Ti0qmhm87eIeUWBERsBu/pFGLGa6c/ZMJjVjhdI3GJqjrs
+WbhOrS7uTMB3GIWDisD6Kw8FaMjZQ2oLdR/X9f1KHNLK/VeG8FWYjs9K8d9Y2rldUtPPynFtMXj
QgucC8614/Jcp5axCfTVkotvlycfp/ieTSZIFES+wHbhJvFucVn6h8CkSja62XoDzubRG4y7516u
v7SSmDaV/DrdHc8LNilefKPjdjiw5V3dc5MqZqeL8M2rd1hMGR4t3kqwcKUb7hIbTRfDfUg8fchv
8PAq31TMkoX6Vp7ehj87/2WYxGLCSjjqRaoP5vIuGKtFVi8d6QzWEaTtwoOaZ8CdRMY2HpF5MQ+J
YTnwk3dyOb0gia+JWEyXfuFF9fV/0JZ3SIiAzcQZaf9ZsFvHOP+GsW7QysfX5wzHFxE/S+IypNtd
7R2+BQbyZ1R+C/CXf1ateIhk7gT58+GmcizEDkiI7KGZbj2nQv9IIs8UO3PNfJYLQ+1z7LMGdJ21
lJG5lhzN4V0s2cCbX0fNKFXoF0z8FIphHPZw0LpU4pHlphNw0dFGBpVA9DEIJtH5uexVMWlhkH/s
YE6NFHpjVyx6G7b4ww1MGOVosmWR09dHk/vMGJBAlznUL0zN8bBWfJRQqTfS7Yhwke99PpmaDcQ6
YwVlfba4nFH1MW/iOL+WXtGNtpMcykwQWMmSRnGBkYIinExiULW05AaiXkAOGcDQnhg4aygLcIS0
PpObzy8eY2R6fESakmdqrFOd3O5hUSoRjsii6Zv0ulXc01T1ySzNdpft4xHWguYeEqN40dtJAkb0
Bso7XwUM616Dk8F2/GawvthNRGS+vtnuIjmGLKwAKpPYVAzuPy6d2+If17I4Nv5DPcyoVmvnm5KT
sv/f5V3uNxTxDoKslepv2XNTGRBBpyeIA/bjchYzIAhD+xKlVAqD9monrfmE8lPS52Useqy+RBU1
o4ZkUQjh2zX/BHUzjVpWjzZLYq/DEJZFFBdSVC22n6d51Z0qZHg93HfAJvM1ktYtU2Rliq9DlQdL
RWBdPMpF7Fx0ykbQeEGQhFO+NX0tU+K5E/9kvKPhxgSCqBfd8EQoP/5huPy6sXCEkW7ZT5R+4re4
IhcL/z25NBCf3I1r7E2c1s31ZX9t/9y4BNKdXEjXiwQu58FDHeUA04J8O0OmbYw/OmDM2fU21/z+
OkX/1BvfnWCsTsCLrh1HRaihdwF44GLlPPxv6JjVzX4+FUJnYOHZXSDcjoLQRmwyddWSn81Bc2rw
e7IuF2pKB2s6iz/zLLkbw8a+vZAniQhrayD/9LH4leJA/igsD4DeIm8oFh3vNvdRCLoY0lDvpJlA
Z7tWJd/M4C+qRCbfkNvjBwNhbUWSxXRhGdH4Q4R8Tdeqwxnc+s9/4jnyJ3P0ALE/zi9Jw6UXuClS
ojTwZtIlQ18VtlYRioJgiLgnbODBwX62Fo/6cx9Zz/Cr/cKYaVNMbQtARSCKmYdcOMO8A2PBRbDO
mjM1pD2+rgSboQfGPSmFJ1dy8SuiUejN91p2OoFeQ3gRS6vHvYLX9Rhs2odjQhbNaLuvK46XhXJO
Q3yqanKf3hl2WWDMr1It00pXeu0hCdFW5zEJ8bQyMSRyyXn7Ka7YD7QFMbOCvpqY+2Sc502RKZt2
5QXXzMtGdbJuwqVGyGs0RAxNDMp3wKLgDYGyysjJVIkojEIb0Z07u4zkebhJyXUdHeKtC+lDHMr2
dHI2Mbnk1jF4X+cjIG5IGp0cqTD0wpwgeX/Zgb2clRb+NMKVshUcXZZZJjph7SVNUfw+H1n9nF44
/EKIenoAluIscx3hNCjXN1sqpBK0gROUqk1PIM6qDuQ/hr1I2NJk8vDbaaQVMJi0TqR5l05fOXBe
ZcNsVn4NizP+Cd8SY38v3S4So0x13bk97UfSQkA9KtdYcZS4bfx1HzQzQ3haAcyqBFaueenD5JyY
LU2bhYY81WzjONmf2cXZ5nvx+uR8DfJhBiaPRd/HBEFAbaT118CyU0dMI0vzZXSQPtgxwxxUc3ou
slJ7M0DshuBK6sI48oXYAJItZOPjBQMlH9YokJkn/Jbu6d/+jA45DzThTLxedl6o+nDuT4IBKIaI
q32j/o6lTpfrkQnmZSDd680fCxVUqSDrt3W8hArmfGpizd6RxUTVXgQ5HiE8oYQkk6qp45IcZlgB
25S6huGHU+QRtAy2WicqEISy+bZJZvr21ywrzulmuxS9peweiVGU8i5knyHKKndGaAc+0qYsl69D
IQl3hJsYfzPzqeH5yLJn/ttXWfP5TRSjaTdRc/OqhY5SRLUp8LQgKTCd0KbykXJS69TNtqSEGfYq
ZhXfFcAIn84+gDuQjCfMBvxiHCiei3tSFomTyKmQAxSsZifvy/riXF3PcxTZoWPN7V5VfimToeF7
f6gLA+5PEyn/AxC23JRmD01e+6YRC8Qn9Xi7xpPRerkdFKRipFbW2ZQ3OuhbVJWjtHgsmtwyZROf
CMdD62+fgrs2uMC+kuy6l/LTEth+3qxUm6XajHuDzvjCsc1bAi2Dmo/DzXfmvjesY9jnavb3wrQY
y6o60fLqQk/6x/za2eFk82cbbaiyBfCC8wq9uOTVoWXOo5WSs6iNlLsPeEI1cLwIV31T+5AMV+xV
6KDnnbxIYF++KUdeDJCQtF4ln/IPA9nJxqXRh1kZJFxrz9X2cn47p5OF0gEtPHq/qLv0brUeAf8c
HLicHSxZnjVrFNcFOZeVi5nYUos7SF80J54a4O+61UbSQTSFDwLRMZRZJc142tzCy55L+PrR/JjF
dg1uQLJd6cQ82WxX9PMZfA9OmI2xU+LIdYqAO1aFxf8UpVTXQRvh++TljYnE6KDMlMc+UkRMCfmP
D+GTE30CKw+CbcJ48H5qtYNyqZcAESX0RQ6wuy+LfojETuhZOXOynf17X6xmGSpg2drEFtPInuh4
/1LRcv94h/GVCunaTXZ2epZN3PhoYbjgI4sjtLTzgyt2ESqoyMPxogKptQmyHIIB4CSpnV0M2bdv
JyRDnBD9XDnYhCwl4WUVnBC6xntW2/XgqUu5+uxc0l8wIrp+3AovVC2V6YA8hilXLjotcBU3lZiJ
dkDhcfdLWZg5U6tChCVFfGupUigGsJqqT7JADIs9aOmIMkKNVn58PtYms2r4vqF2iO8FfOheSmqL
hlzXbAAo6odcYFHnBC6kXh08hxgaIvCn1by/M4HOM5APY/QnTQNB7sdayWy2+svA9E7JsCdntitV
OZVQhIoPx3hhOfBPf2SVKoa943PGCn1IFoa/djRF9E85+LxJ1vEwv2DbUCLLqMqUgDtRkjnrvS63
NMlNa6sj4vds3f1d4dkukTIs0aoVG5f0f8eUKaVS0MmJCfomkCe/iXu3fd0LnIAF1MmiazUiBMiW
mQuVIPNHILONWVXs2YrcO43XURL5Qs/hnao4nfy2y656mJ0e6tARXO3xsC8ihV7INoDwuzXUEk1p
Jw1t+DxeJbS99TA/Uf6yf/mC7GJLaal0VZmbah0wn9I/XWkXJ1ulkgKvrtIy0v5ajC+2vzWb2eiO
DMAoyZ+7vRqJI/MNh5UnsLixZFy7xXlCM/fGZDEMW8vz7W9KertiXc25/2nexfoNEgQ+7zZvZ6Zw
jDgGacKPextrJYvIzS+q862CQYZ+dbtXOh3epv40U+UlC+9UM5l+DSTTap1FCD9By8jOB/H2dtTl
LYFrgEAtPmxc0BuflO06LrL/XlYbkP1sqqE2nhthCKKuz3MpR4G0GUzSAp/mG91Sf3ryIpEh3v7r
XLjpzF5Hh2rGfPJpkyopR3O/jiELpA7S5Za0J1gGiuGczPsAiAbZ+4V76rN1S3Bk2Pbina+rmtru
tTxYiPcM8I0bMCDxUB4N4nAYfBGCzAMo7JjYih8XJxOnustjTwxuwdgWgVeNrlULc8uygX0XOPKr
7iSwq8Xm/4jmd01E8IU84tc6MdZpDmX+Si5nzOdET/vf+EwvG2JGM3lSWZGtGc9Z9Ais38zuB7Ig
863BloDWIiZcjCyCQg4PytJw1zYecSdcg+SfCmz/wmYPpK+8hMm2tj1bsom+cTLclAB6zx1czu+j
AZ++qIkWyRfZgsR/Q9TNr08SFQo2aXmUSX3ofZBYYrHefJyMPPHbyviCKnVb/EIVjgQv3+awrCpz
tVL8S4GhrpMOurcnQiuZ17t3Pu1lpMFytxmuoxUYZLeur71blhW8T7j0JmOAOCjHUegBccpJmUzA
LerHUT2NjFumegdNmzBlCFlDZ7lyV4QHzxhLCUiQ/7ZV2X3LbmD/lVwB1sHhhG7XB5pXZD/VBiZN
iz+4Px+o/E5eUd3oTLvZnLcgvBQ6EcQ7yaJ1fPHO6jetTVeYGBKo2gwHcnrjqnhSW1OR1nDYbAEb
7ic5hoqVLwIH3b8sBU4PAkjnmiJN85LnmKpyYO6RMyTGE4ESbBUD7PlSVSMA30YZqQiJsRImnFlr
TEIT9cmXFnTetCrY6IwXnv7TuZsybv5Pdr2F01dP0nTzH7aw/8SUeGGZGTaFF0ILG4ci/e6SPqdd
9DZ+UlMBdhNw9C1Nlp2jIa75JNeiAQQ1rP7U7J4TDLjQjOugXFnIfI/TM1XoW6hHASAf5HFlaZIb
p+s0qcGzI2p4nRZn6UIWlfIpCQ0X1t+5e3yW9fQhmvsrFYWJXoLCbEN+Blt+a4BY5I7XEHW8a9wJ
wdnYvEwk/EG1Fqb4kl7p1NjPsRRCqBCG4LiibovBpBPZv6+8X+fYJL9u6V0YDTT+kzwNARMPWET/
4/4D7itHEYhNbyBdiTB8ECIakb3MqOcOV+hyAtTMMqGabciZBa1XXWjbyuUze64t5E5wTrliA2Kn
8HSFSCAO3lzUTcgetZbBAsYjUy7fKb/2P7TSS0KypodzU3oZsaRTtM07t7g7EsgRX+bABnuD3HLX
f2Om+GI+hQr4lY7k3kkv1Jx531+9QQU9gyZFpJrs3up32gWT1ytgXo0M2k/kxhreDiodQEygwMkh
VaJ1rmKAlmallUReoYAdFQJpk5YGjj2WLoTDsyhMS+vzNptRH5cTcz8i5AwBRYwQEVCs2Mg3/2+3
9yYjr+FxcgVTNMz0NjK1k8YJId92Uz6KDhwcywL4wWW9vH57HvKgUNVEXIg2KhGco5aW47TLpk4r
QEOj25xMUE/FeYOAeGaUvOAuka/z4eP7Bk9JO6fv29O3bOzmVuUkTH2chdIYPvCaFQY44MJ7XHAZ
GGc5gz7RCSJvEOMiOdbCI1smrf0N/Fdr53ZKLXpxLZS1+/c9DBa4ggtiAToqgBYSEDcAsrfsO7B8
nSVBIs7EZ44CQZ22wqaopqazcH1RGdeJ5H6pd61dVkO1WXDnDQpFuEiYQWxhBlL9jjQKMFIeGxJJ
gKsvB9hUVTVtnmATMVH/hgpwNc8lNbJBS3llXTdIiRvVGjWPH42roVJMHqRB1Ti3/QfDC7l1L/n/
OB7dKeY35mYs/dao/q9W0mYv7sQU80qpdIA+ufXbvM4G8BON1YoG3s2UwJopYKmgMjFGlC4HpjPO
gWbqnsMcMNml2dejz3ItSeEEGg9Wmx+APKsBnDsFeTkcjNlaJkc2L3hOkEdzdgjVRD0tyX5TeY6O
oFEtmTmXxfFyuN3zd8btEZ9q5a36LZYjJ3iNu3UFuAjW/gJ5ofRenOT6NfwI+XGjDsYgoAYH43sS
0+huYSVlAeo8jAe3GTY5zBFKIBCQtPVshZAmOV8l1uvGdy8qSe7rPvOv0/vzvu9uhfCQm7giu8GG
iIO2yRpBkRAaMxknPXGYT0+xQnskZilb4xGZzwIlQD64S7NpJ1MgPTitchVOfvXYh1xz+13YeErS
AW3lFSrpIOQwvsI3kW1R4nZW42SGDBNztV3CsiDD83k1EnNg0cfkI5A5qiHLdP7nPGFOY0pcpgPA
n7PqAnfpiH6DnB//bNUrUJdf8K4D2PrlHn7QqOh+PJdBGFXvziYRysi/lbKupjRULfQSTYHxw0Ro
q9OcG8z42P7g5D/betJuSrmmq7j37RX9miswM15FXL5JlhCofg+qNIOd7vLN4HAyju+sQqwbarjD
vZheL+k9SyLY/mjoK0UD2iYNKIBcmczDcxCBljCzQaAAMJ0uVbVZOQdOWLqz1ryzfPlXlYG0YdM4
/DglRa4Q31EvyfEsePXEo2tC42weFEqLTMR1istXxAV5vHIf/BNe3jQHN4G3+95RTZMj/45OcILd
mW+SKBv8l4aJf0bAJYumge4/lLr8gwchDTjKXrYEQX3htscoZjUmKPpkot9N3k9UMwmvAoj//TT0
CZvpql1YeJecQnCC0iS21VyFgGifgaovr6hEbb59GjHChudBTpaKWFA2SuZa337kymVn+Fg1AEep
57HZDfEU8mflq4LQMQn9KWHorm5cv9e1yOAJVWY5OaFgmsm7nn/aEv28zZ7V8tWuNnc7i/8UJeZg
HB1u4h0VLUVzD9u4aMo3LeahofKjTqWMQ01zS5LlS41Em/LLVC2k09z2EjHYUpH52ih7VduOoVA1
e+WPhuzkuNo141c0bbNKyaOQrfbiJp2uv5+DMtr1AX9xYZBfb2NuH2L8IxEU3chFaZigdzNQ0XtC
NzCpx/+qrKMYEud/oV/U+xbrZXVPcksloYyEQ/j33Dv+5eLf6dG/AtZJxEfaOTQRa6l+N13iZPsi
b44VPK6wNfRXMJQTj6bmuvlxVqHEJLmGcyatRxb0FQu1bECfO+mnnGcLHH+kPVrjsLVuwD5hEHDg
Hxqo99q04ZTH608IUu5oSEBOelBvUsnMIwtzI09ZQWZWY3XJJ6AyG11lPptqM6kddzeQkKe4qAYp
4SaOVx2oteblAEdyMKzyKONpfOzHXLr9usLzoI+DJ6T9K76ISQRXEEiNpvMLhupTGxI+vE0PzEii
h7sjAXAl0HYbvpi61Ga25WK8j/iKEkFlzSDxbWr3B/Ww94pxLxfN8mpcwCjCqAErkfRO6iwscWeX
UbBfFptWPTLfXruXlIdOTKMtIJ2F4qVOOUX1jjByuBjjeMEbs/+FebGETe12bTHYr6ioNvn0WSP7
h36jCN3zJtDwmjQxioOslVD6cWdRmUFaASg1VtnlHAivyY7VBBRUqf47MPgXYojMtSfMmxPRrH7J
HCeKwvI9aKUYNi6tNbWZT25Vtmop8utkClFkcMgWBXCtz9iSLrcMLh+jS/k/az8S6t26EAj5Juke
cahabQFuGx/Ah5K2dSyJnN0/m88uXoeUL9YYGi213P831xh/mSEziANvdAv2xI7WDaHNngME9xhp
7R9q0SU75kozj+plmZMPdgWXAYeRqzPbMm63HbZrojHCezJEtijrOQDJGxbQcjfQm1FefiiPk3Gg
4zlc0UISRAT/rFcyogSDacYqT7aGbm6zOAvDA9nHxkvm+3WbbHGCefBIwG/+g/9OMvdH/M7qnzpU
+69j92d+nHxn8EH4+dCCBWI0GHEzaLr9tlrZjyP/35Cq+73MQeskq10nbRI5yJpxA9m8cxj2JB39
C6bmjJBYB86pNns7VhUa2wy6IvjOAt1WNdIZNLGUprJlZhVGMB0r/Ml4fo6TNpLa6bTyFv0GaFX/
cPZY43WmNGjBBDovI/ZzXAcizp35jx2z5Fm2hymudiKp/SL6ab3Wo1Z91BbxiaqkEzDIM7bSbR2/
CGUkp16K63/hvXPItbgxFV+kgiyUCibdVBYh4KZo/AXq2V/EkxM2nI1/+cek14WHy7A/kRJsBh4j
krIjq3HDxW4gNAXdhnod4jVHrTzVBoAmHI1ftaC9bBCd6WWEDcdUzePT/HKEQg+091ya+UljhQkE
qZbcN7A2wo6zZvv42mNxdobTxFINinuuUHoy0hz1B1i720+vxH1sM1XnGpUYRcT6z387XRBvReKQ
iELtYUJceCRBwRrFp5YMn+hCU3XW0MirArMrDXV7ZpVpwkcfgJ//TtpsOiCh6s/+zEGpx2BkyIJE
RsZl9vY85yV9mLRW5fxuBUxHr6vOJ+VWfihtx2iKpxMMJpxz5nFTCQ35YQkkY/nmEP89ZK6ay9m2
bojLdEZSgWwpsxalIOTCJLJmS/XTbf5LzF/Dw4YMn0qmoc2eioUXTQIgGZWS/fu3dMY5jRxLRiDQ
2nfDybXK+3Quqz5ipEcRot28/dfVcdnOjekkAQIZmBn8u4tovxCnIR/T8ku9op38W2VEAD1OYSkB
//zIu14m1NZ+CRI5V73y7Une+t2yiJjigPo+ce46qtJClcMDK97s5e9/1BLovdF7nK8bWU1uNkZp
1kpMNdmGxm1stQYFM+dE7njdr33qFZrdJFeVapJFIuaa5VBVNVpg/3cklCWzu1vDMEqV7fCxV2VX
0pRrTjgYbUJ2EyCr+h7ReUZvsrQhW2Pr3r0T+gWDyArSxVqQYVkxVOR0BpBVUcBDiJbHwGfRrAHu
N1OXvAGJLSoJAh+lU/VdYknuD3+T8i8a8RICu/97ljGSOMwega0bt+RuPIPTqOLAX99n80C2H0iy
lWphotfje2vllC0DISNg1YyJRqjO/Oq3SO6PootlYT2UZBCGxjmHJYwRs6sknrIDXfVE6gEivMir
w079WcgyXECkJkR8oFe/4A26A08BD6rUmBnVebTOvjnKHEACHl1/xcEgqW9alVMO/iZ0EkQASbPU
6YvaoPniu0suby8AHemz/6Eh9ZLTaqq7Dv1Hy229SdEiFJl93PtbhQug2JOAGxHARpP+VL/y5O1v
R2QMlATf6WLrRCHCZYhRv0+N31pud0bE83qIEnyta6dbqztf1pe+XpMHbV9d7bJrIDHWbPpfVBLq
wUR/hy8GAjmnn0VE571S4cPOm5LnbRApHdTbes2kyZJolraFhSufpWQ2yHMbMajzlaOpvpRna6qQ
4z54VlneMfPgpBCZImxf+8ofT/jb+dq620A9c6M86UvTtqnVLnkm4jttEUHch49POp9Z8YPWw/r7
2pI42iy5Kl/FfSpQ0GQUjBu2s7jlNYcHZoaLOrGOLhGJVsWW47/qHsx06m/WaeDHu92UaiBRRnGA
EOlhXeyBJE8VB9A81Nu7t6apK0ekSKo4GLAnVGk4ZTOGa+bD2GJFhCsvM17oqDICObifj5A58YJa
5mWJ8GPrE4Em24YX2ANGSuEJ/2ObEuQ/sUZ3zEj8rPdi9WhKZAYgnP68YP6E5EEpMApzL5ybG8tQ
xEmESEybdfDFm0n71r3uWnEE4VCtilPFJ5QG/X3jkwzxt2cj4tIzuqifzTEQc1ekpIOaYnLOg8xL
yO1zIRGYwB0XIkfFCyq+WGJ+m3ahvuulHmWxANsz6GsDUQ9nUReivMJk0eCjW3uhN1D4+4w5ro8S
zK9BHO16fNz9cxmNKBSHhx9BYNASAA3+oiCjipV+jn9NcxxAi4Vq4NeMLrhhfekKnHq0KyAgw2L1
1qT2Ixp+37nFBGVHyabu4HXfraGdtQvbwXfabXxBoVVaPpJo+BjprWmuSzRto1A8TbNi2LQZJp/V
PjfiZvj5MVRavPqgOYU8k4MqonXZEghPzAw9Z7hxSTtkPtYmKsHxDjvOpn50B3myEx2R0cCEebc1
MrQDqlV1giU2GHtU36mlyUD8nXREQZt5B/d8bXwo/kunzXBJ8j9djYADYj6CQHHXsrgKbBgLcgkU
/2EaHLsEVEfV+jpLKTCF5sYydpwRx4UkX4GJ7trsU/fIEAkGvzfB0kgnITWus1cha02sNbtDqw8z
xY9mt9sgRoI/oZpDjv6OJiq7zbPvZeRh0zb340i39/AMVoi7tqOW48SC5J6itHM3yJkv07uFTmIL
UMHtuDOwES1x/QwzYN/ARj5WV/IPAMEPFrNdw73BJA1Yrir0jABlLVD0CqpsOgGS3wXv3a0tYrYA
ZSdemsM1vpnzwNWcmM/jT+MkM7KjwNJSweiArHAgrlAouJVIoJsq7RIO1Rbbweiz2r8XeeXEr0N4
IkifWZGfNmumt1QVnQHpsDYFwMbsFQUmiOm3neioug+Lznrn4cINAwcUzU4+yHeQwd3eDswQxGVk
ffnK7XOWTMk0nWMG+dBD0ls2QChRw+G/AST7M153yYEFk9vE/v++TocxCY7ryutmV6UZo43xAJUd
KVtIJh4eKPic6Qqc0tyQVVv5V7NXYvVZDr1BQgRLZdfJop2bvJ6tQ5vOdQEOXgJ5ityxnX2xaUmi
msgf52yYsCCUm9aco/ryINOxWrA1vtlUTafOUKu3/L+6hy6nr/PUQoeKuYbdBY+RwB2nrN3jkocT
ZaS+ceXQmQ966AkRrgPyvluNPxDmvwLVc2qVHcmSvzMA69BBk/ZSmOBmowS21TwoVGwc3v0TdJhD
e97lWiMEI6ugGoCljn8mZ2RMq0S/1X3wSXHyR6pcUANnI0buht4vROaCuxVeds5M2B54Suv/wWlS
Lv5s42UU77xVZ72wtTh9kLpp7qnb8x8+ZDIxaaA4N61VKuG3m2sFs5kMVBeQt+Leo7/T0vU7W5JN
7JdZSL+Puh09acbTTXlBUxRMZbVaFAOqAD1mOnBqIx2t6RjsyBLRBsHQIxfzZzEGKGJ1455CiU1u
NHVBLAMXxe2x2hETcUqf95OUBWhw7pB45QNbGOWZ1L2vRb69B9tlyXazOuhAmF1TQ2gQbxU0CQ5+
eGytHV83ImJhhvoiduvMajuUAERvxKqq7zHuR4wUsQ1hbUJTvdBKFGb2h4PZBbSF26jYjKIHNO2z
boLE5DsfCvvZOB449bMX/k4BCOZ+pxtHYpk+XMNVzOuFJ1gtZkobJsvJiWFC7be5onqQBi3a4rkS
uFJfsD/x0Tu3Q7iYfeRFBDswlzLgG7zS9cAoxoOv2BG4zhGKg8c7MKVs/MXyzZy5hhdZzdWZaJ+y
VEc0vZfNIpufxggQSaNuqj5f+R4Iqezenv4GEvyAk4Tu/d1GT7kndmQfEMrdV//bMwxz1QL8ujqK
VBVNFt8Ny9c/GmNU8u91xEaRaoL06wwqdDBnSzONRxgf2UEj2xKR+Lh5jQwnOa4OScm9MNXBUfQL
T4smFbqPBSneprF3GTXaiq4/VJAMlOTmCW5T6YJU7/jmYh66BXKr5ySDVwYjw1/eklvOKuP1ZVKW
DFYTkw5odIAX5EG8Fj6TZ45QAvcjrnph5yHTwL5mjrTtnNSwL8wl7009bMBpL/hBTOf7ktC+Q5TC
t0lcjKnlAJXTG4d4ZUhR4gQHCIbHB9oBscdwct21+dQrnJ9eukhJ3hHTPCiMszo6yefJHuDrp3Uz
hxG2jO6t3m7V0L9XwSXqqktjNQ0ioa86UagQJTrKsXS1sIwDE+lH+9PDzHMoef/sYkgavVM07EcQ
mjnni8AE4vo+NUf0TL9Jw0msTwWlH9ZSgxWYAktv2AJomNWZjBHWTznr1ILF5HrGnOiT0mZAb2Nm
RfYN/4qfwelMwLvcEmMryXE+JPPp9SBpPLT5Rt9cgYgRIRG+Xk+vOqjeDYa0RJaIzilubNZUSY93
qLhcAihvz1aTC6WPhHr5yAgsTzj3FfrboTh4ftksOcizLxLFRGF8FyFTAyq5Y53att/piSKEZx7B
fOfsTC+jDBRaw//4zSOV4bUBcIuHcKsVHvcKGubAV8xgx2MGTTUj/NkN4hcRMqq1tGUf3vAjGNxm
6h5ZSwMJeSi30/HEQDsZ7bE9DIkZZoV/urSH3t0JtJc4C1GUL63j91N0np9qg2evnxs7XrM2+ffO
SRXnXvgVWp03xQTquPrOnT6qMnFl6AjcOrT14XasztOSwYHXgkNrZ1wH77fbDv4Da14AvGfNWBOv
yttm6N3VLzp9vSl7BkeV6BWg2MJEvsuxNOsGCAdXwjNcDZPxv59DnRJodo4P0RUIKdI4lg1Vm9+U
inuk574dCStVzUPepKXx+5Yukr9a/xcP7/AmU9fdivTzWc2EPw1bXhFHQmZ1epwYg045mGMOYfWF
rToupW8Eli95IRgj7fWt+l7pmzRzAhU4U4bSvXJLL5ETBZ1E8qgD2BtT3A4SHdSmeFbID1WLaKQN
TP7/QDKUIEXAML7g1erVCdiaxwnXOhQm/N2D0FSwDcN2g6PBQAqLqFNkuDjfK2avietBOGcC+xyM
GB85gbUJl0hOl3EMZQ39tQQCDzTDesdeC8ECvyArr+LucGH50LQKypTHo/LzcfXnJxkrAFqVzqZK
/Jm2vhuEjzX5QUUN1RRSmu3nqtXICXDWQpgcPDOYPwTFbzzIAmlPF8Ll0mm8V2mwZUZ9RAeMgJwb
0bJ/WgZjR3zTzpLruBzycz+uySkXC40s7+OgEogqZ5exFTjdjl4y2CuagSA7GuPBA5URhfZZPdrg
iF1aSWOs4VeXogfFSoKdPT2bH6pTMlWmf7+JR0diEB9tq10AsX5+l4Yu/ABTGkXCrMXKoLdwuX1P
gw0g2nIX0mkROTwx4izsmVL+A+RGxkSSzAsS3viWKNrwmtev5dmtjyuPHoCnKhfIcd1Tb9XzEQB5
mHizrtfei0g8g9HtFrYM7giCQoBIHEQAm1nQQiY4Z1+dxpu5dK0l5wWbDEbf3AvODSVn/sm/tYyR
fSiMLVqf+sA6xGFHmNF7qwsSCT2acb4nu+T37ezMu/ae1YXEwL8WZAlsCQoL0j9uL/fItnD3lMeK
4KyRhnpo9HFfduXOkqJR7FZdS1oVj7CoVJb7DbtveUNYHJ7B4l98joK5f26zrnJbQPzKFGX0miZK
W0TQaGT9jxPyIpSN3TXiuzok/kcZn3S0BsNWW2SjygCtsdR5xlthH0xekCRcaPoDPmdG+06mRUXV
o/88aIML8PVdNkUWAan+GGr79158yC5HOPW4Pl/2AXmlnql65+ryVG9eM12g5H++C9IA1k5/scOz
5CA738gx5x7fMXSO/h1NEVL4qTikK29l7Dagqe/ZmkKaZHYyIeoRIBxhJW4wOc0HthtpUnzK1M4A
3eB52miSzVsoVYtsKo7sBbxz5Tqa6FMa/RecYYKOsBw34GRrju8VyWRFCsrgta/JrlLz5Csc7361
whplxFJ89Mg8UMNY5TPj9sg5CY9AzA1ZbGknFZ402kggLRBYuiawJAuAxhmMDAxnCdMn6yNFIsBa
96zMop4FX5wozho+8T6pNztpacrd21/sFmzAezs8hoVGvO0tIxX4dUxvpD1/ZCNt9xB/Cm49VauS
eDoPhyej0Fqezfx8WkyZOfi4qKYX+RqVTPSA7QVg+KrrUe6cWDOshrs0YLapQlQIcbwnioVa7GGq
z1XlAAX1vBEehXz1tlfsV2nn384L25emxUuM0PlYOFrbcjY95M59kTys2JblQ/U6k+G7lWwno99D
/VvBQDRhVXe7Eq2flqMViV2rdudQPm02VG5nROttjY4/3RB5SWVhm0rJAsWKjCK2hxjjSIVnXNem
Q25z6N4A2Wrd/kwh35Kuog4R0A/QqqDGjXMOArzrlEQhoURnbglvaTYkKXExUs8EBMMcKD0dhxzv
B/ur/+eQke3SLg8GkbL3juaGpRngrB/mlzUN04jDv6piNRKxocvlCHU2j1qX+ys2+Rlh59vNTW+C
JgUIHYeJ0+DHmslhaQBCIyrCNUXKG7pwZJoUDcRx8sIZ6ngDtujVHU2Xrqope80xcD+lR7sMyCwB
cOBl4ooriVEs0eGepnKMqdZhRXJWoBypMyyy8s63dB1/9+lg+L7P1X6bVi8zUpcE3arPVcf9ozvu
Ol0WuE41awsFwslZ74KDCgq4umfTmrNymz5PEXMbiHQdU8DfXDNT96i63w5M+n2vOYLISCj+BXF+
ssjLllys9x65Gy7HD3dc7Jk5qYuA47maXAX5w5gzK8eZh9ed8M0KpqdzvK9sN+GqZ3tUAwGIQmEt
NsqAoo0nA3qYGgt9FsIbs83FSESVdmWznGKOjKJrCFh8L7XpfgRmP3QFfvjA3DrU94IeiE7EYlVx
5cbBcn5GmJoWuzqY1nWJCZuQbaJOOxXGr+zoqHiKLmUZRtUFMzrLpJninHRbm5UElItLZOPj+BMV
Tf6DTF9yjwJRivYO1/304t7SZoicSfRrsxFfH9oUqab5N3QcOP7Ow0yNdrXItDwHKZhKDlKQfCbN
SaW+B2s2jP+aNYY83iu4CM1ED5SggBTUTaC3W9yHeaHcCP4Fd5XSjwx0cqmx+xgHc5voHBfytAau
Pn/XSr20CsM9Rac4aIHaB7VL+5bR6GqeXpEXt/ou3ZOynfhA1fEc4KUR24+YraFbIq6dFaXQNNve
SeFOtun7rbvoScoDVYcVAJmFCvm+OZc+/p+GhSy3VoHE8J92IQfCOpnEDOvSDQmRE8TREYQdJGm6
XaMfym6YdBMpzZ9Xfy0fjNig9rhpETY4ODOwlRAIx5mZ5Ti9Q2u7ScMjdRZJ1MiNpewHll2vewIy
Ihwug0w6SIQDoRKKU7Lm3qDlOSDtdCtLptwvbJ6pQruzik7p8u6PY0MlCsegaRCA777OxPezdR6S
mY1ejTVbo+7zDbWZXMPwf8BXIvr2sBDM7RVkRVCKGObUUeNQGmRYkQAOxKa+UC4rSRf8E61CMAOM
xIruOWxMr8mHqX2Ddd5rcqk+P468z2DMooMMlr4zURN2c9PjTEze9k4YQ8VqcgiYg1og3jvnqprn
5Eqtehxu6eP30CKVdPY2XpZVTJ8pNFBCyfCjKK10Nbw2Ft76JStyipOtgeW7OriF+ByCF+uH17zp
Uf6eVKcADUncbsOa8V4zzIYdvios4tjCxARp806ObzhA3E/gnwk0d+bMmAErg88pmubh2Lp+igVV
sUlkDgIjj7KIS6nHljyc8eweDy9xHVGM2oAg+NAQ6UyqLmGe5+gMvD3TuXjAwqBSlghlDdQ/obHO
eJuRxQIM1UCEinv9OZDJggxjBfpMRETaQ78aHgRf6FEvEWUQrTMduUpMLoIPWgE2hy8TJyWuUAbQ
6Cbml7/OTCtYBW7MtCfFAE/lliU51A15aZ8RIxrVVHcQ69QlbjrdDAj/xAn9YoHpaNZddPKQj/ZB
dWxp2pFd5sblaVeSGPWvxJUejl+E4bQBtRfYCD5zmqDKoOtwHMWAgWzAcqipGomsvu8LpLf16UDf
15J7ZNaCDiRQyM2pxFuLUmC+E01pDBQS/i/LYfZ5UKgCLtRXsYaUzIZw0l5MwlHPQCDlgpHpgJS2
EQE0EdDmAoHJTOImMNml1fUUDPutCgJkwrg8z9V1e63xj6CAhxKRxNQwOB6ZTNCVmL9zNQdFDq7R
vHcidHVwin+/F9tLGrM0jPb9yRh61IDBc236LcXAH8oZVYncY4FS3ICFZvkwfJLq/AyrsdMT3iek
GdI+QSjLNzsyzYosEZGT+7LhJKMMWWdFS9tcGw2Uf+fKZcYjh6UVa2HI44DCCMm2yl/dc5rz+ngy
zmZ4p9Tb8n5MZk6kBkcjPHaB5HT+m/7fHHzZ7lXsw83fZll2ucf6pBSg0/3Tn83J94BbYilPmVIS
3Fz4Y4Oi68PE22fKDFqEG1T61T3VVWHuFz4fR7onyWKf8Z16QOFZHE1z34ax80YJRep13/vRna+3
0YegMG7WSfh2+TZSE2dse0t6Ja0JdFk1GywcAjkyWRnYTINDix3vrblmBRIwUhwkNbNF1V1c6yj8
TlouBRqppGrM4Pq1p/Nn+YGXjlVDKKuHXrT71ZlH1HevsCdWL5R8n/pejALuV8dRSgikuj5wB6fx
/mtYENLUW7F6xr6XwjYq/RFAsUrlbqFFXyz4TP+MFF4VINYmpJZ6//3uUkErAg5VJSCU/O2KHIfn
GhyD9gTDKvpw1/cvIDIz77o+xVLjp5DUpWqjgEN9lqQXBNIP/tmp5s7RP369l6uSpThhArOq0zLy
EeVMXQsUetUjLyYjrB9FfdXe/CvY2Ax9U2WuPpu4c3cehaOFsyWFpJbSZ7obUvOLInD5UT4nRl+8
4I3j+Lc+Py/Q0fvshpkSd2xPJRVmMZw6Z7oPVA9IpjTJRf7JtgzqcBXJgku+bZLD7wwUgk2dziml
IqIu/WraKpIm26EOvAOLXRqTH50sOEs5UcNHh9pMv/L0WZzrZd8PenN6zdPnFeUgn3LS/7Gk3pcf
VNeWJMNBLY1PYgFsdeZxnn4Ef2RtMBjfHuVYlW6IiX1kE8Gy51f0VI10eFUJ+A7sukjFlcERZaMH
KZS8NaT3SnTVqE06WxaX1PqVUiW4vvptWjcXPrUr8F7tSrM48vuFQAfpJcYTVdFJZUb8yOtsxHsI
ZfBzFRejLjWw9m/plxgEaA6SC9qRvNIW6CmNt8WS9/3msVmbcJncw+Py4GTFvncwp5eS7vKvem0A
cqzdhdqfGP+d05vCZrwIUe5DFAiNBJDnIdFoIFHx3qaIdLfAisGeBCHobSnK/o8dJE/Bsb0qFn87
EY8Ol398+GRNYWcZGZm0gyjT5G2+9k69TLW1veIfPpJnepCzUvgjScDi2KWRnmIfAbYB3ZVdWJlD
3yjRuAlcYFuJ+Csjvh03GETXkJrTjFOJk0gosoGDifvM9+HLQNyJxkODndPuIytP5oL4TuEUrSjm
/vMaZ3LUPvpOL9vWxwnoXTupINvXEdugFKzxMn2b8rGZm9rpmhdSldhchYYOyruR8gmrd7n7chOl
MHEX8oAunvF9E15luIcH91iZSQwRBiUuJn+83SgeCtOGyzsfxz89lO4xzlyLVHAHTnYS6bSOEAjW
xt2GYB+wuMLKdTBnuaK31wKEPT1rITOPzRdIUNtBB8kiooYVa9tKJG+eNo6RkLmayx74WsFh2l+l
PHo/+H6ixq+SjEorqdCJBnpZwFGByatLxOidocr0d/Ygj6Vuy5gg/MUaP5bJQNaeYC4SZwdn7Onq
fKtW3CIAq5V6tZaHLON5lQItnUi4c9FLeovs0kGiZEORWLH6KOJYR6GbJRV/loUgvJeAKbfEjGQS
mVK/BzSwbmtcHH6SF7v1lj9TqNhaoCF293oJfIKpBJkOLvIGVMsMUQB92+RbpEX+33UT/e4VE3H4
XcIcYT852iV+Gm+0qfY4McfbUHdrE6VbUlf9mUG0PIzVDGXKU2A0GnDkeG3lF8ZrafUHMN0wzbGr
RPDne77qBO3AVn0dOn17gzpL3WCoUY84swIFUmXajudypS5myhjj5qK1wl8mwSjbTpshblpYoqea
2JpmIYBpKNv8iTm7Gfk4LJN971KI7OcYldpBjU4husxWKaJ/qaX5Ni2cGivIGKKR2SydiwUCR8Hv
kZ/hHx/BmruHjSPuhJE6++4g4EWXiO3Gosv/mAJnmvHYu+JxviaHTSIwHvli87kNMqzu7eNjML6Z
deeUhQUkOx+B6Rfb6ZpQnonYYkjSHGdxNZl8xR+/2/xLBGA+1AO3pkiKuIKuO8eWDJyOYwNPjhox
WBJLOfEoA8T51VkcGTaSrF1RCyPN5b3k/zwi8YsQF455dUSBlkmsY3f/ojqCV7sdluzPezv8Vkxj
A17TyT8iNMnvhp+Rl2OIU8hoWZ82REaj4Rhrduu8CqxRDz/uztKwC4eFAnMMOJD/KgUfeal+keIp
HI8Nm7YsFIpclDLReR0JKA7oQYTXoZavVV5rUsV0svzxvVXDTZ4m3gz3X07csM4NW14TXtW558bk
SV8zbilfwy2d9eZWNBJ/gb/R81HYYigVjJhNiMsOHtINcZQX38E0eFRA1zNizu+bcSDvSez1w7IK
KAky6KzBJA29RDkbnrRunzQKrV7VY7oBgZOCRLSzYb7dC1BEBTGJ+hIOvu1g+M9jNL0B0ensjpfR
S5jdxpNbvNw4lclvYAUiy4alvr6bTTamnCYdQardMTbGW9qp+0yeO6f45m8IuF09ncTIvOHRfF0W
qDZpTiMmlwEnJ6KQiEdIATl8cgINBx+rYQ9Z15UdTalrVxSoKdOUIHZ2jTAvkIfd5kf5m1CadwQ7
dOGbZC/hUlHEU11huXNsTIyREzFEFgS/0AGqZo3ODjz+gzKRihD7irEhA1eWAeSBeOEVZHrPrzt7
N4h8AvsN26OTIRSoQ3Xivakw0baoFvM6iTKq/AEbU+INQuXa6FHByVdg4e04gCpTBkBNt2DfCklS
MgFG7IRpNqOly4zn87S1AuEaaKvC1u2rWkQgp3Z9vBSk98huvXtdqD3wuPfxwk6bw/iWEPQGvkNk
t7yJ9mFhid/O49cYzSGfRKmcyzxIxYMpSHuo7zUXeB4pLl61iVSoBHBnVwWzLavShL2I/0Gbkk29
+jTGONon8clyIP05zcuNBhkRagrcaf+cYo9oo3AwKe7MDfPsIiEgbxzvFQHdGTMQy7akIvH4H6qk
H15058XTEX3y82aJ++5XQZeue3ofBDcPnovsGOvgRn65JIW8V86cxdYwbe/LPPoAAyEnSKEoqIGB
8UGvR16kCR9U3Mfs/564kUIE4n8qFXPkVi1AgXrCwjtCEkQ6dBT3ku0Rob2wHdpbNhZC+mHdONVc
cEbp98sO8y/adf8pp9NrZeQTGMlVDjKR0fvp92yxQTXhMHQGx+wFuoVC2giVY2d87izQ+waqChBJ
wVJTw1ykm4PaHbmO4JvnDXetAU8dsHxZp9sTKWQc11zL+b/R6OgXkzKZMw5s9lxFSsxU0aTPFSif
cZJcJL+RENVHo4ESIuNiu7jaqVDhPWxZeZ9W+cheW+hb67E/XQjZRIqcyYiPn4rlOVeGN5t3mu0o
/HmX6FrkWwRL2bCAwRPyq3GJswDZE5lZRpMN7F3ZstbG04iJb0yfLuPr8qFQFTqE88j3ywEnaql3
OllCFF9byB8kdtM4l0lfubJc3wjAHkxHygsQV5WTSuNBWQwkbZUf31SYww8Ih1puIFKTsVv61DEk
ItXMulaZWZM/C77XVvhGA9zaGP/MpYzNXwfdOUguinwt/hiTiDpzeL8npE+xsxxm7Oy+zWZj2Ehs
mP6HMS0Yoe2jqBS+dUsC8NY+1YrVggPRPBjUNFRxLPOSa3VIGny/qpioUI4Fpkn2SNEe5iw2uLzx
IgVnfgu/yRvQNbNI4PSwxQqO8vTXSRmzXYtFREKdfM+bTLYMdKOKclr914y94OGN38WOOilfRzIQ
RwVR69wvvubrp2Y2mvzuoF4on2eQAmO8Q1QEQMbsJ1Gzn4wqCvP+uxUZnWIiJM76GSlre/Zh/IWt
9oue4RutysG+AGpiIslKicSkU4dx6SboBTa0xxlUDmaGj4Mhxx1P+VMGklEmsqfqkNS4Uw+zZwaH
zNFTu9I+/YuDqjEK64WHb91WAFqFvZLUd5Io+X00z2dY87DDBUBhTKwip9MmIBqkgco/9mHPUZ1N
GRN7TGPgoladpXPHdFADBePXO25SZYQw3RSFTxTaclndSMTs2QG4K2JEhZgeGMGsvbbz6bYcx6H9
AESYq0jBS1FKH1RKFrTv/C1qEfqKfgF27yiVLIth+Bby0ODNI70lV2LQl/rclIFrWnf97spaOYuZ
DNz/qkhadxWoiGrjqmSSGRQWnLuIC7e8GpObzl9OMERuSTT4xL809m5xjbFLgM7ObkMLST1aOojx
SgOAPjYhUsRsFO148gTulQBzv2EWOecc2oDuDB9e5pR5Jx/aGr+DT+22L3Kaw6ksfuST2GV+zQJl
PhKvsH1sCdAh6JGj1mHVe0izwVii65LZbsW0pceE/l+WvmX4KPL1+Tl6bcQrq87UULOh4Uv1KTn/
uFvMWzQLHvGTeFCbWHI1iDiDyYix9AWm+6KRnhL4stREdu7AoZUhci38zqulEpGSMcq2M6ujjVEt
ZcBs++gkIBGt6ucukCc1SlUQLTY4nqjbVTKw78AIyprSRO1ZXFZBY7EfsGU4igwn7Z9Q5cJG0vvn
0zW0HCJoq0OtX8ODsYUzHtzUyLgFraPnCufjgqUiX5jnAqpOiyKszvbM7jfDLRlHk7rC2MdE8Mcq
9SGUbFSO15NB7TCJjVdawsASoyCso0uKzO/HZOvlNOKFjTlKRWykaE0weSV5Zm9FzcFn6v2YIk/i
hKMBobXoj0B9T6aWTUQ3GnQeNzdt1kAfoH+1b6ev/Mtu/nLwFefVDuNz8AWQCMhJo+AvMpHMTs7v
w3C9lk8VxgsoPcz1lHGGcjMDPtO1PgPEm+aPmDig9CBFoIUGHxSbS9Az2MN+Xm/u5LTjBmccibL5
nF2VRDdqVlJEWAHm7SmUjTfXeqTbtyxeudyfPuDRf8RuD/WCyynM07U30QDeYSWNCakMHYR6+0tk
+4KEHrumTiI/U1fuXZR++kY7eodoILVX/EKY0TSYmbyo05ZxTxPZp525WtsvEFknuxgGAWFx4GTw
8zIR0F7JccKudoN2uraJc0wUzJtPVWNEIhS5xioFdb3A+g8UZuc50oLzSkdCA9a1iX4MHwYPnzaR
4EZhKYgL3XiS9M2pAzifgjyWz8X3mTcajQGURZ/pCQNQ3qQDLzutg/TZekmQgICpn/5OYi0Kw9mH
1tUPSlqi1T7e1Iq4MnYYF/IFP2+2vL76t5qs2zkCP+Townb+bM1YbZxzmgUH2GEquz7NsaaxE3C2
/IPcEkF270cz3pK8FIh+F2+Un2D/PQhHCPtraPFojms1vEM+qxxoYvffBT81ILaVN+3SIxnOvlKr
u4JTWrb1aoVGCFqmaO2bZ4Q4qNqNgFTsc7z4l6RSoKId1dNf4EYPusrJk03TClmlLqjkmtcs/qvJ
h5nsPy0keKtUpDrVo6DGleaYXiwQdyD2sjjqBZUN+WjeCDf+rDekDh+hzWPIYEPAKhBcOK8nDbU3
N/SwTGni8NRkxZPBgye6eG8y8blJcRUkPtXqiPxFtUIIfzhIS2Ilv7OARqpF++sbXp0Y8FMhc9dp
wRObOF5zAQcL9CK6F64CcnzHMMu6I1HGaysqW6n/yP5XmtBz9sSHHDE5XjyUdgaVrlh6ZYofFPk1
ABXN/W7a0/QFaZal/Wxb7XH+S+IJh/E79HysZIto3DJWiXrr2+6yhN2Rt7dGbdRtlXsHlmTGDQYT
KAS5MNT0/IB96JVWNbwIqJJLsYIaFqUi5x7s0X44Etqkf8lw4pvLLDAkLGs7US8iWcS5OQiY9hVF
BQBu3HKmxG3w/vo3FCwCuXe2QjNeh2ZlkLdPG6F3XJrSQeq7VT06ReNWwvkGAtOiL6tXQYHeIxF5
REWJQE9STQ2RUKm/c/VPu/GODc508sawP6AVqFnhpEr7COmQTEY4FayJNTeMU60fYjDJcfSwtpHt
z4efskDV2tLOudvIuylRLetrV+fVNLnKWP5X7Fn35lEknUs7LxPzZipXkiVVNaxVzCmG48gjN+Vv
4RqhQpBGOkQftBGUSdyo4gHKSRxm7wHaRMU/jyquMDWs6MQio6ElanMWmnWGTZhGtXrGfjamIk1j
9OUhm+rvQ+nV3Zs9z6LpGGTrb4kzj8xsn1dX9c8pUn1wkTN+M1FfgOu2LUX1SsXugDau5FZ+Hrat
gQGKxBNAp8CI5YjGqZhrQOzFWfjZLKl5+bRKgXKO7721mmBrsBTnZVXZRnwn9CCmLT24B60dgoc8
f7M0VCS9r688IQRTKP/BIFH3nqff99Iu8U8UPDL4bY/drGL5YDCQjuI+XiO1Hr6q99h9z0BzlB/1
bDxviIruVzBQmbrIKMSCHTznKX6mBZCRHjz+rmnBGDmiB2sC+PuEChdBRXLjndnJpkYufOM9gVBm
o7XdcMipKV9jOVi4YfXqawubflbJN4Gq7TsVNt1f/y02QO7El/l8q2wctyt971pI0KUYwrfee5/Z
B5+/y8mjeIBEW3h5JFETSI0QBdSg/ST8MnHgzVsvEvjEqZX6+B671zNJmRfov9NbzYi2L56Pukx0
W2lcxZg7JJpSwcjwnwahaH1xti32/qpkW8sd/ZWiE8FcFv0vhadbESdS7JhJRfECjXPuJeoJN274
g7qSYAmVsdClbfEHrz/EXbe3WsvvUEojI9PWVBOx0OvU5ME7/JuSKSKs/EEXN/5a0JbooHduFDAG
5lXVG8u1bcJT1wzT6BKrb2SaIb0xR1fLrzusceJLbUYZ9Rk7p27VBrmM8swlA9ZPA7gHV6IVpaOG
1HjCGqoM0X8zbUDExALn9k/CHBaLln9/+lzfeXd69iEj3FbPreXxOeQ0xDDSMcp2rpZastKr6mgR
EL5Zzmo5fas9AaAM4dBWxcZSJBIlFPwdn3X4yuHrM3dGHXcKNu7U/bHFRbRzLMUPvynzJoxdneVO
ssgLku/8fLYaLjiYcOSoOYtR1Lxi4FfL/AFo6ZDjV6FXe4APkPcPGT3rAXyM+EmnrpRTkbmKe2lW
hn6x0eWR0PykmSDVuwjt71htTBPm5p+FxgEHrX57MCXAtzcKzStkHRK60yYXmvY2ieqHjzjno611
uvQu2fzGAkef7pQRBf8OEQwHpn9gJTc13r3RsRoRFuvAiCPNMhh7kGQZxPE46prm6lDx8OetU90P
L+Z+cdCR060U1tyQKfQuRkOXqVsNghOzCuHrHR6c1WNYQMDSBRxPmd0vWLF/Mlxavt0eGj4q+1nF
oJeQF6XJj0O1sss/Fb8HnhPwcdCO7uADMTV2TwYjbtsp/2k6FZcwKFIdsbrVkc4lAn6p4DSuuQ1J
d5+zmOCR84DgMuqZysf5RMO1nDS4tL3fESJ7h5bSj+8IqX80IMn+WtMhsS3yc8cQp+P0dtSyYjp5
wBaFAukrROky/oaoSUmiqJCMBo5OLGmLk765K337IBXEuKlILS9PCWpyGrl/kXLkWOZMl40vhZoD
BumwrWyPNSsGDTVL8IUXvJbsLoc4+7BumpMXg7WrmkTYtF1LwHeaGSQzKWdB1BsRbFT6iPXton62
WeRPbgLAokKn02QjS2wHTzN8h8gb8tOOepZNF0ScJ/HM0no+mlBPdZ6MqpXZlzkWtHT5KL+kRR/J
psGodHNYtHMgflAp2S3Fl9y4L7NfZ9Azj2P2SMCyjkIddkra5zZkHv2co/ucTZ4TMCVLzTRM4LLD
ecWSfZ8AShHcjP17GLhipsc+sdO6Jyu4UZ5lgNRa3K46fLUdDiaSTrhjMWuAdQgwNmXMJFg3wN+1
/Zy8mwPs3NxchXAkczzx6LFODyohJXDZPkpb+nvBAKHEJAI/wS5WGv70UCnLkXdOI32s+/vcT8Hc
kTrFG+xTP6lWWM+dRJzT34J07edXbUEJSQ01ZgWwTJEgSwQ/INSqHd0C1SYDiDZzAvsyc5Efb4Mm
5cQjXgdgDbaaTTGYKq5prppgLoFL0k7G6mqiKiVouAB//Hc7+OmA3Xrg8nyu0gp3uGXKD/xv28Yp
ODHI9OaB9TLzfq0zVMd1CvH5qepCsHajuZmAa1PQbH9wqUOY6eGvJYG+CJaqI0eRMnljIcZEXDpF
/BrUP0nZ+ygYRVJyoHrQXnSxBlubZ9ihpJEVOnvgqktJqc3hJWbxo5oiLvDE5l0muA4h37R55uoN
I+y+D7klLz9Cm4NpwwjWhNSw/2gb+nBp4sFOW2QnET5CyFXUw5QY12+XxKYUMCeKKOx7QRIlPvjn
X62v4RBEk14nn/8ulML9pCgCUzbaR/+WuEZJG+3hvo6xvZ2jlpYt4uvE+VS0wIaG2yfpMCM8jiD5
xR4q1vwS66CVVmDBYhOAjHCWCpkHb9slXHiQ8m/KBOOOIdqBOlhozmDIncO8eexB/sKXMcg3xdPl
a04jxqmTtG1V+R7jIbV6giPkGUyXSoftid4zABAq/oUhZGf84A9Xs9FKTAZFSmDYiNR3QTSTUIyb
l+LuqSPbd0VfcAvVcJXQ2MgUeFaHzZBdK7/iDb00eCZIiHjnmjv9buxVXpOOC38qFiipxH1WWRZi
4GQOQIaWIUBCJKspex23jz+Vfunm6Lcxo+AOCrl3ciUsdvW2iEM2bkdCFo0U/QZbvVj6ucdlR03c
zoR8tP5vjPY+EwA/ruOClTkRiR7zohFKJASVUutCeRyrYjEvFXgeXRq/pPPLXOwxaVhLa2W2hx1r
coOUVWFwmQDsNLjcC9gd6tOSm2Qhtg1Gpqia5xYTjbO2UWknu/pNlaypaxgUfBVZ2CdSuYLkR/xS
+tQbvoMYIy2+Szv2Fo7vGXVZ3/gxAr0d8s2FkmLf214p3hLqeA4LYMDoOq2T8o21IN7MsmkV18m4
1wO/THxo9RFBdIKga9gTFBrG5gzYsIlFCF+y9RBkYo9r31K6RYskgv05jn/DkmwP0cN7r3zrjA/E
oHK+TUQ01aFgo0vl+NriGD58KCHpkD6YP4DGwsk3bD6ZMvxvxSU9p1ptz5UKJjipKeW6Ed80oVuh
9E5dnpa6pVhfQA03rXDEO6I5QD7BfmITU9M/PSJtJmtIzpAEaBDtwwf1q31MSDOR/3MektcIN1ug
JdlOtOFOQi9BVrNLkcnGhGEky2wU7Uoqx+egLmnlBZ+hHLm+74f2f7DjY+qT3uq8tIWtbOy12F7H
W1LbCqSR+XcM8Rp+vkh22cn7gtZ8p5Y2G+ldzIN84Q0TGCvUKIFy7l93rxOhvCdVeVTmsSncEBbe
lKzty5gFq+WnnV/QgH4PbIY4pjG54GPYoRRpoqDdIlNl1ud8RXiu7VRHp8SbCFR6kcWk6RjtcufH
8Zj+uzwQctil4g8jud6CGORehOXzhiZls199hSkbn0dX+Kkl00LKQOwfRoA4lsZdW2qfOLFmFpIB
5D6EK6We8XUe7g6U4BrIK4iwhhgexQnmtWMv+kPrSFJbTw6jgc+N2b4Az1tXE8k7jlprCzJAcG3l
JGs36xBclmmIVhpaqh17P/MXcKxafkLCLgSfFiKz0PVXycVJDvhdBTMZlzrl1+SSPDxkhsplgS8J
aElqMf6z0i/9qfSAWpw5120qAOuRxjsZ8zcGlYn2iYPV2arj81UtWALecX8ALlxr0fP60dhsn2oP
rDrfygQWdpgZDRPVgcnruqi9JIDtI5jj0oUE3iQBMfYBnIbHi5/cFWQp8bdMTnFCzHiURs++kCo/
xTV8L0Ftj7Q6vliufWfZl4ft/JWcozczKqiiyXAL010lvBH3dUt8F5PuF4ICK5FUd3g+Jpkm1MQA
b52pc5/xuhW2MsI1ouRP7IzQNXMwJhKfoUEQ7Oy1jnJzEi5BRv5JyjE/WlfhgIDNA0tRfOkfPRGh
JkYxP37m3xhxS10jzFoxkSHPnGSi7KcN4hiqRW8AWH4q+q2SKKTYkvj/f9OGEZ3alaONUf3GiOKU
lHz/anZiDxY8/tvv1a2V26JPklwWhOxYr5TVI0V8Etr/As4d7qK2xWUknfIsRjRBzZw+L3vmm9L7
1K8Au0yKTpQkNI6v6gXpzm7tCenukVxgE3sc5jkOEpaVOb/W/ppO3FNIPZ+gJdcmKqZG/tPqIi4v
EhAapV/MLVK6G6me7FG0h6WrCOLWt+Tb9ENo6ajYelE5z6KLP8GmIqJCl9XX0u3/Mcu7cRxIaNFB
8YhDdMubcc9vJEbsHZyRriYrDxrDlvlVWzokN+5rlt1xzBddOQUAMG+EWmrfD3LXpg0+Nv/MYDNp
hlShXPVJaeY9076y+FXi6HvT8sTkl/OxKivvzQPp1ihI9Vlc6KgkCDQ6xFy/2pZAzRyn84bwEhHY
ByiSOo+a1HHMSCZwc+zhoEhPY2tmDeIamrMNN+hWLEWcexa6kHSpsWg0rvuA9J/T6cTZcWy2NbFA
zjUAqNVRsyaGNrC9YqnT1ea5vvI72cSdMeyG0ZfUZbu3EJ/D0ezTreMykzmFosFBZWy4L5IbxqN2
JtqAFFvxPicfJkwIapuMX8hBOOEYkHwyNPkJymqeVB9IJoRS2S50+xblOVlgVFFjYMaWjgP50H+A
r2w1vzMkrd91dZeaWep/sYmOaYR3lO3pVCjRBq7BK0Nz66AWO1xeNdtV/8h5p2eRvabzMp9q7S54
vL14hhZGecal1OWZMcezMP8cr5fQpLr3r2YY1O0lLTeqDhkib1ewPVZTfQ6tm6XTrJ0mA7Pzr6LA
ueAzQ+iThVs9MEwWpJRY+lAe7V9SMg3vDbaie7MGzGj0YUaC5kBOAUr3syhlhhMMxDV2SbNfw+Eu
DjC2WpgDoEKkJB5Q26EGblhpgbFpKreuWLW5MW3KHSmA254KJCpqFuLtM53ZTqtiUZF17rVxPi0a
MJ4RzDHOhgzwJ1H4MKgJ+OX1tgWrCter8ekg/5VV3Zhim2c8W1ujQWjuJrHKN4xo+MJIzvfuDnnF
NfdTQCgZ0ytpcF6kLjkyWk+Lx3015vxc49CF8ErGS6zZwlQlxExC8vZCw2WQRvE7BiS3DVVcCD0B
nrr1SvOnKqeHdaD27SGQZjZm9xWJ3M3NGj1FX4h44FERh9i+DbRQ8wKZvX8F/nrDYmkhObQ3tdD0
rb+tZzrZ7JN328Wh1+V3i2YWADXRERkhYH/Y1E1OypZu7ERYepvynNPPQWECtjwenpiZOTWGStbv
3Slnhe/Zo6hH7nSlEC4LWXSmg1IxeD04kUUkajwh06P7gpUth1vDYGzfD+R5cIs3AXh9d+w9FsM2
W/82k3zEp5BhJl84zz/1iKn0LyEJq3PVC6OYrSj5pR5C4GZ7ILRVreDZ084rChy+hepSYlCZfAUF
VQzmnbjclE4+nWn1ds9GkLK+yXn3MQiSJfGlTyeS1JjWahc/2G6HlMOtM83chFUnuZGWs9YphBGC
to8QOoImNOkWpVBf78l1vnZbEOksoDrKTpGchH1EQeKXelfwnGQhm4r64uqRm0Wne2j9QpIqoo+q
CKQfu61oldiGIw+ZIgLnARdnDzmeC813iicI05sO28ac1fFYNisZRMVZveJjAnIgji3Qqk6suLF0
yKEEGIdacQB1ARIxuBkB0iIpfmcyzOrXnRFO9Kh+2/+8mw4smSSoqgq0wZ9IIgG9HOrbL+NCd9un
YuYXG57vyOxlMVlf2YelHiPJjUtkmtA0vyQxhoOGMc/A0bjqdep620FedY2InLBR1SGWwea6kKLX
UoDEK4I/tr5afkxb7waQs3QfsphmBOjlHjdgfl1Af3biYC6zD82DkWsPLfENTG4YHpD1RwwDifJn
//rJB07dLXjUe+/O+TZ/icRWhSkXbTAKKC7tWWc1vuIHU1UAQ2/asLYyJ6RH7mQodbFbu9FWnRlC
nUAt2b7+Pq/wpMQKg3CSgrbrFhjaykY2dh7PKhlEsmFu4UQXsrIVqEPXGEB5r+KYsnLfGFQtX1RB
8F5z8p1ulDDVibYx0K7D+G5iaIBSug5NK/ngDLAILfumDbq64jwcnh80Gu/R3mGjRtI0WJ7AJQ9q
qeDItIyEP83s3ceRr4OmNrixb2X18VeRuKQxQZid1jYpLpsQt7ZrK8cZ9zibyHmzyOlpkqBRV6sv
F2YA82qqnkmmuITyuUqpln/S00opFAZdShMhWvcP08cDSNg53hpq1jiEvTZaERGd5w0FAfknrmVL
uyvuEKIIciPj24lRuXNw6VAeuxWCVcbOIVpopozzvNelWBBXgrzbOfIvQ93m9MXMZsmxWa5M0Ucd
o3A5EqQGOiBlAo+4dZZECxP/KkEWYdJ6k1nnBtNp039JkPvqtxbQ7YIupMRLTaypO350+8HLrcWi
ggBP8J6lXJdH+TCylarj+XrN3VtSNR/jRB+vecMujbVPnVPu2Vsd5GXSQigsQjn5Z2SGll6U9dY6
oHUdW/FHBL/W8yIrmJ8GBaC+tD8O/kWdUX6kaobskOn7OKBSkGUrlXwvaH6kryxRG1OTXnmP9TaO
UZb0/RQL82QV9PqdaWamOufOvlAmIvZ77iZYGWMNeRyidtFuL2iLth5pcmfpG24zUOF2MMcyQgUC
2Aw+1k4zSz8OtDMSwpYkecTGCS++CNO2FWVP7EbMo8B89bVqqESxVc5cIfhY6VYR6s8fEYynRPKR
Jdizs4uF3oXPeiR3DqsePPpNRwp++EGDan7xHDde6L7NtlrjnaxPQbjHH5NmW78uRJbwqHAHQCDQ
iIZJXxmFkixTvpzpIR9TZHDIj2tD2gB/Im33VVKsY3WSY8LxYUZzHaD/eeR9v+gckwv43Bea2L3d
Z3E2Ou457iZov/O3gjs0R890BL0n3thrFqA0WFomVKF1CwwEXcyUpv1JRjHIpbAg0r1QR7K9D0Sa
j58cxsWumr64DuyAVZdhygWX9Rqj2+eO28C37V6iprBawEQT2f8BleEsvZZ0pSL8eDTnpnPltcs+
LIMMkFaVd0KkDt3m4PpWuS57r84isWEl4dJrA0OfkcvFwEWcpp+JvelYAF0nKxCQupXe9RcPF7SY
ohhH1flNHNhuYYPxWUQ6AsGrRstSmPyyL7yvATMf01oelsFfwvPUgRbmGQ3ottU7qpjTwa3HGKiK
8t/i6LGGLhapie+dcoidZsYluSgqLaIIA73y2amuHc/FryE/cJJLuBdeqnTyWw85Pj5ezPKpKhNs
/OKj/pNp6K3+kNCv7ff1VaZDM0fD7jXVtybXDuo92SCo+aqU4J4IFCwYV5bMrsDzX285o0BZi0Ng
qKtSpFDyXGMgANJllP0nBRfz2Jx12xnKi1v3zM8uKbnUmkM/iuvt1Kl/ZwMjmKplEuNMtGQ/Qp5B
AsCojKg72qIRpBpoIC4UDB7w/0PMR0uISfupQRmzCVLXtLyr/AsC8zhvW/EGxx0VXX0GGDv1x70S
Dr42yMZbDbtRoZY/DW4S1Ey50KlZ25y5Adz2ZorELCAm4T06ZdIBrO3Xdi3ORH357PfoDldP+sGB
vh+npffNudq1tP0mke7a67hmlP+zDwCpGPguiTXUgXwqxy4KJi1tHZXv/u4EN3Sgp5wswQv7jX1i
N8BErBRVPsv//qw5QNmior8z/wuXCXYssx7RkaEXamGFRuoetDp1LnE2fifrUMzhpWypr3+z/do0
QvOgUjHc7ooR5kkn04FZT2j84kx5yZdj85JzMtA6LYjll0NJ4iO94DIfzG78b50RTAcY2OJfdcbw
un7MWnveAvEC6TQdJwteXRkrWSbsO7b160lPoy5BtW8yF2WKvU+oJDd5uC5EIUKzJrlr1TTQAWBy
gW+LzNupfr1AEL9Eb8laFsMkUeZaoSeXQ68HLC4a6QMXiD7Or8ljqbwZTHPvePbs5ucusMTTvPLa
rSlUTR4eQjgWy/lUlVPPzc81yiUtK/bYtJLYIsmNVkvioUgAzH0lkg4EGeSDNkB9bEP35k/jasV5
m6OPO4RHxfsZ0l5aXDabPRQy0O+vCsL3uWQlJ0sudNeAl/Cd2b0YgODpHmzLCnT13HXxyahdOM9j
qc+VSuuGY9UPmnIzl74hUq08RlupcxV4rJPPVxzHQ0k2hfHP1WDatjFWTHlcAm7s1OAqxq9ajZsp
QBCWodvVzQ/PzInXLDVtLZDvR/yTImSTHmJGad/GK/Jx87D6fLh7AGYCazr24c2uf40qq0TjvyiE
+KxS4FHSsi8MlE+qjWrlSyapxCxCJooEBRQiKsfBH7wXR9wdUA1m9ZoyyimyqYAG5fZdqT8r2mpt
g9OGH+CiwAp10QbXgxdAo43L0hBOdedIFVuZXZc1K9CLxeSiarK7MBpZIQPhtHQ343NBql8ZEWDR
dR2Fos2OP2IRx0b1Dszfhqe27zY52NkBC4mRG26iaxQeWfaUIxM2YnbBvuA3ZmvEVEEF6Fr6XpP8
5tovC3z5rAlpk2kRI/ig2AN7j+JN6t+BC7LkRo5GG/wkXfMCbN0aqxN10HB4vfD5WaPX3vOyu5a2
j8pNa2LL1YD9jR5J7xskU2Rvc/LEsX5jtKnanJO1JPr4Kw5Gmwfe8m9nkHUipIWJj9FWENKTP7C5
jiu0UbG0TAeF9D+VIggrnC1lm9yxfVn/Q6eFggsAkm8awjNYZ52iSuVDeu65dFywcJy7Z8W/aJgn
ySDjBuznXLHW7Rd3Tt8Gqse7HxTaziyI7HvT60trttOTt6WN3bzQ0NktWeRC/B3N8zyv30AOgFWC
/jrJlrBS93ZLil6zTiJUn5VedyJ2QoGOWhwc7jY7Z3I24CAb5ZEwKjg2OhU+iKEqDIDKtFNL1XQZ
rMw3dBHhdF64wSCCopU/OkcAOVY2ojL6yvz/pNkB72uxJjiZ8P6YEAF2FuGqKA9CS0bWY5f8HGD7
dbeqoITnNg37iFA0906FjQX1JVeccxmWN69j4K8xhEsa2Xjw2t75obEIDGkjIXA4Sq1AKR7C3bBk
PBPymS5a1yJmlS8G8V+IOKRk1svTAEJA0uSHYHXmBvytVb0OC43LVcngQc/9zWtAsPQRMdbIzfdn
in7atPTmbl/h4pe2rZmWK1JG/BTZ0DhUVl2DqIoGjQEkM3Hxv3/x1zUvP7d1v/6CRnFk2KUdMd4v
ayOnYZ3gAau1YlqvfcC3TnetI9BbLqzjsxOksUscFiAqcRzGjb0Pg9aI4RalLG9xFvtqGglYLC7v
l2CgQs/GUXB+KmcnG/A/J8pfuRy9ZzGet4FwvPZ5Rxr477hNV5L3ZaTx5qAYELz+NtNU3+4Oi49Q
5MhwdDKFaN28awtponsT+iyknnc1HWh40TN0eizMw2oQTyfT5sDOY54LVDmK1XwvoFfE74pSo2AU
faKCOI+ca+uQCBd//vNNAxC6NSxCrHZo5UFtDksWvvM+wvD0At+cNfmN4NJIClH+Dqe1/v7LVw1h
XeHHwxK138bBSICpGM0boQtQy4LhaUqu4LIyrz94I9/cBIUjIycPHNUQpY5pSJ+HQR0JWJyRd5CZ
/arQeRHKpGSCdzWkvGbnQUeohn2cG9B6sdejMOwQgG2Fp5ivzUtPCRbxsuvIABuYSwTpXa8CXqxE
qXR3syONvwxAyJkDtXuKra/6KDSOCqSQ/UzZGtUtdS7fRI/DEJmkZQvtBIIfoi2BqS1DEM4PrGsQ
+tfFU/YNY4zBe2juQh6xPuY68Bwu4W4mp4MwvwqAh2LXA7c6jVr5Vb5CYMH5p8gdJR/G6VfQDvq6
yrzGMmRr9bEHfJqjBxRbM8mjKgykNVbPWQgrl+69M6x0CVBqgsYI079+XUInfpl3L6CQW5x6pfM0
fy1t9l4ahNncuQDb6RPDHqse0AXxq01J4WkxljA/eEMQ70Li9D9XbFqwP1xYFOr7HSHjH9arriyy
yByVgIBIflMwc+8sLLXgLgLngw68cJijxvWc7tEIn/3PPvoSQ6vgUIZsz423jO3i9Cd3owhnx1tW
O3ocPuyhxMMLWNDh2gthrliLU406KdGRqFXma+NAvFC/NSTvhBcMnzaNnEHkm6Ozcv/5OdgF6a8s
xdYNmK/LTzWXCh8nQXJKDeQ5YIKsQxo189M6Flgfufo3Y38GEOCkw5C7JdbVpuw3iZ1iK0WAWRAB
jlKYCzh184hDftBrMvozMHSXghGTn6yieQv6bz5ZXcR0CP5BrmxzDH/0HTeFiwZ8NQXEfPPltYGL
PyWn0x83lQxeQJOD+5XusQECwcMM4UMUpv8zRAzHYXssu5hv122EGuQgW3pMCnM2NNmpOl/KRKN6
UB55Tt5huBwl17oqPkVKCFQgiSA9SZq73r4vUruRlyRETBQ1sq1Nctueq5UhmNDIGtq/FP0VvZvs
+Z+p3TtwKyNo8YTLiQ8qbE5X793kglQz9c/lT4cBblWuZVQEBWoghjR793AhdO+HYbZu7nCcw7s9
wCSGmKlGg3ASeOpLktyEHzo6od0ve4lLJQFAZEfdaw0GJymof3Lx6LUDGtTG+ht5uAe5kfCSxKhc
/WHGbFIi+9mUjY/I1jBICIXrDvJtJYJ+sihQ5qlF4Nw/U1UoO2+tOlqbmFdjRDQLqs+N05+YH3y6
lfqLUSnKc5zsiQKF455xtI5yB70dv47A1lInkqfZWurdfF1t+VfWrg6YC81aeMvXIumkaVK1zzCW
oCuucbmsU5EFhSUTl5kByz7zAjQHNvFvW3pLEjSJ+k+haW0lrbHJSSZehlD6vCCLGoFYHrGd4vCg
BliqbTF9BK0F6RwbitU7TO31txmNkxBG10Jj9hKC93BqFTzTgf3EmjI7X2I+B8lLRvoVpvYrbIrO
v06vfjYdohnIlqzG9xtjFsXZg94hlAVM0t3I0Vfze0A1ha9Zv7p6xk6AI+z2Bye5NPDGjf4W0H5C
BriSQ+Ubi8zeyLOl2Y8TGwSpLpwWmbM22zreNG8sMzUwrbbQjY3QnKfb5EI/+2yeqH3GcMU/SSSJ
iK+IgFm0LvZcOz4PxaPJnp3GzTg2oGY8/aabYgyS6bPnMrlmMvOpqhsmDZu5brKxGTWOpyT4u/PN
AY9ylMZcEMVUYIHgiA9XMScRhKQcRXG2eHCREn2VJ+rv5f18JojOlYMC85BfzKA4JLogdRF8waY4
1+yzwaxOxJf4S2u5NYiSS/M6DMHhxoOniO69GYVJRQe8QGf3qOu+rAbvZVrlEXW5iJMoHcUWKoX6
tI1/3eukcf53hNKnCe+IL5YBEBCxdkq56DvCFZ+EZxiaS6bET/qg2MnjfJjdpnCa1JhnYm2iu1YK
NszWnh6CBSvOPN6RKZu6qUkprHVp3k+tdssb+ELVQBCwheQa9Q+S+3w6OopWEmagrTWJwvo03RMM
SyNK+mJERROoUEtSgpn8bQh2bapi6x4n/N3SWT4BdqFtwNAg05HSpnFbo+Rfg1r/c5JWwDsxGlIL
zK0HbVi67WYi7J5mO+ikaR0oRzn0wWMOvnCusiGMwTwxEM18blx3EleHyshkMxvUCVATJ7rmnjud
OnWEt4YDykGW2WAgeg2gyqxhOL3MgA9q6RBdPhGJaA9ZEZSzQsjUDYKiblrjXtsFqn0zTKpBjp3X
JbLXCq4cxkSXdOebT1bDqchQPJz2rOkhfnq5ejDKrwUJqXgjdj0j15QY0JBae2cjUkFqg8xBcLkk
aY48cu3DVutAhB+Z/geOrd4OWiJz7bWhKZOsQ2S98E20pkG8Ks5DVfhz4TsPxvpHCF+vlQ9QYMWT
dL+l3ZoqHas4IjnHx5FqByA5blFPSIAauot54zGFduaUBP/2eGLx4RV7Vz1fwex19tQ/4N6Meown
K6h9H/z08b3xBfe091W0WZ0TTMb+O83cGJ+WVvmXhCN+r1U2JfxvaLTqJxlzCpugLCrqQjPoYMUi
iyKTJOn5XLHb8nqmFzCY9fgKX9iH2PA3070CiBkkVYLqKOPB/cOyd4lWVlLFVxCDU1f2DeDqbSgD
0dFW99KCxCPM5zIt/wmejq4hcPp5+d51gUo9CqxGEh8Vg++32DbQcGjfXx9ZVa3RqzFVB+bvUW4y
Nbcdto0UB/DPEdtGm+2CMMRQ4wJUIIh/yM26f4rQS85j7iP7yd9ZJRIxNBCcd+Iq7sNVgldi1OYM
bjA2zv2BE8KSF1YI0lrdMOHP9fr/v283ntXX5bCdgQ8EZKtiuea+5QpoZyaGutUqnOwyN5x9rjOF
D2Wh05dP2p5J1gsmkuduQSD8WlEzY2l2Hw9EmBI1/5rEzA0iJnhNUbZQt4CrNNDB32fwmfH70ws2
oirOlP3hS5gpo8WE7i8oYrhPqsYFCz9KqRs/VwmAl2dD0ICmINeZLqQd4WXcARy+SjwYWxq6zVA9
NXy78bNdxSWs1an5YbtYIhnyJ5+FmD+4YBGMcgouVtP7xq4CDtKWSkQSgm9dWXbjo9ALdKgFTu4U
YHl9WnAOR7/caYQknLEBmjYyPOVACu5enTYe2KrKV4LiV21Kq5L6YW8E/3xHrop4ESyBVoPBVA0F
3QLopk2Hh7v/hw860B8fif7n5JShm6Vbh+AZjqERlwP9ZLhSfirFIJ2fpYi8fenhbI1+cq3z2gmQ
Xw8GfW5cEoYWyZ4PB6N4a9HoGUgjXtPAKu2iN+pJq4HAX49pBo3R78CpSBDkm+l25A7aV7kA6vpe
+x/yGQ21HvfcewP9Rk26J4jcT8mXZyBJuUJbHoQ8wJ1wijkFWAHLSshm87l5KJkOHVM3Ji46As5s
WKySZB/FbpQtO/fjAQV03YdMyZE/+lvbDBeitNV8phz1ZefiAq3WHK3Rnz2f2jYwQ5zw3ieBJ/ak
fe51TPsf3xXj1tvipy3lgmoKqjKmnkh5EplWvlHGWinX6VmOml3WBpRQQzLEUUjM7F2ez4kkg/YS
SCQy4P2CGRVky4d4gRUwxFbyPYXQk9Bei72SeFcSNgpNRJ5mNkxAPRHlaz5sT1Jtgo2fc4o8Qhon
EBTuJKqLKwvzGet5wOkcuj3MiZF7qhxxsdCD6XnEjqarfOVwBbUnAo0Zy4M8F9g1oEeETS9VT8vF
jXkquQznREG3yhH7LTMEFFRKejdBmglQZsDEql8ccPjfQTQktBb/NO3os+qjk+pO0ryQlD7F/jOO
eMk1cjFKmCzPr8lWkjFNJAAReoD6u3OG52mLJ+cRNNNiqMyPO2oGiVFmeHpsoUQ/puH74bpNp4iE
zIxKc0M0To+jxnP3dHGZQGqeFxOIx5Xbuk/NA3qLWzkmhCX2IazXYiePIZJEhKUprxDpglfUVCRE
2GjTGYcfd/EIfzTmwWFK43FhFSJZrMW0FaaOk/3ZQUtXg7AQY1aP4jhy/MW5c6Yqnhe2JdjniwnM
ET+CRHq07wDmf45GcpFwVcrN9w0qWfILKJYYmY0tMrPbLNz5XA+9FIkDtObboW033tAlje8JmrbO
so8IkuzfnO2LPYqCILDGWLWXwSiyxpe9LWxH+tbiJGRGaCrZTf1wZwT6DBaY1MGoRWZ++HUqiTmJ
78aDb8khDNZEXwDSfsM5mnCtU8m6peiKqmzF7R/HpbfU6shiDOjaWW9/lMb/SGU7sGzxkSzoA6UL
tPDFXg6dH+b6yM+x31pLHS50vs6adlzMuNxLRhGGBAW7plUStyu/sLoMMCj0qf24dQYlLapst1xG
962KrobsU2JHHlpGl6uETxPHTbFZbi4GdVigWKVd1jVwhC2oj89aMDq2/qCbt9RCv9iAU7hnywKV
gFgqBytErYi9OiK9kOvYdv9Pqg2IxRJy/Vnk9mcXGiHmDu9404lhxQUxXj2z3sngHftl4JzcbIs/
7vbJU7Z60Ka5DdaNgKA06Oc56NjoP6YOf8+0/fJhtWJM0BaFk/5n7IkFB1BMZGfID7lDigVsNXLJ
4MYCD6xf+kP783IEpKQRxITK2eOS4JTbr+qC3IhALNZBxGyKwrN9tBkhDC0p0lo79Slu8wslnIFj
IO9ftbkxSLQOjpzTTLRhK+2MZ4bXtymhDR9T3+oaw4zwaY8uhKBCap4IBbCP5l76Gawab9ZFew9x
oVcPrms/41/Zd+OcGvQ9L98yunQ+DrP6L0rrMl3ok5m+Hdy8VvFtX+IR0KfbHw7FGfWuG0fpXiv0
iJajVLvt3tyUbK8gTTDrvhb/mN3UCKQmwnR/Ro02DZHm6eYhYE7r9+nWeiRde3+1CnTqBrbKhWNy
ejKnG6kfWHzzws0s9goYe9VY6U77IeohvMQBcOSaj0OBlvMxfDGRoFXsTGbqWvMDflQUHD8wb2B1
7cxA3/M0PGlVWY3Wyg8WapNfu1Tls+/UodmeFKVJqgo0lIUkoOsZofF5wsVhF1Tmgjz74ADmYMfb
yinpXTQjuO5qAC70j1X5NenxrNetXgPrTOx01hB4omV97vcrZFC10WwIUbsG6N0COGbFGrjT2Wxj
QTvi2FXAcrWuS15LKfKlxeb4IRhJ5KUcpUhQVqco5ThrS82uLWeIUomY8f4IcVQn/s47LSrYnwUA
z6qsa6JSP31gjKHZmfi2aGiKKiw7aamaarDyCM+bCaXOWO0Cke6IhZf2fyAMh7mM3ZqJ+QiXfgUn
CQdNVEZQhbTojIb0UGG8gjUPC8Nih6bRoUFNZswQUsLfi/s9UUaT6Gx+E9+w79mCVPhNX/dDT+ES
OeMB1BopbbT76vzKq8rJjg6bhV143EDXS54EQMY3Z9xXu0RHqp2nVvq8qLp6JwqNbjCvlAVnPBsS
YAUzMepRROp8wDuc3boWeD20qAqUJ+Tt3b2wF7UXQjuxf4mQQpun0bSjbwSSW0xjxN0e1AIxN7db
mqZOdtoIzuYvAKY1pxRKQRK3uG2+2FGkqnsxfhvbJCwlv52XvN3L1JCSRl4Qm3MDFFVzVIBK5fA+
FlFya9zg9QTK01Xvv9Abs14P+8+AKo8r+aq474LRMgH5LCS/wApAJJ3cl6UhWH7iiu7YUj9tbkmB
iozdO3ia4NAxaaFxEE1Yq/3+YyxY8tm7iSvWDPhm0AgB6bYw7b5eb9/zzT2+JUneJM6Ul3CPev2v
dgR539RoKP5zyjxpykPWE918Xh8ws0m+opJLTloNeNH6tYUhEIxXq8BDbHV6sOSPBlRuB80Aiz+x
zeG/yB1fHR1VxcBAIrQHOvgVLbwcSoAB0W7kasNf6NfdgCbQ4xocdFU38ftDG5HaNmxL+EyaUV/s
a/GyWWCFLXcEfklQ9iaOi7kK5s2t+SrN3ikS3HPVShRULGR1giiIQqgGdX7wBhzwUW0xSVFEHo9A
DiQiF7rEE0fthYujyXfDhnFv2aONFTdSn2q1XLW7+2QLHj9TyHPMbOKPpYUVRDGmmX8e9xzofvxF
LFs+k0BiiLK0D0iFq/BFu/LlI72jhQWLT0kVEglN4MpOR1WDGd3KcJ5ZEZJHEmqB5+Q8yBG3LuVx
5/9CzrSVGCVQo3u7M9QapKgwUjfOfuCeY8dirNOljPBgS0c4/U/sxsB2OYlKIAXQLxhzdyY4GROH
qXKitTybS0diZQTP45icUZU07qGsWawlXQxFC+onsq5KM3nmSVftGYqoiMpwYJIUC0xm3yvV8pdV
V/lugqjaQZ614MVLNXiCdU+jJmUhPMe7/OHJ5UKebqgIekdq2lZKZn5TJ1hIAMrt0apDatXf8MlW
Qv1kkxgyq8+Kqgn+jDDYoZVJXqRqN5Kw7oYR8y+fJJ8M0sU8V3E6agbInB98BDpR3ZS0jVndoy+T
sA+H9SJkaXmGm62G/ND2x+2X3EfX4e7Z0KIjn+jXwU2H53ySBxagxpK4eBoxL2YrK+DqbrSd3SDx
/w6rmpScicZVHRzBNuN/JskAEvPTkA5VvmWpMi0fynjl1d5hood0bXYcC9PNVZaQdCXN26hYTEW+
L9y9+Xwgk2cuzTPqSjS+sf2yLm7+ugjljzCEakteE5T9QaYTk2liRpF/vMXK51Fzq2PPHEx0firW
8+0QxB6RWEgvD/vjtdIlDZzGQscrMlSwipMvU1kLb/5SWlZeF8llpr57tO6ycfH9dVzzkY/1ixab
GQGSmqoiT/oCLSOpcCA5dE6XRLmQ1bhhekkSF9HclpYPW0om+HG6kCV8S6kYLtjz0VLp+NCBVv42
mSeHNZEkIUPk/wGChGQeFCQR32ktunGEbXYy0fQsMunTbe4pHmuv2EVtCAft+tisd4d2AQjbiYTh
YVRp/0WifMJvpZjSINwmmQxZNyYunfcLGp/kO4EDerI/N7lYGOJ2fLuWE227DUIl09Ce/aEeNGOB
HstOxNC7ngJ45gSLMcJa4qlafOn0vwU4bT+dOIYskMKHleycVAwBGwyOiK/xnelB2sJjTH7le58a
PGVYI7sbnbroAopUuYnxP856MPFt7hIsA10Do2uOrxb1PFxHyhSvzZfT0vNAFZ2eb85J9quBNFDt
Sim2CrLqDH1/wQzPbRfcvCxavUwH9vHgdjnS8mWYToXYHWRyPDOjQ7O2Vbw9q/4IVmKoqPy8Dsz7
EXbYXS2APN5Z8uzDiT/rYXKDJNXHwIspmNyDFrbIq81wqJxlpR256PXbu+4OHgP13nPcKa9fEyj0
9sf7nrBfuEDhqf1KHkCyfC7cvPxa1G3KdexNBiZm49xOUnjbSP/JSUpa4Lyh8e10w9rHYiSGmdrG
1rAzvOdy2SyQBPBSc5PKzDvds3gYvPfYDOHYOVFTskT1xYPevWRoD7hxPudeU7MtYIuyCv90pg4t
IGY1Rq1VAot+GWja4e4O3d0SQnvqxQgliXqr/5Z0AEzGotwSYy5t8wd68g+9ACcDvCmBM51pHfVS
H23FI4ccPAtHN1atpM0JD6jqGzTr1vsPkXpmXqniDa+9AAGDIwXBPzILbAnQX3AarXkZFe+GcfFQ
wqrf2SnRvXeiqL5EtISiM7fnpmOPNGuFwFwGik/zgSUQ82m0jPywrbKIeNBAz9fX0tc2KnCeG3wL
uydr8NanX2mlqTmilbxVL0LdPfwuAEggrhLMg2t4lX6zgl+0QPTnPkPie42wi6Uzyh4Ffr0/O/qf
m+TqL7jayD8iHH6VemJsIBD+czVJarka+GUNmSHNz96pAVoJJUUXQusmiri0NVa3ZrzS2mGbupPy
awgJtvqYLlCl01y5LtEHSG+p7aYL2ggD0iabVZjiuIWwyh+QoCpyhEYEL20pEOSG2C66XUW2LfAi
nhPQjM0gRLumXVJLFRYKMySEE4IM+Sq/6s33p6vv1Oaa8oDZo+TQ/wWeDQwf1MOzBOD+QfuffUqG
39CeUhLKVHTdJ/YoEW32+x+AXwzAJSMScwt4n+8m8oWNjtuYfFVItMaxIQMBknFzLkSYV49O8sR7
gI2v8NhvSNT1S3C6Jp7dm5yCPynCdpBWeZ+f2XeRGm77EBPntQlBzPE1glVLGAVtvJfP5PiVhlya
5YXgWpG3Py5wR0zVWxDZR8rvrHUQLG07/yfGYugu7nWXDK1AR1Ut3ZNYOt7Z1Db2OyfOd2G6GyPL
0bhLoGf746xxFivuGH3AuPOs8DA+a4OSZTOL1MckFFU6gQ5TLyeU8bUkSB1HQaz1RE6GACi3Xg8J
Y/WsoPHaBevNE818hRZN26pNLeJh5fUhXHcrWqLCnX4cM88UdBmjDhUhYfaahwwJRwYecmUaZ/Xd
QSl/3O8OwtWItqLqbLe1Ibila+AX8mxVHQWtZELzugWE9eMPkssDbj2mrVBCpYecvKMACaAzd8Py
srZLPTcyjKb+PXTFUE+Lz1deZbmyHW4L00sVzDn2Zc7tRDEQP+Gvj4p6DVDHGaQp7Ovt2A8iAz8I
2kOl1jTJHFXRKt9DetZSSCnpA83I+2xyH36vNz8oOQjObnRNbR55CPVT6xwqSRHmYKhWosbyMbEP
MezeQhHQsEPEFtZrSe54rw1gQLbQHmDadrbUCzc62GQhw+1eQr8ctJWvSiJuBnjazUQkUMkkjjWB
0DOfxVlgDgI/8ebu6QaGL23l+rqnJzt7guXwgjLzU9skXR0EClA0yl1Upo6+bpXSaZX54jtDZ4dk
h6oJo9VliV9vLnf9J4exJ8GPI3cIAW2kaBLvWdgM5lnLf/2W8wfLsBMFD9zb7patM6s9AOKoQGcc
rliw52eWu/heg5z6TpDf+Jkpn2maUEH2MhstXWBoSv2qJXBCzG6hDVQUwpOrs18Kr+SJADS6h5WQ
t1w/Vmt8SGLnxkPe1+eXOg27SNUlQrXVXDqi98rc9bp8Ud8EAD8GawZ9I75xOaYasZGnDjLXwphX
bcF9v2jHy/M8sJsPNYLt2M7KpGCodtET39GRHBdfyctRfbrzeomN/2Upxvqpo428zWpf5/IkBayM
BIWo7mCamDoKZe6HZHJ7h8yK6WJHFaDBSV9h7WB6R4rj8MqBOkVQ+QUmL0idl8Ei1yqxCBjrcDVR
mHELDlKKHQhdO4JWuaCeQAFD0clMWYIBu8wypnaI+XGS+9uBYTyZoyL2o92ejtLaH0pKSDhhBJfN
7SwZ/Q300khmAiwwvZxqmpNn9yZiRS/A7MdWBFaAcj0vnQIhDoxp8wW7DHfClJkdibFBYaNmT4ZJ
7CLdH6j6P7gcudJr+nR7bMkaYiRQu9ygPwplilVXZjFmvWOlwdqIvPg6hX9jXaMho7Rd2RGL5wP/
1URqFOSWnVMEonhwyD/NJbCEBPehiJVYgilYomRvsgEBSg6Tt/huhfGHs/mDJ+NuZWlRK2zmp6ZH
tOa6OVF2jwQDBykHtG4QYfvLiaocQLUuwSDbbIsd4U7SIRA2EYHRJdesAzzlJLhgC3jIm0AT+yvb
nTNuORygqiq5Frjr8cnonEsqad2gHxg2xDF4hUVSxt7XEi9Usvhqj3zVpOXrN6aH6qLUt6CeFOcH
MRqUFQMs/3oLth4xrcCs5Vdxp/ks3negMsXEm9JHQLBoqTbgftYEgGQMGQpagZ0PVyGSvHmzU+j+
T0wSj6CymfRdZvNvY7vW6dL8fFy8nl9Iur3vN4iQQLojIlL/B6/qWqqQdNWj6pNXXsz4UExFwYYa
c3CE5OgBmIap2w4WiLVimJ0wtFmaD0oixkdz4tps2oBKVfohCAt1kdvbvDSTDV9n+y8bn8cLm6ol
pRRl4MIY2T/jqvpfO0Tg9LNN4Of7ivTFkszEf7hde2tTc9aTiGCdhpqITVCR4sMCX21pFchv6SHK
OdN9FEGbTb+dzNlQGzCbwb/gf0hm0UUrhB4EwsPlL9zmpDQAkeRQQSlXNqXaj1IU+Bj1IqePbXFI
wbgI5RMAIBSx0soTQLw6BS2xlO8ajjLfKWzSem7ASz0U0+PF5e9A8lAc6kzCxxOqRSPG6mgK54nM
iH0enqVADkxVC6widUczMKYKCXe7NJ2Mi3PaJGKajhvNdoR5I7hnnxapOrptFXlE5jL680z+rddI
CjRbQXl54qPN81C+hjSo2iLnwtoD2pb0bzQOhCvaIxN/iT2pju4gAu5l3wyO73Q3rbHrPoKJUQqA
4vrzNU5wtvgxW6qQyDKyZKz6pEm16VQMFiYoX1CMSr8cLR3X7UDkiliWKHMgTf7pS/V2BnuYqFDr
cefnOd5Sh/Dp9xxrO+qcTaZWh+jcK/2fjDAvGQNfOhI15O9auPHTkso6z3kHtz+2Gdm+EkJ8UkMn
GYz0ucR3K6CaUfdKJDbebC0EtuEpURK/kPmoRvHCJu2FD5I2V3AH85wXHiCyjZdNwI2XGdDfPzU1
bf40BeQOsPP7yT3ebjZ0ptrbJxviMSW5kzzSn7PXJyKcyFqE4crSxuozZ8peOaLKgptuvNQEMMQv
MUT6bmvqZ0x1jT4h0ASpZD2tnoQwq8sptMfZFHpBe/7NWR+E7xmL7sKAC5zOtFTYd12zx2jP3BQ9
9W+uys1CznuJKjkdNaMvE7ZKfYuG7fq3AufJ1dUeIa0yDFF1rXkqEw==
`protect end_protected

