

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dpj1rsbRiC2XtvMMkZeaWceey8TRzfvuZghjsYUFfvEbx0wxaUtNO2KtH3hQvHr5R05ZRpFvbxnS
y9eflHJ+fw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RxF4+BsurVIN9R6VPOZY6IjRgF7yOLOJFH+DEaCvilnRUUfGXWquiAJNpzEAXSnsWuptbwUxy5M0
I2FA4+Rh4icthIWWJqsNOFS1K2ZEpNoHe2hVsMzmtRpnsPL9VGvgfvA4do7AYV7YhTUgoQfClGAQ
vFYxy/RbXBzM3PrDcTk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OvIp9LkjFoctqOSaxZyP7bYL7KElD3vYsFbzOXm+yqBzueGP4aoe0+732BJK3cSRYLmSREwKo0o0
Rv3hIBpxf0Y7nOdTTISL4pJ3qn/Q9Div9rDMzGaVxIOMLNLxqjT1ZbqCGU0LBxVzmDxHhBalP4V2
XUBBBCK3eeYn9YA+pujel3BBQ67ibuZRmgjKTwyT9B3SaGu2w8ce0O/YfSF/l+ncmV9cvUhjGdBV
Dsus1J4qhNTtraXR3S8daDpX289UCjsNh8krOgCnmBNlKeEFeTxbhmhnNPIAjDgfW1fdIgrmAH+S
tzDecIht4fghpU24F+FmCjpRFfArF8+d7uvxlA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4ZEqShxRoOQpy+XtDUXlHHAe5v38IR2wWpAtAq2KeZ3f4UCuk5LQw2Oc5c9xFXi1a9SsCAzYO6Rg
6iBcvyh5jboOYApBCjz/4VZfMAndhqby+l7lpAzkB6TqAqvqUfdVhSRn9DQMcQZ2fMALj61IBeLk
rnvtNe9XfB9vaA3zmlE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CxLbTp2UMBa44c/UwixvnmtRjPsy2Xb+fkOsP/coXETbFAb6XdUuKlopddrCIslByXBY8SiCzN9B
XnnZENqObWvYgo2VDZVlPu9SL8ZNuOrh2v/bJ7ztAhTSojfY2dBi8ojKva7J9JwGsRtKubJGASjY
RHw8CGw4rdc0A5dMEVmmoAymqmzBjExIxX3UWjtVz457DADxQ6UUgPgr7ysxQXkHN2eTr8eKtbK1
R8VALM11jq0MxZUpiiq5xDX4POkxGrs4QQL6Repo1WUK5V648ZRUZDaWyRJbcIm/J5ref1gzTZWX
h3koqZ0X3HGeO0DTx9nnC43UDVfA3fgk+YpVGw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33472)
`protect data_block
YgMJ9/ydIPotem2RPuFweHMuIc6gCpd9Bwlw8SA/shoZHp/9LWKXbXN8lSJ+6K8c3zvtQFoYcVHQ
OrBchqSqiQ1MReXx4iVFlxy2YQhl3eNOhRMjEEMTP12e3eMWBsripDwH2gwI7Dtaxlde595GKfCh
Xkgb+C/954SZDcv0VY9fKnpRYLF6kNW8aomq+rGeevLa6TAQjGX9EchAzHU3JFOoBIDEdwL+/adb
5DrCSM0rRwIZLlwvouLhxAihgYONZ1ip88f9YNVAmdnvEPwjUmmRt1WrdA6fUEN3hSC4tJwIkP25
7nR7dE88nSj+kztjsm/zkrCTb7in+Mc+ED1VQ35wq/HnabwVqudaFB9aftGYhyG+hoWdhBLPeFQu
+bc/6cIa4Rdp7FsNAGpgu+vSD7e7vq1gpO14d2H1aVQu6z7+DuOauNx8elznTlDuKmx0VRclOo9i
U3P9mjVVxHBKg3kBklWm09zDqKcVD5wjkTOTIn0NtIGgkMiPjtsRvPYuTFtMiIVuM88ydOS1xE2O
lif9FTixlBMkSItlJepdqdrxwgBhWPXthBXm9azE3p4hA4RjWOm1KVjrGfxyfL4soa+A6bsRYE46
C42Ynyxbd6xcPJC28Ixdy21xATbsg8og9BLOTMWrC72rD/y+wfxzUbFZT+DD8amB/8WXa+WNhS2E
dIf3xIPyvRjSA1EHlu6wiw4plRbFwojEx6W6q/9EJNKpw9agxLXKhayFSYU+iSLFeHU8JRtdQ0+x
tas1aSHI3gqotwCgYseSZZVlk+v2IUnDzug88tro7+aHoqJbM5myDauzuyR6EzgbNBDcemkv/2ow
t3OQpv+C96WrBaPfHBzHFghyhmM1DX/U+u4NeUFvD/173bvyFFPeKLd1Vst+nzqdPOc0LmablLRW
uSOzfG3IR5YhjVxFbcrXd32lBhxv3ZI2PGd0brs3k8TVHoqe3prVTBStqkyXvXUSDNOLLi3P098S
id2iLO6JElH3MqxG5Z35wLGARjuIZQKTMO307wBLo9IOzlNt7nWkaG5sEFtGkbu53DEZ1pZyWarP
AjJSwdS3iLe8HvDVAcdTBCfqDHHN4lc+Hsx0uaBqB9d16veCer6HECkij12PHpbNIkhOuoCVIu7G
ZXrFdw1JeqNXN8SuPw5b33IppF6pEXZafFIg8YifJXWSrR6WiD2I03dXG546CRl7g3QL+4b+qa+p
53x2rxMl70r9SRuEJs4dbol53r3gar1E4SxlL5ecAkuq5xORYCupoHUgx66IlwyHc2ojdjQgOXu/
yvGR+gh+RUlvgYI0owandd2B8nWwOKfd1S13AtTU5bsADqoEdinDwzLt64P/cA0doFNcMYphbGO6
mXr7oRa/Eb3bqP42kgb0gE1D6zIiNb8D4WQ3Ifcdf30LyWSPdndnkZDCu1bGP4ja8YdmDrqiRhY8
mC/HMQMUmY5/uIbzDnSJbl6Sw5TlkkiufdcMFMaMduWKqfTTfnjEqFGJdJzYKIaCenc7zEGXkM3+
R37l+QuZ1bKiMvLIL1EkBEzXGpkoU+P2shDZ8vCXm33EjhpaA3aAgbGYrNZHZEjU2zuIjWp5xu3Z
cShHd3gbJPXa/JNiRTKrg9kvzVVWeJ3NywMOTz+gnXiDpxRZNsMPY1pw4F5PHcxZDAoeKX+EyYuv
I6MX2Akc9FSEsBQTFWhxHtzJLwxeNUXjp/RRVMk1b1SFiqdhCGZEuYZfhgJtXrO88WKcP4iZnPqr
Q2KqUwIAs9qLJLVY3MKYLb/AWRO+vhiAmxNZzBxAPcEzM+verVghCpLirrDk8GE2HLchDZj4glJf
y/WJ4MGEVjw4En68n4eecfhalKeVGQb1B/TP/fxfteKJpr8vJI8BaM2qrQuokpis15x+8hOfTvHw
G6ca+5ziJtH5SKSsNGCR5UxJVtrbcB9yLEUQRmy+YCR2hhnEGrNW31L1eJTrcgJfZkl+BLMgjum4
9fjlW2rnc7VH45ovs+vT8T/fdK4av4GqNENw3eSImixv5BsvawzQyG0mULl1uGGCPx/UGbVY+z8m
0vKhhjJk+5hICR9MxBYIo4J9tQjMv607nHS0QrijU1ia44txnl6xpkqukIFSe6vfchtb8k9RDusT
JIwMG6tQqnGylbB8TNK5FrKGlH8ATpZyy1nt81+221xqr7azxQH9bJt1KzwWZ3k2H/CCKMk/fWuU
yFQqcAPH0ffVbGnHhd7gWIRrkIdsnrm/hQtKaPTAkzsrqwD1DKYSoYahU7gsUpAVaV5hNAlqUCwD
SUVwmT2RR3yGcKuNVfALOiBZ01fJR2bp3Iv/7aRM1Jfw7kjUSFxtifSXgQDcuoCsdoqQz0yTUFYS
8lUJ3LSh3oGT10KoK561dPIrWQw4THNcxAjdGj4zweXPCbxiwbGnVHngWYJ1PBkgmGIa1q/nKUDx
SM38+pWqL0ovSSt9cB/xNpm7uelhg8NsiCIWxSrOKasdw1G80wVY7WZiX0XbWtQlv9Xqv/9M1AML
ClfgsuyquAoAE2LHLMyrPN8MnZ2tbXqRnITdxQr4IxM4xWiGdYfCFnlcLPSzEdU4ugG09dzKKu2T
Mka2Fv9au4XFE3eWq26RsKxi0eE/aVXHQ1d2hogU40E0xXRrNrs0OtvLR4pXGA/qcaldXiUXRkJs
vgKvmaaOpK5drBTAw9689JJGo1iY8f5qMTqdV35C7sHe4JvpZL/UsIdfVqbhYCZJqvZlPBczLT3C
5S01kBD5jKvDnZMeUCMeXWpYZu38Oe1b/7+Zkytv4AGahMIrYy/lM7VEDUZHr+SR6PZ3QRm7D1jy
c2bX03U8Bp8Lms/46aPo0rvWBo+9Rhwpn1X3dU/N95dMlVRQRXW6EeXLGg9pxk6L2f95/ehLpdKO
VPgPiMqOLAh0NBT5jqUPZjqcl686l12lcNlhZegLNA320QLc8baJ7FYKqo329u8e+gRpuaPCP3i+
bvLeEfgxggd5JvymAWEhw+G0zG1KSLb8IQP5psS1nnLDcXz1NBo6eX/CvMMtWq0aIQIyKVx1Dvuv
EYXxjwuXncpdLcBxPVhz+KzwWOyukBHUZE3IXPJKhuY+x3qtG1teL5PQ2HbpjPV8hKdmdzIMOwwp
O5RcnR5mHownDHz+O+PnpypmleOdT1llK6qqzmaAG1+7DtMf7k0NLkhsULZt1VDHUnaqLZ9Eqddz
HgJ8sXEAfeb4eeJCY4gz/furM+ygovV+dqsxGtzHnXeZdUvSZmiNdU5bw+aTNGKtKB4Dfc+h+U/g
CNYAF6iQOHBa6vZHLUimILfIv+1TkTSdqbYvGA/qQv3wB902s2IBirTxJ5kd468vAJl9P4s8nmQ7
NFp5jvM+vXrEBudaScWa1otcxTH4DQTPaChO3al46MK9Vn9NMJqhTnLjAFOS1MIb2v2PWJqP/Zsy
B4m5OC17PssPphVOegV4y5uBohHMVd5vzT7rdtJUTPSuVXqaYTJWp/+MJ05quOB+O28nMS0BEASL
jhHXouny3O8OgyBSCkXyYnK0FVX7SYvRfO9RqOank9izYEUy3GEwc2QMFO3x41W4vRjWKcVZ5P1J
006eowEs8BimMalHr7DdPsrvaczebmzsuubBomp6EvpzHrl+qKqnQwhu2HH9tmCJo7W3/WBkOzEn
squ6AUNtyIxnpxdzIx7KAqIbvYYUTH6zCYGpTQvP554/iEl63d0bXvVYtsrkxchin5wFLni9mTNA
CjEYz+CYA03JvLSG1evB7YmXdjyi6cObd6RuaeIOA2Ge4rkV4onqDPkhiR5JMGcLyTnCsU0/WVfc
O7CWB/2xAj9lj61YLgL5M++41lexIpBDp1qp7liSZPD8liHMdGJroUbWM/7GeRb800Pc1G1oKZ8P
eXAXFrrTYQ0q3numl4yLdnPpX4WPZkJtSkGc+HXueR7YBElILcAqubL03gL5fQtSV3TNqBcpytCs
ok7F4ZVtYfK0UHftS09oDXo8KkK8jYUvrjaL1uuSL/GtpzAahE1O77F86wyckL8DEMEL14hX4PQq
9TJQQrQZDu0bu3NxkFCRauY0/mKg1I1/diWYP2UkFCb4x7+xQZkaopHvKI3Cg+uK4ooye0y2/Vkg
08PsRAJbYO+9d0QfMeuQ1Rcsw6u+qqRsbr6QLq0pbEv52FbxrSz/C/1aBNLjqsRW+ntn2VPzjkge
T2qpRpNlEu4C6Cdl8A3YnJPBpNETgU5Zv+l1H+OmJr4gWDyRvnwzup2ojHm/1HDwVRlXoaD5Ed2E
zI7KXo8MYyt8TTH64+z0Eo91cWEo9gB9QX815vi1dI6JTJihjJTpBLqK8MFdxZB+JyA5XI/diWAH
z3PnGN3AZMTUd0B1Yp7PlHiMyAtSHaaZJYaqWdbfSHbhboVswUFd5qKvWVXEvEyFbi1nMs+fk82r
dtTSCxeT1WqUigDjOjJqj8LgkwAZh8jiN2o9gdxe3HEepb3CxEyCFOQZJR1ND0SmjdQNZqkdK56o
9j47Nolv7DhkfomFCXTYl+Ec4RQSOamh//vSkzS5d6BxXuD2L/Gi517LyGHJD42+jjPfHGHMGZiU
XeYum5nnMBwRuxwWyyQUtSEvSC4DFaadpSSwENaVhq5Sz2vIojHC5virduUNO6ihT/TSdTRGlKOU
K9msjlYYjm/FonTyn4/Kd4mLw/2PBiiyxOwxpKhE0/qmEDBjTkAZ5tcwJX2rMwIU2/uXJEH+XTHB
OlxMo1MlAh1DrZd3aTDrQDWeA/oedGygGOEdyFeunTdFGmOstKCENzyvB2bJjZe0EI7NbRvWaHbd
4Bwt716phX+nc3dk4FvcTHgHTUBnGl/4RBrKZ8WtUA+2HVl8g5svyKDLFgr9oCqVhRb5KvJQyEae
qyaUdfZw2vzaYLu30xdNH0aADHEG5T5yj8c1pHRZgFqLD3XxQB4aGzTFrj2UNJhvBYjR4xYZanmV
H5bZSFq1a4PqPvAzJheKAgX9WmHMrjeDNAb9wfAJUfSB5UbIx5UcPX97UVH8MDumyfhofWXrwfJW
jnC2rRP1M4jj50BOIsd5TwA7BfgxPJe4PghqHlSU032vpf2JW3MEFY3UDiIxZl/dQXenrC7zSgnW
QsDObZhrXiuAGY0AEXj1RqP2lKBpKum9So4ZwkT7g6I+TOTCRaNX3aO50f+0DFYZB62g2kV3R1TH
NMIbcQsnq9EkrnVXwjNMEQwoSkyA0JkThg+pFAX98Zq97c9xuqCnHvtjz0B02xb9Ao/xAkaM+diM
lOb7w3HxMvGK/OpHPD3SSsA9bLFOHSFqMNUwCHgptm8jt6M8Xicrh4IyY/AZ5RYACc+n1+8Uv9FW
Uj/l8tFFvVnpyv28I+mrsFFx7KOAZaCemlfEQISfsErWdyP5H9ktjeleseuPVHFUAAiB8hZsJPHO
uLH5D9AHLUPP/svPflqSzzENDO7wNEF8xAx1BVgkVX8ce0Semdsh1Q1GfWXwxn4mVxki3HXEeD6a
LzhtU6g/kYCtBV8SyIikoAl/IVBKZXsaZ7npjxKwwYmrq7sDgo0ja4ehi02Jx6Ca+KRvaILelYmT
M6ql9UzVus3wKctz4d8eoi57RQdkm2SnUi0CN79nF5hrEiUTf7ahdFOT9bI1Qolze3f8LBLioZVw
ILJbw6Q3GEIGzl+/APFkDdUHesOstloC2BrvwyoYw21TnikKAF0+FJ2NBuA3l+/DgS+Vrz+fM9qH
2ovPp17lQR6m/T1MRgMb8xs4VWD1rWdaak4YTAmYG3J6Ar1SByi9q9Q++Y+ASjVDkkh1dLDhMhjQ
heDuS1+TTPfrWuUmWX9wQRedra6b5b1kfmzMvDf9KPlhxWfKP20SUz6f32Y9gwgIHn+15ElFpOID
S1jg5Dj9lbi4zSkjFXDGM5HhmAjadBvaCM4FtR+r62tAMYx5+u38i9SRXBWONlJoGLgwIghWvR7H
LamxxFWvPHGe/l4jAy3Wl91LMQEjaSdUpJWkne3R1ygxWr8Y2KQxRDqcQ2Izbz6xQF35VD4Kt0NW
3oA4l6YEyL/5j95EtImYpgTgscYRRtB5D2fOnbrQRyCzJpEDNsJnJGJpM8cgrh0ZB7/jfrziPcj8
jit+Ysvjg5i+NzZ7OUeN4I4kQnmAkF0zAF/cFSAwA0eAUVgH+x1UQEb4PESKjnmQleYu6cCu5ad4
/FsQBW4JI3vbjwByq+UApgwEHNcvcN0dKWu8GqqfUrdZxzjfrUvMPpkDhIgjPCpw1aGmbAb7kvCx
kXagi+S4Aq4BQpEcTwozkX77/20d0xKwbtA7ptXYPlOZ+0LayfuJsLetZBkDT0qO/Yf+KxNUbxLM
/ghSz7/URe0Waz2li2m/zXAZIXiP9sZzGd3tsif+u5nRTif0chHtYrKC6DIrx+/3rnMZBgj7cFTW
rHGuLzr/TyyeWRM35lRAZXjM61I+PVpoF4NXby3Gtt2+WnwvzY9YnbP/tzu5umtD2p2sNea+5oxJ
gtjBOBKIRDxdbNY92KaFu66wwjf12usZAG3aOOpHpRUzJri3EVPaZFaIe1dwfnRcGT/D7EAdufFN
v2aLLZrrkuHlTFzSo+75jRoqP8z3mDnVH/o8zXUPQ+83KP9GiCf/EmWOTxEkI1LRJgkJVm8G/CyI
WUD6rPPDtFQ1htg+vWVIqmi11jP20Sjr2WL5/Y+zBq73v6tLPcigigPcTOltiBRHcAeb9HA778E2
Q3ucWFWx0c866O1LjOERIOkxK0MBFg2xK62RsSyIB5FBUOOwYSRwlg78yPPVfGcOn+/kUxdGDF1I
61csMmrNKuUs0Gsev6sMmy7D8EgavWXLPqPqXotx/XYrBqdhXMpECxz+JyBRNqobc9Axcxn4kql1
dMSyoWgRyjdMWYCrAp50FDacM3WIOSLA5U33Bl3HrIkzg7IEGSsq3FjHICaQir+LsLpv3T14BRlU
iiriZm+sbyJ3FFHez2dNKwr59dZG60r5rSUTM6YglMwFazPn9euKIoOD3KjyDFLfeDRJ6ucLMR6D
tO2aLzMyez0j8HK5Zrt9wbNkQhhIz/O739aq6/rM5nG5RYLqHOHejSMfc5xzxunK5NY5eJKa11AY
2LP81zXgab/T2fpb0EXmosBg9B9T3IVtG62TgAnWSLedX++/ADpilfmbHjMVqvuKJ9HOV0Gar4pH
y+EUuwtsBgmJxHiP/drXTNVSQXNv6nXAqFYGevCgvSmLW/34NRqHpIzDf1sikACkpNmA1S75Tzs/
oxTq2pAOg4V2mso9CmNhmwrHNBCdV2wnzF++x4kSGp2Qvaabc9G7KWTs1x3wk+CaEsCo0gawJRzJ
zpiT8prvSOfke7xtapBgfSoTjqmmAp9j0Z2t9liWUwEdbRL5sezBxM3MVtefoW0cjJCgWdKIsgiK
3G3kfhlNMO7ffMA0SSyGtXXHcnvJVfxECG16vXuBOC6VcSoi7NDhPl8/3RWWqm+9WvReIt53ijsC
bBq/Km6k0MkNeG8yv0qlkPnV/2pogHK4AcR5rMy7oNW0+RGtb9qFJxu3pCZoFn0Ef0wTShTzwzgx
/A6WPuLzB+Vjx3fOO6mNKaUWNyqcgrtQqZYnEizJ5ng/OorLwwTpCnrU2xrCfbOE2j4HYHIP+/mS
9Ua9KkihtnKnvGY5tsVraTgs9UxfENVAMWCzz0gdkvFjUvhinS7+l0qjQCHeOHzX/cpq6RkDIV8n
kFejdXdsLkYavLFyZn68pMMUkZO2IbW9g8BPb+5nbyBabH4950wyoqpA+Fp0LydKDdPHKDxtG+dw
Ntcw7EJv0OPE6aLK20EWHmxwRddvadSpNuaBBjd3Q0bJ8jq8YI0TOpwxzW/wIoKR0rECvNAOzBWI
34QGx1hzoxUIHHPn4m6eUOxQ4dHTp9b1JpZESJJiqwOTmbHo99Vd8ODIDE8l9TWBDbmwELjRG6LA
ssNnhDCRO2Nuzdy4Y5umP2qFS/Dd6eErJJJsH5JQOmUcMRQBqicczCY5d1tR5RZfvSYqtQuWkA81
GXYuxwQf/N3daSVVRHBNFTzdkMXM8eqcXtdpLIWuYxuuMtR3DvGTQ4TUK3NPqrbgrVs5EBB4ZrUz
gLETSzQAjHc2tygLaJk4zMVptWKHEoD2sNADZc+1haIIUVIPwWIuY+sOvHjSBuerth9u03MKBvMt
NMLVgnlC8utUNTDC2DA2ejIRr07I59dCuQsAie8O+6ivfPQIyVerIGPHlKGUOlEq/PttBSMWgrof
Up21bNzgkrMAxV7x52hlh8E9j3PnyktzOsouOZ02lUdOhn2j1Klu1ZKdQJJup1LqAhoNUrSxCNKh
9jNptTs8/ViWdtXHzPFrJISk2sVDjxXvYHCUsOMm1TzSnhHZ5YbjttqMLpHAwtoF9/PO5H1Qyc2z
Z72f/2NeesHuueSrbbWM7c1KJv2q8Ie5QhcHJBxFi02/KcxV8jau2cKuIcBmHlwAOzTdzp7jDRki
07SJX/t/qdx7IQkFO41X2pe7B8q80MOf2uswDxJVK5znfT7a2Rs4ezMPNt7JkNKirVmwuGEgNrk9
FO17X6KXrKlws5hXgQideiFoONRWcp/hZ8fGjmjj9BCcWdGkC3m3BzSMGuetazNpFvrVTm7SOQLQ
DZahfgJ/v9mtPx1IFh6aZlSBMjd/2jchpkXbVJFnbCZfidJ2dYb0b3OfHxhrubg6nTu1s6ubcqdb
UbVS3PHVykupzdFI46+JQzbabrVEQzvFEyHTKM3Qaq8DLKl0q5RlzxLoP08ddxyVxQvz6iUnMKZP
EiaLubheKYWh0LfA778RVRLsgc4JXNKAorFZPq9OPZVO8UDfiuR5nGZM8Qx9nzCLeQtZpNShgIp+
rn4XKkFFOeb8PJPY9UBWGpIQx22riLtYY98rJl2oOuDgr4O0FGQfwxGuibtxsxO+AI2ItK4t2Q8Z
9vkbL62hKDV1YQq/1JE8C4pkli0lq5LbrrBu1jBqlgNGGq4CJ0QAkziKi+9tPLxArMTDmCF9CXwN
8btKbR5GybXAjFn4eLeafWcQ9mr0KK+fVgYX1LmCEMb4p6dysdmGLBlIVlVgYSdE3ZQ7gIAbf8mL
UktmhLigfY975t/1KKAP6Fux+ieMOFo90aCoF+GeVrCxP4ZyddJsW6YT4O1BkxJwHw9rzlSRhl2f
aHMkfu9o5N62FTDlP3dtTKtbdg6GNJWvnfR6kn8+vvvylMJg9E9FxwX/cb2mbqMwKGTyxuSd/pgF
Npxt6BL8IybUV1LvixABH3SNsauQEd3V2KqUZdQALWam+99tioxSNVh0ietbN8uq2nlaiAxyCK6T
tcQnboxF9zH61pS47wFxSrn1FH/2yNvuEzsJ6Pq84/PMmmZYtI547zYOnsaQnnymRScbNSfGDya7
Ciul1GPZfx9p8H0vd3B2rSj2TGt6TbVxBVjjqTs/JleTR6eL5Ydx24po9bNyqnP4xnj2qRlfeOIy
uSmyuMuPR0y0cqzfGVt1R/CqHm3BTS9Jx5/dGFbV/+cCc4Za90Ek91Th5tZ6pgnw8unTaTEz8Ljv
ItUkHblICVjGcV4rmH7xxqwk1EsGXe1xfAd9S7Aem8fNIt06h963KZBdtu5MgxJX5tKPOSILd9ep
Brekt04E81BDG07hcgqPQKw16FmC70LqpLbKhUrrU/O17xHO01dQGvwu04jbfjyvaTLCkh3M9DsM
tPJrKEwZFN+Cv/xxpKpbR1Sy9mnN4TsmEn2+0iInOyEpQKnPYxFurxRsX4qfx08IfF2gZJmi/C+r
br176umt4JKHlTrJm9FuiQSCUHYRf9fEtUyPm+8teK62Zsa3rvaBbgpEjUBk0BezdxIyJoh5/ZK+
RZcYjd+P2s1SRePqAUQ0Tx9aZPU3s+BfEnsaBaNqWAHmI2DqReLO0LGLcUaZTrmhQbbekmTasPjt
jaZi+3J02Z666gsdi3QpkhZaM6XjVxGrj1oDxHn8qexS1zYUMX64HG0Z1LLoTKkx0Qjz6USFINbi
5DvaXkHvY0W3xvNnjMsOwOl3wvEk0bfWBJOIqXURmHDOEYKv4RgSsCQhA21x7MEQBbcZSSO4u1/F
PtM5gFdJv5CS0h9LNV9GmDrw6/x0M5ToQGqL4DniWBjmMchbHB94L7PdCaQXxIRFMxyRyH5OgSK4
2tAiuYh2EupFkMpK0IGad9/UqQls6PoUVcwp6KvMapGnARh5iauV8Lnm3uLp2kElFgt1GsFEYKJk
qEG/M7xlXWK7GrWa9ie9p236ooVb8rMpXjTgtf3r6NyY2xpMf1lA9i9sPHpSe9FecaNiE9td1E8J
0VWDzgnjykLxZSN3eTX/tTnbHU7XuqSc/uAMNFaMqOxhBGzVIq7WmftgMgS/+46G+isWLl/zwht4
zBRm6TFrW6fn5CE/ec9IJeCttkeIz+++Af0sL2kbo3Da8XRPGvck3yYBVPKd3Kj3e6pprivxsBm5
2QN5e8eVpVUG/s4T8R+uKmfVZkgX7Nj6Ff2RorWmewIeB3Qy2N3XieB5CsjPYVpwFAvjSxdCLyKm
DT9oB1IPQio2zE6P0FBaYdRhBs+eSpK6+utEidF+tLefpKDeBFaSMxcdnRhioh2z1PU6g+dRoaGJ
9USvDlsCpd0KgLhiPw+rkxwNkEqp1lbXR1YWG8q+rdpZslp9ApXGv2XZ4xV8m44akDccF3rxBn1D
gvfkOiQY/mJjxh4GiUqMGOLaRqO8TGt1dZWjvHkh6wJAJoJ7vPEwgsSFsM9BNlZcG1SL5H42QNZM
7A1ugoQJO0j+0Y2twJLbwWnN4x8T/WBQxEaZ2Ns+b9Q2izhwqWbPRX4Ed0yhD3w4BWpG61oekyAU
gsPJFdnd+YOkMjGhgOrYVxCgG7h1XdVCyP/ZsFmz7mJ6siblxgZOOFFO2qgRA80jQPn//NH63CcL
6uO4g1RFO0IPuomK8vKAOL5uPVCg/ZgYJxnMARTSdzbD6dlwjCQu5wNFq0CJ9SNEecuj7Cg4/8i6
JXkwUTcNEewv1o3TVJgr8yyU+ZsdMV7M33/B6gcF27L50UUbkK1TdGSo6aaIBL6LVMpLVX5jVfAB
l/mMB3TBFtCrCsVk9w5WYbeeFGP8f6y+zz34J4jaAEcXfEPuzrAqpB/92A6J2Ix2PwPwiY3kEj1j
j06Sg0Q/5epLW01pMeFGxtq00EQivbZzDhKyF5J9H6hN7A5jS8eShCrhLNmWxa2e6mJwnmm8g7hk
yxaEY8wkrs4Cjok632T1zkwUxZtkVQkdmG75tJ0EqMrW30PzS++fbddy+tK1x2cwUvHEXTBjYN/r
TeyQQAvAaSXmZvbDlIM+CQaf/TyNWPMcgpjMVJNTeui1JAktLij3E2sdLYM1XnHgvw1TNQh3Dlhx
Vz7kLEK+VV6hGjn7wCghLs4rDSX6ox1x5h8fEaNih3B6UGAuo4LsOfFMgfpmZFVIsBOCAlw1Q/Lg
SYaB17RUdhbh08tkF8FD/1K3CyOmlOHzP2HnL3DIOOAl7EBc8c3s7WbBM7jcWT4lkRY/cA5f3efV
i9hyeGtyr8Knwk4JkgKpW2LLqphwrbIPkSN2dKjVgZTplLOjjCIIOOo+fAcCAFQxtUl4sx787j+i
Q8mAco55cp4KoZVOBOwo9I4MT5xbrjevVNToV6nkEM1MxMt7B5R+ewZQyBhxmezHwIHzZn59iLxk
XiEvGZSdi97+7JPpW1qP/QCNEeyaYj9LwtyWIqyLPScaNNR15EK84BYh4SbGYQ4jetwzmQr/GP8Y
R6fwSGQSS2lw4CSSNbpmRktFmj83xk3z0bo7AK7YuhoC3n1WTf2VmzR8J6uFhE+vPA75GtHorbot
lhxn3dV0JDYBYtrWAxUcNt1hLOnDzIa59riCUa48AFtd+cgNu0kjnAZzGDfko8BRer7fQYwijidw
ILPXkzDFjPnDF7slXFQT95UWfn68pkNKjqclEWcBuDxVJcK7GHK13iMVHF0JLQivf9mK26DTea+c
UAbqpLnKByLYI0hjc/zPro/xtuJV87rIgsu5rsSFKpiCbg6TUIKJJmcp6biqMiqnzFS7fnGJvX+f
mW4XHG+kgkViB3SokiPSDSmZzRmJTRz4nTmLsn9Qy+BzTxsaUowfl/HPDSr4qKAgGAIa4S5JT2l8
dL7Zw1zZwxxok7vxQCXqMP4LfQ0ei4jTQzwGY1WLJC+lMLJT9bYelVNfON0cAdq/NUWqd/GsTiSY
2pi/51QH8ustPhOCCUvOqKrDgZH1i6Gldrfu3ZqPDotQa9hBtvGrkabDwN0YNROuYmm/+fZp9G0X
sgcuqCGKqeEqfufwJt6Fy6ZLTObTeO/mL2n4idA1SLSrKwZGuy0r/YKMCWBr6Zg8c1vVRG0UPtuA
PTZ2zsZ3jVrxSymnycQnQNaWpCH2dX2MfZ57y5YkPwc6iiNLmX0HLvoOZpngUTG+vO9VffSA0sm9
cdEhv9JqjxuFcg7S8t+FKyMp9e7CmiCMeowuxIe18um05htxphe+93tPJF9hVyhUHL+Ghrc8Zb7f
Q7gryrOvU4/gWTwGjnzMWBlX+CSxE22sfN5x461xbNUdiHobY1sgtjQR6j3newRbeWyS8tUqHkmk
VhP9C+fI4ftebWkLtFeqQuUC8GtkccsQnxRcNidityoLHMnfVSVRxnFnfCBEWIdg2Cv34/hro2Zk
Ctob2KyBm/nKPMxCfIXrTO9gcjRMUbRH15pVV3EkI7Wo6ooTYZ5p8k97uGo6FP+DZkKuBnDdPXAW
sOUhRZTM3qps5D4ipBeseorXgP8aLz/Y4vQzDT2RTUTkgoTf0r8aWBg30+L9eYoxlnzrIgJQcg79
zlHkosShQW+LcQwf0IEIMfRYnajAURTa7XUzhPSFTwcfK8yePMQQziQPmOu0wdqoiesATo3Kz5zf
6LM8dAE1G8xgdNFGxrgelXJuzccQh+GW9/3yjUhOOLBAf08QbZdworiDT3bYhTsLa8ZNBxQCUC1c
o99APK1UaBc+H5ON63MqvImsHyoUzS77gBQvSXcnH9Wzv2Kj+3G1VYxWFXvIGazkoaEvwKMi1tTz
dGwxMBPSYkSp5s8tVhejTddezfkSIknC3BCLT1oyQsgklEBLc1XszIsVz1TIMGWrlLBAVIJYjOo7
4SMu288/TBCPs3QvU8fzZpAGnmz+D7C9lZwsp6rA5raEnKQY6gAZQvxeTL55V2sWiNNsNlcPzoXH
mFJwIyuEKTPhi5ZdnXI8DdGhAPPeVBxA6KRLBttYGd9dAC8AoGho0nm0Q6o+lgCJufioogKxTI2l
FCv3pOjstnrJ1F6CWDtu877WK89R7pRIdw1J2xW7V6MH70nCVCNh7nSppmyj6mqhLuyxcu1dnccg
yrEy2N8g22J03hy4TiZ2d9CqBJ5YEpcL4bDIVNfbudDjBUCvPv0xzxiHyvuTe9wjTYCDUaq0A3Ui
I8rBFPACKsLEKE81ydeaTF/YlGm35/gR9r8bV4wiHgyBNWvnbMsYhMVjv+UKeSHxkW9jVKl2gNUq
wRq9vzuP8PdvWyZGlJZ/KHFZTZwOvCMR0i9kHMNS7GPZO23dztYMIvXOFfz1kGWaycpVCZb59JzG
2dXKaY5c+0Ys9k9YfXQAI5S/QVBZuqbJ6b9/D4CdPP8BPIOi5j4/TzfOas9oEfl13Woijt9+ArQw
soQKo3HSMJlysRFY+NkyXUgKnArX8NsL9Q9GDrezJRetC8D+46xMGVrKiAkPKXREQ6NR8c7xj3DP
hKTHrq4u/NE8IDQPbcg/qlj2v4Qeqhq+0B8RQ6n20HuA/DDyRiWbq0A01vRwQakv5yyPKdEFd58R
WAICRgo5hCeQxESQVNF51Fc8HxgkuiICzloZ62KlDNAWPHYNJ/LdfG+A5P16rCYhl3ts5NrK1DZB
lAYmIvnRL+5ujrOnQS9Fy7CjskGCJQvdMhIaOo5MIswIiRPYPmMc7FsLqRw6cZZS9kHAKLQOFeDi
6fau5Wp42dLgyxZSx/yoYB15gwX5RDHU6pBoSMNuwUpynaMhQlyUGzGybcO3QgeQTyJwaLE06FOA
feh2yaGYUycRNL19In0Fj0DXkzXVhBKL0cZXkm99oFQlQ/5YkMupH6CfpoNtAv4/g//9Vnap2M0Q
60THqS20BnqeKvhSeuqzJwbxqErc0ODp/xz4uuIH0RP781jbBKU0wAQ+C/KsCRycoG2DI2lVVnot
M8uvEMHz+wxRR6EwXuq+VLYwvcogjJoH5Hzu35CHF1UedtGKoBfzH2n1Y6jHEuktUOBy6Z6MhZ3x
XeOUOQs+HEr3Dhe4SpPO6MhpMynF6KN55v2JDa8vXN3S/WyO22n8HK77gYT2Ads80RHjcTVLuPPa
d4xX6lQXRY6d2XvnTMPtQZ9BbAqNwxp+Gna2KKUYrBuQrlQpzs7QMEyx9uA/UtQxi2FLCNVXTu2x
K+KsUEnzF//RyjlzS8CmfOAoZnsxOBcvf56JojRt7YTgoSfNx9v8807SFIi9IJHt/GQWLTnftyP0
JO/dkZ4dRaxHTBoDaX0ZPc5rdPHppDvJz3mKgGR8oTg6YUDiI1qfXRuiy2ajOmmRwPOWnSiS4ntZ
bCCBsx+Kr2Iq5f08OZYiG4wrq4c5sB6b/bEHBCRtfaWQ59AoyO1GT+1EXYdjcoWgy0G9ZaJY7S3X
Lqj8LRZoNg7HgHUMG3qsTci7IOBFMJ/ROI4dwxZ9VWjloE34O2kwZtv6mfXTA3Jrkp5sfEY20/Mc
vSq5ky1rV9ivIQCRcRUoEiFadU7houco/wrqLytLUmhi4Mpq/wx/aPTzhzDKbnZ2FyvVCOibHnby
HkTZNbK2KIxSzY7N7DQ64Z1AUEL9dSQBc/7HXrsfUdvrvh3KrAA8ypnDrXsdvcidPNP4/BsarGod
eRVHFAMk/OoUiRVRntZrSMQnYy47JXgW0qJjRMlLIZ7F+V/zy9uP+ts8vLTbrGGQ2vFtMCDJ5vuT
N1nQNa3KOMO7MC3blTSm9oR0M5hREDPc23EMb1fvAT4MUgT5znOOD/kmCDhAUYL1E8xOTM/1Zrey
QUl3ZfCRPzFWsXQCzOuIHvmigXXd2lU8m7YyXDvGCcZ9Df+NEM5d6ghtUNq5C+lYVz1auVvUS8wX
D1BpB+GKWngckar20EvNNs2xTlRFTQjIVt6E1lh7TrX+6gC4GEGMEy43sGR1nigy6KNdRGCFCb1R
cZIvnvhYYMawCP7HnvBtzaCF2BsD1CBN/537Iz8c3A918zQqbGt6qEFpMqpewEnoPTFZ5EO9kYEz
m982RbdtcShYU7sRH/Q+H2ei5n4z8qjcPhTPCOqXQQ9TobDDkh3I0jsjXASTHEfucd0XtHmOM2gO
IRiiYawbnr9E0hcRX4ZujqJKrA5Shapr1Cdmizqt+ehnIaSibGK4J59ufwwgYLhpzN19I8qb2TJM
NGtp3381aJkERT06dTR1coZMgg7Ayki5MAS2zvwe/VL5fucG9AryA8PlwAjsU5b5mtA8Xxi/9RkW
3WgxIKEItDu3rioMUIMKtU+FSVSiD7L5MmnfNEjDUwiiKVNN/lZIu8TZw2PepzmhrFD5/AbOlvjR
mwKK75eihm3gJlnTssCY+tQjicRrz52J2dogqSb3yV/nZ+GCZ71gdpWNDzes4COXQ4/BBhQPJ46F
CTqz+TLDxto6ZZFc9S28ZBs+NXcWfOdUP0OVcvj9UalYy7lLra3qTPxJwQUe1JyjMz/kAyaoHS2H
kkBD31w7QyBbna4ywK88GsWsGFk8bIGSGhpxk91Qf/svsLSLzWIlBNUHADQqnFpC6txAm8y+Em7J
qLa9eOURawZs5iG1pFSCXoRMWCX6RzASmEyEMsSnaIJBMVCYLh9ywYGLg/jCg0gURZXIKNSbSRqC
PC1OhfLR2XxPx4cBF0NH8r8YVsc/o8wCkdMUwh3k7SXOIYOxlcHNtxUsLnDdBdOOkWsWf4eH6n4g
wm2hlAApFgYi+NrL0MUlgbUTRAgxUI3xSIttVYeLWrYKOslH1QvBYelOhbTSCdUGxDiGhOJF5/Sy
lLbOI9YtCfzKijMjnFaDk4eHbSe/buVz5SCoaz27WPnq6J/KBYZDnUj1ZWfS1qgqSLMVARM+RWtr
clsvnrVk+qTaB707e5NYuedktBaGt7fELK7ILPqIonkuZZ/lSeqPBUqof2cowYS+bhdFxaVkDAcW
rCwaNXfaUMdrYShZZ5kb8MJyA0ceVlXn+7tRqMDrRs1mJRoP95WxrmduXbAl6ZbaXBa1B2c4GibQ
vgwLRzaw/UL83C4efJLcsCAdei/O+/9lcI4nb6QwoQz8ZM1ptyL4aIlxE2HreteHyt1RNZ874Pmj
GGSoxrBkYm4kKzjeb+52nMgqkI9YBTsZH2tnyui/Ovw02vznGIi8pZABGflNXMPVSIMNvUjmaQot
FjlQObzEY4SsNk0ifa2pzwk83IJnGCDA22gZXzX1TSaQ7x9Ps5DTj4W/+7VCj2SrCI4RgSR0Y+VK
XnofOh4fDA0i510IJYvnUz1bzf/ZhNmedAk0YteXBHvYXxmmLcJpvfMMyfr7mHDJKPI9nAvdRvej
hx4Hka2MjNPGIEcxJ67lU9ToQYg5gvj2/MBXnACCQc0qM4K8bfAr++e0aj5vbSUFrz4HZI0JCxa9
Ds8LpMyYWRO5bUUtiJye6qnLDe9T3uxMd6P5v/nNt2YPmtaiS/IuDOMErRrJNEzzkxThL3r/3F0X
CXlAZ2vbsquElAROFG8iVVrWoLUa0WjqUNTx0OHtFmZ85OH/AWtEbxVxph/oLp4b84Seqr1LUXH8
8VBrLjy4oSRt2LSlQ6j6Yxw84QrWtKl1xaR4GipyaEuifYHz8FmOItwy8avdPYuPDcoN2y8W14/8
WtrVx9IIqAZaMUmtVlkihsfkk26S/dbScoWVhpWrMJp70h3qymior1pKGc9XMYqZBsyaopm/rprJ
YZjgVFhBLHkmXwmGg8aGZkQHOS3xjw4ajORRKyUBGZZK0mZ2Q+bWoTPWz8jp1vq3/3HlWn+d3rqF
KYVQxrGTO7p0/y76bkTPk9AAzLkGa8GjQZpOAdSDzsuQQI5x/mNnIt9JWlHBW8Rrlhu4sZK759S9
mIRYE7vyR0ucBHFJ1Au9I5XbGbI+d8fSFmPZm3NQfa3MC0JllQTlj80cGmavXLUgB9+pV3Iduz3a
adxL3lRVLwfRQdWn3F9C5CBXdn0DXvdZSPSwRh6sIGcJkHam3kLunLDhTWZ+/1H24zfa4wYtpQ+c
oWGwmEX1l6f/dE7CiQsDB7cjKZaye5t+VGQ+ut22RnSRRd1Zhov3dHwHco7GBJv7acNS7MaUiccc
h+vN5omHI5spC5LOOjWeSm2EDUaCJ4Jv8ccSzb7sxS0Pm5r6f3ufdDB2jnCKhqDVR5zdwSvR4aPE
PgfIXyObuW8eJbFTvg9GcPv4w7Uvy2TQMcrOlwGkz1Ef7EhUce7KkAOs2tkEyk3Kdu8bU/qYsVGH
lyNfXry43pqkASH7eRqLXl5dUYn9aMJLPomvKSmdetKuErcKfJJCVj/GFzQo0pqMxZoPYWN+VyNh
iv8xXsNGQWpUK/qE0URwac56TcXJt2I9kydpqAZRborR6VBJn/3m8iWjuMFtf/qIgg/eK2if31AW
0Jf6Lvl7asP2e0mxWlUkjmq3WSwJ5XZjzIIXOo0aql84WKvSJfSwAl0Gxh/OeuKRERVXafDEYOTu
o16fMsfOoxTAC5pycfvxlDDgqCbTT6NAfJFyrGGMimEcpQ0NAMGTvBw638mRjMbBhn+KeQLF17aO
XN8/1b69xDbk7hUr0QOg2N0rI2l/+qkoqmaVv9tnFLh4Xr0YZMfdQ9al2mtIO+W1g4XExulPM/tu
RM+3s3Yx0fWjhsNcuiTTwEuoXN1CRKAjZAWwMwr9A/7g2hTCcQ2UjQJaGXkTxrX1p6qpIASbFxYk
yoKpDF8hqiHEfOFqCgMOljCJJ2b0A86mcOWRl+OHqAXq56UfQXpAdVYDX+mxlPaxC1Q/KevWXvKZ
Wv5tfFCwl+lJMadqy7PEXPeMMYMhEd9U/rJB1GGVqtxHrqM0MJqxDrqKoEW6VbRkrjWqOR7rZa1x
I3YVarBRQOShdMw5F6nqi4BDGWwwQq2X2CXNp88CO14xeB7UeFPbp+6AfsmNzilLJjbBxk1RdjrS
sq35oegLGaOPMi+A4nlQP2DMhlGy+ZXlrQOA0Xxj83k2tYIvOATm4E2whHUz5xzd+HnU9tosLwZm
pGBA9jipmEeCfa0n2nBkKWeMZQhYUKngepuCOixXMyCEocFuqvoh1n8eGMJMMttqWzDHP8CkGYA1
sOmzGcXvzYSSq3GVVJw9EV5TtTNFQ1toP6WGTc7uPr/vM7wflzl6HoTS+SGaZp+jDO9aozcnZDFf
PPk1Vjdro9DxxQhj12O7aafelsgIeQTCXti2yPaO8/uxAnOB1hHc02+ts9rdT/xiDtlroG80rEOS
t2rcO6pk559CNNOq53lLlyAAC+ZgEW8B//qUOenY/8NFKCjiOgt1PfMEGv8GOhH5T9ZWBBLnyXrq
AsEAXERAMmKeVdULkh3eiR6ZJPsL2UOI3qm0MHgp2PsIlZ9NL0pDIitM1fxdqS8/LO6Zr2HpxVkl
VUsoH2Uf/XBZuc6zhm6V6T+gDSYQnh0CQOJmdTAKmcIG8uWRRv285qxtQOawdDBo5OumuStFogi4
u8t7orUbw8MbPHiU2Ck2KNhgZuJi9nOzk5Qi/jOLltUEw5kUKI2RJUW3XQ/HCoJ9Q1IkvGNojyqe
gS6OTpTaaSIdRWw6SHO1T5X3NYH1uOKTnZBAwXd4TMFrL/uWjjIs/uOSUcgF0oWBzHnAOdXN6+mB
2epIuXXhdSjvEWxJhgbIDylm3524ijNbwcDRUbJ/5+95iASTKhX3be3JvrZ/sPbnu/30BSSzGvBK
KvrNjzMfblRpsZ+vcnNXs/2btGHEwsjQ3F8seWZOq8knaxMixaP+SOQItZNWaIJsMcX7YQGWFIBo
ht4qvERqxlTVnG6AQLKC5Ls+zqZzvd22lGz+s7UEIRGoPpLRXY0sQAtPEgw3+NGNP0kH228F68Kd
U3hO3lzE2ITh6/rs+POZJOx7EaUKnp0Y4zqim682ddrnv3NFAyBDVMannoqUsfqT5v8ifH7aRW7d
E2KwB6HHhN7PXV9m5PlqX46jmVHCcQYyLAftbUQqxun9KwCXH3fO+Rg0aozkT8SDRNeT+PsLPyTz
9zmu6XTObMLhFjZpkIcNgUovT6HjrduCy3WS9F8xMQEfyLNf4MnngIAJE45zmuQGmZgBA0poF/Q4
x2R1PfAobyMoDHy08SUg8biaBxuZN/hRVmMNCUS0ohsrot9aOg9Yg9nlrKh4ih5UQW8wVniyQjn5
VRG/B6OZ/2HNw+HLvMX+zgW577uaooWRxeh59mXINZKPV/GJR6mslo/3vvubCsy6DWuEYP4G3vb3
3jZplVp8P+pfPajC/3I72Y8KDV0wLERvUAc9EQxZtoThC7AbrLsrkBaqBzllBk1excOLPAPRm8qQ
UjjGaglwU6Av5e1e63XtB8WJreIPN+7T0SUIXXc9PNmmh/5uaTL5fgoQP4cam1Xgj00vSUO5ih/b
EUAq1c7O+cehBokIqkD6Ua17HJsD6eL6LeA9dSRkfa3nRdjVFtmpHo1diAokw8+GgatwzoUKIq01
qwjfkAdHQwkCZt0GyIVYaiqOBrk9/CiTgS0AaJfpB2gsMVic4nd70sUnQOK2LFFjGSyim/zRnt5e
GKAk8qCAciX6Zn5p+oXk/OUzEqeATPu3Kjvak+duhzljlFj4mx6j5IqQJlXU9a9GtnCmXPkF15wR
LMcBb9n4YvOrIxn5rZPqPoue+MVjVi4+xVmFZ01ynqTdW1wlZm6p/El6HKLfmTiuT6z4rVmfhglw
UyW7aiC/ROAUN+6QH98RCMPzTUMV0vWqU+HcT24HB3Serk0jgmorHLO0/QfM/KWjXgl6LXLQBj+h
TkwMXyP6rJgvDKZfeZl+ibLHywJJ7tf8Og8Zl3rt9MNwI/Q1EkcMNPq2eda3/B58AXe+Ebr5QkSV
SZmIb6YutrtC4KNbnuC4L2x5whlcIdQBd/ZIT7JwjbFXaNAxgyvtHU/MILABIbmOqoNGYjGJjBWI
DjiF3MlqxSpvfWaeZ0j4j+UAp25050qqcttPoKOAKCIdUUBYVeBOuuLnGnjninctgszaJIESOwSU
jDZDW4j8wH/wwSKJG6AHMZar+O9hRgKrwi7vsjcigaH1bVArpZEF2cVnxue9pBtzkcafgbQz29pO
16MhsgrPHB94xqqEHZZidHgW0Qp/tuymgHREPj9Ssa4T9KHPL2X0R/vB46YuygmiDyZV0gq9dKv/
+39HTxUSxxV/OfPgyxCE6Dm3kU8NbEHANeeWYPBUO6Ro1LLP/5+N9d2GThm6cYdOTNnBHf9SYguO
Drn6jrAA/deYMiDncqFXLzw2hFE2To3ExAK7/ecXMb3ddTbzYMKwC9QKqwncJhD2aWmv0r0TCNHB
RdLCB2HYTYVCqyeG9Z74ZXzT43z0hI5UoIlEqdf5e0+CPDTkI0yBNumnIMgHbomeF5iTogPGvARh
Ldmk7sVSfTK+0A93D8d/5l/s2BA1l/fEiiw1nPTziiuC0veUp9gjna+VUJ83/kmHp/vljbUuwBg/
B4b5Eh2/0rSkzXoQk3EZOErj8stgbOxdrR/UT1uw6cqWZBrETBxw+r5vWp+3Oduxr5aCUzb/fyLq
zKfX1dQpUv67Kg6Pv16ap+fWZMyZEvZEkfNY8X/erlPW09rmT5jgam9hFW91FWxu60lixGEeHvns
9M7b7DR71z/eCYpYCvxEOHK5w17nDXz6chs51e/PE696Dxo9/4QsW1vTMJ2AUhxVtYedfX8xPoXm
HdyQIaiBaM053JgVHv8TsdJtJJTVUEYw+wOZU3e7DjuuwAZ8gR3kcVw5n+8DcnfCdGzkBDX3g5p/
sZT6icLkokE6n/SXyfb3iUto8gl/o23R8kSBlkwJcuS9yknwHX6exWETWcVzb8ktzJ4jJBLt5NZP
zNJNE26ek++/jME66Cz0Ab4K39iq7QXSY4CNFVGAM7KnEGBNBsqajmiN2GH9Yjcgv1gAXsuhRLuA
AGSrjRKKZk+DrxlUq38H+o97iwhjLTPQq7XEr88Cax+8K3gxBuKHQvEe2eBQk+ePQ7BU7EBU3jrj
XYQDXcTdTp9Q1Q8BWzUAdDCMI2AnYcBNjBtxRtIdeDEcCwbmJWoUvseCJz5eLDhG2SUtaaUOJ2jE
sHa0Ndl1feazUXewypGTsLmd6VM7gOOVb8/z79TPt/J2tdsskyUExbgbVNQOkYsIySCA2mZ2sBbE
crWnkjUTgxrBpZMmdUAqw3YC3IBa6RD6SGkcLTilKEOhLa9blHu3F+XUgUJP+raBMi9Rq/0czacf
4aLTOC7cm+lWjsdufwd4NpHIlcwkGanNvmS8elpNrrrlH0ZdXiwYob0LpyyKAO8c/97lkS631cPw
z4hOv19TZoVuoYPXLameOkZdq+QkuTaKxLi0BxOC9f+0Wi4MV+3UgFSxEgOwnAarmeb9uCcGbKYq
VyO5Axy17B/v+iDkp1cN3zTFslDHgGpmcObnaC99zFTLuVYXp/Fds553Ht3PDqx0TQqIgIgpx+rr
mT5thZEKhMNhsTsREgvXaV2BMQrue5wswoT6zVJgIgsz80aI2nGGV1cbZPFk1A4KYDopfOQp5xlj
TlpmaWbInAggdYhItqJz96b6bxBm9khhCc50X8p1YwtZPHiDK0qQLZz31vXMwajMn83pgyE1oEyM
gobsE2zuNBHm6Ff5/AMWlBH9PZOrozz1jbTBZ9wkDiDOnbDo3k79AAbZ03eByOTyHmbkBRfF0Tt/
h2QlLlrwogKvTjwlWcn0dmEe3VqbJ2TyPUGWDpczj5dwVDgWRt9SiApCZwimOdDAUknZVqtaOcsp
N8NUhPc7AxJnAY9kP+E+yfB10BIV8EUj+Kn/GBJIlr+gJ7t82cmqjhkSPtja/I+muPxe8VV/yy6k
CYwosu9F140neHZYvjcp3M+g4qF6Ubr/EVhkiB+vZcGLxUJHIettli5K9CDI3rrp6j/aaEVZzAdu
wOeZeuScbsWSppkt+8hegUbKrlxs3PZVJjPnkfqwioajnVwZtxj9Rm1uAwkBcnruNqmVbNhB++51
As9OUXn+v1OT0rSQ9j7GvyNti8F7v8otPh8R+cGNhNXlgCqD0JilBtN6kBzaseKv6BRZY4948Ieb
TCx7q9bONr2oZViWBmbLqLULFiesGRXnt7wEF9J3GeGmSLtzHIGDpQHVOr3sogPnSXaT5mRmUexC
1GmUJjzkVvwbz+3wABRVSdZq4vVeIRoRhRbjADtlidguC7z90NMPbGIh1Qt+Yw1dn7hLzylY0Ffg
BVJTMR5FeBSuwTVgHK8iUAK8XDfwfiZu9zM+xMeEc8IPr2Sc7iPzB7ns5n63ix2Ni++BivEc3tLR
Qm9OkimROpeel4Qhonufd6fT47yGdF9+kmmPzaIR+kBBQ8fJiNASA/pQYJZp1OzbJ7T0b0BHhurF
emfMoG/8LwH3ylhjLttAzaXM+acg43t+OLMKleZprVwJXnRT4SVDws2kIlt+sXt4NWp/IGKzQInC
3HbWYDUWSW0STFLIxNhseCritMsQB8GoAV44efP0jxMwCjRYRd1PKNsFIyqpcWIzfNoZdHbksIaP
LL8OTuwr0S/lfLmQSsWg8RUkFeBapP8ztQAEcjLZswtZUO5Qy298xRKVFtwYOpyv+EmWuV+wdRc2
oTkZKxj2LkhFZDyG2911rUkHrs01CvK221/CIJGwXLhMJ8VZzKUZRC+3bDhJxL+C4XmQxDexMj34
HMR2NHH/F44UcosZAFcUn54XsqXgCAEIN5TIKSf9sQAUE7OCzMYx4Kb42WndV6n8DyqiYhZW/x5v
M4B/TMbUZXFObS/8cgDHaaQ2ldYc8jTDsTcC9InVk4XDlwBOtU3aYWlFqWPhbkDw3e7OxDGgpcJg
Ce3J+nyDplvHsBm37HADhsn96x/zDjCWN066u6/3xXQ/2U6VAHvSqHL1wMox1YXKFxxW7K9AI+ER
cx41z+/FMP76XpgmV8LBJWXbDakNnLCkmtp7kbwPcwUa1sYXZge2ZH4Pf3kIf4F1MVbEz/LnLxve
WXoUFd2figB1s0fQ21QhkT/oKoUGyUU0E/9F0Ble+pl3v3Zu6EepoTzINm98GLGacwBQFk9QOTHb
Zj70OAx9aqey8RDnI4sljvEMSkb3AP4jlw5JT6p3XUMPh6UKCX+oa+ZRHBfz6DMOgy+iscSK0hoh
2pHtpm1/xNZhHm923Zt9iDQFJCHEDEPOKYTP2t1l55Y0m5cldjWesDwSZs5GkcuyTZa6XkGPiWRj
XsVJocd3KBT2izIRhnqn3cMs/uBu2FKvFRK0YdrTgByMcp1o4lrErX9uZeel0UCVujrjMHuTW2B9
0WEAYBDjNPa91a7kJ4o1tAvDGWu/RLJtV5jQ9qLj++K5JITUpDN7i6Ua9OxLNIrL9A8JIisjDnmk
QNjGM562yyZ1DFU23RnvkWm9tgS+3VBwysMfD0ymnjbIxA2VjFIYMH3pVZsDQoc7JM7t8Hiolmwg
Ld6WsYIMPVM73UCC4QrMNPVRWEQi38bHS8oQ3QvccSaoVJIGPvh1BLDDZMN/iANj+nzkVP+l20o4
rhMsluQb+T4YUocxMX+HOSIIMwlm5ebpRWrbfYVa9AVjzqj/Oo9/NnyWUM9MXzV38PDmcw9fE3VB
fckdhwSfWJ93fNgqBOzucsWGVkEkpXYUhUDQb7FvPyeG/e+wJrVV54qrdTe6PdJKa/vgQ6uKMT36
ncVqLWetvaCvf/As0pZ+A/gKMGHhwGmTXfecyZIE01bjM1AP5qJfTdD/Bz9HGP2icg/PlU9hI3wG
UcbFifza02OCg9KwPNIAAw6+hm7XisGY+itfMZX1qTfWVCZ2wxGAjGSHanvIJi1osTc45tascSkg
XrO7+GHsQY7XsMWsj/LjTGL+hT1fKZ+fqNVxY9h+INXr2L6jaoYI0FZndo5R5J7fjmuZEnMJJ/4Q
rYPmRGkY1PfiD3Pq9WCUeZS51vT4fcxU5efMiUtf/kwgsYJQjGOxHEa8FOM8EWy5tXdjMwlyhtgp
/oMYJrffcYO1Ifuk3ZbwKN1Qon8LkISTQ3nFbROmtSVab9t0/WG+4gSnohYm4q+L0nlyx9W7Yb3w
Rjt6TKZx1myil0R5+lD71X/tvNBpZT29bjKewnpzIC+7Br0oj9u47qdhXhtTQt4KUNY2UB8ZnsDS
sgYf/8Opq7pvZCl4WzYrajjcpvYd81im7leF6gZL7yAkQbQZcQ40+S+XgFsiwFat0gOkROc58VWa
F3NbCFTNStc5PFgmdO41rIo3OjJyhz4SuIyjW8U8+zVxQsMmFSpMsBNAkbHtdjS2HevCGGANCHRk
HoQy7ONvKy1hTlST/y6b0rw0zK4J6MdJLjK95Pmm2cB6sLpzwU8C2/UFgb6wcTsxTKl+HuMRPumc
kFF602T2Ooyg+j++wywnStMG69P46tdQbk/opW2x7/k/VadtirX7H03N4t4Gpqs7eEiKIun/nf30
27JtvNxkrG99ljt/sEZXlL+QHtStC/tMXNYu8VJSMUlhxJvNHFEqSZZnwrp/l6dPZtJFsZMgA1zr
3Fqp5ow98IVODBL8O5R42TIHF4Ps0/uLVxwxFWNey3uEJSx5JSkC1CFNn+bNWzKq4r4+F9WiDqH5
6VH28bqzz85Bc/rf5iKfTtpc3nOiVKUhI1wLYJLKmU5b/2bl+P7IOmkMvbMNJxmZCTwMtJBHKmYg
yrbd4POW9o514lbGu4NZ/6/LOJfAIyavJVrrN53TPcCwS4B6mbtX87Z6U8hVm4rCoYyw5THFcKIe
IAe/u2YmPViI2xGrUUuQwFYv+GV54dQiXgfumwul3Fn08JNi5UI3mV+3lKYwt5+GLIvgBra00jBt
u3s8/NcRtWNX83NXeJje3aFZ7/sptv3/E5CL3S7ttP2ntoaP+1jA6MVh4qvr8+iVpYWYCoxj3laX
B7udjUmHh2emM7AoGBaKYDSGJoYBZyukPaRuQ+sam1QF8H5ob7rPcYsLb0uURlhnj1lpLf5ffFGN
1n26DQbgKO8HRB3kyhjaKxR599dgyTCI1/TIruu/HvrcfomGcbEoA3tpTTtWy7wR0BfA/49sMvQs
3Ki/kSuppgLUcBjLwvABcGo4Y1ogz7nu40133UtCw/57IjDlgInLOVaODqHp4hQqpwIV2znIcAID
F62pjCpq0hjz/kgBFow14Wp1yyH4vFadOA7LH5mAd0d9tT2HHvHJjKd8LFQGtfhsHNZsCfuKXP7H
v15cIUuN+AXkiwlNvzn6ZHYripzAsJ2R/EOtJ3kZHDP7DJyKX2pwsrw42bjY9K94SRoRgo6EtdH1
bB7DV7uvf3YwMm7h4UoCMf1LIvXUqS1MCRoQkoBxbgFsrKmOdWEcDEzeaZylp9GkztQj5tGmKVgR
bRducXwqn4FZ00ZEthr8q7J7eWaiSO9DviYhhxG7VTTRwHBz1yE2IO8wWHS7gEUdfhWKh5oTeE3s
1WiOSbVlhj0N7/yi1lFwo7BM4Pyyv5c3WPRPNaSH46Wu004WNphHugdOf5n6W/hc+6Yz+c7s/ME+
ipt/a/pSn7B6DN0YVU1xo+T2u4L8Wdi8DWFLeWZw+zOCN2Ftlg2l7bxwwIkTPxq7j/DUzXwSuaSA
VpLRCHf1A1kvfMuJTbzWXvQR66/6IlujvnNnZiiry/YzkbJOz+qNgA3Jso5615KwAXjNZd0+oYDv
/nPJSfficNj2ahdXtccYHLG4E+4R7qWQqX6i5d1bD7o7VsCuHSxLgsu0jyIbplDoLiPi+bR9mg/g
RgaYa95fCmtH6rH5+x8pXw7+KHY+4YHZnrWoG7KGhDOP34Nnl6TAt5ruJ/jcAeiWplMjoqxvFA4v
8IFzJW7HEaSctMfoA3tKMb+MwUcKX2orAReNETUpzsO/ndbjeLkxC3SGQWel8if7fR/UGgKZEgm4
k41KBlcgXrlc7Mi0LVg5pc44sgKaet1u0uqqrptat5+rtS9fBB9jGD5/h5+2IwV2EqJqx+A55dIR
ue/uxObRv32mAO4BPt4uhXlXPSN++zQTz6T+decoUOXki0fsJBYKQdxw68antVCQ674FmExdqLvn
lO3A1pOdSVdtJj6yz/hO+HVn4/QKbucPRjjm4YQejkrx/jl1Y+7SAyPTX4WDVsNG9vFi/MhjUFF7
PFXpI8wP4Mu/vr9N8OiwdA3qNpNrXUt1LVkErNbGtu1z2c9oDoXpN8W9W4T/jRpmUZR9hwXTrJ0S
i2h7QBPyINIsklg17H1nm9uNzXtNnVGw8ay961giCiSNGRCW+oZCN3oynT9P0gzjuIvrfpUf3CQv
ioHaSzIuty9eqAX1MHxUbeQ4j9PRMcAeC4p94x3L6ojaGzclq2z9GvJvJX1ptYXI2z80wNCY755F
VAx6iD4iN6rDs2sxnbnX51kgQApocE+Q+kquzjukxUBulFdKK+fGxl1579jgQ3VjrOJ4rp2kHlf/
uDM5kgcKYBa1aZboI03TLilZXIQiWSukjy1nY+Q3JyAMHbHHIS4p+Pt9tmQZQH0gaiNi9/+Zjkf9
WS9Opgzie/iDzDQqzeij5uK7Sjl9cpr4rG4+Bm8p534St8VZ9AcaZgy9p7dEFoqBMM/nPo/SZ4iH
5U6N2b72tAauNuL4ikrGNkfoKWh5X/Jw9Iuk9/H1IYRfM2bhd0CIL3uzjFkJE/6cg8zvD+B2LsDT
BYyyBHFHfsEU6UfW0SY5a3rV47WQjrAV1PYb1lxlVaXom7fF8IHap8LYNn1qHTDBHMWZOp0/z6yA
ALt+rs1rNBVZwH60zd8rfF7OvKX/qD9kOmpcLeflfb0QSQTMZrqB6Cv7QCVe1ckOiaw3NaBtB3eK
P0NuHreEt6akJb+sgeprymhHMsQz1JqtfA/5gsXeYCzHcOL3cdGqSssZodDAjRKqRy25oLiH/SKh
J9pdYE9/S0FtThnB9E9Y+OrRGcR2McHXiw2YgDEWdQag0wPKu2GU2vLyiCM1rxMq46jIzA2rVnMs
fpTX2cttAY04Oh94Zh03memi1t4dAobvbYR1oLnscw68mHfBBelNAkOFxQB95fvhhzEJkdswa3Np
IUZfRcSuXbsRafAWjjAblQGzcVGv9Uw3m0nDCNnwzwKV3ck8hetZ1vdd5W8ei8hXvXis0Gl/lKyy
Y7cbNTeEu9HUlZtrB4nJmKyC8sM+uHmZI29pvBhByKzQZ2HmLQCQOu4F0XFvBWMCrJm+uXApFUtl
ur6KpDPVFOERh1Dxv5UT+pB6PmAgK8F4HjseKjnTPbv8mNUi7OWJaCHmpVerhS9TV7ZJ0e5GT9Pi
3o4OIWxWYBsaCCWG4XMGrffMqb2NFSTm5T3x+VivLBiKxHB6XNRDp62qbnXYd4lIh0HLr+iKycoh
D32Iw1pcxZi65rkMcVuwj9Q9NO9CJuvJhRRPDct8Yihm6wCD0B3BRdPHxndzpVgHmREG3gnnb/KZ
osBVhcl8eLM8zZFacZjGW2T0APbhpKFLHwGI3gYb2NtEqohN2qyNvzy/agjr1iqk6u5JaklYZGhl
SPOjDbguK9vhll16LM3uTkC9GiCxqzotLrXupzGGVYinLsrQr2EGGuXlUD3V0/BtOGvKVNDzjRC3
iVJDkBf8G3pLb/l9QZn3Sg/RGq/kk5iaj7YTvmWgLpfnnhFw7N2WZJ3g8VUcFqrb7c2DA6Np2fRt
1Jda4Ek0cRCKrmR0igRAFHhBG5g5FkeXdWLwOll9jrQZ7yUsQjff+QjrleZKlyjlgwhuuMiDBiLX
W69QVdcR6mMMjGbjfVTWnoYAV3HgG812VD9AST8COjqaEwifAAyweRuwTn++car24SNeco2HKzaK
aHXMQBRcXe1b3gY05lInwMpySqwHOaPf5+9ywlJE64JKE/RD9EWY7R6Dhkt1Rs1B2XTDwsX5680O
e7Oi6axhyN42nGdeev0PkO08ft/R8aBJ4ciueB/IYQ/Df4gbZZDpqpYHsggxCLKeFdl75H2eoz9q
xzEBPyb4UnyK46gynmKllYc8X9Hz4/vy/Gjh7Ei4d4piYMqUHQ/JzXjxQiqtk+tkaDandX2YrI6w
lDHDaSEAyoZkY6ffKuFgnf6oTKYN2AbZ2ZrpNOyq6mZ8b59XqPe7lcN85iN7ruMwqMawtKz0o7mF
Obwehn1mJHmz/H55o9Lb3DaLIPKpTXK+i9qGzUzgNTjKzkslVQo0rq5QMlXsVhcAGi1A/dmU2dZX
9HHMfVeZb5PyfB11izfONgxWnUmMGMlsvWcuu+tJxDiWNgxFJknxgDHDFMtEq8UyzPnZH3fshcXQ
1J1H5SjCKEjiKhvU87Rl1kLKnk+ZbO7kvo6LkXJh+lR0xcze8jO3M1wTwmI4CKPuCCNt6eOIDIlc
HBdGX6zmVEaThEgvFD0EG5b98r677FlygDLZ1fqvBklD7CppiROlSMg6MrFBdqwD/1EEpFBLu5Af
oJZUyMZi0d7SY4nw3MGgG75NUYvrkzGd6v+5FIRkQaIGQnPsFHjqBiR/otKSpd2fQ6Uv3NzKkqm+
wDytc8Q3bXhkDagzjfcy7j6jgfhe1a6I/OQZ+92RBqOiR3AcZjBaPr9jo5KVc/iql7wLHN+bTxja
Z4/ivtZ/aovihD6urkKGW5zXC/aWSO1nYQIise7qhudTVmR1itUG8y6i8v3yKZKuapSjuPcUAA0B
BKI0J7q3+1t8CBrYKDRBPGaOMD7tvLvgqvczwI7GjBritT/Vn39xxg2Ty5WM/CU4bOmbebzARn96
vDf6+QYfFILeiVcMbag+hQ2/WVQkKEu0tRKhl2NlVEBx7JCK9xG8rnTOSZ94Kltbz86tSUlmO+fX
hpPf0hjGvjNzKL13KytC7fQWvMaqz4WFPJDsBNt3zaWJd46mO7Nu1tf6WHp8QXMn9X5tDNlEkfNZ
7zFpVrwzWUpdrNQHnPAcMJKCxAs4pEzACee4o4LHIa7pcgM7cK4u8Y+75lj/6FNYDmbzm1fLCMQF
CyR2SfNOpy2qOjZfsMjRYRd38FlAOrNmkX3pmiMGmnuuFvfZ4fHqNyMrcXSv3jJX1yatUPKlo5BA
byBU9GqJqJxBF6QdcchTNRmK0n8cj3CTZYt911fjv6VatK1On+ms16AVj5kZPhSoZBmg1RQjwea/
IckC/B4PlbRjP8LO6p1lS2Om4UcKu3dgvumquyf6mfjwLAB33w9teIqliQaVjYOEJU84pvX3xZdj
E8rhM7HOZdW0uyHSg1VLNyAOtH3PjaCO1d9rooUw4QtE2zD8ybH2ggtV3lrD4jutJPYlCIcOi/5s
4eqGTxzw8iG9nSxBX+V9qmojyfOhMluXaQonsd/Gs/zBQKzloR+u3ix/dX9zzhusjo3Q+tcxlB0V
2Kr/i/CyvAsh2A2HyjTLB33tLyRYFU3tD5fw/45L0vPClG70+UY8zpScxZwGNrMw0ldP5lTuv+2M
h1Wubyla9GZxtsmGCFHq8G61oGWI03y9YbD85CsXGG7e8tFncsfH+JMOIup+Z8e1sak0Xu5tYbZv
FKaj1lFiTq2n3tBTQ5rkHgkEP3GzAI6e2xu44Dx6wjl0uH1KB6HSDea3EVPOqRfcSd+/DBlfk0qR
RGHlG8jJ35oHGK8l2vsocw8+miKY856QM11jlf0VOdic1/URb6gQaPgp0eFI/iszb5+b+hvlqtBw
Qb8RIJBZpT7/VavSydrCewVTbCBrInGMUimkDTEUciWjmpuKxjgo7WqkO3eD8fki0ZgbA1Ecorif
3pFMVquZunPw/ScZ+FIHOPmPUMb01zRn33GUeC99N9yA5MJNdlyH4w5Xf2axdiQ+Z4/Z4H1XkH1Q
XTAUbtZPzkRadZVwxziwshaTAe24XNRVR0O4PGSdQomLNLr5fIdu/vlJL6Rvv/Npeyq0BzsDuP92
kwy4pYD1JfpHnSONc6cvDS8dAhN8vCfmVR5JoOGINX05gWor9el2j9xqty0MgZvjRXzac5+lnx60
zRL/KhvIkk9F+hYuUgXEwRdZceAwrvRkl2Te0bLRNnXN9uKYBvld04y3uLpXbMfNh+fct5xyRUvB
M3yVeKUODoxVqVXDEEAt/b5ZABoGUbYHKTLwo/MEDn9B+V5Ak0pdLPseVXmsneo178DH8XTBeE3M
QwAo0iNVDJCf6rCDXwtOoL6Tr8g+fqa2T/U9gwtEzZM1UDf8uuss8m8t9cknbe9ty+lvyvRPoiR1
ybAQt9spZSd7fM3bkx5LhUf+yXRoaH5gxrGMgtZ0GNDVz3bhimK3K6WiVqYdziSOMQxBqkto115J
vu8B3Ye1p3lZdzk3usSj3PKA3JMO/d0CJlmRm1vZVp7CAblLTsT2wWPRs2f/VKNHmtjSeDwHpeX9
E8UqBY4Y06QsRzPxn4OWnBqo01z1Y5y267zlRSNpBDPAQwzT9xzYQnqH4hUC2dl90ZNT+xHDaeb0
Ir3Xt/3gFdA/YJ9H03beLjG/KXKmIb3/sd6yexw9tDZdlmFbsUh4kA18TtAXLLEkRuPmXt6B3Y82
IGuxUuul36uajMhez4mBaylOMuLtUoZqJ1Lg0ibD+IgodrlegsTraNJApnEXC5cXH9aNn5rqJ+2z
T91ta3p3HvTjSYMTjG/OPkwNxijvid3kKLq2qRPwzoFasAJjmt/qWTNBrUniHDhQyEgzfYQO4u+D
0+1XuquazHW9J6mDWW2mF+e5zBxDrqnOsOkoF3lZKJ0lyQbg6TW59lQdB/MXLZc//zi93i9n2IFk
AaJSImUH/e1RnKjaC/YpwyDDC3p7jbbNpg1yO1iN79CR5t7itv2S27DFp6+6V/IdsN5zvEDVXkrs
8YdtJG/C1SYcGVz8Hy6jRvDWnEWZq+WCoZokcp8BBEj2q60tlc+NCA97V9uB6xTp8+PvJtEHti/6
oTfWfkaq9BGimbrERHmZClSrlc+FPJ4ivsdoCkuTDuFqhjfxPVOKa5oo4AI+Wf7DKg5fN+7H+VOa
t2a7g/iaT/yzqKRxLGfU8cghSaEd7/aofRGZzXQXW+CROu2CmW0hd6rwiKkrb84xXV4NgCmFa4nk
zhuoNgF94At+esg17/zg0mtzQ+DPF88nGfHoGg4D6pmnb5XeggDQhqNZ0DKMLoDUWfneL5FJ9McM
QHSsek8XLCfJHa2MzuWYkxDmJSKp6m8Ztf0L2cM3C+EbK6mTa/zSsD38niEP2q7n3gXn/VAjHMBf
j22Ocg8KEK4E4NJ3B4ywr29CoXjFm47tws4V5ZMMzVDrCyvuwY1pw0iZT9Z00BZOQWCSavuHeLdA
f4mEj9F3ZzjvP7HXrqNH4AgG9sGEK00PxemFt6XNxidbtOi9pWIrdmSsBGql7ryR3GcUnmcSCTlv
cLJVfLiXvvj132ulr5zgnBIOHEZmTcyXCYlbTf/ukyyxMxHMyuFDrUj3O6mgme0q6ajv+HdLstrm
j0IF3A7NgSp+I02QQXGmCEbW6oZGwAdBuYcHanX1jnub2Y0xFb94dCteGmOKhkP3rp4o4cNddA5A
2VtBVrh//x9eOTq1mGSWNZg61P9I105jMpebxnEXGGUpYZ0u54ZibygglP2OkTtaRv7eZIiS2zgX
5jQptjNgq7du7CBJLz3WgLb+erdEjk/8wUnh0nAyyw4DHKCCWP2bWmCuvCXwZtREUy9Ux8kgom+/
yWeybNlXz4kXsP0TIKN4l8FOnU6ent+e+LGD96QjPIF00iU2/7eUYCzeM7fOz6Cb8QPDf/nna5aH
hOqPS4w7E8VC0tzxOnBlbowTOSe1ebP07JMsfWs9mIx9K81b++3zDG1k7lYLNMznCUh1M24XH0Hx
6ymw4Y5pNYBAHuW35TbQRH7aYeWMCJ1pGeBTztENY1AnB+4Wnwulm8S96Wwk+cKnhxx+yT8l1nWM
1PIcANYGntxkkORaPCsboAIF4XJSefFlYLy5twGAEOvkXzPQfbsaAXXIO2Csyc3N4m1H3EZAxoya
M9LKdFwht/42kWXwW9wRuq+MqiesKVS7n0OxbIK4R8Mh8mP/TzmLVs9APP0z4t1EjG+I2VdJJyW9
CvHC+uthHTuT+qRtVEi82ochRuVifDViz78x47g8lo5DbwK8So+BaoSP7f02RXj5SdfJA0JThmmM
icEz3+AIrgxCM2xWBLGIK3Nv1ScXrqYFl2z5Ph7wsj49R+9FZfxgaXedZgq8mg5ec5LgJRuFKqgb
gi6OgcuJdbDlAxEtX7/dIXT9HxGKCBawErzO4JZfTK/DEWYOvtwr+ru7CZDDX1qcZlUFgnFCUP5Y
GoQDoUuhy9un07fXlkffRPgLczFhnrZqg87PV6B5RIR4/swnvDgUDt5pFSfE/PMCmh9wCT3hZEge
P9iKD9ZNfIlV+HRMjTWCm71NpICUYAREP66Q60mQuz91oa44hIrokpl091BofJNODR+lCrJTl2Yx
747Ct20rGN7/9dTMG2Rnn+X5K4dfZkrUg4sgLSMRGOZsMYFXFI7HQqD4YE/+/xPD0mXZNN/kIf4Q
trjFTmX76Xk+WMMEbmJbGM5oXGij3D1/CzunjQiF7LkOB6FJ5n5eJmyRLYcfX3EFA5mkmsQ57Ye1
r4fIlh2uN13mgs31PHoZi9tnm7qWWMSxWE05HYQ68je/s30G4ZRoNmQ/hwsOOC4k5eVHoA6j99Q8
l9zKEauqNvI+keO8GjwuXnxFWjGbEfDKlhDviGaXV5tM6AMD2nABWQzaQe3u4Ouo0hstaQPpgJRM
Bomu8U/vMagO7gHrG5xYBqm0mcyzhy3hvImIoUBHoKAIN3mfXaOArl/cUr2jgVw07OvohAX89mAV
4Fe4Wsld/w0m/KgpaMjvPkuoOz+aN84BXMECMVSklWXfphWeZDtZZwSSLI88E2a4+J7Dm2hP6MXi
DszRFOZy/YWlENKF3or/TPYaJi+gwdJD5CojvspJb6BTlhEKYNlndlTpd9Y4y2p+ttbUTsewsgI1
zK/jL1EIJzmHigsALB7+Ik2ZzMw3IgixASPMbrOHJBJy8GFD9bswcstO++AFWctHJ5RKCI+c2aSF
SrZzKUnGKjh8LzRPQiJmT3aTqBRZvJEez+BGZsAOkf9AdcbmbY4gba5a+XULE8Q4FzXlHvXR1DGC
ymI5Sf+fiLF5/S9j4ELbba4ZyHoS5cFZDaQqkcN3fLTqanTdgYLDviIIUwOeTZZnVjGdVYwBW/NJ
wgRv3v087UkJoC+3gTRXX+qsWKxryLZp5gggtBve/WiUZieFnsmIyi5Dn2cYeBjCmJRbrs1vyHO2
HUo8eggDzF8JFHI6pn2HbpC7qjkbtQjbI5XS9e64p44JiMqagwwwhPLQ5O5+x6hcg1/UxxWLBTpV
uBONT1k46UEyDrfK+6zq4ZcR+12ZkKouIn67cRDgKaBejumDCGAlgYYBTQGWFN4jtSwdVuaP3dwr
2toyzateiai0sfnhwpg8ouUWFDe7cxSLszoxIlAgt3utCH4rcaBhkp1nodk6P1DbIRYUHfxJUZaM
jx46SOcth+13IYOochdrSW3FHwHmVZ2/Cs3tdQvGeX2kV82Z7GUw+c9azuqY51Is/Nv0Tvb2s0L2
QLtahje4EN9X0zYvQ6FLzb55apOHAQN75Kw3gSIpO8Dg5KaKpFT6iIRMRHrvQ+CA4DPGfhXGqZp+
c3mEsYUW9RUipZey/sAWVXuhZgYvYXKESQaOPdN6RI1eiMmLNsmtaXWcSg1iutcYRqno0/UsNXuf
XKqY3VNTEEac8qtHKz8yXrNvBHDT2dQribNsTvFqMZxcaouzN4FdRhueacfXeWxj50po7U9AvSZs
h3XmR+MSzuBRY4Za5aMZc5VCFHOdJkWaQy9gzqds4qGomPDUhrxbIB1WXVaVp+Eb+46zePsOUNaJ
gHY9ODGBgObh361liFVUX1Zr496bhEF40+SqxHrPhdkrAos3+L6HoxyT6nEHskYzZJXsLqaZGDBI
YFeqUymQKoZR9/2P0TVTs4hrk4SW5vHp4VXoGRbpyFmnSq+bZdHQoyj+CYCJEDGGoT3we4rL2HLU
MUYUohbybI68e8deV14UgRIYZNg4NRanGRZ5AGhEq/wrXOKb03qdSaUkSlTE/qDV2SAqP10zbM7y
WUMXgX7cdqfyzw6HvJS30nO++W/WRS7tZMicIzrc6u9Yqadgk77X69DLc5IjMW858CX3E4N48o0k
Yo+zff935urNc+2JrPj1+eajFeMnvEim7i7Ljuat8p5JHJa0zQzX6jd45DCaYTKTf5vpz8kIfH86
rfumYkpxKqQkj5GCa3QEz6G4MrOf02szCjx184OCA8xQRiHGv2hO/2tVWgR5AHRVO/2G1R5enxmc
G46kWq5KXAILEIyrrv/oMvXcavlVrWQGmG4VR5zzscA5mDlhwpjxsHm3a0FIVx3YiBRV6HK07RNn
TSIQBaylIUK3lyAHixFghdZ1+88Qwinz5qvZp3VX3RHa1eRH4nwnEfvWad5OgeNYiH6mbBf4p8Fg
DJMLXpheEdZjgS8dWbhx3klznK7gXr1C/Crt6kXqZyLYR8t+uIpAhkXvrKnPbygtxNm5RB2WxJ/e
25iyf1YmKcE9bvWR5o+Q8xpW9XJKHribdK8ywxweRd+7I9gIoyXdZeGqs2tgv3x7Cvez+pIPvLbm
C2FOBaIeX/0kFeAl6bMsvkNnljN2qvuqQs9LeL1VgR1/d9bKlXvxzA5ZhKM2h54oqfwKKE8hRz2/
4Tsah9RuXBwiP2w0mV/4J0/ElGWyhlLvWyt9+xXR4f5XRZinS7MB0nEEuWQ/bITQ+C6HcGPZyLFx
MW/Brr6oO3HWBS39Wbfn2RglDGLTAmT/glSUUG0aV3SgX5crjLJiUVLamlPzxNj5sYA1fremKwjq
i4nh99wfhGzyHQo/1tFci3VFigzv4p1NLEKAp72+QnrLNNwqq7Xmk51VBmCFtJxWDxV6ubU1lDcs
/hmqzLAV9B3C2VkPptPT6vBqZm4WYK24+fQuINCQAaz3kfSPXaohhhd/zhHIpDZWWOVHWyyBgDjY
I/0MY2PqWYzPB7l0cMNR0HKGYDAq0h+k40GdmNYyaAM9T9v7nQbnNwItozl2g9fOMJ4J7dsmUhvK
szRkbEWo0XNlZto09Jy0CQ1s61mdUTUQiEnvvx1umGJEKnSzwB+3exkxAu3VwGx3QMxYPSUq/vtp
I7r4qJHvSi5QRfcCCto9QXUCOIW132ZZJw398mtdiVajf8wH/WxqT/mvuAmlZM/4PQMfRXkhhq/F
KNGdbDiSTDMbJasPfUt6kaKtEzWqj6QPPWGGEBSSG8iCIjmkQFUzxargAX7ptfdn1OWRbX3N/jAU
F+krLd8Xa0qbcqwaL+tq84nO1gnpV/hArkfufiAdoJvkTwSd9AcTBo2V4IOQfEPdqKNYckwyTD4D
FoshOIgg4diyoio9hAB3VOVVbRRwDTbCvQTu1jMnS5FeD7v0k8zAeaTerA6jOwDNRXpRhTGByh9n
XGfVsrVBfZ3YqzgvEQkp5JEX0x8T38RwtEqlKgONHerIM+8NS1jEXZwnfOe74qKhqaTxZH2cStHl
ZYB7NVUcLAzpCXesmiV64YFmV5r6/vsCXJtc3dQMiw3Zz/7iONiJ8sI7FPYinIrufZNbajzNjCm5
iX+SdjKhBpNdDVyadCl/KmlInPgM7yFBDCUnPREC5W1ikW8VGEzvEJsexBnTg09OrmpB6hdT6g7z
uVHnDRX3x6/nTChq5KQsJxrXYjLFsQMuQXbAoytx3F3JU3r4vX1AyWAhALD4lRE3vAiLP59SQvjo
Gd+uf3AKnSpB3JWORhjxZOeI6t7smUYe0EU7RDYjIypkAlF2M5Nqpysxswrr4AcuqZQO2oqNRsmd
3oopVM4jT8GaX/VSnAm0QibNz5SlrmFXNK7KzUGYd/dlIoEGVuLCqsmQBH5ZyT8kfNEuNUgimn8V
5zfrETVGSy0rKtGXYTqCAFnQ39IU1ZJtLlQasX74bsXNIinM7D6rPXsXisdMVHw5SvsTgb37Rtmc
/bvtOlnL0JAXTlLouun2PmE/qa4VMcBCRcMe687II4pQqlpIGWdSOWNW5NPF9KzlNM0R+8weXD5F
AwJGKWPJnrSy8Ly0qDsMHaQXKlQP8xYutLwZ+CHm1wSrrj+KKnmssW9J9fo9Si+brDdbNwrfp5SO
NTeQCNwrx36SBjUgfZ82UADRczsL8+GETqA7PldYPXPnn0lq4v9PBuJGZj+jmpj894btbdJBmlnZ
2o6ZD6AmJcW4CGyVLnU279Sohzv50+MoyhjRQ1JaXbSwZbzHt06b8onPrHrHagwb/artg5lLtxbl
jt0qVbDFHmJO0pcAHXcpSmGIjv8d1g2snUMxhpgXhvEY3qIetkq0Lj8FnEj23Mh6hugm9OUd7ecQ
UJ/+WAe2FgV7nbNPiGmB8lfRsja80f5R78aVr3w9sGh2K3NxyYoeZGvI3IV0FQgDmD0EKFSTwPOo
VLlDABvClR0FAIkFrwZGPHxZkPJGsmMQhl9xtBzOgY/rJnBSPam1JmbcXPd/VreuSM73kaogXfc9
4waq7lP+j+H3NuWYyt2SVVmiO/ZFQ1z0VUWTJRoiezN5wp2QrdntYwTjy/OlPkpDaJ9zr4+14Atf
BqcYTAlcTckW0OSgNQ30ML5duimsqhoDXw5M2nRbbuvKalKXOjYOnNcL1VMlUSx+Xjcdu2m0oZeJ
bcl0GV9jjImjDnAu/IKL9uOF2ApB+7LaB5x2yVmBhVypWP1dzvey8lEXBLoNhHWqyhkoBn5zKZ9Q
lN28DXiq2KpOHg9Fcw9CkTOQklrKsIhRrNQhvKRulLQvwIe4+6MvBQCTQPwJovqOxtTnt9PAHR7w
oU5PiUq19V49C4mYdQwsY2AmGEOdBnI5E/hpJgJl0QD3q974ZSehxIcQeZOTZLB+4wpDUrA+alRs
tQRMLE7Kn7R/5H6AWtt/2fUZoWs3RJcDwUpPFYODHVrk3TTwKMAb+FVKUr7INbSXM1XE2/QGIYV0
lkup1xJfpikno0fvhZopf+APF9S9P5jCAs2ALanxn1Qmstlu8t6VjIBQjE7Bt07Mt7LjwYi7AYHN
oAZ/kcZ419SJ0/K0V43OVpxSOBI+S8evWFOKp/2E8wwY5mtXMHZRxN8k0rrYv8XApJTITJd2pwVP
ECtTNaiiQQW0LWISpgKF/qt8hI834aMT28GhL4CfV0g/2iTmaqmZHa9NeRAZJm2lOJYuwNgtoVuM
8xhbu1sGtZyJZjxH1bOZdXXBWMpRe8niyFcE0taop7SCQ+R2NUPYMIywbISrSsw2Nj0gSn7EZkJ6
p/Z+fl5tCujXgL8FnXzl9c1j15Id3hGn/9Xqsk6FSSi9y4HEZd4mEZJR4MEMDuXphHqoakuoPD02
ENyBuuIIeEdsnXADDE1fqVqfi6T5cA6JE6s/HG/eQqZAE5DDxdRuqsjfR+isDCJWqzmcEvoREpws
LqV/Oxfcf193/aJMiQ6V65FXNtUcWQ2nYkSSUZZEALSwHUpNdD4CDkCjzy3oWggWb4iUnkVQWkJL
XqhoVT/EL+YchgKutZ0RWtKcK5qh09V4Lcep0en3HndolhSrpIkkQqAL+yGjyRwCH2zX7tcx2eqL
cfA8EvXGmKv16c3/7WiwsB59EcoPusUEFl1HtgHjn7yYfGLXU5TZ3Y9vOXRIuIrqbB+vDfOVd8vx
VtxRgFq3fHw6DujTI9qByBrHWryBPYw9UHCtXsoGUMLyaCBWgz+Xw+vA2lNmDA/kGaSS2CwJtjH5
MtYpM7e5hylxFdZI/rrjjUJ0kggBYJIiigdDoMnw8L/9nX2TCHD2XsEQ+H3DBOr5D/GYOiIRfYPO
4i2M7Es+X8L/gJ0MJPzpKbbjhEWzMS2rFslCUSux5Tu9CKb5JmFx8nV4WOrDRXKVtDjbVlm5CSOr
a0vvkYXYRoWMa2dwCvzWMyQeSnXcNr3B6hawbgrDCvcf0TG+g3Ovxr4oqMxnZQzcZKonnuK+HNQp
q9wQoZCBKJ+dQd2AnhbdCly+I+27UI48tsF2UgfgMyXyAiR80ZPJYsuETQyBoKJT48jr7LyFTH32
gI88+QqQG7lbzWOFKi4pD6R7kmp6Tf7Vbc+CvE0xuY2+vmesE4Pc1NAhYsJ/pF8PG4G7ucG5XrSk
5k1iAUxa26wIXZPVS5XBVdBEIDG7B5pK+92NCwKIPLaQ6F6ocburYSJ+Zpt8su3bAfbyQslmd0hL
D67018w7olU6GnOh7qO+fQ/6IalMwOCcjfUzQ4tI9j+dDWJi9ajwgw1sDBbQDRxF1ej3RTUq+WLX
Kr1eojP+bVFofwaN7nnuqs/1PhwSl3cXd3Dcq+9ybhmX//ezftXx/2j6YpcQD/gyoCCo+Eb4yazL
jbLrV5CWPN5/NXOmGKlP0YvvQoBPUvUtyptlrnZVDh5FGzVQLwwp15I1iWjumV/RTDkL2R4Ie9oO
b7M21BBm8ynqcg5dNZwo470MNrwKdaTlX0lmR4TD6oOGIDoa0kpbrWeLIGlwtH3sc1aMFYwDBVuD
/drUeX8NOEEga3zWL6FMS+ZSE6N7N1WzF02eNGw8a8C4pXH87o0ajzsJxDQRZ1M+Ot2jg3R6iyO4
jGnZgOUha9RVWUdzeM6A+irA82TrJ3SqzH2w+5hknNmoOeNihpT7QWlW8yd1BojY8w/zPSNJ5nCO
rJozlptYtESRqbqIU2ci1uN4rfOT28fbCOwrnhMZ4d2cwoS8OUU6qxQRlNM1CqOTtVYIfM5Q/FUl
ukfegYuBjO2hI1wPwoNulqBreoFUoQOL1Mmyx9VRwY8KcONie52bSs8gojTsU8ih/Ibzo0hXPaDr
VSZZXF5Ao88j22lFcdRZn5YtnUd0ujvee7qB9OWCUhZASB11rm8Xfj9RRYeoXXS+bsSBYfmKUYgA
PlscpCcRHzJbvpVsY6/oboo/etPmi+3TVJdWhkWtkz6ZgibIlPpe3KnF5etZAT0L87ZbKg1ttzNH
thIY2BjcY4eZJiJDOSqFf5zfv1mD73KuO4foxekOGjYmh1hoL/NbV+rOZ/C6iZV5vHEoSbzD+gLz
O66Bp2NJG2OCFblip0M1g8nEh2t+d/IdfEyU1cgso+RAIYuh0YRsFgO+kUGNcfFnSMVC9xN2CwFs
AfWr89I2t9KtMP5/Ug14xWhKbTQ3OhRQawWqTxFq+m+/8w0z0t54cgXiwz2kLrsPA5udB5II7laS
j1nEVgMvRKD7is/z9jRo2rk0BaA2mkOP7gBnUmH12wc2JoY0V8XwRREAvkvOpmzouJVyWWX5QPGk
exNepQIDGkg2veOgJtGjUh+5dbHrj/Dn4K9nADfbBqJS/ia+wOQGebfyvSZcyLlxheaA520wjz91
MgkhjFV8W+aj5JwKoxO//fxfAg6dAPY4UrofPan3bel4i1G3WU7lBSNsNKFcMCOTuzxZtC5arUUG
YhfhV25f8byWjJfU9ZyEUhGcddyqpyZHT0YDzrzb3wHLQSEy6bh3qcyosjQm6byx8pNzd7OiRMJt
K6XtXpoXZFVdRD6JUlkVDRZibm4yFdKUhUDkZK8KEUFDYNCEJarU5Q+jGKetA/1oep+8N2r4fp9g
r28+C9QKq+A5doMav80Xuck+H1f9HAd2Yf7BnzWWjLcC7XS2F1lUK4wwwHh+BLJROW11+W1oFgNW
A9kpnz3sJ/1Emwa6pCEKW+lTZvreExsaYX8LqCwFmkT1AtKM9vwTFcAgjCTZKuQlxj56Gtr27M1v
X9EK6SQG8jNmjd3UbnZ9bGufuVuBiAe/iJXDyEcOxbrziCsrS8SK2YX88Amo570f0x1h640wU/+g
fb6z8zAQFsCyaXYbyPZSVUyJPWi2a5V/sVvJ6ooZnC2YixwJwDvUXOXm+4wjZoydhg1ojllIhUqc
sdwrBz+iRlCsSp0lBHFtriskowv3l7gLBJe2YuLQt8uN6a+DhAHTuo4ePgSzdxTQmx0xTqA37qvS
ft/1zfUKGV7yRP3fNvDLWJ4hydZfWdfmTyITrr5n8Bed4u5zFU78esMp27Qwp7tYK6Nk3cpXwuSP
seGDtyaE98e4pidpf5c1baJDw1UcLabQlafBDfHUfvhWcH5u7YbCLkRCeStlblRCQVIhZvZuMRn/
tgDIeWxM8RnH6sd7v2hTy8SIwmYA7lRy0fXrsIOPRUnT0jJI6zVzxgPE+W/s9sZPKgn1bvUruS+e
626O4HM/ziYUUj6/V+faTkvK9n0BFakT2CbadprYdsQhE5vZ3/OhqKo/NgYpwUIH1Z193/eIDpzk
vpI6hpqpcisH+2K6Nb5Gb4Jym7U62wfuxg/x5mBZMwTsgjsm05QUU3dgScVXP30rJwbZSLJk3sOy
yzAbB71QL3+9Luk9dnMVJMvqxln06tlxZF4zGnvvdVQ38qHi2E3fSTL51ooF1aB01rK01WHhUtuZ
qFWPh8z68MzcLtuXIxoIFg2290FWoSDelGVdW+Zi2g/7eod0MDwBpPkC/F3zpETVYHFKEQoJ6m6B
r+iaXE2bpkuX58la4DTjVgdIzXvsh1YN8O/AT7waamhyLKtKlNK7/y5x76421hxplNwrape76+ay
PjLOftZB+x4dim3EUMmDmVroixFp3b46rcxzW/Y107F9Z1PxCbbBaco+lw3zFnfBIc3prN7gA0L3
u9nNJ0/CPEQqxr2+2ga6ptlDPAX4DOn2T0uQ2Y1dkpS2f3KB8uGykgDPkVVWr1yVsscgnXZvy+v9
OCeip2DWBix2ZVuaqA7haHdsiC5Xh93hv0MJ+OzCurxyx/V1LNueTeFnvX+4Fq76+k5l6+ZST52m
Q049XWyGmD0NfQU5jUL4VqusZMGodn0rXCmSILLbXA5ZhBrYdt7ma418+FHY6ylq/joCf+rnpnTn
NxEjNLjU2PStpp7G4vG6NQREhyyGgyJFW7h7NlrlpBrBNUTQ54Q63ptfK8Ye2ECvEvdQxMiSnEgR
wiJRixnNAHnzk/gKuIcy3j/7K3VluV17GpUoojF1qWl2+6toIEwV5bKpXKvfDDkxR9YL7bZWILMi
bhzxcmPYIbO8JHg4pXlxyMxDW7MZoPziyVn8dsyVVhN4Shuaqf7nt270d4IMcQ2CH59UIAmQLvw5
dsxPbP4modP5TOgi+NnbREh+NKzgWEox7AK/eD+93clrmbMEJNdvuLu+S53vpuVblTSpQwBBfle4
gc1PpbN55TIxFcUfg8+b9jy6nQV5o1e48RNgwvDpci11YEO8NVUePZN8Xr1b97YLJUHE4y2v1HEu
JnUo+WplkhDAyC3yxqkU+lnIaxMUjYqiRi25hB8+Ou3WTo9+f/rR/h5YJRfPkxF++o1T89Bt4DKh
rY4IMJatGmTiR3C2McZQ4qME3BuIoUeKwXpCWr+7h5TRmRAInojXO1LENu/pw+rzmN9mUQ9wNxLm
CVE8Q0v7jfh2WQyaX8N9lklNgRAXa7T+HfmJakInBn0srUVlLfrUQoZOxsi4beTOL0A7d15u0fWG
ORb5R04zuOa7rAxnP40KoH98x1mjOZ1pf8C+zCBu0BAZQgBciRU5AsyBbWK6iyZnImZIAwT6m3db
9id5qhAI6SoYe08nvaYg1wwpjw7vKNeBBmky+s6wMOiy1i5HBbXt+7xc/lL2QHDSnhBdqxlrCPcM
6T0t/s/r2t2CwkkhgBymy9V4VL4Fmrrln9WgvmWEB49BPyziPeg/hh4bODCKizThOhJ0a/EYfj3K
iijQFY4FHquBv+hjXY6cxryPEhgr525A+ApKs7bo0WbpwedtHqDu9fcwL1MnLIVr0NIxXr0wjcRL
GUV/Qc2ngrpUnOoSF9k5zyumIWHhGMoUCcMDsudxiHT+iWYb2nO1lSoiO3VMN451wuHZ2HlR4RXc
hHpCbgHdXzoM+3zOpqHIB55Qwwy8CTwhIGtWYsCkLW/wm2L02CiHJ6W54LyndgN9Q6y3zB+kLEbG
Vqc22AgnncPLdlNoNhY4HK+9kPy7KUhRTsVmOZgLpfJeOs+nZhrwckS8Bj6KtKWQns7RlOefGqHu
bn9d5p0EHjRmy256LGJQ/VluEcFqkwzvrhlelLXWiajEeb8W/8m2w28r0xGIKbWi5L34uh7Yljzj
ZytNHl/QvCR+8KM1oUo8fCb7NlOzJUoNRHoqadYOZcq6/BdEYsXNyJkGXDdYlRmrQfHOYRUXdqhf
/gn93vhnAEq9m/qRiNPXP6U0azavRqLE+LlMRYrKc3gvKXxTYR+tedbIAq4X5Cjl3g9C7gC8/07e
symsf10ex2tEbZkdLp6qNU20D8/95aIV/xhWFLmyuWJhT/+Yuov1qL9xWNhamiwl9/SEHObJR4wH
SKGoTYHVxbV4afH5CDz4oPHjCXDFGhmkj70iIsAec1a4kXBhyhlgb9hKm+RvHdzeve/gKX88LgCH
DXLJNFP//ESLdzESnS0AbuM0XEfzQJ7Pc0H3gN4njpsjuBHDgnarmQ3nDJJNlY4pTgetzIo2uJpM
wztgXruknuOc7Pkv6mr1V5++eH1vnTJv0jun4xppLi/QES9I9KXLg0HNa9jLAhre7TwVTP4knzfy
PgDZUfjWg4FDonfrutD1rUl63tL65dxNFyJ/jnip6ZXqook5Yu2DS+wFbkqQVZ18xzMIUsSjd38L
esBR8j1rVi0q5YdQ2FFbORqb9JrghQMGLZPDDQs1CLxhVc2gP0Gqc/4UlW7sIf4aHNkWLJ201CJe
fmlWybXatiV/hIjydmFFCda0nNvmjBm0R0tpnZerxMK/cLxZAxd9cml63wBPRlV2uA50ATmUeV4X
g1C9ILm1zZ5l+uGUAwe3l33BM6Cmph+Mx811Rrg36+dEwGTS4OBkhxHsaWe1LE4YL30dLSOPA/dO
9EtpEyqYN/fSKN7UlwByiUERjIfQDoWBp6Z+KScArevQNLeBnNs4fXB9U1Iz7yo9H74oo3uyL6GJ
RYe4Ete1nKve6CjFVmMlBywnEaEfU74+LfGWpMs/xqqCVCk+kvm5RfwRM4vLIjHSE4T2oB9q/sGy
v32Is/jVak1sRpMJwSCpkYSWDvZng3S3v2UR4gTkhwt+WeWtlws8NJzK8z+TmR1GTveQuF56NjSA
djdddBoo8AI00iCoop561GKcCGkK20W8OlQKGHh8FQnlXRoNEYRYTKja3gEyRwhkmkV5rKIPkaNn
FhC3jXfmRG16qsPLitsQOb4SAZIvlb8xBlKnWurczziIZDlkckX0tp8srnhugQofSop5QME8RdMf
VJjU4QvwguiIUgZbpHcnS4pDjeAZgFuTvXPlXASNnRtOI0VOVjRe4NyCjKXOd/XEseQCLPWWSsjq
JE7u0gZJsz5UHfmO3IaADiDS+KE/gA9Xl/GLomHfcLdF8k4+yhYbMpIuSgp455kC8lQK/InH4BGn
DbObN2nEOTocVHyp1M7DskM9YC3PkXkPqIM3pLLpm2762WW72r6UOvqXuRRgPYq/RCAxk1b1yrU9
wDoGESu6krX8/msugcO0SgjmBY7N+iQKje7rZi8Vku/CDU5TRUuWTQzz4CHLPW6ukwwJFPi9dwbQ
VSZ8iLz8NsakexbhWmAWQgFHRrfTg3n3sSTNJCvoNHV900MvYdbhJ+XWdecCIu8LMdZ1N91s2imO
m6yR0g+X0tgbkMvJ/0ZSeCJHM7UFph/ts9Q1mpHM3k4atK82vKDW6ltsnjLFzy58lzCgqlWKbj6J
1mtTOWFLaCrrbbZ5RL9cW7OBN2YpfhKDzZIO+O1rfecQj4hQaFOnzoShE5FQ861waVjTK5fbuZJQ
0YOau6coPN/e8nhymY1taHFh0kUFe6n9aESy+/rxQpkSFfs98PzB3px9lTJlAOR/C2XMCE3Yf4c6
gUttR/X06kx1tDSZCyQ5yFpG2kk9qIzqQp2syw1vDJg6L1CzKRxLi36FQAPldzb66fbAn3ycYiD0
UZqnrl5P0m2uPaJxwJ2FZVQ7O8VcHmgTWCl2XgomNW17IXMfhXjEMurs5CRmQIon/ogLHlRX/sT1
T4Mo5JKGDATqocCdjyHW6Za6PZHw9nf9/qNMU3WVUSQNdf2IfYd0+dqwVZ3HCnL0TcwuLqqKsxwQ
PjDImeWKHekBLxr0YjY40+wuQrzAYinKVgdzjPOy4HreqX/r2ck3mECKeGjpdF9fkx+XDDP1Ltz4
NvHHtjbE66BRlYMHR9OdkWjLaK15EXcL048KfwDLzBzY8CRkR2bexWXFCV+66s7faFRcq6XPF+Sr
LLwfDZrNqVPjY92K7EkkY1VlmaAIq/JitQUXOJ6fRallg3N9vFkuGUzVSmzTx1ODbrkZng1dPCl6
la4l4/507VieGGpZpqbh7IHHQhcpEHaKWOGWVcsYa1DWJTMp6RHrX8n5wxD4HZ3+zi1wTA7bG6kW
6KsnRgMErxq2cLKXobu7ffGVTbuGlB0mmnAF0+tg3CjJ1RsHFfdOFEMgkyPcBWx0FbE3rK4VlfAC
TwiBG4X9nKfaxiX2RZTmYIu/QPWFOVE/zxe9EPzA3oLpBzlwpHpOjxHE50KDqOs4YVbGoISfB9sd
i8aqe0bPw0p2iLzdhLNqXxFtx1FF48lCsJ3dy1YPeEHIoDimECYDbWX7+yWPZdO8Jfe6EsbGgZOv
nFXa2rFmcH2uWygVWw==
`protect end_protected

