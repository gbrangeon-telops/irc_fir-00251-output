

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IVTcVKz+qqR6KelbIxn6hKss0fyLwIejVgwej+TN1ST/vU6syUW6hxZyGugx/VRu65UT+0QU+88C
5SDN434/fA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W0uuDuJZlgdtFvYMz+doOP0vwnGc2SXfLiGH2a5FulZQF1GjNx3fjKnarWbbCm92Rksm2FFSGof4
SgtGKAeCq4Yz/Vqm5xuP6QHmdBwou49vkKDs52HUud9c3EaEYtdNlkb4+DCcueqZu76yWN8rf2DJ
ekmu+LGiL1dmyzv30tE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Da9hmR0COgf/nsNRjZU5mrjIzRjN0/ufJQ7crbPh82WrNgInUm192216ks1D/Quh1gQ5TieAOChY
26CHNdLfPPmjLAo5/cOIRsIuy2JD7JAEIDFhFO2BcC4GrUAhSArSC4/9FyqXrVJUKuDybwv0tWSf
qpHjmJw18CiVw84ne90mESBOJ0fW1ujayfbI70yaGaFjJM/DPm4Lq+TC+TFlaimxpTFNrAUzQNVF
VSkf44Zb11D7if2jaL6ua4hPGgYpPcisaJtcEYpURXS8Lw+NjmMExnMpUW39NqnMiTEPom3YBwag
JMKm6/EZOnBvVc8SljH7y69fXiGUXgw6Z6POkg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1/llP5a+sEX6Ky1I5ak8Fr3e35uMro1bXNqkrntPBRVTqUhQPFl7wfr/6Abnu74l73YggylsZJi1
1Erm6sC9oDhL9IE4pENErrDQRZHuFnl4+DlguLd11swTlNfBwauGoCBXbTtZ8+O70UI/sRzXqbZc
NDH1RywyQLhMRmSOjCU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OI4vyCtRzSCtjYNsCqL7rYkcvPw30aumOHoxNPQx0NU0Kc5/zvGo5pjE7sDqPsv0b00mAjKXUE8e
pVllo+uquegdt9Smrq3DaiQC/9hKGiZzOG1rJH9JbLcfPMXDGpwm1inP51BNgkQwocfUEAVndeWo
GE1Y28I9gt/5q5Fs/OUAX9cAh1VoS1OcnYX2wbgJSlzuLqnGWRIxOHl4+NkNkBq5Q3Xm589bPnnz
m+d2tBEPyqaCTvb13xXW7hqIf0ahuv0AQTuiClY+KmF0GjLdJTWJjDWPuRd9WYhybCp/lrgDnhAK
cnRXJnAOwP1Vgr7EPuoyVc3UkNsZTxEr3wrouw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11680)
`protect data_block
8m0k+kC6MWaZDIKrH0eHKwtrubY5A+rxzKXlC847EUl2mAw+r0BncJIfBna0wPBthV5lrS5bU8f2
2K/83+iZhO2cJEW77c0mYPRkXMZTCNZ8eBkJgWhxZamhMoE/h3af/N+XqvcvpHSnSfm5ULrZoBJX
YRrVpo0XCFuLN3IJvC+Z9XW2VVElr2pT7mKU6UyqX8keLEMXEKwinEsWIRyalK1g6p2EJeTqdoa4
G+sixQa1xx19aKDMNZ3Ir+PDw9RnU75T0zsY32uLVjcaGi4R/d6GFK4o+5RR8DDY74xR9OwLhnzS
LiPfVytKVOmRkUjvYC2wqL1NEqTuWs2YPm93pSag+Oz+mMDnSVhH3G70GGBqFBRPepTxoLPSlvcV
710hzgwGw2tT9/HuCGX2eBs2aNtG0oatNV3vOhH7DgLsPQkaPCyIox+KnO3TYpAslhXuGj7SVY2N
H5mQo1sVfFI1u0pPtlOV5DXXdZbIpRVwL15ozWxLQPMi1lE4QYqVJ3TOZyKmegVGD1AK1ldhMZqm
trr7+EgtmkDtVBKZmsj6h3svuOu3zS9ngI1jce/CCgRzbckYBoHgNJKqGSgZmxwEm8LRPcJeT/51
yWhx2KomNwu+iGjWCgxgAqcNI++cDmCbI2vKPOb84HEgL8nHAxfRX+vvqeHQg/0YVT+5THPwjC+T
Ma7YrqdtTQDb4n4nSdJSEmDCLGqhpLCTK1WGU5I4hVW+JCZMqT2mamxMPUaY/TuE2pqk2zYDSMG0
31ga2+UE094Z+Sx44n/vC00DlE9kjWDHtmZoCF2L9aG/k7572U4bl2uYzw8lrGLIO/gjyuWPloCM
xma1b3qggoHH93kINg5S566R4sPMd154+eQwv3PiIvhxp5Cuq/A8xjAhNpITUXJQ/PvbNjXzXGdc
lERidwGIl4Nv8lfonjp4szfD15tpS7ZkmuJW7gZZch5Je32jMIYD5mlnV9vuPIHhw9qTEArpzwPj
TSrjRpg/e1dFnIlKiifPwto4NC9VWQ/wz2PZl6fdM+StUWtz2PnPN2WocwNqAJimuzQAXvovMxYv
Qum/W6zHWWngDg3tIN1aFV0323SuV0E3EhWiLFsa0iNjmGhFO0C4rZr0MMTFKooOoeQnp5AzrpV2
J4d1DZf3lKHZlr1qxn2UMOlL9wvrqfSQmCo5HqTM7aOK4PdScve+u0M+ZcKZFGSI0SfG/XQNtX/+
J6ouBjQPcfDfD/IU04tNNiCeEBCOCXJbZPRmQ026KT1QrCoHz9nGeSeIkcLmJWse64n2QxPBEdIR
bM95DG1rFy2lYoFuw6uCS7XFSoPSzyoyhzxjHrhWwEC+S/F/PzYgBLO1YvVgJ9DHARuSOjxMEbdq
h9qIOiTyC2x06qNgfSn559BcylY1b6JJBemoODiTojavoWyQxTkfG61P59AF5jmGTf+zctiy+Lc+
j73cZmW+f2cMC1X3lQjMDr2j9OVWQlSPpEkmVjSQq0knOKv63FUBxIsZ33UpXLbadzwDM9Zn0b6w
tr7+efeUNn/SE4gAs5tR8lOZAjS5slkKp8kri0ufDTidLifsjXm3wI1Xr4iifbz9qR0NfVThHSEi
6iyvIBV7gQZHFrr4wCkKd8EjXNXoNFOgMrss2GBcoaFZDMQNVN3Ie45/OFFdCBjbCmoeqav456G9
8pIULF5alQAiNGP0ZIpW51CXNOgIH/Hg31JRHHnZ+3Ro1A8FPP3xX5xl8NSvlKHdRYYriWUc2jqU
kkje4kswpXAOBEbmHkb8gsTVD4GLwYN+SWdlio2CyeGPjzMPkS6PYB1eshQeBgK7guZUi8rDYyqV
HvZfPw0wCMf3KlP7KyNd+eRzwgmBI54OrJgsRqyBYHBVc+qq0MxM9mm/L1+77h3dNubJp3m99Wrp
E8YHewaRGzrlM9uPZ9cFtodb5eJKzHU3UwJrTPqGQo9lie12y1VO7LXGsYfYUIcL5RmLcFE33CsR
kx4bmgRJMjCWSeKPbW0KZUm2mgh/q5xLtBZ40P2R5D3DnEOVzEtrnHp3M6Bn9PbYpkCnR8xGbCYk
EISxMwUY4LKiAGpeI6qhtg333kDG7Q/M3iqgsZM2o+jX1sfi3LocVnb/wFtiT/mRCW59HP6oXUva
XOf6l3TsWgFdEj38x8FpHg1i/MWyJmZe+8LW3shM8Tk1yvSen35Sath3h5HJtFF5J6dJoGboyont
rKfu5a4afuIPT67XvP/XOK4OlLV0CzJENazK9NjSNER0Uk4fe3AJiUPG7jacEtxInVEHKYKG4vjA
QppMR0oSgSCvrO8+VBc8fN4RgoL52ZMcil9dZsOvLux0o3XjCpuEj2VyNY1WqeqZ1i69ojP7uaDC
w1cLJFJ93dplQicvMT8PPn/Nh4oG2sCNRkNpDQC3UrA1SOnAOnjNflcLZkK8nmgtkpo/vXWg+uR2
TkVSVUMqtruLIaCGweUkdTAc24xKhJrouN3GPhnnC6fafpqWER2hyOgk+zO9nFzXWJ65OUxJTg5n
BijHg81j8Jc8fOdCeMJqzCRYdzGdjjzIF0W5XrSM2Kl5DhJN7OXQwlsOlu4QqL36a4jWzwnua8Of
1TAlwKBaMatRLRSL3UbSg1CDokuv+fHM5mZ+l0fQ/D8h2PQed4ekzmAUBRxQXL0AVH/LkBYBaxhZ
8qe8qqH4Cvt0jyIQDxmHCnPBEOWitYfXE/0v41t/k6oM1Y3HysFyTbekTfZxkBUQQbfVqi/Y2qGb
2RbusttkXIUdPhPide1oOTWzKoXFzEbr+5DXZ4cdagEK/JyaM5rMrbHtY5gMCj65hnMAJ06baOfE
dL4mQvhUaGWBMm2zu8k1t+pi22NxIvNIgX9ryuXKDfZNhzM2NNSnJYC3Di/l3VvI2gkIcFOrK69R
hkpB/350YOoc4L9/sb32N1mTyv0rBD3ivUQ7Oh9eZqAuKNyJoLpJDPRmAaOsBtFThUyzjqU5sFny
2G26Z1e9861ILQitpqUkqkFadyGmf9TDDuApEwShTPdR7tHRCCUZQAkv56TBzS03yxLUB3Qdlxhy
nm0B7nPY8W50FfubAAXo1Aj83MrqSFLcT8azPpU6iXiRys6hmN+7vszpE/350vJAw5MhATBWykoD
hvdJFO7GqvbKmpO87tMcQwBy34l2umNA/nb5To/B78EcLQFetYY9swvqOjapM1/C82g5ZGCVc16o
/ssz2qtV7wmN61NJx842gDhF8QO8dbl9x8kOR73lYy4v5B+Yjo7VaE7kXAu+//wftKiuT4/tcztL
CpGIviDhxrGKXPMv88GuY+LkannyU8XsVRClILb4VMVk2xEHnDl7qiBy5mdk4PcHnQPFUtelV5C9
nkDiVWKK1wkIOmjw0Oy6nm5wuB6Yb4g7ozGQa5DQN/lDmZqjYrj0s8q5MlEfAjR7UusyOcHIBlJ+
jAzBUeaUN55x0rZWNW1OzgmDbML0WAtgWZjnCZYqShVMfqqXcha+tZrlPfh5Zg0/2QaOXSQV0Sop
K+Tx2OezMopn02ed3jL4TemRLHvTRjhG2++wO5PowvCPp1E1C6LWgr3/NiXNMH924NKnJ1ElTYCO
UOgdeQia5aYEH+S/aZ2A1VLGtucBsoMpCSAh90KbUdtjObFv36rgT++OA6SpBxaDnj+UOOeATk0j
70xVUZlVw3RW/5OC+MRDX0F3r8cBRGYe9IORLm86xCgmDRSihsF+I3TEmzN/2WrR8LLs2evKIxZQ
PIqKxuLhRAtkuCLu4JAqdjSXFATZXBbybGVl5Xp6jMzx5nJasCIiq9nvacXB5Zs0CD1VNbSV/A9J
fdkTdBqp6rHKfc5iampsqvf2UvyNf3XYvLDSjiEaXU+jyg9TaucJKzCKi6nf0sVK83kHJ77TQiiL
cvTQh20y4Pd50uDyvnfyGMN/14j/bePhkknUgRmN98Z65txx/JDrK81MOt4+RKI/HoOk0lSuEKn6
GC32Fri3KjKFsE0/aZssk1TkLVY0R5i5Rh3caua4Zn+E8S+0MZfMVlS9sVz2UGGjiY8qoYXDfGpZ
c9PWvzJNq40/y6VbgM0gial6OwpRfq961aaQVyBckJbniuavSFULGc4oj4K0AlStRMHt0mHoItye
0rv1qNfFa8KDhmsqcCShhoOhUMDRjL+bC29vih4AKzGJYQh2z9FvtfygvA/6zAkULSRaLX3bVdzZ
5dAmeuxbkwwta1+Nxu9QBrK6NO1UTNmJKujKoSkzkzkySn4iav9xGLwdl/CkazX17guWDqyZKKiS
8lkNa5A9oedzm+6uuIWGZNmYr09S0Cm/MjO18VQdaReoF8oZgOyyaOjwSX1+LI9dUq5vb/5mujhz
09onUP2sgLLAhOupriHl8NoZ7EekDY5NRUCKPJk6CyVCSMPqUh0Ss2MrX/IfKwbQgiyk/72YgKRr
ewoX31x3BBhdFpqZOhcYW5BHRiYBWazfAbuvMu4QuB5nk4C6kdMytt8dBo7Q6WpPeGT/gvjUsfd7
tzcSXSMlNhIq44HGPiaTloQCBCIcwdYBdSLHKpQiVG9c1TS/euvq1WsOFhw1s7/HlSY7M//jSrSq
vpShR2+cZb21HLOSPB2aFKq3aCGLpbwhZ6Bq6qhndZ2d25YhDezM02E4NwtTz8SNJdDTQpRz1Khb
3vreFy9DPW67J7AbMTUml6Oa+Eu9ZAh1V0DEFBLR5Ij03RYCi+/NaIvFPNABNKJK9DTLVNdi0a86
MKWmeGVAllAZQlRcrMJnw6cy7q1EVbEyNWzOaDCYm+sN3jtGcLap2UFrUHRV3vUbwA75h4QIbZsK
NC7V5Ktb9dExcHVTAlxMIJ5uNQ739oK+eQ6pXehpBrCQ6Iop+z+KUwGelRptu3LUyodFqtQNlg/J
aoD0QoahISMOrVSvIgPQ/Gf+dgSMNQ6A46fMje2tvVgN49NG7qhdopAaoTnVhSxa/brrYzxPPjbw
4rTzHTzdxdUvftkiYSGE6B5PM+lIajpi3dxVLFbFVYbh94Nzhu0F2WtxF8aFI5MC5vv2odpjUoY7
So/Whd5cFdpb/TzcvKA0d0YMEza4qRivOTuE21KhRN7UHGEhKvpeapQ4TFeadXGu9z87aej39+eV
mQEHC3K3iTgL/cqbdYA9G78koJqa0rI8uUn9wAOuQrbmSzVU0ARssDMFf9D4Q/STqiiP/ow/qAhv
QBQm5VuHX57VOtl6RxUtIpE/GUuZuqDHHSzC8BMgTMZzIp9d4dfXXrNZVuL6eQFLzgFH5gEbaRlP
ZOljq01N5HY5NnOR8N3YlcsMhVwgmVxjc++Zh0GlmRHXZEwVscQfT2RMfAzjAA/8xBTVWUKYy3E8
hpa81IiVhhizTzDNjziy2K+supPUbamVPMMIeAqTZkviqYnqmYqiRcWZpVzjfovdkry+Ug10m3Zt
4QTWTa6pyWp8IGupAY6k7FdS67qgYgCI8LDzxjVcbYJUkPQNYlZWbQyvv1hpfvCeaDJNom5pRXQS
47CfEHzvjd4C5VLaHwINzreTMg38w6cQb0gBd2Lu+nlh/mbebFi70SMTWyJ8fGl2De9FTx0CJic8
FqiR6uDF0jBeWrh7jD4xgBubkG20+D43IBn/AfkopfLGm9LmJepaekT2jQw1IUnn3JKtOnXzjnVX
mxv2xbzW/0A9BppHyXBS73mQcmE1nJX5TAhkCtn4y/cMcq6Lm9gZNF0ns5jlYAyNBB1ghZ3sw/ZW
73jkywJtBCZ99856BhqsKZ/JkfyE9541sZsEEiuumMHZfNhonMpYJyerpxO2ul2gCR3al1FRd+or
M8ukJ4SoUhiFaFEmKfCh15IQsgYHSRsKsKC7rRazDvIVh+IujVoKk65ZJSsswO4fXLNnij79NbyZ
2qJexY7ZH9xDtFSU6vFTi6BVYGT38LVq7Pj3k+a40H1g6LZFoNAJxXVgbrdUx8gEZzf/hJEZh72N
tt+P+s5gxMNq5IsGmchVuCR/JYfK3UuvNq/hsD2V5I8TEU7glb9h8vyx8Fl5bCwFQPe/SGYt1ZgN
0rpxeNRB5CUL1Womo8XI6B5M0MbM+aLFZZ9emE53YOyA9BX35S9NDw6xdkhgRtl0Jgfbtr+1ishu
0Dgl+9TSahvw3Ay+YDF/ZEHAhpL0ZrnicNyUoyvVoVjuVulpv6bVcIA9PuUraGz8MdkWSmH0BJa4
b8bEJxzv4tpHUiiQWuCVsnd5EteZ9GPjwjBfiixRCp468R/BvwtEuKNbnlg0uEz/isOXqajQ+ri3
Lt6GuBa3i0zG0r4C8x0V8BnNG0ru2LkML/yS5BmzMpAkk//RhqypMfW9y0OoEUF8VZzg84fEQ1a3
fhQH7JiA2vXKntJ7SWvJPI255XBqwLGwAOSDh4E04cJQd9jH9WGrSF29gG9nVL52HKk00BwmT5Rd
LTLss1ZB8qYEjWKjybc11zpz8waCON6kirx8SsPY01B5QrEqEfa+luv2zU33SJKts3xdkoETlkTP
C7o8m3RuOfk2gxS5CzHV0VCbMLzbf7tTxGy7gZu0NHgN8AzfAfPgNbIrR7di86xVO/LXBfnHqduw
WsadITDDc4CE3PhdBLod5u4iLxUS9pltiWhP+X1/oTjgGS5GONpQ3xZtTl9l5jC8oseSEhOvC7mK
HfsBzcOiQ7ZM003qBCzHMi7ui5pS72hZiGsq6/RK/3AwdaFqipIPLCC0W2j92Llw7vhF9tFU1b5U
oaEK4BxfjBNJZtyXsAK+skFq6rDm3NY9OqX4iA5rZeaFKbeK559AimOWR3+IBAB3NMiA92ZwGHYr
iaI0mw0nuKp8Kl4h8FCL6NgkVDcWh7DCPFZ9bBS0cQ0p+z27iJQWQMKsuqM9QD2kzckGDaLlVZA6
DseDRFcGHjofnVXTGmZjD+eCGXXXA7JJorELgxJ3JUuVtb+zir9r1WQdFquodG8MywPCR6Qg9Jjb
LaMv1GYPyDBbRRXb3s3qo6YrZYk1Y7emjBq1xTY+ql0wZEM2UoZN9J05yVSQ4AoNKXME4OGZ7DJa
OkjKC4UQah6L1qYbkLKbUKrEXGArwfGGcz6ZRMaiPX0+RmvSZdINsU9u71M2mBsmKeokJZfANiSC
UzOMkXSapVsC7x0kDI7V0HUW28JrQgn0UcukDOxhmR/3c7o9PkDwaohTfEbADg8tisOTwTjYvC6J
Ob6k8+loOB8UxFLVJxUkYYr+18BX0jD4TjWe8k7By4XrAX9euC1k0JwDmdZi9aYgwd2F/B4Ty6gl
iWZUwfi7K69O2KYMvU2aJOJqVJUmPKwlZp0IZNVjlfpm8r2ekBcIT2aO/fDdULlwamT33AU0fCBL
/hQ0lE7Iw4vqIpt8xiu0PO/2VCXZrW/TQfRWqfnhoVVtGkilwrJLEyVABmTsOofoylxQK1FSqIXM
zg2JzMFIfwSHUCpaGa9bsAQNAqo4YojRj1z9SBqbEcELdJ7CCm1smk/4NBQoIvUTd/fYL1pI2n02
k1dPKxWAELXk9Ryxkn/UqdO152pT3VJNirPC8rxa2ZsE8jo1bmQ60/Ua+BW+sQjHGOCV0NBlbyvP
wN3htsMaECcIGeZCmI9FFzrlnjLHVYOfbr4I/YNV6VQGRiwY+qtFpPBw5pmRO9RYa+Pjz4PwCcHG
t/PI/qAfXyQXttWAK0gBqNUxz8KR7EDYTw58igC8U0JLUSsRwQAEePbjC68B9IuLuFGtEvv/3h78
eVA6RdvNrUp/rkP3ut0l9pov9N2Vy0i1g+KHwSjokiKB5Q6wdALhTLntkxW53UfLfFQPzESJtyRO
jr/AtwVE9e3x0PG6jPU8xzI9hmw0jy8oHj+s3ZiMJjwuPNewtAgdSTntcADbOdPmEATHy6mofwI0
6qnNKu0vez8ni5wY5j935UC+mHfIs9gAtZU2MgtAxe+pzo5Zma7WHj3vMlUp3wGl9aGoeZYwOBrW
sb9E+mZT6UfuBKoTrZqAwfHsVGY7X6JLl+kWxP00YCcBOjTXRECg3Vri2RjtCi7mhamfCWyeB71Z
x21+WNTrBtQB6CjUXOueg0i9u7EfQbOr0v/yc/KQRct8BFXkDLoXFcoB3TxeHuiXdJoIM6Z566Zl
2rQ5gkI48OEyLYX4Hlpn5lAx15iw8rOWPWF/ld1WtSHqsYHxoAKMkA8PnqrIEgqGZtZeuqOcJx9+
HHBLYhLXpFZVHw0vsnLvpCNDHBNsKzv3QQCr5l8RlAGtfpqoOQtRBdBT7DxC5GTCewmU6SR/b90W
QYUE5IkoB/ZdMMRGlAU7PUeI+aZHQwkbmEVl0H3K64xfugr+JogCQTZvrvZ/sLSXuPfOiA81HQi4
HalzdfqCYIQsP5ds9pf0PF1rOZjmgRB/yg0luZzOGxCOawePxuRBAK++WjvqeJ/maT26cTc4XldZ
bU7SAHykNlipkZzLQqjqJFtdosKp2awycTkzl7cPKrJWIQzA/MJDTiTHUVNroYQx86Ng1K9RyxJV
lZ7UUloSt/HdzjhJXgBt9Pbf5cxM8nk37It2Xo+9qr0coCb+VmVbfzf4X8TsC8vjZvfrwBctBCl1
7p7Bxlm6DMAby/CBnh0ANwv/pAJzQV0+p2lmaehGeC2ZIqKR8NIqY4Ngpm3quGkojVFTL51ah5ak
C4FjRy9bLThP3QAxkSK3eRR1zP8zmMUAJe+5qnRZOb5c3nhScK+HUaXt2AqpuNXDLYG3EpSU+Aol
6dP88w/87uTkxWFhDxET62bLaKkgR3Hb9kcefVcHlOpdZH27nG64HSx90rgkLIq114Pr5HQPEd2z
L0wODxAnXGApGn2SEY+clSJ/s5S3g9fufRrWyizTHLdNMRYldM/zh4vYmoDQ8p+HU+AzCTV4HsYR
/xD2hV4hc/9wPWYmF9HfzLjhGm8RVYetIQAfZ9irft0tdMbZcjcv8Ay+Cr5Knf2sybPpmSRusMov
r/DewKe5/SRtVEJwyO+IXCvJOKL3yzrhp1WK9/2+BKErJnR/ATwfgBJHb+iYSUF8jt9fc6ghZXQn
WEnkthgucAAbUVA78nB8DyKvgfpCHNhCAyQu/mp/9iD0AOk/HLwaROQC6ZNUqJYPUgtbXCTVqNd/
fSepFNycRzyivjcLYbPW1uoRTRwSCkZkcKpWuMm/p0mv0lzJIE/RVxoRhMl/BjLXUjMWOHtEh6DF
ocatltzGaQ3rLqULb79zHTKnDYZpuJipKSEdcgy5cyZx3v8WWPIFUJIdg3420+VPEwBsQkwBC8eJ
3D3GSE3y/rydpdaUtYHlUxCid9GzJCuRcs7meNymTIjQ2kkYJPAkJjZsQMiKsNQ1u0xC7uq60zaB
f+wosOVLDWBqaIIrCh+N1zluQXJDxmC/RlUk/XKAH1aFPdGb2p/DGYzHTxi2zHcT8wmV/AlPGjzc
IeaD4iPDNeITAJeUJSbZoNLXrjE/ntr6idAX2KD50W7ABLNHlNjKMHVmw+yxOXx+4jdUes3Mvx1Z
YVTQVyNZbCKT7u9h3V8itSfKU9RrkD1wAyp3uUtYeBIDcZYrL5P61/FGEFVJeMvYX2bIIJOXIg/j
ZT4CzGb7/4rjFmkBNV+zUBlaWhBAPyn0fUe0UzKMO1L68E4eApC7IFrFo2f0matC8CtuPGMwf7Ah
TAlkY0g/HW77pKfvs6KRTz48/9dfm1rHT7j43VNc4ekdGM1DbaPcfy0KeJIZC/9g3VARp+xZiSUp
IAaV8Ai49m9MyDvKHWu63uPt6hdLaSvt89qcYJhxqNliyaL8QnllVG9OU6jbmV4OkwwBsHJlI+3M
W98CDBhNrp2iMp4jNqLiAonHosjmBGHuoVBS9eNWNpqcglot5k3kKxk/Xw9GPl6ievRBl+dYhc/5
Sqz6xY/N9rp3I8ZiyWobVxu7/Gx1tV49mDKRwUWPlzEEGtd0unP/y21zTpKuuMLWPjSNfP7VdTp3
GZVQvgnIaR0fllm3Na4bK5EsDnVTUIKOp4tNRxojPLaAv5wvqJ882p+8zOy9p0k44YjtuvPrv5VE
FMrA0pl5oS67E12qYnE6ik9aDJ3SXn+HiNmPGhSF7s9GJrloa5spCL55kDfViWwtnyWtnrXKzJMl
BlwpWbvhCyIsbP+93frn2LthcVH1iOy5QfSLo9kwGD0Ag0tfVA1rhHOAMkA5NBoNEj7BG567qJgE
1s8jzdjOnh1kdSd9+GeY3ZyCDkT/WkW7zr7/rlM0muzC0Mk8QXLLPgKLJkQ1jYTW99QGoVEttwLY
vmEVk4R2zzRgJQylZszgsQ+mZ5LyMF1TlZWgnx8N7+G87XZ9h15173eYV7HGvUaYz3VSrNPEdhB5
wFDNObJMrsg9MP14VTsyWJFY1KFnlc/o3jfPGMfPftWBDQswkruCHuqFH44fDd8ouSSs0OICunmX
6XXemAucqDaOVqgwrNGNwxzQCejKJjaZFo9xcpRIGAhaPuEZbqPQbVbOVgt8JWmAS5iyMT322VPi
iObgTUDNTqa/K6hyB7KvY1KjKkj5tvokeZpHDmWbjyP/s/db/pFz5UaHQ8/K+BKaU8htGsJdszL/
v71iGRGYZB4ZDmoqEqepA+yVQ4eVjeUn0x+4hPzOAp8KAbucNBADSlY1gEUZkVHRruPg1fyYsiP8
Cp4tK0Vo6ryOEqWPDh2UAWkM9SM10sgYrgIctyG+DZq5BzpQQ99KSGGFkN7QMxtwtXyovtQPVQ5m
tkANK1QWLUsjsTOqVvDLY5IJMnEnbblcDAgOfrljDXfyFnRrQF4+83om3et5vvchqGVHU1yku3uE
E5GbpkDKLPv/rmsH6/ZiFWHzHoeLPyENM+Gww79a4HmvlI/bH4tZcWReJQJAZQBOeSYUxCwvH9RM
xdMZmRufUKSB/B/my7PGRhQIpSrY1fiT1UsiZ4tJ7gD8i8wEKxtmrrVqTnvbIm5q3tzmMFnHsVb7
6LYNLq+Qh0dTXgSiFl26HyAJ7N6KVHbLLWeOqCTTso8pfolGSYn3MsFrMylhZEl0/fBNai9sqZrt
mwb/OYkOmAOFF1JCTN2HuYeBWHfG5YgtwaVAlGf+jFSVlpRBp2gFf3LMllcKyVUpTviZt/QF7Y5i
uuJw1T3kVPMapnnzT0p/2dL60KcKMwifN5tQoFNaK6GjnUWgpFlm/0aFMPQfS+5+mdCn/95Izhmx
5Kl7rOhXry0DpvpA0VnwDTj5zO8YOcQ9c6ENPq+Wa9ylW04YolEDMXMYP4u+OGKVZGQUCTwxTDmF
ssJFAnmEtATEE8kxPrpDMBm9ZySENInEkOMo6eFWqlgGb8R+qZz10PJ708ZTq2QczwKX5yfD33/d
iCjZRyIVv9kW99taN3W3lCHYeVcMG9AANBqmy7+qMEgahSd2RVNYE4qxiJALrA+8voQveC0zKewt
favs1V5rtqdIw3P5UL0ITgH2T6DmPm6x5nJYs0rcaAXcwAe+fLn2CqaiW4kZPISFeksKJK2Suu/T
ttRg+xPB/aOJeCgUqhlgIVaHhuNMw4x4Mo/nfqv8J7WvW0vORAdromfx9enOCqwVD1hbEJqaysK9
+WP6IKmRu8siC2K+u6utUMKg4uDqK2gCG/AZ12FTYVccE3KM33icJfzfjNqnQKMhBZ7wKtzYeMNk
4i/MiBPViVDv1Y1oGtJWC5FxQpVvrSJRRhN0RileCUJyWcMDWxJLwu60Kq1bxbAuekVwsKG7fy3M
/DzeCO4EBi2SJIkcVpZseQ+Kk+zvWd7HOHOLR7cEP+eBAgi70vve9grxoAdGKkVomY6mkuOv9RHF
Q6h+RZyPbe+QQA7bOqM6FUYI9I0Y7U7oiW0JM7CfKFXkRBCt44c8OvfZRZJItsCDg8m8C81C9deT
zwAe+19doPFBg6N2du0cIePpe4PO1bDwHMbQ1jrXtQ9R21RGOyTd7WURB6QrMn299No2UYG+ubQh
T6zaoqYXgMJOabbKbD8UTHe7lMgXqaqjVGE/QFJSMNeQ8VujWWHGRWQVIZb6fuIgdVFrOSp/NBK8
H8ZoJOGbOHK3R7ay57xvlZNzjXjLs6cnCzG+zk0lm4YHjbFqNkbbszhCVpy1/jFDA+Ur7HlmnAFw
zo8Dtfjuivg/w4S5kRmmjQdBKmfepwJfVyvhThLWRssD28yH4QnN3BSZ2nV7+tR5iiTZldKMb7zj
zHGAyOAa2vt1wHmp5zcQXOlJvD3XLRi/IRT436Ej3tAnvRiSNXu762kBtSHvsMiqICmNov1z3Erw
Na75tSiFH8O9QYXbm9syOj5WoJKoXtlT8lwx6OG2kEUcb94cCRDdhcjvSFKApb29ucfEbtc9p/FY
/iSqHD328E5qu3jR5DbMNRo/GDwqHk6dI9Y9U9ZWh+LfYsgJEne3tNj72/f1Sy8Sizt3GCkAyVse
4RhD/7FBqtVroPxALrm+oo8t8GstP4YJA4s4+FPbn/rcL9oSm+H03QGLmIN1Yh2kCOTnb4ZdPWp9
ZauaFHBlycXHM34pZYO+AztK7zGBwHJWXwOXkYOeWvykI6TWF5GKSkO9VzCCa/t1PM/HRB3T184o
rmz7ACdEaL/ypiYGWB11DAwWUo7g/cOEgVByTCqsymENkS10eM22XIsWdgxDPIKvb6r6p0blzdYK
di/MVCDa7KWJJxEfkms1aDgyxxbqXFN0IRFDqgFGOikZbgTsOhdAZHo6S1dAAK/JUrjNg5DmvTAo
oxolQ4IvoUbGTYi5G1LcbDm/tLOT++xyv0cQ4tniXD3kCzgbo+XqC1Vn2GpvfqIfo9B+pz7MRdzt
AI7/zhn7YMvdHHA7MKShzb1bPbl8tNHQl4t41qQ2gnbw3pnmg3MiezP/6NDTBTByBDAZyoMrKqCX
MSJc1iAk1YbiQqy+mZtS1a5/UpxmjTlGwoI6whM4MgTMdNPyOel586Ke3CBUyEVgUXOyHN2W6AaW
tCszxSpwu+Km5P4yva98b9ybVSRbu1eQO5zlxzjfLRHPxG/mDHF68I2qkNVCZHuZz3Kyv6xzHee6
ctydx4f+qT44JuV1Nb3MvEngvQkSYELGuHkK3qYQlV0skFGqRZIZ/D8cbR0oNfJLhT3mC9VyHpcb
ncV2FdPo09sHj5R2pJ2UTp7AxU6hUza+gM0ec4Hk9KTUXSq+o8R6KIrqZpfNMQpoFrltVxnSHwz8
jNWKt/xfnA+N+1Vh0vn6ZJkSWFdEwX2hPhwKjKtZHODlMPQRojbIJ9EX3m/OBtN0BwjCyTeyn1sF
PrZ9ibO9QJgKWuBuVksGQRWTbSNnuuSV1HsU85DilYCL3FAJVhe4RHznKyH9zJ8wnZj1RrR7tF5i
DBzpuuSXtgj5L19yk007mbNe/DnnmmiMcZ7zjaEWib7BVSpak9lmyxPqWna3nmZGQRvRlGZHAGV6
WFSMTt1ZEqfonuOJIvHbGvTNpH94SaF4nbwhj/TOb+0yBFcA5CS0bnSbT/lgp1WHQ1NZQueLWO73
FObD7NO9JyFCEYC8qz9RhLXF/N2wwudzz2CPFRhPM7Xa0UbtU9yzpKaD2Q+17wGbNoQVI2I5eIVE
o/3TDerLimubBr7tsm14iFM7096bspObBYp1PgEnz+X4j9lP3+RUUzLEe/mJfBuiEtxP8uixP8Mn
ocicH7WvUlTV34q6ndQ+Q1if58+MkogXVPCEvmUMd2bEikScEiaSkHfLokC7K8Md6VLiS+JmmU6+
osJFpJtez2DWEOxLWAzl9v5yEFOCc30GqyFkhkCKc383RURY/ozQi+qc2yYx51ib9Gg72Gtkm5Zo
GQYwP7wrLLWrE3TfwvFCZjZNXSqcVBWJogQy14JRy3DHXfPXB0atwoaePA+CYalgdF8J9VBlqtww
pD0BhCYv4XWBMVZUt4eJEK37kbFCqgu3sdOgQInasZ8f/QceGNVFXEj4S15D+gOeh1vQv/ac0Bgt
m/H3jCsX2MtLiFph2s4BTF4UDwkM4dYLnTXo/3u/PGHw/j3M2Zms+Jhu+jsxJ+LAQiv+QvBWDPip
nVqI+/rqraApDlUPj8KoARmUd7qCGJqw6HElDG0BwiZPqAhfFb5IaSUpihkCY4e6mtv44uBXjpEP
RC6NmqGyn9VZQ1hl/zNJyVB4vlpBR9NkX7xrzk2f4AxeLELe1Zrq98jLkGCCc7CWvhmxcOI6ND1V
OwS//FZ+KAcceABcEA44XS3ATUQ8iPHUwswxuhJNrTg5bhTH1uV66ALsV92M3eCksOjNuFUq9NDu
FviZCRbNKD2UqaxhLgANvTRVL807dQXPEk+209/VAFRG+vxZNYfRB9Ldu4mV1tqj4gIrGF89Cz/4
IMPcZg1ht5znBFfUkTlHc0LPwKuOQpE52If6E7sNdX3c8EJnw7zV1ZGh/wyl+tZxKI/At1WM0euT
nRtMrZxob1gvLjPiXtPENHgSBVEboJut9/LrxIoNZ/tS8xrXE+I9A0tS/X5oO4kw0EP92Guoq4P4
cWV9xs6Qciy88zRgn3QfPAc0SWNGXRp+7jg/j82wQs4iSFYbpwIZjmvexfLSgliDp1OO7j5bW2Jb
HbKvLGLX3Z+H11nrm5y/LUw2B6Gfq1/5JXoYfaanb8yZtqmcm2XZulTbTUf4sAHYise4Fqip1UzK
OOBGc7rL5LuOBw+d2ECZeE4ekVnFzNXugZhqKa/IEym9kfkaopedo+xQbplrEMR0I1us9g9+5X/l
fMWw33HipPNfSp9agyIcnE5bZ0w0ZT0WnQaGfSYLJmURPB9cwhYmHh+zq4ZthjK+ZdigY/7IMpoN
Z/9SiD3S3e4LdpajQvGi5v01hHxzBYdfhhfiGGoVvvrUWxdTkiZCm3WVmqT6fOiyyCJRAJRVP43i
mdf71cCxORS4frQHWwAdPvS0cdZa4I9duS58KmL+ByF001fGtuWm2DxLcnP2BLmuAFWZKfejM3VS
fxn/fXOW7eBXytR0Ufru1JX0iM9yN/K3x+OzAtt8ZmXP2bHY5rMX++Ua6jFVNFkbrPpuLipmUWG5
iZ2SRZUuVkHErMC5iZxF0Cum9W6HYz0AcL6odoS/ZICPRoA6Xqg7Teb8++0dRqDCXyLCEhry6amV
m6Zru+XvsAWsjxl6Vg63J/nzG4og1g6Iry4/AuUIk7DBrEfj0mQjp0Dni1Yb/bFatflECnYbfoyA
U26WWWSOtoxRbFSoj+TF9bOGxn2zU1wgksMoE1XOELcafDlI6uKfWtJ4ddFJDdPLbTkM8AajQXgl
MCmReHJniLDhsNxagd/rIWJAmvtqUZitfygibFwyLAgTgFphgw3Nl7voUHJqC705FWMcwQYOzGNS
OUeM0I+7U5F/A4/k6JyM6aX+D6tmkyR6mUTeDt8Ixqt6WQ7UZH16h/upp+860Z6k4kmdqOcGG+dA
+ChcN/q2FlKjKJj41zKaEmKUicAGMIJdm2NN3Ro+QNfwYB3TJwWz+1dVRhkT6NtAa0sfdXtNZXXK
IjpRoz8E043+oGSZGprI2BcGpEFpkMCwqUTVkOAZjBTAoJ0z6IMBmf5z9vg9ALI53QkSp3b9Cp1K
Z+vaB0m6l39PBz6fZi1rqtjwHlSHGN1ExXy9VAKkcaIuzaZG0l4vRFL0G7D9zr03DZdjH4SChOcz
BW+/wJ5tYBopiT3/kiQ7IMh+q9rRmfEY4/n5LujKOKw19qbsHjhlnWq3i8n+YwMvbtejkw==
`protect end_protected

