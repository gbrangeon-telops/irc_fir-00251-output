

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dwCKj5yWv0+IePBqJHT08eVU+DwkTeU5oOrKTCm5D5dLE5fjKonyT8s7ehOuYqmaU7hbrj8cK+dG
v6Hkf9vaEw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofPimz6qWDPfdZmLTvO15AJD3qAYPdAcnxW7u3A5HKCVeJi1plo2JwW0CBkFgjSMPqG4mB4Hkwjh
aser6hfQcfNXvJ3JUWr5ZS6ezr5tSrAVnAOcpabYJ2vlFEce3rPTiHxnx3vwSLvA9frZJO+K8rqA
zTaVjBo7aLNhP54LcX8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xVx1mMvfUwlXTa88EF8IX42tnG0cXSGFt8ROQqT5GxjYzkciIVjF2lg5N/iujDWrU+m+Hq1jVN/S
7L9ZrnRgKz1GFQOxHGVlrNSRcf8Ej88lKuK02N1SzF4b1/VUH6ht92N2p/ROW4dBYnWVBpIxhF08
xg1QHd1cs9lodA6VBrB5Eo1G6aluz2m9EBGHigHdWN9RnmtH4Lso1/y7QElbZq3E4/diAxIYh9aF
1JcFvli+iX9S3ENdEluRyVweVryo5jTYqJabkRWFuo9iOs/Ic616lgSVONZ4NUl4ItIqkTq/gP0J
z13d7iJ5zyP7sku49PKKDfaHMGhWx7ug9eg68A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mm3ysnbGmWPGigjf3cW3nqCJ7td02DMWAwGM3y8Ir0JjWwms2hUSloczYrXXwus0KFJrOvbcp8EI
afa1rxF5AlIKiPd5moyH7qLa6s40f+FTseHQnAhUIfuaGWVSTafXnP1rMlydXotX0OgXaf8ss8Rn
aesy7+qw+4loCzosrzM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quGvQtw6SKSqCyA6Sp/eeM9Ow8TS12WLAPu5jebLdqM/ryW0A17A8N0thkaJZco15r7Owh4nFU5l
KZcrcDhvn1UKmGv+3eWd84UW4QDpY80dJTTq1XGSt54iFPTL0Mo21C1hbrKXm36H71Xi6xWsaAlk
nLsOCKMEHsujeF1naPb1xFZWSlnfCp9K2SB7wEzz8xUdktOS4rqm8CvHN3HMePG4N3SsN68l6nRq
sed/9GKEvYzA04tbQb5NASiphn6udoZq4W1cZDMS1xzdJ8v00rtDdh9Iinn05spY0CrdzbMqalEN
NkRAqp28PSG9/FiSfEP/QtuVq+XzCkevSe/NZA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 83872)
`protect data_block
wWaRatsf42xkCO34Zy6jgix9A9KQv2cG7NUoklNo7t7kK7qpXy14A+XjzxQ3Kwoh7MYQzDy9XhXJ
nxzIbbTDkUolrgpMtBJ8h5k7RbVgw0jOsetv8g3n59ff5BLMk50kEXEYr6IG4Xq3SfwFffVTyOOy
qU1PHZt3yS0pVPJchKOCQCxZXPZ+2Nz1vz9YN8g323uNxTFVr7Fzg0jAazMMZe4W+3NN2xgIIbO3
uALX7XF2eYEjrDrfhBS6+1lnI/rf0kp1Y5EM8NEkuChcQ76kHsYpeh82s9yyAoBv3RnCWjCN58Kl
Ofloz30ZTnONA/qe7WZPKBU7e5vA6uf/vnsdrchYMwTH520LpIKTyZOrTjxZGVSc/+hi8BZlTQZO
int3SA6AE3Xt1hDid59WnGuYy5VT/LCGaDgTPMq5tAEOCl//u5FFlrBNUme63Wf95CyhaF9Egyzu
YbcXeo+gi+QV/51taBpPHy45FxU9v/izGDLTErJReMFPYZ4lyYKHZUmcUGodh16R9MtrtaDGyH/w
8Isuum+U7DQP2Yxlk/LhNHh5DwxJMTi9hjVRZlbXnM3skdKpj44oQ1eQa7MODRjs8xwyyieOFP6U
4UyoXvP/W9ClddS87Fw+XFiKkZBksG45rAImif61v2xv8wR1CKLgmjJxRy6ruVZfEC2NklV7NfbT
auj22RiY2841ciHgfMSWoZVZoVvtFM8012aD8Ar5LaIi/bouvFQ3faZgHg2Cp/RcSuuQnqV/8YB8
GVh8LA3AS2IiCI/hVJXln7mFaXj0fpITbIEbhSyPaEUeMpStvzODH9IrpmtghrxRKs2bOycZbMID
FTLC6+VbOZhEQELoe3zp6famfScfZKhZFCBAGq9r+K1p3aJxwT8edUp+cO8cArcfejTGlSeBhMbs
QzfwJ8vbkKWQSdI7gEh/PA5E0X/VtB6gdLkNBfEV9YW8u2KHv4TZkIH2kojBGTtjZdfi8jxJqwu9
BtVGB+oYSlr6il7ANfowjNTfZ9yO9x3ga5fGwJJff8KZJJgAKzBD1m9tY9hTWes7A2WWCVFITPO2
ViL/pPRSvR/dI6YFcobXIARp75X2KHN4rZXVQqecaeDJQ2Oc5BCGXCSt97TQSIqZotTh50e9WmY6
wlNAEYYR00PDlSd9NY+9ShsoFSXvi6xGL4j/8HdblLDyOHKkBeL2aGDP7FsIpR0aKOx0CzZjnkY+
dUf7Wr1CwbY1nj5fm0sykryh0rvTdG+HhFxAkLfx33+T3ChoZv5fUhlruxavakkXccxu1SjRxMrM
cU8kwS3IQKD+QXPWi62ZOYZS9Ql/GmwankWqgdrs82/gG/gFimMsuvxTYEWP1UozuHxQ6Iqwmam/
OdqBFOKUkOSPR+nYGhY3uXwNQOBnk2h2xSHrKannaXm7ft7K9/ifc6lbe5vaCbLrtZvzTulLfaRW
FF6n4rzlWvyVJYxx81LLkGSdatyvPduTyzzRClrpMOOxVv6gbtKCOKfhzy6Jiprp8ZdBM301TD8+
QEDIwUfTl7pXOniwJm8H73j+N2pDwIRNvCBzirPPyVnr6nEef6BKXUgcKP0/0Z7FvHcAaFzto7l2
PaBS7IAjVPlN2Nl5PXYYASHA8m6Ncg2ntqZ8vQLOw82EJdIm+220YxD/hLVh3Ev5QsCE9Wo8/wGS
x0+pbjKpauYtSrHo05OsjLUEWo6pyTbDCEENX6JmWYOZdfz10A5j0Nfz//YzcjuO75WUxRyncrYT
e760b2DShvQF0o838MZU+2uIcz/klIpmSLtXecxYgJHM4cqczBxltC51aP2bJqpaWLTjvgQGwBrl
8kOWYvGAc5H7fBtN7C9ib/HtHadlWxpZQGoYSHY1M0TOCvh9LE6WrWConav7pdywvdmw/gm2dZaz
3PhlgP7Uk17pe512YtMDV5iIy4afnPJj/5kN/ZVvC4sJoioPOxbvIv5L8uU9x7DnJMylhdMQxjxT
uN+J3+drIBrfkd9c+PnNqm1sZ6/JO5+iqEjVWs5UlySgJoRvSb27fgZJb3x6RG8iwXkpRdIbcs7Z
Vl/+Igw4w5ph9CNEDxgEo55ohYSw67Mx0I2yZtL2M5HZm2PPObuZ6tCOFrRIyPyzqLoaZhtNipYr
ijvhnAuHwuuNmU44uyeQ6EsWlUiUP+lGjOduvMvc1fu+38Md+C9R6CacWuxu5NPKW4grGleWLk/3
NZjvDuUUqPn81sFJ9D2QY42korMT7J08X7IeB4IN4g5Akf17avVBp/p6cxv/NFhBl36iP5goQmg8
6ZIukZO0PdUEZ2SaAjn+6G4CzScQVvNrzDzWJXXty22EtwRW0V1KE8pJE9n342vIy5JAQYlGot/g
Nm5MUhIlfivkDplbUat7Jxh+L9z8D40HOG+kn8tjCCKVHfGyesNB7i+cFS9hX1JCxRVtXJ6L+hg0
ojijyUQQ0duMdDCo6YrbTt0yuDLwctq7HzIiXHJGuuiwFZ0e7aGh/5JKkc36va4zFVPi5NA5nQY7
D0rK34RFD90zbG8YGpHZGsCD8kN5R2Jy3XX2jljePhepPMro5IVW13SlIx+o3M/2xuxW5Sk5tFw+
khmYF345yvUpEkBNDndVyx5roQSIWo9ogc57xio0eOTKUVN+TuwtdFijcPOJ2c/jK97MyEAj6zJR
jQ0txkFw3ovI/2KF9AxyylkpnCSW9ylrg3TnadYZ+ZyiLvmESK3g+K0i2Mx+7h6yFYRnhNcj1cEX
vdx67aYfq4C5XSQ7WOlGR07Aj2EcC17CiZCb1YpHZ5biMUE35fhjfiN51BtImShVWakFVHxZNyAg
yXQU1uPR8WA/R46ss8HfCm7IbSRooNIBfVZYqWgIWGbeWKbbZruqWlCHMxFREI3i1tNKkc4xFLDl
HIvisJ72B+9X/326djAqzXMCfbqUcfeWJ58QySvVsAocTKvvUS5UuEa9GWeg9pNKMAAHcgagnO90
HXz2SfKBeiGQ68eka+Jf1rdzRCVFBoYXKJD+iDiMo1vod/wf001/jVfQaJDxWqX2nBnW2eaQgYX/
sDXZa2uCs9Lj27ftv93ZiN3NafGxvgHdn1KLPtSNFhQsiZedXxSh0yng5mnxilpThIDlKRzOwDeZ
Ww4h8QYdcqqbMZQYK2r8tuStJkd8EoqLcUG9V0pbUP2G5pHaztnZXnw9jHKm10SIk9wSDFBjUL2+
dCmQrhxZuCu749AARfgO5B9kBi7DogmVSF2WnvNRWy7kdf6cY5LJ/+BZ1j7rVpnVuoorlKBr1aSm
pcEOWs51U9iGJ8MMsFxafWnFZvkjaygiGCYyKVm7c9dT6nnDBoLmo+eGUFmUOgqwxdDmDhqoTEjU
QxDz82mtLrsdY3g+Iq3xdUUl6Yl2JD1X0Ta2SLpbywJdetVynf26+l19D3XDgUow0IR+dEFdwLQM
pwHzczjpMujSaPOPaJGkYRX0nClSeJOoNVv8XNprEi7p7QjXI6skXJI66BgfAVVKY/mju0ACN6Sr
AyxO3tC+yJEjwOgHDFwu/C5PRCYyPxT5Q7xJK7I3xS3e6UHJpotmG9RMcY+q4OpiJPhnahofsJCz
Zl8jdYJN9P49bwQ8/h+Rmnr1w+GDpojlP4Swz2r8w9YKXAs4kmkQzmX9HW/2yLqzu8Op4j9FqSNz
Lw03Hl6JjLso2qtRpGToI9anUnchAZ0LHrTRozKHL1M4Y0ollQjUgiKW1GBp+61pb5zcPySh24dY
3XHJ0qQ2R9ytDdxSwhq6iouAXy2yFtY2CoZBAKkCd8U/SkZ+iSaq5h+KLFI9xzsM6BCmggcMp0Uj
0PCcS5OQ1XGSlS+oRfFTBOj4DdWUnOZSrt0G9+t667xUXgsjMD7diqUaXy42VNbohALhMDv4eY+W
1IJmnODIrEqQCJrpBqOKTWO+TQjYZbhGwsULP86T+y6qSEhImtrDnJapHDnqF2kn1YjHzOYQNpn+
bsxB7pOfmXlIL1wGQeQp8mJZE17Fwu+JeR90UbcoExeV7Vz+YIvRMQEOh1koGFPykWAZ3ULdgki3
o8j4DE6dmf/5p+np4Srt41uFXwwcG8Rg0iE4ESXKruqNsKsjq4dfPioJzohFMtiekT4eQQE2dRWT
Puo8S7pQkQfKzxRcmlzCVS9neHm4yWlIJRX6o98Q5vwGN53mVtqoSzQyzm5kXf7OC160o40wMAPE
mHn8S8FAfZ82/JAnnro01roTQ8a8phjDhVgnmYD+sqIc+huCP/UH4eSWIf5RIaTroZTBDtsY6tW5
hBPphfPV1tvK5xMDWG5ORYPGcRdHjAWqNCjuGRDeSgh52ACDDDhz4hrPaZm3ShWBxJGpyJLOKI/F
6CkdUD7fNlJ5tp60PyidbhFyIa8hA1NNAW6BxnEQcv7Q0xyDd1Dj9eDFar4eCkGGsk/YkQ1R8e/2
B/q1rsIjJVlmtzJYD4qPNqenEYS+aCgK+dmOmxch+RrkPZyPTX1YMbg/VF5Kuo2yvkVWQ08DTIa8
ivn/JHBJJas3rxfhY3EBjPg3hvWtqbztFRZYk15rW7TofStTaT60tDwjqC0GWrzGJOS3aj0cXeR9
sm863KnEl9+RPpoop2pOmwRo0ejedjfMuoervJHkCR3dV/REQ/pSVMMWivEE9wEpnAZXKy/PUXSJ
W7Qp1TwF6S4Wgyfo95G2dMXVjMVQUoDerW74wgOj9spLRuIC3bFBVq+l905dnrG25IefhQuzggl7
ymyQNCTb40wUKBIoQItb3ChxwxpJgm0M8/iHvhD3Ye9L2lqaqdyMAAMBwVyOQyIo07u5CjZJAbHv
+zOmt7wr5KQI5kiPGex0EjYTIkW5av+i2pvuwrVqmzAA5J3o1KMiO3IDrHpSOclSjgpVUzRcsr8m
FSXZJlySAs3vAIYlmFEsv/gIoI57G11WxOULgjJOEbc+X7eQXdqqUGVGOnYML8TiFI2bYNE4MVMN
FJ2TtsZcwnEn/cnFbvWS7mmqYsFgimQwE62PuH65Kf+sg6cuMctPPZO4pTQWEt5kC6owFPbL0DF/
UkSrz2ILV8njTzD47l798PFluf0WSuAq7Tyrlwbyrq+Di5LGELp8ZKBax7Wy4QSL6LASuX03yyMY
iURodfKpgPPUvj8PIyh/Tg8EUxEYfgGOeNaYJ+tYbIrc1eaeeiHABnoAEqoskkzuth/KwdLlfKjj
mje4Ag7WOOuNOKo9maX9G5zskZ9+YpjGiIybotrxiHfAERrt6SyEwbk9cUqL6KTHMU56aE8dEBOl
G81WY5pRKvamj9nQxe38F6xpiLLwrg+jAVyc7o90M/5UNugx8jh2xIOcSC8RSKGKTTD/n7oVmKx1
MKITjlMigHCMumIf9lJpyj9fEgmIUAkQi9DBgeYNhNQaYmCcLi0D/HnlBQo+Nas6PcSMFpJYq8Ie
H0zdhOd4f+nX84ntNf3/If0kP5QYQi/iX94eaTsFgTbQkQfV9Fpm83HsX61IpfwGyLhwi3SONwJx
WCh9WLIVXXUgZ0y2I8Tvu+dO/qdTLf8TPtTd3I4eLnIBuBzDcvxm2jxUPunIdPCDmpfQQ1uWidZu
z6jwFMhOuZuricvj6Yyi57be3JAcyOhneTeDAlyw61uoQHFOlKiKO95lI0CIP8i/u1I8wkMI4crF
KVKx+NqmizjBkesudvbWLXXZWICBE58r4QqjtsYapl4A5KqD+I9F28Lb8YJoMaA1YINT9R+5GE3b
j7bVHhKHYucMsOCo9kBZZHEd+wPo3haDgs6/pz4/EUVSBTvVErJxwT2SV0gqXbXYwIBj+Athu0NO
dx0F8s1jHdhrdfCotiBv3mhpsrwDx9HtJZk7UUyHE9WaN3BOIHdRQ9vgFubAEuplcQOZLnhOKunN
bg/inVKtOZA7ikaPwn08CRQEbM+KaLJ5+TluqfOO6QaIbR36wb/WWtvrUUmYzPCQWj8zmqO8FbjM
ZNCsDIdb3L8v7XPgR6hKvcaERaJ+VPnERhkYonw7F0PKOzyb2PU7zZsEg6raucrgn5PFjoPeb5g+
v05tUgs58scsnn4Wl9RWAapuuvIx5dmHy2n095iOaLmucy15czBqGz/jlE8A+9M8WMPVEnShezBI
yY0GRjuDF+Jt1AB9ZrOYuIT9cuJZDk8z7ibQD5Gi71aMtQB9mCIF/lYfeQMOXY0BZ7Xz5rO+ZTMc
3B49wU0inTgrgavVX+hPpEAqIqbBXW0YnIjpwKFhoSuNjyMPfY217G0K7iVFBMcnhArICDTjbQ5G
lRHaic+EqTQPbTYntYFuw9MkeK1Ydt4Y7voV0aHCNa+LTitgrj00/WbZt4X/TfEbk47ltFgmMlHv
Nau3u46NPHZg7PgOpN+wRzVaJrk+Q1dNAoVzhLlUb8ExlFtoWOAsm6PaILmBYDZzRzhHRE0D/L7H
Zpay0zljM5k5dHTyZTW9uDWlWN9Uyni4yLSrRbbiW8FEE8hK6ILRHcwwE3y10h+0zs4s6/xs9oUn
pcNnwqQKsUCfeJlpxZMTmAGucBxRLMBAAwpv4jCKemhkhRzw5yjUgErO8pFcc+otPqLsP+0KyZJm
L+fopfZip26vPOBTyl5No3FytrgL+grY4jLziRu8mzMwue8ngzniUPJYGESjqTg46NKMpqRQqvU5
bSwEUVyZbxf3UpTFk7T0q8ctrA+c0oUFwtBwUF8BC9mLf3S4EoBJqJcWdCnZsKouTHpUCBUdRP1l
5/BcZRhbucK4zBXZ0Qx4o6amfMP5AXsFH6wEDReOMVEK9rEuH6Odl0hU//dfBKLerrAMOs/Sr3tj
9KOLOsfSF702FxFK7tC/ta9trnpYHmj6Dw0E+zc/bk5J1boFOl4tdh6kn4hjlKTKszcM2Mq6w73l
ImpGqwraRej7T5r0i/nmN9Dro+qX3xpz3OI8o8qmfgWE0bC/x14oaJe0FKwsDpNWUyNFFUXEo7TB
tJy2zb9meyWRUjgpaHaRXdN9i9g4Bny4LxI0ea+E+u7jhApYRxazNOSVASz1hv93h9ISwJiRzlnP
C6s7t2i4/ywpU3Ranz2FRjRuAXZhMlHsgdxtsR3Ji9PBkXgWng+n3aSzvLTxvCvz4K5y06Rmzmsq
P5iATm03Cjq/tfGu/m48c5Kn4MrCdYmi9alokf0JuBVFSluvA7FIQpf7gp+UT/Hsanb/Wzh8Fm33
e6nr+geMFP/lF3S5SMpGBdgsl2tO46BEgz4qcNP6vnXdU/tRaRHHIFZqnGEu231jXCFFKiYFsNlR
5IZe75rApHxgUT00nG/xp6HTxv9yGJiT3u9zFB5atZqQ1pXF0N99n/KYiGqkBtZckCxrfOu0mO73
Q29GNg23QlBa8t0ix4YfbI0n4q5BMIbcHIE/xjuKBqpLxeuOWtmwpbIshFPsyUoQWdTFaMZJtLMn
0XXpf4T8qw1I4PlvMPl6TTwA5PElPIjbIzCbUH0ub9hKMxkFCwxfC1OVS9wG5HYiwN4e1i7mwk30
LIILgP6XHNQVj2MLTKljyuLtv9OrEb+2N53+8jMW6WJ3btShHZ3jQ972wTDBXBDH2cy2rvqwRpc0
J4vZicCOGfZ333pqGtfQe5LCUvm1kggmmQWcgUlDOy/050AivzHEWsWUmJCz9HhRYz7j0YwaTFDW
AHuGTHlhj0FoEv5HyARUIrq08zxLXRh6I1vSv4PECmAmkh+rS7vxoaSnBsWLYTm0JkO9+9IxGVMn
SxWuHu7nDEZdGLuK5sTF8/Zq/mKDcem03OQLO02J1PdS/RP8qk0o4FLDYaNdunYGBVvDh5lVkhyV
aP8p3/i8qB2yyFLuO1XdPAbZmT3+xf+2YnayUs98IxVDKPN33ZqSH1gcOEIur8kJh4PHIyFLM58I
llW6Ej9plDxCngl+T0HM8DhyzUNhLep4y/FX2MSCIXatvLC0ox5XUb/ec033pAJIx/w4Q1xxwc+a
CcnrgwYF1MpL8kCByAURk6exaerL4UJwTqo6qPdyXOMXO2gDqMkDMn/0EGjbv8wJiW+6xeL1A8jb
FZXrhtye6VkcFzSBwErR3CN2kR1ZV4NpMT6ZC8GulsY4FOg9nfxEr2pzlcPTsZKYuaApJA3Aq5fY
rbrRSEUBczm1jM8ChbCD6Cpl55cSqu+/2pjCzItdHtCG3Z3+XOWLnvilV7GgekIh/PFcBz6DecY7
TSsUDtMFq32rrq7W3QoUai/bV8GiBXSzPDB0MSL5ahMOFwWzrawM9v7CkNb0/8DMQgr4UnN6uWnj
uTu6NFMl0WieXvwfrHBwwSCF9PIW/TB8OMHBUOw8qW90B/NjKkg3ErQo895whScEgl4i0sVWdB96
LZPC9bHkCmnP3bEs1GLAdNq459lCjvzN4loVzI0UZUpkDGTTUuPvlq7G4QqyWeEEAGwtXIjEmNWp
UmRHt5vkR0eVenjTPdaOKoSja+YAKd3PKVFAYQcRSR78jNd8DeLAMgZi1YROT2kNncv7PNAwWmmu
Pe2jlfcUn/nAO/g1CrH57B0J/wRc60kRc9kICIwXkFRrg+KFCAY0/smislmuXJAUdvRZkom4cVWN
tCqRET/h3gDqlpLjIpPidRzpbDI6aEj5SZCx5ZEJP/j/wuXI8o/aWWu4SS1SzigFhfr9Yrq+lZc0
v8aVmLttyKImX1UdvkKRE4biNmNYYyp4g1241KuV+HRYeuRXrSm+sQQonchXaeHcvBDSFxv7uENZ
NTfMgGZtPeL2te2cQd6JjhmVXJAIP4tueVQSAaFLusi/h+EB5orBcsPu4zgtii0oG9rSWxiadykX
nYunQmfAocT6qeufqdlnjOieD6TCAxeuHR5oiahMo8cRrtQMkQHYno2aLlnRB/WoRtUKWXrtR/uC
36u9WlfRvGlPJcWeIZvX5Qr0ty//ipZ4XlZwDYFmG9T4Qde7NDuxnPz5ih9ZdgOPIzZWOW3p9xKq
jRXUFp6HnoXPPRjv/ci5Xh1vXay5TLla681nUvXHO4Q+ycdNH5F4dsNyc3D3Nz5wchfhoB3VLG7l
Pmz6KR8TCRKl4s1viXqYN9gApF+gQUpdNEaxvVTIiuHULwTrEYVT1rIjiA3v0b+DW04pld/JpF33
689sE5SAQ/FEhIArNCO0Ya2ZiKHJxoQjjuPuc38f4H+6pXnCYycKhnMvSpJZr9JfRUVjGTLdNN4v
Ifkgm1LMT40U1M9xagcSyOCnXD8RU5NDdpxeDdCmch4Eqem9tMRHQM35cYUuu5LfLSFqrdg76Xfv
KTTQGfSvgMmn1iyVpaFTDT2cHcBmc+V6RNkS03i4viLluzFLToezVkPJpHBatHxNm7wDMVN1tdAG
SGVCw0l4a26NxpjCTPcrrKnuU3T/kJ8nxGwiCxjcivA+VkhpG00WeptlHtQwlknb2YAdOWlByQUA
ZIRb3WJPpbkGbFa8907i+7yLbB8A2vJGP6cvclNJCPBGiqK8R4d4uUBeE2tf7tqGlJLo0uOksoQs
OSudNaPqQHno7yGvArpZXgAYyMvrnAlzFUut6XUdhrc0XC3lP980CzJp0rLH4Yy0biJ7zJsSB3JK
TotkpTz5MOvb5NawLqvbToaCHwCakWFgUy9sKtnVR5W8s27xn2CKe024tfLbXh4Qrer0S53QtCDY
8x+VPYAc5Ga4uYpg0O49jhWMWo59JKONvFntEOpyNCNRvmKrkY+v1vGiIxY9jepeBZEyuFoc/puM
6vFp2SfzlgWiV2UQZIhizdDoJTyk+nst9eH+kVh456ywzwRMfW+JsbE3x2uQWuYtZ8pfgycq8HrQ
armwYmkQaUzt/zJGLwRXPiDRmRbrwHidpHuz2weErZ3+S+1vi+aTkuJEpZPVRLAanSniTWS79eDY
tBpQnjGxQr6fzqYrfvrNXHFtwV9mL8oWVOhAeMT/GOHG3zqxW0kGjLnmsltSoZTyPqNMrJZ6n6gp
d8kr1q3ovuGUUQG3leD5Er6s0m/P5j+jbgC8MJOhhZZBYPU3ZQQgN/6iHtG0UhWDlyyEh6I9QaL7
EcrQxbzKACvOR8P3O14/QS+BrXePXokQUhmbfxWkiMG2BjtlxT1P6ODgW9PrlSL0ZhUVZBBDEemW
EXJwefgygygcW+DM69Cq7fFfHXsNqpQaivTKMO5rChDJ/MdiEaTWgX28dsL5FLWwme3BEG1kmeU5
F7cs7Mm1xmuOlHr8pIfLbuV3QH7gAnIQVpx+RuGiJrILgAUYyCHV1LhSucO+YAI+ADap8GrSKdcM
NxwVvRRamnvH4AjZqfVA6GQHiigNqW/DiWvlh2Ch2hNFYaVEttzsCc0Vf8aPVuMFvAmCbl++fttE
1zI0QoJqnfy6jY155xMi5KqG7tgyUWY6p6MjaiCSfinpfOCHCUI0zVVJJf/NLdHXcVuxAM407I4V
e3UP46y0iNTQKiF1PQCUTs89bX/Qs4rZJJw83TMw9Q4Xii0yTq4dosyVZ7vVKpG8mBnBj0TWCV5Y
Q+wiA1rEzUGDKjFHAlw/gYClycVVi4U/pRIqcuNDlwvYArRQV2xjxA52xvE7DdPYqqN38R9+bSVP
yk9MpyVRTrGy0gCoI3Y3KtMnPwibHQPatKgSJG34IpRMRFXg3QHkAK0ZxUqd+sxWIeG2kyYk/QRQ
V6j/IRveJCJVxw5fBGOrthjE5UZkFpmyinRJxtpOFZDDpjoCJQ70t/bs3qcEYTi88HPVhp3RbyvC
FIkQ0IvfaTyqQBZ/x6xepRvhDDrwA3mlBHRXHvvWpWGNAcRPlNiT+VQwFxIXISpokmTOhH5/BmsG
SC64UT1v0JwVr2mi8fvVA1tiY7nHV6nkxyuwndwx3Hpj9/qn3GIWqCyjs3jAdn+IfXFRrWQLQjJF
NmIVwQTNAWMr94L0eFPwBze2rUHXJVIpKMkD5meKW2rc1orkAC4pjnxayyTtmq7MH9NJhuu43KGK
3s9dcJv0HJ572/4rRyI2kQ0z0IuWNa85QgoT6nNE4/xo+SPU6mmYisPTs0dkdfbViUjLZovv1EDB
lbRBmBqiaR8GkZ+ITo1GqpY+KwcDYFXAG0Ot4ZhM4BnumG3Ng3MNhjG1qgsmc9Z1oxmFKXPDEpV8
QyFjz5mc/CgMNt6l71LwQF6VRird15KtXMMf4wtNIJrWqDEC+cUSnB0VY5WFbx/RzeUW3hX2CJ6J
5LbckcVJcYfcVMdvKy9EBx29Y6Js30fsF7r44MRgORhZvKJcwfogMcbajnOFTuidm7qNLu1y6Deu
4D/IZ0Q+9vP+ScuiLIM2/ygNR3ZleHK3xb4TswBgFJHISCSkfDm1G2hHK/+Y6ypvJWDOA/q+vnia
zqtuX3Nam8XF7KhdanvH6uDV633o7XDhrGGI/A8u8hcHWGDuD8tzizVnoc5Vzw2w/EBG0GL8TyqJ
YIs6YgkLC6B8jJaj4enluaQ74WVXE4F4Szvb7j7K/r1x1ZEiRKwHYkMVckukWKUFmJYsMPq4HJrN
oFkhjKTkqMuJxfGMtKRkzp3EDM9e8CQejwj/+E3bgghKKN+9Y722e7FU9yd1rY9qK/49y/JLvsU9
tFlGaL7mOOv+Zv3R3mgkDC+RegnWQnX/uBRHD+OClIgEbD/7Rm0SUdslWLCycl0zwNb3eXfDb5bv
YzqvyIBqIBBLNmKrRQwAsc4gZk9E0lK4pHqXYsO95PIiRQmV5+S4FU65MplErhtPIFuMrFT67bYH
dGD+5JiAxcL95Ua9cy+w1td9PODYlN2Jxd8FuRZN+WevDOkVs5YewNauBF3XBHd0qMz6ZhSm0oim
xJ/V5r2gIaFusIGiwMsUsgqD7Xu9ERui84DokbALMD23vsp79yqvtKwLAWNWN8CsQl6B/j+OqJTf
ZWbBEluKDmyre551Oy8QGO4UfnnezPMhYL0/9qNkOErr3GtDopMguVdfV03yxjUSMrAGMIqwsr+Z
efJQzR/ld6hh09ROGxDTzupprzxyLVLAcvZOn8LheV6oXktJoSY5VBAOiJ+EcpJUvr/oFJdpt6e1
xC+9gqpqoAoHBxuLBfCQp9QLKGTEBulovGKUdnDs2yPwfRLqI9+dO2W2miDYisduE7qjWWWLxApE
r28uTqijHwd1gnTsmA7PflPRUliRvRPKb9Vcd7G/lfot7qjgH3xQSj2IjfJ2xpax9oVZMcF61FPH
As50FISaNHjdVlOODEwVtJXB251IW7uSXm6305vMd5mBZw1BPePFGfpcG4Yecwhe4geQ1KpYiHzm
Nm3R5dL+frPPSLcamNh3fid3XOt9vhopVxXXEg8TOZdVI6vkxVv4i5/G2P7NazB9yQhjZ8hNkqyS
elmCrxl5vRvuxulnMzsXpdhvrZGmwMTDtZ33EUrMBhw0SM82q7sF2nOUQ1QI7UW7UVSqkmdtBVIH
SMy4XnZioTaD3NyHCt9T+WBzOxyejrIH1I+Yz+C69CyXJjRKrvzZRx9ZYln52eTnEBWZ1E7ObRoM
JonM/g7Xn9Z89jTjTgtSPMEROlyKauHTEehEeAwGbsTwYdjcIIHhnBDvgWv66NVcM11/y7Ie2cHq
mlgLBHJC7bbbT0zhdzOpt6Fzu9he8jdf30r3ffNq2xdUQaJgWCaC5Bje4KT3UBVxuH+EO4j89V4C
Q4yNk48snUF7WJff8ERD6fMMOwKF/Xcg0NH9eb7JlVztmhQ4nWhqfmrSM8t4rJ58LGFi3o8qMEio
s5OhzY6Jk0VTsZBeCt+mvh6kMMDKvAyJ+UoXn1/OTuY0fsmfX7Mh+ApG0LeTtyURfuV3iMDA0yST
SeQbfAHXQCo0BKHyaMu+tpS8TlaD0cep/KntT+vmZGeqmdx4maIWOIQqpKy35O7FhLeba+uSuUAG
eC2QE39CCaO+IpuyEBoc1jO9+bZiSWdSgyjB2RGBsA7Zjzo+3CPOYneoda7h4qv2F8DVrBNRtvMm
MBJ3jOOQITVY7HIH0LMyHPByWRmomOJsE+NmijDsEc6O+Zfd9WKv3htVqvZV8AZtpPBqe2xo7jOG
wgOfl/udvGMGwPmSsRs1CIfNo7fdsVsoMnxsCVmRlqvOGWzqIwgNbVmK5s7KDF588sjUUTWg3Xhi
2sj1H4vjl0Y2pM0zAQxfmTPfv32nfpOLCskdLfNZOGAXJ1X+YwraS9haHnolPnQys917npYwMarP
Y0keOkt5fnJ+wWDGNy+jhrGQmvjbarDkyR/jFR7EPrA4LaTZ132YqIuyrQKxENxKfhFqN4EWU35k
F3yz2+XMvMRr61JbQF2yvQPJBsWZNjvBL/6nvz9bgjmb/NPuoMe5oMJshX6Z7ZhEiJeb4084CaSy
QvQKOXVYZdXbhEGdeOI5ecn2M31KBC44UxK/sAl3YwqksKPqP/62iDn5/bt9Zhmox+q133ek7T1u
EOfqrNW8wiC6+lgm63m8gGFpvECyAg5Vza24C8ipT0zBkbG/k+Q72xhGPqQ+fGsqbrULSFKOf71I
oIFD4BAgx7zRuSitJ0heok9cSMouIYB/HB9m5gpUp0HpDZmjQjdtg/3fqLYihDvCEscY2dO7brmA
iabG/q7lr5/MhY/yEEqWUvoCq4MABK6y2n8J/1xyadYM3u0Pg5q86Ax3AGhEOIIhbbQl6EIgJQuR
HH4vKTjRulZRBtpBeNQtszCDs68ShGhpfApVSQv9pR/vfO2NXlw4bkguLSdZd2qTLRn1FE8+2Jsa
MhNkefbxYhO0kvBoDHUyUINKXt9R+9oUdulkgfWijx44Ag8NPhe2HRFnE+L4jtkWVFVXwx4Pao9D
yGy96mzxduQo2Cb4PIdBpSHTnpQJ+rpbSn9gmJZUBdBNtJA+xDwc2SjMCT0BLKB7iG7Y+mP7QQwp
3icmouHaja5MF5R8Q2F9LPTmsPvRRZsiJFqvPWjtY+Y9Ci11QPI7rcUG0HXZnbkQgO3Kspt1vFcj
QV24Kf/bql2Y/gNsVB29xdgrbd0ppUiJjlEa0IW52hbin8nKdDIrOvb1OgbEtkTmbduv+SadeAaF
ZhRXUdo1eT/hQ55Ux541CAOlicNO9aKhps+UNCpiWyQma2C+mzGzFKcZAWRuYs5saGH266RO1v3p
Ob4p7n/ST3A1aS2jbfxs6hLP3BzlTysS/YGjDqovons8WA2jSyRox/LfY6B5GBFQkVoWMMpY4qpH
yld8azgatuVt6jjNT0kCzM8/orA9slKbx8MKdYhw5D7Z7qMhgDhv3ViqP6IucRw73qFz26+wmyff
G8dFQJK8fgoYTx3xMqAPi/wlCHl3WFyihbMJ2SUg/aUGiH2UpltaRCLOrzk2nVcY2FQ4E9GBvf9g
i0VoKxYrlGrU8NLL+ni+jxKn9AfKKEreZ764R9bGM425wSv0m5hcA1k1QBfG8gl/BFtOt7QHri8H
LC+9kWNrgEERilydzQAgAUsjkfACeqSu8eZZpAxzPGiBCknJMQe/eyzFmOEq26EZFfobLQSkgHHU
kc0CLw5m2hytZv8R8lvhQIDJZCQhTrtkSlF6XvVWKomql/lJUWP7rONCQU9Egzn8tfNf94APVYWW
N6PvtsAJEqH7k8qTsiJ8Z+WcvG2wx8ETrY/g0nAkufSbo1zbVTdkxyrmo2G45y64hnJ+BukLBJ9P
wO9KmmYHp644f5ZrSVKOYZLauTBvIhalFhmwBYIvQFoazhCPNdSijmZWSVby1MFLyMBB3LsRwXJN
1IyXJdnG4pGPl4qsYxmbBWkzlyodOpG2qCtvWsvmdrCG+UjqFi2yq/2grpGyIf4mcZMUK5FxVLgS
KfbaynLDvspONmomJdf5jCmqOH6lstuHyyhAVaEcMDqmMlcUXaHflw+SXazuXXNBRuvbsb4Da1tx
WbCWpoWO7QqiZnBbHMsvNa8NgbjNhtN0l+gw2AxyUWvbIV+tzdkY4Vw1XI9WuJZHApZ36vt235Av
6BH1CjxWj8Gr4R+QDN6AUV6jtlkv0ktItCY+gXU+1CFF8GuncRZpUYwyr7dSrIvGer3R/V46N5d2
INS3vGhtE6/zUzaihdkUjd4rxykS8oFkf+K1BjhqYZyVHTH/46BuKLRvBR8S5f6KnVq7BHjO2o8F
kwQxml8pa9ltLEFl8I8XsIIJtMNWWCxTwN+CdIk5FWmlVp1BuvF10gxgt3R18UMXNzU+LtzdRvtv
CWkmIxnJt8ljFlvUTTbxwiS17+uN8i/OaOP+vc564A9j5mCdwM6c0S+jG0E08GjwlSxpTJMeBoHi
k7fwnDKl4AVeOyW2bIxm9qIx0mU74gj0TFg27Zdn8s1bqTfWtiBeEm9sfF16Xxp5DqjJk68R8sT8
thhExr1hhIMp4l0j2r35+T7kpjrVn+ARPyFr0i5G0agzo4AlQJlG/OmFIV3ZUI0P3b3mt5fxAOZj
fKzFV0cfR5+OKUOvG0dps1+hkjwLvMnlJokL878omdlsADZPw6hroTHp0xdglPlaW4qN9ceUWop6
Q55/PXLXXassfcb8LLeeQzqjBozd8BE2ipNpGNjd5V2WGwiJsBLFN1w4Y7fBl/hxHMlcLGGIQ1u1
CthWjI2mf1qY7V6uw760ja4rAh77rREw+/fc0leFrNOB7Y5KotEE+MG1BO+NST/+tsT1pd4TbFZI
cBS25+00CTyv6Z63+bdalcyUS233eSh7iCOYzcCjSVktw7lG8Vu1wLSw4Wli75GI+qWrjYi0o+qg
0zQm9kvVH4aFIEz9V196Mf/Dow0ijz8FcAZjbgP43LtIDx8AKXA4u/4o9Sgat/pVXRkqt2uSF7yY
5jlE+Ihz/zYk4DE18K8iM5KzJ64jM76qhypYVRKaBx+yycrz38deLHAD5dBDT5pC6zZckAGbHqq7
WRImS338MVlcJHKe1Z7ufcqdZncphY9kMYXR2dYXIWM8leJdnKhIHOUyHsgDrbe8tC7rsREgNMMI
RKnPTUB0zbLAcX2UyrOR/5ueXyO+iEpbFVF9A7TzxSxhkg5/35cv78fkBwglK2oWVs5wrXbRA4aO
uTy5ZqE/+1YucEGKOQcil8WJ6wY3MzPTWYTMSaTtzV64fIV+/4cpAZjDPt6HZUGKhSXE+gVtf6jc
c3YDlVdjmDREdu6XThhv2+K2sgLFgWnNdCNtyfqPXeTqmM3w7FDwWbReo3S7P+vaccQ+z2BpiNhg
vjHypaRd4ZlEWKRmFByTefKKQrC+vU/ILfVqrSH4UwkdFIRWJ4njVUIx4w65QsrNkPyMUOa022gn
61MwhchqCvEC6tSqNGoVr+4ST/BREhrnVHs/wWQBN3+SaqRVtz8/wW49m4e4RWPPSZb0T6bUAHKm
0VAJCZnNkfvymwn9iGVE9hrOSkaqz+3y2v+Cauhn3b2tGNSf3PIYSWlAUQtVYck0GbqRcfvsuGP0
Sto7dkiGcYo5zkeLu767hCE/1O5med4oJLOp0Iy5o6wT1pxs5Qxwzc/cj6neVA06aBFYFhU0VqNh
1KzkzLrSVpt+Su4QTDR0paAeAMDnJ6/zItQOc4rBs/5OXGuyrmGfnLTnuPeYluEvRJ0TXu9jZXo+
ABRvmH+jWuER/5WrQffzqzFNiU22H4WGSLN5QvHSr6vU80VKNe3MbaUY6e2jylt1NZkviSFdXWqc
1hVO9QBmMkxb9QstZtpvBfmx5qmbQfkfvCrx3aF3HhdMQAel/tezhQKxLZr09XIreYlUr7KDjzed
pmiJtiOWDvoGvOK8kfRe+e8jBTlfX1kulaAB2QpmlYRhyrQPmGuLjMVhQlszCAMVKQMAy72Ryfgu
m1JRtdqZgeTZrMqH44/0eXy2/2I4HIVmLoW48gqFDDuB4KxbsOZltonJ/g2mkQs0fpELo5eNhbQa
I8OSvaX3FZ533lP2TKC4ii3LQyWTr6wZZRwaFi6ODrZ1N6v1ByFIHsWOjpCBSBUNi3yyOMYAkP+O
76Gec/e6y+McusCvdsQzsNntFRmbywU0c1zrNVFDX06W0SV+cXCtzjC9t1xlX1o9JwavnUiMKmvV
EAD+flvlWYg1OlNcMJMGGAj7Ipto2PLq2oUxE6ZT76of61CwsVJ5q1o6CDdBZwgRrDsJ7q13V4Zz
6/StE/G+UTh2+2epOQadQeJQJ0sX4ihWtI8v+RNV4RSs+qRuv3Gmyh3iR4EXL7hwMmUrepQbd7tH
uWHhl18KxNN7TmltBKaohuwqQqm/wTzrliQcem95I2JICv+4LmSNW9Xh8VT0uxWYLDYMjBiZdi40
5+3NdoTi9XTwv1RaacrYBqcdNtwiJHMe2SEMIaAatljBtugfDNdL7esC26BqlPc7QXwF+HamnCR/
mYmaYg9WBgN3lNYYAkeDD0CupCtS/qw5V0r01kDiRpU/fAJTHT96HB4a434piivHhLDNG77Uqwfq
YhoeqQ4l1+pRFWWzXhn2skgPOH7CisLQdeR43LEgstINqqgbxpilYs3GQuZ8YDhV8+Xhvq2X4xbo
iU3lsVMJLdjyb89uLersL0lOSGMcFcakhw+7KkfJY9gVZpVQxsNBM1rzRa6ApxWn1mKwq6VFhAVO
A7aKxwVVXXQUbQzqFJiWwKAtxLxo/T2idMufQSHxOsZjDHzh7Yu7M4ABnndZ8A2F0j4cKm3GnvyB
ftMIXyKA38yraZCPO+oXikAEtVfPDFiMutKetdjfwhWiw/28BWb+rdr87OTmCw3OkX8/xMBZiPxD
G3AC05eN88hzl6PYuuE5eYDbVwljgivHkWFkNwAp6UTjc71PjPXjOmAqvI6Sa6w15t8Bamqb4ehO
Ox/6M73j4zxkwVKfKHQEkxamSWavFku2yhRGbgoN0z8uw2nL8PxKzDaM4vOPrcZbxyjG97wwxM84
1gvfYRaZA4u5CQU5CzC8PhryKCZqwdaprHxO9m6MmJ4clAzUE9bZCt6oVZ9NkuPDue07+31N9oFC
i1agdRNYds+Lkch9HfvrEvek8yAlGHroelPzLhtC8yr6XIfOYNv+TnIGx10JSSc3ElRgCAUJBRFv
3AjBBFPlzYDj0W0uH6IpfAT+oRLqcZOb/8vogDaxQSP3g+73y7IlXjZVnKzfXlxQJ1WyVTi6ouzL
bUFLUVxczrQMlpuYz1vG2i0tpY3AXwE3tg7zQEx2DGVM1jCfMdAYad9p4gp48P73/+jb7Jb7Pgxz
NEwEhPTSmLeLxeXE6hlPIpVUOomRB2uoYNSpzhRTvtgAncOopAyPSw2nXJvx0mizd1bwxfmOEMlO
AdXStMF1LirOdSB1bW/HKkvqr4QdvRfgUckXPyn36Rz5W/+sHQFlPcbinGWmi2T4MFVbWagBCxj9
4aB8qt7C/0JrlVnl1kEqP/qc/mE/K8nvL9PpvuGxbhF1xew5PxyG156rK4RgDoTqs5pq1RPb/3V4
b8lY2MlnBkJKfJg5wQtFWvfnxIQK+wcULxfsQDPwIZrjSt9lU3NqWf75nOQIQePIJhIBFStLxFxd
04LevKQc8O20g7oNcCtELRMnwawnRPBFhNu8zZJP2fLQlM8UpdoRL74Ec951dYuic0LtIj1v0aWJ
91OVb032phV5FxY2AU9PqovXgscREIC+J0UDrlQZpKe87xlhxYUnhzewmRTRxDWek9G58yj6toIP
Iw9O3WXbMo1q5ZzIR4U70tcLF/SrXr7P9zceGM0vQjGTorQGrMDIOftm4H5DHNWfTCyq55xHruFd
EYpVsmoxv8AJ7BQv7oAV66/R1aGvAKmk1RD/x0CMEeSdhFePcI0tGpIrRdha/1BX+R2/7WW2jPZX
Kem9ycvrhSDe9GtthhdLY0aH/NRvp0XprX0TGtak3ACt8KxMDmJm8F+xb0xfzQ+5VB4OgQcSsJer
hv7dJm1PxUTXWbmj7G6h/PDJkZPO3D8/KzHxmUkHghVjFgkqSqzZw4sOTBEklTjNDRNs6/RAA9D4
hL/df6sSPwC0pI8sgp6mDkoGJk/qmAAXJH2PP4t/JycRVAKD4DPcD8P1d5ZfHwuOh6GQi49kSfbo
SaXLUlSaiKItWnV/4sI6sqwrhj3zp0QQpCs+KWLcc+k0OGhzGVRMZC0XdwYbqfCCIooiUBadIAKq
N0YhbM15q6z4/L9aIY3xn2iuIAywMy0gnxRJRHAlCMBt2CUw8vxeBulKmxfzC8mTZ/e11UaUlTiB
2UJsTDe/cLVQ1vuHWzkiyjP3VDzEU6IPAKfNKd8VOyA3bvkM8Drn6OTRbrXeVxrxC97qGYn1zg2K
1pouGc6be1tjjIj+hqHUJQgHKBOj2HqabId9lLrF1+aRTItLzRnmRtL68gM0iowTztspLl3g1Gc7
xzXbnMiypOl2FxLg2wurPbwymWZXE7exxX14mo85HNvW4FuSYHvr3Jdqfuj3tU9PJabe7WxMtlFw
d8E6D0laZ7bYLdHADWys+hxVFonAYcQfTv+0R0mgu+A2/px6H0XgMAQINFWBIkO6fVzuUEaojlUk
Y0vwphDMG/11J26TsBIMn+GajsDrEG2FSopDKfAnHKMtH6amGtskUukw3IvKvddgJi68JYGi/88l
erclJVWVac8hXDIvVooNCbc1qozScETm00DwXNmFymN2UH8FwCej8GTwFcDPoJc46Ai12Bep8TLJ
heS1M2ttt5TdBiP7zv0OM2ynje1Clal8G2teKYxt8ohkX1K/cU0aA6uTH0tCrmiVV1SzQ/CaJUFR
aQE/f4OkWI+1zueVVlG6nsQpW7RX9Lskgt4oI7LvMPrXbRZdhyp5xP26ylh2lm8uyGq1OV4SSDlf
OHyXdEfh4799DiWfRyMCMkwZrJ3XOOeRmwGtcEDVKqgsozrMh+C50qhfpP1Mrx4aMLxvuRjEGRTF
Tir7qvO1tllsPWGZUOE5ukTiIDAZbT/xGoZwZvoIHdJWGnVTsbq89wopq/hqL5v9hVLvNPJVBcXA
3UrXaNc7pV8IOaWBGs3bR+cz9lY18OLCCX/1NqNOmUfT9GcaeULYKXw3Y2XmALCU3LzUow6XQ5G4
/3gf5qTclqezVFkLkM6R0lcV82Ii46zZ19pjVQFC9S8EBmg2C2EB/LCMVolw0UDWc9ltbogGCmR8
Thdi7MNIO4pjfxRitRnsJXMLs7U8WQBlgShzrf5T6c18nHvmdIuX28HZfy6xXUm4FrW6ShXzhZcd
vtpdf7la72kgYBydE3s0+YDnC5XlTcNavcX41QstQjFw7ZtnjNhxep7paM1jQh7rfwR65co5P16H
TH99sW8kdhR0osMvNtjBPqZlxltfnZA2ndrWb7cD+JvxmaVnQdPrAVIQ6/Ru7DAafZjvOpqKpbsX
6mhAfZBefv+NkdPX0ZkLLNrURoV3VtmdruNeld91Ft8RBBiVQZ2fmeL5hvmmVGhRqSIkH7sAj0tO
3qJ3LUWl87pd2AFVoEG5woRAHCnaXfipOWdjJO1nnHrR4a+8/kK3wfNah7VN1H//BirXSf0X5CNx
/o/hn82Njudb0VnbzK9dqT/5q7dwYWNIJQp5XaFJe3YBf/xykRM29ZU0BfhGeCllEtWxiw66Gmwt
oMt7eXipo/DvmdMeasnAMX0cyN7iqNUxuKRyoL4HaAXNugtF72zTdm6puR2mDMLHtrAzKizOaTba
22d9BQCD0S2tSa44DxOG5g6IFMd2IkEQPTDxruec9QdCila8BfbRsDxOR+elaLHdHItheqA38M3+
X1c/M9Qf/3TvC5Ib8dcLlTJbZiMmfGhs1P2PUmqGh6XeP201v1iQdl72nhKwfXX46ftt4f9lILjf
NqnViEyQExkKpVEHCrtxXLWZC+ByXhu3UwsX86HnIzVnGw3OKi7g+fvEHU3jLpl+Atmuq9YXPICr
XV/iPiQ5+YVxmmOEEitR1Yk9TG9B/FoyEwyMqI+8xCsP0DOyq5s/9InIWjrYS3nOWMNfgAx4YutH
2ste69rpjPPVho37wcpyoMKeJba4SAVKpd5KKny8r/erDOaf3vo8aik0lGRZ3tH+kOOc+HKV+gI4
JkV0A+krANE+CFehQfcc2oBPzOPwSms62zL0+ER1iC3jK7Mvp7bu6Fl6O1xY/joSYnPGBerj0syY
ABaCZeU1ozUS5LwhyERAS+kneOxHne/1gXbCVOLkWfj8NYN8TWImeTy+ljNldkaVs79DgGQ8s+qh
HrHIwxPG1ePTRwzibUBREWHC7vjKTxt1UE0DoygCrEnvQf5CZZCKPlYhD7kRxAyTqwFyJoanC8Rg
dwnRJpla540+FlmJCkVZ+8J8h468kZ54HQa72msdZoPXgNk6jj3DF/z6/pOI2hVUKhECZEqjdny4
86TL0dzxhRk6KsVLofCc1LkgNvZS+fCrkwGNZ34imnggtRnpZAmULUq3OUVYKu5CA2Pi79Vo4NUz
L5Slrnf9IKG92Dy8I4yApZD9zSGrzS4+K/dWHiRr5NICb6rN2LOYTdpycoRuHMHPVTewwzFNovhQ
HwbM46VN2YI73BTu3Xl4+eK3s6y6Saf1eO4T6OAJUY1/ty+4d0XhaVjRLlaPtVMFRNcKlnC3RRBr
IR2ulU5I/WTZ+OHn7RntyEtu6cG/oV1eaikaqJfTzFbNovjU/HQZpeCm8gOVbsLpJwsEnjm0918V
OtL7Rj6jLi9Nv9iXuOyZ/86ihMNeJykpzmkgiBEA+MBPFVUZC0WRJe9C5Y7mBu8omzO7ZUgwVdYN
hhsjdBqrtuyuN0gR7zX9bMTNLHTRRhQzIimBXKgvZrFtiavzdA8IzwoYatg7UQiG/zFKWixLhrlH
rd/JxwsI8UKu+FHO4BShPIy12oZU4NXNP/4JMAIoz4pdk4I7m8g3+qHQOaLZmwRAXbbFsoa5P+Hg
fu8UTo80xDcF/65j3OQ/w916ZYF2PMjtIPdusHqk7IrfmSqj4kpQhoqf5OxhnbpZwsYFZRTN+UO4
QaJX0XBPViuRnlmmLwFfSiPXBeDzJ8/OpDbmOJ7ZTEisleYQiYj3zzeqJtrl0CSNUmYxAwCbyDnY
VP/308wMOVf0aq6isj60Bj9xXU2Nn8gT6V6Qy/9A8nRmZNGXJSruuWX0Pd/3SThDjBHutwQ4n1uS
ThAXwPZZ3nBAyN4vZC1kHIrqk0hdulW8lWd8qX0HreolNNISw+YbHf147b4qBxQPfQS8BZEXeSwA
p+1NS1uBvo48TvV/H5ddf2fwD2X8e6SXsb/LgF8LjCBqH2ghKtBwQxIHvwNlFbXPpZuXtHyX8ms+
Myd6S666VL1tHNIG/8ICXimX6hKUSDedJZ3Dq9MrTSphZvs7QHS4+e7IY9Ua1+I9XlTaYI75t1M4
3krJGBJs9WdzplzJXNdCpJ75GgQaUfhOj2NdPbYfiVU0yEr+Lx+5eRrvGq0oAPuyrChCvhEUE2Zu
KV+rVnco99zdG4FWT+bykIHb7g4w12i0SkqcDBLyD2wa8fNcwBLuWACIdB2sAAtoYk3TVjk74y8j
IBVUyjqnuy+Djj0/J83QGKwiETTZyyeZSFG7/NFuLB0rMcMKLBzmc5uka1t+7BzNqe9pr50/UL/3
ZTZgjtKf8j2TBKzBxC5FnK13V7ECB6uyBinkZCu4aRD+3YLzZGL++9E2FwgfTxnk34xFbbQvgIZ0
EpUR2MmTbJiRabVkSg8WBYLG/i91weCWlVm4Qfsv18VX2tQzDce3OsrjYY8qpdJze61dxYE0uYkg
ODo1Yp0MrAYEhnk6DzdgTbZnFjP41nqY6GnHs/MifRsijRQi9erJPigEonM8FnxbsioHCQ0TRT0V
yM3S3lIva9QdRsSuAN2MmyuSTUg9Es4Nscqmg1gVAJyCmJP0UPxQL1SiwGOH3VAEEYLDl8/ZHj7i
moRRmoiJC68wRI70dSvZLvKBpCupMC1pLsBQ4DWjMeKv91jSTw0NMuTIwRw8P0yM9tVYfpHr6bS5
uc2bBmh30/vzZ27fv7G3qfkv99xkY0BJiD94Av78B2oihI7UkJ8NHSSBl7wkmQBqG84SQdbmg5Xa
IfFm20/NPPNoDoUEewkjwEHMtnINdNCNWwW58Ym2pHzgEqc8TmvBX2zQTX1h2TnDu+y06q/fkQ6R
N3Y8BQVy+5YkqJTHYO+RO1Aoh+O0NZ/8vacwjRjmHol0v6Wu9gvQCm603hBODO5rGhkpqoeuVgKH
I+83OZkZ11PrTA15Z2BWuGGowLT9vK69BdXjzvAY1MjUBlz6KVTEZhy4Z5kjaHs6I3TTEKVvAPhX
LfljK0m5avQvMiRaxAO5i3hjEARkOHPWOXs/hI6hIjk1a4KmgCUk7tWAxE0OWSEEhrKUIhoK81sV
XJr+5lMzrEoOdPJgFvlKdv4uPR7LhXD520LN5DKoz+v1eW8I+3umdmujkFvYosr6dFx9hm8wNyXr
Pv7HOm1c404h7ibPz92Hw04itRWaCXyZlx1hm+iQmkHtO7+qkSm4RHZZ0B6aso3xNUnnzEB71T3j
ekQRFGN26h1jbzOlWgfGMMVtvkEo30pLe9GFM8syEKSxD8otKdq7681hGrhG2yr7mGhwvdHpKi/V
rCYdkg3PXnxgQZ6ttnWcDkO+rWSoohsuQg0uW9PuW4xOtJq6symuPmvYZ01O+99JwfM+u+sO2X+O
LXGkKL66q3H8NlRy5hs58K2i45DLHbz78G4+naOk50r7+gCRM2zr6L41c9c1CaNDfbL0kZPG73o7
i3XppNobr/Vqiu9gtayg6NxCgOgAcn5QM/cNMes17OCuBpjt4asK2trNy8eYyU6iN9+RlE5xe7GW
Tct6j6PYCT5S7hMAHYCL1GxmCRd9BPQYMGeb3FGoKStrJjV5UCiMR+ojIrFqkK0YgVSNZ+wm2qX2
YWXXuGvrpfCGRjPLTXVv0J3FCCDyh3qeRrB+OSRfMMZooLwcdhqF8tIlVd6gYkNYSEjSB3WV3x4h
5cGHdBp5ULz7dPHLcmY++aDBwvINBOlJbwu+0kWknrNUP5L6umm0v34GWVS47s9QMA2ObVWgdUB6
DNKbgEPCS+Ej1Vd1ygUx6iXoLz19woYG9puL5dvtFaLrSHKQRRiNp7TMCM9Jjtm+xB4fOQFCQcZj
E3Ubt/CQb01QKnxfclcv1IMynn9RscbIVPPg1S9D3rbIi/05KpRNkh3cYWBSsqd4KjC8VXprsRjD
cGwOYrcFqLEqu8Sz5IuDqKwB2CZmg62xKMFn9pGrurUkXHYPiDVeDg/gH2b075fBIjNgKl8MV6Xj
pM7FQ8mWZQ7EGsIaOWiVFgFKvquu9TWhDksI168vd7mdUhWZBXlIctL2nFGirt1nLQbCioK7LyN5
eMzZx8OKCF/Vp12WBBFbV4etjARtZ6hRqeF8e9dVPTKQgHV/0pcTxPY+kpZJZcwrCxscrKeXcza5
+WJRpfsgh2XudKIW1G6smQqTE4UbPhbhH3eOewF32ei2Syn9aZAzfXR7w3d5/Dv/XqprPmiKXEv6
lj3mo9EfQupSUrtpl/qOEX9il8iSVCrTZhmgbwcguL/hKgzed0fy1tG2WK+CbXmD/tvAvCCrFlsq
ZF8IEIDM78lzRMZ4ICIblCuI8x9KilXVxYOkZ8jwe1svFg56HEd66ADtieRscjgmsj6bra1DfTzc
6xtsuNWuHi6snrD+JU8vvIs+/LdwlYm3Rkf+KxcRvp54d2BSQWalT+aPwSdf+33Lo1cXJK9FC8bL
65CUsEFU2Y0aWTK1yKzlR94DKRtPQ1WE/UyqhhnVw4VChFa/TQt+0foFL9GGnf/25YtQuhSbKe6n
3SYG0CcAXobfrm8vVasjNm8EQ1Aj7qDw7tPc9QBSVPyGi2o8wBzzcngDr6sNqqIxOdaY5avFs3zT
fLLwx4cc4ANmDZdo2OoW5tdTlVkoGIU/wUSPVnJmYRAkJAVazBe08Ejc56IKxi1AqYrBA6rjch1m
2t0E/kwAr0h4+HwWBqRhQZoq3/227u9UMvnhtv6MZDoM0QOS53eswnZ9wvo+RgQlck3aD7aqL1+Y
EE0bZc1Wnhn/1QnXzJZjquDrjpbT0huMGusaKVP/KDLw1JF3Kj7XUzNMB2TCF0YnAS0fimOCFT9h
iDho97M1J/5r/MmhhIyLrLKCPezFJqTc0Pgy53kZ7TUgbZuAadbbaHr3IyEflZunYOGaw5IYHn90
ptjN6xqyWnzXDOXAcg1nSya5iuLTnG6crcrOmjKBnwmzfJJ/CA/9/43bTPkcpzrF6ow8RZSfkvUw
bjjER6ADdihevA6nGk+3OmyH0wHYmiKZlAbocEz92dtVPiLhCHJWHnDdcT64zFyQ7zhiouA3SUWg
k4+rp8VDCmwnu0xSeidtAgHAZIXHhMOUsWXvqkJdVHyE1fSyqVey6Qq4VAdBeW3x4HoXnJVY/j/e
ruOIY9YQU7IAJcGI/YJbB9q6krEAUrJfBpOVF1N1K5BKZb8980/7uMczBfmQqGhEybPoCrl4404U
X0S5qdMC1O1nEx3IkRzg5+SMS8Hanz+jtVn4UwauZFYj27qFiKlEnkb1MKKxlhehSHrU01h55b5K
nSmNmau5FvrdEF7DTi212LfFFUrpGE2xOcrH3ze3ft3Iiqhw8FWNBT+2TakTJGOy9VICM8Wiux/L
1p6D5I2eu0wwqixBWbtFuDkJ3gfwe78eZ/ptVj/4ArAk04jOQQiTCXjq0ZXyDASpqH5CYHoYwwuL
rABNSXBF0CfiMX2ky2VJfOqXLrVCFtiIXXlR5JthKPUaiieyN+O9fVkEg81afcvV7xcmmPMhZwW8
Zgll+qhFjKlCdiTQoIqfrJxpWRvs6a9aY+R0DK4lmZxaWI45O0v9impRFZNRdOKpTCBIhf2RZxkD
cMnrd9dBxjOJSFVxPa3iAmvr1wlfquuIvxC0zYQueWpgq6RRRD5PmUnoN3GmU+UrLg8NkYxmnlDO
TQ1zOo0ykcqTIv6cqV872E+OPPcbceMmc++h794oi8+2vgMEzN/IxG7RNhsKJDYvyljW3T9ridDn
ms5WuCL/WtsWfpwt0eu7zZrejuFBVXatAzlJddUmxSjecMBCnr5oguxcpB8NJvB6ftrBc034GH9V
FOSGrbj0NclaqeR8C3T5lRYjberWrPz7LAesRMDesFwRqBagSa4yoawviOaOTeqjjG00p1V0zd69
RWUm+J555MqYC7/iMRfmWHqn1P2gP/1M3Vu/7vINUzwPddUtteYvYBPnHObpz0di+ZTQf5qAZaqr
LzN7A0aPpcMce8Nf1/Cvt6J3aq76j/E9O7c413sIcyDg9om0uZdfrutjOZuTzOwmnAg7jY/WsB0e
I/DoFxEMGp1sBXuNWdieCH4NfkFkcw/AmbuxESbenu2DQEqxpzwkVbCm7sqYMkVk8BcTf+YBbDL2
1QA2x4PR3Fmnajk2rrGaMbeLk4ZjpSDWboPBJbZqR5YJmqUfKF59HD6skIua6iDUwGDpNDyzBAWJ
i26DOfZN3rfxwMUQj11c2/SqQj+Q+xM5Wa6OLNj6k6Db2LuuH6aP1OxSdA1oVy8i8qTVgMOcEEGJ
AEa0u2teF7j2q4fR2ndwxyXm33oYsZy+9whrMyvuTWo3EQrTluorE/VgSYJfSKEj/1KnOolubFJM
PXvsHqhhLKsF0bbCxf6dI1L/cjFE+eoHuRjZSohR/BdAD5+TJirZNuvQkl8RQJ0vP4meC2iZ68ag
wCamZXvhiXHYb+Gt1Xq6cnFzE+ChazAdpgiY08gKi39y867CGSf30tynSPMpjxLgKjv56HI2hEBU
aFRZ0hae/LjaJWLY+5DktAY56pHzDA84S3qM5A3tGhOJdkGEvUzdtmDwMpAP9wSr/1REgqr7jRPp
o9/vCJ7dVsgsaAxLxXMHOhxX4aJgmIffi7L883Lj4xkzuzDCSJ37XppsJUNZKhOO/HBSo+DrLCZB
EmqxaDh5ZuNXxCjLIoAupCNMhdL1FuFBQ7HVdYtiwNiThYNMW2t0F2G1YWB7hryCTeww2hD1LkBR
n0QsXgd/6FdQRHUWnx/w496635OuQmVaaL1bai5/qb6O0FwvMcMVIqrqAoxXS1juTHs1zY0dWJG2
j6/6PReX5eF2GuKuXBW6wNPndf1+j7iKr9pOfQe5kp743weC1XY1+Hqkf8A6yTUUPF45zdYklSgR
tZRlu6esGkbeIz064iMeyvh5Jr+w1kV2JYJRbOBGyzsPU14+m2q960ih6sJx665bNavfFYy1boBC
K/jF2YaNfJEqSW3RUC7JAeIOcbF2N1qCUi52w08UT2R+UdPm12AV3BUMRP9+FS/UsprxVBY+aXTq
J/e/C74BIsQqhh9pTyB6+T6EQMO0y979k/A78fjYmnK8j9q3g6fukMHJgchJazWZmOlUjHUQqEoa
LZccDoc/yRXHn7aat3nRFeJYxB/zklbmCr1w9r48UHZWJLCNpF/6nNvUNLsHbkTENxuMViRRdsho
tNtaokd8FOdjRc3uhGllITVq3G5eRxtuA9gH5ZOVEwvKrxkshvAfZz6u2rXgii/6IKAbHXKmSQVX
BL9ynYwhN2KDoxmPGQcF14IJFgEKaly1aI0Jlx7WYXeyfpR4HIHNHn9rItlOkIk5QnOxTF/kQLC7
ddqnxdMGz2PJsV1Oy2UlTBSu1MRDUVw1rmpw9ZWfOt4/bxsSlLas5JKM7wMf+KJDlzsINPS0hqDf
7ZurdbuZvgeC7PdeegTJ/DBCs3QOxPvzBYYYXLJqkgEGXo0IX+0rqMKRHSq8+xtDL67ApMMVYiz2
xfUbF2LSF0l4EgcOn9mDzs90ejBHSM0wFk2wOHZZ3M/VGNcF1iwUAZy3FFbYFNJkPGE3z0MT50l6
K79H1Q91RyLVrbiZgCi5B0zmd6jlpI5XfwGoYGDetv1EYhKjlQV+vBVqrTUPOv6XXlf5Ak/RQL3l
gbdQPR5OCxhOG3mCkt/ucQUb/Zt4gCy8ymqLQZVFe4Y4PM2L2w5jBURMHYR7qNk36FH9o0KrSKmG
itOl6fdS3ZJxMDidE9/R+HUiidUp/Rzlff9HI5AohMQvhoyYpY52GsuzBZwhKX1QvXhRoDmK3710
8/2F+ke9SihDnRVWgqgAzf0VOuCngT7Bn14xZl21MAHCqiXeMK7V3h/+gWIzwyveJOG8LHj5ePhz
kuazJmbigd65BqffZ77CJDbRBnQYJ/yI0A3tkCVO4Xc+TAL4cldtFbgFeJxgQX2BkLckHj+Fx6um
kCWTNqLFz3LtZVNaPkVeeNCG6dRLGxD44fmDPVaaXezip7HXz0DLzrZNvGASq3hUgtLqOgPoMu/J
qyjrfWxDmJQxd6fCjEg2KPjTe9Fu4+e9TsReN93sRR5Lh1heJump71uRdAfP9pr2xv2vvGZ2uknH
3IbXPZUquXXJeAbCZpbniJSK51HmK4rZ4szJsJEvlmOpRvcrJSm8rvuY5DzYn+apdXcL6a8toW2Z
XZ3kHp0HW3eX56ovFOv9r/ygna8F7zhK/DyXcfvSjZNsZSfpBludPrZ8+XuinMu9VWYJOB7v9+9P
NLjnW8UlyA9quCgRnYPFrLwjXr8q6l1e+KbS3/n7TSF/eVQiMkM6bFtWz45gaf+RYST6B5r6B1xm
nX84GX0rNYdFxSH7yOLgMhuK9JvvCUjg9jYdN4pYiGh1lq2aZpWscxR7isQPIpserMLHFGrcmWhB
oGcFqxBsKa0yIvP53QGsN0AVqiiQ95COgijj3HfVGzGnRwiSh8yAXdCjDkw0Oa9vqB9+0NulXqrk
kE7iIrmfbS1ekm/UHG+BRRHomtmMJywFYIMOnrvOxn/orNk+XHjex+KaV04vjKuFIA0aFu6/CPI3
hxpFVqEhAwEhWFtDzv9SJCDT+t5hw0dB90eCwptJ0EruzNzsYblzEW/R/j99Ubj3D69h7cxsHXxG
i3GH+gkiSM9eTtDtyFDozOJOvYGBmxzBC7AioJ2s4hcZYXVDMTYZtInNuUOebk/GU1uHELtVCdj8
V66gGP3ctYiumKY3l3b3Ql+ajw26haD4BQ9lTDe7w+4vKrQZH/PmsQJ0bRHSwusMBuro/39eyrkP
a52VhO22lNsMAY+4uE0GhzeKh0C+BdW7D8J9B88QgrcOzYVevOX3gYiWIz076bv6sXCi3hwqMC4X
8CGFDEmhi/cQPNTsLkH1ljhtykH4KgoyuqREK8dLacg60eLQk0b/M0mtTWl9QGDzcq6IafQHmyGy
Yr2IZ1AnwIzCz6xAm3Fh2BjQVK953lApyrnjUnBXrs2EoLuobt+XDglPwAzVFFDjCmg01+GLJ504
HnNAyRwMLCj6OcmlPTSio4dyyjBw2n1EG7Tqp9/X5rAbZRQio6ycUPj3obcxe2zChJ9WSGQRVKNC
u4O1wbbu2Z1sumF/S422FV4ZUXupeRG6Gm2AomsW1sCiGQ+e7X5BkYMSlM/8Xq1RUtNwPOhJHZxY
6FwTUNKgQAYSQIVGeNBLvpPLKU19fBKR1AUEPgq1FHYQXA6t/u/aarxOhk8SiFRK87eMEO6zJ7IO
Tng0rSs3TWm/Ao4xzp9F8Eat/5JZPhaUbl0N9k1174/cpi6E4PiznqYtbMjdJEb/OO3mPbAsA4KL
fEuQQjG3qFmC6x/ncBZ1DTB19K7/o5v7h/XCysysjqGP+QIiCFv2ka0zBrFetREQciZxOQSceaLW
9U5HDjrCgZNb8xizsTqxJRG7p+ofvhkLRh/2ztE5wkqboyX9bww/PD/+2CKkAZSF0Ze3tpDu4Kot
0FmGsXemmlW1YNQkCxXXAjSUHyIsUxlWGIyfrQapuTFWtXhqS/Ujs32VeA7YuzyPqL17yvfuNH4d
j8mK/0GquGzz5m1hklRNsQVd1j9mcqAi1GL5EwBAmr3yDlQTgEBaixJU+JLOJUkqSPCv8iyvXXj1
9t9fpl3nc2me5x3DYuMCTJWPxlgzQxmc4jEiS/EqBaRivZi57gpbbLGEincTzvsrLIFPZDXP8sBw
dt36j7FWKVjSe3jJjoqdGzGoH87fmD9YWhL6Gg8Je9n8wT98PWmjgTVzs0xY5/o8JC5lc1QuZ+XV
znJcY6NX8rHk8wAgvy1Ga7uLzqPXovpVYCKqI2EysJbmyXj7ninOVfF+LdxCdefV0Z8Yk2y64/5e
cSgNTgQIJxE34dAv6c+/jno7qsMG7frgmFc3MZPVpGK3pdWw/HM6tjzWlfqq1E9lbHazE9uff8xt
Pio18JQ9i0eYynQY1qisvqz3HhzSw356e382UR3j8czSP6ho8RmE9i3QVvb2Rt5n8yiBbLwnIHF+
fhB/3q/tBS0Z6zSSOVVA9a3mYiw0BpaKDwjdqGkK9nlYDPDBD9PCszxG4+Q45Whmht+ulrMcnsk3
tA0gma8scPmLPhREPJoIe0YuRGhC12AYaqL5M/0BtcZx+Vs6hSlYF6NpoY5qD2Vegp7lMX5ZySJx
yCyux+/IBmIAzrxWlZ4Pi+Vf8Emc+nlNFeMhs6zlufYLx1xj6YPWvJjMdJ2o90RsIkinRAOTS/Xi
mQWp2eKBBBKfR3x0vPx12uiWBy3WlzZjkkz8ws1k3Eug+YecpCNh0U34WYAxKMBj5AjHRE38cDR2
RbZSds8AIo2Z037gH/21RRhkvL+ixWhvJVO3mhIsK6BaftQQ5SUZO029kH3rE/U9+B819iQ3+7x8
SBRf6KpfvDPZciKNULK7FxvYLP3DOpEc1nGvRWdo/pnDMXTJwYRRL4mCC1rIBp2aDbxZCuTRn1kG
4cWHnGHRRUh99aiGyF8T3RdVIYFTYz7ZBIPUMYi1rI/hxkrKxdAO+SWLQcntuo0H7xyHMI5zjSzI
XajdzG/MLj8M7jPxhtkYcU7hqmErpt9UShvaQGrlytCwaPuORvui3dmiX8pfnIuWu1nF7MDe46i4
ROQ+yAqBsQ4rTDOCy+BSPmkbIJtgDA6b8bjJ1YL5XhxE9JpegaGuUsnOP7hHgx0On1QgpyygDBcY
s0xbGPUfnUFY0hCx0oswoEQM/SmjRNyCAkfJwuHeYeMoJKouZbaTGpUp70PYnHCn25aoN1mFaRUH
SRxw40Xoq8IuGGVzccxjbybNAQRuFeedQ8FpVVe0ZppBcSIw/9GhHdR3OtbBsz0znus662cZFF6m
1KiifwSmmS/a5u95+0IeOx7bMvp6RKbSupqOk4K9smV2ICFjWFcu8yAH+zg78SP0M9dSBs3VMjbw
PhRYrABptewVxHSsUaI+ASNvUN+4MVHzd9jVJ5LM7CF1sMmzxVwbrxLv26tkiSjUVCklTYnfxFmU
aDk0x//+ItSVTh1fGKrlOKg4koWvDoNexA7rM2HeUJzZiBHb9QE+71k+HpUz6MYe0nitMf0XmFiJ
1d3Bq4shgLdgxNQNLlUMrQUVEnjytMApFFRq5kIwN3mw61y3u0F7hu0lIwPFprDH0L4pOfNZn+v8
QPgxECXGjNlqzjfcV7E72jE0ME8hjUzYrrshI58nXgHbGKRySv6hV/5u9q6+931iaHzkddvnsc7A
vYD4emP1sEftEvY9epxbpXUbJheniG4RfNR0FMCllcwyM2rAf2NldAn5YN6E7LXuVBGBse9q/ssQ
F+CePI9xLFiEt6EUxB8FxPw4iYGO/1YOP3da4MT5mUSeVGjoNBPwL+KX8/Vk06/xbj9GmvGzrKIJ
FXjHNzUeQY5RvVVfkDrDXPQB6iEDdMDZQ689KdjoHnS8j+tIJX8zQnbNet9twmTlQj9XiG8J8DBn
IG9Z+VGiRCZFFoiv9f05aUueR1Q8aSCwUw2Lnzj8cL3YbW8GoLkX8vQtbqHtYJzO6THKykvrzDsN
2xEK8QtIBSrH3RtdG+vCW8Z7Hg5ifdLizghdmI1P4/nJaBDt5HirGIvcouETV2vLSKkBI1ejAiH5
aMJL0ushS5xsWwPqpa7n5ORVxdd2sRPWU4ubSC1IDhH0Wh4l9UedxQTo99GHQC0rIJFnWluNRYZp
cHoJ7H8kT4H4n+ldMeGq+7JzRGSi2qbMs8PvMXVwH2sRqX0w/1ePBxMZPUr/1vBSs9KRk90RUB/m
lrGbgh0CxMN4t7/SGEKq/ML40xbaKNaCPdrSXD+xoO45JoZw3liE7x+KSxOmdGxoFXNhYOMBYs/w
zCmH3Mi1zZ18SsKZLN5k02GFy5OYToaJJ/K7bR29nY/yzg3KS+fBPttiUvp4kbPKwqmSR0UdXu9J
Qj5x3ws8Sp5x2VhLf9kTfZGUK5xM+TYMEti/ChHK5hIEEBuE5UycDMaQmt3lyaMSEXExV8tVFgNi
IfXk53aSMFYGNz8uYEG2CPqSBGeULoFvqlrtgBqD9fGz1qqJwNm2gFLrfV0+jajAkUhDHyffQgMk
2z5T9pV7oIDtkIn4uCc6hQBuIbcKffbBvE09ZyLtlEnIsg8upeGZhp7hY+ZdLiEByt2Wlp8tSaTW
NRLdjpXmuFG6iupsaR7x1ccIt0irNVqnT3sfLOffqBuE/nlqfwshGUXQMhaRYO83ezVQZEp34wT0
b1XUORBxLgNpdCKquc6je8tDXIDMoGv0nc3zJPxqPt2TI4tctUXjujNzPngeupLQKbluksTtu1r4
/cjVmgWNvu83CwStzTJvVjWxZFPiUH2It498JFiTdZ958eApccCv3U3orIuwZC7o6/MqQEOORW5d
bFzr2G/e30vV9fNFfr+JDcuzZDB559sDgYzuvK1J0OsI73iJSfqeFwW7rOsNjpmjRF+Yjb5GkhhK
n7fLGmqQ1kdjfMr74FE1u7Nph1VV+MiIP4u4DVUAdHU4VymovLZsM+SfS9GP4UXQ2ju9GnUQ4tuP
LW2zxjUwgSUsX9dPheMGn/rE2Qs1OxUqlGZzE8CLOIzi04mlnvagtkHwvF7RWmCeouYdIbLX4Vy+
HrHp1yrhQKECHNKTybd/u6PUDIm7jCgApdaXxJrp3wEQt0XVvdcu60diEmaidzaEFlv1jgIA2Crr
c8NSyqBWfL+y56G4cHsVFQ0YgYEIClxP6t3WojfMmrxSrvYxTlqI13T1FzvBRUmofWzxfT7yJn/N
ZWQb5hrq69zVf93TW1pZNrmzWxxsLy7XSapGi64baMCcsSVizCeaIqeywG4Vs12rcGRIXDUHzMVM
5jk+sXMja5QyP5XcqzBCwIxCaauF/MMAUu8E/xxOx8N3rIuLWqkbknLjOE1bhX5dDupUplmtB65c
I/Q/fjUDA8If6XvJTSjTcC41Ijj7zMrIulRm3ezbgEydzYm6gzD1CX+0ChFrhe7Z+qv6dy5HNO6i
xxtrik4cZOH6c0+8R+wTv7eHj8gKvZRSVCPM55A35qANqPGMAzwA7ma69JaEouP4oJpyVD1FTD9Q
/wIQe583jRBZN76TUoaNjv3A4ot9sH58pxB4IqlrrjrrcyJd70eCq40pXEgDmZAIp0y87Gybx99W
cujl6hw0WQBcBXuLyR7T8LsmILmzPbvQsXGjYEEjRvajLBlZUwxVnbizOjoMiqobRVBoyEJgMBTy
sdXlaORZcI7ktyF5sBpeQ8aS95zo/JbuyKY6bj/QXNOBS0f7XIRJBvMYwnmCyPsQb/NvjZFmPDTR
BKxkfoX+Lg3k95pI3KEaHHN4kIcr+nst0lFJHUMVR8ld7L8T+0IOYj6fzrU91rQODBDPQvxabcsV
8HX2mF9GedZeQtkNmUOcmnB85BtYb90xqgQOvy82De6glasfama/kMmEorzVHTxzXCzAnoFWGkey
zRWf0Ma6xP8AxFQ3XHeTXho9DCW3tYpcWXJYdil8wlLKZ+VTMTTHYZJniC33hWQ/AGNbPCPI/EsK
5J2+gpWYTRweA2E70YO3BNDPez/dhroYX6k8feF2qWwvzln+1c1BRUJ8T0C++AzVDOjjJqHUoUpA
iFXjj4VRKGrDwVd8F+wKL3HWlfXotU5thnRC1mU4aAFmHX6ODHOPBvpntc1m9S8x88PdS55l3yJM
kLmLe0UxRfrUcNkiLSyW6a1KyJVtHbCrl+anzyL40IlUsOH803tWgKKd6UZQmKA9IBYuw4SBzfpW
pTlH+OUdeG+p321b8mTlx6VoHMhuAgyBS1ZXetwnctEjgizB15OUbMYRI8qpz8I4qtvfXfTFXEWj
81Ur+ZaaCu8R8wLXT31yhIlR+cLmmCB0QHp98WRpaVlw8g1dsoSLYZ7/Ld9w+l0fGc8eM2B9hLbR
hYSuk0tcLD0MiJxEO9Xem1k9t3a1ma9sSm7dXoPd5wT4RyNhDZ+0JuQk9Gb7duXdtS/5a1zNYeiw
RF6PRlEmPrQY2bGoC3ryUYlhtiDcXbCs3XTki+ZhyITYz3xjhEjXaM2v2rSpLrBWtSUJ6dlZUBDd
5XT4SnTq/YAtRSn9Zm9nlJgNzRJwO/l87Ysi/S1K+LHyh8Tbg5FoMlvfrnhiSf0V8AMPuBXCum2f
hRBs3SYVbs2Zj/85DNtJfE0a1/TxRL3qehYaWg5FwZBPNiVvx9aEuEVJUuZfM4M8+SZYhaCX+eh4
6hVE97AYtJjdwfCXnuaz5ARKAnmTMbAt/Jbha3l8daI/t++gtmwqEWwD3otikqsm29FDWELyjajZ
XB4kfwZsZH6bTxbavJozQuy6LpHUu2am5ge2ZFMAEr56yftvVaDrd+NEUreVm8QdpsPAEdbV1MLh
1aWu0kL9bm0M8GlbODyPMUrbftUXxr3MbT3E6lxY7Ywo/d8UNJpRccJtUEoQpqmZJ0zYjWAdLKM6
2YFAslxyZ/OnrWd75DTkiFHOe5O7WUeg5LbrUBHENdsPupb3K66k/aKv8gSBGiimfjsu3ify1VRM
K9ABqNyovm1jMMuApOGOBGGciFyBlCnpdmQBP4GHohz0n0q0pJiIVDdswiUZf10Ht5zK/OELiMsV
29bIcQVJZTFhinnaeNgCMlNHcW3QWn7WJF3h9DyI/SPWV80BCq4tnKl6Gb2yookz15wOZ/0oVo9B
UDprqQ0mG8b0FRjhZj+XT8VcdoJfCVB0Lyd6sylnF720vBKk2dymBBWfeHqg8jk7XOiF54jk79JG
QF0iM1MkfALlAVn/OnZTdP0vuSdZRebHPuCiat8X28LfjlPmfLAeRDu3+8ZeZ/jvbO0VouEaVzVo
YXuaj3AnkX5fK4pz3kIi1/BjPGDQiJnMrW0EHyEwe8683WbDnWY0vl2cpY5q9WyqTrfkZxvQ506Q
J4pSSLRVK9RB7FyMMnzhcA7P0blC3/zCYW09jl/6t+9DY4ArRRAaEu89leLG7Apfi4bAL27AzGnj
Nsmfg+xCPzuFqVpVNCExID+OpkfuV2XbCQC6pNZA6ndM5Y2NI5xk/uidruK92N+e+G3m8WmU70/G
/05+3rdMsc9+l/sLkes1EL7X3J6QCeEBNmxzmfr3zQWiBO2iXi5HLFeQaptKi2WTGNJADULtYFNX
ciAZdEAoKpzxt8/N6jaLpe8XPB6C/9LJb7H5Xc1hetK5hAKVWLqHd/Yw/msOFxWpIv7ImtIdjSCG
L27d9ZyPP7UBwE994ourh2y3FWqd6TF9Bc6qnzUtOccroZzE2WX+fv5gach0Yv9WtnlB9yvUQG6f
nK7lU5axUrD3G4uXR4xTbEBBIQ9Wtz0C+10nOAUajG11Wf/Z5M3OkSsRYusCTON6QnaKGYYspBJT
pDeRH/bYM8afQs2/RuHX0kGT/rsJ+9Eph1JYmEHK2yTKWUo6pYo1xVGtt8h8584C1nZdF5Glh501
Ifb5vG8z1msfpAkgyhGRI7Lfi9csU2UfAa/Qjyz7xSGBrqDVqMHxPSWxnaFPEN+6FQZuw23CdP+9
97mjzqFFdRfCvIAATKtdNzO3URqOCMJdCGp9Nby6+n991cGU8toTjzfncJHHiRshJDxM4XsbkaOL
Dfw3VG83s+V+iiZKUSG10mB3KnS7P3pyn2aJG4AXzpgtgXhv+McH6Hd1uam33NWfCHAaTUQqFwfG
A4idiUnfgf2y2WbEZGDWkcZCp2WX8ed6fp9JruBBTx7/Bl4SQb2V3i4tuRKY9hlvhCR2Bl3sMHhQ
M1xiKm1xVcRO4XjTsL+KprcwmaOSpyhSljnh29s/kVqkL51X1rOmnskn7MPcl3KCwVG0TV+r9S6k
VF5ppmjUhusx3W9s3rb3OcscZCWDaYZFfT1mSTHJYPjobWTUQr5OANNDIH4qTToYzr55J8xAg2tP
N5jM+asl48BuJ2+B9Xxx9WQx8OklDLQYTX+bkYV/BJT5j68oEjdjkT0V7/DRhqtqmsramSVy6CGq
ziW/N2zHCSSuuuhfKVs6+Av+Jp2CD2ayGC9WQ/YzWLimDlqxgO0er+N2sFQX5SntJYMPMGGJsxMW
QgKmQnYHuICSpyicMU7IjImmSPSS8QMcn4anmWB/8Z69vBdepd2hJezXRHFy46xYTQ07bd1LaQiM
1Xx7X2gqcE5k7xrJ9hNmn4FNPTNUfCm5NiqBdpp2ZsuEodPia+hmzGYkrXYx0ygVnoTbwTUaogHd
pbUI3BSjsMA8BTjSnhi8Log/gavHml4eKAAWN0dFwX3FqmPR2fOMklXgDAE9bOnfwSb/ZoPQrXaN
qUdDqaBdAnEBDrkvR7LsVJ5/7LjyGGjEcOV02ANfNm3UsVyUnEvVPJ8HIz3QctnhgEp1ZB+0t1mu
5+a0gEJMBI2plaExruh100U2Ked57BxsTQvC1YRHItlbbL3xK+qVay6HKy5ZaoFlrM7Wc/ZG9+zk
0c7kbfOr5CgEcy0HRNYuHVu+AzQWy9s/V9Lea2OF3Vqm1lXFcKlo1Vs7tv6lEB7X+xk6vRnUHauR
uRNvQ/2ZSg26uWv03K05hsPtJ08mpAWCNpoyJJFsYV0fTgo0Fc1eDuSW43jimuA7JBcZ/2rkTzJP
3BOy6fTRsJ21YzhN5w7qKZPq7fmzYaWLecetVQb7M+sdngQkyCVSfB7NnQPKG5vKDjLK8lHHv7Fs
GSgEDT/hombIyNlb8O94LNY6nlAVaEK8efJv4DXPJ623rZm4jpaUOAAAet6rmF3yZGd2uLYDNlBl
LukGtckIuhuXP2W0UJKvEYzopI5qxv3lT0O5X8ox9xRR/WSe8w4zYtCj1LpXLkFYOcqNPM4niAh1
fKSkPYG410/3DaCHXgvse/i6Du1w2aRo96XvuZGiSMMAP2aQn2dDhKMAiSdPtqdx5UcjHuYJJC4J
NNS3Y467RI4fDCYXOQNJsOEHRlUs8loDwLzgK83XFvAda1jXlwgT/ZewoqxZ4Oc8nqeFQRDzPPBH
QeCOWgGNsWHrICdWSPFmFNggjdsDPrsx32j/uXqF645r26sy6kdH/mdU7zi3ltpmQX6swGFl9z9M
LccFgCd2BMAwje0yVJMELIu3PuvQjKWH+zh0p4VluEMEij0Lw1d+uB4f999ns7v3U82bgBLlz8Bl
jzdnhzEPSJQAUrdu4vROsaug0U7xPNbDG6+SSXvKMUVSQ8A+sm+DDatqxHbqWwDYC7Bd2L782Bha
eymn4CFYionzJibju6DmZP8rXwSozM+KPyIpTbk2X+iCbhvTnU2wvbMB44d7Qt3mlbHYsfHZQGxH
lzWHqOKxtgtUra3bu0RAUHQbEYtcVJa+4b3sCLBQ7BJ3g/zxx+mfcsrs3gt8wuqsbshmUpkXZjXp
yx+VHwGKVJWPiCMXCfVkzZl2s6AuB0XKCbTgYc49SeFAA/LbmgGaML9kkl355abaq960GRqSgSmM
SUw2c8OLtecXDRtIJc8QS9Ij3eGZ5eSMgUyiRr2GHJIH+gyKJpARV1BKXTeZtNLiNUCs7yzKGJot
9PCLCcg5Ya6V51BbGj6fH8qSGvRYWEjElmCqkJ3e0fBr4LOLcnC230BHBl0WsjE3QlRu5QKoQCey
lmni+7MmxbMULd9/lFSlDWH6CnQWSC9HdXPP/n/uGX8ZrsY/6LkiHCwlIW++BmIK7cIXGQ77vCKN
FzF99qRW3+AhRfHYxcfJ91QYjfI52/ZvFU8+83zFX2ruJtyCFKUwphoZkX234uPHBbfv8WXOgYvU
AjUVpURY4R6oeHO8nKgkwu0Sy2mIjev34p8aasp6Bmrud9/fQULEbsdZ+N8uw7mQRRjwl5VV4YZL
Ve1trVLJJzTtXfjE50FdQguMPojOUUilWCzOLJ/43kvoAy+JHNimCmDj429XvdxrLtdPHcI2BuI2
xaSIMZwCAjlzEYw/dtzgqk2zKE0hTDnyCHFMdrOCuDQVlae3RVr7AZE92R1HbgDzECSzlD3+BFAW
FMguSLcA8XEZ/K9p+OzhVthl8buDxeilJ2DnnPaQepRu2ELc5PCGWsTm52nsh+Sz7M2YdxPCsoEK
PbiFdsYjtEFNTWPxB1H6TW1Ne6XRGs17NiXrBZjI7qXWPL4Mo9bfOywuslY33HzvCbIAslwiVWSm
2yYVghSSM8cu4IlkJa2OBR5wigAOMInk/koNlseRe1fh2AsY65AVjr+uSQS1a7ggXGLjzJsGqEv7
Z2WCJ+fubrTZNc6fVnS/1BcVXn4rhqBbTbUFdGNeGGpnrm9QMDy/GbdqmOwDREMdngKUoaOFJ6uh
7bsGFL/04XAg8rz/gYtnfZ9c7evDjAcm2uwuPJkTeYVqJLwChLXU2R1oh7dtxIRWHHct3BthNC3S
6wfta+H5yXWY05fOzSG2YimFWEScb8fOM4nLVvWeTy3vjJql3TMUH9cqxPhNSa3SVN1HfL1TyWHn
rQpRcNxdmX/O8Z0SspDTepfoZQIaPH3g2FreGIAXkFL0mAm91HNfwO3FIcQunj/eNzZ/xyVc99du
ZFl/4/5S2WIhWAAWxDK9vH5pzb2YcI0hW+oxKwe6IIjnJqyLqNJYgi+X9tEXarr23nKigrcGGKcB
5eXtMTOpbScC8bY/kSRKsk2h8+Nthjh2vPrbx+gBCVuNWwCQY2yTUHd2mykfG9TlfMrWEU6dR9+T
QM0EaGVXvCnsiX7tmoPT0uK50gDKf4V3SoUc/Gbwot41UbkJwSvFjgEpB64Bjd8fFXkO9nrQFPuY
pZQ8xnR4F5sO87LsZ17lgzXKqukL+BxcaeCSxMveKDpT0BqIT3OdyR1kwZCk7reED+4Ng7w8QKKA
fWaAASou59tmJQN3zFvCk4FRhOg/DCMI0UBCMukxHuO3TCiai0HoJ3LUdPNhL9yGTC+ni8k+NEJB
sYOw4UojgdIhQlHT0fDjr2imGv4kcLM/ShJ93aPKUIT2sOXhPvc2CGy7OKRk1cLZrH47yslUOpRr
Z7lD0ffR632h0ZnOIE6MaS10VIoBl+nmkP447VnWuIHV3+N0lNGd+xkWylM6Q+ytZRNKXF8jVuUa
RZy5GYO5sjjG1UaNuVWO0qC42IkYwofgi2/oQeOgViKwUhEYmxHz1XkEM2LygkK4KjTd/V1iIo1Y
1EE4O54oHRbtnXq/2RET45pgAf6vv+SYRB4K2uuWq6UBCLBY+hzgNSKWyGi+PBprzJNFD9sZPWKd
pMTi/YvfEljf8F4Vf2sThn4aY08uw2vS0nf+Xw5rxyRzOIOx3NjcLF5LBxJkeaCEaO9manQNJsff
xpKyRzdqtat0dhtBrUBaQi7ZhfL2GhoRz76AQOKqYGdEpvjUEHJy7abGUG5mau6Vy+yVUKKdidoc
gw69tTONchXDKBR5Lf2CRA8eDmWcK9rpNwAQ2KjK+CBT5miqW94u8JnWae2BOIfVf0NFm4nGTIej
6BFYT2AUbDrNXEeVmfxp+E7EJ1Hyi3zN6vLtQnc/8ve5B8MoOZ1COHa6577nf6H7G+gzJdAVHZNG
peHUUXH27IaeiEqTZEuFY4sWs3SspUKKpx4jT3pS9/KQSWPEmmHjAVSk6p3g1JYsFrUQ7PIfMdKB
+C26vctrtY3onmlzPMjuBXSVv3Y4NHEdXTvoxxlrwSyBiy52xuueeMvchQEvE2Qo0z9S0tA6IO8d
uQ7mGf3bike/QB+yqNhNGKoSL7oz3guPdibKgmcIZh8iEBGmxanNL4ua1/CGJ3cF3yhn/yVrvIu6
McN97FX1xbb7PBBe7Ay22k7pSIk5HNvjIaz3uu6+14lebROt5qOWE/hsTeA9uS6XoLRlBK153rw/
KlWWBQRBtx/q62s2f1RDbXx3PVviY5A3ifCOd1uHRKR0DD4vh4/xDXY3KUQAqvKi6R/4HezVikQj
r97Oz9TonucOhHwzKWGD8HHY4ISszNj2sD/ZoMhvbhJ8xPrUDSS/DJKeoB80cqFmkJHrNV8aZDVp
wvRt5SpwYW1TGrCqR5riRcF/D5TPJGhGQ1/uVEmaG7KOZcQBCIuDj5iN6/XKlOI+VnRWpxoq8lD5
tfIOm3lhjMIYCX/FGvPBdajcjovbWajbfFSXb6uR1hl42MytI/OuCFjMloijMrdkynUqdqf+QZ6S
VmkBV6pEi9ZkoQ62IlXi0oCFHw6XxFhx6KMwAX342lHmPhH8J2ihEdMJ2COQNSwiyhsdWVX97qXO
PMBZypxZK+hyFa7HYu9e2c/3LSCB4M1T7jEWatavg4VMzHvtb6ihm8YI6/bIgMJaXf9kb8pmHziE
Z3nA6Mu6QsP7HLW3/B95s3Z8aE7SA270V4Vb0DyBsn1SfoV3do2YEadMDhT0sphexvHQPN71M3uP
3sBdkM3KDibC+NcCyf24WV7EQkm5TnD3CRpyASogar4t8x8AQomZ/L/YZNN7TznZMqLQEvpp9pBJ
faqAvik69Wi4YLWagFHkfCgKl4GAJllTJmCVY+OjJSiadZyMksBNvxLWSGIM9UZj9j083jVdvkti
X72Gwb4l8ZUwTKxZoPDIA537zHkrMwGt3GowFNHcBoSZ/szOEt7uR21mbeO9UqtZd9iFJDspuOQo
hwgwt9HZu323dUkEW/PMfSa22r5I5Mkch0Y2HAC+tViErUBhuq8csMK5J7SZxHbuY5Gfm6EaD4zc
jDEwmqaQrol72zBpD2I4Z965pO2m0idUnxJcwZ9DsGkexStQusOxfY7HcCTPcAkO11AT2pPZJhtT
lGGTxFtruPmohF66fVrLbh+f2Hno4G95kx4Qr3CTmOF1x8nyocjE941auixctqyWWOlV0E1Keljv
sm7o3XQbWDZXB7mJb4Mf+kciO3oNHhRQ7clPizBxAe7ADWG/xoXNGw/5OdTePwiWCVpsvP5vTp6t
qcxGIemc9miA1xbvOwuhk7KE8WFm6VxFxPqC1mEuyzTmroRr/mRkPWquKAKEe0J4rHhc7v/bbaeP
rjjFz+C91zUy1joupMhLVePiHmOMuFUz0761ek1ph2k/XCmFDftw3oF+AjGkSH16MSDjTL9duhFm
htFzVb6tsnhL1wXaxS4B+A7DalnTOIFz/+TOKQt4kNVHE/EDkxZDKU3YQzhY4Z125lUWL74886JY
rIdsnPB+dt+42FFFIINTXkrf+oQbjnEO0pZZZvmRE/ueLazIrWzFXmp8qVdgilrsi8bQatQixvTp
cT/g+tY+2AmxR8ZVPYf/QDEaFvov4QTRQbVTVIqulkUelhwY7LbWEK0Dl6gYAubQ2JrKnbv/P9SA
1lo8uoaH3ElQVPO8r7ed/jKJxY+NUGlkjegm/udlf5ccG+BLWSMwsOMOaKebt7jV+WASMTauxYJJ
WEWnQFLBPbCPOnZ9uWJgSOIjqENMjtQQo3UbM5WYrnE8hshpzLhd3bv2Zd9S0iEV/BUWkuM+tQdF
BaxpB6m8KdxFBn+mf+YJLkkW+NJ196JFZoTdQTGWvDIUeVuToNxo5NXUyByxysBIHISEaPvUovm8
lqJNGGEpQeAK1n6lJVGJpHJIpqEi44w41ez8vIguYq70Ljc45cu1IoKxoyLRWjom6M9EMHn3JvGh
YWpsDJx1pU1anEmNvyna2R0/KTpbIksv4A8vAL0+I6HFPZyveKI/Wxw62GgBOtVM0eKGZlWT96Mg
NUepdJbZlLB4z1x6IMpJLycuFg1urzdLf9zcY88rJewRXsFkFutX0buv5rVLmb35Vx/B/s9kNPK/
R+wm5Ri0BHNqyKwaH1pD1TgLmsAO0DUCDqe8gZ3B+tzvk5//9sPUxvpaju9M1VMifLBwh7ch6sQ3
z7RoydkLhdZ12+tBikFk3GFsBCwYiS6xXr/MulNzSejPyMb7AzqWTZnGV/i9QBJtdzz7la+GwGCa
RLJyoBWhjtjX8Q693dWiVPJbjlYCOMbChCEz8R49l2MFi93FQTnffZBFtwADKuCd0KPUOubSj2lH
LyFQCDl2j26ecelPf1OHpw91Hdt90uEGxgFH4z5usplX/kd5l04ooTaMCTMo80C+F7pKUXV08P7I
DZQ6FYbOndg0ZMBQUc+8DPXH3SQQyWHIqxNjFGi63Whs+SFABBx6HGHdkN2+2yVd5FY/mhmynen1
A5yX6cDQwYVkxyaIraTMuwj6cc7yEyGHiiW4t9Pdh+bawGnIJSuN6P43c7/5fYJoOwN8EpLnhjua
mBqmajoA+RTDbo5BrzFYfexRicNpJagNkeMLoVjcZC5jabrE4LiANU5cARvoOfwuVIWFDMGgV8xi
UjbL2wyFlQIO8YOoX+cDKOgNbSjTGAi3U5Re3GHh/P46826ZNg4WQLgb3vB+uhiQJzK/JCNoVLd/
hR5BEuqfLDEJnqxX80AZ1GTycXUFQXsoG3bT4Ms60u4lVq+8PJV64xJqLdEUviD3NfWl2GTVc92Z
N/hyPZvWdJlb8TfhmXiLvWydrk3DSXavTHspm/O7i2EZnCYndbTTZzSB0xGrjCx73gn/eq8LU1ih
dvp2Ke+izrBR+N5gKPeR3cuLF2Pokq1WVUWzhiojgn4t1auQ5vv30Ru37kMlpIBaO6WHvKLUH0dH
ghTnUPsRxejAy1YnCo1AvJV6qFJPPiAGHQtzBhIAxQFNUmsR20B1WzdY8cBfIa6f3jX1Q6mjSuOG
oKHYe9jkjVeCNGNeUKgIQDu5qxJCht0nWcjAJrsYUNaKbXXXwDdAbqm6rxAa3N2dNriO61f70rgQ
ufZkKd7fUDfc+8GM+oA4B1R6e0cqdNzDkVFoQDD6r3e2eG/HXyji42+vHhF19SOaD9pGpVCvZhGj
rU/k8t7Fy+bERraVP8FotCZ0b87wvlSsda9mz59HJYuJYwfMxFxL1VIfMxwPsA5VsgnU56aUsTIa
e214oJgOFd9dHzS5d7nkGxgCK2W1B7oe1B9maTo8wN4JDsPtGBjVr0o0mea0tkju3JhIF7jEre/4
aEgBieTLyxAIFZrdu+NqFeid6uWUGaeCu5TOJvFJpB3d+8gZOpiKTMIYYMFvG5BbFPyobjPPNMvq
7ONZRqcgfm4K4gQGMri1HpKGtqPS1L2qIB/ptLs/bSG6rqUVeVhduZ15SCMQCo6KALStpDCjMj6h
wuFV61kz00S/7RplAKnKEwVfWDfu46pVZzjRpGfQ7QTn5Wme9KPu/6BZFPDykHSJyBAs1O/pHPHh
aI3Vx4C9z5i15hrH9M7PKsCr4gK6ZgJogQrKOli8RWde4mDlrnusfJj3PQxd0g08QTr8yPElAWE9
d6evxHN0+7jeid/s58vjybTaDmUDwppvBNviBkAd6yZK9F6fDI1VRxkvZyzErtaK/B2EG/crspYr
+h4w9USM2Sxi8vrtvgk/oR97urL5aqU1j16kgDvr/Eyu+zykBg5Qd6SU2GskwOVwHaNm62SBb6Zi
H81kszqbvX2Rs8LXAwbLTisxRmdZwqIyHjvYpmtdrRnZXHMddPGeG8f2ckPg3nEFHEp57v4EFpWq
3Ixd3WLJMrM8+kJvcIb/4gfSOc9aGEncgoEA2nAomHgkDFY6phZShZ43BW+JyYrWfMIdHW5ZrQOu
QKY3QIqnOGfiBZVLncQIc8UNn8kQvHZciaCEquZVyjtpkTTR3p+/uTma702rF2lZAiQcnbmTi4wE
x27uELpQ96Bb55+H5TqP+mEYVEOw2iLIdK+iC0i8Yh01Xr0ps0lYXlxM/cTrVHn8yD8UCdMvt8Bh
M8rdD3jilQdDw6eoe7sAZl42rE8d3jiFhv/AohbJ9YahJo1COonjcBLHsSEaO7mj8Bvs3X4nbG0S
D1N7v0QxaOCxXRDyFDk7U47jW8CXVMBZCRya5IAAR4MHPsbUcv0zGZcnnNEnljohLXIk5JIPi6kF
w99IcBa/C8ghn53oRxYcMErRMwJoHIM8C77J5Lk/L7D3aJZmQ4zpC3lo3rK3LgUlukdzvjxKkQ5a
CpAnARI/cVRXYl88joc0hzZ1sGPcoVm7narL6NLxIN6qQVNkk6bfDH2DLw9WsSQMICsy9ccLtzz8
lbosmh4Cp7gGr/9t/ibQJ49RBMZqjn7/xyJmW3G30Ul63wTqHipRdO2OQeB0rDq3sQaiHTezjDSY
Y/yXMWi0KVXzsmCnLL4W6Xo3KR5IdiytFCGeWag8FCDsxn6w0UctuX20gjvRP1BWTrO5t/9+aGC2
N+re05EqYbfp5Vv8vKiFHaeivXuwYzYDPAgLzOGI9AcOjZqzyER0As1/Ym8qudZtNdSTdI2eLxI2
jQlCdj1b8nGjmgqmLcIdh90W/A07X13QkgQEzNSW9x+a7jpD9OFXpVEWMfrs8ZGHUdwl8c8pCQs2
0TCF8BNGdFs93BRdtIW7HSQXMMxtkswUsJnk4yK/LemVN2XWQbczkee421wNN6DCv6zu0OgB9bJE
aK9tdi1SnQA1Xy7tZtGj97IOwH4D+UxXcU9kToLEPRGxpg7t3qMCqWbpMJSPDjAFozHaFCPmeVB8
bF9UfSeGe3IFRt4Nm1g+XYs1RBaNz0TbL/RWBr9LUrK35H7EqkTqvpoQL50OvqwCrSfg88g46Mtc
aIV5OQ+fenV4zvTTDCboR/0CgQBalVmdsggq/LMTZpIG7vPea1YJMB1Z9WA+Eg3QZ8QGdp7CJsL8
kCC6EXEyT0m6ivFUW7q6jJptROC4eLnG16FGpGO9fyJXQTYdAeQIoakFw4PZzG3B67Vg6SvZg2m/
BCNJqET9Vuvl7+IFI+IMO39Vc3UTOhQxD9k/jMGtfNvQjnhVjqzwyMds5fBIztTe9WZQkt9M8N2D
+J5pD1KyPCY37IDvIifmfVoDOm0mzsVk2fDgbJdnTWVnukMc2WptXe1rgWI+td6lotzCW/hk3kNJ
dkaEP9sz/+fV0BHFm/8aVcACz5LttkBOpxf1qiVuOO2eX6OIIPTKekZXEqGFTZSdNs3xtZrel/Yq
hGtZxQQMRWLjGzXvTB1TgWOe9DnVRE6AaHyWsCbrEK2ZfS20LFhZfeRpKNDNOlP8K7FyPFgl/Bj+
MTyNjnJ0ukD13PUfnuzezYq8B5fgfTj86HQYRI3EKecCtuCqajbtEnHjHO9igFkOQvowUEFJE1lp
C2Te7RpdR4J4Kcua4vM1kUsSCRraYgv3+l6Iq+sjBv0tfuUzzMczY8i0jUSHeO2RWA3nyRL/+rv7
NXtz6b2BLhCQm8LHJLSWYKkkYe3qZ/A55KTrPcW8iE4H94rSz+45o7Q7rtZMOIpoGiWXOunkpB4K
/+kEvfSDXpwdSCcL3z2epUnIGkr/GdS9V7qZsLx/sK5abRusmJ2//OFLYGT6i/N+yWRPI2brN5SG
3j+nKjWjX2dcuqXK7wHT/8OO+I4tTrekpHBrCYjCICMF78JGkYEh/5ZQqmoFA5w+H3Zp7hW6gnDe
gVn2lcfpUTI7PKDSvReyy2EEssJajZ7wvIlAdjlmUc244EQdnEqWc0RzBXXusHSIaSsccwy05IX7
QDnJ5BKfklZyhIcpsyIlLUC68e9rzM6XtjJINjByhyTWqjJbloKZCn+CaQqA5jN50vTBCJYQJ+lv
U77PNq+WT0Kd9TuBnBkaw8SRBOmXa5RlDB424XT8vnOgs23aNfbNt7/T8zbcgIa/qVyz84NnnOw8
rMrQ6ZoUXUarm5VNqClPBooilxMjIZQOsq8qXbKZRdh1velVc9KfAlrIzV3pqFjD+mP4DqF3ajq9
S5YBtyn44e78NSDVHJaVhahUt5rNW47DqFLAbAFKh1EypiQSV23CofuHV0EgK8KWUREiVG/By2es
e5xUYsDBwV1rH34eLrOuLQVs4F4lhv1S6pNn7Cv+DpS7eUPWTgTXdvPcnJr8odtGVFloaNEacGh8
sUBoZ+pNCsGBu4d2jIlT1zGTS74QTU/E4S64ZOokdqPW5CyuwCvhywkSs1l4G66iAxpAEepPAMp6
Dmq8v45tdGP7VoLZSZMoHTObhmKNAC9SyyebuaF5Tb5LMFuOuwqDlFVIc90lLD9BJJyAC7wanoBo
IuRd0v4byf9OB9Nq3c/gtIVviPyvj4BHbCFd8imLJVzL9vIVLsmvXYOWMf2ESqNHV44N4pIG0UT1
snN8itNHzrexnDJo0rK5ek+y1e6Xp8+ONDSZgPqeg1wmUv7FiXOkEvd09KRKbLso3xJNYCCi4uf/
DLqSfIC+Tw6lYEvGsO8KbjnNB2FyRpaXbYtF8xlrIkjQglMje+UYsVNcuVhXEImU8OxIJ11RC1YD
I0M5DVWuO+UEoztXS/aabvD1fLj3aYwEiOFDXY/deIdAwFR6EUu9RHQXdWuxkwAqdmjIcZFrVwo5
laHO99udoRJrq4onLiOzXuPOiZBNjRoOZ84Thjz55/FjSi02Uy4OM5EZf/1S127h0H0khi2JN9XR
RzOjJvs8IOlwD8aLPlcK6NMEaBUGmjbR4bq5wBtVeL1yNXgqOIvUslc8vbDbxLaIRDD7t4jq4WyX
vNA5IDhgI3pZxyKewZIlxZ6GB7DltX4muE6BRiFV7YCZjeKV8c9rbR8wnRNwC7tBMqWQydqzPYoQ
ttZOiYWCW9xnLfhvqUyfqjpL8NoTPjWLJRbik58sFUBleLoftyUwJXqIwwol1gJ5bzPc3j+RbkHu
n8HkJ6EKL763fNgcNsTaxJff02r0H1qw4u2JA/FZek0JAeYMSp0tzbop7FDHX9iShSS/1a2kqNWo
5oar0zkFGEaF62BClsqx1YgGdvwwHisXgddYvl0zXXxm6OERwTHivJVJn2NHw+cwwb5+X6q1LhR5
zDzmbvBMfUTQz/vEg4jZo59qmVFe+FTuZUos9LMAhvfrlo2EsMSW7fNs1RL72kyDhj5O4NOm7sUe
gfUrnDxW98Ha9ezYgw7zn0pCdHdC1nr/2bMXTpAGxk3ZKcksbvquwwAMYaAJ6GJXGU+FQnV54nVW
SKR2+KPSu6d6tO1nhv5i1NzK0rRHVzNrAWAltyM8zBGDXu5RfkGrojbZEdDFCP+cLDj3BWjwppPK
+gzJwxQHYyvfwOYt2Bm1baokQHFqVLXsjH4nsH7/lUAfgL/XcFkLCAg0Q1iXpZXPXswgqYtGZGiu
cxuqs2vAiJsTDM2UXYn4rEhaSwGN58tTlzK0sH8wKASEvCIWSM3jGqqb/Omj+SAc0muLTeCE3JMR
3wz9+3pRlfXlJS6318TxsBOoHK5ntYDI1ZuDJd9WHzlIg3Owh+4PQ/X6h/T1c7pRl3a+owFeAmBO
nLKv5EfbKZFwhUsO9Gla2daROxCsjCcV0Ic9eLPPj7qEtCLSHpmh1XLEZvDX6FEKhMt2w5DOCyVk
XMtCXZpMwYPI6jDhvo+/VP8Z/lwYi/L6Ko9v8F2U9DaoSih87R+WyfRGMb7sPag0KZe1WlQ0PqB8
Smn6Sd6MNy2iR+MclLG+3glaHH3Zq0QCNjUpajdODeP6UpbDAneB6itOwA01VghaLVI9ee7mdfGG
4w6gLf11PCwaZPMnu/DdqM3yZwKq/vVeWJ3HTMzLp0e1hIlhGD05q4p6Qgzy2+qQfhDa0If9ciOF
9VlpxE5XN8Hd43BKYnkUD8P7Iz/3ahCemDM6vWtQhFmfQQW85/k4rGv/HJmzcQVloqWOTgrM2sA8
SchbibmYWTSD/ig/nqf/bDaVTITRJKZdbzQkixr6YAtt/YfJD5ymexNSexdGI+OUQ9NcrUqJmHeX
b/3GQQHv/QbioJER1UjuO4D3ibeR4KZlN1eZ934FuJwgASQfGzG9bzA41syv4tW6UV/T/XndEpd1
n+TG4FbZqphvqUEFfRWsoG21wJDxSOC7X622SAURQ7xzZGtQxsMKbYDlUUYMBZaj7xFFtRc99fGi
dR+kyYBUFaVftAm9XJtDA14wUpo2KI7OBDpwaE8zTLc1lFJ6gXQCGkEmGgCit6w4/vX9VToBWYMQ
cyY8UnSrskTevjqyxiocr5Ugyl6okF7gVBaXnAD114LzMHvHD4Q1epheG3U/JjMQkjDt8zaDyXif
t/sVZyHMnpqXOu0jAkdewbErnzi2EjyWDrxPxbtzX6eVVxXB3yoUJ6fP2SeCGRfaHGLNHC5NiArE
JEovFGCWXbVCu21p4APCI1ZaHgIuWPsYifN6SGe2DII7FDbQfsQcGHMP0a5W1ew382D0WPsn66Ai
LaErFQJtUMZSgw72kKfuxGn0mWkYEoB3jIW1d/QuuPIi8yvh3so/m4iSln/Y7iiXuy5ajkTtIG7M
ykwCzPHsefJLJMsmqD1gvmfth4CNECyQBqBLS1/KowPJCkdSpD+s6uVt9kYHz0UxhDzxbfEbTUR6
kjmqYOfcXkpKpheTAvRwkcYpQ8lBV7aDK+SkXveGUCK5WM/5CuNLIuOf9vRNVRMwnCS9kkaP2eN6
0LNUOy3dkh4VrSNcvdiEnbr9/tas/u9v2i78GN2lqayY0iI3p0LL0z+n4t6akJYdDjW5EY5VzJi2
QWDWPF1uriIqqT5Zbf3pMdADxJA7dwDk8Dks/j4nGi+8c6KQAnVwxtxdLkGPjzNSAqp5vonTFkZ9
UTA072FVyLxESoUp8XMlx+gOKcwFPEdLkumLSkDi7tQxCY113wbalEwysHrVXfsl7uFTiuanS01R
8mTWtl835rklaHpFm6SC39qmTLetL0MJcID8YAy/SGtl6/J7dR/+UwctXhEceplD07mFB/qDj0rp
jESIHB04TrhlisBZ86wIo1va5SJN+ZRWtnbJI3FaorKgxC4nL12eXlSUBv9G0f54qejDh6b1mNOK
nosALjt3nGppCBuQXobXt4v18VbDh2QvA3QhmegW0bJsbEjSkzsGWDj9ToS0zQeC8o2cwjqF3gqk
Dvp2KZaPYTeHTjeuyj2/SzdyPESxHAfXQx3TfkvDTM4wVzC/ECrSb66CTK4ekhe7/nWqESdq0vEz
3kbl7r+Wzwcy9aS43K0Njpl0+4Q4+PMCFVTVVzKKFgvm/9bYl6nGpZsioSRf9kjjoOjqGTC7R0QS
9UdGvOcjx+4PrsVzL0xSoeSuV7vCbm+mbegyYzAG4sWdNNsIUXFM4GBgMCdRL1N/xPiNsOwYwSOG
kBr9yVWuzYEQJI3KzXiNmGRnYj3Dl746Bk2QTZAu2pglswnoJdCqjeAcA8HewiW9KlbXNoRzKAw5
Sn1jzcbKUTkpLfKpsdoAwsS4/kAvh/mGu99IipMBLK7mNQLcdMnZ+AhUvVgOUu5tndp+qJALdu/f
3+pmGGWHyNrTSbI9TyiCNkSEipWnpK7yJC/0lVJdo3T4nuLyijYzxw//zZFmY07DQpYApcfLEZFM
PHMHHbXYj2S9dW/z+MTc2LhO0wtsuMhNPLaIRKdcXj2RA+StnhaKYT7dP6SpR60WLTVeogvbplrs
y11fIWFg3msRR/RyK9jraPr+Bz/rDywbNb9OowsQbsezNR7QGTPO52WJRzaaNJvsYXnAx9CAkHAA
fFPw7+J3+9mXW1xvp3aEaHtc4oB2KAJAQ9eGwJLjJaQtRYECpBJuYarUcv01QsHvYWksbN7IkF3i
97hTH08Pm7eA+TL86JW0Q+Nc0ABCr24fAwgNciZe3kDPEMbrgKyNvgqr1EbouwnT+BHEEw/o6Yqy
aeatofxugMOY/bBB+5SAGnYr+M6YQY7zqMP3R2jYmSrtF5CS/U6yBu2qSzts9616jYzVuFiOcBSU
ierFQxwzgjjtLrMAkcZORY1ja4v9sjeiMN7FS4/cvgSNtfRmwuCb3jrjUKjoA9C5kez9+1ohNvVd
5vpreye7LFH1G+g3xM9kOydaDJ0IoBtIsSWgRYxTJgKYfEsex0SD5GK/GYmprjiJjs8R591TN7fM
dG7nRgv9J/yn5J1y9DNH4okLB9CQPWmnUUVch/f2SVUTVDLQ7jdfr7SolECOul8LZLK1spEoHZi7
2NZuC1qF9CphCOVGlc8DqCzx1YQoOWsSuUWRS3F68T1P4wfQJ8BDNuC/hs+ovPgsPeshJhn+0D9q
xXg1UHdkLdMI/TZwAE44otqVqr8VM5SWflHtfZI02OsCsGvN/5TI3djoKr3wJi8p82CwF/9FcWKX
D9iizrnVne3xpCl93/HBQ+2pqvlTugLtRAKCDfbjk6VFr01/i/fxLSMKyuYn+AcNr/YUempoP/XX
5MLAUjsCMuGYYbvSb9BHlsFmkfmNLINndAKTBiVf/HZ3P2AysKrDT+MbJejc6zSQSjo+fnolINdA
pWtZ7Ze4u8jZPhHyebmD8HuLKZxbmekBV/94ZXhepNNR4tVlyRkWbg9oev6nGvtkkNw3bySzWp9B
bZW+4a+t65mkfIlkPnz2PH68epViJVMwKoEM/O+41+ID5BdNDTJMtf3Cj6hewYR9ynikG16s2cjL
bcnHJ/DgWcB0MLqCIuQ14QoowYvd4z/pL5Y9HEy6V6bfkmYdNXzv+Xgfo4sIauD3lm3ix1el1MFW
gY+KY2debwKZ1TXR4L24YowgAq+Smz0jExVMZ/+go8suvbiTFIbfh/w4S87tKxtLDJgSEJmFzoRt
gP0zfRD+/zEDc34U4uLadsal1RPtAkf9lrJMyzaFYxfognQzQXlJcs+NX0KvjS6lHGs9/ursX5JB
wqV9hYIHWTEi19x8UaNdIiNOLzH0JJAAFOuJUHxNVNvcO3m3tVgG4+OxexNcIdXD7L8VlIc9TON8
ppNrIlE/oQZ0UYLs8YeboYxEVlRGUlMVtPb3iFj2ABN5p3TQtGjHJ4YyCuOygnKHXr4OBe4yKWBd
ygGuDo4OkBZFa1kzJ6XQ+wj6ei5s6HHvdGWM817S1hfSqTYoOVtQS9b+d8vCd+M/XDiivVlrl+KK
Qww688tT3JTo963f27bS5PahP717/5JD/ofbNzX6Eu+akiWmbeuiyt8bR5BoFxgoMx2rfVU2QraI
bpfx+WYsgnGXzGRqrLf6Zvs734krOMRmb7MP2uYKjw5DI0cY98CLFmrbpRnpzW8lY6CBfK3FNnKy
UBWJ5Lyz7CvVhIoOepQB+zaOB/V3JrZV9zuLJGalkYbF+/TioFFE3RN79yzk1HKtFos2KtVOjdiO
bZrOsBC1VS1mRjAK1+3JpINbnesXOez84a9UHGo74zEdR9aQdGF6PEJaXbR04kwLX7tZiZySFyHh
+INB0OOGXvqgPDet4qFXPR3jPcpbJ0xhNgosQK9VFzrmkalx4pvduN0ie2PlYXFLWQTjtxdhHMaR
SqV60ULMo2v9XzigX9Y2WKC0TNYP32WHDv1D5I/RF28GLJuegQt7zk14gUsp8c8tkRx2Mmv2g9Kh
OGN/62cKTGHjR2Vya8M3j02FXWppIKMbntyoCK5OGGl3nM8PV/9/4jIw6smQlzFBmpybQ+HRdPQG
0WRThJD6yfHqkzgZbt2jT8nfplJghLHnYZXzxLB0wJD1jz0o1vVTZN/a7TeVEhejDPQfQ5dx7Gho
6iyPDWOd3ygppGy6kW+FYvpiUBLBA27UA69RVYp+9KT58WqOWXuG/6nH1qDRtvvzFR+kDZMK3wSN
nGy2BfNIn4O86ppg+sj+H9O4bxL1D+lzWwuXSVIXKutbQ7sJXiqa5M2XsRvHjRIJ+IFbjWRQawMN
heP1rlDd1xZn6/Mpx3TTuWgt3Xj+0W280w8vXoylxoz/LKOJHkQADjit8+b2ieC2K1eTiYInoRoN
mKFhFe9Rm85ejVHgrahudIyGGmxzHrRKueTCep1ynxCtgWpb0+Y9bEeduU/DrkqcS9OxWFud7J9n
uqLMmHjSXwPYUk5U7Uz4l6BE0MzGdzxVbMlcOnnlp5HYBNfuwkEpv1Q0bZmgXSo8XcOfUJPYL+uG
oaVfDkWzGh4NczwsfC7CBKiitzC11V+aYzd/wvbyhl89fw6IWlFeHB4W/eQNy1S66LrTMjLexOXv
efOvFXIE/WyCVof5lrbX4ksO01MURaW4tekYZX3Iqf4aTfZMLnWa3VldK6+0AghaO/pYRxyNE12S
frbm+pIwD8z7ZTsPvXkpptFAlgWFk+TfMPS1wSm7PG+EIdUFLUo1wx48G7xJ9cV7YGJLvt3VqnLI
VQAAPtt7qnId6isftzKRijmBQbwL+XK9Tndod/Ylb9yg5jyvJ8p/QAtyAz5pGCrTZYVVBvP9Gtvw
b+GfgIR65lnNCy7ZrkmHl2zDThDFE83cTDdFsoR2R8zEB8N0PDGze1pWuBRqrF+bsI1Um3wV/oZY
mwCH5f08MIzmkMfXoupBwbztMmkQPBwhBFr/Taz2Lofp2RO+T6YDPW38+1mzHz7A5PF8zq6MqJFp
LXoFFzgMvUR6jK+GR6Zmo9V8MxdOooaGPhV8sRwJhEx4m78dqnArj5GSKyQcJShawwhla1Fso1qv
uUyRi6jXb+xfQm6OkBQplePqd5045f0zqTz8UBbW7ZFrKMps0NKu0A4+JDPZqDaemSHPReP5OjbC
9c6C/ddrSO5LntVlGBqsYTkuQFrN5EwA+jGE38FiI+46EpG3E6PuKiUxmOI2ZJHkRz3eRilAWZiL
X3yFxuEDx6xD1ZPUrQPLlOBJLOCEV/cfCgh4hwUrTRJAXozEwUYDf6D9mC8A35il9mig34npm71I
dKqLxcfh2QDwhX5wHxotxJtnhGxN+6SLgTz4Eui9SPsF8A1KuB3xQ5nUGm7MXUZ9j2WsWnqj4odS
Yz2cjCXOSeMB+HJroVwHwJs5ul+TocdsbA6XVEZIfp/An52QqejVCRIBOvH9s8r3Iagj37aRDj/f
sbN8+WYVhnINb9ln6lO42Y3NCgnunt7x11ktkup08pGPxvlcw+8fnfc8lxp9UV1wrMkopcI1hrFo
naMaF1dOAnKi3/PjGegXsu7x7nlnInNLTehP1BLkw5xWTtng1YhQiIvJN++gUo8dQBCAun0E1ZLP
3ERJsYEwhfpSPqw3Q6iyQvNZ5DrUwhwHxpST3YkijjdBcW+a8t4aFjPHVoPdp1zan+Gzfgraeeit
RFVY10N9CHoh6x4+qnH+HoUr0CzeRYbht5i3lY5zR2T+wQxIbNU556IgQ4LFqIFAXStK24ynsaiK
ZD9cLUq+sy7uyBWE9zhMSvHl36n/0k6AJtC66guHlgrmukSEpt4tNj7E0CYjzgS8PW68jFla8WS/
sgjJF+zrL7pKaWM1W8OxxUQl+Wj6bbhm3lDANPhkpRwFH6JVLfEmym3nov2Xbg7MxLnJXuxquBWi
3luETOaClzMCEpaK3LjfMUJ8hX54xtfEiPCX0QqQVoLRTw02NBgmT23R7GjSLFRwDLhaXDRpk59n
mpZTqANO4devYIDuj6W59clqKzNkwEqGpM/HoJQQi0YdUt4KfdbkXm0Yh48UeZ7En5JACUqX3PSB
P9aW4BdyuIaKkBYSpPNAxuKTl7IgU7Q95SZDBpz3tsstHjAN7F26sRilxXjn4ALIt7CoE0LfsRwC
mseQKomV6ZqdMg/2IUQTyzM751sc02+x+C8sLA3fDG8KTvTPc3fBUWe7tfJZLU1GrwYrPLBO9MR1
cIhL6w9/6rqVW9uXFvqJH6WUGJxNtqwdpXa/8huhufWAnKHHImyJDoiE7PIiBY1c2pEANo5t200N
rJ6XAgd8H+kyFJfw76oooDmPR6HP4NNmN5i9o4VyWAkh+GN+ptO0rnXC4fezz3o0ktcGBC4Nfgew
12BdIr02FwjgCJThhwnkpYrldv0c7fBPhAufQbf65cmFtF+P/xRcyKWbnvT0PRjIqrXxCTK6Yy97
j/Jl1qqi5SCq+URU/UZokWbWKS7eSpi8BanLjyOLaJoyrIRNDMTCmhRkBEkcihK0RheTRC+M1fWF
T7dN8ndy3axUF4NAk4h5FWsf6Gge3rMcZb1t/KD1H4ulHaCLfRll8y/RcTvObDbkgxxNQwNPXKF7
MM2H8CKIHjVb0kcc5DuKJC1w43eSe5Z+TxJBRo5Yz+MvtHon2eZ2t1qgnntK5yg5DcoknvfbzgDv
y91UFpF/2pZ6L0boiTOQ6s4NwgUTSLg3Qgb9VDspd8aR2AjXRpeW/fFMoak60HZuRL4wdHGgNiwn
zX/1GDcxn7fKN4RCTj1fBbfBdRAW8VVIka91raZbhWMPPQHX0es6WUIV0SyaCDoIL0AQiwgL8rm7
hjuA6XZRCykNuHikOfFOFkPe/J3v73VwDKs2EQrp+9EDNgYywpGnXWzDycRAGuuvl29H3CshEFNB
ONVIj7SPaLmmnAewAYiI+lcXc5BzQU2kUXvzCmmzlQptskPg27jmn+e/5v/6e8fUKul7YQG7aY4C
6rT6I06BbMLGInc29Ae+Ka/1hNQCBLka/l0oGTCj90Z4OB4Sie9ye7tHiVN6guDmX7tBHTlJlnDK
1Tf06wRGTqKJjcu7H44t0ZKZLAkLwnblNDvJmPNjF6e4+BwVvemKWTRDVjVOuUJKhYAs5Vz3e026
W/iw7B0sbptEdTr5bgJGHt2LVUmdRbGK412bTByCVasVII5y8DcfWYpqLq1cPB9RTS+Xa+rlSsVm
3rpUM/dmX1E4Ywflq9hKvk/D+2W3C2yiHS0213hPRknro+s9bZRN66vDQYKT504pMZxMsh1h90By
23ULmul0cCWhr6fybxlwpmgKHDv0QiorEAbKuQeAhmFxpnoFvL5kjHdjeyFdg2d+RqGCFEVkLtuQ
K9w+f/lcddYDVTR/Bd3TdiO5gGI2WYsE+AWPigQMBgLSe4/9ylrLRMK5aeejdY8t5NbVYrrCH0NM
y3PLwlrOTwvJoORa/cALLgE9t/YEVWyUgw+knbzGyCtpJ5i7AD74PjzCGRu9BqUP7YMF0/tf6hGL
uSHL2zTdzEEotB/5tjAkv5HUufSANj6gHxWGD+6cKDZxOttNfCLkGRsF8lYJgfhTGjuMJkjuUkxn
tuY2u36fxHULcoWv9xApjTEXxVpKOJw4tQL+WuxwyMWEVUIqjk7iD72t77XRBOsYPGa4vmRENVY1
DD9ddvHdTGE1tXuh+qb5DzMPxra3hXUSs0KBdnQItEK1Cjs2RXa76JXhXWmQHDl2YBWIEEb/H7gG
KjZefMSfQoIIBg8aNEQgHspzJ0/WGcL5kbQ2efMVNVOL3UKHV7i96AwvZrkXJWR6ttUn4X2ejid3
UZ/dJFd7r+RdywW8L/XZjNUfYhMmBfETeF7w6YdsMcbWjT7QkT+s59oFXgjyN9OPVjmrohcaONxB
1Xu9memHTzXgtwOhfvGrWh6Br5Zm/5BVrjfzu8No303d2PeSDkTlvsg48s6rG6RZmwcFhO0csRAf
nl8c4B87robFXTMo+g2IbGT/LbXtRs2gKQ+vDMPcO9VEYO/Oc+aYjLlLzpZ9Sa4vUDNHkvF0o7+D
sEj9LaLwAsEi5GPocalSFzEqY2asIOHTIZHLfqtdUv00BQDujBTK5GpDFT5xyT3De27jh52gVyvN
8ALB7VCdnMeSYprbrE7OPjm9cFcuUx77NOVFDjGAJoqnEs+gGYHCOOSyqbEuGuBr0g0SZAmLoxgl
UzCLcbp1njwjwJvkUPoOAS/DojZai5QKzAEFzWlaw355+WAurULp79vZDcUoT0b4lBI9z4cNuaQi
JujchH6NMDE4C+dkdxRa9Ln3vyt112zYXAgsrQU5kQ2ChchNUKjgR+yABuTq7lGtDzwWSD8OE+no
Aqq6fIVKLxfxWAy3/Gw48lKdhNkvpIA7y0SjfZ3xVsKnM9tThtgw7VzGlWWCc5DlNBqhzEIzs1N3
UdWtgZ9ZY79bC/FU/n+BtmIdVTX5KtNiwbnj7qXOMGXSAJNopC9x4dh6LxhfbkEsnOr2G4utiRy9
dqZjlmd8wLKJWa8rDKVJJWC9pCLAZVFbLu/6ETGH3Dccq9Sw7+rVyReteTOedjj2PI/7kEnKxuA8
vJrdbtbxf6mzDLcOyFSaVBLvvX71gSoSovnV5m50sOUngC+YmKDwenoqLPrxuIVKB6wXFl4tseWt
Naz+IEMRIfVm/RmQbMAbXwiOChe9zB0z+pPOgwqULgDEAkuAr9nFRnH68DIcQQRcaDQ8pdttQb3c
/+FI8cTgVR4uL8gNOfyJz8n8FvoPc0p9QXqffUn1Br6wMGYUVw0QP7VXeOUDpiaj2AoiBNr313Kg
0paXEvH/HAh7t2kLBVBmt13HfOQ58MEjzUWO4HJ4bSmhVwrzemEZVQQlVv4dPSKqlmqF6Oexqn/a
UO+XpytRLqOvNkxbbCKnl0xQ1a2+CkZsK+OaMoxP59xGz+I39iHYQHEqEuRKpf6b8RC7wOaEmPMt
rq7bbBqe3vHyBXkO7IwVbUVudAJVavkJrmBmmg+feMraqMrmJFYgvZMamJoxip+fygRXJFTPtc+q
d/sdT0YmuIGgFBgVb0KR0BNPNNEH8IeqPF+0WTquLyaqZuB4NavzIqf9cWCYaNyBE1ttFbFB1rQO
RVZD47uR5pgR4CYV1C1vncZiVvIqZUXoIDdhs8bhCGV1CEjj9Pnk4LkBEhs2jK9pBBg/JYWJ+wYx
QFTMNXtsBC/PILhMkcKopWDQEr0K4SEhGQhNkn5HcPd6phQd8pxY21dCOdgLYR4VqbbqeBAEo+de
yIGL5gHgxGmQK0/nev9aSadS+KctAWO8pGjJCfKBHS0abz/bB5GLal0ZcPbDnR0o2FyUWOkEbDIj
fwu5fPyaP/TTxUXFKbPn6s0uo6GEM1jFSfvjkqlE6uTB2AJ8pSkaABuFh7NJ2LRHMQUv+eCykhJ7
u6IFjKsb6qNs1TPorm8xAHnrqbjpKPkeUZg/LUe9oh2Okb5Y44wWlBZH0a3xEypFTMkhlBXIC/9B
1nA/+KilK97ZdzcvuPni8uTRouEVehoV6V8jPX5+iMsbqlF1xIV7oPS0/sFJFAkLPAbnyuc8oCDl
1kd4KNzMKZ6z5D/jS0yzaLPdTIQWQeu3Lzl36XV+TcD22g8Dhzqu082NFF/T+2UUxWwlAteoXt4A
X9d7mXeFB7MU4w1ocACwmrNMKZhhxaf+imDrUMFNZlsaPgNZm6hmGSkOBIPru/8PK5fBrgg0zABz
DTpjOy74fUBMV2EueQzcCVkYIaJw8AaEYXsDfnPIFwcsFOuFX14taxeYcxZ9H1IrZKqrc8NmMgcP
0qRcPTeREJWipJ9SvYo1aYAt3yg9gb4bXhVHmR2BsupKd164c0I4O1wYEg6iHf5eTqyHHaP0+757
3zYXSlSdq3SfdRbFGsXFh9m3+/1KCfqc9MAFfKSMdqHBF68yYIcjRxGlFixQGy9xqTovMeAwxGOu
zXbzNEd/zXHCivS0JuZkD3DQGMKXj3B+l7BI5gK2l/d/8qmcEbvpLz8SFRw1VzBEwDJ2H/NlB85x
OJVccXnytlLm9NnNpzkylxL9oZAk/boXnH+TkMqsSNXq6DBbpG5JIasCZQTjEWOquTERnid0yc0h
q4/1I5yrLjLuLN4DhlmaS7V52btvHdUnohMDBcW3kXSGh5/lk3//8j9WtxTvRm1Iw7U3ua2qMTkP
CuN2rWUhu/Zqr6WkyfJHAKoOsklTrY6DDZTtHYU/CVBEfQDtYIM7XdIQrtv2n+l7NPZKdo6+r8tK
PRX4BOcb85bYq9kptXFYVGs2zy1KUc9GOqaK2zgCpnExAN5EtiDuwL8FI8r7HXCp1vAtlyF8ETjm
qkkX6ELywY2gIt5v2ZIVX80rH2736gO5peFJAaNvC6wdHP+r/wi8HmYA/JdJq3mK+5mrDhJWSf4J
P1oqxroaCcXrzNiqb3kYmb/vqg77uMJ9Eoufv5R5NJIy8IP4nFS3jJn/PR3hCzCYENBZTsfl+0wI
/96ZdWf3Z1Vk0B+4oM0/diexZ1HatZFSLvcwNi4Yhc6gh8KTBDjYBbMGWt5XeyZuUelGAhQZComu
tp19RUpsa4N0t0RzmYi2H+t39Ze4xAGXIAXDRegKOTyUGcY0A+rELqkh/Df+EjKcELWNLcD+5RLb
hx7xaIR5D/pCM3IUDb2qcRpuWPE0+FKafw8sqYxEfDE/NoXWToak7L5z4X+aSMkFZREviVBTeuWI
nuM/Re48iTvJcmqi2la2ZZe5FsMNbtoGkz+vH1pHbLcM6c7t+W6m0j66jko8nYp0RvFK+bZJb7AW
/HoF+h/dNb7Js8dHUqglnEUIUb9tgPMLYadkI6ClD5rEXSBcsoJntwy8lNVL31Sf2kFDuJZGnxxR
VsoJffRgjLzS2wPSahS+7bIoB4bcaBmPMcuI6PY0c5U1jsYq3DUt8HKLtD66ebSwF7hzTzKsMHDH
NsQEQxnmhu1spmRbftRYHaBBHFZAVDQN0Qy7FFVMcqR0rwRMbWItpvIDEodMC9snQzJgD3TLvrT5
G+0hmr3BZgj+Hzy452wmZmTqwpwcfAMASHPpsoTNYN64MQDRazNGDmmee3BCVIt1Ym7kkvnurqVY
+4W23lmSmM1LQLa26pQxzuAWqVEpvKaUWmKwSjpBnh8C1OLb/GJ/+J9nh9Rg1IlouFpDW4pp+e+C
ut038pIvMaZRBBFJzX9U534NeEThP6t05W4pEHBvBXamX5D3vkImPWNVpvpYCVklH+049u1ado9L
RL/QqODTHpXycB+0WmPeFEoeFYGWmcRMylzWBddr1u52/OFLpYYjxe9UnARweztepGuujlgSJL1/
nlq0l42slRihl1qkTgBGqgTFvPFpPUt7VVqcOkK5ARumiRDzqXElnlPrDfw7dA8CNO2BByeWdXTX
ez2JvnOgf1hwjlOfNNV599qQ9Ltfubofp/oIri7MvnSPklP9cMEaIaH0xTeSb7OsBrAo/jUeSQyN
t64tb7f2Knz0YxuddUu8zNBz8S6kzDVWeL6YR/eiMc+9tgBDZBF6tIhHDixQUKeV5RZNAeBe+AZC
rAaHroUqggIqoozJ8jNOn2Ubn7i8pixuf0wtXQR41YLJxH7wEi1OqPhl2L47PZPn311Ytl7kZkBy
fofj/VcFGt8xfcD6dUc/dQKFYnpYKN7jZWaKreQJmvhMX8xyfrv0qmq+wJL2IGrdQfdhJmi2lgVW
mbJLk6zicBIk+z/bvZ7dqmL9z3RsNgu4ct+IVOa+dz1IAsS5H4mmneo0sSFTi28IgNWnnfHUi0Cr
XO87Aw5MU1MkEjEzcMyKJWdxbjv9Ki1YzCmJrE/oiSoIU8di3zZ9jZN4wNK223NtXkVQCSdxLiS1
YsF3rDIOV3JuF4OStoQtGRKa1Cvs2olKYP6Ig1wMjdA0L5pDIi9ZEsO2x7ymuAw8Mh3V2Ce+R4Q+
c3jnNLlEyVNRfQbYWPS112dXVQ1XxCJx5Yc1HSDaifejZbM89At5sMCu805LihI6w1SJaJl98LS+
QsgtvDLmbhABJnnTzdTrbDOiuQ/j4CoHS0x044aiO3SqwqbkEG8REM+q5lbdbG22yzd/UfUM+shA
K5ei7b2wiCEbakR2ShbRltE19hwFify+22tkipYFbfSlJA6UXkblzVqoQaKEZWpz++Y7jJk+sdfG
dvLa4LHGrl8xnu2G//ls0sz/48wu5lO4IQOZiF1/bjkIjoOSdKWc61M0MKFzp2rQUA3G1SKI8ZRz
KfEdoSXRwerykxQGM3bhK+aUCW4TpmGWhhGnDGFCG/ag07s1yeM2bKSyjRDDFAtHEE+a0JJTBxy9
YwC/zzETLwkmo4cLdNR5nkNejlRibfH1jfqu4rOhfjvjmDZGXeSuD/9LTu5QS5oNi09PR70fGGfw
n251Rebw2la2dGfr3RYAyLiildxaHXBeXJfvRv+c9yPmGXSVricol+YR2St4FbgY/3ySjH/5t/j1
S5RFX51DHOys/WEXfAGksNl1LxpSk1T1K9fNP/SNwYNbyABglMFTIqRq9Weu/CgvyQEcGuSx+Ids
yiORcczxzmrNGG0AXg2bEwufnSMw3GbY+qfk1gU+rfEnsSp47zJCpE1+Zs3+VOEba5EWo8+0/30J
m+tmJ5/voR2i8Wg+apJABgWJA1vT8X7brMNCBwZCHhv6M+EQm6fqJ2Np+SETDTlR6qFUq8H136hv
DsXejWWpDLkA4SE3FgP2y5vA9LYr1bNVUFs0ApEQeiVUolzftEjnjIW104su9CwvEtVga5HdYzcE
yt4GbZUqGQCfr+oJk7Xd58hj2/8HSpfos2L8l0OiifImYB8j2n9EyVXfWINSkreaZ5Eq6q1pMUDl
sXe6HAXrRp0ciK9+O/jE73iHkI2fN733ctaUDK6JiqrFMhGuiQbxP/9/rYEq9hkYPQ7hwv8utC6j
lLpgssNh9LLWVZiINiaYce1i5EnWWujaob6r8Q4HGmNWSloD3pUbU/7151r3Y1fqvGx2376obC/W
PHzpcPRPxADq06OYum7qc83BdU9zdQAVZ+cftlxa9CUTP3VIvgxtMs0NIkjykzgF1l68qKSY5Uq0
0WoOqBN3lnQ9i2TbXpefcMx68Y0cw/vHQPgOg63ewFc1dgNeAiGZ438Fiadkh+dgSf5054sa4rGs
voJUd/6cp9C/LWbYKRL/eT1wsRNvEmZkAOnY4xno7g+NhBkoLNYIDFa6KPmAEwfu2R2c2EXe/zLq
t0Nev2696XaBZQDgJZqh1DxMBG8yy8p/waeLvtE4N7ZL5nfKzm3O2cb1w5JkBitJa0tJX4ka5q1l
KyJhiqTq7H9+I7KTxGHejXovei8AAFu2pUYXoHv62zQPJdXscBCKWrjGxGs54tnfCI188ue0atay
Z++yfWYqvcolYLypn9ajBJ3GmVVmVBOPdcD65VjICUJNM//69/gJv6motMnRLl8/lSO/C9BNzx6L
iFhSRsztGgboO9Jb/tm7RW70y/47yER/CW4M2Xwfq+QTC5RF5cx6hbFXk4VDVSgZ1f2hyAX8Bdw6
stGC1IbR+oPt7dn+NkMhbjTEtvC2TOuaBdBKkB9tLbNEXr0xkoBcvXn+0+zhSPke5eSJM9tqQPAk
LXKYpB5RPksEFaaOtIqBlPKj6T2jPDPvAiA+I0ybH4l5gNnbH+N/vFwMrQzhS8Qz2volBObRAcRs
ImdFkl1Q5zZ/nQgJCddguje53fuE0TKv57dsE0W/3gcL9mepKSq0gZcpWCtDGfiL9xH2hk3/de5z
b3cBYImVt00f+af0U1EBy/JmXddpah4dVL2rCBKOSkGcDrByVchWrkeoZnGJ/VZS7ScIojK8eL9J
T7VviZerkt4THS5NegsVOGSRoQQ5MuBJIW2LyDtmQk/cRBZxT0ZvMQ7P+JCWdOEzwSLERD/bG1us
tX0JUIZFIg1MMTe5O8DDKH68/i4Xs7J54bwNO3JZwWcYZyHNjZuHgZ/3KKbwiDHgtzU5+bRCNDF4
VFJlzY48L5A4K+SlVm2EMl5e+t/33msvc643humNGzQIeg2o9a6eXgHP9k2l+Txh2RWzuW+ERUj4
uwbflZD3Hi+VKtGHI6vxk16EVCRUcHtOtq/Ln+8pSYDf0xxPsoImWSC/1cqEwmHSRAaGDS+MIeK6
/Xf+GAvg2ZOgQkjbBejS647O8mNomBU8q1qkIh8isgo5fxbUad77fE/AA5WlKoKjdO4eg6W2ICwD
hKqIGuu1omqFVBMam95ZNmJW+PWdxheHOwqUVLN6Gn5xoICwA4JDLDjVGwFq0m3hytr8vsgS9OaY
gWAdAoS+o/5mBm5iLKh3v6MBUCTC+U3t8/5NfXPijnxPyq3ir8pV+nqvqTvo5uXIi9MyMjetH2xO
VcyVSGfW2XRT8BwY9tom4SB1nT6FXVDx/jNJpnETs5IIa3crvfDyBBplSp8NX2631CKk7GvkZpdh
27hiMDrKLGK9bQ+iPs7CypB22kYP2d/hVhtZHPX7Ie4zuHZ7Y6kFofXVusKMb1OszVVTQr8KRGBJ
C8Fr6IAa9lfC+RiccGqLsGUqI9n9jArga/a2bClujRwT8uZ0FFjeoWewEF4dmXfj4uKrtA1KFh1+
AyPE4dsqwZmW7DDVIi+1rm5OaEJgvQMff6ew1uoFE9W/aNZYidrWk4D6shknKELJ7Nrooi2Hf+i0
z2fmlzhAtWWniXRYVrGEScBIIlxZK2YnvaMlwLVZIYIylHEkiCLIrJdkTVrKphtxf238xJCTvLrM
7O0hJGx2fZriOAnJS13nw6p6LKbRqXJK6XEsCoFVinBLsCd1+310G1d9Ffu4rtM/uS+RLkWo93Rd
ZbG/oUAdnj57duX0vAhDaoKDr2w9cYTBDFOiJSGUkkDhdRE79uYHwcmz6CUUymq1H3HwnmpVy6kM
aegpOsqT5ZosSSBEjirRrYOqQ/zJe3sifzHqQhC9+V2InyQdzxYJZWt0OYfnyrgoXA7BOhHWa5bR
9Mndx8rzSRPJuckNb1ft7J+c1Mkx5WtWbWOnwXRHyVCFQMkK0aetUZccg4KGvceISyVnZ7ntCKvE
tz8TZzaehJwt7ZgraHDaVMZhka6uIYBD28fbc1aS5bu6lgepsla02LpPjOKoM/v9B2m/1pue9Bkk
hCdJTH7fW88H9njahq8vEugqrknJFa9VGeEw1PwxLX1WVU25vQHIB5sR4FIJXO2QM+jk/oWBIzfX
+hGdtJJpND/oleRJepyDO/nOUb7R981C82hbpai7/PVQT1cGYFfTEf7HUNfs6IPSMFr6l8whHsNX
Uw1rBLIwz7w5FbhoLCeWMtZG3wRx2E2CEuxXCz2fCPoxkc/t3pSGYHfRmbIGcIzPZJaMBKRDo2tZ
NvB0BkYnGtNAyqD7W7OEkQ67LCGnkTmITDtJ3W2COkMOf45Vyg0G4e2pLs8K7hedgxPBuR65w2FD
CXkr+IbB6wgF86n8UPNCQUgqGRS8pDfmX3sug0GjOc/E5wTpjKahDzd5DrOEg8rtN6l2sEM7d/2o
Gr/G2Aow/bkDZ908dYbeIhRq+vI4hBXdmtlraHeANy4FU3kjX4Fypm0t4LItqptO032SXLgLJQuD
c+pRP3wEF7kp1GAT9NkfdGm1DS5Ay7G9m02wan1KpSFaJSrF3SnIdPwpCoTA0TSUd2wOR8qVebZE
xy7mlQvne993+i8T6uzeBOo9+7xPm+LEy+XdLkk6brfuL2ocYb84r3RyKCZf8KY0x/iAW4izqbI3
pkDYEkyZqmUYRIN1S9DTthJou/42rBGSiiYHiNlSJqHzeGQQx7xBC2XWpFygNUmwtBXKVOoINteW
2i1XwXoT/e7lTbK2v4Yf7dUUz1NDvOQSlsuQmw2IYHeeu6AYfzDbh2mTSmoU5ok27aF0jW0dtmrk
6xSSpu0w80olu530vmjqPeS5d3BApz+wPu4JUBLVPDjSiglpPZ8TEBmYzVfWai5F7l76RPbCvYyy
omCxODGOmyJryIiHxmEgMFhXjdf+AaWh5yu71mUoOwbgUVnIXB37mp8ZL1cC2OSUJ794XXqEmq54
29YwulfXfslrTlmBEbgoaEFxByO7z4K3GBzwK1TaAQsj8uYuaySJo2nl9dYvS+fcBRnnVSwoYAPL
HFuKUSwL3/DvINCUNnENr3QSOBurw4AvwRav7iVeRc1GTOeRv2tNXJ0/6yyFN9Oqu43urPSTe12n
m+/qnyDsa8bSOGHerclqnJA/MKd7/j4chBav/r1k9DO4AteaxZYY18+a1uatshyzDIej74eERR51
Wu2Jza5i4yzQtrtKPkZXqk6n5ceO/8RtkglzKqWAI2EiLUStF9AupPB4qEbywz2AAadj0H12e7GJ
RBodMc9IT9s4lnn1efDT9fDXyZa1Zz/T+fEDuujRiX1Sv4w5MKE849n+HT7eNG4SwOqIEh1P0Fwt
xrCeEA7N3he2oN2bAOsOblldljsWKVOQzHYl0gkSZFqj07bAxQc5FMz3ZIsgCvZMaPTTR+Jps9FC
/Qmq5eauzkfHJmgsWgDpkXDBItR59mmVR0ZaHZ9aGIfvbBZSTmT+5HxDs+GmL2DZrQpHr5yWkXZv
VHyitqMJk1VYagd76R2ruEkLFBGI+mADR09o42F63APH0nBpvHqwkZ8ZPD3CL7d5aNQXhIFobJ8T
rY0T4z5TSJeeXqUMXRcfiWLspE4ElA/WAS7cyne7tCQXWr2VdOm8nc7z9v+F9Y49BMMP4no6sPDB
vQ5mxwjuqpBKnsOKaym6kRG0b09vJr+0d2lnzXub2V4VLniOLQe56t+11Z8Pnuqjz5kbPSHUECrB
REnq7VFFXAq14qncZiULb09CFukZSoDKdxFQWS8YqdX1bmZUBF6ByUvWxHl1c1rKnAWJye2CbsOC
2uPa1PEXGcrw5kdIzw/ubZPN670dLypGR0N/Qa1L3iQp2QrXt5UJNdcJAgjb20zMM4X70/RyMJ9S
uIOgx/YJ8tUaLmBIG1Q0mu7O6baMDzXWv1qHlpBGbSN0SmHgrzC0sMyEXS64Cl84mwxKmweTA1RF
eehThjNMk8s9ewrIBVilRXbTW0hokXXAQkiP16GDkEMvGHpeMifn8mnAOCRRBjNS5SBmF8q683eC
PIAyCUFacivbfde41zgSxH0lK7V5dTWMQFWcPa/mccYMxE+DJcudUORxu2t1au99AijAucX76fiw
v0vV3noEO+/v9dzks0pFb7u9N6LdPHCdWPlmrJfrtzLlcFpfTLyFAr0tCy83jpwbigFSnCAnOkjX
XfDo1DMGcbCO9DAO/V9A81TzvP5MYeZNFNgQ29HDjkT0EWD3FxB8Qybahf9VC6YmLx4CJqMnf4Tn
DS/aIGkPrdXkAyIw7GnAN1g4JBJpqnPHn+e1Qd27mawmQ+P3bqHSN8FL+ew27LgEoiuIXR6jf7xV
NFODX93iGBuRs+54UW9nAc8UX/NPIf/PMdbVE6OssEwycZcJpxCm1cOgQt4FUujcRAHGIBRTYgaw
+OHZCPxXAT9yTEQ2iYKygkiR+aapB2Hurk51wCx098oERj+Q9tACNR+Lstjxol84HCKmRqIEFgoI
vA9g1yeOKTChS70xeowWtpW53CUnPkhW12Yo6kBxa5GpQ7GX+XihWkSOGC8Ru81x5fhOaABGVt8o
Klf65Dcy4c9uSlXBL5yBUio4CtApp7Be3lv90BroBvduPvfjDPrtVUun2dxJb9O5OAvBAn90/kMY
xUAZq3saIUSr+KG3Yt+EYx+KyiCJa5fGPYNsyw+rG1LTtQF2akpg0wXfpaTZ3SQKnMQhfTZWiAl4
zuXMcUFPIDLzUYdsIm98U0x8Iem8amBBomTaOAASYZm+FEckkPVzGmGI4V2xOIyim+6Vhl3Az/a6
jUs7jgMLpXu8ScrsJRexvPre7/nFDED4maRGw9pUfN51Opu0I5d+rE2+sxdlXadZXIRFnSUn+EjC
MEUwccspzy8go8ssR1mD/i5O2iint0EntUhsALT15Cmxz2mG8v/qdiHjaFSxfKJfkz48GsvPzE//
dPFnv5X2kwEXnkCkLEq/G2DP4mGnDILHO7U5yITcR47SYfH0x9HEnSmQ4tIaIq99g0bxGHtnexoS
kIByK0TuXf0zf2hKJJdOpPe+ojLigKMKw0hAphDfn/9OfCPkPvJlly1vea6N90f/EpfVCpjdvD5+
V1jQ3hPbx78/Ejgip62Ycy97G4PbZH+II6W+C4zr2q0xe8ibvxM96aQb4zMiT3XWWNRWnd4MHDPZ
M4F+Zhigt7KwC4lOSMmm5fz7CgcxM+R4b67CWenoX/Yj7DDP7bv8OIEQcbtpYDNSdneWyS9pgprr
XWqEhI7gAzx8/LjfbrF0I6xtV/+L4FdHjyZoJqgr9LYvkcn9lPa+wui1kFjQ/ybnL3HAVer1nFwM
WfZFHZEdm1iRUm88Awq3gpevD0DFqae1JybDpEfIUHsfrZaE5jGw2oZFSVcGj1YNydnrOxPdLNE0
3jT5ugrNuWaTYXfVgZT00kmi6Hoj+RrooFyCSrQ6nOrQsZuVh8P87iGRaQsWCylPIQCdHwyMq7el
E1hP09Tbz7xGvuApejwZIvSJDsDFt6i2W3eJlIEc3QK2eV39flNzZo+H06cEK7tQoPHbEz6LGhJc
LMVz/rKOLoB5R9F7BrwVWr365NumCdNJhDvvKB3NrQwhOeIki40N3LblzxJsJGk1TSL37lPC+ffd
V+xGQgZNyisXGL3LCh4WuSMBxvxs+82o8UrYNH8OkQbQfUqjYiJuFaslr3spsk4RG8cL+OMNrujX
8cxat/pvrumYHaYDLcRC3BSqOlLRGIrS/0afGq9bLnubU/DHst6irLZbRycaCSX3h+Gq29aPoes/
RTFlDUMuRzclBPIe07toj+qa9gazhFtNES5pefwJI7ZcrFXMKhhOIex/HCU7KVab8Vfv8GvVoAJF
4GgkXB3rWPsj5YAW7EnEJHtptWOff+ENa44owfFqx5cxWbLXxJlcXdfLxgOxS1SBmsRQ0ivLA3Rx
4OTYIHVIkoGB86r5LKIF66uUH6TjGX0Z/e+2gWqpWhtTu+OgY/7Q2ZTBfKLq+QU8ph+l9wJXqgZ8
AmfnzanYx5FxO/ZrWVTXz3EjRqemhxyO9RpJD4oY7XAbkMsqRivuTpsWAM/hJcqNDvm+KThzwvM0
qEOdivdMdviGes/D39837LpvOCx4h1f0IJijJ1I0x/+/PSzeZGBviTsShg2qZ+Jwsmzrd42Iafqp
8srAAJKnifRvxu/1TaP7lQIQ3Q4Pz7/TXHURYSWXP2S74Za5N7sTfHmj6sURxkpHgqyQL3nq98wk
PqbbvWINHIoR5Jv07HCyXVRRGjKSWgEHZJQ4veN8VK9PMeHwUACDdKO2LWqaYC8iGmao0eIB9pnI
2hGTTFXzITce6xuLyx9d5mb5E3sAkFuZ/6vCilCUyxt8xV9nPomOhopl+4b5rIrahqEJ6rbMjz00
OjOPxw6RLp7MqmPD5mvQk4xaRxBmzRjjD7wQhVTTAqHSWOPvUK9B3bBAPGbVPdi2HkIU1Pu0JFZM
/X7KOrfWXGQqeKUMH4A3TwIh1YdMOxRrO4HSxBUnJgq/g6pFemwlo2jLKNZmkG5Gzo1IhvNfqWgt
5A9NZhVN+mUSoL5BZ6SXn24H0gC0vNfGvclsu9aOfE4Yhr2uyRoN38ibHO3t3vH6T4XQM92wAw/U
c7jtIOC0Ml4gr0+EUJwg33CM0lj1WK3ONVy9rUAb/ZmIuRmibBDM+Xs5tumF8+s42tDZYbgyYjcY
CBbK08dCIuFecblg97y8/MybCGCCMOu5KdCD3+nMmDgOVGd0IT8M8ztelpvnmv82j3mNl5yV0zQa
RkXAbst7giX6ihxlne/Av9BVb4C6qsPdW7Q4snhf04/h2NjPheFVD45uAVDkaIUmeReqaxQ32tVg
qe8+c4MgOpmMNq2KwnYAXGsZZ8YZ9rnnWGsRD9+Qd5NGX3GtluqHYttZW3sce5TJ2IHbU/Xl6Jdb
/z/eq3T3DLxTOufdTThVSFdi6l9xG7mFMzUNifGZH2RLRMnWS4IwFgdyIFWvXFKv2DTSp70Dqrxu
KJws+StuPZJfsx5i4RiAR72dZ3B9lstQvjhUMqaARz5GMGsGZ6RcNX1zRHjVCvDcqVe/mb8ZrQb4
GL3HhIVF67VJISKwoR8u3ZzfKT6h9xIUUrxfYTc+P3l3d4Ouc1vg2BZ4tlA6XnFZy5VhWud9RSqz
w+eMCIEy7sNVUVcRbHY3oyEPeS+7RGPbO9u0HgBPMZR5ZRpHnooCG58CpP3WFG8UlgfmfiNGLsiY
BgFECLKV1NZJ7gyZ04wz09xoI3NcXwQnUfTEZ7RjMqVhx9NvVKU0agFly+/ovQrdm/KPgS0TV7SF
9jEcmsVyuDTwcm83FrXo7Rrx09iMxH0d614OR6P2LeSQD3zSaCAGNLIuut5yo61bXMMEvPH431bW
NcTZj6EErfYwEZqGQqNBfhNfYF6vAxflVw8wejl6cVJM7ytTgDfhK2b3GMrtjnVF6RWDaJo9L31w
gwimRIbDK8qMbNXPfdMCQIH3h+SYtTnqCOu5qSEPBPXBSuek0FFwx4WAS09gCFX4YIp5VwMUYipj
cCsjz54k796QlKnDHbUwW+msR7K9QljLeBL1kuvvWQeJzzy8AC/QUQHrluaPpXKybUE3RxmmnfhK
3seP70uCoa2wS4TuocqFTbp7wrBK/PQ184v6dnul862yGsbd1/3KKQG4TD8FDpmbdXtOgZ+kFfx3
OwFoDYBwTyBFPT0iCtcOJ3KgJ6PrXDtgVJ2pVImPjQIsV4LSJuNQQAJRG+qeNJj8qs3BflAc5lGa
JBvLtYdCwijijnPHuwXRC5jKwHfPXXPfT27QR4ucooLnSIiddL9g32Ec2niPzQ8NrlvpFc3KiXb9
Gq1j0q20gJ13FciCE7zNvCaJgwCzY227c1p3WUbqpoprYQjHoRjhZCL4wNoDMBo2ZwzBiinWknu6
RVKAC3WBBa/C9GiSIgtAzn4JH55BrzzrN9U1lq9qoEEfHA8KQ4lc0qV7irkP9jYXZnW1CqGt6U56
qcYkon7GGWDdsHczzl5HQgr9Mw/RsODfFHqBtOmlAHzRXl9YFNvviE8IzkZTQTQMpHrrDT6KIB0M
i/doAPtkeMEB+E+Rr/65W3r4DD6cQQEp0qYxB7ufFkDplzDlTwdz8ngW1SskVAifJHp1/dTzAy6r
imsUSsUSzobxSxr41YO1s0wqv0G7b2IqAp21n2DO/6l63BvRTefPUMbpq1tIcRfO1NOpoHu/53rd
q+96Lr5D2kZMsNODKy9RzwisoOSGREKKedOSCBxwIYZdboR+oV3JS/OqAIcaHOhLxVVj+9Az2yqE
ZzRY8KpBSMLuYqIsjx+LZHhL/Dunqor7Vlv5xqKWEcpO2SwuZseg4HinJ9Rg3K6h9oQhVb/1TdWg
salqEUu8p3w3J4dOg9TRHBxKNLnz3gqjTbPHQViqZ+kmoq96IVCmAEv9tbbMeombQOygv4dw7mf/
AJ/Uxjx2xybgLeDb1WkMyxprSsDmekSV+Qs+aV5SDB4JRrdFf3Ekl9yGYpxW3zwuj+wDuFLtQc5M
ttkpdjKxKy11+3OuvZm2xtpks86wWXVQ8yR5qdIkjGtAa3fTdtUmXCZJ2U82VSgHy1Sfw/EuqkT8
X8/rOYqA0W15aZsxR2cyUYIoQ+Xz/OdUM/q6eWGsZR1+wPjA8y6voiMUVeBu+SYQYxjZiCXYjIXw
oxIC5YoRJSOplOO/SVqpMasHbbyz0gpt2zEa37wXxL/c5Gif2IuI81W2pqnMS0KEWYmzIuLZvr8t
cgH6peh97BTq9eSxyENzdI5vLbrRv91K8CjwkQkV3xnwBrBdbkT9GglGeitGapKhocJtQTbIXWsf
y+AnveA/EqDOxEgsx9ycFCgRUocU4ouD+S3GEiG3uGSjiF2xaaGMpiK//7iZ/aDmQxzVhur8+XQK
ALCdwdxsleyKotAKg7OXFsIsa2IsXQtszcl1boRYP9ePUGADL9j1AG3CVigLVwulFlbJwX5b2+ZH
6Rb/ZB6ahTFRONmlBYN+Iy4e04vWpnujjBmnQ81YlOYh3dj7rN+oN/Netr6OyjKnHb5facoDV6mr
TEmKd7MxGQptO7NX7kitHxq+DQtWoSD5WBHqk/0vkI96MuD734NyJ+TZBJHrLe9OOTrNHRr1l4xD
CdV/cvMJeMc9KlASJ27txUqRGsM4xHsyS+bG8PHMrOaLnUbtBqW9faF6qx01NgFocYNifeaMkpaW
UAScpKUib+aAqE8Rln3ZlN6+wfzVW7LSktEZxUEU0sSAjccDzv6XKi4UcPaGYKtX+j34XRbG3X9q
yzBxuLlvLOcj+GfoI1e3XK0pkwChDnZuEUG5PDe53b8d63c7XtG/dm417KP5Djw9fT5yjjXupvjK
6JVdPHzk7+udvGqA0n4SRBjrbfPo7RG4w9Dk2evsMpq3txjvOMgrc2UqNTKWJv6uPL/Weln8T4Et
HIxoBiwCDTd3abt17ysTkEGpVexgk7nDESZQlPJhwopzYQlh38PQrpOi1rtYP3Z6nYTmLPqUE/BF
a8gU5r4bxv2PZRvtgmrgs1VcRrAXq9fZMBwROnxxMYDhMr/sx6++1jAl+Sqhkwa+uZG16xae8MoE
x0xPaG7vH0qGgcX31t8h9i044xvYu+OOehXPv5NLPR3dKlNz8GIsubNzdnvnyZ8PLzeMX2m/UP4K
hLrHZdFGW1vaOj8yyckiFyw4qT0dbqqKAxPZdGP4Z+y/u6eUm3TIYfN2XH7wDLhJ9vo4+XV+llew
cESDxpnf0hReXb++lbTgaRJeGi+i4LYZS8rreEotY7jNVfOxqESjnlVY+4pWDBEyiT9YkvZmBr1x
ODUPYQs3i5pyAOeCurJeHmCYDXVppK5t/00g2Z+tmUSmmJBrqhTXn1tFqqwEn8UonmKeXJ1uUAC0
xv0XAl0BlH6T2W49u3SIYIujV71lS5JhXS13Fbb1uv7DCJuy7jjtvHX9UZbic5/SHjvbkouTtEZo
20YsbjcdiVktF/rw7qfIEHPlXKD8LSwH2XnOgINRWmHeA9RTGULk13r3kSG0lOoNkB/A0jj/yGZ0
JY5BDzUPfQYlul68HKsN6N5ltnzHmeR7WEEnM0xFTSKF7AXrj+Pz3jrivESqG8R6Ecfp5XVQwasl
RymvIrNPS1jeOhxsUPltjUi3HQ1LtDbb0RW9MgUyxsgvDOyjtLTexIyjZanZ2y2fU/pbQxqw5W0c
WeFZq5Uk0HfjqAO5kspBz0ePmpM5rTiKAlIZwmxC/0IyHW6kYqJ5dLHEEwKchIxyrykHxNcjYms9
J69qOek0tiGLxpIyYFjSvukdBiA4JYcScEMLaajbQALdoDNdu93a3ozaHxRI6Kh7QRZ/sSsmLcDD
9NVGF6pALpTUpKiQCLyFeL8GkR0Xf4NPtbwkuSaInaXNNe2FUaQ3PcD/Yzw1iLBzd/Yr2CYZWcUo
OVC1dgdRRA0veJmTCKSIy1nfuhrcsxyALuC3hwNZJLmqLDfI9M8zef5KHwwRzj/of49l23ygVyG/
rd+CEb36gtN3Ep7zwBUbJ11yfSH62jQaCMwci3x5iI/RYex+P+Vsz8qoDrsh5cwOT6nbQD4bkU6g
pP+jJFUcu9KTdga2WAipx1skUEZS/Zx3n72TSoNGjtyqFjPuG1tX61LPHDfPpt1t7qWc1wBL3SKh
ZczvZ1I6o4+DIXK/hb6OaBQnTc/8cz4jC7WL1GSoyRmfWN3x+dvkm0GREF4lcdHjC0+eyUbwur7D
WNSUHvds6S5XvIauEQhDvFQl+EPkMGmkNFHhst85tRFuuxFyjmtPakE8P1Y78wcsqsWcwZZQjss4
/CD4+mi5BjPPPqlBJqLy8h3tHp1+EoSv7ci8CK/xQBUwMXmyjw0M6dbq1XWed2xG/e4hA1/DvoN4
bTgP+ug/w3VRz6JKXO+czIkDLV6zjYCMHsBxNVB1HywK7nz4J8++zB401WqASLyxOCWuYlt1wyOW
iaf1L2FUS5WZIDmjiW0eSa0vUNJ1V+fa+A58qdK7/h2XvThonCLu+IGzkr8Ls4f/Ubs1GzBToxaw
fvErTnpeqaEpcRMXYdtvoep852AbS/sxexD685W2EyHD01d/zW4MF9LYZZKBcgZoI+gM+Kaq3H7G
pHtkuv0z1dNpSQgFurFqhJx30dGcDCgomzNYmlkwKhgnpPJenn3FHcuvTjEijRqRo2sG7t68aOHn
u0kiI+bQ3KUPSRZVATeVR3xC7dxg+sYHYZqnwBVnNkDLLaPspFe0INSqTCs98QbNbHaH/xCItOUY
El8Q2ZTdr+bYPLT/JhHCyi/hR0ex3GzeP+v0OwqpNoAlOB7nP2xeLj9iHiQtgCn70cUpNPIIeTFT
D2im2WjOf42BqA5T5zh5XWYi9OizdhP0KutL1Wvlp12inItRIlcsWqKX/vtyvY9szfTfIAhP+I2I
30/y1SxX5PnyPmGXlk2l+/q9QeL2ZPE19agNx7PxZZDacsfJtHVXa88CsHVQ8qv3MXFO3UgFXOyb
QA7WdQhGq1olzpIwxnfPWseKU0ZYQhpyeKRnYUCbRSc1r/ehRDlqK7OFC0xezT8J6jZeqbO1aYLY
ksOMw4HVj/xIgUWsXWlzQ+asYofSf2fPeh94U+gt7kvCdc5lhPrdlFymMc0VhiEOWwtd7q7wBS4v
y8Z8mxzJZkBeKBW50kKXuJuFnsCfTwoxO3iXutqq811Wck5L2JaLPSRT0ZMIzx8jPjEspwhUJz0+
poXoYUwsGF1V8QHAaP9Pi15pvNafmyx3NZSC1OSbccVMM4PqxOtB0AGOHTZCchE9rRlFRkf2HLek
bKntoX1qO15zQGNAKLUCb6HOy5dfU31TuTCrRu5xTvE28m/m187hdZmb5LMn4Y6OD/mu2ty5meoJ
UEreHU0ByyWZqJD97O2raXeKCCV8yXJwRQAeISBW4GmZXVx3Gfi3ivME+4KhzLSIysWct+6ZQOf4
dwIQF3AMBXy7cSDa7281awL9AQpE4J5NGoivH1WchJogwAzuP7dOGr4/G315nyg3YhIkMj+9ZjG8
TVUddFimIc3o0dpiNjOln7EgpxL/W5hVkrfqtZjAMWSdhjtrpxaIC9x/K8+MT7Uw8SN09sbdsLlM
freFmrLbU+bruVYVTlYRcJgAHYMv4NiZXyTChFsr4m0M7pFkNhRwqcSx4lhFtHyDvBNYL7WinQFj
WhhkzymPMg7ITD21jFncpRetbhZVIMdMwiAHmh4B9FPPjmP5prJ/Xqg3bFGczMU7mVZIQx+RaOMz
9Ggn+301eG8G1EibnCWIXyLHHZrIY8405Gp/9PaNrGiYSqP5y7zAobiYWXB8iCTPcn/cW6KcyXFw
Cr6Fs6v1VjJi4IYyHqj8ENZGs8ItzR2kdZLg1J0nmEMnHVq+P8G2u75QimJOuOkQMQWKofQIMpdS
h1VcpjH+c2us95qTY+zyO19+675SAulyMmUG2CkNysL4JxsZUV6jWX3vzDx8/fxTHqixB0KYMzKV
CUmj2FlT+24rnpg2s3pTG1S1ULqlM0UuKKFKN6984x5QUk/JnkA4lZVNm8sgCNPRu52SgR/sacgT
hT+JVNU6f53Ir6+FUGXxDaz5mP2pCFH3F9mzkKvbqCzgAXcZlDToyWzcoq2M21l8nU0ld6mc7DN8
KPc7Tw19tRwvfzV0RO4yX4BXKzmEgWahz3gwKqPyckpnmH4SYGMdzZM1hJaVm6UHyrghWHlz17HO
WGf9/zN96uyw3tDstyuOXzDCfm25ynUZY1+A9r18Zuo2Jl8I21gu8e8IaklmPoguniX7DQr0Kk39
oUWZ160rKtBnCZpfnNZlQlD4967ZPcXV3Jd8ttGIbtlOlOo3AjJRn3ljqVuQqMEiTW2MfXFZ9lyL
Rb1vRpG+Zw/fKoq/nuTXikGgPaoDppihJkqF3Nr3dfZp6wopc+SKk8snMs+KhWdk/UqT3ayDDkIe
o7iykE+f9FkqJu7wzVFR0+yM12D305c1g1mpM/SngFTBcQ2C8Hizb5wbOxJ/xXmPQDJLjpxT21dk
DNTJ7KwkhNvv0xOrqRHRDe8We3u/FIyCb/m6qAJN7ATXyCFDujL06b4JzHOvgpko9bCtllAvB3nd
rzL0NBz3OTj5RzmQpT9bLnsRYeJ9hCkhPjQQZHMF99n79CKfpOYCzbm+1wLeAKcJsWkENQVM+rWY
UZvHCxKE5GXc/Lsn7FGEiDYuNBaUH2hzHN8qLv4huw0V6Gbv7JUQ2G/cHH8NFzsugfJ7tOSh4HqS
ep918UkVmR8TdfVZZC06lZsAjqn9wvcND2yz6m13WoCBgkAy5I7IYPnr0wRjoXlMkvP5W/zp2nly
xaZtGjCjKqgKBaa+4+ffHb9dW5Q6XYjfGE++zTfbWZHjj2anpnZoht2gqpuB+iYB2uKIBXafvJyd
Y5ez0+atrLeta8qkS88cP+PKUBw3hIz9LbDCi0Bk9hyzOlM/M/d/w7grBgTzNQYjGwnWuQBbdNY9
pqZ/Yh+RJhqT+7pKz6PMxWBYabHbyJ2naxfCRGlH8VfhCxIwgk+Rkrq+W08jnA7E090pdsH5179c
onL2XbBicfjXTZr97w5Hwl2pCIJmnS8OE6rg5Hg2FVKlmCffLZZhKPSStgm/TAAu6obFUTpgjgQy
uENppc96cj86O0QFIPQAagwz+8swYADQr5qrDYkdM8yZhregFPuc/BOYpiyR0pnWfAeySnZ4+G75
CnslRi+FgNq3OQZ1zkRZY69xKUKonLiBrotGroz5xlJypOI2RQluOZ7lS9XPINcxrcAknqdB6NuC
0hS9xnfHp53W7AgNkze5jsv/hXEj7Nf9wJKd2I/8P406JEku2u78BMVo8yg1z8IaE6s6iPUjNIXU
o0/C0ud0rXV1RQrPPRXPflYz/tF/F9xLvespsk6VfyIK0sr1fIYk4laI7xm2IGyv/8iG2y1p5Ihl
VRe4vdCComq8WhQIi2va5RR1SwH3EOEOdjDOcfm9lypU1Uavkuh+wEfepyBDSIUjq6KuYdhRMG7k
3eYigBROzlMX/QXQbaPQEILVF1uZb9s0YtTU/d7ZvTIhykXO/3eDhwSoVGvKqGd6+46xW+x8Rras
ur7LUrfj4uPbTmJSU7lKCQqqTpith9EYIlzWGgDjZLboK6lZeBr68HsIAiwDLdb66jpGyUtqIEYv
d2rz8B64YIf6WPdW0+0c0WBdOAglpabsqPZvq4t9aGG6NN4APdejGLCPPF0s1OV/D0e3X4cJa+Uk
eTbJQn1oft7Goaw+bm3tDRDXHksX5BvJfZYy1KgDUJGPuZWUlBC6ScKKbSVV1q7NCPTTp1ZFUcMz
+O4Onl6oo8Y14U2hsVYuColcmaqhHPbNhBlnOssBN1M0kuG93GUn/Tz/M3E6tBvloEUkfPBx9jnp
uaDUX3v364pftOt6Nf76Qn4fjNNR0dF4jt9G/UjUUTWk6sTDcLUW1laLPi0842dkPI97hSZeMf9F
zM6oteRkhcmOYIT2+UClSAEIZi6qitbxxckgvcpgrQFeVaTnmyJpUX2nDa1BqGDoa+rSF/tSLuZY
kwZ3pkAjA64mHmJGgp2Tqz8ugOt/a2D2U5/HGQ5LPn0F2BMfUwyuPS2W/cQwjYhmBBqbcCbBE9K3
U7O2qgrFZPsUf9vmFkBsWz7o0ASgCtCHphg/9APZKuBoS8WbDXH1n/iGn0yxlQKz2n8HE2oKN6Zw
wrG4DebbK26Af+aOOdgLWsdvjUEXZ/gWb24Xj6WqqhCsrixpTN2L0U6I/QVafDLC221sy27YObjp
hqVJ5ZqOr7Ry+OUXLda2Y5K9XPTQ2y7HtS3cGZaq0+mTjpbZXXZr2uQbw8D8YrDSJNxyXisTegue
YvKZRw6viCcu/iuLTicuGe/Zq9OOjmHwbsiR1jES20QJoA+vsyX+ZRfHJyjjfHICP8Trbiv3VkoS
AH6ITmKuWREQ+6b3pchNU9bkxFCID9PslfhZSUnkRtws5zxD9yZQr8aDIe0twJvpoYvivCd5vVMk
n6/7+QUVTj4B4xMoIhv2LZi0uoPSoeD/9VwXIV2UUyu7V7kWgZ6F67AqSObcmDpeSOVlV6RRUb2C
D+dm9KJ47wGVXqsuYW99nUa9RdiEyaWSlg0PGtcf8UkIrcSGVljC6VpA/9OYj1j0aYZC+3e727pa
R1HuaLa4BpeeVh3VUtqt4KLtfsL7gV5D/n7oL6Z514LiMXEslpPJbLuEu0pLwPk56jfh5Njz6gMD
yNDhpAtx41B84/kh5Oi529c2IhXPM6uDD1JIZrWIii9HC98bcN2Dq37PEd2Uu0kY/DTPSl7/F9jB
DLhnNK0XMTs5Ohc8aSPWc7Torj7mqta4fHHqnlK9tlyftGljYscSy4qOL3tuzEH2AoeoTTMn6jaY
8MC9mpiJCmaRz52sxO4VhggSmPBXnL2RgPX//qnCwQa5Mv64KIJC5jzLe+5RGhYkZ43+Tuz8LJEQ
gKar1XIW12n3f/wtRhnKDjHqI5jVP3eJckeapDnPMX4IzZpAWdDhxiGPVTDP5VqW0EksyDoT9lBX
C7UmHSkvKj9IdPTSGDvXAZBlJLW8fwB3+NUWwFkAX2vRRqsWrOSen6lXbNCYrr6SHM+Sk47136z0
PP6ea1UwnBoaH1Ojki6JLIX0GUHsxT+vcIpqAIuoezUgryGK6sW61hu7cWqN1PEiGDdsIru7xobv
zZsBw520KzSGtGPKjwDUNfuwL9htv3FB6wi0tGjuKyjqQTMKOcjR5nMXwutYB9/n9BX+xm+V1597
LIC6ehd4kJIBAzyg+kNYkcMpVHb0WaUHms97PLIn5qYNfZWbJnmb9+zm9pEFF/mVpOzXK71o49aq
FjJxnw/mE1o3jXkBMPRgWWf+5qxbA+GhTTKuxcvmh46DQkHq1q8fO4bDI4npRgYLFwkOQqsoLiUC
+atdkSUla/sosoTn/TAgpMNXqtbChjrKEzJEBGRG70s9GPsJHFfZPtXlSeuWPpyZh7iZN9VKuyDx
0ODMxLWW4q8z9qWIaptw0vCAOI5M4cse8j0Ki6Rt30hRxd3PGUoi3A7GOLmc2p97XpTuWQsjaExQ
9uSA9zyZ/dB6WoEQyotN0k/Lo9E8Ic3Rqj2sDuo0PYPk6a80NPd3L6cIsts7Xdezomd7c9YPawj6
7toKYwwtMfns3dMSAIkdmGa3Yo9YUv+SzcFZJIjxgr5k8VycJuC1C9vgCdNR5pADQpqosrFouDlR
AQjmacC+ZXmQS0HuqhLp4a9Zw+Wovzgv9wGNPaFRkg1/X7SQEeU3EBNzIsU1+IK/7aVjwIaH/j5g
qjzMtSE9abKRiIPLLeE4CUOZjCa3VgqMNzzHsYkaVqBBvbFUjk2HTasU4TaRx8aMt6WMKyTpsGqj
w3D1/9yqxgvhdijvfe2Jt4pTxhfRkgrkYYqbic0pVpm4Dgg+/D6F5MZXVfQ9ZK8lhSCHjC+pWFs1
YkYw1pRXRqNv0aAxHKl8ibwgcQlnEA9EVDHFsNSFPC+mJEd5yA0piIxQ2qrZuQ4115TcmdJuaEHC
dBDDIqNCsh+Xrl2DufKdaVOCxZUSe+3UNcJ49ws16t+AYySqzMf3xzLJaZB77UQOVAECCEqTcyCX
XP8sasjgmhWAFBk21N6N5e+RJOzF6GUnq2qs1A+m72AhE49vTR02bPZdEGZuuqxCRKrwV9yIfn+o
0Z+s/AzBn351IfzSroXq0Lejk0qCMYFLAOT8gPXxmNmd02KX1clJjaPPSiYg84kvJNTqGpS3kbPf
Y0kZD/9QBjoVqfYYdvqllnvxYohVGe/HwCYHw1d5Tp96nDNmPJFxYNCmyPYSyoOEEtvXKF5YpO38
s9MpwCThaXHf7aEzLt84DzHgRXnVQepd5d60NWkRQ57F5CfhnvF+E7q9fqJoAArjO38eRFzPVbJD
Tvr3yUBxr+n+DNfPw88Ki88ECU1Zv+JZv4qMoPhM5SvwADneDRvYjBGg0YMyrU9igeOLFmM9cyJN
9PL6g2IJYmlXdOsdS421Jw3qwva0LItCG52YCiCIggdibLw73TzCVvuWKVWxX8dI0VIwQL1VS3at
DRqcGKduKYap3i5AinK7OKKaOqvZsJ+TxIZgnwxAYIjO/PJPJfZoQ+mw0cXFiSGdxd0TA6PXZlad
AI7XiLafC6OEqDfsY/HJUid0VrFaci9Hn/M+B3EY6IEaqoYEac8qLphiQAp+JYb8yiiquDpkBYj0
XS8zlanhNnwaozkPvcsBha/fSu7ekmFGy4tpBVW1f4kY56KdEU8wHE8PQIbB5iGaqduVi1VZcZwy
s9Upli2JmCCpI+bmTLNlzqhx64U2nR+FVxuad55oW+cQlW1vtNBQqcvpa6qMbG4y9+qY2UUi1/4F
gIi5QSUBR+oNR9jOJp/hoCA1lUmPP4Gvl3kgtUVfpL6g5c/ZGdb+t5Ooe5dyOc5hAN9VD1pRj7++
y/hcQemVbHft0039tbO4nY4YMwz8pX1lqWoPga958w+zTTh/agL6kvBsQfTVu550MGKkCIuWY+6t
i6msInhJRIwGa5ZaREq2BrnlotGOB5b5uBv2cs7iCph2L69DangbYJnCoxrOVkYZbxFI8VCoFvaa
VPJxDq8HHkr+iSTqdF+YGFpVSAWvlOQjx4VTNvpqb/1oav+N/g9scQ/VweW6LaCs9nhXJ5blOvSc
dnz843awTuxQkvkYCJsK1bi5gaJ0Xv9iQfLrJpvOUefzh2jQD/g6AzkAgcFymR18lwLz/hMxiYqd
ZMSkBLQx6bXoJc8I3XPbGzwK5irBl1ZA7RPv8TNKf7rrLseS9rGfAdX0VNJWEUfDQTzfjB42H9Hi
vMXk7BdF64yPeVzV5tam7JqJ9tsf0+EOCOr8G2qpSVfrKgv35Vks4Ac/2LVsFrQzm9qDgqZbptZZ
BJJnAZi42vPUUnyDY2DWDaAoOsOoX5IJjXSbhQkEO5Ggwxmi1KMO2SwXWl0U1/w62dE8/ebg/C81
sVpMAPs4okKbyeJzjeUDIdt4XhgOD6MeziJ5jZhNK4NCrJh7acSrMGL+xtIwBqZR+5qoaCFla7AM
EBRlwumLe2WJlX60xb8bSt/LHxfgfFZoTsfEg4jZISwNC8QyvWo7pw6QDSxcL/mlDrWzP3NVMQiJ
sUmdk4a3qbcfuTzOmtaG8Qlk46rf2SkjfGiSZZfFUugS46iwvzX3rlqHOobzNBufRfXp5TNYB7FO
LxnmdO0wyN51aMoS2634/E0MKSDLaPKI7KB3PaUQqKa8Um1xhlrOgEBGWQO0kgZejnI9TC2pEDFC
8oswlCSS8czwGagcYwojSCVveDwDtuUqI1ByIJz1yMeQb2Pof7LWtofgbP183GVUfroq67K1lfgf
bE5oEc9p4zatLTkCx8U3T9RouMm660fI40FPWE45gOcgtdKgTNyv0xMg7gQOeTND8GgFGfzpemig
EggrJ9IcOF8Xal5hW6JkcuCQ7bCjvKkBXmQoj71q09PYyOjzqhoFtpq4CPVeT0A8840ATo/wa9ml
eXCQqkDthe0C4otGLLsQKeMeShOic1zUumAKjGpR4lD3cbXsBLkJnHFhecb3dnYZYa53HxPlgjiE
SGPqW+CLlCGjfOlheAdkONLJSWHUVklFllCbIp0XfFbT5W3ayA+OStM+nDuUVGxmZLjDQ7JHPAH6
8I4BLj3HKlDGEK8uYn0mjhUdQjROW3OGS/5RtjaUXVgFMBGBLNW58CuA/21PL5TnD4r/jN1I5eF/
IpE96BmHtpcJmfVLwKOwf2yJ4t+Bw3XF8NDYBWM7a2Wi6PBVsNWyRPMAjxqFDvjyQzuo1USdG2Cw
YklSfvW9PMugvaqmjdTEP5mmtByzcDUHXd2/bidzQllrIZ5HwRruJ8+G23hbsJm6Tb2v0A3bsbv0
gdtmJAQuu4bPZV/V4WmUVkWbb8lJjhuPivpWgsyoEqJWdu9Ba5t8l5qdSDxv+QPSWemWytW+jjE+
LiLKy2lCI91HUHE8cb3LcnO6L3gyowN33tqd1ZOJEH4PG62K7DN9W4ZGuPhDjoiySjjvEnZButN2
JC820OPDdaVBuvwzqvremquswTenDJdn8c/isUXnOwygWGZpxn5P6GGhKYPqx0O86Mz1tooZYf74
s3pxMfY1C05duMGHvG7EPajpDCh95vi7EZA2jm/CJYhdcCxb+4sNzKZw2O6KWHRLfwA4yXLW7Jv1
vIVZ423uf2wq6Y77/VmOOfANpilu+SHroUsqEIWhDnduKXHzF2NKr9H+3RJIbs+broOGtbnL4JxZ
7jEzHYKJQHReRE3WOiTCNXEW1qQ3GPB/xXlVMIPgKMVuro6lP31AB9eFpU2wpMYfiYpFhH9LFRre
BDfaqtjpdlk6NSSuS3Mw+fTpS9332k3wagZXj/3pgUZaKuOPFjiDAnF9qkk+SA9JonaodYYkEzka
a5RVPP3L1/Gv/k/wQuSP09LjzLtDJ2JXbnGvQwf7NRBUIeQVS/FeKrZgDjUxtqEDM29D6RnglKjP
iEzPaCxxNDFCNAq6JbFzSIbioAqxIXLAaJRKbjl4PJqJ1NMYnfjPFE43zX6W7Fcgpq/JS1Y6ZC2l
NhGXLGsKVWwNn6xgkz9wOBO5K99woRl9Y7P+ufPSzvAEP5j3qnpszSKiUnAUzcPv2SpWNLSMubek
dZkQssk+b15TM1/7h4M+wDa7kCJkOAdHIXSR4VvCdnNaQwISmwpFRuZBxC0eOQyJM8V70XXOyvSw
mjScP0QDzYaF5HjRbHWfzvYdanwL5fwxIrHdNLnOYdd/yQgFjo6lyf4uPuNvqRsSkHqn8aW8w3Q1
pUbpASN/I+k8bWxUNFLbCrSr5hkNahOjJa2EGYv5Nb6DQIpw61RpiRTgdZpBss+Pt2AG6q0BRyJR
FE36XkR2ZobMc8G8F9Z3/YKUWars6+BVRWlVYSX6avFGva3urs6FG1J54E6xfPSgdFh9BDYKLQ/z
a4XMvqMVVpuv+BL9uVo7bnbhv6cr3s3cguzOmsxF+q7ivyXD1Hw+jQjXKrwUWPfMzCHsikcT8QvV
C8FumwcXglVlXSTJAyYNNpmyfDpPA00LoHR7I9nbeJHKxI+3jiFtush+LTaSChmTIuvwRQ3WRGSp
f6WGcFWDj6x58TzH2y7UMj70Lger+vR87y+d9kGt9hvlawH+f3qC/KtlOTicErv885wwCVmoNWbJ
EJvubS/BfqNds2nUXFMTtUFTPF2WDEDuZH66vhHI75LqbNAM5d21F1X8nfqjmFHxVv13A36elnCU
2ueWAzThz4+bnNkJwwDZSUEuUseB5ZkGjE/HGWNgNTnw2qBLWDrT2Z4+qu1q4H5SbYnZjnhYscEl
HC9mBITgWGbSmA6gKt46QxXtTxvSTidxotr6lRe0H3ieWMBWuMIcYAH+mTSC0dMpoDXGfsREdF0Z
6yLQ3BnuPExdtP7wD+0W8PX5ULEoq3UHPHBGirYaWdQYqFDfxwZN+t9WlSS+iOvSZA2AY5+XIgap
5IYagSz/sfmU7nidkKIQNVtmhe3oQ4KWG5Yam3JOrSqbDmzfmTs69k7mnecyMWF392QdHq4RxmYW
rSCjuXvID0q6341KhiE4zYnnIvgllBEkvFZTre9Zndux1k5QNVncDX1npcy9f+eXRxyzf0n4gX9u
TZN1PRWR5vPU2a2GT79nQFmncBbAmIpPoyDdvWAXSQqua7r5oy7A9VJuy1idbNSdH/ldRO6zSdzv
p3D1kUbGv+cIOElZNWURF/WShBTJGjAUpP8QFXDAwb826QJTBm5aKMKUwICIhgYeRuNpUo0aKgKh
DTKAvn75bHpeH91tBLst0Ef98gxvZzhVtCSF130v3grl3dMpThPDt5nTDvNINccwPSunOgjxZrFr
uFqEqf85HYunTN6Q2jJ6tDOkzTXn/cvQE2t8VbNWfZel2gBCFRIefKKqK9Fz1VdSm+AgU8Ac7lDf
z3Y/AdhL/UwH6WKG7C9NlFiD9fLuDWpRVZiv45VmjIBKNWoV1Lw/HBLcAd/d1bkhBakeWJsKYR1R
mde1if4kKCBT7pKFqwnFRNCAq5qON3yJDxP0j5z20o65s/a3l/0WWX/qdK6eLbtFPm1UynzNwiHg
c5GD6JVhfTskIGg88yWohVKCKXiVJb7Ki0X2+HYmYTFbMLE7G0H9aP4ULB030O0ViciYh6rddHmA
+ObCo78nFd36KEg1iZtajozMP0WVASu0DESgWQd8jGZtm56r9UiIPDE4RKlv53wjjOwrRJY+LPvY
I6WFi5g+IT7PdX2OHwcDlb947DlKEQg1AGvzmvSKMZ5H4RwQYFFXWLjEyHTganGt9S3ISjlIlRgW
U3HOcQxiQMu12zORQe5t0gMOXsGisMoYke9D0B5YEMnp6uO4cqrxP/GrzBhgUgYlltcepGNTa/ov
/0L1YQwJoef7VucoDicku7SWfLDWPEwQQz+Tei94rexGB1EblorbQ7gdL8AnOdGuwh2WfkMlW4J+
BkSFIRveq9UTb1baRRSpRQCy4WAGE8s0qJP1uT6yjFhonB5FrlfG2R3X2ycRw3gMqRzetl7x1Gtc
eFnMu72IOyxtYmiSmOjaIRT8fdb/kKRYpeidUO9WVrr7szcv+cspaXlAMHAB80GJpwxkYlkp78Zf
0JowHnPB1fNZfoKwD6iJIg+ZuTmVWJEBotMHTfHLtbzaDuI33JEkgJRTwTXZzovD3XFeVryB6qc8
hxQ7m8aK3+lKvS0439qSZ2KfjJRJXteu5sXuN8cGGWdXyHnf/8CHlGmWu1lN7ifTTLzBEx7E+xi9
ugvtzEiWShLvHpRwAxoc3I5k3NDvzhd4cvUTVPJL1pNg1tIRlIh4aWXZs/QjJt9xTNPSy4RSRVNJ
7VAYeCLm0kr9R902qW+W7V4NLMnG3rn1pgr1DCGGTTvoYhgejXRTP0z5gDp6eDeM4oj/8srC1ozU
CIwo7+IF9xmpkMisJSRDVlYCBwYP77Rs0G9JQxBkve297DsU6LKdKV3U0/Ih8daV4kN2Ha/j1OgM
JFH9PHjiBERSUFgsd8uUdncv6Eif6A9wUiz9kUiznPURbm/ZXEJMxMPddbPFKL/EbOT/LqgIF4jt
GP1E7T3GdVH+MYQVjPgCbrJs8N3ERxMMF+eQ2moS4PoCdhEEnQV9m6ToNNxSuXPLjPOoaP86dhpO
PkFgh/wnP97u6eW3BfIEPz/mvUkJeDg1o+RSj7XjhcnhlnRTC+IIlo92o9ie05F7/tZPSqc8BbJt
xZX14Hi9x7asEbvrDdzRla72DujB6WOVE0Z3mkXKQ2oZ6q89IICycqgZ5E3e+fiXDQ7V1TVwJjM+
2No4u5FvZhRJEYu3TxEuMkMPiVQOIKqsVdKCEJ+gd9XWr7IqMaczpHrbskwSXnFmeCeAHidooe7+
nEW/lUlHtU67uLIKf2w9vFKSXxPdJfTUzwQTEDeyi+YF7t1hF/HjzwWaqe06Cw4z+0pGV4PNmpxK
euCe/g+1SEUCM+xPRSefN+JBJuJauhHf+kTNE3+th9JK4qZziiTglZQ+I30i2HnylNcpWfI4NCMs
8dXNYQ63IQ/itFCrq9SSm9Ydtnj4DkY0RvLb7DWMeT4v1bcLbRAXoCmHqxDixouQHZBaZLwBdE7M
zxuocWW4i633ULz3KtElT3FhJnhkOjQfb7tbGnM4kztetDk/zyzeqaWPAGoWkad8RXBLOP+ZEfAp
eBZyr6lC9BucdbyQmlAn0aPbVWAUhn0F+/ypfsEM/4vExLfGmyxesxnGUJtTprMHfMNILC1IdT54
NSke2rfaY4xsoYygEzYEsDyX6PuWdOgK2/mwz9DxBSsxqoju89CHF6EAPXrIXI/pFpeXA/uNI0Bq
mTWGqqr+Amfpy3Is6XSVkY5IwM9KzP3aWB0ZbkL6T7+wKe5Fuj82fY16i759AyX1lYhuqQlWtEmR
FTvtpMsv5Gir7SDv+sRqQ2UmWEkv6YN/eEZdO0RFWYOadVaVnJEa96govoyq2FZ5V4LLf46KRacL
gWucBoIqgMSxQYm6936g72VAol6JNM/qcLszr06FOaU5qXPUma74XF01hi2Xt+er9K5KgNKyCSbL
5TAcb7jZS5upTFNRPVfYMngWe0kMXCI3dnNOR1YV/0SgiGvIB79uULoNw89qkCXA7dbjkKe+Dp4/
y+5WqA+RJ9Xt61B6MYCpUhJK9SPlfof/xxJUYoH1NDao9nAI8eH7i0fG8fLT6dhDy7W8h9NkKyTg
mE7FGwSPGOAwMXzJbTW24MGzw/zrMLOh803XkLry0WeIAwi7NvKJTYgEG0ypsghW+GHiaAVeEH6k
mSlrU9mKd7UZOo2RTplc/6EHs9FattVOyA1agxxHgPyiwQ0BeBAZXDpASEaWIdKY/YxD9dPMaazq
o9srIvR5XFELgbvPvdx26BI8u+EE2vudbbIFOvr1suNYwBsW+ADwr3CLVCr28ZRsGkEgvinVemPe
9TNR5OwiZjXWm3pG8CUK/85/73SslkntLGskrovrWYCOTd5uOadmgq2/e4pcmjn1fs+wK/CUGcKu
4Pc5v7/MMMAusYSYuBEjyjcqP2MZuXcKeINJRr6uJc2hL3Tqqpmp/yWWHVEo1F5CeQ4j1F9DcZt4
vhSMMM1z9SCjgl9xdqEZ7afRutOC3wzycqIrgUdOS+tSGBqS/+wHDTR5TPvXi1QCWw+m/rdO2iXt
9snIwGB3p4htYojnyUQyMTk9uaYxHLeDxXTtVJ5575PifshjMRU6LDY3KsGxlR0Jp9ioUtgKRURa
GiHFBORK/hSwMfcVcLh524uCaKJAlahAmX6NSEyrjbPslyD2eFYRf2C3dJlQjEXZ3Cks6u6EGRhf
FZjof/Vo7IOrkcF+Vdc0Stu5Wt42fFo8vvFIzksr3M50dqfgZd5Yde+/6HLGZx0/M5iQZUxJloMr
3mpJyHvEoYX/0tmjXz7AOiSJzV0ysyVetedj8CpU9PUWgGRMQGPKj+QMHoZGF4YJDd13DCSdX6/I
c0CcYQ2Xvlj/CJ5tmeIWwExQihK5Ida/nRbZsraulNb6Lj7lqzhf2lL9ZH1LsCJpfh5FLL5j3QSN
qDKOWJ8jrd2RHaZV1LOVR8seEWF0dAqTogebttVQT/ZDodX9+HUY4O6udEnJ4flaB8zH+XalCtq7
/9JDhgdpvbCiBqVb+/ml+IgeakgnLBJ0cYPP9l8pOLH1SJytjT7rhX/JXmpoTBPnAFaeBBjbwbdC
blHyjumDb4kKADoHQ3JarWTszf8lYtymZpX194NAyLR6NdovuWNCmZtYNGcfk/S2quMxI//8g+E8
FL6I72JJoYXYvNFuWkZmYKLD/wHpNTT/feWZVqOoRG4c5MElncoFTrHN9Q1jWWYMOi0yi5cbCRwj
wx4KymtBTHlK2CTe2XkzUsZWxasOG+IRdA4OGg+R+G+N4KGv1AZI3mZXDCZdXZOapLHn9PWIX/vp
4KnQhffksYAyaPfdreFjeoybw1Pvq6fFVzkVtemOB3OvFHbIKY7Kf/tVajGEyozm/ZN1fUQ9FLTD
IX9R4bh8w80BVShv361yzKMgHkKg0CxeICd4EG1ZTdY6hDq2QgSbDhLsOZcFEgN8GCK9rtApb7wz
AYB3O1B48vHVzXrDuJcTnPV1qy/OKlBFuiHFpsoUlIDXmINWNzMltoEDcNyk+N5NCtme0FXjSYA0
rt10PXKwpgR60HP1yV5rzL1q3dw/3cBmsgoWPFaB7xhSVOR1sOOlSMdGZy31Qn4d5cwLIAZ2TEl6
UYMMrp0oolqCqinFTu911JUurT9hcRXOW+/Xxe2miJ59vhUP9fn4LRxd/2CUH7YCv+05DEU1z/7k
sapZ8shfI9IoOa6hfV9MedeDffdYFeoJZbLaX8TaukWywpA0hTty4MVZGn6E1wsRU0hlLnRLQ7cA
OJWgvV3y9b+rWIoFmUouVyZMvJgalNwYtmmkcuNCZQV8tQEZ0lBK6PmkMSeRRv0RhthOGN+u8BZT
m3k0DqWuZrdv9fJd2glZg6RGnASzywsLStHf0wPBFpUT8LCcGBImhVc9t39xZac3+39iJvdXsazD
QjP6BhHyynSxjvyyq+INPjeigG+FeGbbyn3JROZJMCmVXRvUvn10spHKQY3t8DaCgR7PvV89Uvpc
1ZrkBth7qSfkxmxdv1KZpJr4eVRoujbKOG/aY9VU6DDcnQfk7AWMEf6Fc9oH3DlDGnVYKR6oZN3U
Kg9JY7pWxmqkF/I2rX27BvDFDeW4c523SrtyROUkSs4d5RWZ1hRqHm+2N3EFR5dHu/OSJKog+0PD
nR103xIP3fyo9vRxqiIj9B9nT5+6Pw1GWb9ZcZos1IpDsFe2LYhIHnWbvCdNy5taW3d2q2+fuilW
eG9YQu2pZMxnGzJHbX48g7qd1fg28iOrfROo5n0PSpjhq4wm0HvrdL+02zpawAzBNNFR+WzsOM6A
5PfAQIiIfw2MfC4RLEInhbAzDg4qK11ryCW6AvxMuhXQL4e+ma7tjj3iXLEsrzPDg01dOWvKR2Xq
KCVbLD3rov7q8C3GDrz2bGN2dS/ZtXB/6LfgDx6Oo9kxNuBnriM5gbxP48gzx7nflJmnlo09YqCq
PkXaiB2EbSG1UGCHixThQ1sFaSFtEi51j+GC0ASQerq9MA/q071GbGw8INawemm3BRMaRgJqOteo
B2CdtGFrsplYhs2LTBlLTfk6YYIflI7QJAWJKWkOQBqgAwDOGnVB9gexgzi1T/uz1wXYMxXkVQmH
fF5a3m7Apgu6kGyFdesNc9E+JtNS5AmS8MlP0kmQhlPogjdpFYvfH4EwMqfnHmjgGALCmpBLdenk
iTtgKofoNmzn6NqAxfL75c8BkoOHr6a9yeh8LYIXwnxjJwQlI4erKwqC0iErUkZWzKQuvJLme2Ap
pjmDnRNILIYuYKE2JLaUAmcHIxZzlEaW7GnzjAEEmkXqlQNM0I2X6P9q8ZqdqpxhkyYjUY7Qwr1t
UZbG7t5sOEVy4KFhsXwCL0cKRWdM+XNKo+aYbjwk8UwVDpX8yrdAvt9q2jA2LidK34NiP1TxSwyg
qjCOGtluNXBqIkbzA27bf8EzRMEpgyAUxUTO7ytW2mItCIJYeDNnC0EjjMvzdprDPij9nGJYdWVY
BC1BZAWNsiy5x/lD2LnbrG3KrLRSi8qvNsCcuZRUn8H8fEVMqjiXr81BY1Chueu4VnZ44DMJVllX
DXFNcRyyBny74yiOY4+xIOiILOYCQ25LJqCgSoL5LYQGiP9aMZmtvfH5RymWkzGW9Z+pUNl+bAIT
RCrg4IiZpPgzazrE/j2fXfoCqTYMsfMzIThbyNTU7bg5j9k2v5M/3gsNjcVe1zRjai5qGtw9nNF5
d+20eehgDhkj2u3yQdsEPoUI3flnIEqdUdtWnhHFL6MV1NJdFvOxH2aApSH87RcpLzP5sqz5bTqm
BvE8HVdwR6XA1hW0KI6l7hDez4qAzy3ZikvmeOfOY/sqbh6WEX8M4vHvB+8yJbjz+5hGYdm1J2aH
qtpHQlT6+5f8dAHedNIo1vELlhIjVv2MxOsnoYdyYSZv4oJGYfVIDRYKEsnUzWUsOq+GHRMpRFYC
58yI1DY6Vpe/dm7CjhJZvmJKdMtZiqg/MU1x0vrnle3OChdYOlpFY5q0xD4WD2OURpXDGRTM9bQA
X2p/uWzY7kXUsxlO69n3OgEA0D/TwiYPXu47dpOdWDat7xikTGvhRFnlKsIbCB+RKXae7df+iQA2
7/0cnzhXsSRlgbPaFZV2vTrrJM0lUno5/LJTV0Cbqomd7xTDjJj2Kkalp3/OQTiUIJHsUJOkqcoh
6vgjBoqJL1dWP5ktOHjQDj1O0UQd/gfWzsUeKLQxMIb4u5RQf/ngrwDNB2IGJrk+qvV2BvkZjJ7J
QKB/iPTJpJzC8J2lWmTayVIabEbxJTpW95AatoBzE91aZGslB0OkDe1CqwisQrjGqnUAgsEl7xBe
/nCseTztj4VK8GpEeDDNki9BN2GUiSPqSJFYzRoOQwvp5Aw59CgcxpSyKAcbqcStgflMSwVmMAOM
n8WIJUa23oUE8Xp8Q0OFp+J4ai71fthu+CRYXuBfojhsvJxAZM6Y6n06NYmGfnHKh04GvxqsM7uR
Fh4jKSJYt4PetlmgAEpwDmaEYHka3dF0Y7xYEsbwJRuD7ysummofLoTGXJTHqL3oAllgMZeKDKbb
+IFxK9YlNuIXS8y/bQ6feXeRdZw6f0cCHA8b4Wpt3WWUMovSGeGZf4yLSHGkda6Yjf1Vy43Do+LO
ao/d9yQCVyKnYROys8XISFd5p4dF8+bZn18aDFMweTJ+I/EwKKeZdaudVU2dbiDMkK5FaeMooQYP
1bkX1kV8RV31ybKsfeHni0X7MowWguRoK9ritaFnNDTK+UxdG14JY5/FbtSy5RhYZNkbeNs5Nl8I
+0qSchWhALGbh5uspMiv3jOm7JzuYD4dEziDCCn5/14SMFj6jF7K704ivyk0zMFpyX011Jdhvsgv
iN9sy6kLmx3XJe5pCobcZ1ysIy0nq2CQ1p+jUfPr1NQ3rMNjDyw9+hyOiCpWsDB1ClJdJ/VZsVuJ
k6/ionhJTCWxLZPiqA8a+Rpftn1cJmQs17ldeNoD6jv9uS/Pem4x0G6cxS06pL8Lo5aeajI66sfA
TmJPtIME6aRA6Pl05MuVTKfCOdDsjY/UGp8oev5L/KFTISV6Cu8KyiRv61rScD5fpoIzYaXDOhe/
1nB7tbAfqwgi/S0uHdVfFpwsR7ULzjFPGCMhxE+ZSw+phlNb8QTaUV/lKXaMlC7AMT0b6LkXVLYb
nBh3w2LA43fwMPnozg65Vd5ytAaMtcjCp//AuCaQgANM7P9uCG2bmaxE8+6akK4QsvJwqbMSQTQI
P742jU7qQjo3Q2CHfZ3PluVxxQimBz+kqXLWZ26rTCGF8QJxfKBxqyoNX97ycLjyHB6k3LbaBR8d
rQdojnqpj4wh4d01b8Nyx7Om0WWTHXLKwV/x8mMjVwvGEoY4+5q7GoWJ7ijIcOakv2Nggfepd+33
+UC21CGXUJfVDVcwfSXgR27ZAoR/n/cahhJMG156LRmZptW5wvJHz6tXjzATYPvvE7FPoajPQFXS
NDpPzro/uOTmtSU5DYQ0r+O62fYI9TLW7nbj6kGRKrWLIrsN2novEK1zw1kfuneoR07Kw72QD5zv
UE1UZYzIco0wZJv1pQxCrEIdtkDw7vbRYaiSmODgGEGXOFl2Z9bHzPpLPYTcfA6tPs24BgxZUp8C
2q3zJnjxTgDNAWH177E2wltcjGXjzAfimR8JaxwBJiujqjli5NJ+5qyqGUeo1BRwnK0FzLsMBMjq
OkpInhogMRc8Q5kOeWdHko5Yke6tx6BxDGbpy+rHzlt7/X4Fuv7XwYqSnI9v499ASBwLWC3ys2RO
WZhauYqMBIAuOeWwIu1pwey4DaEvkjOWESES3bTBx9Qr/zZwryRZKVG/bww3xVOX4NmPX4sD1jaa
5HOqUQ52IRmjIcfn/tj6mD5zvIFSZPlkP/mNN7mB0fGQkuTedRVAhZVKYByBuHjV0pkrEQNlIzof
mMjx7vMiTvBqEdTEe7T8XzWzLkIKsEdaD1RboLU2og25lDqF0jBEN6EQyzoxGvRuHznWriKJiuIC
b5V6GINrvNeZGUJPbTaowK0u3HjCKEtLPuMKR/ATSg2WIvrBbnBkQLI0Jbhru2UR7IdtqmaYk8ft
gztOplVgNBbNsC4KSU7CyDxxjR81n1dYldPmGXN6KpYYAVOlXQpkleml29638LbqvsOkiZDJZzMA
LWJ/mqokjWlLQx4WXY4P4vmQnCBNg36gIdb6t/F+ktCEN5w76RB9zlJz+fLkm6UoX2hJND4VceeQ
W3zfkCH1Y6zTjm4y77iFJJszlONr4TbH8k7iO/SBa9z6lsD2Hi+yMGzYzgNAhi40d1TtRpHbLOtI
aTjTKKfml9Lba7WJcJijZkQ2QE+kK+8kWMImBot8p1+9gQnUWJo6tOeyWfkQ1KsxzyqKYHuEKrl/
HkFtaH58jG9I5jJ2gizm/aJl4X8tSpPKRjd5sBxleIdRnweagb5l8/np6DlruGOzce6N6HZar738
8l5u+p12K8ny9PaqYaUAWvyDY3XbmCeK8pQ9cjeZZ/GTKmSMtUtDyibZrAaW5b0p3JsOSuFr7gqx
r5Us6G1PPIeBjdXeidoGda+RcYa3Eegz4EBVi34t29ww4PfOqP5Ts5GvNn1LPOgBjJUOxWciJ4DI
hO2PHjtfx4/kIb7IpaOscJ37fqbH1c1sPujVY2oZBRDABpidVsJx3VgYF4jCf96Umh9v8yYBawnf
Tz1npvAq4Tuu3S78zd1x9HZTI58ctJzCuKdj51hUxjJcT9Nq8x6Z8aQctuS1hffDKSx+BwBpVRic
OMuE2pxuUcGHqdnmXGmvMS3N0xGV39fWgIne49hudA/pR4hS9JXUEVnpm32uZcOGHiyX67gx1TsD
NdBWVKyu75/PoKYGP1/nlUp3s5//jfSf9BgK/59g8XGcsX3nu9qlgcjF35CrCoxVQ3cdh2D0Wd1Q
kRw5Td1kRq0EYbRnRI1lLqIz5HdmDdiHY9juqmvpB4c8C6/awsKmRmu6z8RUP48UrGihq1Ge5laO
OkYiuhV/yRpxFxOAger6YJqRhHVe8ZVIRP7UO65ruGXhxCEjyyIJqdOYyUnJv4nFIi6f4jHKZtEj
nEXUkNiCKJfWWoPg2hEA429bpSVfP+Y8Jc6a/HtNAX1slvJmOf5bsbWsEqoa0wMTZ+wjJxlaqStM
xboNQkKER8r8NYZDFKQAsIMW4CLhiK+MbiPet48Slw2mJwDEXfQEJUt2Lqc0OdVSX4f42sG6hCGs
qehMNw1E8FjuVi1I/Isg+YjdsRhUR4O94FI7DuWORE5IJkYkfLLhnwaBICSZ16v59KskSiMJ8SRW
ltIGQTNZ0m9a7uzqOjJcYEVLqs/q9NKCFlx6fBDHBDWTr7NmsRvf/Zb7+HIhTR3HX3dWViyaVE5B
YUajlufVES6HrcXA2ESsUDuNwjUS6uVpozy68qWpJxvdjv0Q4I/wRK6hu989CSHbaoAUr5CK3JHM
FnjuqgzkFbPVaKJYBBoG5gK2KHBLDe8M47FWuX3Vr3Wrm8LQ+1r4xp6ZGWOoYESYStoPqDDI1Jsc
1447LIeWzu4cfheyEvl/hBHKBIIqpNMRp8jPKGl/SFr4Heh7TQbJyVzlLxttZ4bgucvgxRj8EA3w
6OAPfQSfQCyuDX+CHFx1MPgmAzutKiiLEFZbNXrbYknOuoB+Sld1MotMx1O5XYA1v6PISeyVLgeS
9dZxLVaQo4MaQHhWZr2EGY6EE8zGPSUvG35c5RC+WhgO7NuqTgOX4Fik67TNSkRVusCA6Cq1LHiu
lNbGJ+SZWLx4pUEnoS1kJD4aWTxOryB6r8hWyJLFK3+Pg/4St6kXh5TEZ1SwLWPMORSeO9Z64Tre
p7+iZ9qOTZafZRN51D8Kv3dPO37nXsjvFRDdSPwL75I9YzRAwudbozp9/o0P2InBALhszNaahfi2
3vfm2ZRJVoSWF/KKVFZE8TmmvFziMpgawG35S7hyEbpaxGayDpmncBbpUOXst4z5PEChhlsPKVDk
4D3no1g95OpIe1jCMliG5RtuBrU57sz6ktjGKKvhC+HlNGfwOjtIoUaHe2fsBfXINq4ciMapGwnO
eaVcK6siN7VWt3L2K8SdeAiFPppmA8pm4QJ0JHX+exFcjdy8lHqE8gbyML93e9qhwQ8EsTTmdOol
2tUQoWToeHVBBTXsil5ZygPnde14OoAoI0QPOyx3PjZlCyvbBpEScJKuovyXMnWoOCrKrvVPEwJz
an/k25yCqsFIE3KOItErjHK4cgL86kQ333mGXuKRu7f+wLogZM9hfmocrnofk38iaEP+jCifHeth
3LtU8qR5EwiqT9+EAy7TBlPVCMJpGznHZFl5ZTGrH1P9MXEAbG9oJosevmnFq26RobZwDDkcnLYu
RH7mRteNJCCnAoLRamF+Ga4HedB3zpeIWSiwHPztoWe2Mk3n08TRd5Db4JdGwaRvhtNtmnFvjLdf
DxoZzKeiJW9XXnV9S7KGAQGEBtylxjlAXTolRoT8DlCWfB7xdgTdOnHfjUS5bV6cfGrcRQVroOHT
2rQZF1lowPUpXzMMYJcn6MkL+94fw9j0CYHAdapPqC2QgBAYwIMEPy8rDlOtq2QHjLXi7JD34KwM
R4J4cQb1tHOoHGA82GFlGyFy6M6ZmVzF95e0qTTNWZBcXNor2jXEQeSQCyXe5nasMNRiANhIkhvQ
kYB180a0l1flIuYONSYTgOkLECLg4tAfiniy+2A+jPxe6JxAgkHPiwg10IFFomQ+O/wc3ZmixP6T
9v8IWT9zCXSMbhAECKR5rZ4eUiqiEBB2S5mxtSoz+QsKr9fV/3iQ+wHpQ6VNMUlOTaSA1vZcCYi0
MtDVDRJyiqIW7pyuj3r4GWUAspmOldfMBw6S9pTq9+u7mxqSFl96GglvySmUUwA2Jg6SvUyf9UwP
m+Ws/mUuoqjuX9m8r0nkTcHLSvg1r907vFIgPs2FaMVGd4jNGVWKGDlFbE4ArEY7SiuVKnha9IUN
I31bYi8QRDIa7X0eQHZUDf/CUemlxXKPaB11AjlEzgwaKWdS49Tkm8hduRiOrPhzZXBvPfEGcbk1
b4wqMHoqJXIWOmJNv0QhgaYVCEL9nyiQrC66cLfTjtOHyiSCiJ/mJoLo7/p5dNzGk79K/sAVMioH
AczY/mhDODzyF2RfKIboI3eGhx2Mo4z1Ij3ujr3bk3qB+uyy8jUoZzd99RxqZnmHg3u1ZcHfxpKW
TyXIva9aRcDltT6jl6Nme97n0TbQATNVYTJJyl9FKp8FqZ1NHpAXB4iW5tZkiKE6r0aCSVgHK1fX
CKOTSbPkVYCyoNLWyB2No1XQVgyT+JVoUOc+my44C96dogT7Lsq92NhIIpV8akpE9dWuAz8WRXyX
3aTe8M6+FOlDsrutrwa2T9hiOqt5zjJ5cy+1yPx54Hzg3I8HK/d26Ift9GncKWaI2HriCX8HLGmp
CWqp5Z5DOoQcEljXT7HFPVCgMiDy16ZXQhCk7X7IzrMY9wAft0UDbxLfSZ+LFUR6uKx6xsM+EqoV
c4zHuA+E6DKA0h9xpMlJhJV3y5zb0MCW1XEQPcJ2K5OTUjqnqSOzChzaIKx9WTAV3uXZqwjN9+8F
0KNb6LDQn0BOmLG2m6eXFCIraBRX7G31ZPE9wybm8eqQqC5Rvo33GpLQnRReMNkhOk9X2WbdwMiH
EAPC2kwgev+GL0DSkcTXD6cH2NHwHydghdcEh2+wRsqf3IME1q+g3LNBV+DsKi688LsMd8jGU00G
cAW2AJw+LAKUqOy0kAar6ldcgCDvg+42uTKezXwagbSC+Fm9XoqnVQf91MU4jjJpVguwod3MVorp
lHSJxSnLWn445UlTON+cBqk0THRjOiAf4jVmI+tvsWo0ZVyIr4e/remwC0ZTUrbqvmrDdJ/HTBUY
n/twI7Od978sZGIqtupt39dqGm3P1PihMQYpSPJf1USxjYu112ok1KiAPRBSSkt7CGMmooAJZr6L
bEgxZFYRT88aP4uyRgNmhdh91LyHXzA2zCi8UsRH4JdbWRCdvQpti1fHO4Ef4YNOF7eAPDZXd54j
L3CQprqGLwR31j1f5QHt9hXcBtzdKvrdZOyNbpG0pHHyXtLLk4CG5dy9CGEk7YmeTM6TzGuEOV4K
omlA5EIoswolOpKgC03XbsYK2KhGR5/A9QbKrxqYHkOUiUmI9OoFjPmOQKhyRxMSKDgF9Q86H//p
wqY+gPrwU1Q31WHhaQW90TnC1egBTji15//SzQU4E5pgjuyb7+rorYQQy8NHj31dPosM6FYv/oDQ
7Bj2x7NNqTT+F5fti1g3ChCwGqjkQkZ4kAOOKQGIuBNG1pFjKcWZClr96I1RpQyJBs2BvB8l1KXz
UNgiDwciDw7MEG3rXxCcUm1prtI/I3vrU8JCnx6UwWnvsawBCsVRBhy4ubonA5T7RydE9rTTCwEt
w6mWRGe1j3YqNp9gmekJD0BR0Nqqhkc/0M50pf+8Ku+xhPtpIPkObcjfqfolSZ1SJ1lmIEf8KWw5
gRY+3BsxQVppnHWTAT2o7NKUgK1JD+2I3SlIOJL6wL9MLw7jShg0ImBkZPBr51T0cThM3FvIbfF1
QU2B0WTbLVBrnVqTfN0x06AOUU49unnDbKfXZ+owKFV7bf6zBLfGU+gTtAtlTu8tb2vjSOCJnMC6
4B+HCh2VAG4EGQL3I0fZAJJpvqsKCsREfy/xW+i9WCRB5HzlxFBKKbeD0THBY2h3+cAk0+YP8sRo
dvtuxgLxmTh+U3HrXsozOuy64d6nqJkGuPhme9QteK0MZdG6BH1Cv9qVL+fcJrD4fg/RXaW3bWhJ
zJHSgkaNLtZ89tpT2xre0q/GF2BSJOxuFVeEOQkjm9uRmp7BUVNjGb9Va2gjT7TiJJgzfBEnGoEB
k0GdB2fHigLWC5XUYNp5uoPr07uMk53Fb7uDWNfrYq8S8PBu1Bva/IBQ9zsybIPMpLgHQP+Ctvpl
ebTLmhaapDCU6ZF1+zL2BMosyurgv0C91PVuq36I7tCp8kmNFulGIxydwduSFriou+yNWc1d8OGy
cGAHGqhVV87emirTfuPdIjUxyyvlGsXxlRkLx28i/XllQrH//MThiopJYgLG2HeXYgby8xZztN1e
U8hAOAu4KVBScbg7LQ4KzdImY40/Aj99idFux6sFe3krSFn8Tym1CpMoZQR4g91hp/k4QARVWCps
Z6SiUe5j3DxYTt4J7gYUmDs3z4lD3GZAYppDZTXzggOPri4CuLv9BPnHd56ZdR20sIOOidq54Kkq
qEZ7Q8fIg8GjS9xW5mdoixvJ2BKTraSBNoWAhLAnxQ5PVlku6O0t9ZIRGJ0wbDrpJ3cC7K15dldr
WjQEB9thQQzF7P/OPEk/o0+MKeAWSr5etz7GM0ruxiIOl6RQOEXXJebY+oWUl8A1cogB11JWm0Md
HvwcTiV6fHXrlse/Rs3P9v9w0LNuiExkGUMKvDIinNYOEWBxaCb54itanQfu/FIyYsVs5yUQxTTO
2qnlI4v8QsphndS4NC9F4dRJDnfiwsP2XKbRNPVol6gRVN5d8w7i+qxXEN5BqAGFANACOm9LJoO+
/hg/JERiP8bjxuhb66lYTB3Z/D2WNnthIKSgBU9dDtHe6nNhmQPPTO/32Rcx78TXvcs6tO5MpLLM
eBQ/qMq2Vzg1wNS+CmK1gLKX/U/BS/1CDSCaHdLEWfFdVPsp6E/FXxw/CGTNuTz5d7jzUsm6ddtL
BNMELc/JyUSi7g71OUu2FRKWGytJl8KtIgS25nn+p1Bjk+ZY+V0ajLwtVfA5eWSAYR+ssVlDyvH1
Blcbgj77GeeNvg7PQZ7enzFU3nAwjdDVNv9AJzcKV9WorD6payUjMsjqWpH+ra/ToT+4LM0S2vTi
WTNsStMMhrsIf6qDlHXZBefBxZM6XzYnc9/m2SLRkmGnO/zGkW3MqHWkC57+2CAq8JQe1pjpwymA
LlvEKku1IUNuI8bOfm/B5Io7L2LuFHcw+MaQbn34nTgSIcZu4dbz72xNHm2jZ3z8xGhHPceDhZ2d
VfklvlV0pMp7llh935ahs1gc7zcJSQ+2dsRTmLedGsyV8+EAfOY3a85OZfy2pLvb4QFMOiMbXg5M
1JjNcBoo0yYRE/h/awu6lBLX0PaizaWL7nV169z9olxLhmCQVL4LrCnVxIUoJfz7JHTh+kn+gQFw
ahEBu0wRhCRawXzs0Y1rVS+u31GW/FSYMtVo+YMgNETmD+KjjyApmR8gHTG/tzunXYUSJ/PexlGu
nL8Z1Y9iQ3rM3ROPgbxieuxaJ0FCFpZMPCbGiDnMZgChZSQQh5CXROssbMyYfUkrvwKHpfisvDsN
fWG4hG6WIWrVb+miAuVxHcsx8BPxh8vVAa+O0AHy3JpfcQIBcjPJCt9Y+mpRK2V2Js1JFlrp89QP
v0KinDOYyr27O5Jmr7qwJpp/tncydWpOKdZMo9FDdXFlczPd7C8DW7Et2gkhQpncsO6PrilkrX7G
MPsiuQiCv+YRAIYymefnEEImvv4SJMlAdjMJ/Ao3qgKYzNDaYr+SjX1oqo4JNKuTbM7C33G3khxS
q1axrGguAIExd5Ep4HdBBuWElJVRVTXcOHOiPxyGVNHAnCI4M4toY2gGhvX/O9WclOjhxLHBaNOc
4mbXDzBVJc7Iq86xhBrYr0/9B2JB2scqdYHvumZ0PyguL1V80bep3nzUAYDDOTqBZpt902KmZ6GK
xMOsR+OwyRaLgxFXLs5LqkhIV0yZE5/VxB4iCSgSXqAw8y0MeWA5FbkZrzfFwKfBJmkUVObaW3lO
GG+lLg8UW7kIuoEYWNkwEZLTw/3zWFta/Gl3WU61ITKjYblHbXmxlZ5mQ4LrYjpfTt7v9nY/Sr1f
MhjFLsh6CV8t3MdnIRvQ4eT+KX0JPRn1ty4XyM8Kjub6Ke/f0XDMnKk60p1sOfSgUtrRCO55pmY+
dImfcOsQnQ92W6bv6AEsL+IpTCz55sF++kGArhnm62XVagkFHmLphY3nzmKBcmQ33ORs35qS/biU
SRiKzWcYB6YsDo/JijTv+bm+JfMaoFBlCySUibKZcHLxgmPLVg9ThXJTHsg99t9jjYTmUSx7f6p4
rNcZO7g5efd3F/3F7U0bbH6tBdK5Zsz+pFg8EBcqNgFY2+MiaCWQPdXqfb3Gimsfc3OiqY+o7biX
eCtjC57Qdmwv7IAInsFORj4hFQcaYV3ZfBBVTgd2OIBHxPpBFd0ezESaUcKGvKhvOJMlogMLO49S
sNmJ9JpfcQCutsM7/91SONED8BuztHop/vfOvEMAjxV1e2WlIsF6N4MN7zNQFo/GQn6gSiEZGSnF
5ho2bzs3TSrNkSOLfHK4ohU284BMJmaf2be3dzOkVPPTGMnz8yTjWzXGXciGx3K31o6LIAe9qF5W
UVH6JP5oo627VNti3+IuFC0tPcbCczI387wc1nTUJ6lqUkr9y3y0t9L7wDYl9O48qWR6uraSqwwb
AhyH8NefWRY6tgbWoFTMSQM1xY73VTdgUhdDw0WlxA/u0FhUCSrp8bd9dqcSve5954TIGPO4x+ku
PZYOAPyhQpc21jd3b7QMd92/n6STN/+PmszJvoFguVKqhOd+yWRHaNntm6hBI0P5ABTaQZge4MOE
9qdHnfY8/0dSp1Bq/HzsTYmRLsrkkv8x72Q90LaN3dXTpqlLt+lhQUwa4I72Kt2BOLAXgG9R/8xa
BoV+eWsc2gVexL9fratN9B96fCdijILuMHdrZShSTSZQIcND3jktXo/7DyMQjxBgVOoOJ4F6Gi4j
NatLfnDtOcMomOMLUdSCZniFmjXBd4W3a0oaTgv6sXxbePaiTwMmVzX0MzRVUFoJhOIDZfDS+r/a
iHvknxLJVRASWQ+g/z5Ad7FkFxI3eTUbUChYvkJrLXmabbIU+vrghkhafrvd71qi1ps/5sNHhIyw
Qq5Tm9myVugUQFYjZE08yEgkKEtFumWt7W5DABTjuQPqXxpq6Uab50AxQkLK4RYFJMsIjzSPjJ5K
1/ejGhJ+eKw2oufTLXyXUSITEfwAVG1fVWDPqsH41Z4y0+AHmihL1p64fuCFwVIvuH7n4PhR2pSs
x4hcGdIstIax74wVilkLIvqu48B6s7p9Z+0FB+RR/57YYMzFOlHIn/x7/9CHfGKtY+k81N84NBG7
saABjZndS9ILZH0Fbzz+HoZXSIjEG8+ZrkHLtIJEmFKkW0tiyhqfCV0I8mCyGxCvisfUvvjIT8DD
290RKe31cbC0ytcP/n6bLgQmYiTNseJv0XE2JcKENt6xnhtjAbZyvgtMC3+c8iMHugMJIGFNtR/V
sCdgj128ebOHVjQ+H7yCnjyqERYz38rVOYvxKtoPeCcXn7K/japJTE2CtvdK1QSN4xei1CR8JBAS
X0AJ83IMP/gjxdRwSJZCzFtFfOyAihc+rRio+tR+DtteiT+qWHnGBEzr7LAaMTt+4wvFa2TTFO/w
osEAq4krFyPAFpGdllbjpOtLfm7yoqs3anNrh52cJkNrtWxiQvH+7Xh9nplNIwIKXPFi4ltaSbPn
SEGuLL8Ja+E/fBVR469J7yg4uHr/lUBmXAegJFO4/64fAHd7VMOqJueKBhrzo2wDoiS83h3MULTr
CCIbeXei69xeh294VM8TptJCIhM9gBvEjS6uncbZj1a0Ql5b8EhrHDBcn+mWknu3J+eaf3Admmok
oB7bQK3elcZtRFW7V66/7NJO0T45WtZj8r4T+ToYHnxNZGr8cLdyRi45xSfg9BPumtfhwLlfA1Hb
Cgzfr2YnCYu5klrK8h87ajDMrGONQD40Y+N8zNEjucVEDSS/FEP2vjYTTf5ulyxbSenskhn03rCs
YTlvN5pFcrbMl0PD0BMPjK5tAuwt6XMBDRvGuexWEATOXlL6Bd9+bvIA92RZmW5n7SNbNZW7VGLm
1qTjSGkRIVY0PpPJc9PLiAQAzvBMXZI9qqvalpbn6bhIGUCSJP8vnoYmYw3vIYnwTMnf/l5B3MUq
4Xy8XWaTnGAArrp1KbvlL/svdXmxJoquOjrF79p6UaaTju03bf97RBBiCiUEBUZRTdo3K4sj/ccb
PQaQqO60T7QiZqJI5zYBYSR5i4mhNegBRXXr6CLSYPejQW/ckJv05pUEKzCJKOig8bkIArm4cO1w
FL7CsrBZip+jj1Ei9lsg0wimXUOcTu22az72YVa9PCx8D5aiL8HO21OWpsDon0CpvbpcK0cSGnhG
lgcQHYTDN6EA2F4Tm8NtxB9TiWD35E17tyvJ71GFpCxo84XmjIKnzKOHvEjW4IE1vB5hiXVirXkZ
8aaWddJ9nC/oopY49eV+BAG0krCFwOL01KYV8XhAhiJvbIAvuV/LpVgflnphHV8ACWf3DKxlubqP
k8twpyzhJ5ooYtVPubfd1ElHgXcHixCXrFxdq/jE6TtaTcAoQWZhd/SWVfuadCy5V61Sve85p8jn
dg/QMpBQ0OMwb4fTynmYvxBtpLKXim+/s4WGCYmL2FbZ8EMksVGSVotC5zjsm3QhqwTt06vpVa/h
W97GdlbY02cPsuI5aJTNA9uXh8vqmyaaSCy0OQN/Sc5kd5xP37aVJlp4eC44o3ujle77KjFmt/CK
0gSOvY05DakKey7NJMu1hUv0OpssRNun+uFPW+9+Ws9+reO58flnFbNeQHB3dCEZXMClbDPQqAUd
v3pgG0eNI94jxfjzzcmECECBIcxk2WgKsB3yhH1FwKOZ+GsIjYIs1efKDV2KnB3EqS8Op9Un9iXy
EBStFjKhloqbcgGTN4ohwfkhqIn0FgRhBqNVfppq3Iyo6EsK9SQWoVdDadIGR9hggtj7N8nWJXH8
aw8PUPWK+YQnJjuHXuaGduEmzhTmz3iVFJ/c+DehbsejJ8xLjrPptTyGtdewHFzlSI1FwLM7/G35
2Y0Pxo+gP0GRqsFZYUGZni+zP/21CZ6hJmXRL0G7tov76NOhBjC26F5NlEfBccfrsUWqYRStndvp
nZO2iLx44agNg+osHbvzl8RUPc07QIg1kAchywFWPtgkQzzOH41bL82nUvCDQ3RCircdN4ZRi9G+
n0qOWpeuBbkbO5tAcNehJ8hsFKuy3/uxeefs8AZhVDtbYFi92igRCtqcxhujZ9pj3fXpWwTK/Hf5
P003hayYLEwpuw+BcMe8JNqfpLyj3ovJAEuLrcAgHs2RK2cYFulI/gZgBPuFSw5/r20jRo4TQRW4
rgTF3GP3SljHAeo45DLYb470fQpWKAHRwyvwJaQwDm9ZYFWtBPle0SuPRSJmHvENW2lLjlOQcXRp
FAY3glQSHMZtxjMbxCOVGHyDA3XyOgfpjDmDVEhbW01aJA1Jl3VwRigeOX9m8rcUbf/B0fwkEd5U
+a30eDcmQLNBP6JgkpR+Sd8ElNrd+0AxOmxvJ27BlQ9uUCxHAZGnfPcDBlH2x8e/edYTzXEqLi9X
JszHeu5dNOcsny4DUhSN6mXXANxxunGQlOSG0rOpgH/1CYZ8I8zUIj1ZIC2HxSgruk5s410aDtiS
a8aLmbWJxsivo2Nuob601nJlO5aHRsi9J5nC5obYeo4CtcGdFr0sqbAhCsb9+kkeZR8Xgko1zjtV
QZv6p+5BOvfUxtKHifU6S0bxaMWPPVnRXShGkEzkl/ZQ4BNyPOFHPy2igObVlX1SHVBavoOq8V0i
GBo6muT83OALbPigHUGYOnbmM/gi9EbEGppsioiaHrboP9COo0rquHXUTH3n0GD2Y4JyVKxXZpk9
Kl5p3JqQfxxWjsFo0FQ5B4qMU6bUoaszihCIIQtVcjXqdhHP/0cw5190TIb/zHpr59Q0LbyXSwSd
XKcDaZ5RQL0amRHhPciTNnFUjd11hNGlExHbbhVfThZ9BksVVNWM/+KgWjkUNGyNm4pdQAX7K2a6
0gj9oqVOWdGaiDDyGHtI1Ytj3x3Uz2vZPKBgQql5JIkF0iK6o/wxciox/QPRQ2vM6QcAWetcdSIw
zmOwzReLmZrCrC3rHO8F/b+cHd+sg9uEINf9821Ox5Tn4J9TNV7KXgl3U/JjEflR1H+kC5reMuBr
F3Ndy+tTj8mMWVv4bX7AvR5M004wgGby34fZoCo28a2bf8gIl2xLHmg+1sADXPkn+tsjB0J5slXy
QmYsp0kO5isn6Jy/maSmTCCZ6fspFlgZ0CkB5GCmS0C2q1rWTzfyasIP+oWMnAt3qEcCt6TcYgVT
HmCZbcu11dB7eVZxB3r5EJhUsrEkX++Cpo4NYMfK0avb0zsnMMGv854akhuMQxEqSfBlsECTNvve
NYhv83HLrIEupz5NeAad50SAevgUWvAA9kT6tYMeIlRYqT95vMOT9kHOs1DmUtcfeNmp4jabELXE
8pabCryw1//Bh79ntW+EY4PyK6LC21OyNeJ3hQiYcIgAh9i/RiJyYgReYf3raAdZicvXcfaMSk44
PvC2nXpX97GOKj/K/fNBWQAygUHAH5CvV4u9pBPW6OnJYFPxypDej+g+yAc+v0Kno+siaw1Cr3ya
OGeUf8vwn8AFvJ5k++LMydcLZ9+qqd9I6uz2Bn2yOSsl/Y+2ZRzlARb97YSJaqTnvRxg7PU7dVO4
VtzS1hSdQNJQN62KU1g667TrLo2LfleVybmXHEhZbR4dWx7j4hk+UsLhDfF6SyXYlJhwT+QE6XL6
hNv61yHcU7LIdGg17cZxnDbI+j1FukxOYhuCNo38nCDxv2wRsauHDZqDg4u7xoz9jV5BU+GAforz
Ee/wFBX1ewEVKiFHJot7SPVa9kc1AZDTIsZo0xOVkExenwwFNZigTc0Gnf98mpzlnOICcOislxgZ
+pdmuO86bTKuskmA8YbyO5hczWvcZRIENymG3Q3Pez6aAPeqBAT8SRqjwqSttkDsRdKE4XvKSEGe
aiEsFSrjhALi6jQl7kWSChb7eBAJ524b9YSYjVYHAvpVscXyBwZ+vJQHPhFZfNcFo2NaPyfJTzKr
H/ysPCbLByeUmk+0qvtoj0+enIpkJKymPnVR86uzmp+FA8c4AbTDlLPzaQG14FCho+ByYPnR2rYb
z4XWnqZTt4sXMSr022lmwGgIDVmG5OJfwPC54TQPiTYrfbHkWOVwJn47uGwLKFRX/8gYd/WHvCSP
BwIG2dZYQc3QuFbatd4wS7Ohsdk2apByYl6AriMxvkskx3tMkX+HlU2eDaRVgdrofH0q6XKItYQX
/SOcEsekwu6RlMP3awMQPaX2CuZqv2Q15xw5u/RPe8B4qA9WzdjG9aF/CAP2TLK3BEBQ/4Zk+LRh
PD/TEy2qM7qSqWkuCcfSKFT67eaJorA1h0tqj91ao0gnjR014t3iDsvhGZUTmqDoQhrOoWa+KV1e
eF8xKtqYis4wR4NMWeL3PBRTrhb84SKsqEJLA3vppAdkNRIA/wYiB4pbIrYXPJiLMxJCERQgjAdV
CX7P0ieUi8tStEqzAWdw7AR5Qj3NIRdg6vUwmFHU1QW2wpgYwnq+QhtcGu9e0RTSW97gYZwo5Z7c
0JjLWTI2UtL7Pwtr4Zl92AJPdp43g9l/+8olCyTdx+47fSiEZoq/vkwDvrAnDKnQsewzPBm+yiUI
34fiMnzUHjrV2qlDvnP6V+m6bJRjn9tfLOB/0NCcjGUoZFZwuWM+coOkx50aAyygSZ9de2Ixpxwn
ayeGzNqF6d/aeQK1GB8mSU775EGMNS9uePaXgTtxsuaMScFX7G3ENvX7YB+NmXXbxljMluj26HO8
+cXjTsgmGjCJbFEJN1QY4OAdWQmqjcAR/w1SRyRiT+CUwSWyQs6LcTqFl8rzuytgt+a/w8lw9hm1
bTMcHpFRu9bB9mrc7wsR/2Y/DIOUmDdiU/7cuX1l1m+LAYSXViltdPEtsN4US12lfU11/zJUy32Z
7QMM1eaNy8/uLh9+pSIcKoFYFAKeB91hkiVQ/zuGbifE7Zb+N37RR+QKPFwKfppai9U407jpDCG/
0aFh8ZOn2ddNoM+9jRk6nW0trhQseWQWVqfHB3cTH3Grj4uWyABMiRmYJwR5TjBsN2d3Hkq4XfFT
SijJpcmcdulqFHgLhoYPL5qN4KzGUvJbT9rVy19zbb/uXO/dPvlqJ+o4SDfk67l/mfvWMHQEDVM+
aAvwC2w3vI2qQBNzal/LIABAPelV820x1f7X/URc4sr3nnDdj5utc5bdWrNeQwN9aknQIp9dWKVx
BfKR8ReyjzcvR+TVEGZvuj4JgT5lYHNX1qLz7IGf38Mto9D1yXXeogyDHR6xwaMFpEdf/MCTgyNc
axHMH+AMYbOPCh7dLq2NQLTLTmkLhtSE/s4mP+F6ugNDfFsIb1LHnjH2P+zWqYt61B0YyWdzFWOn
5RygO0oDr2dcW7UCb2Hz96JMqmPYUBo/ok9rDg6KIX4MmhprASkS2H9nVzxNF9I3T3Gs6S6katn8
Nfz31yaOaVwAwP1zbspmqdzPXl24g6vCp8B7Neu+iIZWzfsvWp6an0SO3mwAbeVC03PK16UQixYe
nEX1Dzcjct184Ma62M3fOdBv3blk9Q+1oYG+gBKRGZhJj+kxbizDZ/vllGHFA/YwgAKXdMgUYbu2
EnxP2YyUut8BGBXNdN/mHUa3nkaQAFmTXdm+0T9bvYbatHT4OOkaoCusMaW5WvGSlPWZ0+/XLX3c
+1Ffr5o+bdj5tWr0jV585XccHoV3F/gkE+DhjNyYlkYgkVAd4OohbOk9H7gdBAiTJQChBXErIt1c
lpBEWPcdYwct9Ukcvk5bv+W0dTPQ8bxz9SGlYEBb0RzlgOdzHK+PzXVjBNTmY9BZYqmA/rzSio/m
RLu4OQV3MtWnkjnnoMaKgP7C/7ymg3snJmWfqGgmSytC1IxN6f/+swrKUk3zSjtQEqgEVlh6Binp
YKyzZhwEMtSV6qDbRZfIAooNVxUdXdgdiq6NgM13aKU3oMCgSvSn0pOsUi87Z9lg/Qg+O160eBbr
43NEyPq6TbBp/sD3GA68c9jOWJkfs/Wx9RzKZgkkNrkcDVGbVW4cWvxwUqQkdiPrYwtK6/7mD+wg
36/WkEVaw2RZ6cZDp+G+zJ7GXofjcXNL8gPC2oGzYikrsR+cQIBLHRzl3ddTpvKFGtmH2+tp5Ib2
Y1TMIsFisgdHXUkHuNoSSovptlFwWa+l2qiWk51jYZP358P6NWztIt3LsqvZ5P6f2Z5YFz5m0Kph
cgAKiiY5cual3VhI8tsFiuohzXaF8A3tVErc5YxUpeOfA9pQ9+sdqC/5UREI0zNxdqDlYg3gPRq7
dTazvhtvPmi4q7bsyBVDydFuGaYYap1sujppfPtR3WvuA+WR+/cNV5vfC1Y5NVxg8wyOwcxridLG
fLM/KCFKR+ZqdtrWbmd1KAXZl6pr4AXzWyEiTZaYNyV/iTNRR2AfWnL+mOpbGxgikcEmssDA4zGb
ZKOuxx7ruoPlTgMQMJArRIsCs7SRbUSRukBKduvUTg03foZ+QgDpsVZPzylp4q3zed2xPH8CFPFV
lOqCT4Wle2oQxkgAoX9CYt1AGERhdqEoJxQwzrhdS/oxPdmUosbF58EuxY2xbVptFgIcH3vZ85w3
GNjDql0PCaBf2HBvSmzQF8m0WOfLqxiFoOc1T4uWBbqvWtxH0hAjlmUs48lwyCddDzrDZrmOJT86
Wo665dTtO58aHeLZc77gQxQsD3O7Lx5O61lwsF6nZnt+3oMbYTvBcaXnDPfFjFi32HcSC/Ex3LjJ
6naOlRAvxwkYGn/BH8BNOtj7cS83fjYLvUTI3gx9rKc8h4WncXffByQ1Sg1QUv07qqhZox1PmqxR
dqH6+MhBH/OyJ8havgrvqDr+NS/SXal88IvYmalCtsIKwLcN8WRdcSCdY5PgyrQNaZAhGkIkG7tH
/WLYMh1e6jyByYKFxQTZWO6DTjt0gnK20YtguhIGAcShtEVNnKLtM+VcPm7Fl/C24pyjT+cwpUJG
EhroxPAtkwAybvC/Ydbk88srYLUOjKsM7z8OiJzLhpZA1rXSzw/+MpiyEjbPKhTNSTi3sSLkVKE+
XDpaKcL/iTvWl5Q/XyghTYdynKTnfJhbNQBTWxHl+L9/YZKgrH6POQ6oNbJGDBlmXVbj5rEy4T/b
GYkyOKP1QbTDvQfIzAWPjFaL+HVjZ+Ae0UK5cjSrpK/GOptvMW02XYYvE7ImXOnSSbZfanqac20X
XpOoQnMdrUN1extQX190bWcCtEGE4t301p7LsnfS2ZA9YcN0ItIe95ixli5oel22hAjv2MHmD52Q
GUXCS6g17169TWj4XqpqIzyCis47dctEKDLjZAWDGq/1LSUonSVNQfJlyLWksKO7omntKjZHnhXc
wx42G/rfDCuXqgCnDhLHYGy7nWvUR1cCn4xmWok6pLITjg6QYds93/QPjSsRMG1JyL3MPtJQ8BTz
K5KnMYuDxXnWqFVN7RpBmkIOjj7qRYwuL+LKcKuZ/HdOJq5/QUgT5IFKPHFVQ9J8POIOEuaxfa7p
em2OIl1ZwI9knZKaM7zbN8tb8Gmjjq664S9ZoWQrgtlpE2Q1dOCiEsWgxjjRAGaG6+X2AYO3hlfC
uFbgthmu2pcddW+KUzXF0zKVCvLXtguwyPrbsK8BWEVOaylAjHAFcnCsrus7cHeWhk/K6pwx4nki
0rA26PVOYQF5SEtOTSzoREdO1GhNNjmDz+MUViBCKqGk0rb2IfQzifFXPcNVV4EQX0lWaJ8H+/Fn
OB4QLPNBHBpu+A8laN56iihv1ViFlVdJEOUz39W5Le8OtITJDwkQzlKbATby6kSI79lH9XAA8OQE
duU1Eie78x3gM+N3bDSIOSJhjGzHgDAXMze+F7ugymSG+tpSS52E1bvYO3piTHkNpKygK1TA7sA3
jyjLugduOJJHIe1w2++xwSPvW9ILJ4ImZodI6IZX18caSbk1B7xVyjjCPGwzEWD+H7fO0m3SVQjw
4g/50ZZWx8Wl5PvFm3Upw4Z2wplBSCQaUoFu5ysbUQ6i7lP0ZfESVZKIsrTB1f8In0QobOu67paU
uDGHji6ki8PTOtue1rjahOPXEsOeg7gG6ky/ZzyghwJW55E6cPhNa/sAo1Tj0EQN0XHo0zts4FkW
yLKzDGG+1mPO3oHG1s68PEDSL7Q5y945y5bSDt8AZv3wogHBaYkaF7o5eIVd+nppqfCr+jqKsjwj
HfQ0xLKdxmkDBU2cgcx+EMzt7IPuH4StbFq/czBwgCmpeUaYERG7yi60jyaoYFfopS9wjUahcARC
xupdp0ngXw4cD7yKt7qFGuqlaZOtUTpvnhMZ5qH2W0EzGhO/4rrNxGRoLJBzW9lNLLZ6NDYpfk8R
STKhiKlCMr/xLpYDLQ50QK9mD/6AtCV1mixK14A2zQMg41Caa/jC5xE9Ee3h/IexZyIP82QGsbCB
ykatj6rzt8sHe62sOgNABYe5Ts0y+rk1IoVQ0hKZIMPaGAMVEAeokDyfxzdpHbgozc8zMG1SU40B
DQlKd4tAWHGqNsCMANT7GL0mXHG+bvkk5B4+uvYUlFtQyKADBOMcrM6vKmpwEgRJCkIygDmbjigO
N5kipYvtacT2h3xRkDs7MgEkZlEc84Qfa3rx/X+FgUXNDoDW5m3oUTy1rd8iwWThocCTpgNgEU+N
GhUkviFs9lSyUkLQRRWkd//MpXXYVWQ6TQ393yzc6xAN6dmM+pns6KJ+SPwqrnPA+Vn5GcpSJ2hI
9+9cTzOqfS75t6PGg5wh+MVRKDy+wSszZQghFc31Tm3vzk1XOIc7KTcTrZfJeKkFlklabn6Do80j
+BKtqWs6bGI53wZyw2WWe6AS55WovE1osUBsOhUl01WsKEgyroB5fEdreAljxA1jzbKr4nZ6J5RP
vSr2I1tbePOk1MwP7sqQ4svH5NZsHvntAR1dfh+7C9yOTCiuuQmk4pEuScriyjiPiHDWvD4onKhb
Cr5Hwe0uVxb5CYDyFcpiOIvBetYM3WJvL/wpnLqb/cseImxY3Srt02PLG1c+w0ViwvsbbHaFYCI/
ZB0Xj3+D/FjaU2rDyZRmVIe5wgG4Rv78yFCpSB9yyGoXPyoZL3tDSfLT5yxIgNPFIvrmu596GeT3
YuQ3mVewzlyMcZUv+ov5D0pzmg/lBkmUa5C7d/sQQVdocTysOwzkO8b9LxavimEihYYhqnzEVdnP
rxBx3/76u3lgORrHQQGOOtFaQg+MJCfWfiLaiknQnfcN4lqsVHwMPYNi+VlGRTq8NyWmmR3kAMVE
6qwWwIi3/YrMXrQBC16FTwKPItrKnguFYoRCsmdUs2orF4aPz3ni58bK7qXcGqlEQNNxBVTqPZwf
VPHPqZN+kJIQl+bvC7sssEqUaw7B01j6fqiFr9l80Qpiyu/KRXWPbtnemapWgSUG78Uxcz2ls3mY
QPjMhatoC0o+nj0TDyZaYAjLzg90tCGWdwHs1G9ejOB8xRya7k5CLl+RWvqMte71Gzmbe9ghNG5x
jXpJSmiiIpCrYdvE5/ObbJtfWrgqKu6/DvQ4MB9+tePFDCdiTQna0sHS404HEaFOOnNHUO1q9vIH
XfiC95uFjRiPPHx4yUsd6p0Y4zFweo+WpBl5IyEF4QUPXDOZYl/MVHIxlHfMOiWQpoOHBLjqDkvi
4fB1hhSDQUBC+AD8dQs2HRf0Lzk7u5HGKje/6C2+fwYaifenoJ3+QBhelseG6pMeWYL8gG2LDSpc
4VmdikbJuZ2LbKSm/NkWPZAB+7Zq8BKsSJS950LsUUG1AHHqEY2EJkEU8vZl704AHaTx+y93roNB
YKO8BMzNnH5wwRw4m9F3IsmFj61Jl998pwu6aL9MdxDPXfM19Siq7PsonEk7o+p54PeS0EXtqaNO
Utnvtny7VvhbIZHJobzp3YtaESeEmrj3K8L+R6p98c5bbDAAI5c7EWHYwT5FuTaaodaZSmaXd5xa
APvVp/gbtd0MXWsR8AVbwPDBvIIdYe6k5LJiJr2n6UY9XeiGcJZyZNvfGITXuXXmyS10Dmil2fYF
oZb5NsE1aADt6wF7HO/yjUaxMB8MXVjKHJMZQDFY+SiB7k8zKp0mskme0TV8wrwKfnjnytJmt+hQ
d1ep+lyb/jWVVk98m+Bu/b19RZbSrG5DyQsC3SdXuguVerJekf6GXI/r+3yzvmecC8HObFC4yucM
HN3I1I/vU9FA73MMZi1DTbeapD0IIJBpyRawOq7ME7Vu4PAVVin6UO0/C+TrkkiRH+sh0d4BjXGx
DXf3YU6PiTHVhT6ugCwm57zidRdA6bbvXsAgu3bYO9MtC9FanvYGcDaMEmJrQSsk4muLvZXzi7rM
KYrhIsr54UVJvf+r153cFWBvVboQ9amV5H00fQ5YFB4PMOAee/dbKwEL7xrx/irWiatQwIq18Z0L
6d1lvL6rCWJyzG39PNhE02TAqcLkuXTidI838XoHMt2RILVahBY0xXNaIKgiT/hcJP3zUsb9RHt9
51YxSVgchOQtBj2x4tEKZpxO+AI+fYOHXR4Sgy+pTra9yzMKVTW1eVgeiiteLLQaM1L8MkPOI+oz
BtBmfDZSQR5hoYCt8Q55OGJCFQGIvP9ncFuLYiKv6FEUnN3yG9xnW01Z0aWP5vSz3H43mMV0XYhD
G0U7IqoxFV5jsLu1Tv2wiTB+iMpfcdIpAcbMB6Y5uI4tCdL7cbwOBztAugz0XheAnP5mdmG0U66s
UPVzuV67wpfWaNKg7MZcubsSr/lVB/gCV93doJRd1UFe4m90cTWNIeNjlxe+LEqTqNaKQ3JdY7al
Gbz7TNHqYEubh8pqBHN+TuGzFyrxnb1NKxve9XVPYYWH/aIUKX373TJXyXgdwK+7IggHNNPPMOut
VzZjAe0VPGA9u9nfYqreK7/2og1WG2RFNPY5Klj9BMAduIK1WXrKDFzsS/pDc/NCnJAOEfLrhrE3
XEO0c1txXDRSvTPU2CPEyH+I4J5K3uoSr62YTGXwUY6efWR8/9fgXT95LeS+hr13GdlFhdS+taiQ
2kYd6/rX0PReycqt+WdxA6PkMtnVISCkpPhbHyzZh/R5DDEypuRr+wTxpnz2lHfFt/xK/2XwFa1E
oYxuY9xab2iE5+x0z2xyHHmiEdsGMBu911xWMUbNKudvTxEESHE8mCEqg+jjmrwJTGJ9NzXFn4PN
2942N52LyeW4SCkZeaitRc8ei1nDwaKmLfpzyB4chck2r9u+UjArGMMW69IX7NZuslsIRh9qDlym
W12tSDlgAy6W7pdyvS/GyhLgd9JpPvR0P3+iBMLQ5GIL/d45ql8UfBNOLczqpAlReRnLZn8ZskCq
7NipQcy4hL3ZKTegtX59piTLiOQIiPaBKBJjHNEz89MuIAzsDjp/RI5rLK5K0vvC8YLYsaJbTXyo
imr46XEWeY5yo6ByuGFeXipSrJWzvMFvP+tWPcA0VXxZWui+p7Z0z+jgCsKGWJUf26sXDHBcbcqb
zSvzp9ydGEyCRajL617kadhiuTV+ssr6lVoOpBYbTPYFw2/oafk/yrlFXx1dbZ4QPRM1mb3s9521
Wcyvftvy0W0EJV1ljEDTxyfTjDePh0NktAA9AoBMYB6XtHF52zWD8w5EAnb7GC5K/vlkpVyG4pWM
3nUR+A9Mmz6iQdIAelrKq3ghsXfDk2ltGtG3AgzkHGj7bAdzA/U5ySfXOLLt7fzqe8tl0n/g8nwQ
2M2QZ0yChkmohhhEDn+7tp/Q3iwPxotj6GSwU2TT4JIthcHeaa/RfZi1lEsLLitC9UqVyCue99+8
RpQs5rlE5AqcqHgWysQlhsmeqpOEiPm+Wh/OEHsNrpBUbxU1dy0BzxpLIiyx/mJjxEN8KweQleOg
xVC7ixfCl7h3X6qRxqRtGqjAQGKAHBDrMP/5Xqagmm5rjcCCAvUT9A+qNemBQrQbnkBWGcZW7qE3
BOc4IJX5iNOZuekvFUvWqm9j0bIPoAgQ3BWxqtjpzYyt26Z1rR9WmDkb9ngLsgbFaV86oTtKK12r
GQobgaUECc3h7lpkzLKffcqTO35ubvWm8jahHKWUMEqXQvclfSi/uZx/xNnq9EJYEufcMKR8dM+f
dA8XrEkGypeB9WCzV0xvkbNrNeAAZWZ9TPs9QaKa80Vm1fSxDBDbTvdkss4QJbSKqazFC/UOJ7OB
CpLsDljjoRGVcZOyECv8vG6M5Htaoqgl3EQW6z16W+Tuk2zvBanQpNeKp7FhF4uQF3dlQNyi2pux
4nCEjTgG+e422sSl2Tb/5+Q/GUt3ab5A/PAQZxRUMHM7Zlof4/2Pc+Th/yw+lCu8psAWjtyna4SI
8udjAgKVMRELdM6ZC8fL+pllTZfHe/63G3KeUQsu08L3cADx/Q9O3G2ry6MlveLOta2tMdQm45GJ
MZvf4rODDKkV8KMdx7j/Es90f/WidlLuooX1m95tHP90GAQ31zYmgc6jI0d4nn80DJwwJHnXXLXd
MsfEsdkpX+nP0rt5VkDR29qXRkWboM2TVUEL6WN4r+P5QlGeQDP95ay6ZqWwTnR8SBK5STn7umfj
MwQj9IsvRgpshCrGYC915zRbV9arzoG5j72MNVN9s88qKsWb5vy2qYb30/jJm1ODf6x5QUh9lmoG
ATRROxZPeJMk4L7zZgE4TNCZGW8lUnxKpUD/oLiLuLa+srJafRP/bU0eq1ZQZnorv5vR9o79SHRS
ul68PwLwHoh47bsSYrZ59yw0goUWPNoQFKrJahS8Agv5Pdk4vWgO2roFwogxBbWcjWCxD5I32Fd+
l0OqM9sR6GGm4f4d0Rg81y00xr+ucU7gTL2e5dibE2oUHD/QR0ECj0ZqX/4gfExt0SMaWBWNkciD
X+CKt2607RvD9pXyUqCqlscZTfBAeST7pYII+RU6HctKQ/ab1UmP/7q4g8XJdxnykVq6AjYT5CGl
Sgy7qjp5sHxpgFxTQfCh+Wg1kH0cEKdBIWDzGvBL/6DEHwDYevEXgBN9LcKJKPf4O7Tlqx/hB1Ty
DBRZMIyfsNQSyBWBjL3OFRonQHBFhYSg8DqmDxMC+RXXw7hvizggRdgDRcNyQRcquawtU2j4S0Lm
UgpJh9bUQGvOfKDX3gmrHkqvB5/qzUd7vNSAhQlMZJF/NirKinbcR7kkQQleVazAw05myC2MFqAF
nQUj900w1UNenh4F86KgbEZYFI8gACATZU966pAfTpR7yyjIpY2mmyKVCZg0p1xs3dR8yBkwcOek
OKPvQspx39L8wZOuZ83/E6w9Ry4aP1TwF8fPa4A1RlhMfZsC1vOmlaQZ5LzlvwCFgsngXksGuk7b
85ZKrRClEEnWMxbPg3D4aNRagp5ZMabZJSAMudw/d9jQnCvNvA+tGhJT8eupdquolh1Rpkw/ZMrX
5kd+A5M1rVOnKJA/htEx/pUSSuw2H39jbZJxXB5Eg+EsZTAM02362GTTI5nsJ2RJxUXWLkhe7Tfk
tAaduD3sn4xe5GacPzxB4cH/jf/Wk0wKGobTXuaiIYcuCbWAmzszPzkJCqocMcd3/breirYo/Nnz
BNtPpV9yAA9P/lMfZ5JeB5KaJ0mfFF6ifkNVCf2KqpCG5M8AGaf5I42geBxtOZiJSv2ladC6Vnkw
MSLXqncwDV2iHjENYhKFEincgGiSdzpzN0ac46MwiDEFSE9VY+GzhhCRjxXaOfykujQ6DU9xSncP
fK9iNpgrfFYAkwvJ8+1cy/11tt+Rtiwg/OenABt7zKEXLW6nvWqHQNYEcKuHD7iROQ5k9nRgbqV6
zfp4dh1YJVeXXLk3o/K93xaLzsy2hm93Z0AXsoj18qai2J5SiPUesfa2cZSx8/hqa5Xf0uCQ4Wd3
CcUb4aiDKqed5ygaJLG3o3Rxi5RVDkXtj+vX+FVUv+RJK7E8Duuu9i0TQh6Y+4jQ+Q0CZcr8+CkJ
85s6S4xXAF6LQHxVPpCOQ9MnEWtUWMLHqkVYt9KYs+b8sR8FjMQoSlQslMEHKxPjKKhgYYmHls/q
t8g8PxBeBHAd/91oAoPVkKR4lvW8KCFK3mI7v14QMW2PmrUU3UVyI4RVIQKF6zKkj1xtDy1/0vvd
W+YjNouoe9C6IP5MgwU+H2hpJfGOGIaQXBcL/SH/i0k76ZDKnVU4LGMDQo2zcFMYmpahKyAW9rg0
nqP1MxneW4zm6btBzD+zjG+bXavytUBf13h59Mm8SnqbapZqQB8u444qE4LPmL2hodZ7fff8FQ3q
3ctU5ezYd4L9e6w4eDpzMKEjn8JMkIrSXovfBJONSRpfVeG7ECM7OxmdNjwiTGkp16O1FcinruiV
GUdzAYVF9SixJnOn+kO7MaD6YldPvm9xcOYkX2NQIr6JK4HsXbUAZVP74MkKeCFB5oZrXNQhxD+2
vLGeqA1xvVe8gI0NMIVmvqq+J8a46BNGKv3KYysrfcIcb+2o0avDfPaY6/+fJ+7fsuMjUQeXd2/5
2DGJpklfpuLOruHVW8uNVB2OAywe2DYYo/NwUMP2L21RUGthuoU815S1K1C/R9KWHCNYk7MswZkv
tamdG8Q8j52cO4v5+dJrDRF5rNoaiUr8qf93pj9kcHExWVI+zt8s1t1mQBp6cOfW3lFslIcyMSZm
Xv2bs4FvaAlBn6vsS/0S7MRlRADwmZuOSeqpFKBCWd6ITPv97FeYaHe6C6nbDuxClGzNpAnZDD9X
8rNwDMISbZnnPUMq3qmGHswC9Tg8uJMG6a+lF4k85hTDFtguoNrCjdnQVJio0jcr2fac6tuoYXbh
4FLxVVixJKkaeJud4r1nfnNV+B6hG9H/OqT1wfvPUT6QENgEvqJsH9b1z9ZG3L9swZfYYbD7nS4L
AuFXudhr56pP0YEnj63N2sNJyjUbMG81PmGxwGS3/+6GNAM0cL/3uahJzatv+8KLWXG3Ommau8rX
0Kb1VnJQFPCejsIAoxFbX9xtKAB1mv+uxGof6UxwN2pd/0YdyXMOitPgcPoTL5BdVuJM/JB6DhXU
7qxksR/QSvVOq7YrOXTwPw3WwnBMlvSSxdtJ2hfIOWh/8oIGUFaY6gyOEK38pPSt5gmdwtck+TWW
fXQjVKX4J31aQVSBaPBSyqbeWMryPWenM8mv23yIt0SNDc82X6CuwtLSLcSKUxQDrX4M2ZO8YDaW
aSBnZTJDxld+TUk49lHtMnomAy7+7TYM0A==
`protect end_protected

