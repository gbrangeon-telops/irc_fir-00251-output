

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Gub1VXq/9my70IMNYnI+loF5VZ7ee86ZBpAGzL5j+jwLQfPXAWQ9vuaGimuQWfCvI177d9QCmrcK
lRbHtdPXqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XCHJyRkscuJOpjxAlpPvd15b2tV4+cleGX5HVVJ/2Y6XWbVNSZsCQSUsTkLA7IyKge516I1wj3zW
vSbDpitOXWUELSO5CG6d5r8ZVemvSn2BJybpLquf/4fVeS1c+edRHNf6tkj5Q4P0LsQat4mBIGGY
5hCeyo5aPtqLWGIyMEw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RqwoFbaHoCNWZ4v1HvZQji+hXgCjT1Fmm8RnwPGBKk3/N74/TfbSFLeQsQ92UsPWvT9gifFKCg1j
7eGei0ot9ncWAfgeoFsw2zoynofNtXpuT/2o69ZZvCyc9OMmSHilEDslciAlUOrRZtsCwGDHNVP2
rJ/b+v8vvCejKLtIXh5C95/DXV+eEcsjEVRpSeKGeZ1MtzbV+fZPJnRzoH2U025UhnP55OgE68T/
nVfgRgkiVFm7ZUA/Q4uTOx27LPbQmDFQ6plepnrYm3dIFbr3WOiv7AWG29Y9MZiC/1j4MvPp1qqq
xE8dCNkJmOz9uD4DUQoSIb5VP26bf6BmGLvFDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uV7zzv9Zx+u216Ml06an9UEqL4ajf0AMjc1K2s6n9qbyEnUVTSm6yFZ0M/IFYGglaG6jdDDlz4rd
W4zdLmcu66F6EUQtwXBmHtk4+/Am3fKB3kIu6GlcyUoJhx3DF0omCc81HS8JxypUZEAxz3C538KP
dZmq/6pOZleIRCziFs8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c2sM3Lkice55qsGCUzeim6Qm2yWa4rXMhx0Gil9+l1mRl06adQHebvNeaVnD5l4UfTgDiNRnixMg
t4I3MixM5k+/dqMphg9yh9uQH4HJHJ6CTIPJ7b0uq0QUv2e+GjaxWZa47ZVWMUHJwpscHTsz0hs5
a4sgfCiRr4cQxV9i8u9cWFqcZ4eu+RYLEbH+mYK06INaK4Fg1vBkwveCaGhKFtvHtOBXP2o42BPE
2i+HCKN5sLyGLlDI9h2MogiDBJsNAtjJ9geF4nPG0e4nijR/pyFXErJCeKppN9041em95AkpK0CN
GYWuH0jkznlTfi9EHnlKl7cj5ibz763zI0uZLA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10784)
`protect data_block
5lyxam+8MmLQ7ion+XNw2V+/KeH1Jfk3AWwa3j0r3H7mtgdiMUTBH7PXRgFvRUhNaHCGjYLF3H2W
WTcuCZtr/BmDqchkoxluvqq0Z15Rs0GuBY95JbSalA4QV+vSxzxjf7YcLpPgGDqObXVyApXe0rSU
DazRm0FY4GguHnEs5hYrrKt0uvbc/rq47H3ZZcKDJiAW7iX2oqgg7fzPmeLhZ7GdfCnceS/QAJIY
OcopA5lc8LS4Vll6zlS8y/T2qToEq3C21sUWlcpLa6tJnTXjOX3/nOmxZnC8aG+KRwVFODh5/+IX
Mo/0xz2aZXm0Twpbz3hTn5SDo/3n5yYKznwnAMDfQpUV++WWySAnHZLbsXL87jzvByErlCCuTo/p
4kjGxNMCB+8xsLp7agVKeeaWUWpUaA72ZJDTzTMiCeMaBZnmUo9WSZqyDVZcQL+DHlMKK1l7u1cX
oZwTNOHBFE83o69RNW6GZHdu0ydJwWKOefo66ukXAyr4smHYL2ucVOxFxV/JsAKXx+S68j9PSSJz
5VBN4wlCnwNDO+BTPXDhnVi493UVBeIDw25b85LWef9K839sgDfxjEuGoP3tIS8yKA38blJd13nz
Ym2etmdB+aLt9SyXmIy/v37aKU2KkZ/elPaVdpz17I4sstpvYiWc9O08V9koqArFLRA03ylht/ro
glK8eISxVqOYyaTUi27JeoTiteNCv7P39SDPuW8RKB/UUI80NuIWk3NRrvHXxIbNW635nxq94mQv
37Xy7J2tvBwcExtPkp3X0VD4I/HBk5qiRLynMS9U0kTZAC24Ysa4pVdAZN0MO5OrusdHkBEfldSd
cLxMzktNgHvMxYW0YVRiLlFHCwFFewQ/fK/4H59zfgm5Ct5zz3XUcnPZPYqT0pkOn0FUlyH5pQ8s
gsTH3o/HQFH3ILxrPFEerm/JJa0BvGC7/3jLe81zxhtWuEmXBGNwEgMA6eoOqUTDUfzqGlTE1yuH
eBghM761aNrloHDj0zGu1thftPi6M75paCpNCPzQM+bweN6sGr1bFikQbYWoJyMnmhdk4g87g43p
WJNTjBRq6oz6yT7VzhUPkXmvjwgqUHOFT5k14ziK2VtFSzpJ33AVjfqAJo3uglgBmWSYvfhcyTH+
j/W76vf2N7W1yL0+TsPidjN2HfbGJ31TjOcnL7EaJHU7I98QckBfsPrw+/VuWe/TFRAtyXbT9Uln
NmQgBAQTB26NVxXAekjRibCYwdLvWp6Nzynr/LmaFZm52rgBJqA6v5QrlDIsQNXY7+gRmzFJ/D9n
1y+js5Wz7/VYaNG0Nup84V/OZ4EQRDIliGpg0ApfK1QURmrg3G0vz0VsCW3+EcWHrs+KQEmAhhUQ
6lRlFLT9A36vjRNQmzI3olXX9wr6MA0F20YrFR9s2RrF5UA0jzUER2ITSXLbxwkUDgAf+X0qcgp2
YT/y0AdTF/y+yLa6bCGE/Np40fH6xrgjRUXtLq/+BMXabTE6nMPsfEIzKkVBIMHq3M6UR77A+HW8
07Z7b6VQqRI49n+l6WDx2WRlcopxpHZW13/4Q3ReESrw69W5djmPFOW58UZxWIFewdYAgnqQphJV
lUYQGViQ+rbQH1WQOtWD3iVgvqU0s9dly9Q9k0zQT6AKo63Xmbs3vtYkkLbeIDNSWp5iXZvXe4Ev
/D6VDbKKjLS2taWS0BHlcFcEH+NaAP6IHxpva8AA0HLNkFkdnXzElvXkYk3miNhPk6RQeOGeEu0/
5HX+uqYoMAlCD8iJmV5ooYnrnpC8BO8HkCG+qBQSBPq5XN+ZR9cu3edwP09POICg0O7bwHTpz112
5T6m0RcfySzTMmquc4qCMS9UPf46UYX/hsqnJ6FojFzl9argRC8J/mjMZjxrl57fg4LidUknViOQ
eXIwJ5n3QPiy8DHHBDLVKPtUYa49jgeflHbEQKoooIivjPoK4Gs1Dv4plDh3by6/iinj9JgRTJxJ
pwGGkPz1ik6KlA5BB7LLmTBdu0F9ZRsqSoFFrFhOkqNTha/DMjM4C/XkdI1r2bOITzwIcxggJ0q8
f8+Q0BBJLSn8h3L8R8zuVNq3VaSGV+eV0hZXrKU57lteinw4gRuVW7yaZMeT2hvcx7WykjENCzV8
AqHSzvzaBTUbeIa6xCOmWNDOe4MbstjH65SesHVp96OFFkK2o8cZonDUoHVsgp4AAWFjBMbysqcI
Eg/u8LtwhIBGWsPlFOV/EteaEFFhzCv6qievedy5j+uRTW4b3Qe2/2s7BHIL/wnRoc11h28G8F5z
+wHiflViatcild77LPmvJLWJMTAsbBZrShpVWTcjIc++rpbr6FWEcsQHkSBBhd5yu2ZqoXkiXEQu
ia13fxmbAMPQKRW0eP0VwyQ1wsjjt//P9n6svy0hxqGxuVK+L/kPOB7LGuGRrTvJnZPonaLj5gRP
dIwzA3+t3d5uGwZ7I4BB+FrCXX4l7xJzGZQn9M966EhQKwhDYTxC5y9z/AOjquDG92wqso3JurU0
/4CNTSA/Mqw7DhtwrMDdRDQfc+ZJT5l5E302IDC5J7KCNE9RkbvK2zfmLqzuol4fyRcp2Lm19SLL
4EvtvaMYf/8DGs72jZ7lrWZ6fcJU3JOe/ujQD5eS7PuXgtAzMt5RVwGuuNMmfYNNkYJxPE4mQqxm
BtcX7JZCLW7+yesDzWN7XoF9QwJSQO+eT8IBO+3/TtwatFkUE8mheMbPN2SV90L2Gueaz523/VIK
CHoqtcCaOxDT55YiWSHELE6gSEuALNzXxkOZ3AVTFrvaDKr1jmiIUuT84VY+QDS3H2++S+goCi5y
kmwEkA+4s9RfQuhFAT81Ba3uMTnAQ97L1Yf30Og6vToQh/T6eBKuMdrqIFr1AQmez9o2EsUP415e
6oIRTvY5R8dDsHTGuLwvAIm7EYh4Gw0pNhPbAHrTZiyqgpAswVtJkpEw3aSmgD+iLBTWceGrBCvX
5dZsfwwsaVEpKGppJnz1ad7Zub8orlsYQfefLW/jZfF/L72V44nb2Pdwmwl6qf5KyKpO9F2/FXKQ
VKhHXh73bD8AoID20ynQ7GlMtonV8W0IzZRWY5xgKUajTypQpJMf2pj54PDEu34D4bvwCejrs+Np
11WfqZ9sEMMfcRuuU5qpGEfkBHfoz1DYVZnNcfo6h79BOmrTRxFP3Ufcziso1ya74y6vkM+j3gvH
2CfLnBmHfOP6b4Q4fGlODuUDLOam0HxgRDY/GlMu9NVIS9HW0C6VoqYdGJ8wjgONiTzK3H0JYTEf
60PgOcXp6DwriHQOf+EDihESP4E9O+dcdiOvbJJ/hTUhgxDN0Ks6WoxvW6kwCmj1egC0YIXn3HpF
L44lMUlDvWSSVlMqpVKMB/PmF7rv7bX07AnC3sFuIxoDm2bBfttBB5cAw0Dh+1H+BtdISHfQ0S05
pmKu0itnTWUSsyPUbKbRBdnHqW3YJ7g/8i671haIdpUzO+bC/72ElMvXRKbkhlLkeg5i3DJaD+jP
0GZzage3aHMhApPrM9Of0AHEQRymwLvkCSS+g5mPLQgY0YShWA2L9sp+xA//O71gn1vvV19ApIrT
0QC9mF4nPdpjLc50ZIfwKGMs9WTf3XDSnceAbo0NiHwRmq5SkspOI8MN7p9aHcg34plUh8woSmA7
2FHmdxx+uymq8Fh1WfRt9apXdK6deHOjiqz8A4SPYgQisvTF4BX+TBefdVETy5JjkQhgeYIoalRF
fzBDKu6pXRc1H6bqFfntYuM31wq86K6jrdJLRbWvJahjkIwTFxnD/IodyUc6RYBpr3G3XLUyLOvR
wJN3ZlQ2kqo7Cds/rIIXJmDaATDeOcfRjOkHHN7Uox50Py9eanBuc0rd71ltkkUdCwP8N7L59d36
LQ5GpfDNQxomc1QfJQ60Q9TMDzpNleq13F/vPmUMjKs6qe8ku+Djh17XKtYAKmhDi6l7iqgDqOyo
usRtapNN+0OZCd4rco9LwjjFmnHltlqHOfcceR9AKP3z/QESK7Qb/LcYDmJ3Rj4rTBzk49b4Ko5M
BTyzjnVIZhlQcT86VuKRi8vFXMh5IG8Rsv223ccFiIrW/k+xDZZN/JOPBU1n17WM/EmogSeh9OWP
cDRZbuyUFXHePeTryZSM6henvEY+mDaAoR5N2S+7PnHnMDO+HtGUEJeB5Jm5VlIWEosiEeJoBe0q
QFfJg+bRMAgI2W7eXpJfp0nw/yg/uYxX75rguEddAvm4dpVUQlsHqOnqwk3qRL5T6BormPPDfOv+
3gSFA9A1e+v5lkVFXGNUhlktaA1+47AAPeKqH2gzncaaq5lD55wcOuOxvUxEomjbLnwWoxmctqzs
KqOrAL3NY0y3XaSb5iWNWQg5sQhS4nXD3AHnkEmxgPNWxGrui8gnev7RspwGKHTa7sx/67hols20
MK7I2bwZb7iRrWZZTloy5M7FeCO4t9UlBkkfIwXLEVFESrSbC2+LQ+ZRVFNYOfEWqWX+tVdyd11O
emCgcLfR0epkrwLTF4jU+Esg4Nzw/W5ub9OjV4trtGHuAExVBBMpWGLkKKCtRJDjdDettXVIicSO
Dw4fgWosucz+fpm92wfWeoBAuFxYD8lNkkuOSVOViE0MRyEfo5KeIO5Wo28lcnCKAxRdNpO72Z5Y
Me1JI4tJcSB0f+kyV7qEGYCJwuWuhupwBbAuvTMP1ZjLTV7AW55fhqP4bkeKw2rquz4cJlN+wzu+
FnhJYDqobge7I0SPv+mBG0zdO1AzAYNFzFGfKblczT6ulWYHxKBvtKQ+j1xbBOukT9/aFSqnTyZw
akdY8PdLFshcXiDFHprelsivSgkdgD2NSS0e6SdahxZzxUuSYl+jSn/Knp7Vg6L3Vgj2SanYZeIR
sufK7eTazT7ZF83dbs4OhjUGamBLL4gG9ngcSzwcvqGIc/sMjj72u7Uw7U7/JkDrc8Hb89M5tZQv
DHO1QXg+xcwZKHxYlIZTZg9ddNie0UI8conMQOTzVElN9EYjLPQAp5ubRegi/HD7rOAUlo1OFdp2
0ZZ/5mJho2bEzuyuFWQVAwVj0Qf5cLnZ7J1Q1FO8X0I8ksuE+DLuWh6GcF4h+JZV30lDtppdYWtR
Xl6PgRpEwHE+RhiF63VXGIUV7nyQ+HERtQMRrXjCMryNGBD8aSiMDvgYK83mTGnHJDdDUEt6A8IT
arbfmls6kgXXlqITrbVipmTLjPLp1PxlDDlYRNNQnhnrkpEx+DfAPFJY+JoPoGoinejagDs4mdSf
oD0YTJWSeMxSmx7tgSmCuTp63q9YBWvAdknJ7R6ZVwNjFYakNAgS5bzIqlJ8fJ/waSK3HUVdi/XY
wMN2yV/lLInRu9t348TyQjh5MN7u2FyjK3xQyBygZbJf/TtRGLXQRZHhq3siC0Zoo59/1A4BTIpK
4a22Mmz7ePnp43T7buDMoHZhdR+n2Eej3JiwFeLfFTSFqWUQKw01OoopJ9Nc5lzh4GSFWy6tgKLX
R1+s/X0LjOsER4ILa00Soi+Uab5ZdHoJj58Mg8IqaUHFlfZ3Ix9XZFaVNM3J0ftrhwCqDgGUWZoL
i0vElcCizAtAzN6RB4u2lCXmCgPD8eXhfmsjELt5D0QR+XkUr+J88u7H0CBv0H1ah0g/30sqYSBL
/dg1iH4uFlzHwZUYJsjbApsFZ1ZrC5ZBzs6kas5sbBs/QTQzWb7RyTTBXkK0xW5p2nWW6iKSWnjA
YlrVdXI7DVtZSOZjCjQw/vIvHulCgrenAHYdGxQO//kjUtg1FHjvOt4GjW0zO3Q/gVsNwd2kw58j
VTPz0Y8hSKgXkc+3CPx4NxKHhImW4180UEMKTb3CrGh1I8UBj/+xjqz9rFN5rml3LDxtKn1LT4+l
jZwiYBzjaD14Y/Wg2U2K38qLi7Ce3B2GN3+LajGK8Wot9wDSlVzwS/dcYT+kE+L/zF7b2sLrNjUY
OWmnJ7Clz5L7c9Xf9mp4hmyX9HrUqW7iIeTmvVj/ga90sbn6UVQNO7N+opa4oTiFSKD0tAMimwLm
ZqSDxn+V7S8xcIXmyprtxNB3GW3RBG3+YDEQX9/M92HIqzfFsAXgmIdOlR5+7WVEqENp9aObiz/T
9hsMffQOsDyRvJ4YU11XdmLT2whJFZ2yfVIx3TAMLG4z2tLPsP0GtKA2t+WOAYi2b51WpAAGlzh+
OPIxLP8OANYCnx7yPHAZJ3Uhy9tG+lE0NEErjpryH0z7Y0Wzxa/px3hz6kAj74FWKynCNtUJY6iR
DNkf9XQ8cuwfSUbCnSmEOTiTWziJ6OvqvHR40/hO07bQW8S8WBRnjIqOyV7DvYCkPs/U0n+vImtx
GQdfyudMDcxY0hHW+cg6wJ0Z3nT5NBl11RIKcs3HzFnRO+ytwvnz33q2oKqZSnm5ZA/0z4+XyEA9
M4RZKyOV6IeB4ZG0IG8nbTH8nGA2XIbZc65td0SDxNCOnjf70PYjyEQwcvRuKx5VRwi0w43nyW3m
uvArkqk4zkNVKFbuOTEipz6FKLDXqmE/8nHMJK5ahL8QXmtxES+7lKobdklse/zongGmv9jRqsZI
dSPVa+koasKh95j+w4Roet3C8iC5dD1hvdARsyg/9vdBbc2qtA7PXGWpQwoHIdrNuSRnAx9clN79
YDNJmrfhOKY+I+dXM96ymhkOo5OjH31Hi1pUjxqSUu862AVD3q7DlsPT7aj0lcF/7j9rd1BHE7j3
f3xpwEXCaNS9DraMhy/WYoPUpl+f4/WlrYR37NG7SOSZt8o9HsJxBoYaqUCWygkCZs8ffzxUxdIw
5C2CugJ9uZ1XXZMc4DvXiItIa/MyVuQuL/lAkM9O74ggw+tYJ1KXd/LQyt2BGQlyNlU1HSVchmr4
0T/9ZGJ6Wm7w8o1Faq++aeZfn/4HBXXzN6o2iJIXRER0vkf01TlRcjhqJcyRjMN0iqFjCBi2KaL5
gHQ7z92ZWQYruOcZHMdQH29hJWz9uwQtYx8ehRsWgvpaSaZ9+KFQy7BHjdgcbT2qwVPyDdsWuMMb
IiiHtx7xCti7v3oCvPGUd+b3ay4dBNl4UGZQa7jdxD+1fqWYRw4ZclbTKb8B5RQIVp9GjTyJYzlV
Y2JrDgUh6XBIjHx5tXWLhhx3vUDiBLfyVtHNXvJqrZHLLTKlBWKjgtRH5LS5AOZnAXlLpbESgM0d
otkwVimPWHefYvqvpITZzpw71lhu//Lglj8TdLyijlM9QUI3UqGEA6ci/ZmF2dfhHTJcI6Nsb3e/
1usvd82bovbpLtMHbMyCeXa9MfZFnGNYoYx3X3i3LL7TLL4FQl4aigzFKM2BS9iYmP1tEBLyB6FF
cy/Uw9wZLiFP7WWU+7kxnfntyHa9YXC6A2DfzmGclDY8CISEAOQ3a1tedejOEeaI6d5J50gA3YEv
M3WTLA6QntUTdqcWU2EJcquYujCdfo84dQrnjy2ezS1140ACz8iovnqPOtIiCeRi9QG5yKSaG6Yv
7j1wFO/oUEmhL5MnB4Y434uzFOkSOD7+EolHf/3SX57qu+vaDVSHFhlzAgseTkJxnx1IhlPqaB5n
COUCCmIYqt9KPtueGHpU5aUZF2ogh4AsI40K66X1e5CMXVbI5SWk8gWzJ42Q7ZWSo412c62sdMcC
PiT240HHGgvyNKHRaHBb7L4UEX9HkCE7GPAyaGaRjqj53Rj5IkHNqEc5NH+qn/NwJQ8bdmdrV8Rj
SEmVUGnQgMkzs1DhzQ4zioyExTR/yxP5WCC5P+Iano49UIKeUsGF1VuBfuWrTc1nevCOvUcwKQRh
kQhLR0m0ct7aZtNHtplJTBpVydgEIWRmCysknup0G4DIz8B0JScoNkbqUJzGuucNN5Xz5+7fai5k
rmwrfkAj7jExhPVuuQ05NCwfeT2VYkZZUmudBL/sHHJmVMh+6wMN1dFN0CXIaV6dpJMG4bhCFKZm
By19KRTyuU49X11tC3cNFdy3kNNpf3Y/p4Hegkz2xpqCMOTN33bJpMka4Lm4MZhfUQFxix4gtNy/
zfqfDO9HXkBMsOi8odgkf2vb7j0gdNu9+Ru4O3xeqnsui6Xh3F28f6PFNC5XCAO6kvLKp10I3ZdS
FRFjpeK8urBm8SlcXfsFvW4YbG6WhkZtOC/AU4WKsxmracMjuSpnp8zkgyRDiKJgX5k7Eehb+keo
L5WD2fmqz+XhUqOZAnjJ91LwxvzQkWRbNoHcjGIuhbCs48fnl/6zWtLtnb6e3EhBje3G2nXCBzqO
c9ytCaul5MhZgjMtKVQCltNaC1/ObwJAepizkOvqiDWdLm32TEKSTumHLL9E6tA/2mVzqb+qASeh
+KL+sDYZq9LEFInluWyudiBWNoDwzywFCDmzaLXEp6IhSN/Y3uaERc8zVfvC5x9hkuW7/SQVUDc+
j8TgzY646Gi6mkNyQ7ZXMlP+TZKrDcLqTv5Jt/7QDLycPtEyEkrh9ebJFRuI094zNTbuDrFpdq8j
yKiKVTxWNFo/ayPreGbNVtNCG9oCI6ROe1POoth+UgjSsBWo4GLmU/2KSo3h9+AejACkFjQ9q7YZ
sgobJ6n8l1CciasJDydTMaRp5DjSLGW5LEIxyOGhqrehwT7fzBtOrAKdd4VMI6Ah8MJcIX1OrkG0
kfGKwKm8WSgAN/4jUTvN//1RREJzdvgwt/a6om0bif7bopq5rQ22d2YTryun08HHnfzHjpQzQzlp
RNd3vQu28YaLHCG2aX1nQo4H/S0BN+kAT0/BvlGCcTFIEyy76ji0709G9shIa7jNl8F73fIxOqPU
B2reTwYqC3PZD9qKaTnIcyCj9wM/KLwandFkKr7PvpQf5cFLIzbN+r8B00D74sr8khA0Yo1xRnP4
acSegude5TEF8kR92i0IiBEUbEiJ3h41pFkT+cH4uDIGgvZiMZfDhSDmGtDYoG6Dp1HkplK/wTkN
7q3j8a47M4ewY5RqFMyr1qero1Nn7LAuEHjSSYpmO1JwqH2TsslzxY2XluXW4bXDlZes5N8CGStN
I31ignjhLdqkHZ+sUj7xlLcQvTgDzy5ZQaPZJNamkxTwgjRLj4fkk29b/3Y6LIlzyX8GdZBpx/0C
58PORn2D7uj2+LjCM8T/z/31Rk81JLjmuLaJotC26uc8QzN2w7iNtSaIVQXG7nV/UBA83BSacjGA
wq57RqNUEml167KGlrLEwU1j2jlNgwMsDHi7Ge/bjBArTy7GZ3gd+6/Ng1VCeNF02nxOJGhvYiWn
dIFkPobzK5mykue2GThL8p30U+mQJONZzPyV2jpPOauyUxs8Q/KQpArsGBaOTehW6uvFvPrKzSkK
olMsPeNZVlmo4reLvjpsBELfpD7EOXtCU+9vvi7bEOKSGxfsRW1nFAPN7xK+XMZAD98xWzlC9akT
2apzbw2h0MJe7mNqINQh6BsZ+Zp+i059a8coLfSLKnRliAWDMplFLcmyvTGzJpmricUADN4ahNBM
yvwEEJvq1BWGmv+VZBC1r12iJd2ildxTHvgWHyr7YC2ubu/IPSERiyVnqxJDowkQsx8y9DSSRNRb
RlMPJ3iWdBeZL0RjZ+jYaMLzCDTo5S5g4Q8LzSALt6utJ/0Aej92mN52krtUL5dTDsxPX7x2qhnH
PabvWLEJunjDirJHr0x49LbcXt61c+Vq65sWKY1NmD5vdJgwQ6JE4xn4O6LiGsk5n+QKTDZtStpK
ACT/zq2rMTUh88v7jI8BwejkeYR5jYb+y3cmv+jzAk1W4nYSH5xOicM+yxrCncNMoRk7zsVTZ/X9
kWAmTVeisgAzghGifezvCuP8qztz6O2KqJ2MLeBjBlNw76Si5Os+70mFuORaxGWNd4Xe7Jlp85F8
CjmAl0u6ROUZJ/1pxVSwjEs7/m463DGBMYi288VAB+ELPGE85ABaBj3cTyeQUeeJUG9oGQx21WI5
PechMLJtvS3uTOMPaH5y/WlqD+9VpKPOTlI9oYq2HBwBEG+w8b/IPZ0R+SVZQ8eUu6ex5C6ovBk3
Fe4M8kR6K2tkGplb8Hw16NmqfnzRWGtZuobV2uuI2mPndAApAmwHQJaZ3FSNKAWTB0Q14WIkk4Bx
MFQnZQBs6SmjjEc/X+jHyKBHJcJwa8VkAIDqfSKtKEMW/Zg2G+1Eux60FOW7o9TFqOIwCx6144DM
Kzj1S8BKP1WHcGCbqh84nj6n1Rcj86egvOLJTTJnmVLgS65dSB/peCLvxZ/i9MxwD6I3UyN16SqU
1OR8Lr+Ay3bJObF867thumeyVba4NdBOXc86czlKn2MmcvzVBKpFpIPWRqiDCnIyJgfR9i6NpynK
BHix0wMBuIMlY9/6xM+im3z/+kx2Y62HzaC4ekXOMFjyRjSpLaB0W6/tT5F+p6JjdoxHKb7ol7aJ
zSxa7Wsa4jsjHsB+EVrVfXV34peu541R05Ji84lJvrwTB6w9cxEUcKfld9tHIA23JJT2OEKGGGGv
9N4iZlgySzpXAJf3PIc2CmcwQ387PES04MXk/8FD+1rlgSXfYa6zlaC5qETUA3cF0ibCZVoNFsTN
+iZXKjGWAlF6a/ebQ06FZ98cu4qpye1lXk4k3ugsAe5VdToPXwxOaraa66ok9l9IC3cen/MR2IsW
k8dnNYkyoH1hhcngjk03mcJgc4yNkH6bBMCAkicWUd4Ahsu0OJ+VpZDDmkpCBjFsMTu08RcVJbgb
3319ThDDGlkj8QDp8SlZj9bRQIr1KV1KSU/ntTgkW4YUGtZQ/0LzFteco7CWZmzDk3LxtdyOLlf8
Q568mqztdW41pJB6fl0xYHXPYebkJ3Wf6AnBlYj2Q2UC4SYyjEcZx0RGniGLX4ABlXqyZ6SOiCo3
0nhv8YCzbKOHnM29SkH4tVfNB4HbAm1ilON4kNmJBXnKYvzh/V0knR04ZXiF5xDg3yYrr566Yqjt
mVKm64C5hFJnMwUuLOtP5ARq6oDIRds9409wdwzs4swYHDoDturVTVy6rvTvPuGnUjDyDK7ybwY5
QqUZrq+DQ7yU16U9Hbfu7rl3GoSDVs1BX5+Wt9RAnfibLWTCmJ97PSfmYzu1nHiOn6RWuFf/9Umt
8pf0aSuuowd55dvRIuccfSN2zdA7tkEl2uYoOqxazRKp3aU81geGv2GRdUR6HHyoWsfX5EVt7zL0
F/3l7TJlp2x2pmCSSeI+e30wU1J1TgXdIh6Du6yD6q+/ilaamgHxvo/Ub/i2QCeAiXMn4m819tDB
og0Udha1agbQ48v4PMLOumey+X/eCVr8KN7lxe9MHDUi8npPfHuG4FIHeerQDu16Wr7UkkWjr6Ob
P/IfHX0Xi3euO9M2eYFThqTsKe0nWjlmJVFPVG29sFTa4Db5WC4YWpa8JGrIK/SQWFGQGH2mUu4w
ObCcVPz+wcfBFUbLM7pM51fefVnSF45triienrUAdNgcnAUmKf7o7Mhq9DnplbEkPrWwEAEnhUVg
MtnOVtN6TyK79IceiM9hywEbU5r9Xd5kjnYVZSRYtZhnhjfEvbeCXT2gL46hXkn8LQs2SKair/ud
X9piMXMBcCM34X8Huxzir8cRcp8tNEkrCKfaf5XJS421/ivccRvBuJt5OSsg7wybBV1415U4PmfJ
/Kt0VlOIelcosdEZcNUehNrrNgwTt8fOzXI5p7ryRm8AJYOFP/gs+/avhg5iAgQnzcZWE30GpRgt
mC/bXtmWsjRKtFFNu61gw6KdQ5/ww1iMTU88HsqDekxE0Gn4OcmBhnz5Y2OasNisWjoi92uCPN7M
iqJXI30wxKV1Dqn1X6NFSLJGU77GMCL0f3V893nL0ByJ7GSTIJEPafOf+76cB2amt+r4smj67Lyb
OC6ILeEJyg7/AQJBw6TDNd9tSVzK/ONwQSvwZsHOF2EHsJfTaecFp+KVYhdPHVw9rRBXj5IKzIzX
fzvvTU1f+GdOa0c8u0rfAVR5n9mnUcx5OcxHsB8gMGfiRpd8N+y3w2fokD1LA5AgDXzqsonLXvoq
UyZsWOPK6Bj+fq6tCGVQSgf9URxOpUNpkgXRFJlQCifIct32TcyFK49VW90E5w2IBdqhOc2rSg+O
Oley/cZ/yvzEG9lXImVy0ftJ06LLjtRO/m2uKW8ERZX5ewFkkWx4PoxoAV+BFPll502oLvn2P+TG
e2qVB54gGn7CxeCOsPEVZAFg9oJls8gmsw58tndgKQ5xS5UNgWsY2Ni4PlOy1JoeHkvvroN9xj5T
00uowBCrw9sgmSgX+JFK/RJlkktKxsF138FihZvmT+4CfuFF48/+qjfE+e4VHIrlo3HhIBRpJwOg
a3yUAEJgUyase7zcOnseSl9uxRZEtvavoJD4nI7zFSmOC5srpgpj/uAPI73sfBmIhxdtZpQILMAm
tf0x45Rpd1TpUiMVWnWAXtcofKizF7wfZeNpzhaMXiuBtBwURhhRHcxMnNySWyzO69RXflQPdLX+
dzau+Wy8atlvugn1Pl3BPwW7HZlD0cnQ4sAqBDfI6EuRBWtzSDAJIatNcgK6ChvaVh+m0YHJ5NO/
OXJoD7az7zRhil4dJf6DoaqTeNRnZ6mGFXwPSY5Dax+/Hefq4/aK+LDzFs358IdeJsvBx+e466sW
VEZt9aFUEsHdGnow6iyFZCwV6FWxZ4ylnNrkMDAx2YjY1hQnSauh6dZ8GfpWlSVNUvTRvLoq3lJL
eWjRqGnHlIguEVJkoBiFyIotezABBS10wYHVGrhfdx5fyMznKmnsM9dC47wo07L7OBIOFLGXrRMU
LLftn6hsUO8Ix6YzOA4r+8OUgbr7RZF8ueubg98A0O3mOPCQLV7iLv6RTMs7GIlX+QUFxx3U+DnK
no52ovztHVUmwJy58gRY2LiOLH2XWmp69Zoa0HMXSor+MqMVEESpHLNPdRlBtSKIKXlxy51Dzufi
n7MTOFHXJUh2q2orDnhxuHPyC4K9BKCBPW4lMS1Xu63xpr8VVLNq339D6qCNwpvf8pkpfzAPFDib
BfCqyyNXck7tfYIkoEh2ypjzmNl7sXhLkCH8kBKwnUDLFWNc64UACPyxWaatg7MdOOR34cbSQ1qJ
i0+Gs5XOXxOehXTb9SL2a4sUsKAqlyAks/o0OMdMaWuwmeQIwPvZKE4dlsok5DX4PIrGHLVoLfWM
DylVs5CHqTUpKGuNM8ciHtFZiUFx0raBB9X4K0s4lHKd63DRPA+4nWLRmAd+/J3lLxGzVWJtCEmh
dNkmvZRA3axdVmR8JMVE1q5Kkt8jd8Ulj5WizSzOreYMevoP+rolhn42wXa5psOCg3I65fyoNVBZ
oIPk/T2n3Qdk85B6B+StxJv2kA3eDPSLjHMb9sqD6xBSJJVASq6RoWjB1ZWxmiVrMdrs4XDBmxjb
c8ofLviiF7LPTeslG6FHAoQa+e4tXrrZE1OiInVzY7VF1O0Zfm9MJt7iDn3DPnzYShG+ZDrEXHHo
VDWxx1QzowBykwajtMdxvTwe+/syTUkSPAK94RcRmpjhjGLJ6uQTcOS1zv8W4WhIYdqP72LrIKuP
Cq73gdRl04XvbGH56MIoHTR9FmJSvQNrQSwq8D81LnIVCPMv1/UlytDqZvI6kPknxplse6UkbsPA
odSN/H2e+MfkfxN5aLivG4TlRctQBb9N9uxvOHYrpovNuul7Tp2ODg59jlCvAJ48LWzo7gdSINPl
r3Z9AkjlF8GajXdbiY/5DN87Dnj7f/whg57MNUmKQx2VJs+NKze/MmIO13r6FF6NmM7unpumk0VD
K45QkbdaVtOl+1gZvLRAtq+hCxi9JoMG7ZOk5V4X6wrOJrnzXbMjJy9aI4t1vUkX0UCBlFHAXNZK
4d91+Ef+uIe3Z/wW2bncdo5GJ+/mnTRZ0KqAwcAysL/SmU4MCdIjpYrWqBMDC72eoXq1yWzFhy4v
ckqJdWz9cCbl52b7mQ5lOUOzmwh4+UUaes8PdPbMNv2sn8mysT9qI0tcKNIlNn8ygPqFp9gNQdrg
CZj2VZohMmWhs7SnseRHsRDY+kO8UxvMGZHUGjjUE3e4TLg/9zCF9c7a+PfVY0F4SACewhryVSNE
ZlaFQUYGIWABPtiCTgCT0Zj9vhSVczKxWnm3o9hZ2MY2zYc1V71uZpGQf47aVwCZCILgiuKLrfGd
/nPGncetzvZk4h8C5RwJQqmlhSqQAQE3W1sY9mHm1Mj+DoNAttsDO54BH7Wd1z13jbU0Co598Akr
zb3QvTL+oB7CseFrmS6/FlW4NLP9OU72Rwg5mZgmbJGvYCWadjMOq/hh25P7PZCOaiKbS7C9W286
i9nyeWJN7arkIfPnnt6QK37kPF+Wngws5pGn0QO83PHK7jaeBOSliblp7zOxZ7RMFi7FmgPJ1eq7
+WHiQHJTfzMw9MTL0RPltO4pngIEyYMBrHL8kBUCnNK+WRnVz9jrwZa16aA0Y1CsnOClTSuiCZfz
twq3xXt5u84FehU=
`protect end_protected

