

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hB1MkDF7gDUjtp9+r0pYANUYTDYvtQO1sWNXspOA3ppM8SYB929/qlOMzanhENZQcOQ3aiyEm3Wb
ozapXP+k8w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nob9JCRq6vcsk9H9VmyBE86hdNvS8BGq2p8Ka7dLN2J7EaHNc5IAaDkHipJixlCbGOjVeeUZyKme
HUzNgZTvjzVoRv6O00gQMvGJEhPJ3XxSJAOF+OM+ukp/m/tTtC3aiC1VdkFrdu6+fpapkZIb8cKo
kmCmWqIF3vlM9zcrSOg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qx+ritZx2pDvnekLOZeaFDvpDAtmg/hs096HU3U8xSeFyrj9v1CUwvI97hgO9fhp5hx7CLb4dRhp
iabDmveFs8T2afhIu9MmAO0ZqxUS0SV94sOYT5DwWoTjy8BTwRuP8Xrs/EEWKwKuWJp/Wjv7M9k+
wpkev7gSf92vj7uOWX6J6ECKwgIRjUGLc/NIrHrXqaq0yVd8j9fP6cvhVKR06OMq6U/6hMqO3Mwi
SQI1xdCXs2NXbTiCZKqVDbSBBvTJTo2cH6JXLB+E/g9NyF0e+z7oxCuyReCUVFJ21DVUfLxU3OhZ
gXG23tcqWGm/l3ZWHVqrETjEni8mwIO1yFoO4g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IXrSnaP8yioZkxR461AE2w19esRr4/fF4dA2RHFQL4fY5TpvMbkL+7RQBJ9eOLT5OFH1DsXcS+My
6KW+sTOsl2ndsfe3ttRCDI7Oeo8joeNZ8xJuwUGdOxtV0ae9PUAaVjkgDttLOomzNLph4uCXW202
bI3eFzZlGpn1iGIKiFQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iqW10+NxHcU1vbwMjaJKEOrgcrSi68eS0/IgZB3xPrIkkojO6+T2kz9ISwjr3CN6PcPo+hXCdZn3
Q3TnU/fMPFYF96Bkmhtr7AtYZE8GinVZHXJyKmm5x7dcsR8FyNv3nSOE/XYU/dyZhfnBj9H8LA1H
EJZm8T3/SQk6AB6tpXwh7kVAfE+bMsPCp98Fijzd/ynv1FX6O6GWv4CZpIVUKm7Fr8lIGCex7lCq
foNktfSIPTqF27RC3UxvVuy2VPf0Ck+rGl7pVu7l375TxqfmSlC5QxbXyTQ1NByeHr2LVJZwC+Xp
5uMCktl5vyr3uh4gEJyZSJlJ7E+uSrhstePVYg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37424)
`protect data_block
6ym4Y/M0ht8QlQcNG6PCRphIFanGOaY8meT2vMf8/pWYYONpNOqKn1zvWPS/GlBi3EbybXlkFdir
IuJyXc+W57LofPIoHlBWCoAvkqbqP0MLdZun3n4xny2eheFBMz6qbWNHkXeCuh152sYeHsG5/Y0d
z1ENGlL84EWpPPQ5vMJpp6JUdMojIiIzGcvXJDVqYb+vIkME7b7bfp6zap9xxNyR4i+HnybgfWuo
tOht5H8Mey6hQk2Kega/hMIGWZimj4FJ7iJLkNLFDzrUJfIYggZhzCo1dFiAosFqEqMIdRu/qT9S
TTVrqiprAYex9z2lY2aOfVhxgnfclk8WwmXDhQSzTmbcl2uMCWfHp6BCFRpKV3QlYTx7+r0mRgjQ
sSmAAqSuaCNmyUtp9EtTv5B+6Np3w0M4yayFrIqZ7Huw8MyIiNrLLzXM3LMJVJoFXPawDU3aoW1o
aNfVo+bDhTmGfD/P647sbDTaeYFsOJwHRi5sCOMo0YrayF4DE3i/QfD6yka7TayO6xXHal0Y83j5
bbKGsYQme9W0Vz3jv+ATEGDj1k8r2Bgzj84WBn7oYF7Q2sI0na9kNmE9/sGO3syi/GO4YMllxCki
CPJOvmqReF11AumML0hA1aBwvLS2JIw3J8BfMGybDOPoaPU36bwqOeB4UTmYoct0rybBiCZ5R3Fw
z8JDQYujjwyb9DF8+Y2gquBBsJS3o4H0NUgzhFiefF1NE8Puya6YrlNsS4ApeGPU54X5FxxcMj5C
pZ6ooGNuJk28j0KHOwADa6nyuLGKwIEsg9auOk3XmpuMKb4y+gsXehBGuAqqEX4LExR/H3cuZirL
1ZciFn1jSn+fwpe76lXCEIrZRUEmDMggVUXpWr3XDZ5SmpvWrEtIlbkv+/RfdK7DUbIypTaYlGRq
8gIi6MxtWXM2Vjz60G/Gbt//XtAetDVlizbGvhDJw5S0NqHMOumeW7f0Yey4Jm3o3s24h2cE8W63
Dw3RJ/W5wd+plwR2VlIWxEH3afZoXKSIhlpqK/89Dx8m+o8vSMYfNmXgLNKuMWThBukuquRy/D8H
hQ08/lPBx6vENPhW4jGCdPds4sjgBRTO+INoGyOYkFcYDay2MkSoJnX5RTZwRkLZqD75OPl3ppEW
BuzSnGcnIGEQlDcc0oirN14eC1C71y90/3bCvyrB23z/hsCa6bHgGG5N2QiI86+yV+MLPxSv0e4o
z4CIv5lGIW85T2B/ODN+heM4J1vSnUe1eC0Od8nvV975dzvREqygE7K+4r0cssGa8yOB2Jv08jzc
bUz9Lg/gy+u+qvXDDYy1Q/G/sAUUvZHoZQSBOFBymWzG6w6GQs0ymje0ixRMWaIZ+av+q1aK1y2q
CwtP8iy4XJ3T+beB7rbb3VRNwv6Fe5I8snke1QZI8G2vNop4cuHet/zkElFcOkRe7C6dLZ2adtS7
Q+76mR/5wgt7fPOGyQbv4vni3/hbUUCsfbMK3qnvjR09qhoncp24MNHhGIfpwhgDT7pl7eXxuCe4
hb/Y5mnUAJ3SuYmySuEk3Nx9gYtaiqxizVBLfEqIt7BptRJ/Q3yNFiTFkY8SVSKkUTgLdhwM6+z9
dOAMrEaJo92vQtoCe/inpd8pBNdyv6rBmJH9xd78ehjCOttgtdK/+6RZwqWwnM00NV8WmV6tvHLS
hhUwkv5XP6wUdDUbi2BfOl3jr1aqrksE7HNax1RWl4kGHtKLZp+lWNCLGOVZhDtn3VdjySRACcZ6
W3YguCKcPiTq+++lGFKiRvYLQs7fLbExtC4aFOzRWrRChJHp9kfCgEt5Oq6LXV603uTsCWW3vbwv
/tG2r6R7bYY3v+ZVzckOM7pqoQLJtY7lDX91AT/FOfFHnM0qI/VcyesfZ8pmiiFZW8Nh+wZesiMS
eeJBLjILAfTl/QMSUQpIU26Id6YfHvnWITVjyxrnkcSQK5DenUPryWEV7VMCsg28Sv8C1RvuoFN7
KFd/3dFsGEUQjKDsZreQHItO/zopecvvEdr7Z6TDUEaSnPFeRE39U/llFFWACJqk7uPCKA2OgrkY
l22wCJgxLcUAUjzykbzKJuQcHjYfIToTUZKrSb5YmZLiZEzEJhaza/NeueGroQFV49moKscKjy1r
iNsvbkgE++kWFOJehhzy5M41Cy+6ggQ/NCB8KW90B4L8q9sOhxRRLFTlrLBKCXZkURJDaDhXuV/c
MkBLnFXs4u9pxiDGgeyqkTlhwOuJZnhgTGl4rx/+a3gFIkqiqDqVvlkSxjFDKGQGWpjO8hGoXIGj
+4vT0y58de/J2W5/0qja0zNsrP50Ewa6muRIsKr2Mn0gZGu3954lSY3HJ7GvTvF/12JNFbo9FRU3
m3VJHi0GaF/aTXBjM260VDIzf6dnK8IabJkkhDKxJDDm7vij5GeDcUMdOCYYa9of97FPzf7kuXoS
Jh+7SJJnO8wGkvBYJrldgsh701fySWCQMFYmQpzVxzPu6FLICjJMScxr+AmHyuHcymW1TbrZpURL
oHySUW3oZCGMgzO/NmjZuD+6Itq/UM/ykOGsZfqQJUg5h8bSd6DVwTh/w6DBLe1jsxlopkbr2tzP
19h2tplSye/D3GNeHgiV5/7Yh7D31ONSB51Skdvf6bjPDeecaa8p8g+UXIAIe04t1EKswU++6MLH
WrlcYfkE24mOg3qBnQX3ZemojIB2v0yJET1sFtydXNvCGwij/xl7Ti/VItyio/i/EDF8fsi1rynQ
pVwzF97I8vzUMe0Z557vTaf4QGEvs0jlFmyXozsvkBm9S8pG1EUPm3gMu3FLK34WOPg6x1Oc7TGQ
kTY4wrVNvOhOCVoQCryj9DnOBdB2Ggm0f7vDW2/n9LID1p+j7YJJ1hJUqEr7U4E09bj+4Ddi5k6U
j8Li8XyiLm7xnErJ9yaM3nXR5BJbAMDskOc4PjktNx9fQKIyTMYmL9uHrnPqmPaBJqSWgzv5Ge2Z
SA8YvrXPX3VbO4qt/V9E/0fYuXCOMxvuJzTwl8JL2lu8O7FXWXhd4zuqfZ5i5Z9FCH98vam5kxg3
yi9HPOFGkYNNGoEkdnToOdQv/8upQLsoOJhqAYozgDR11aFp1P1XiBeVc2vcREMAURj8ZKbZ2asQ
3N9j3WfkQEWaoCY1PhmhRKgZpBeStVNwffgbD4v62sjLZg8lhgYU5KeULb3OZ7buwWBWaoLhOcOP
LFREOydniP6SK31DFiAjuwCMa/s5RSpPJJH85PdIy9qBIFDtSo6I00dyFF0RHtl2XJaHvu93cHMu
1row2c2TZoNGqvtsVL2DMEYvFBtlK4vRI5z4b2aXb7x3UrjaTB7j92yWAm31ScKolkfKyon+kVmL
szqxfKZOAoph1xaSXyYegmlGV9fI/wsmlg87AA1ELGfdUNblkqxD+zJy6DJoOov80uN4F1Wf2xFO
kkUF2AVqafJqnvBewIAsqXKYTkjH4NCcl7++iNvxW8mMOqZk60WXlijdtjs7qhJwRu0Ah2iDYQAA
5bYxk/0iV8to0eRaE1h7YMZ50iOmbpdrFuniqLyiZg9mPaw5HVPuzM5hnoV/6Ry8Grv/GXfUuawe
+4V4mOPHSE9w3Mv5MBesVGrv8Ay2/bOaPHk3rZAcd6iLRxqslfdc3j6Ima9OSVsbmQa2gWtN1vuA
xHgW2F3w0b0KO8cWrme3+KiPiWLn74DG46Pv0lJfa1srQvTkuwnQvAla1gZz/J3+0lLPCnQ7WT0e
x9lVKPPc2tTiRu9nCq5QwiUqBXjG6Xli2mMURPLRxjBSQJVVyvQ7YgpnCvoFA+DBBl1Kfpsrn1F8
LMQQLTOnyS5/Ied8IagEKjPMzGo9w8Jn7Pbc9gR3UwRX16KR37r7AXZWCCXEFSIZPos1hhRyDfVd
fJwE3dyRqy4uxDx7JIq/e8CttwbzWKaMocGphWArg+5X+H/WmdInkgsyyEbXvKw5CE/FRTKpKjF9
OGwu4/U/K6zp3B8fccA6M0OvXoX/pH5OjLrHavuDAS4NqeJbyCCMCkynVa1V2e/MpYVXlka1KnrT
6onmsTIKsDw410TnV58oTmz4UYWiesWHlAOKgsGWo41UhwltPs++WTS+fkZ4ovlRBORmYRJg8Rok
IT+fH/W/JxYSDwbO6Q3uib1SgBsmZ8uzJ+848m+gzE7FqyuphX0ry88PWAck79BnkQ8Jjt3UUxbO
Pfy31YOj+C5lChUK3uVsoXA28CAab5l8NOwmGpyHThjzL8dfHZVK5OV1l72Vgts+5jXjgRylZw3C
DJoCDwybgW+XVUvrn9zccsnha22v2O5nNCskthu98ncpfMCzoXc/dPBe0/qBusfKv47/No99ARHm
PNF/RDVZzB96yrrz1i/95BlqUOw96Vq7v66glmwqUVZDI76h5MzTJpV45SgBLZMyyCjBJPRdnGyO
kfYbkVpnK9CMOE7vhAdeIAABH32a5XNXlp5Pketc4v+p0oazFbhQt27kX42hQowQI8DlfGuN+lnJ
dVuk1dJuLzus4aboTK6fxfMVLAyRJjafvs1DaFkHRGhOUjy0b+YOwR/VY5/LDjjZSw1XHmRponh9
r4mjUwnSJ9EWTJBMET/zWK+5+kB/YvY0Egg+JTA6NPQ23bRTdYuiuWuO1/ouuOAA8mX+GqBi+jiQ
r4e2DcINsVgtTFAtRzbbQDQmHTcGaQ63KZtu+2qjcZ0NWST39cyo10j7ziEoEkl08M/fYOZnPRrR
xRKYumgu0nlnR3Lbj2pDOw06GkQMG/YMejfagjShUumM7yhnSefMx2Gp1Rr3dutRj7Sjkl9VkW82
iceI062OMB0u9UIHPijpkrUa6xnt0zuuKQFplb9TGP4R4lQutk2yDv+M35u4mYze2g1Tma0Vqosx
pvtSWGpXgFzocWe9ukgjG9M9VXW/y6HBerBKkQM9ktGKnokOtVbEfTJHTPJFRZTRSY4rBVAtUm+4
jYraN698S4bwS/2elZW5suFInimiWKcEXEuK+EwRbsyUaoyXfmvM9ytoBeVth25gBcFS+1ilCVWx
gImbaiWkyKo8R2QbkkMRzQcIgC4VHtm2mGLeFt/PNVJ0B1CwWtmBaT6MW3+S8KYZWLNxQ3B3/jns
pXvoCb4fJLW+7s0J4+6aa8q94rsav2eUP5m3avr20we2t1rlMmr/DUdMCxpQA3/sZgsFx7QbA4+f
Q7s9QNy+jdzk/5m7Ez14rFeQp2uyDbqHpRTY0UlNi5AKk71igjeN4ghomp39A+IUDXyqCdldjzE7
X9jBFK8XjWRxoPgWfjC0IpxDHNfQuIvgenVSY/ywz2miA4iSYnYlGMICXYLTzjRbbex0Nmaj9g47
0p406mG73hHU/6qh3vVsMn1tK0Gsop0Ntgeo+lSl3pZdzCl0uwft6tbxMCtlMgWLQdLPibzdwsF4
asUTadzqoI3TExLFQ2JdAfC8p1T0HHiPXuvtoA/zPmLrBvz3XseZkZY6sGYHNoWE8tSa9dRyb7tL
+r3TZLpddxRsb5G9pcJ8TU1+taNRK+4/wJXP/P37K1iNP1NbITR1rQ/LbmvlvMa5Y8J0r4YxJkt2
eom7z6ltLt3Y6h1qRlw2J96BWfAD+41OqwHSA8TodTdnGHf9NRhynLjN7oywSvq2YFGlHCcRpS4a
q+Ccd23RqBJtzBbmbEeGqpVyYYK4h4Hr1TKE/HdmN91FeEMbLDj7om+8H8SCSbS8Nu5SEBm7UOfZ
9y2TRNa+TR6VxJdwogn0v50VbQNosrrMWbI1bOI//SCg9DHB7+FmslCT5JNWqRP7BZcjusqAnphB
hknNYHmQTbmp1MoKkMj5ta3AejXqvn1hwLzaf8trOjBvWD1kx0C02Ic6puMPVCiZNn+z+KX/jfIv
GFMlNSA/isw6qDASbKdVvYwZHMmu2ZxZnx7ZKCEbogx5wkALYi7BRJkGLGWt/lVW9U0FHx90vU4+
jSnoocsVbUrs+X9An8mghPjGzDzLgbaJJ0JdmDsWSeggbLLXl+LV0okP8OZMUq+yu1/cIRqD87tA
DfxczWxUofFxPQX+3eiYZp9LMd7f3VcD7z/yAMWxicdgKh7Q/vbTD/So28bUbskHGGNYiWDMKlQY
pvRePqlFm4mkwE964FeiTkoZ1uljN/yGPYg16xaH+bt7nOoVRqSNkbqfcP9ApRkxuqQQz1CI7uKi
QWnuofy5/quZZPwQXXXQXLgUp2321OO8rwXdRWdOsf/U6bOM6JyXINciQ8kR0L8eqkYncc4KJ7RM
HIBAlF4OknDDbBiDcBDM6hukm3MmY0vzQFonId49KXeizY7YWCn7OEufkpIzj1Uqs7NGXQ8DqqdL
UoYd0fuJwnxRZ7K/vwJQTIR+k0gQ7KYGVG8ZG2u3mZQO5k3bOgFUMknbOzPKV49sdDqAXKjwtD2m
v1ORgfTs9mtzt/LHwwCuQZFfUorFdgLB2VMhNs6Asm4mPMzKlm7QoMg4DSzQRgtSfcgDIfxo+x9B
ymO00Y7wR82OXgHCYKgSU/aDWXXCJ2CPen9TDPFl3om/2a7s1rN3VSJ5XHIJCqMk4mq8uKSe8VqY
MbnzHwrWmIeLxqw6LwD8PvnXfaELQ9gPR/I9uCAXx6oxPZj7d4GCFOkdNsQO7+t0xgfBmttQGNNR
89r1O7wgozSWHIUS/5GUm6K1MzTh2h40yEx57z5aqvi3oxgUZcc972+9C0M8X/mSh33p1c1OU7/n
dXeDSK6YAosojaGbdn0qbwboV2LECE7/+bs6apq4JCwWVPOzjtZqxg2DTJApiZOReMOTf/fVpeQE
Axl1d5g/Mg6QwISgBM15QAzm3N8pXxkjDRs/k5xBc6Mq16OX7+XqxUokOj/+/A0HUckVm27jextU
Pmjy7U5HvYVzGZRa7YhDwB/OPOV9Z01S8wwswoeO65DfakQpIPHqpSEIWwibnJgrk1B+lAgq21gO
vDf7DlF4vxjG2abuL8l0LOdXoWL09TRm+8js1k5pLHf4ibb16nZgtzkxYqt8t9p/krvxcwulM01V
d/UnBLVeeBEMzTBGCim/pYfb052MPsNoIcKpdojT0XB7L1gt3ffpJTJY7DJ39shHKbFAu7buKe4C
+0Z5Nn3yIpoy/SgZpnRHLRNYkXBxAf8ChN5j+x+N2cGjK0hxa4+dAIBAY4Dc2NuxrWRA+UA5WR2j
UldtvdjHDg6LEh3J9qGWvniQTHJI2pG1OLPUTF/KXYixNBq3myfJ2WTYOkspiHoVz4ta7X2TByKM
ehrlIIAVv77uTlJZQekiRTQxuA4zUSy9Wbp2+2pRIOySBsujf072GycKTgPGKG1iWc02xWpr8YSG
ZaoEIa7Dk7Rkr6qkuQ/YQuQNXha2xQrsLiz3Cuahw1Ukl47RXPzccuzRrcS4xSjmow65TsTNqw7y
QNYT9XtLiAHANcNu1iFMQlUp9tBZF0WnaO7tcf9TrWCojrxp+DiLMjTsjEZ1AXKzAIy59154+OSu
kYNPYE62glRQDtZZ9W//htZU55ZFJPdgoxVEWY+Go8a+1W9QPmRBXD5TCAveGUvzuuQ6vZUJcwih
zWYkJbZkXNhxDJR6ZW2CncN0/3ArbKtG0vCijevM5Tt4J9bGjizRJ+Uglv5u+1/DLhLrZCNtY3FF
U+Tm553YB1RkBC7vaWs1DetbUMiYKvbvSOc+GXBpxC8l0l1eHEm3YN9Me/pYDiZ6Qj0tex36FbHr
SDq19stEL2NgWz7Bz/SALqlEXah0qyk1FRxpBEiJ3GEoz6fFA+mYEjzzMh7hjkBPfFs6+yK/Ey2I
GmAI0mCTe4ghpCdEoLYkXmXFmHInwd2wJ9rkUIG0T/p/vTr2Lqu5/GO34pMmEuaNCLqyhXwFlZK/
ecGpq9zUAt/2p+l4QLjNvrJtfRgDOTTGw4EQhEa0/jNjHW2PCgTJpKl3piXFy05yBqzoJ6o4ZjH5
THVI1Zc7e1azP4m6duhlzD/5w4jY+dvKWJZWUylcdhzNmVXN2hGPqgbxx6QQeZnu6+lk4yFdI+n+
v+dQMQ7j0B6sP/gs3OvyFcBo03TYDEBQ+tqPhJBN6ijrrgfUaGBl4yxmEx20Pcb7k3kAP+Cay27k
bUmQ5Yr933r3IyWSJqq/42m6qzGQxLVhefnIk1WOdXWz5nxLIzf4c0fmL+oc4X/3q40176CKLmbb
q+skJNUEKFgH5YnnD200xjHun4UlFaZ9J3XxXoau9A5fLj7emlKBnbKSesCzXLrhZcaJtnmfSdF2
riN093vIUNKTSe0OyOlb0SJt0zmrVT+cco6nVS9BqXGAOY+qCC+PNN7VI/PsKrzjc1kGKgP+3/Vx
fHyZ3PEo8gwm5Z9nFFwjcgMaF2vY9KJ9/WHWtAuF6j1reVEpy+7yOT/qTjXDEE4GF70s17lMRgzN
IK1QdG7tnf5Jqlx295trUEZmascFNCQisOtW3AeezQ8Wne3aq5PYoaUqlKr0ehEKT1OM85ef9gyl
7wh7H7YxYKTMA23PaUsGlm1QgAH2VGq8YT719WsvYOmp9z3lB807Bqtcyxp9zSq3IQuV8g/hKX7W
Xv8gOgzrRj9Cu8wjzqKvWovoNSVas38lJeZQsxHhwzC7uv2u+Zr4hBPSoNzgQOYMNmEPp7oJ4QMU
4uvTPkg8jEDK8ddzaq1iAADgdkthL3i+KIEi2Hc8Z9okduOYU3VHrH1O6LIioXmeytpnKP4tmtXt
uhJUiqBGjJdsppT1rL5rmhMypKlN/ebvjBNsuTkQNR9ANKB0yZWG9e6zVIcXrRx2GM+gTp2208uz
NBEcCVq4SyAeXegJ991P5cOJ16mu1atY7X1qyJjD3GcXPWTZG67AWi3QP4rgZiJwsyLF5A9ZOOKn
p5QgNs0G0bjSLtAtE1PLvPwghD1XaOBw2wNKiuLgeUIsE3Pd8TW66WHlhM2coo3jbgNqquCU7ycb
KizhxY3u4y7S0Y0b2e+8Fw/s+jpCVCeqDEAuKkbgWbCYCmsGPys+MB1VdiKH1TBJDfnfNglCUrfi
lCd8tlZD4uUDcaGIsEG8OtbHfQhrexOLjKG2G9GN+ryfrKjb3qw8vddV3WKDKt9FTbBtNv53BOOs
tgL8bIiFGh0FCGaZwKNUhcGA520n24ZaKLYv3Dsu8oOiCbXATjFUcnTJB1YvO1ja6OhBoidnCUHS
Jr4S8es6s7HXTqc7daQIchjMt++gUPFuZK6CGUXAr0Pc3OwrArCiqiG15gIE44p8dh7aIY9347D5
5hOY9T0z749hTYYz+xsYTesM6dV3NESq9r88pz9GSuGILgvOaVqGKSOPJW0EFAsHLOyqwBkMgb9y
0WDHjeixJPjyj8b/VhCQBUJVB37b4SQ2mvQ1V9TsjhrbV5shfcGAWDEx9QrFL/7NgTLhTftLdqCt
qSdJxC+mKv4TTQO2MCufDqDH+1a0aUyutFj3mirkZKHvPxKOKEmGgt8afwgKtLdQxumAxb5Eo78Y
1pj4POj8J+n8P4DJYaIq5dptEhV2yWYQmTnb5bwL8roPKHDS1shPyGHQ8/RYH1yXKUR4uPAq7UvO
tl5V1PicOMpkwr5TFuvMXAlEAKhE8z0HK/895ETrwSgIkMZMVNAgYqidaiBCNIvp7IMQqke/eUzE
dz/Pzlx+EmscM7CFWiKkxL1f7EUjFllLLECtcWYiXVK3RniVf4NagpoaRV3skZbEMbLhIEw1gZ3n
5dF5LAvvuZxVfi4KsLiOJdWx/bxR04OC+q9t1AZJ9Yhg6VD+IkWhrmo3WIIihUgvnbDu4PfpPkfx
rasx5/YmTfIhNOD4B2YWrkpEIOWPwb8QVLJvr3TVYO3R1HoBC3Lpdaepr8aXVC4Lx9/g366krTWs
6JzD4ssxEF+8ZoTcyqr323duoN1JyIcWAk9iWfSRnswKRJVb2bc8kBf8RfZCWIHBtKq1tYr+C7ss
+8aJ+LDMN+TMtFETxclkOQJd2SfWiTXv0uCTpM6TcBqhf8zVzAsP8V12gHKGidrhBmeeCAw2O2ZC
2lvb6/AQE3NIf5LtQTRwjJLGdIKQ6TdEEFcOnWxuAWmQTt3WfZxOrwyHZugjQ5KHFzQNIlGUBJEi
L2M6Ai/1ngh00PD4ToFgy+YzBK0cth9CLOHRmHZ/xc1gEpSEblM4KJGlWeNkEB4kP7IJD6lOAsGR
G8OfuNWCeMi37yrqsBAQLEl44GqQZLTy68uUctVmMAGtAOlTsCr67BMMkBv20pwZ3o5WWjNkjZNR
nv9nTJVFjtIT+hKY+R5aDjEGbJzvpXHiUSzR9/759pryMutjJNeQhTJuL+5JZ4FDEHZOkI8UDaXa
gThhdkOIbiDJAkZCQs3ccbYsTKmhRsKt0KKLKIpyDGN3DglGpRUMFfomhHQpcJw35okwC3Qg+54f
fFc+YmrAkrabUmwScuJBD7XqZgTbJGrfZ3iy+YKj7ee5pirbax2GCimJ7e+W9e0Il0ddheVn1rjJ
kTsTOHQHQmj3U3ZUD6EyM8qHJru2sc8pp6wf652e3ieY8xjUF7L11Qx8TIwj1+8I9DPAC6LV/Mjy
pgiiNqJYjQCq1V9AcRqe0QH9qiZfPykjH2Kb9fdLZNFx6vkhTO+xJPwHKC9BkUV+zEGXNbzzthY2
RR5qwKh9xy+VZj1GJyJTmKSlGTrdeM3LfXW0Nmo6slsgRsinYJJz1dzjYKfyDP1sSplZLqThjtsX
AmTyRlRGar13lQjiEbBeFdc0JnmU4HSyuqkM1F2LZHxIiL9j70NjiHbW6kZ6lyfgr6Bcc3O+joN9
5tIK6am0XBlKIOewwceCzzBuhKa1I5xH/B/twfIubF8AiIe2w4Y3lGWsuMPxnnX3Mhy/tFiRKDR4
3hLmR4KcjtuBraYIranXyqpkPvbYeYwRuRank/zNlI9oIXpD4jZQ4Dfva5m29P0Tat1CGTh/HPRJ
XehYwW/XT3Am7GJX7f9GHXpzd1KB7E7btP9CKZqtslde0GbhDm0sRjLP71aMw1sl4l497HZgQC6a
0Fb8aFktavrT89+rHreRLxN27EK0RRDibNRR89mMp0+j9v+naeD4qR/wVYnfr3hYXs3vwSvLTKEt
fN81hqsz3WCpSoD3XE5HtUYuJ8A3YLs8CSHlKanYj31w/BSKg488x3wpSL0YmF5ScRZQia1aNZ9n
THj9ijYTGQvXF1CiwsT1OfkeG821NV6jsYyb7aVS469/rxFsjxgwwEc4hqAnolj+FHRG3ZMDBdN/
2SGN30iwqWR7rUTTRkayfAvhwW1zr3XNDO3MiZ0Qm++gpeeUrkdwGnB3dHAvp1RmBeZqkkhvnJu4
j+55iJP0ITKPQcGChz3gbHrer9e21JYDzOfG3C9u8T1COqFU10RewEFw0HA/+lOYyr3mjRmy8iAF
ET9qEX/RCaeFNhbh8BoqZmMuqFKF/DppIQOPaz7cce1woOhAgtBvUFjnY4V7JBV3A+TiJTogVkL/
1+QIHkYzeTWvQprcPOh4/tTA09tSjNCaCTTa3XYLoOjGqZZhCgoQbU+c76SwojnlfENIjMS5y+Zj
/pv+NUmPxwKzkqIiiJReFRZA3p9OYnb6T8s3SVT35wEq1d//ndBDCLBsgpE6Rl2eNhBfcgb02rIu
Ljz5hi60fTbqMamqg7vqJ0y+3IBtukU3Cn5ddQJgLbAOnTCNZbvjfj9pFY3WSp1Z7kfy2kywEvMv
nuC4SR+L4l+BbiT4q8EN4HIp71GpwkXAH//2dcUdI5LzPWB9afcn4NQ74zsotSrjQWTAQ2zH5gNw
gJHZnI6CSWZXLtsmJnzPIwu12wvNp/mx/DnlJbUf16Xg2TSzj8iCJ3eOqxf3XDnEfUk30B77DHHV
KZDGwDrApPeofNpBHRDH+B+WIkSBL8r1YPUI/i1QPTWC5WhIILlWkch1AI1mV+f64GBXIh0AwEUl
ZoehHP8DZ38O0wkG+/OiOI61lVROVj/+mtGXufdwHCsg7m8+THfYGKF6VZbD4qjaHd89034vJqrf
gEB8p+nCrYeGnqjHR2orZLsAI+YoAUaBUBaLtDqLffA7T1CQlOCOlLywa3M+g3TrK+A9BFuoPjil
xK7u12m/CX2rwTSShEKG0swlWSi0XjSZcNPhQpJKtOF3BsbuDU3oolyCSzVjjWEIVdgtxTFV6jtX
9judCN0YZWPvqL/JPZOYjkPbSK2gnUaAFwgr5hE+PKpztb4j4nkvZaghiNDeWb9kID+kKliLH40k
eZw1KF0Qc9CNUiLEwD4J2qmQLlM6DseUTZD3Su73nkw4UeFyXocEDYZJcvyPHONwx3PJ3iOO3ZNv
0huR/evomvRHmyMeqpG4m9ak44iIKD+SEO0L9N22lu4Ae1zNUWUdDS1t0PNn9QNfXn5XH+YO5Bp5
2VncO4bWAYXUFy8uYy0NWwjGh1kY3CDKoEa1O7kBzQ9mcfpHdL0a8xf2hBrRDhFna820oemsI0g7
68RIZsDwOvvxiXMYBz4ZCzfln7FOH33pF65RUgy3KNzQLznbytwj+m67ne35JydLiNdEOANWx98Y
GVyH+qO/7+/jX4z0m1baDtF99QABWZRG8GQv4wrsmxM8ZuzFrfMo51NkTMso3am0jZZYOoqhbOYB
SXbioBiaVmy9ZY/aufgX5xhO/meb/aW8FaoZtkAjZK9yLS4RJhnqceRyRigWPmMfePgv9TV1Ahf/
uj8sqbkqvBlYqybpOSw5l3DJ8mKLnXiMskPN4EvqzlEpb9ItEJnaKML3qLEROqExHC2zb6D+PaGg
3sXpmQN4lw5zky4VxgFNwQVmafm6Fc3HBfZsBjYi5RX9tVSeS6uAZr43KYcUVcaD5YmdlQEnz44g
02o0d+kColdypKCTJyX7VW6iObZ9Bw/kTTO2mfSinbXlXv3fO1x1fjwM0ECYrHTBo9ZLkm/vfdy2
Rdxwh61mcUVtZ2utOBn9z5wj2z5UjPcoDNM0WiMHfq1Dp9g/UD+AZlskrGoZbMo5mjyR+OOgDhNi
opyxhS0UHE18FlwVxZ1JPAfgtT4lfYfe6KacLi7WtzQuDMOIfdQ05NWG5QLoobqgieiLTeWWs1KV
fMJwGGICU8ftyPm3Vckf5dcEfKSThpTt1ab0R72K5RBZThVoyuFUjWnV1yiURqJMTk2/soSEAlFr
ukPpx96X7Wz0P2IJhnrbAnzCElzsn9j0RpAKke9Ygb7Uvfw0RKR9uFNSwpxrWX00OkY2MhZTV9tJ
AnSNixn1vzWPdoGd25Uj8+aE+K7kricGqOnCKvQVfW/RCj4bhcH4SSABZtGGCIZUyrKA25c6dl94
EZ7ARmjtg2VZHp84AYdlf4vpPtP1EES/eXjPTb1r4nikdqQ5oNYEWJClgUom+k0IdJfvIoak6YFF
ffiDoid1595OT+JPKZyF47LL3RnzHT0P8wucSph1Q34Fy3cDxivdiMD2rV/72osWOCkszNiJFClj
MhKXc5N15zyz9NYyO/umJlEdDNhwZ+8yI4IcremyvHCGCbshChgLcuEC+3WYTDrVE/XZk54Yf+VC
DqxEpcYZfLfG0pjXz1Yzn7X3vboQ4zUMwetIIMlk5amFwn01O+nL6tdUlG9G8Lg59DBYL6qjoonT
3OUU9x3y1pCmZQzjUwAc0CLDpmEnA9Q0ezhaBfvd1tHDJVY560k+rLPDDj7Ywf3JHMtKGpv3LDe9
XfxKu0x8IiZPzu36Q0B3LahgpJpatBCVcfD5Iqbbmlu/eBSoBrNps+Iatl8WmVn9rTS23MOVvycn
6wFESbcmAhbXwpdbJckQv2+psNGHHwonX2kU3WsX1TRDvmXrdIpH1fz7/4pXe2K7RQbKfNzo0UjR
/kUAjrlLJW8X+fl0FK18usQGVN1bLVqqAPDaCIzq7VgAwfI7FQ8Tu5C1uMT5Ngk2iZxPg3Y30RwJ
NzJfLf8oA1DzAMbzM3lji5aDRY2Rllo9yJwbpRop06bakvefEF21USBV4zTW7wJyuADZJdN75dCG
eF9b0JxH/xJDVK34AbcONBmx9Ao7FiPblbYCtTK8B/c65OYh8+iEjBGrTvFDZMoKSlGrF2i1UVaa
72+WSU+DhUY4zwT/JML9mH5OVnMS63K7WvXWwjd1R2TvQrwPPGVYlXcLkRFSes7GRSOsK73pTAzi
CCiIWDZ+aIWCQOzAYYrQcIbiLG9VNUlXnfkh8gHP6w8STo2rIiv+oLmNU/ATk5pPWdUwv9vjo5ZG
+ZfZf+AXo2Fh5xG5rIi2w/sflximQCuR7AbNT34nM5T9PQWgp1rqyQMuzSkg9sWQQdoXUK+9ZSP1
vb3kfMPT41n8zuWZwOQrIvgsH1tYeD+Ob6LtePivH0/gw7Wb3S3S29IsYvwDnHxgGCWQ3j8dIVFM
vPr9ZZCg2cSfE7BJL/6G5UGKDO5GHJaRdev13oJgTGXXVafnDfKtwZVb19HqXXWWlisBw+CA2ja0
ioGjqOz4ik+zzIZYnE2vEYOm0mysP/L+CgJZkTW1yEVfJZ9LMiO5Mf2ZrLSSdR08uLKkxRj+FUVz
4J6lJHo6Qlq23eh/LMIIYG9fjX2kYJmhqB9VxMsbldpstTeAQkSQv3uzTUYopmIaGPvXFaQ650Gs
VMy3vJss6VQnK+l5+kRtYUbU1/fwJvrHMhFoP4Qy8cOeqKdzRXu5YRDOmNYHcn1xrUiTJ/3S1rw2
NL6M+qTC/TJrpJojO2dxBQd4l5N7IYHGTW5kD6yi2qCBBdQLRMQzsKzMKT2irKI+soXz9Vt9mtpu
6uh/z4cCZfzAZhuJ5T/IgUKD2unuWeJ75wYjaZ4a2r/WnHZMPRmG4B4N+az+/Fr6NbLT8ckOy7gX
v6Wq5xZtUHNonPSnJxdA1FE1TUVdaug3PEvuPbKDXzvH45517H0qFKPQ3xkxapwHego60QlryX9A
Rq4nbpMQoeV2v38c/mSUo9u/236cNQw/3MMJSfZC3v6JEmrTvj7wy9FNRBt9NPLIpZPBlfQ8h39j
WGKkzNY3MeHU5nr/b9pyGbbD4sQypj9eXGWu7QxykGSEjya9mEx7Rq9GEkCopP4LohyR/kcEuYWg
az5TmL3Xsl1cmObsTnRG5fQ2Jfa6y3QLbv035uh9s5JhiWSo1LZocNuPMca7bGc4ecMuLioAwR95
+oqMbDc8nQHvQV1Zw7ite/K9+2ANwQ5mGlWgbU4eysil4bWO+gy3TVgEjhsL54F6RlQXaCNX8HNJ
ZbcfPUuIXCNZbcrwdFM6s+S69+ce9uomsr4gkpeIogIqR0yk0Fnid4jiv+URW5bf6GKZYmRNtD78
9GUq36QDs4dqdXjVnmyjDY35A9lQdxLG7vXeCzAFYK3pOWGR+gIutLx4xp7AcFqTmDBU7g4dPwZQ
rYQTnz6u4j3U5mATm3bBZ3QqRTtNUPTRrezRqZrmro5V3RA6HheYP2SHeaIkejol0xWM5+v+dp4a
/pHghvt1kqUN54cCVpbKsFlSwoBR8gPStpS+yAa0bWizAbmTjAnqMnzE0vfvmup/JjuxgxgGMQBf
X5cAma6pXAOp1OG9XqCrPTQqBytn1E3D1JYz/wOJwbDnVYMscycEMVsJKEx4210JRj0Dw4NV2643
n/PwgiQK1fhCPxAQNr+tgPkt66EeDR2+kG5GiB4N7j9oC3+4WK/I4UY3yiPT8EP48keHYVnrHveD
CHiVDeQlWZBh+SPTim4NScRg7nzYV1M6vFQZMicIxCBhS0iz7U9/Df2lCC0JuyMSuYWBEiC0X71l
EpNDpyMfpo2pb1KwK1d12ftV68/CVZmPoHRHo+lMbvwVg9eLPmREN2UhXOhuFMpeqIS6a8mtAiha
cRNLdvQWr0dXL4nw2uEa80xA6b0qnF7XH0/oG+tDJxTF81AaHeSOG8ojz2D+7n7AQMk8weYSQnNx
cP1lf74D+/ReCqHpJbIOh9wGRHHCuPlhY2/lmYUcrOEGdq924rArVWdVR17sOmotqWkFu6dYiD9f
QtXhbm4A4KvHKwABQU/OuX76ZLN2RELv9pai2bhzqbyE/pGczTDhwUeYGHE89hsx+GjOcpSoRSYZ
FgopRMsyISiIgY9krHbRERGgV3ePV718knr+HkrfzYGqTa1NYshPHPxO49UVjN0Gbx437D4lusTF
Cz9Uyyc6duJI1okJqKPVNP836qdhXHSLy217nLnc7nF+G+jvR0sJAjpB3C/kNGuL5pQeaEhNMlS6
OBlektGoe7lpJEmo8DhODkQ6+9tddVkcEAPHHGwWW9ictr22/AcK1ncd7P6JBShA6fn59kbur5V/
R7aKOzBoDjA6MBDOTVtdjeunkvLCpSQNSSY8PGV7KlMLkpl4xlf0OAbmPTk5aU9Knl83ctLEkaJ9
R3fWq3xfPM3gbObOfUA5SD299+6RTkaSwiVkb+AJFOeDCQ6JrS8vd7jyBX1/QITZe1aEChGRJ40L
TfemkMTCrAYSTR04ThRN+UKS8KuQjVEiNXgbLHzbS0D/eyq/NQFTCF7ZfHbZU17OhERqFgRVf3u8
oZ5/s2fliJdsVuszmPLyILyNsqTm57Kb+gFKqj28r0WhTYRtzqC5v2GhBn0I03PiRtaLivy3l+SS
hwv0m0pTtmKS2Et4L12qthXPY4vKRaFRkZvR89MBsbDJourXs9lbTdDH4lApJzGdOJB6CvppEwhs
3anq7jQx/K8hWkUn4S2vbsJNFjMluMIWvcrnKOWc/voFn5IknB3LXd0F+BpDVstXAUnHbeTLWpdQ
0yF7ZEjQzILesYSq8GIYLX5wU2XzZ/91Pk2u1JxGgLiq+VZUvb0exL1Li9kIMGeqLCM3+GiFc+9M
liCmOhBR2xbDc/SHL9+3vgZDNBKWG+ytctFqqPWuLXN8s4/2izvPJHqgieny1CG0CSsCzZihcJq+
MdbG+qEx7d9OZ5YnFcbSJPrhtoDstBjnoVtjuDgaL8mBW451DfTWvzRKJ/TERUpdTr/WtFLYJ4lL
ChqZrQEQyeSxS5alh1MtPX63t1nqUBowNvGlBGo0hXNiFRKoQcOoBzx9QA4s+A8gOb5RjUVOw6gu
RbKg3fg+sZ8n9KLjNSdol7PmBvTArWr+cw9qUujvCziVKm/D6uTE74l/971gFbninV9PlBsPTOkm
Zjdbmq8PbEmqlC4bHg0LKuzdvwMk7Sa8XXuATauN2LlDhcequ428nrGg3PebKy1ybDFicI7Nq1c6
5tKK/33TBHbjYgr219iBSCH0zxO00mcTrYWZwxrc3Do3afbzIJhAAjv/FkNXPJYmmec5oYmUgRJv
RBu0QW9N+sxHWpJR5s9jf2iIR7ihdf0BOIKNfCnBDCQD52lOYWxLCV4jCPMzukzOSqel7NmRb2p5
aUwVciuhAK1pmSiOM91ayfzuT7DObOzdNmo81gTaVa7qKcYExVI+A30jji1BRzyhHV23lzv/J6V6
gEL4VKgspQefQ0TZbKJg8TIn2OmDervnXNTzXnopzCvitp5nkrmEDDyiaGnqKBjPlrHYW76oZZ3d
xnK8LToUY5TjuVThN60UbzrFOs6RP3BXjRbHUNPQl8V0qpmy4WudNPewivxPmvtQrpOHswgMRgEN
Qy0cfVANLw11LMQ+Y9OIfTzbhBzbjpCSCWFI4A7wL9SglRkrA86Ao7/dBbuxIyfr8gI/nSfKMDkl
fSCTau3xh0FSDxXS3vOl9Ijk6Ko+teX3tvJvV/UeI8vClKQKf3jHfJjcFEWnAAfqhvv0mr4wzKYt
xEalfYCKfoc8YsSfo+M/5hypZelPk3DFsB01JCql5q1wCln1bMmx0Kkzbe7wrpCpkz71fra5WPPE
a2yT8ZCfaki4PzQ/h485WSCh8T/2x7z8WdWXzOpAUw0IjieqRP+KawtroN6/gHCPkiGBehesaKDP
8dEp2X7mV3sBVOVf/77Eev/ZoI5RNZLlpry/tyqL2ZR5rANWhtyprdJI7mdu1y5G0glc1z7bUcUn
Z8H8QS7+5Dr2uuXnnQLmdYRqioGNMTSkN2vcc4VMTzpRMFIylq7p+OAH0vnj5H5pHofOrn8C9Hdg
Zy3/GTDVQnAaTLJLuEI+WEq7RLiNTXPEi0nAOgQ9NpWSUaJVpMen9CHZbwnW4togFATFHy23naAC
jfCE3Xcdxr3sO/byAIrQbPQ3j6Fvl24/ykO4dyrYFGaJ8AmY0YsIqxwShtDkDjpSoN6hrZ2eYL8p
DV4WdahmFtNpMHVeVvg34ya9UnYdC2VwrhGkkICxGlvFIDva8SxTNdFckiyJqHYpHHSU2fbZSf6u
ZZ6tkWYRWOJph1YywS8yQHmbdmzuITqROO3YpgRoQv8R02wdTXKaasDePqYbTd8mdRnj1cVmjp/+
z1ZOBT+iuLgAXnyxH2d5Ld4JvuRScHNHs8mfZxcVT7vu6RyGH12iXWaBgPyaIHPm5j5adr1U/tkN
MvIbk6dvFbH9+vWHRITUK+XagVm2ge50Y7yPjDTmdf7pHy/hyozHaQaeMS//BELdXHO2/LiJ7jAj
s3izJrG9Syt4yxIXm2uptvl0a090TmFCHgUIjH6V9s0VycAnPmG2vcHzRnEHD2PysqUE4s0TX8PK
Vpc696SDn0AJtvoqVHmeFzYdTDzJWTMDWTfV/rAmIPXhdjI1TV04x0sPVqvtqj9rf0uW6vEOyNYF
MiQ0MFg+NnHl51l47i+EwoEQI4N7iegx8G/RfWxepw96FLx7IOq07HGExUct+2ihijTuY8Q4GsIB
4ba4z8hJVrzNdcQmndNrqRkIFWqyLK9Rl3SOZdEii0EEbAK16szM31kzxShOMv4zY1kPjMWSvh/J
BPyNM2AQJ8xGIzrfEojXIIq0FHLPtae2NF8N7NoMlKDSN51NoEFq5UD+uo5JhDy1gQsPkYRUvju/
T/H5OWGR6QepzOHu9oBOB6V7iWJ/Wbj41anWb93HZRPcFvIzHsKufmWBBruhRsJMFbpqUM5YPxr+
KElV3WBOnRDWxf1ujieVGITfTKsMkIGDNV6l6rcRatEa+/0NPNC2jjvcxDFaaBjCbGR8qcZZUAdC
r0eOxvDYgCMzRpBzA2+Ea3dApaA+bnwDaHKGuc8GlnGr6m0F5xUUF7/Uh+xBoPmXok2g+lxYrlLe
pI9ZInl7C/IWR1rHQfJBEGuWVQIsabnTSq5BTnnsifFFhlJQT0f4p8AGzVCxQi1IKtfiZq+XhDdE
Yfci133tkJnuVcUMddxGJiDk7yQyO8MeJ4mO0OeDCrDFrOx5fCcUZh1td65xE+dFNIxbozxZGzLP
NiGBDRRhcIeqLFyebMItQTUO5oadsbbr4eCzyycoMlpOVXL6Ht81765rYnkIPznn8fS+JfFo7wBS
q5ifZ7KC5A4Kj4cTZo5jxmf9Frm0sD6+mVXZ8SSerso+3gvG2YOFTk/hFe93FhtyQ1P8y9idV3b2
rUMJCLNtW0cRn6zdl5+582l9KeGFiqF8q90tRNyTKMqmbTPjBquHy05qlhSqNZUEvuR6lx9+1gQz
AYhq72VQSgDJDBKo4XCYxKwTvNoctEos7X7WMAmruLsaLNmAk+0UYNra+X5Mph3BCR7z9xN8KiMs
YAtGn+JKPxWt06NyDtMY0AcPrGuFG9nDnUIcLviTlu6v5jMwagSjLis6LKw9POIoHHiwSUDm8cf3
fK8OzbeKlWQmBZQyUrOal/i9Pifu2ukCtmlEyyGaAM/RrEGGK30LW9aDs4nzIqTa1xaPDVGSnUmV
DGZ4dmBkUCqs4mv+A+oPHgh4T4gCfqnPv0I9qMNjCJjkobdSfg15RneZYuGc1C1A57K14qp3nfIQ
iZbQvNGlWH7qVb4GMJNUGcenaVlflfzcOJUTBqHMN1IB8JGAG9WNSIhnqXMraYeSAzo0gujw0Ugn
6IHZws/v7YK52wyUsZTFsALSlEfCeuADYC0cM/Ron1An2JpnhZx6LIl3LowSULfqhBROLaMWJut9
l/IemNzX61shK+sRfPiYw7v/YOL6MCEWYTxcOW/xO424L7L1LmUYyFBF4Vq8hZb6KIk27WKR3NmX
82j85+QdQmZE88Msquj2JEmOobW3RMMEF49oyNvO7os4IaQFcbp9Mu/ejj0WhptFj8AWTon27F+H
RYo1O31pAsywT7u1joOvWkC5xLnoERLDjyzgsYiU5F9/T0NCNuhEYNJHkJmMsnPBy8kfzhkjpkZw
HhQjxqpxg/eOvdx7+1u39oqzQhyiv5F+XtfJ34BnIk3sVC5JUu0kvpEwLyZzj+DFIUHL3QXyA0vk
PNRl3tRKLTZP3QwBoUusyV2iiIeZvMf6y8ZXiCSJE9LFaq92A7g2zo82tBJ4AMm64xctMI9KQrWr
gQEx3ip4YRzd3clcR5ZQCKW+9CVMXeTRcnQMVwAHug9U1n4OAARyfMjsGf7yMc7jz+0YWJDyHiAp
Q2cuabnLDEEgseKjHnWRgjRV7qbSNguA9wHapcTGC60SrbtC1DC5WZxM95K0/sdYQvCOPEnax4hf
11Aalv78bVzhAuc+ks4qomqwIqlUlRa17MADsUC9JcLHx2VQSFd4c/6WKcZG7ygaFgxwdafs44jF
/1zjZBKdTj48xUppxsu3Qtw7PSW8J/Nmjb4PtxjWVzVMk2o9+ZZLzuAsP22OZ5XnabgZVZMdudeV
PGFP3hGWbfrIaaXXBhpkUeCeDl2cj33e2xW9PFDVgrQzXHXNuwXID79c0kATFnX4ikHVf4LNQK7y
iSLPhoOgLsdoEao2Uz+JeRtHid3jh0Rd5iKUvvqT6sTqo4/zxWYgQVnsrt2CiUjBIvXYFVYt2Kc4
NqDOFyi7W2JByIOeG66NJrMnPexZKwC19oTh//T3PwIcG8eP7DBLTCrKoff7LYDhD6jOBfUctROx
/BhA8Zk8THKPyRODqJtXHGrD3StgoSkE3MGI99ZbrPt/PVNiNhMwEVZiTHLLRy18OL0LsxMtiVvd
bh20TOPNk/otT/LUJsKod+OVa0fTfwcKcCHCaT4EkV+S1+UFIsZuhnhVmmnfvDygW54aL1KZbhlZ
l8jYl1kdwYQDoS38iehozUZ4az8g2Vs9DxtODCh4t+MasnYtzZynKI+qXnO7j0I4A/+R7uUP4XEd
XE0zwjU7QxW/xetAbpEfijKE05FQ56frsze2nTSNnU6iUgMnIkMGaY+h8QcdEnsnAZ+e8VSbPgyC
sDxK8q1X4F1TJpVwDqy2jVFzR9iZnhFOJaJZHhxXL2dO5ENm8I6IxdcpKIxM3G3GKXsHgfzrpExJ
wnAN2Zka1CJNugZ+9sgB0QLi39ceSwDtsrIAInn5vcMPliBGYvtdgYks6XbCwS1cKkBQ+SfWcj7G
rBkxQAtAw+v831O4WDR9z1rPEv3Uv0KJB/xj3N0OR/OzolIAZNtgZ44ZTDuP7leNpOJfzXnsETMT
poA7KIKCefHH7Oz76pWhVDhhvFoYYNA0X/y+QorfTPIa4EzRH3HSvp77wvwazvHpkYm9rLAKwo5W
+NEhbz0tyLMz4OQBxY9o1q3PNqMf3Kr1IZM2p9HD0Fhay08i5LVOZJGcDIdFypIdfcAUtDuJYRQI
kZX1aybEB9kDKo6iwA5xdXhLpBvVMd71p6ltPP6YS+TyVuie8qBGEbHohFFPxDJm5kKLus+L+kMJ
0gvN8XxFS7jUyj6LjfToyTy8T68zf1BqLO0dAKfDlvpa8IpybOzDX+T+CMrkVNlbLaMO9/eaB+tb
hC4XxFD5Eo0k5CrOMwcTiQEOx7HUVhFeK2yFWLanBWQ5eE0Lgnbfgr9GD8UprWHpMDd4tvLzwLR1
ZHhYiXiXRNLlvn4cDXtjiFPXInqvcK/A5ozF8xs8MPrBfrK47JZynSh/guGGOKIgmPx0bbfIzxba
bhBbUsgiYBeVpBqH4lTfuPtLHbEswROWhTIL2Jc9UR/Z9ewU93XVrRxs2w7iilstKxrob9/Fcn/G
2cKwfuCpasaT5aKDk7JkOwBVoueIyZUCqvQkkVQbgADkAmEAwERJR58H5MUiUQy3u/oEV9UddlkY
Wa6dUamFp6hHNVDp3r5BMf0ZHZD5juLMil7yu4RDYflzb2Ha92eGL6CVZW2jiSj6b2tsuLHheUQr
ASwIlZThB1t9ASHYiM9EhE7pnVH1GHLOmKkfyWGSCauLTVEllb+4EHMsJ6PQ6GIavhVzYCnDgZwS
eS/AEUm0taT7KNr69ATQ/MyfzTQec+1Sse2ierX6eTxY7edt34mY6GVEcp3od+vDmAHxILfDJM5N
jy/at0r1W+BtPSZm9xww7D2ultvaQTQHoA2rCye5rpk8vFn4MN02xPOvGxSObQEJ14b/ueeuBvl+
P/lvaVy78d9wJCUdtBqveitnm9Yo27hirpv0iNZWdTImDALTHyoaRtI/xmq87eN/ASiggQAstjyX
NBqpvTawNFt9cqzJlVTzBkxfCM+Zz3JCCVBqT778inKySWwHrn9xw2Q59t91pEfWixwIWCQ2qbMK
n3Q8UM0RVIK9LUG3qGW918UD11WwGHA6M6a2bHQn1s9668YCswJSJ/b9SHmE+Lp6q9jPn4qAvLzH
n7bSMlQJKk4BibfFHPRCeZvwUmPZPmQLLzpJiDr1/LHwgVGbsTedc7NEouvvh5Rr5/dWKN5+MJnr
OObYvuaXPi5e1aS9F1WgH0YSTQ8ATSe51PMu5TmC2ZlYuqvZ4NoLcH3DiruxMJtD7lfcTpBl1kCI
m2r4W4TWx+3Hfl1KG1BcbvPeRUgCwK9k6ZGPnBZUiiWELebqdGiACfzDcqjVHKBUeX8Jg+TIvmuK
o5yaPj3eO009jYsZZPFwPFhT7QV7wB7nx5zRqBSn94Y1oIXFA8ijyNy6NPzMFC2IhEutKDke76iL
uBfVda8zvDbPs6meM5zuNNZ9VRpuZfm42+5Op6WqfLhh0Wu3p9LkSn9eg7wO4RnU1cmNQEF3YZ/A
mC/KyAAbVTWmBbk5k+x5X+1KbMkUuZtiqHE5Uio+5MuoXDAj1g3AtDkV8tAi/qGU4qj2LW7r/EZP
bGkid4U6WYzcAonJpCwXeD6zPpaMjhbUUybK1ykcm3RtF66tPGjU6nETpnv1KJh26YuaR06rLFs/
3pO8Zxy9wHvPU6zPa/aNE6Oi8hOPcpFNXH11JUaN2VW/cHcjyqem+jXIGip9UB934xxvKQLdaE9v
+AwptWUO6raOxvy8l9svgGVOW8OfBbOjTBgABCxWncO0Jlioqn0Q5s9V1KG2wxZe4l8R/6aL68L4
XOjljCcn1YaJmwJd1saBloiMsMsTgZ2S5u+3r4NDXJVnnaiYrlag9pPsIb9euJ5C7TgCdIqZJZn8
GrOlkXfccvtGArLvBJd931Z5cJQY63Az8OjVB5vSc2VE5ClwRYTg3SJHxPMJ5MLhrEkjrdtx4MEl
OhoIQ73EOmiUDmyWO7KOMLqfy8MJqd1x1u7PhhRoqT/Q1z9bdDpjstxjvn5fRq+LjzDNg91ro1vV
KzfhXir84JdzcX4LXwcI8C0weAmf3Od4IzD8P2TRKv/VbKeyTHUqHoJZaOC8ZqH7pNbIwb1Kp8RI
1P9LtKRcIpiTut1fzX0rlUagKoduqZ10BpRa+e+obtRsh5fn632GA0vOOBFa0hWG7L+39exGKiqh
EH4w3MzSa3vCWvX8u8ecoUQwrbw+xBA6fWgn2mpw/YP5LaJo2fMi90yvzrHbz/IC1a1fhyoK8iyB
rteHwTVKWhF0ASg8Z5Ai65SYDzs+nC2qYQ7Q5+Hd6xOOyOOFsviLLyZgaU7ennf9VHfpbnECMnF1
EDHd+0kkzjY9BBdqEKIQ+LgYmMXiIx0qfzc25dphKnp4JVl9QWceW5veZUb19JHrguS3hCgynKXF
P2qGHUbFdC0zYVofA5kv8IOXwcY2DZMGZUktxHbjl01oLy5A7SstECbmCkQ5AyY/TrTvl/t/0QNc
2sKNi0ZCHZD5GdN+c1mSs7APcmfL8qQ7fzg/PMjYRZpkvolU9EFDdjJKcdXLiAx4mcK6ZB5am55j
8RlrujOQ0Qtx110KxKVsDUN30j3lhhE4K0FU/p3U/y9Dl98eBDMIeBYVxXOdt+uevC+aMgQ5ORZU
pYwQkl3VY1XLQgSYc1td7ib3cSVWpMWXr1z5onijGeT9ljwnxOpHC5rd5Co3z1BH6l36izIkrjbL
MQxCSZg9Leu0JYupylSayegYvYS74qicGmnx1URveipVo+TmuAa43aihbqA9rrGZlrf5SS0lyuqJ
8Khz9q5cu0P891Tk5BmN50pWC3zmETv2M80hTx1mKlWQfemiGv6wzPjeJC9LZ9X3di1Hku9UrnYh
4FgtdRkop63MrAa1gMIYjm0MgsxZo99Q7cAfBtrw/JlgsGSBeBNJb9CLCPiOAPIfU/uGQK5MVhCU
Xr+Rv1cqZNYI1pyPDaciIgWhGJAXgQnYJS/2rpdKQ5QIHsVtTEbzSa0ZvoUJxnz3thR9+BF6jZNL
CN0ivqsnTBR0x1pIvb/p9VN6Qsdx3GVPaMbkZZMGIx24u/BkuP2w1UEtn8GSX0Wi96FnnY3Ah7Kc
DKOVETBCZSsi1WNeARJfIbMsKRhBy37hYc2O93eP/Uuyy0f/jMjvHWgW8foXEKEsBfk7BrMqXQcj
Zs5uTJMoSxjm8BOioDEBWRbC0X2pCgFLzG/7U69ETwBb2dks0qmOHg5ol5IMdEo2V/wFY/I2IY3g
cUTEFEPwSBRV6C9gLzRSqseAV32BegIgW5aklj/S4/NrrrVN5o2B7DVeT1laYqHSvanigbtSJEnX
hhp/dMNQeb194tWCF0GvHYiEORZralDDP9fQtBR4Jzpd81wdkNLRWjbRRtttJQqNX30cQV4P/eM/
0aaJE5Udwcnl+Y+rCn6pSTiFUmpTmlhO3NBG9bhkc9oduxuaU0pD/eAuD6A4igui8xg1ZJ3jepFe
gvgO7a+81AAJGXgLMQOtJ7lWWqwIeQRhc7Aaml7ab7J3GKtTdg+ROTOCLa6VfRCVchXugaxNWKSp
N5mxQaCrrGeHd7MrPqe1aIq3X3/01nskgRHzKHJwM/vRWKL7GRQKEaIyB84hWeCgNsq5VhVCRBz2
EZuoDaODlN1rmASSQ45FKMfIxXU2LpFoVQfAWz63HUlEbv+IAt00FVeaqAjQJ+Txczl/W7AV7/hp
jvxH1lmHKE78vs1d9tZpk9pZ8ga2Y+ZRRTFazOm+jMCSMzuvL41Fnh2EDYTo3nPFU/OYW4gPVlYU
2Eu8EAeFSJI9ajsx77PUMscPtoTZSOo55/WKsY0Y/OrnfU8M3t6e7UUUTDRbWmFboGUoOv6gCHUo
fa3iXL4nz7najVObsPV19MB6xMF/tC7QBOjcPalpHUzWEB0Z/jJW1oAB1+UAeucXqTdXYb11+ge4
XX4dLgtnOXcEaDtP19dtLFyYxXvUm21+rldhHRBnbVp/Uq9fyEjm2zwx/BPCm/5mo50dKCZ2jTXi
HSNRoQTrw7HZWRulwJR1zqRCt7rTUhmU2Ltk49tJOiPHQrx06ydLgEeGq1ruJcEFf4P4YKnDBHlh
kRg2W3cWQIQ0mM4NVUhGul93UkAzK+k4nJ/xGdNlDLJj0pPlIGaGUitq6AoLsEeF1Xkp+2QMnEo/
YZcD2roaHqbbNg7HprbFS9jWqtMUIwc11Elzvh6Vn0qXEjLrwwTMdshk+L83k/pSpinplKevZ9jj
k1BDi1Gon1C25IPg54ak19SUIqp524l7NUROSRWE2rIt7SHuVA4SNr4zZEUtZTpxcfirmqWrslvX
0XxMpocxb0CFEP1UjEJgB4xwWvRYVIOncfBXkIoO225aj6fM+j+l3HB794YK+TJqg9Czcu0jMJDV
0tSRC57uQ8/kyBLM4wnGmGEtKRDLXBDrHfok8ujonaecHA+Z2I8+taJThyrKvsi2ntUGs/kY4b6d
G5ls10mkL0Oofq5SKToix9pqmBxxzRJoeDw7NjZOYBRdqY2dvzELH32Z1lDC0+PFnUDmSH7bX68f
rByhCAlbcdeLOeDlG+fSwN0KHUAZQ1lVAgcqBWpruT6k8/HYeEVQECfEekYqo9BNxJCRwJpv5UOF
RL7eGcTGRtgL3AmW4DRX6pnjYBQfI98IujmNiRIPjUygNoLJS4tBnf7bWB4U+5L2Dht1JbBwaZmn
jX9TlLND4LFfpXsGmaqKKoe2WX4SkdOr6gn2p3A+ZiHM+pwD8Y6fYDLTV6uZVHsxiK34cUmv0aKy
T2b7n1ZJDeiYC62nyLku3/Xu0PRBBiX8NYlCFkziUm3n2xIn3mQ/eR7qnzduYbRuPyPH7wZhI1wJ
j6uga/6XjsXA618JMIlWPL9P8XeuhFtEsIPmR4uc4VBLpJzIlS0wT9SwhR9+ULEnZ1Oc9+REKrKm
Ygq+JRHDl3lBDbq+NOd1v9jnHVLIzq0eEzHcSmU2g3jYTCVE+HMQEeqBUosVhCWGgh+HXdL7V2WX
KEf4D65iSL1Cl2tpS52keWNW4rWwlef4XeKDEzUdDHUrYKyKkVQ/riqUpZpvzAmYweFw8seoYA9H
QTjtyx8qvvfC7Vjxzg86nRHKjCV0fiYS7v7bC6nDlj7Fa8tKVvn6/cWwRSk9CnPiu2TDjdG6Jgu1
kCq4tUdHiyfZKsm4HNjlN0y2ZC2ADWPDni546bJQiinuai0FvsCzp15OLGNxYRZsykcehAyqgf6a
a4EICQhhZyCrAueQMFDKAtUTblQX1v7FAKjZiFSIpdB2LDj8P7dXBdJRPc+l7DDlymPmDOLdh08O
p0V5U5XzLTTtqYZiwAntY7gpx5y4FJqmtsSuXV6zdcuolj2ESiQoXgOMCVnYIOUDprUuvUif9P/v
XkvD43Sq7ZtW0/iTYpHYD/lvTHqVDtZm50V0PjC25cuC3KSmQxT94uyMkeNQMNrk116XXfOPM1o4
DUYUXWOdlX1/AX69D6emhnqLZFcBFFONf9Y+iozhSVxPBDKpFyVGzhZO4W2nqEUBmuTVtO8qESDz
nLiN8LxSK7ZjqWMdNaKYsHoL3/8aOimOa9zoOS1S4/XY80S7NCl6ixjTZpfL3R0EIt0cX2HFkUtP
k7JNYuVcXek8ARBCJVLDCD8pCa7JP83NXgKC519x/71PJOxaCg1dPFeHeaM7QJIkVVY/ssXR0bXs
+d7LqcF87qcfDzjwHD3S8XkVE39j0nr452Yt56lhilKUjZwu7TMetAUT2ZaaN95JiUTgJ8OuxxZW
MoH/HxukY65KPO0Wz5nc9YXsBhNYmDIs9uTzca7ynzJVemuS1YfSL7TcuQxnMbvU55y3+O1t6fYr
d+wNXpId8YAm8XETvIwE3vmsfClRBFGJ1AZBxA9Y86JjE4uEu9QT+R4gbm+rAeoHB5HUN3dDSFE4
cwk7k3FyiSY8rdRsY9AH0ROi3GiODgEUEOa+HkEYI2GEd3ot1gG1Pyjb8RC7wPWscn7OiaHroAmv
BOQeefe3SIdhq9hD6Qx79B7ni1ggKM2J3QGOjq9LQCm8HZX5OAmVHf12CMVIpmJVT6sFns+nCD8H
jaT8sUbL9wICnLzY4/kEo65tTIJNRBcaitfQJo6cQhtboncv0q6MxAthn3tWrxtmIXB0nik5Fp8v
Zi3xanamGbCjlH5FihrTzjaoP8aJoxDa94ePYkRMAOn3PvpK9woMKpdJ3SNT9BWLSyY9Yv7KEHtw
BpO23ATrGmoREJgECJWAEM57TKfOP2fjVWygPq0A3blbG4z+HTITcozAYPEMrO68p4qnSnZ9K7N3
q7ZrdlcajNZeToXW3XL6biCS4N9sxWYkwYsY2/DTCYetGLqLyyap9fIz7ePpG9xfieXaMpQYIdu6
uhZy/5P1KRC36sq7RDhlozt9ttsCY57huKwkybxN7R/5aeJsswyr+2zkapUWVhuMp/k1l4Z5Y/jV
9f26vD8qFywuAPd0pu6ZiI3ECmwNd/xDWQtWu+frlNnNjdtDnRXthUvcV0e7hZZcMwipn3efBlp7
08z7UxLKNCW90TuLGjWqIIwwasJ0oyGDO09A6vz20Czl/clEFIqMAQfEYmTzA+LU/zYMA/7OPMMZ
jPgcaN4kS8sxY8Hfp5iac+tFNYVordozLCoLJKyrFd6DABXwdGqrjZT6YCTv5nzEfe8N8bDtE3o1
qT9/91QMlKX71pkwQ0U/EiT4bB5ZGlJlU2eDNDj1w9keOIDuzw1cIyX0rmblorvtY/6HmHX6ei9P
ku9GUUMNQlNXNQ4BEmFwOHpLTBQSENgMkVmavnr/CqyZcJKEA7L7Wi4n7oubj0b2jSqlOnFmYS5Y
LsbLjdJOjF6JMuhhB39Ed0AflKJEFbJ/XtPwnCU5OONUnCtnDrX1eHaA8iEtrBmv/yvwBEVMiHE0
5KUK9bRRQs9ulELm4lgfzRSVETCkrjymddhjcrSR1W4ozdlDc7Xr1Ug7dCgNccUdcLbi7TYxRd9r
l7W2tvuWC+gghz8O8ROScOrteT8vypk8zjztaY/ZP2yDPZxM789JdIZTjB6ojDF6iP4ZmSPzzacw
3JikE8dsg8A5j/sZn3BBYZ2ZaWRrSh7T1+jXQzZ/aGitz8Qq555rQ5gaa7zrFBDjcA4x/TSCgCGb
8U0RXmz/+MEo2lVkotodJ19qJzPVP0ZjAxP5tkGfnz2QrRA6HvtwZxFOHT72rLvgAeRV46OGaZTy
kVJgdQXQG/C3vmQf+dlykuJIfzenZsn1JrhXrZy4zFruJAbVnIp6tUGqwn9yLQ2/RTE6ep2bt0DV
EIbOW+N50NlNwlrKjpTYo6TXF8scYC3T3JyXNNezCOTFku2Gv/1SJRX28fo2i0YVnSHWp58Yc1/h
MXu9NLOLiTZAaFpT/MtxNPkEQNOrxyydnH4oRuxuVCUA6w7D/4ooDeD3b6C44gd60Y7DwCjx3SsC
SZThgQFs/gjXX1TLBJaccs/KBpBmj6nLyRFhPNpaZANgLDQWjk9AospVWt/jK+Y4v06x/qLZO2PM
n37HHfz3plTNvDLNGIhUH43v3JMa0glQhdAC4uicYxUmqh5UFXKefia1Y0k76EJYuWC0MnQgdt7v
ycPgv5KmZuz+Fz6vv0QfqBTSsccWMs64lrQXylypYvd/8CEILOrTSymbia5N2YR2W32UM2Y2fF2g
pu3DjpMf5ZiiLfioTjL/C1/c1vWjNSUOCypo4FvB20eiUTe66GrBY6EyBtfsev0UqkBHuk+URM0/
483HITRHl+wTmOAKSWJc4x4EjYmxbQ7sDlyeF+NrM2TAxbPLW75JhQ7nG1neIOxreGCx9GcoVd6d
EyPtveceP3WrlskGeoSU05KpQPFfq+pHBL5UT5OYie9MwsfO5GfV07lSiRkMpQtgJ5w9J4j8v4xQ
U9ZoD0huWZtLeSlYvaTIRajKsgYQrZdfTaWDOXLNHyAXlu6sKajVbomB+9HPb2u6mjLFekpiTzvO
BtGqQW+hIJFB3v0X32xwsppT8q9ARidXvLvEsKqB6QZV5jEdhTjRGn2SkRI8o1lH7RFE8+H8AT9G
lXJjfITjBJu+3YbFtrXvVw2nGvrYCjV/eyxXXnA7CA3L2nkjYmIesKlND/Axz+XvchOmV6uTfRn8
flJ+OGabECHzMai5K0EapECFrlWe/mdx0ZBkUYxauddggSnUFiYEPHCJVkwQIRBKWw5mNhRhGais
fXsfRgwAnvYTdAZCn8sFwy1VDRFQJE3MZ4x/agjAMWL0Mv9t8zgzqsHboCjUu615SKpabs/SNno0
g3Ba1ZSkc7AyPnJFTauOziurs+P3QOAvNV1qzWNPG5i3Q2Cj1rNnPFgqJfwLxSJeV+W2xyVXl97M
/XojlyJsJ4EA0yyMafkjtpc82HtfPM1tbAYUi7nHG5NQzKkZp7fmZLeY1q+2DNZPBinT6hTqxx1l
LBq8Z/ZGOEUz+pSsqmibipqfJeJqDd+eHyVApfMWstEiWz4dr3zrJ9aTccsRrQrI4aRf5LKTkE0T
Hne5c0UUFY+YUqJO1UOF895yYk92pXbBwZ+6smIfH9lpU+M+ZgsQwx4sdT9oF9xg2UjWQC2bd2Gw
+OyhBDbblswzuyjOMQbH8U1qJGJb7GE8fkg3HTqzB2xkGPKiAxoQm3tHG70K9thH3yFPikH61kBh
bOgQGt+VxXmr4i2+FSig0OnvplyAtpPSjCP6nOlI4Af4WuCWScMNQQcL1NWWHhhc3VtDP17ZJ/I8
6dpEbS5KC7lGGZrAF44wD2IPUNBBYHtes8Ev1lw9hMLkVqVPe7Dju2pUGlZbEh8/uQBJC/nFP4An
VNVRH14IfkB15pqe4ddiJzkO7tNZQ1suHeDTpevdOIykeZVeKvJITfj0hMoqyLB3sN3R8SA7aL2k
6lSLq4wy1bo+dnGjdP2AskzZI1GyaQHJmujkG19P8n2/dGqgXkHFLNf1zvLXWZ6t4K1HK6sr5nx7
Gh5T/6VPNVrAHPXVb2QHGEZwqX1I545TZvDGg4YcJ0aw47MguK1Nyrsuey2c9sSrvNkSFElTtsYU
+WdISSsJNeVxt4WOcApDWv4lBRctWDt+zWLAMVL0LMGZc0+N4otEh2pcoHXMMT0jklKqHTirVZOx
G01LacpPwtVUQBKLf7KfRZwrftvLRPjqn79rE3vM1QcspV8++yr4WD/zFRgY92u2VV95ZqCNIf17
a9MriwKVjni0GBE9/Cz7FoTK3ecsrDzq93oT6bMWlrdyZ3wFuKvhDJozX0Gs+T4ovltAF/5trKDM
KozskwxrPyHuweDDYueho5IGMJ6eLbIIu/ME7UNkTLC1lSWnBm0OxPxN9V8arlZCy0Eckg5m8dJg
ZUZ1+gTMZtqn4IypaRvnDxm/gd1CFBumrpvdV5GFbju9TSePiipg6XO6jHkuw06E+MPskB1AJiN7
kkTinYUeJKxtJRq19CEi3T7WJQBBKlLi66jZ0djuxm0AcYKGWEDqY1rFehQ4y0DDCYY+tFwkR1f7
A0sMbJ6oBIU/5PBW1xCN+JesxBs32RLifp/qkikWWo9dsmlXBt09yTIzux8jF5H/nVASfQetqxtj
U05u8jkr6gkqVrUjW/nHK9FcRKlJ66WhG9ST8dluMt0IaSblJE9J4FSkbvYoVuUlPL5CtY/zzzkt
yAh8ixCTr3a0Am58SfcR6AY8cQh9OnOBAGzfKmc6AXPqkqALZXt5lGlLe2ENa/++4xa73YHEPTqf
+kQO56i84oVZNx/myoo0luAhR8+jpofGOamP1MgdIilEHJev4N/EF+nRl2vEEGJJEIk9FbLHzT6m
j60GRIGFT1cjlKLCdLQc7b/xvmQs6MOguwjzmu39o3P7eIc35KQwMWinxpB3ZZzftgIbpUV9fJeq
7nm2tYRpLoSX6HCmHM5ml4PwWxwBnxzN4kdmxcggZKQ4LE+BEigT8prP36mBj4D92nrdJhLd7D2p
BFrrwpWSYcOHwgWF0znDhiVc46S68r8Cxjj6PWf97wQQegC75PmdB560pq0yAk8lHCgGAiwcxiN0
7meOk77MuQonqNrsifia7EmFAaHt2lAlYKT9vd26ms5NuhQRxaZno1AVUadgrz2ahruRs+4QzPxX
5ywZqes23LejR1Jqhdb8n7XQf/lYqWpwFiY8nf0Smju5Tzjbg4pRCwNtZVlDWsfwVE2PGPgwj4W3
AE80YBIQm90fe+PF8wVu0gIUWd9QB9Mmfo8UpxnoHIRRFJCv42wjXhL1k0D/8v9Bq7xBZ4Y/xE7F
9jp8z294IXLpPOLfCtGpAzkcS21KGyTPZ+ItpmknkoF3PKetJZ0cqplr3wKPTEsSnlOVKl+Ee9rR
DNNZ2a/QOE0fQtCzmpPZsue3O4F+XA56RTllNrm3l+J3Nfoq+Jg5Cls+daKU0d+h2eQrBFcyusHF
u6IEOPdqNpOoq+BOJL4FhWrWDJCkFHS0UkyCxHMHXFPQn4mCttoqQRMD2eI/VCyzkcugaFR8WKLp
qTY1SEOmAEONbyUTA9Z8rM+StcYxSFJQhwTMStYCP2yknyXadIJ1wP94EFahfWzDExIBSJQAn6+f
xUkpawhONvee/4gqexSnkgFqtsoJTF9JLmN+AUsial/K1ar4rejg/GUfoPQTvwPfd1nfVkJMQfX7
C+S5moxiRmPUZDtc0ZOUhYUgtVVTnTLC1oZgB3+bYjBpmjPRVZWhXdx3NGx4B1cqbVxu6+0k7oea
C53wWOeKtbo1LT0Mo7FrSpYaUH5XU5VcHF4O4L/qulfZ10LToIjPJTIArQogRs9HpY07l0GluCHk
k96S5oXqF2YUxLDqNT3jGLxMIBr3iO1lyRmhzwGkxMTSuO4Q3fhMp7lQgq3HO3lp+3YkpcWN1ryj
aFzh7qbkuMBMNP/gj//ZidRP3oA59N04WUd0mjPAD9AurJYoa+FNKUGjhwgRFMSjhX9RsqkMpfgh
LeOMhMXh9B8U/4YJaK8KHnZLvFOLv9Fz43PxjVIQxkcr53YT2/18mHWNiqLmU6sevCabqtrXUb5z
z0vWOx5TBt6Mus6CgVubMzGhkjwCqi3I/f6d/BJAcj9/tyMDpYO7H8yTapG38KLAOT0QTyg2oOR+
1Y89cJGP1d1WkbAAa/Iwjso1A54Ok2Xrns+YYDiij6wwM3M+LRvM5fLLRF4P2m+tfpn6g6MmwV3W
0rsZAC4jArnawslV1Qoq958WeBKId4pNIRXIRhKBRkN+QpMW/931mK+3PM0CIx3R4hNeP9/8tMwY
vCx7iXr9F1zKba3wHDoXmv053+H3imepfQ/idRPRrfKYcLmpmWhM6ANuLpDXa9wv9nvrr2EW3aP+
6LAHEgDQk6M0+bPvri9Olp12vcBLB6+MMtX20eNgIWJmKzozKU20Ya2bGm08Otky830dbWfZDIrz
Bl9HpZbUGiQcP0IPJGnWWvTWVFFtEQsfUVLy19a5Q2fGiI67JPmVr3imFE5bT04Glf7Dx4K91Fmz
kpJRI0N+2IHqUQDdJEMJKOoqN2T7Ul1OcLnLMEiVY5T47/tMDi8RQKTQ6qVzSzv9PLNQ1QKUifvU
DvqIFbPehKKedNIBOGJcRfGVYjMyQ1mOGzk0K6nQZ2vJP3ukg5yDjpnvJwoSVeYXKKSE4olfohKF
z3yMABZr55GzV0kEwyHyL0CMqlvAJffx+7/VQb7Zf0EVDcEeFmiajoKYMeoLBf4IHAyjRdIDUBgL
FOHXhwfc1AL03j/qOPMFnSPAfVUu92ui5TXdlBmiKTXRz0qb/r6C4h2ySobIU4/6/wtidiMAxKM0
ENP4bAnt5Zz3B3HTp1EzntBD5VyHvb+Sak4oeg+8MVRLaQ7Hi3hwO2a4foU5YWcyZx9zhONkBOQj
tyIOit1/YBAL6Tu0z/f2iMVkZEOyEEcZmWrPFmBjyO4mg08BAnZYrqE+M4axxqxVk+aeSrtELXFK
SVClo2TSkxjO18y19S1wY/j1TLNzKXULItWepaEcn3y6gObOwOTEHiHQ+kz12oubBBOhe1HYjouH
9vuMU5zvmosIIJNrotiuFaeaZ5nCS4XhSReU7JYMPhnrjYikYJgGQaPckVxQgyugL2hxdkVbDIuG
oI0PoPmvXjJ/FjArlwunhVzyL5Ng+Odn7saZ5HeWRjjGXMDzuWcT6/ngz2CNifiEV/znmLQzX3KJ
G+eaiYNWPs1/JIn9DrZR3oePBhOekWYimKkdUswKfTKDEflBz1CIE2JHxzVkX2h/6dMysVY921Mo
KshtMmh4N1NjdteLV4m0YxcZY/9rhh+LUgeuy2kUuMqRiBpGVnBOcKeESQxw+LWtt23hIO+TvAFV
XDnOZ2YNSqpGoGAD7OUzvHpY8gsfS4jew1+JpWN/356+/n3pLSm0rJm13FR4GPSS1UaMscmVw9FT
g9wkvTBh+W6WyknvLcLoDpxK6ubKWWDdioWKtoO7Qcm2oDGZKNiKU/dFMyuesCqzCtM/uZ/3mFZR
RiTCOGpmL82tExyGF5y2K7lWMxtGnE7ZoaRsUNi/cl4xqittonKDZVcht2pxYNmtSOL990yz+jI1
4pibS8PtRlJG9ql0L9fSyHDHS8sxCG3I3aDCUCXK4Yezral/3OL8tDJd/DJALw78XNuhqp8La+T9
AvNnIZFBTXu7l+MyP2VwUh7A9ucl4LmAE938SKTX7Hf9yPWsu/qc4xiUQsNgwamMzhHS4eHZ+mwn
+/vW0OQ6DFnc1fS/ulUWN8Re8JiQiNxM/RS3zeKL88AB0wGaVTDBQ+OilV6VUSwGVneEr9z3MNdS
yhThoLaSZ8vvqm1ViPPKrg3GizRpbY0bFs2ZdepfbjoP0+ewCt4bnCeT406BZbAaND21MQ1Q5Heb
0P4o9s2ewANF1ewXynvpp7Y4fmXeknRLZ6c5RfA44XvlivGV9HfA1e/nabPS8ric3xj1G3PxMsh+
b+HopfhyuPbIqp/vrY2KFZgkADSAlBJ9q7pHAMjw6sUZ8hzxRAmuTPXPrP/o+xtn5A4wxClXs1ok
zpVsA6CUv+TZvf3xny6zcC6hW5woUKAGazZQ0wLJm4YSruPqdpDQ0cHZj394HHcv4swMQ4C0t5VA
VhEx37BSAynFyf+XMr6HihpIuRHYwAh2amiXJEYAM4bV/kjwVTMcmPlP8cQSNtP36JhU9dS5t0vy
cuiCT/1uOfNHh4WUGUv4SMMjmMSI7ENWn0nPDWbfLAhTJzcOZ90UdSXPc1ORqWtud35NGSAVFqT1
ZoyFPAmtUaIHOMEx6rAzQbsvmvpWF99aUlQfp09THfHLnUgHvmGCDklpOK2nWhlBDIhUdT4r/yvF
rBTjvIgRuuTIngt/+x91kWYts9Ykw2Foh7yGFMOgQIx6bryQhB24UKLrHk9iyr1abbYIhAdA1kgy
CTyvZNwdd5TRHcevSqveP0pP6cN5PzLZcr9MfKVHqCC+yDJ9DAVHZ8jJf8FhJMSLQJ8y9Otx/3ZS
3DRDsQ8VWKcViG2Al7iCW6XACO3W4ijMsQp50BmDXP6GZZPYDzUFKrG/aeJY2ULjGeQ+8B4cJn8z
HKm+hiBxMni7FgX6Q7WrobWKj9At4p65cdwssV5qj8Lmbw7xG/2ehKcYoo+YpQNUJDlGQ0bj+t9b
L68o8VetYpI4Yl1/QYr6GK3RGhpD4hipH4uLxvlNtx4InRfxKedWagxJO+YRvEyNkRXiA11bhJpB
7ZYfx92DcjDb5IeOMXoo+R8qhI7SNo0lwZTN8mfq1B49v3Nr49ZhD5kjhsmHuNb5TEHi1lPSy4Z3
8tRwSI5Hg1DvO6rw7O/tGS+/ymg8PqeiL6CJ8+qaqTw8C8VFFgi5W4R7bcqfBuickfXN228PvGx+
SqaoCvVKGqFXs5C9Y6MyLTsTtjNOq4xdBjqVzmXtHEbpCy0KatX+Du5hU45aR0dCbZsmrn7gVt9W
lwYRZVob5LNBgX7NnnH6DJWEQ+Ef/BRXZVYTPtleqqx2jMHOrhCdkFGgYCj7gl8hLf8yN0eL3h0i
Y2rBmwBuOumc+xM9hB+8P1A12tgncwPyLEuY4QOcVd6mX5sAVVBdyAzKnhUsHF558nrZXctuHMFy
SamiizVf+gxAlnvykEUTYICVgNV/SxcG8Mvv9T8Kj/KMr2NeftzekHIbSNTruwHeHeSpkvOhvw17
2ASrefDuoUSxN0dNCD+roMglR4+tIdQ/j4rF6tbSJUOqeCeFxx9KTo/B0+CLSGWyOWYYdichFzVD
bmjptqeYVQHmC4CC7CUI8kb8f4mRFm2LRDGIj7AHlkrTt5TlLwChZNPo+WKb/xfcDbbrZa127Rby
kQIdbyehWwBSK0AyU+wdkmBwYRWbr6RqPROcNv2plx/JEhMcOksEQ5LuwedqS/+ekYL9Lq1rz/1M
JWA9gptG41VQCG5h4HEQFNky87tNxgcZ/D77ANZc0+CVk8I9xSuatQxEUGHN4Xz6g9PC4BBv1Mlg
j5OE80kJ2hyqEotygK2vgvb2qPbkLPsmOOThu4UeW88e/Sc5uFw8cC0Zu2cF16AHg7aE6j0oafsx
SCcDPryWkNg1Ln2EsnkBfv+ckPF5n4HRmx7kt6BxW8YVA+wODL1/xkEn+e5hmtudn1RWYwjhgfXH
I6cCbJ7jpAKSv/1Or4oAaSOMhtS8mjhaITL7een3Kv39N5i+K9WBYi0TxETHPSnkHyVc/iXnlXip
dhULrTptw0cetL4T9xdUaSjRnzWdK681Slp3H8GZmBu4ZhW1ZlifIqNVegM7y5VcZ2vVpOdSKtKE
BtkdDaJj2OUNfri3LHrIFPBYSlhuW3K00TQhO9HfwYM8j3fDGuqruQZSU9sZvPEVOXdWuyuf2JOA
AmN1w0af+NA6oW+nSyT467k4U3ZU5398jOCI4Tv8SXArxLlk+FWaCsjmT8e8iLWOVmqxo4jSmYK7
2AdfAxeny8+actbdhNM33m466QvzqdOMf8M+RDAvVmjqp2QSoFN+SxxTuU3h9KYF0alHOeDgO2Mk
dsbsbHKGA5SHBkpxkkxcaD2D2W2NXS5gJQYNhnGxTmvQJ3Z6tiVI2q904CKerQaigYD6P2Z6nTgi
qfEhNssSQYJpaS9TaeeRxUewC7sTIMbeSVGManPG4e049zQu7Tb/raurA8V4z5cHYqYf6cHdAoEw
UqS6OHBwKFSdvP3h93NSLdfg92s5y4tLc0vl7Qb+b+23hL9FVvEGVmDFoZICthk2FwGBeqG+zWhY
arRrLr0cjd+FyEmkyky8JRXx8ePRwJLEq5L3XTkIiJLqK21uPY9NtTmPpbkvgj6Zl8fzgqwMIQs3
GXsVVc6ZPdgv7jlc0ggS0MRRNHhpGbn+5N1+d/HzdMHErFW/7NWVvu+HMM2yn08by02z21Kz7awz
FYIvjHjkEGAUmjcOTndoOjIRcMDDMm154XX5ouQTLHlRQBPNaVaQ6S5DxpDQpnmoji06Ia8T1ASY
g7a/aQVwtlXw3ySrd3nMX6C4qIWUoXzMKWnqjxS6AysRXpnsjJT0a1GeXQ9jxATJwzFcdL+EKXDv
H1zxHHNm8BJ8AsrGtUlWYFnlSloi/XwCp5Bxj3rRxd0An+J/uStQxQF/8b/IQflpoxDqfcm28PLv
iR0c8jDl9s77/aE+YbkX2UY6mI2WERUtCB8MGR7AmL+4XYoIqdjB2fZtt/+6zD4fXySX7EvvtNSI
XoUyKGNuKTa0YwHvk6+QRPuD9nlSmaAYzJK5gf+6k3Ujf2pORKiDggGIwpQU85DO4eYbtM5FJNDn
ubMS5icE0WPRRlRomGrt438mQUtV8SAbptd2sr/DqdQjMBP6OLWMK8Id0wlF9v1PlNEpRvzzD5JX
TY/EFlvZxDwK1H9kuePKi/M+d2VqAvjZFoVIHBu2kl3ZYL/PNx3TiY70DGp7T3dB6QVG8laI8f09
dJKCvrOFlvSi8UhQhGI0qA1AyK2WkJkk7qz01V4emZl9qyd80k81VVOMF8j+yLa9OHOrsI2GUwQc
KGfcSghF96iELwlRNPA4kOR01TP/qD6E8UB94hKqsMWoxOcLRdqb6eq2DKd+ZsgLNupSDgo4yKsx
tjJGyuNnQKLW2oTz2oYC0TQI14Jc5fRvT08s2qHKHTW+066jX8MGwl45cj3+rFlOB+XH8W0JYBQb
xEwtdgZQ4L7K4hJr3OB78jh1d0cf9Gt4nuSLXFOr21bghjmIpl9PtrT1c8YVsCdLLCvO2BO+u/9T
OhIv4OAhef3OIksjuoz4fY0Qwm0SxDL/ZV7h/SgGoV9ZHLcUFhYMa+KE1ybr42rAYapi+2uuvcVu
A8SpWmtZTcSygX5zr8yDN+BNeq15yuTxC9h5Q7VWlJHlrYjjdihCYBNFBAMJNLCBfzurJRefuQTs
QVxOkcH1ORKsX+jNWfjj5a40EcqSb7exECPxUgWGDZMMHf29OgwQi1eYsiJpS0Lx17XwMCozzp1F
Bp3Lkes0+ekI77TRutYNRfWIOY3sHiFCmPTL21OfV42yJxdKghAPcb3R39bPlFcazijyNDMnC6ou
yQgjUxvgs6wUjMiWuHhTtYMlRnVlES6SHxX50EwmmnQd0j9HLnC9efYNc5GgGgrJGwWsqyEcSzPd
tYkxV9BD7wGIZ0nZLQqglqWlsd/K3ksjekCpJEYxrqnnUlpNWnDPixkjR/+z8JapwH3XZ9sRlG6L
ZcAoh1SJW5I1rtoIsmVMlzIRqrIdGnEl8nQkg1n7U173cECmX8zqj5ibOZfpTtR2k0PvHk/HB0YC
OmpRnRLlpdsWaTp/9zug1Mt1mv4KbmsKuxcC4IuQa6GZLDzBf60GzK6TJobkOKOUJtHzU5tcd0+A
q8i2z7/keeyNXgyrZ+tkGAWOOtreG3Qyo8K/izfqdiWbcc4LQeBms2xQH/VM1nw9JDfNVU6BXKz4
sgh2qFYJBoLCWZ4pNT9kgd9ncIImYkeyeKg8lcJPSDryvPSeuZGPJrzTsKeJZNn4n1P+G1jjMYuR
b+ey/Hnz/2A3QR1OW0BV6+gIE6C8S02d3zACjmQgS0g36fxCqDx7B64PNVhdGV001aGrzIBy51D1
jPAT6SV6GRoxR1RCFFKg2j+UE/N/Fq8MvA4D/nUTnzSP80qRHooMvQ1D4f1bd3H3yNUgjUpTKWx1
dt6VUfhNyzS/Wxs8ohBD+natBNOoScxIKY6oLnBFcb121gEO9JuUfpcZOfLUoU0Uirks3sbtMPNv
YXw20AZ1CdzaYpQVeB2sxET/FkcoZfnnr8t92UXdL21cypqOpSBZMTZsg3oVpLX0ZbFyN8JRDmA3
5dVpsgSJNeRrtG9ZhZWiT6Zy+RS0My1gK2af+CVQD+ahm6mga/g7FrQQ2MTX9pOhJJ1w+oAgkRYU
g1vulNjkz8pUnp4ok7WJfs/u+vugiWkjomAmLgl0490YJaUJsbKlfYIZkI7BIGW3luJ51NnvvTxg
P0T2Z0lZewZmYsR49TQ0SYiaRSIMe/P6DcQnJct1FZ20d78SkqdBtV7kH4ulkylcE/YwMdtFZqf5
8zHXHWG3OEZxqD62VTqI0fzxTu3HYZtiIzYOuxkRyW7ZnZ3Kt54jcugCvbkIZSkDOWUUXt1nimLQ
ojnqkV+YeJcGQsAfKlNFn0XCBY9adKkw7tM9JKFzinMNiVslws9AWSo7kGve1m0p20nrguWL1a8n
XQJcv6Nj6bwXVZfuiOzwdjghKt/knqKuYH481bHMfnF1JroMj0/t/G0hOIcBtXn9zUVrAjx9pA/9
TMKKQeWi06FBD5vCE+OkOGYiCp7oL+kyHL7ZjwS753GEpYzsZqukqs/mRLKW4sTxa0C3h9h2aAbu
rCOL2gtzdm/uW8TKF2IUCCmaKGNEmqoHEAlCql43LHm9MGgWAT6rOBxp6OD/uDCIBJ+qL1oEa75I
J0AsQkro5SicW8bR1TGRWY+ysrBlRHqvWLgX1QqZMX9VdWFbXRoc8DNGZHhKdVLd3SR2q8Jjrr+2
ayt1maTctkjTmLeogm0O1tBXXJ6eNJ9xcoM29W5AkXNaeoKXp41f0jlNMNbDGhf1o1kqIuPxKWYb
bE7kj8mQKixu2TOJdelwoY53fdwBQQKEJuqeM8K5MaBhbfwKmwitdOIAhKLOBaQfXDqKFbjfm4pB
MzgBm0428v2geP3k12Q0nERipcOkuXEHK4CpGwQEaj53BbYHPK9VvC7UeWavmyNGQCFXCNF4avVK
/76bsk2T8vBhpUcMrJnQFaP37VHh0yb4+t/MSisJuglp9xt6yhAEji2cTWtReGLBSSLofwuusby7
a3+WJSh2qyx6aGt+5c9K02qqrHW/Cz4QFYxU5xsIkhalUSpkmgaHuormcqbNY3Qv1w8CJHQCHcId
rF6kECwH1spcZVWOEKQguYz0sGo2U8Rbgc5eErwAKUCjINKT3iW1PDkWRAmb2KNgDkCKLKyk8urs
rDjUSIX0UPpRhDsch+uL3GXqHyFsJHz5s+8K0v2wlJlzs3rakog5OECg7b1E0q30VGyoX7GNhuln
bzQxfGQbXBz45Q7aGBi5j8JQ6OsSr1yExlCH28+Vr2XxrKyOeyzv1BXL8rYWZ5KQVXZh4a3nfI82
l9zDcOIhQbuTiL7j7LGyndLipHGM22vPnEoWMptPIy7Jt/HVYKIWsBU7IKYbKZrBub7KKnBEXjlH
A58v2mnttt8iTtc5VhX6bOftcP+VCySN8unYAs8hnmWrKVeLiWeL4ZiEBwLxJ+1nAM5/xB6yW4Fz
2ZepfHpPvJKrRDEoQ3X4Nu8/eRlOU0AgDVXBkb9uGtXwYiFk9EW+rXZcUZ4Fg6m0xdniwdyp+BlI
8lwTfatPF1O8ZeYbDh/AOqLCq0TlfT+PBipMnz/w9zL1nAjUAauCTz3DlBNLzoBHTQpru+f4PA7M
m7E+Qj/ih2aWm8I+TUC5PIKAtkE7GvHSyiKxqyugptCxjquJPNvDh7nHD3i33BvdoMZLJ5M/APPQ
GuNZKrqoEPdkTp0rZGEGcLDrcMurgaFmU8SA9SK1jjb6VKLvlKCgt8AHmlKFdYmoSnqYOU3rGnY2
3CKhSsJhhrUDp8eUNs7UkfX+LAdhS+JvEUO6Vo/3HdU6hL1SbDUlbunMN6xQbm0m2g2DswaOwbuL
UWfgwafS2dSmuod1wwya3QiFTgsoLCsRk6kugKHg87PTvuOZcZTQUKjQL8C+/0uz9ZZ9EsEKDovr
I1tYDCNNcHEJTqGCdnS8Ase2MG1KaFKUW7/A6QGrCuk6zDJ5r7TzWYz61o8/9e/4DaiXl3QK/AaI
R31lyG7QxfU63SrVxr02Prpjq8NuVj8qrO3c+Sp9Oe+G2X8TirTukMA0r2p8eFTQ3mMTMlKUrv6r
WDTbLoTVROB819Ff0ZR9QyRY9RyfmykazdUC8Gs02lqhCYYdMwMO+1lY6k0/WvIcPCnO9frOGRqB
7L1fSyWmjTzFPN3e/SB4abwUzHMeDVfPqo61csG15uYCKhNp5WRy49+Gwd6JeZviXNNTi5J2xuej
aDJu1xfb7fW0qr5gxqBzEt4qOcfwvR0dHYF/IFlKUSBP/U46OMa54YGTAsiWibrmHFXs6731zwk7
mkFsRJ2zzYPQirg1sdk1JRshdl3Ez621VWgryQVtLq8kM+5e/BbWfYfCEtOTdqbowrQa8iCr5qkQ
xQkxp5urDLWC/ChEWQZc4bJTm1i8tuZ4UMmuYkEaTxDaYPZKA5zUNJsWeeMZnxz3QElhQN0Pv45Q
O5+9bxQ/1x0WeELCziqY9IEtcREtIj4QFNr3Or6GV1G3Cwf3EHzjT50OpnM4bnwdb5Etu6XHyiQp
t7ZolSUBHdivebMnKjTI2amD8k3KRlcDClGNrXEN0K6Q13MuIPOChHLlVDIZJ0sh1yVNtzepyqI4
z9ueG8LLcW46FkvO//hIpS51wnD8LkNXnfKSw+rez5ci6qQxE6WjpV1NC3a1P4pf8/GKIEfrpSpo
EWZQ9LZyXaSV9NPiEFY/dPoCGO7nf0WuxGaA8t5tkQGW0GZv2ge/81n3bKlsiIDMCq9ck069pJwv
GvsQpZLUf0iVeXVtI4mZGGYOTO/fGLx8nr4Nvq3BeUMEF8wTOLc/zO47yyJzurXO/QX/fqGKj+4H
GI9cgqjBkuPzdW26U5qmm/M7oIxrudYzTgJH38j+/mNpURp2jrYWvXWXZRuXvcoWLWj70tNpiGuh
OKeJ3KXa0zUiU2y3o2NNpTKuTbzqJC9p1SNLBjRpoA40aMUBNUrTcdeNVEGwiZIVC1Hfe6aiX+Fn
r1rEJhprWbNuydd/eRnuA5SIx84PFALkvOd0uOU9Er0rYZxW/YBLL7hyTUbflxEjXqyu56FT9At0
tLxHUg+MMYq1BKvTpuvKhMX59cfkmFd6ENZu347cfVGwKfijOlgwlyPQlz/1sYURTCdZCeNl/LFv
Nn+PZIcS9jdqRiLpyHzr2REEIIFtaakKO1aPuJA10dWX1IQihrXYU7/UzCJEXbHK5sNUbti7tSzG
fdwi5K6ukZXIfmJSMsvu+ws96X8MK0KjRd07kGOASVixIPbnB3Rkqm8o+MZXDQPiX8w1Q+qT4trx
p2Q5mNpkDNVeie4lPJD+6FZJTtzGY8/R+NhBDCjYkQqbt9dONSxoNA/L8MR7k48jvHISucKAO3kx
H5oFLRci3ZSPJa4W4gyrTzENxlQUut0IP1UQ89XuoVutRdxiwhlsrXsfk1+gpDqG2wVBYCDd0iZM
/skKBYXYC2fS8uZWt70UH5q2KBlfH461tVGqDeSTRCeZ7/4U5E7dTCEnsgWxZAndohQUpjk3LN85
UUVMYj18UNTaFEmXMCEMDRKll8qaPcm74Gx60gSCkUXB6vaBSG1Fg12ure7nRdgR0VZU9w+a7CN+
tjq/wNTCORWXuUo1axxd26zzJ/xIpw/h2XjA19TngdwiqUiSr/5knO2V1sE4a5oQWKC+Sz0BousW
QV4z/xLBGjpzibe1wfhq0kXQRBZzdMQ/qDrXx2LaRbzUGTNFtowLrGciZ5OQqphV9yldLTFZMT6u
tuUpboCzzZj9MDthV6vsXYczeGMJxnFRaZrZSDJurtLvr0VRXD3UUu4ORVLQlC8XNSBgMq2HywKe
3jii9PDvYsHrZ5yGvC478CcWes+5Xpu6UVC4oD7LK7VpqHyHiNWU8UNcMsKHAJXy+tsMqtXfsqxe
SRsL7d8GesjrOVbV+oxnz42MH3ADpAdYJfwKGiHiv+xqpPxIcXfScR76lED5OtOSAig3J1jFrifj
MfzLzab8/JO4Ss+Wz7IIVYf+M+bzLAvooS4pSvpIUUuV4rAaa9VcgJqI1swG6/MSkWnNftfIJblr
jrkfAot+jhuVY2FgvoK/V8FzCLF0c7zxpVKCXPWRvVv/nE8PCAWc01nZY+dMVYmzEIyQ9U6ly6wt
01KRsiScHzKUqh3bAgdMKtBBGCdcjzP52/9OWQvZTB8MZUJ8peLChoEn93XQz74ZWmVpP37Ej/mQ
NNskx9hwPQ1fCk68hUXsqhpyP5jKJubAuZsrt3LSbFYbfE44GFt36ZYOHO8SbnfMyQAbMBPglR9u
TgYJTGev/AiplbgE1YtqQl1ijnsb7I6HZVu2TW8C4wIuu42lIeY8jwLBp/ei2WCSwnJGW8NHhs6T
jxfuFH5rthncYXPcWeTt17zOLkZVZeQbrXUZy4ge+jxOYKXttnHQCnRhL3jNkSrN1advtwZeOLTN
g3gXS0Nd0u2CMiDRrecKF8+W7Y4/9QOC9wy62U83hvlVg6kCQBchoHfWlWtUqTGHh0ZmQ8wDwt4v
rgMyQTem6jyPVPCmgWP8cUVNyCzHK6hOFH2rxGhYsZXwy9TvgZ6LhC1B/Ce9vq7zbHpTW7wpwP/D
7J4Tvz6heyvbG0iBbTJZwYSKfVVfQwRcH1m7+bMr86KGO6pHrIZqDXBzltpzA6dgkpfn+Vfv96Sf
0OuaLCurKbyKe1dof178zl/H0GczIm3ZzmkYUOjyjFXxeSkp4Ip2/Xx/otvt9rsTYymGXekCJeqN
S1FY13u48dUs95u6ISFppIfeE4NeuxtECTn8Ccm/3NXryMckzdzIjePmKUObcWIIBQ6ZJ2CWIHQs
o/Sd5ndSNZnAsXXJQaemADd59njQqGkZQS/O9bRSK+JWEzCa2tcpOGYvDeNcE6iWvSXOzq1XFdGV
H2How3sEyHdHLBReH+dxCRRw3Iy4urTm/ZGV7ec6j23dZNBpWibXyzVL3oNiAypf+K/U+iRKJxbp
ZUzHhe6PEGygHNwpbTRwCN+9emsJ6tZdItLhrmNS6Ub/WwWdFcbtUje50KXkQb/c+n/3Y7kgRwzV
C6L3aZGqv1+ufUOA2Ij1gjnmj6Ec2rcP67huFtIvNb3ZyehBLJhamJmyx00tdlmBnHdZrVyKROfR
DAHAxk8cC4GLePEDMDGfwXykKBBGbJOHNqAzO1fG3lt0nRQgv2JFq2Yh5EMbYIzNtVn+mIWk1Jw2
PWRSXOb/msWCnxCDpHomOWSqC5U/MuP33kfVIvnq2mtHU4An2kMrXM+cXsQaS1ppTwZbS74Sn4QR
QETa7MnjsHB+MT7SlOcXKJiqBifQH6vFB8BVPrCvX3y+4NCruezaqfgaceq2R8I58rXA54JfZWRd
Vscds59H/WyZxqbBooIwU0VtzrkiwQJotSvRyya+tL8CRcLu2irIqjoanO01Fenj0w2esk5G6IZH
aMHzks2CVvL7QbqY1h/xFmdGTd8UnHvOCn/zDJVxAz5XWqwGhuN/ZcSGhzxVs1X6VaQ1scXeHyfG
74cz5JuRJOkm97zmDJVREHnst6pjwQUv1FowG/lBuJ+5y/x+5dt5os3ubPBUu677TCUzRJ2BUyKx
TXcQtsPkLQ+YBsbJFTniuxewVrW9/kUKsHCXHjbLVS7CyEoOkOwtBRSImHs1/5NkcxcpZCLNlgbc
EAOEQB+64EToBmWlc3X30ilLtZ8RG1R72WOKCIVFkOApOOVO4ubZ9OS6cO3xbg8IzTGJO1Wq7bBk
p9ES5NjzSm79yDiuwKe1HtYTv1JkEdKOkVwojLIUhQh0qHdOUpzdV7f6WM4tAxIbOokIj2V4h3Kj
3F4PqfGTYIy+2VLoDK0g1Ut9su8VNalnSJK1AEdXuxW62OFWwHTSNMqq53XM/TgXl3plVs05v6hd
SBtsQKLs6M59gzIRWcPENMhYkalupugMWZXr4zjI+xTb3O/56EI3j9K+vZfWrfGR0HeT9/SZReFn
i9Rs8COc5kRFPyPdbAepdK/cQfkyzUrgUiynW///AjdSdx5evyN+o5t9LrTkRpFB7knYpJuTb1aj
miGo3Tl9SYDTupgxt/EVJV/DdRe18hs9cGXjA9lVwjJ+Av90TkID1BT160memkkQJQ7q5yeAs5GO
+2dyPRFtGfyV76kN690qoQrAJhFMlRf21VsMyV1GKGXwJSNYip1tZkO6JNDvRFSOhvAOqlXSoQUL
p9Ps09FvWq3T7qni1kMFVt1lFsuQiQ8gZp2mAoqM6N/zzNJb1FqYkXlr94VB2w/9AiluCrizh8Gy
ImEGXXeN2LaHIn9B8ggceBwiY7TC9r1vafKY2LVkTwoueiKCjr1E/uPmsVcuKX001sr/MQ0ihIVs
1b/1XB+QrWL+yqWUquQcL6CWm6Q9/rUcXw6iHRuxcLWRqoHROChfBNe35PYaFXxqmNPtYL44rPVA
iTlGPEHLqi+neRrDPTMHFZ7oVD94L/z1zKu9jmtMwi73/7EjzSBnJFfXXLKSPbNW0uVtIBA3gs8S
CehT1SXxYOKLVmiECAljLjemmdacEN7Gmm0P3B75QTnWg1kpIB3VaZD+WSvVdNNMo1d71z5Y2sFo
q0ssKncZPq8GDofc+qbnNdcTGWF2Ky+8nsuLcoklBFnosHz1eJnrDswpkC3rUEFOSiI3fMUvu8Vz
cGjGV8kE3M69YQJ6zxbPk+Be3SfvXnW68r+PooA5Ca54CNOChJn6F+pViBmzW8dvNaFrCbqYxlMw
tU0PjFrMO3PwDQlYCGiLCP7ATJZXtrThyXyLflI4AQZa1alrpPp37oUgJX1SN9bgGljpNlEfbG4v
l06ejg3s16CcdeXMuHxi0xLKxA5NvDoqQ1UqEcKYGgK8Y/KwaZegZb6a0x/sFrusNDEradf+crP8
pZD/hexyYCbh9wX1w7TR09xUySV245cobij/53qrUXZ8AYdfAKrvfbelC+0/t7VHEO95DprILIDn
k88hPPtNcygTKHuFh12FEiRIYTdSH3o04vJPnRnqVuOhlUtoq8hZW3y2xuII9ukxe5LYdPWGsfaX
xPJ+lDmbz9Qf2xL89YMVXKkfVkKMIcBY98AEQDFbcttdBWFhWSiJcmFnQTU7Zsb266DJXS/PmgTJ
l3a1e0X3M+aCM2F7vk4VDxnbLiIaJPnwfgnzV1jHjOTLNX5Wjv2ARkJmT7wnEJ/FN4sOzKKuhjBT
KPIBuO169ssr4BpJQtcQpJeBW/KgIO7ZExKkEDtk3/MGTyJS93DY2iYEuQN/19CJShQbMBphftsA
eoorCP9VbJp1o4/u1V2oyOLUQp+H9a2nMs3LcyZ2uTlvSdYoLKLC2wzAlCd2fJPHCoapOf4YcGOQ
ZE7I7jFyBZjqryQn5JHxd+N6q9F2KTkupGpgK7ctDaZEi+H4y5pCgctlLt/ZHO8Nu+mikfE3hp34
Dp2G2Q1TmfN8dtSufcHwBxUQsZxtp3HW5y/J+Cd7qnwQ1KxrlCSz9vYzkraVQQE01Y9RF0edRXXv
tFta5qXbdaF0CQARXEaA9aW/uxYt3l9CAUPVaGIRqBPqIqbiskTrxT9wx2GCZHqpulnDd/v5IQgg
083gVYKGEeZgsyNrjx5Fa6DVGoZ0BLYCqd8fqwyccfJmLvWFZRe1lk0sBhlnwezSjwxotXSfLbJw
ylqa/1d9Z/KA/vQ4XmU/jJ+PAuhlK6QyO7HmxmA2UMk2oa0iGxzRKFFj39XciM2R9iYTsCArsNHB
suk5xH2syPfKat65WoD9M9vdF31D0LVbnyzQvCribhfA1zLy+AhTuMte/gJ3CGSAbO09/+3RCCVd
b3qoH8botOqPx12bQ0KL1pWqlN02C56Vyf4Mo/0OwoOjv104jqFIkmr+MT3GW2j90RHGyJWuSUGZ
Va3YxxdrN3ZlpFJrydCtz2kYRjMc4nKns1OcTHGH6WHeYPOLiKx7wrsO+1uSO4PMxAhWpFspygEw
yQEMa7zTOID4Mcaxf7o0wyeYdhYRIAkmF4kkY+dfk0UGu65VTvZImaDVTJILfPHTC2+czs0V2tcy
0n3vpenNI4YKyS8QBWR4PFGNL+OMb9Py+wG/0sqSuuswIOgA3m7z+5X6p3mJ0fekbfBVtbQHC9kV
i6K/Ce2O0eVPDcsEMC5hzeYkHBy6ozlgjschUFHTbMoTFb0czB39EFYq5YKE9LsRr86t48yDIC+H
WSGNUuI8sU2judsDPvRXxZXfsAs0KgDeut9VnNl4C1oJteQhxtJNr+jEFa1UFfA7qEr1SivuB+0G
nYW5dfaEGw84xC0WuuS51xtpC8Zq2D8G21kebtyJKpMZiqN9wjhjlHjrOct0Yk1wZ6ATkAR83YhV
R/oPbxZ6CYYq6LLTPZzNYoZOhl+ZBoV8HgqY/Esui8enX9syYLc9Nw0MbaqhtWuL7UcJmw99+kNA
9mKxTiJZNoYIaDVDbXZ1CIOLeTucuwJztS+jD25e4ZCKn0IKdsKj6fO8D4PDIYp5JYTXd1fIs1aD
lQzRbV/FUC6dgo71DNhKEUaff3SXKwxUhH+19BdKdhq1RW93FyfoWYQwqJ2z60y2OBPmEje9sEK8
U0ImtoYbobxYcaBnkAxfkuQJUEeqvcGAjQDxV0Nwc1VymlEJuwOUD99nhBgxNfb7qT/yD7Mos0ps
YekyD2MzczrbvSZPVlN+Wk8X7ct0xZW6bPsrrYb1aRu5x3voNlR4zmLgsoKsDboU7blKGmGtgd7S
UQHVSAEs0phbFs5EjquRBMGlNNfREFs2847GAMQh2eWfSMzbHxF5f2X7mgfhSvlRu3CjPs0iRsO2
+u+zQcg6b/1jCkb4zR+KTzpBx4sEA3Yk9A/z1YZVUpEre3IoWTni0az4s+hRoflA3pZAAPJYf4H8
1udJVayAmjf5FBomlOUL9gfhSknjgQq7n5CYvxLlPa5JG+ExCDpQJodu7tHlfQXSgGX1Y+I361ZF
Dh5N6PtRUed5id1xiszl6pYDfepPSy6jmRGWZ9jf1DQKBFzLjXmPrh1DrWL3T13vzjbGyYvtziR6
ZyU+2wMdcUBJoEBFrOKL5WyarXLcQefTPN4PToTQDzTf6Mi7HtKLhJxYmHtl/uI6CzCsbTSUI5im
nOhZW3EJuaZZokhN7H4AB9YwNbNfxeYuf6CwQLr5mt/5V/rXuxiu68Ek8QPvZxl+J2O+ztlPMZbc
Ieiu98PHkDVFGIBVZT8Evb8vsDfSwqVpnAjEeWMkVSCaic4RSLwnZUIf+BcRAJyZ+NqZWr/q474v
GNydgfR9FQru34cC2Mlty7zYY3yeAFflncUKIXr1c8y26YoW9fpjTQPGv3CPmTg6DIo3YkyA39qX
rsq3Di2SoCbXA/JNLF9ZMLxhvXAqRAvYcnTFYSrd6VSUgCWwgSg+Wozzq9MMkQHDejgyH8KvcEcL
Ux5DvT9oN6qK6iUy17HcRVsj3utOyktc7ad24CwZwhL+vPl0Ny4hsMmk2iUwCzU2xCJk2rIpdxar
o3iBSvxP0F8NyB4HZslGhp6ueheNZpsxSE4G0GkwOee/Q8G82QX14j3OLC9gi1sR42Tq2XxvFqrZ
aYehe8zqH49/+zscGa11p9kCWpUuJLhVhbXWUqU9cZWguJzlGVbQAfxu2Ucgz/N4hlLgJ1grRDfU
tce1V23VP8pPNFNIEERS8b0ChQi/c50oGZJmlZ2nJpGOcrVVTrik4rmIB2IdOOZYNvvBRxoq285T
YGiMh18ScILx3RJFfaiijFhh+SdCOTTW8lVxVwhLWVV0axf/qtr4k5O/Ahqe6SfvNzwcTzD6Mr+M
PaBuu9KmfQO5xp5Kw1ZtJto3wbvbTF8A7sBtK+We0fzMVWHF3MNDMrOZuzbw6WvjnxFhDq+W0ivk
PLLPvJXyOKgMbEVfALdSuJyF+5PrXh4Yl/MN/dkl2mpl8vKOUFiS943D1rPWcjRtRhq41ozKOPpR
eLq7kvchZFN34TOgnNSXddmTwomVVmmcjH9AC+Ll12RMR2Mj3LoPAO0AnVpY3sz5KwQmmN71D2cJ
acY5N3nHy3qMUj2FiUWsmPuEK3AKZiEPquwwpWLbMkpQ1zM0kZ5sG22MhbVkwrTWTLKc6ORoJFh6
VLIKEmbMYDniEwYigBxNXIrrauG7/SKvEI5CRivq9dv7skGcIwV8zbwHqZykKaevChd1Y3Lj8Ci9
uJ7a0jRVVaB2lAPzSXE1sPuEeX6Xcu7M0r/icR/AhGPBiXtcoH/IEWCBuQrBFWpmHjx8jJFAO5kX
RzDO4V1ZQKdqJn7beQQI6JVNvD3JMeHAtcPUBF2lHwIw4botHhJIUI41mXCypO9KRezQ1jtowFx0
PBkHwQurOATQb4f1OLDnm6IYLcDCWiHJC0wq1+I5QmqjOflbLa8s2Pyv3i5c3dDAjZ1Erf8359Lw
sQPopj0qq2D+CA+Q+a5i3YIfwJJdIJQhDoeYLyBNZJSp/4E3OOMOszxXy6STXYfUhznfkh2cPees
ALeBHsUUQ1w5QTx2lbsfS25X5cmKs9T3aE2QJkVHo19Qzrim080Cc/PtCiBx4TiuDz8Ld/tGFE2N
5430qsPoheTK2bThvezFliXq1+fCjRzmXAkVOj8QNVRKqP6jSxiS0ju3XYZn4y4JU8Ozfhu8SUXQ
yl3PI1tdZP749KMmnvLKMnAlvcVZprLefo5AzVgljKNxycMHM2jXlQ1cT1N5HVRkldXA3H3873CV
fjNrU5XWtcRR8DSM0seUE65m3R1durtSC7iYxGC/jW2L6GxlPCTwg1acslCcj/nFvzh8P8cPr5Rb
vGyKtj5JyysU/hLehvpQMPL4kCthl+VFJrvJJj9uPLUS1SdaHUenDgZGJIUh9eewRawYK4nWL4HM
zYWVAwyPKTf2ZfmRRNQNneNWjAbISQDLJ4EwXvX5kHduu12qXWz8W9fcPkgAhmXZmSpDd4++bjeE
BhmFAWtdKYaDVuP63JRsCDDC4+23Ge7pSJyeYZbQC/antEH7zsLvR/+dcElqU3syTaIZpFK42pFD
/FQFxI+grNOgQUR5KliE2TbpSZHobTlMSRteO4mzqg2ULL7kqjijKvVYYSQ3gU3I/VoK91unHyEu
vPo/+YiAA5aFZK1275sl56D4aZjVEPcecxt8A9AntJH6g9j9SjV3b6q2jDRrI9V/5ZlBkILUHC5H
31gL3r7UeRvxh2nL9/xhOUCot3gOn3nF71t2J+cUKLksgvOpqXeRpE3KgKWiGYrd7mcDrCkIYm+5
IP8KFG98BuuNeKhqiN38wmK8KXK8uF9LJut8drMJ2RMoqsPSRfaoxv2SAMulyWjjeVWrbnmLiVB9
chJi0A0v2Mml1HkFJ/LQSJ1UX65AHdArTrYgw/qt5WGpVnuWuA1uTT1jvyKB1kbaYppSdQuQQxia
inYnBo5KDUTyXyJt2AANmyBV8boiWuN9CNQ8yjtiK98=
`protect end_protected

