

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DYkUg37UnVRJ+X5v5iFDmCWObMw/mUCrJuxa/Cr9wGl4FgcJi6OQesLI1M+aH7+emQJssoNWrh+N
iL9trwbpEg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vb74X6mc2H0e6MLiEAhBKZ84QSTgHhg3aAfwLeb5H8AGScZ7UqNDKDmI5IhuJ/LPpdHQCtOent5+
I1p5tELHTH0LzN6BILTKGZBdaGJ2AKKoofyljqaR51srCF/ZJLUOrn1XUZMkdlutYXGikghh+zK5
6+/HFEYyz6zhpfFGpAE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DUY8u9eRLqeXCDG4E2/8OtDIacK06AysbSio1XfMMKnofNQFNkb8eAjngrn4u/YZ6G16ZNMG7YoY
jk2Rx2Q3M5GrNkHLNcW1r1FM93KBIPYna3s3UsOdPXI8u/gdrTwtTwv/xpFT5pO5KUummozg1ol2
CfVK4phP0ptL6RF00qSF6IA3NotRdVSf39i8Abyti2fNqAeVQtQbe8y1/1WV9RrHHqEjarv5sqIY
6GslwJ8wdJjPL0QS11gBEh6rDpndqUhWIIFTUrFMd1tEU2WzUCNSxtbBPYlWfpU8e4/l9e5xSsF6
weW3wzZvwjgR473vdWcupdpbpXFjQjfOA39+/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
p0GGQgjzPW+6PIUsMdZXTQnjW6BUopNyvt7ApHmGMwjrt0lKkYFdeq6NnHPNeKi9xrrloGAO2Tha
FhPoK1WSUQvFoRR4uKVUk0OywXYhciTgYL90XL5T7z6pvP+T2xdoDnAiUPoqzH/Ubhhi84EoGyo2
+zIDCCcTvvnznOBjfpk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m1/kaqW4ETEcDTOeEJMS5yQHRelnhe+7sXgpcKiP6lTf8NZHj87LtgfMx1Oh7TGMtL3OsgLwXKl5
B/MVSSTPV7z0P/OvFd/MWYJqIMAVI0yV4hJ8dwWC7KK/kawdL1h0Q4iS0dxjn9/392LJCmqkJJmj
TEThXH1uoH4tMKV7xRRg0/MNNOk8hPErcV0Sx7ZxMFsvJk/PuOEi0wzy6daa+A+gop4M475HPjAb
iPZ63o2focv37v9R+NETZc+LyDzZAZPFDxIiHCnZlRMpU+rYc4lLu+Wj7afASerzvuIcVvlJO0R8
MuDtSunchT2Nxfc8io8WUTVsWpkmP/zQb3BvSQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18992)
`protect data_block
Vtx8XMnAZmKOz6NrvpVC0UddFRh50gcfKxZm09IBdqQjytQLz9g89t4Op8wwDdFWzTYrPQzyvcZ4
nRT08FkcgsHeOxIAck6svcrAzILGdFJSUXYn7tA+LKNBkb7mBWy11vBOpyFuj5nBcOGJ38di8G8Y
zAe1YRT2Vd+bDjZmgENftqSPVMAfH6NeGiKtn0mPelPEr6TCr7q56OK1h57KRKkRNVepME3lpgL9
m5hpkBfa85WYX4h1nW/w021S5tbjbLpnqbPMTwSwOV96Wm+kZWYErCfmU8h1L43p4sD7TSxiZXCQ
GnlVpNppN9qwY1g/MvF+LeAUjHVm6Q5PNsfdrl6Gha48OjNV5asUFdbwCb/1tRjqrsgcdCT5FUNu
YF+zDtuZ9dEGQaK92WxzMC9Wm/xefP8Tjy85A3uRvSY76I6X1gZn7YymTFgzW1VJD+QIg8s8d/S3
64dmsxRZOK3TSYaUUrgDcEidFGBaJXSDFLyX2V7NR9+EisH9pA3pVclb503HxiPIzwFcRdTF+U3X
kSLR7vyvsCOnY8QOfP8AECXHHC0neU3DXvdK6+WPnC6qiDbl14S8jR3CjL/7cQ3QkFoGsOCgQOYG
6LhHlHs2/EV8fK6/bN7dDT2LuuGWVZlwWuj/EE44xcQ2VNaLo3y5FwkoyDKyWU2+SV8h13AwYA70
ZibVed1a462b0TeeKkaYfxQkwh79QjD7oUT4KJd4c6TxfHcw8w2ACuRvo19K5W0yxu8VdfP0pDwN
RPL5XTyTVAK0zEjWSPM5RVUP+skg9y+pl3YKvoqWKqm+hlibmHyCLjJHQucIuE44SALt2GmT1RLD
Vc5JMeS//eCoKWU8YsYbIBo4s2YJNSvkWq0ppzOpve4XfkmTIC/eZFDauSHcc/kTQdivLxF5vdMz
m8JMer9l3fLJrFVHIxTTNBAhYHWdoeRI3Ul+JIJbOwiu9NbWjp0FnSgFPYdwZyJapELH5uhwELSQ
M2gXvslTR9KrbhbV78FFWm5UOOGE7nF88fbDbzVXAnO3FO9I+JMaMmMnX1s3aqAlKlGV2FIAmXr2
u9iK/kQpxbKK6CcpDevMMHBI89jc/mrmNxaL3TR2tmG+x4JHe4tCzWGOlnyisqQHG4twXww3frBx
wGl/e+cGtBgEyc4jqRxNdmt+Dc34bxiWV7v2IepLj2aWvb3c0mviNyyWcT9qUViodw91NsTLYehd
Gj7mf+hePH8EqUMjH0Ef77CRdNA0nYRIFGBlpr8waQyiLqHJ7hDKTup0+PXKbxK6HQtRUN4ig35n
ZALqy5ybxXiTyyPRX1wbP55KZlSQgl55Xg+VCkGm6NC6HZUFDl5S3m3++uGIGujzSthbaRvjarm5
j8nsnrqyGtqj60tlXCYuFKudNx5BnvgMrHiyUCxKjlUHuroHcxB6GrM24sZ4ALmLqAOTnNu1dkZM
5Y02silx6FWht0mZBlP45jdIzjHpFedHCkcwRzVNs4d65dBCqINwLtiL8xiJ6w8fVetY+Zi1NadI
V+RMTGTydH/x9ZrQvcrGTfqJgNQAxAmuq4oSAmHJGfsYviA7OhNJWfub4J+b3cXKBqgY+C9b5Djw
tgu6CdL30tK2YEroYh/yLH3DJBC3SW2rzgWHnf5pHNE1nSMAADsPB6At8ApXHFjkcPZpiX5RH0DP
BEKHGqYIPXLVYDnTHYDq1J9EvHV9Gh9AC7aKXHmAUfOqTntRJBJ00xb7PGcpzVkh67OsurUciBAt
1W9oiFCs1MC4j3SVAarWcT03kJefkOd6IqnPzLaDn82rASjGNhmbMFAEgiHhLHn/ZXz0oLTPSiGM
68rzeRchkUvHQY9FZhMElI1z0+4ct0Dwdf1yPbEJck8/V2lNEP4H0OfHer6HVn2sh0XGXTqlXRr7
uJIGYs/XoD6/sLyIhh77/QSmxkNKQHaxr+5LEPbA8hS136kr8G7TxNtYOcAAXCDpXzQ05Ppqr3Fu
LxPNL1WhrEPR04Gs07CwzmRxi6RvmRsXsBCCm+eUyhFa38KwYnANrT7aKHcZhb9Yta52Y6JxSCKG
XSfAkAX5j7AYTIAKn4dCSEzXpAjB0J65Wsb13AquEkAxJbFesVKrFOt/qWueHW2WIJAIFx0HL1/Z
ZUcz66kfiLW3lDq2KEoCSoPsl85vNndjNdiNEueoTFfWbhilL9CFKBC2a2aeWa9ug7Ln4FkEXjvn
7swIBykrXnoQx16nDgtgr63iniqZ9s1az0A2lVBUpC9Lk9lo8W9ODBffTBGLoUA487mIIrXD6VYe
2Ps+hv2F3xLDucWjk3FysxTOzrkUgCLa618CB1BKWJRDBDyoCCuP0olwEG7v0zJKnVMDkYLKdnKj
+wCgOLNGSdWfsMworeOe+WPO6f4tRNrUYNcFeL38tkR8FjFebWOljChe1QOwoIwwT6WgYEaQ/4PG
9jiPOgKWGVoYlLDVCXoWU0WyJ/HKP7xnteEvZ++4p1YMPDghyeP8iGq5hjZnNOtUjmMit+Z+SlkD
JU1+xfiaVUzfWl7JNLAi9ndx2vGOeyIDp3LVZwRc4G9ByfrRuglpDxyh6iM//sqx1ngW7IR5JKJ5
R6goe7pjMu55Vb7dXVfhmFmoI52DzS9NEcRCIzymHJHprfODSBVYUOUxA9IjhuAZAkeHrHsIut36
OWKK/yElyem3MWGYiZDNVVGcYnaMg0iV/t1eEMQP7NqpGYi3sl0N5G/W/ufqQ6qbmXZ1h16Ajf+/
oDrDbg1tTLKsQEsubQh970i0Waar40y0pxrT0NMkPyvGYF583Hpg93g71QGVK0nmocXqfptSSL1a
DoYEg/vqPwRIh2G+TrifjtvtDBJ+mBG5JuaT6VXiOYeJNUBwGqWwFSMNz0bP3IGSkvwGiCsxjB8E
Wtwl0nSnR2U7XibcScpqrJgp7cyk3Xa2Wfvl0iONvMCbkhJg97xFKlRzHo1n41Iaw4N7bGANzj1+
6Z2k57r8Aunko+HNNAd8iAzYTt8LTjeGmAX3SEWV+BIkjeNBWPuvdPnLXp90M1SSKQBAENkD09VL
dAM5RrhAg9Fzi9xS2DETuu51r2Yh7vf46qWppUAIxFdia1wc2QMz+P5jC61dyMdefrRRd09/U0+S
fJhHpJkqZ12BGH7hsnGPiRCPVmnnfv+EhBTeKGbhO2yFqBir3TcgG6yTE/c0RdGuZ5EFRc0QphvH
Y4nZfYCszzcn9a4Y58yoUvCpbNTUPpj/4dwzi8svRN3GKUjqEIUp56/W2A9Oegjdi9PsZiV96bB7
1ithijz4hvHoxZdCLl3ghsXLNOfRn0Dczj/NE5yV7FQai0IEw6p7DjKqwOIHCNDfVgl315bltb4+
gulZk8R3vRuV4uiZeWsqPuVsnZD5tyBkxu2rv6hf6msMIEpUJODoTh+w3tAA2WI/FBZ+JXIXNnJB
dm3eqx+qdTt9WldUTJbA5Co+aP8nKl79jdoqquVfLwHy9oeZV61a1UABchfkOW+WBxwzmnK4Op8v
IQ1RhpfhlFlorOye7G6Ee7nlVj8vaBFIVzEC4xsTPrXreRVZmqN4/xBqmz8dIqfmRVAFw1i82qm5
pceEuHB2wW6A7D6YPBaecu626Dg7wdyyagjUx6umNzObNfMJTm+PMpKU1MZWANWA1rYrGYuGVWh/
WCAUo9FG+6HqwEpQo7VR2r09sBSHgSgyC43hD7YPJkTjkcUcZdXv2IT7Nj4C9uVmtiGDwtyS4m7j
wHdlFY32jmJAvKQacAznxCa2GWvweQ1Mifvb2NLbXZLTbYwubrnMpyZ2hfath+IAI2k96gnHpB4g
leRVR37L38tvNCLwBgGEUx3Z3FTkQKFO29XBx7tGO0n5qdMAAaG6hI/M65JtB8oZe0lC1FkdOoPu
cQZqTtP27CNoHuUzSSsgyWfdl58qXtgSNRQ57Dc72mIdC83zwi/IQurTrcGDIEYKUNFXzCDw0cGu
LZsibXtvIXmLD49XhqspVefNwjdfxubdxFYU2K69EX7V4ohFuj/kX/DxnwGalPaVky0lBIy9VJD4
owLH+Rz16WUWA7MpWjeIRn7v91oul+Te9bN1kBOr8utEcSpX5eEasqn4W/eX5bmp2/qR4SmyRQpP
OQSAAON8L3BxbbTEn1Iv5GkvGbG1styGeoZHtJzY8qupi4PttIsfo25RwlbtTF8W30OUgqNt0rMF
YEjsFL6WM6Tacp3vlb8XD2MP7Tv2kileaZf2hVMpwQB8E5qrBAYkcCfGtsBHeyqa8tQrOYTXjd0f
ySm6MJb9jTE/6h7O9LWzF4oWaWO73IQ+Qc0RaPtq/gT8dYUNT/KRB0OMZBYufhZytr1OTa82E0at
A97VZYq6BahMZwOtukQN9dQ0gaogTINQF4h0vp7yEjJd4BFBiTFP9wZyrf6SMCT7w3N38Kmmjw9J
UeIM72pa6reb6u3VaQiOrDFnx+gjsrpcVKiVtbXkU0gkD6KitzmXxOKAMl0FoswvitqaqLKmiUH0
j7ojQfoNo+4VghThvQ9TWNeqvaOArBaDl53BSdh3JJWrO2D7iQVwlOow8XoM0OB+idlQ5eJ8rAa8
lvFmYF5sEK8/E32SMLf8UIFoUp/QGjdSENzbS0CwrwWcAwsjSD/b4LWjcjcM/SnA7FAIUmM0XnjF
C11V2E5lTlhXLiOJxDKU6MJauMqcg48ihW2KdnIhsmhZzgxliK19u78uj66djcOyg3YUdqiAnfN1
SMipOxiOc3o15i/060dgucEeUROlIut81NYMRchBDDnD2LLcfq7TBUaVbrzWuzBXp0VTxG/utFEf
1T63s9yWPZ0nuFBMIF5qfu0hD2Jzz/0uEvRVK9AE1McrUCXiZFzdxqLXr8DdbpSZ0rWXsNqVNeYm
cvXXcydRywlONkIDXAbTvWaM9JNAMPx/MUnYDkCWSAV2g1Ph4yOagUTt/BKrE5nYWHHni2QTI5AW
oN3MT7G8AmK08GIfgTkHYc5Wi2V8CLIBjJZi6T9mQ9rZsVei6su7exy/EBpkd/ZNfket2bXqEkhn
13uHe4DqWykjoNEXpPMp5Jv6Th6TasaGXuytUWet/75utyjPBxrllZ10k0QRmDGvSK4JtdqXr1Zd
LArzs2V3xdxxcyTRtU7sK7GQtXMXwIjc/hHT2TOsDStfi0LaRYMGoLcFFP3wqCV06cBh5jiYsgFv
RM2jDDY3zxH+CiR/GQNyzB+c4aDJMSqX6AN0wqUEyLeg0upBgYZXQCNJrBhjj1jnMZTY57nDgLXj
w6fMaQXql8G1BTrsAbmg9iE+iyPE6+KGFapsd9CfL8EBpr8YNFk/m6t7O5/ltGfKcFt2ePT92po/
wOOMyPc/ontjq7MoUfOC8SJqU1n6ZFdGHqd6aPzqcygUZa9vk4hI0Os8YVUuq5wNvx/V+5jErBhT
xPOGCNeY4WNLzO4xWyY97h1iCg6X/Lr9jJSN0aEa0vwEWYvV8HJbDb4+ZKosE+FtllXFOJ83KzXc
8kxGaI2dJFZvdWH9YVhpjO8wi/1BXHGOzi1iQl3rfgD9P7WlKpgIxDEmZNtrcQi8P3d/f7EirmpH
QYFAKwFuuVkr6Wicc5yNXuyFjw7cRELqITt6f74IertK/IMr/PQTOResBQvquPgFbTbBcScTuqaj
VF2mQd7UcT+tUJiQnhebPI8LoOzL4xZCwZE22lCeqJgaypImR2aNc5tKAqHPFaq4RgaBOpw2/dY2
55qCU+SYyhsFh9oPaaXkB9v6ylMMAL0X9UNz0+5fxFpwgIflc1Oot6BGiT0Lrmh9XVgttZ0TQ2S2
j4mpmWkF7z1T4iacr4VuwVOXHA0DQo+/lidS8JySZdHZp3BIZKwiv6pBCZhPXRtJRcgtfuXPsuK6
3aGPL2dX5jGaQD0mB2iZzBja8MCMz7gM+NmhuUXm6bU4ucUBpVff/zayQ/hSM0FiRPq/+kVCJMhB
LfyyTHOJ9naC31MQ0KRyb3YJla6bkB4KF+rmv+X690eIm51AaTV6t0NKD7hEP0nNXjMzOUvxU0I3
cSKJpZUDHubTIZQf2L7w7mm/ipX0234T8jfC7xWRHvCPhHlOrIB1zWN+GXWPexxEzeoBBAS0GZvJ
PiS4tvIb6YT7PTUxpd+Tc0a5rr37gj+QAkiueW4Iu2QVmbLHkkiQJ19vlXs7sXqjG1hsMdmiOQfC
4yhh/nt9L5n3SQn27k4GV4N/3NBbpjlExZFuroZaWZCeWkT6OwxVQbzkepX11DNp0FdPG0AhGdQD
IhHc7YwxqTjYcZFb+Z6MynyCac1kSdeqc1L5aFvba3HEDxDFygx9iGtsigJFUpjZTLI4qOjzizcS
6c+h4YjTf7Ij+D0agFR7XXsJjqZXEMEcgnMlJWJrEtnQ2fo8cgFEYjIoUSL+sRmKE2cjJmt/t88A
9r3BzxAl8E6SSibHM5snwneGwv2/1Tqpp1xMiGSCrjU1cfd88eQFUH+lz371dYxk1DjfrSJ+neoi
BC37IIQ8tvw09S/wDJb+OPoiFQ0/2wtjvjngXHBfyBVNH4MtiyMdHD07Z4fYz1thv/mKxeTqXnVr
mfWFcROnizDXTIVRzPzv4WeZrEkzQwXg3RWJk0SojcB354AC5QYJj4YrA+crp1/Ak1Sj7BntayCq
HXw6s/kQP15Ta+CE9Bha3uCGSI4MYHhwAr9ac1L+EvrdLda0FzY8hu0batIhMi0isrd+TV0r1G0C
HK7ojyLVlGYsd+lpc6y+sXl8KP/+BW9PnAVHshlgNjQ0frhyf3Q6rE4zXBEAER8EWtWtScnamUhl
I/OR3yvvq+PQorXJp36yEI1dw57tXUBEzE0Nh3+eMPtB+RJ01+dCbxCjv/r+JVrczqNpywlcIMRN
6RtWn0bLeqkAXqjPcPEikUUt/SvPbUHjBt1VzHRVs1cVpL4q4mOp+G45vJ2wNsdR5g7DdUIhoBOT
u5HMACdjccdzWcdziT0O40CeGkH6twBRXGsnFDHPK4P4ltbtZF4rywD4kR1ZuIO7kOvAiXVt2MlH
k3V02hdXG8gNQ8/1LUmkW14dtBav0VmKihY/pSxpeJCRU8FRxKEm//xb70BEDuzyFz14n36pCniw
LF73v2NZHOydjvzocSF+ZiU9fE30Yeo5wxpLTLdLAEHlFRbwUaewM02sGP9Wxt8aXa/gCV/K3Cg0
DfxlCRtoQRSpt/v/gn8eoVr1CzJOLEZ8/9ZSGMC0+QwqAbpz9BDwitDnUxs6371CcT+KsfyldVsn
gIBB8wL6Ku64Fdf245rIb3vneH8deXFAZ538efv49ZoJTieZXZxnx3yu6bIb91XbO3YaaICifJE2
suRTJBO46msRT9AfUhp1ZeKvdSevfEGLMw+4ocTUVknOsIsvJux33Jd+hwIcqK3yENKg3OJmcDN1
d7oTcLtKzEaBfS7C2CH54MslET2Rbk0aZ0ZCtTOb/05yJGKsxYXuhrLEU8ON/HqrnCYWKzT5bI1h
b0l6u1+AiKJof9fedWfXuhbIeCpPABnKXpm6EafsSNvJn6fEh3+8Mgc2zjDssaml1O8oTmh/o103
L0J3GpAjUOUVziA+Es0+lxvtBsp9Vz/NuuivK5j9JuTbexv6Ftcsoj/FH4OmxuxOAJXj0eTAwUye
o1KaAfRDy0tie1CJ98/ykYMFW3jVZ/F6yT7LT4FfGW6ewAs5953uwgNjCdt0y/zGmbPPydG2IT5J
M+IjBy9TTd2A3zSXgmHZkQzgecaTJx26GmtF0obg4FE82+vYpwpUVfygHAkm3rbtO1CFoh3O5W6J
ilYWB/6rEDSTsxLqvAz0aGyxY3O9fReIoqqfnHCmegUIbacDSrFBZEufO8A/cGmaH3plUeRZx4K8
MPQsSY1S2UYuBaPJsNHt/5EMAJ8Dv2PsY2/lHnaOtaLQxw3BMilQcDpk0zsVltx1Kk0pofSr/3wE
BSOlaAlBbuZ8ic5u6pUI+2FTxrokKaog1uA5Wq872QzP2DAH7Y9Sdmyb6xvowUeKZdfnCH3n4BcM
bdylVIlTe5H6APnLsi0bn+yf5D+xVHIyeOomBPbRtRdQNN7NZBki/HOch2HuV2cZ7GNiF7iJa1u4
dxWN2vRda3+yE66jSFFA4qGx0yt4pGY35hBxBOKc0VzODamyp4qIgN6IdF//xZ3LXTf7NGzQ39Rk
NOKXGuuz3qzQJE9nHYXMfKJ9ZeeLEPRSirdZGx/t+rIBZPsgZi3D2VEv09l0kaIH+PiYzgwN+i+A
lZNMXTST8sc2tV8UzGY0wzCr4uCq1q5TIUrzXT5avl8HR0dIzPnTsPkVvXyKljES28dLlgcNYqeL
MuC/RMQrxnn+HklThyDvGZoy+A/u4Mqt0I+QH66PCa0n7ljnziuf6V7auIM8mLcRMhHqN7+x+Kkk
oO72nEWQdLE98yQtsarRwQMx2ayFBeoUNzq3MEPof+CxhvSXVyUREdLNo5HD/pFvW9tUysV69Y8B
4oP7XIAs1N1fn7jflaq6MToLmEFciH9a1rVkrOopTWcFFdeV6mY2pDwhgvDtl94m8gqtjpZmlOix
3BwiKaR1ybjGey9WotpsOClWdPtvH6YVRLZCIabhFprW+quL6Yf9lJ6Ul1c8bpuwsnWOFxsTKYH/
zskoAxFk1cnLqYAaulKSOIHRqiHDDqeLAxxHtUFgNpevQeIZccq6Erug1xMpZmjESUF0vHgUFSUF
PuHTzkCPCuwLx6uppoOpWjRiOUaKi3q6VfFP1Xv/o3UZkGYO2ei6pmGzW/SRUYsKwFBefd8nxgwM
WvR2IYmntkxOVM58PyWdydEdtS98CzlNOO5PrkJl38lCYzdaObyQYB17UfJyKsI4gtYcs7p1SDV4
yf9vSopQbM5vQmHEqUYuQAYj2nur7xgQye88WHuQGUJDEhXM9PBmULyk4x/AM3aH+gieXC4y8bei
cTswNPEJyyQNEKmFmwzeA+UXcfe1DscQDiFf89yiW6HUlQHteLTwgvdE61jv/1/fZrABCd/dkEdp
aEPnv8vQvFsWnAcjCRn/h5VtAn5GU5OIvtwn2AjvjekWAkZyhUU9tpYi7qez+CXvRvShQ6zeAygi
3f2jCqgiO0H1FmA3dic2MGxL4Q5JJIqSPrqn6g7Fsz3LcLFlOWWyZf4OptMSicH5t6Vrq/ICJafO
Hd1YCM4ol9cmG5JBqlDfO3qqqoFV80MYnTmA9lTufNEPIDdh1VPfXe0CxxlicmzC2/duRFkgB1L2
Aj7+Ky+1ggRLVV83zDV1TpOPx+TkMReHzm94HRehl5Y5B0ccJTOgDklU47elgTIA7HRPkwVvOKU3
DZs0bo/cDQCzHITcSyI80wgh7eSRPcpxlcb69sScwlGSwj5pQTKrLkTMZsf7iqqNNXIxlYNfcSMD
YvyrEmFGP0D3KJJTOpiAAs5kWl6+65DKQkW674xPMR+Ib0Z/7r6kDdfnY9SEd7/wRRumwNgclMRw
crHrnQW6ZkxLPTZ44CXa5m/932JdyPtPC22hMzU7vDGUVHeneIL/ohko9XMEYhKx4x7/gmRkKlCn
Yea38FYpF6kRiE4BeKWvxUtzj+WWlqY497ZOQ1zgmYMBcF7HYIyCyzd+QYBi1DEoGaDdweynGtbB
MDyWMgI/4JuiHGqXFyFk2CsvtYKz56WqXhn2hfRUY0jRslWiqNxmMeWZOL3Ys6gecXQvhqBVxDCW
+wQ6V349BYaKfIk6PKqlFuMQu73RTaLyrfuV/XB3GmKFnNyVhXmXTLE6L4mx9bY39YmQVGOiVtdA
PCbvR+rFM2GIW/3JL1geI7A9bhdYgtbB5DLa89bDHFIGL3hQ16ACSSmt9MXCii7dLJuXUrK3EOru
fe2eexUFODmfXs96hhdCGmp2t/KF6nOhRWt3cbQH7CQa3ThLvJa0xOkn0msbPVJ/10/TpeSyR65H
wxE0LMBnu9e0Sn6JbUK5OEhr9ssSd3cHSQqUJn5sGVNuJGgLTcTX+IMbp85CDj9aavK30GsXDOAJ
DRY5rIrjr9ojE+4AUWs7nqMtdkzKDliq7WnAAJRvia0pyWpCa7UGhAc83ymhdAW+GA+WY8sCUlb8
8C8enk0Vfn1FUqSYdcpW6fWBfyC36rt8bdhI7sC3OWkFdIYJ80CH4Al4aPQRbY7nQKsG2avG3EpK
rBnz8gKz11JWZ3q9Co68DxjlZhGDSmm9t06EX4O8mPkym15RdkYnt0qM1b4KLSs4AgieHKC1Gul6
g5hvqda3aD7AuQ8er4XA1Cmwnp4huvsF9PKYRdAWWA2I/y9W3CFXiAMuYFvER8tXOlbJOdpcs4vK
vao9pTVtD2fhzm0wJG5VC5YhOmwClxIEftj4vkFkbv1gkW9I68rMcqhqEL/t6yyXlnKyUHsaAe7D
Lvz2fH16S3rcfulEv3WBmTb6n5rwkEcWFmEG3l+brLFa53QK1UwifgRhDUMRX1xD0W1MyZbodtot
mfEt+5YpZlBVyDJRyobuOgHO2OTPrPjOWymVX02QI5ohyNXGG9BhyR9BNH5Ns0lxCNF01NPZnjEs
5+71XjG/zYAzQMWzRXl6VZgfsm6BfOxEexFQw7NifoWYlAk8N6Plq/bBzKAYA+tNsSP6uXCTJzBJ
BMD7Z5EdiLQUri38bRdlMDEU/tsq8S/TXVe+SUABJNCy3k1rvPJ+n16EI6V61d1Zo9gdvwET6kG9
lQytM7HNaE4q1cD8Uod1HjK/2dnV1aypiBw4aM+5l19DQy6F7nx0+bjbI2oI2lwx3jOVpt1xPFjR
YeYdOYV3S+51RVhI1W1/TRnGw8GOuqHwkksK7TFelnrl7WpHPgMt2dQ3DBraa8S2/v4U+G9VO1Sa
ldYioRcS5nFGaGv7A4/jd/7ILiXEQ9bUeGqZkN0Bi8MfL1uxxmKNfTIS6uLKzsR3jzS2JTvx/QMK
G8w1sSS+gxZ4GKtNhRegvqLE47wSB9iq6wN+G51qudt2UFzTp264wDNzlpG9DicnUTalgSBmwjJT
8gxQceHDgfERtfuMHbBTHwd4gd0+kGm+ZA5Wj41iqBdNBNPeriI7EnKi1klYERIoQfO3qtBZ63EN
2gGvnXcdLtOMTglSy11aOzfGNTxYDHaKDjuW/CyEyEpSqbpf3VGwkqPhzqYTWf+B/wsaNHNKkCxr
1+v3Z+jYCwvzrUPoKOxXF7MGxdofpoGdXMr0N5uemV0SMQyJDFerdfngWk+kSTpVZzGZcOPNvVz/
Gzwkse87NlnFnRx0Mb92LIkVOmI5vMPeAfE1wV2HxXYrAgzX7zwzYtBCxyM49540GXl75aGVOt8W
FNCoAEIMFpuBZsxE9e/TrfGRGIUcWa+S0HIvx1bq9ULwjCW6RCwIP/hTPrWakmx37TD18F3yNFbR
8NbwQ1ZotM7BzPfEk3sHTba4dU/G/nrveNbUSySKFnXIijFl+WyqtOF6bTiX2p59ZF1pZecfuTwl
EjSdObHOs8b2dOe0YKBZybwIVAMilCExyR6JoT//NOPf5Jd/UBOZmuexxl8iEPBYjRE2PJzm03v1
zGZWqly81ADnUgQRJdMdlR+huCtE6PItI5DPx6+wQZV2AvoEBTnww4MiID9nh2f70Bzjd0uBKy0+
aEqtfKIycVEFMvzkJGr+2MjtXkIcVE/dSQDriFNnskykZF/zVILSxrZkz8RjtjNSnTYK7nQ/Duni
Hl+3UCsDhuONeb8fzUW2pTqoCpaURX1RH3NekA/uMStYmt67bQtSTz26HVI1aSldVmPv84ySE548
KeE3tYBL/8ta5SiDDORISEslSkvwRSo/BiMbkqs2y2eFOn5yjB9tfyEebz7bG6dZ0c3nC/slE1DW
8GwT77xVxIBdtNhs65zsZ2M6bY2WwyYwfbe+HV5Z8Nc5HcSkuKdPyIZl4UqwVVlIkdJ6u50ZlltX
izUBntUllvFIqvAZkojuG7OD/IK2ApdNPf2JoulAlwWOmByJYYg1xE+z8d83F+tEfH9Bt/tK04Pz
7Vedl4oqjhe4zvP5NmqQJRUyskyf4ZxRS7mQJZ72zlCD5t1Jyq9gUJwD8/aMoxaIfDE/CnwLRTG8
UdZ9hn6rzFpFNu9vwnvd7f9OKjArjY26gjSF0jCBf9Pm5MOe9yu0Hj/lWafOrE2i3K9kjzOalMa0
EAQKn9ZR+rqPIrZQLH6IL0te5mezXAFKIt7/LXnCIZAJ7YOetqSk9+2VLmqY0ZERVh3zzI+T+xiS
MI4ggHbbV/mKKPNOX+8qPpZbeLM3/LTVmlw1zNx5xpTPakE9+kNCg2Z7BNvicqDbOdAG4jNTT3yF
1jloWJAX03ZOOcvSejWKXgdZfVmf9XUC03BUtgrLJzc4b0Y2ZvboXTeuarVS264zpdz36jHuUiNY
qgDszO4Ack3qCHqz0I1NA5d0OIzSWXONf2SEocfYvJTE8a10WSWmSykhFFCPOcyke1oMg3ISLXs8
52vrjtx7e7v79r55M+yQK7wABroAW4wNifh2EoOoxusRrA0IGqQM6jSbeg91Ig1XPQVQTKEg8Zx/
7dNPSGwyb3VCmbYFcCieb72e8Xj9Q+R5dKB0jm1mehkdiDgwaNQO6fQvXX6mZ6uXrykayq/W2tLt
QxMKucsiM8JA49nWA854PMzcuMLRS7pgoTrJvFzwznLujfOAUSmju3Uu8wuCe8M2hkfSk9Ulf5pI
Zv4dWeOj+DkRLK5qNQiTu7UPp3R8YXO1qhwqHzHhsNNsqwxBzGnDJLJ6wHqoPbTGUi+rg1q4gfvV
bnaQ4oi329cu6JAA8f3jtSE/L6GODq0utsXyiimVxk6TSEXjF7KmWLCh9yJAzvgbYo2VAsIfCf+3
H8G6KoBwMF8agQ7T5jAqEMc1RkoxA61aG+FblfUdbUi/Xrhz3WHdlCexrE9Qw1oCxaw9PdxKEtu/
UivX77yh0hxYuUC+rbp5b5QmFnzLDmmGRqhHmfS9QlJQazqBdtLRkKawBd67b/Lgt8ww6Vyn8yES
+zLDqbDGJPIgYxQNpfIQWopwuM335WLwRO07F+z5lDTonX+sTjsDyB2KK7sK/usBH3/jhYeqE71H
XYq9Zdhi8/Jvhp9iOjHnjis3SyO9s40wip7FMfrVOO9CvYROddJJG1y/aGJqStieofoyNyJz/8Dw
C7/NLdMsq8DBpJbjZNUEoxF/szLrsqjLO1Wpv4rx2ImDgkJ+gzAo4twE48ugn0mIBmUxIiYhJrJ+
duAg3ag9WqcSuwUvJwauJ3skOJq07AVbFpeU622TovOPUJis7JnDR2MJOHWVYaJb0qdKtkocTJFs
1IcMKu1+pW5KRK2wRq7LVcjFlO2WvNtMSXnyi3lVJDkQTH+DjlJu2gqCtrJnO9vPwSRXBzqQf9oJ
y1xlS8S15tgRy5Lzo1AgoM3LGEsrnDrui7uZdYF6pnH+fTwmukH5UvjGHuKd5jtwUW4aI1p8gPbE
lLwqj2UX7jpgwp/Z9PtITdRNbFidso/DAI+udhsPyceq1jPScnYOY828Vvk2ZiQDABV8DzDiewZ4
BW7W9BtDAklUs4hs/FeIllGzExnqinPf32OJXQJrapaZo7wxapTK8j+Yt0QnZKnwHETemoTTMzzv
io237QaO6YOTx0PM1+I2snrBND6wbJrOZ/7AYxORuEJJRR07K3iFbO3kQr+EQEr/tVsd3vYanPRK
tmOOfjq9sQOvsgxKe8giaDSWyR+cIFFSaNw3qutyetfZBNPCmRPBqS9CgWTrqS5fw5BF22ovL0vk
aVfeQ6XXro6hq7Tnoz3GlYtSp6TxOke4EloIqbDci/xsVGdSb1Ht2sE/QoThnE6n8riau5VjbMsp
JEOoJYDbhJtOrnqKHKEMdobDAx8hoUhBXOVHmHSOWxWRd1uqxztRbhGiskms9f3PXXHJAIOIk+nU
jOh6RwlWHdursq7zupdk6Iuk7TySliBYfMYX7hYpTGWXCmhX7AL5ce78iSKVkVFxPSxoHqn6CUWn
qIcXOehuuuKEGCQCziYxrWrNuUMvNv7WV0LDYvQyT9TmxGcGJwycTSQ0H5ov1Xzr4fXw1uqmNDxL
H2QsxHKz1c0mlzr5P2+dXUvIZK9eiy65pqDowDSDa6ewr2EagS5duxHsoGlPrI9sJLy/ZUKUhcf2
2VpLm0x3cP7Wx3WxxAEs+P6licCQX5vgxoR6D22hmL8HvQir3sgrW+e8RwR5UYvxVB/N7xN+uftr
JCTWM4LfWRSPcfd8Xa4sfuPSiMQpam5tGvqtwl2+4A3D2Peor5mGv8I4MNcQxFVAr094SK9R1Et/
4bzb9bQktWq9jYUU3FaHhwvJOGMqdDgDobqVusKCH1Qr8cfTQMIOvdGPdqDofcEEwm8l7cC3nSvp
vjPQVM/dkop7VZhk59ytzdRBMOr8vs7p4K+LZ2SYOIiafQzo+W2hVrm6W5p9+tlpuFZ91KfEsXCB
0zylP6wAQ1VVrRMJ4K26CzTrEm2M97DZAvh3b0+aVDVb+kBBmDIAWn6I2Rkg2ijpZNn/edKoHkTt
ELyRcvFldxAESJBjAHEkpLAZj2jvuBhdMoXQKC8tT0z3MuOXThehZ16YUZVsA7YIw/a+2UZrYCTo
kFBjwrKeznddS+WatBHtIbkldAeVhhJbhKHYj5ymbcG2/lSkzvfmwmMI2r1Lr7NCPjL4OKE/Wkby
hZR48Agf9s43HNsXCn1AXD1aHRT+CHAWfVTRQXRng3fwv48W0rCTgMBrVZkkAm6Z7T69HgvVoYJ2
asJc1QBm4oQ0zWOP7jb4eZ9uO4nvS0GcgAVmzYwxtuXOX07QQ4ucG4WBSQJA/Qw9PVeDgWRccUOs
ZNGxwmFmDKfrOVRm1JKKBinHLxL79LMLTKIbQawkNMOzYAjf8M4TqGq6z5jKhC/1Tk6T2HeXTdad
nj2oa0RZ0BNwmAm2mGhOU5eqzuKYJAPQrW8YwE80eaniiDXyC58mOgW06iH9VnTlP+Gqop/8DLo5
rVtoOlM2wtu10EPTtjoTV4116sD88W5xu/c8KOtuj0mHpZJP12K2R6+0YVEBP4Subhgono13+ENm
gszYxFAEpjxjMwqcq7VnRL8PZsn5btuEV3g8ltMA5NDANTv8anCc3rLZhD2IVHOLm0cW73jMdctT
O0AzbPr/6vfDcl3iqWqevHmmyCR7CI1jEg0bgAH1RejZ9OtTOuqgFge+dwkG/RGF/GlawKEWHvMM
/UNv3fIgRs7NPdYqsZSbd0FIqQLwtOY3bJwDc4T9Hs9L1te6QBmkhTANK5E8zcriRM5ERMhuc2eJ
++x1QHy4PRHiZDMG9750JwcmoJyr+JYvszqr1TWFG8mS6ij6PMdzWLTw/nnXJrOgaUHRhyPz++tQ
4BqYfiBEsySCZfOiYpRXMQqPccOLR7nIYyHCrhGj/6m/2Cizn67LJs8wd02q8HJ4As/jx77+aU7Q
xQoseJNpM/y/+LIQOBBCgqqlkZP0mF7s4oCdLgstVrDedoaUamjUIkcJ+OO5rEQ3HrymWaTx48a1
J4ffoulLP1C2qbhyvdDg8ToeIL2dgiPz/c3uxLyCJg4ZEs+igZV4ZDjoYaIppGIq9dDvtDsj6Y88
zA7X4Sqj2aHYPQSITkvQ4bvg4axaOXVkG43KKAJE/Wik6V9MXVbu3RpFf6ZQdirb29Xrgch2sF7b
0nZ1noopGkAL8Kruwb0Bt+zJ+38jVRyuRVg7t3zFnPvs6OO2SQGBGFq93Vlnt5Utq282ERXbCzC+
M/t3PynJ60yexae8s4tCwiXxLLEBLcgdySPPcegv9KRSAbt30ad4TAwdc/v3wXlxePuM9vxmsCT+
LAPffPV1w6C07PCFk0LKOM1nDskCU8BdubAvhh3hEsbqcEswefvFwQ71JnNwIUyTtBJ0hkuPoFDh
lOwIpGDGCGv33qg9kifFRwNogs0YiqCR0c53tFPppty2vcqWNJi6AI7SFdaEO8ShVTO1EsLmnPEm
/9ktcKnf2SnvdDAj3+9vvxhu3ztqh++h/ZqJEAYGJoBsOqbX+8EV1j3jViXjcP3E4BydUU0y8rHJ
dft79gEZGoEq93kacBu9aSVwIgetImhUMkyTpXewnOaIymG1ah1HYJRMMPHr4wTPS5eNg2HunLJg
h9FZBvMJB823GiXNfYKZlKc7SNJZebm5f2pUSKPU5aLVZaAQyTsJu7Ypm188z27sbDlcC6yM6VdZ
iuyPRJS2MiTqwk1BMeUAiu8myAD4SIk37hY8YHOhk65k9c4Ei/15gcy1FufddHW3HtH2+vaP/4ZO
lR8S1ZySdV6BUSlsDfqoeGZ9VojWr4jjs5QPYNfZcfAF2cvYROzqJUHaiHfC8llnkSejtQuU+vqe
UB4SNKM4CMKyr3maBB2V87Yq4neb9w/ie+VQZiWncLcYJg4DXLelnQsX5Gv474rMmq5LLPxMmnwg
JmPenCSN54Aaw5Gmn9d7P/rt0OucldDPaJh2dkcHTz1yoE/M9abGYsiWyYpJTBu1FbWWq+yFDipC
hjdiyV3VFZ+wpUiRAG4W3G/38ZL7bY8Nlt8erR3TvULD30YUlJOyZnrKmVsR6T3pBrEEGuJLj9x3
K0aa9qZlVjhPOA0Cpgju9uJfcML7+tHTc59Q12YRyGjseKj653C3SAVAZHefBqw/tgUumFcsHhrC
QY2LZ7uByyIiuEpbfNWSZfoZcNRidjnkLg40TmzPhehLF1UJyRhvyG0iziuatRxI3rENjW8sCbt4
KgV3cHpVRGgRkczcSeH/IlTtXAbD45lDa847WUpKMVGPAi15eAbZQWBZX2dUTshluEo9eyvojlkR
DTMDEWkBOnqNc2Lpo9VAWFuVdHljDBraHhizDFPl087qYrlRoiytN1d1t43J0Cp347utLfOEB6Ir
Q24kGVwnjpYHL5dRS5/osOT6x+/Xch1cF1wlvgFjKU5ltW/iEeZjNKKySEXcp8NAoUYFVxHjAnUd
F5WrmZJYo43H0/OM7YqGUw9I0DVnn8h8AZPLzihLAdLLyRN+79rqu/Nk2eUzKpafBUVNeMbTKKBn
xGLeCI3lRLyYNBv1JwLl03j/ENFl3SFZU/L36F3q74qijtJJF/lep3HbjLDhdCRTIVjYLiKqGhsS
fSrenanqe3szeKGtOoCs2rSvOqMlyn1QRHfML9syvn2ytBSzTxbuCpbA8cmMEvg6lfy9mrOEmmM+
Jm8iGfY0P9r7XF7VOb386IQmiYVeTurotCC/UWo+A1LN8I3AFZQu4tVUt8YmXGO/tZrH0dfE1fwq
/7YdfR6cfGyV3I7kLmRWrz6cfC68F2pqEnbesh/6XyeY+846xi+Jt4rwG/3M8rwInLvt6jtH5uVH
HWsYuDrSGU7BuF6JYp5YSJAwFPj+F9wyBm/4UTBLPY41KRFrp06Xam0mOEHPr+xLgFlB5xEqi1Tc
dwdNGVd0kceMy2ZYlF34QDr1TKkwXf0Ier+JaJDJErXhLxoExooXkkWC7wMtBAi4rFdx05tRsJSO
C5MD76EzxOCqJUqcUshiQ50zK7Lr1LASSLrIOm1/o4lB5XCmGwzSwXfKMZmUMZ2XVikmF1rfRPyX
fp1grSj9P6vfstm+UU4yB014/M1jBHt/CpHepu7Tvfeg1MJ9o2eblhyWHdweOM2wwo871PevnHAL
wkEKXschE8caqHcPZuOxMaE6e4oDITUQDCaSAcfZeEVX3c8G23Oat+nw5Gdq5ogfq7GSjQ11+gXC
cH3r2HAYnXIpnEYUUj5UtRsXoTdX6bWefx0lZtjAgSJP3vu6NhE4gurvTmrh7Y8mcfBow3M6Eidu
8IsCZfkzXNVe0Rqhqua5JZSqMtH5GXGh3JhH4590aejh/G2zbQ0Tl4SPbvw+uakyZB2jkAaZnK4M
UcPtiMJUdT3lISyJ1d9t5Kfe/1WHE4b1u/iuC1WGhKSuKBzTddkVw9or6zKBodlOHNjuIzwANI1r
Sc214zbkIUofmFazXYJ1NnUH5Z8nDcV3PmGxZxSBAvfLgh7qOKW4T9g6XKxNs3SaW9+z3OOlb7AI
E7+5FedgYa7gmZdJ+N8Q5HXllTU+aITweuPJA2DnbCJo8/HWC7xRrVuRkO/cotEwGDJfNd+LawJB
kbUv/lkHMZ7OtQ4ZoewxumO39XdYevpGEHHFj9YjWC0V7nbF0ONwuDAzwZyzoMaOMZ6qCKpWxoWZ
TN+4PZXw1j9G34w5Lgg9zYJ/r41w1FNixXNxLZ4pFQB5pizx7apejWyEUgXckLcy6v81YLb5Ar+G
QCwHltaPz9QXxvfNu/ddtBGyA/rnqCimDIEPYDc2cg2LjRVtrw4gAU7mAbCHN4i0Xz/RlUkCJCg4
TU39L/tPMLIxHRGCyVlBPu2pPjsoHSZopdRT+Gho2aDLehZZpCDhApWzp/vq9D1wvDqQwb7rOSLm
SrZbq+DP7GkX3bcRppQw+3fvNm/9xp31GoGyPHn8XjDeUHL+gC22zxvbgCLrbVAXpUq5x2Qpew1u
QKsN+ih57ioud8gBnf3Xy5rU7NOBtq3GsfUfmKfUYmW1Jb7wT4lat7NTEFjfG3eyUGhjKPRuhlAQ
c97CKfo44jh2AdSbAmb10E+PQ8ujUr+Dk4ca3qkO6dUXocA+lDMzPYSdhmYIbQR2caVZjUvO/wlV
hmMTJYlgTu7vI0c3cqwG1g0CJmT8+/QXLLZ80gQkl6gWS/OAWT3d+FQaMvR+5SC0dgIJHEvXd/bO
4vFUgxmtbo+CVIfAV+OgX8hAMm1RomHGZCiDuQsCZpid/5IuQ+dImsCAu4Z2/jpqKETo0d0LiVxA
elyMqcO39sy3h/AphnI+3R5xrQCqPn6j2VLfUo5mtVVt1tNi0usi+VGOXuo2bFSgLyxtf2k2MOhB
cjnSC4+1JcxhomhK2K22cZZnng4FdnKTIa7Jw5O1Uxy8elaBFirTERci+CAYffSs9I8/t2Lrs5Qe
W5vWH+o3b4QvZFNcF6w9AtdY2zTk7lE9KqT111D03+/SUEuIsyIUyovA2HfYqDFe45wrm6c+3ivk
jtPrJ7thN7YUq3BhyscT9hzG2jg8dRdDiSsRBo3RAylxcoektaHe1r1Af+p8sS0sMZYadtkMZSA9
5qYkpjcAG+tf+y7WoDZCBvemfdunOCuDpWYImboK3onDfq21/jXuezKUh9dCuYNTwev10ocxBKyy
ry+K6qtLctSGzt85P+ooQU3c2/RPIPhAVy6voNumh4sM14BdIvpTdqLeViPRQPaK8DFLkUg3qpXy
7jr2Qpde5uAha0AlgJSlJFtCFa/7oGWNRwbkYY7Ao+VTG3l2cE/WVpOx4ULKZsZUnpz7jYcPkknA
9GEJxamdzdJ7ZbE1H2PfcUEBxVRS8zIZdesPf8imY1vXu+s5Y1jAhssZQDEnOfKYI5SF2V4FwgIF
j3yavjgneA+pBbIg1PiqSIRncdl9O3gpCsMclIpJi2KfObdV44HuAD1fl3E5QOjeI3LGgL9KPAIN
ZFiQiWljhWpqwsZsVB5UCM1DGWcLpnYdFjK6ohLCg/oHBRinR64jv9KGy4iMlJVon5mMODE/4o6e
EE6/p93yPKLiGr6tAgNnI/pQD56102CtyxSvgpCzG17mB/vq7/WrW0EWdIbXed921um9z7lcVhYR
FOss8+MK1pRF6DsrRaKBtnY1ClZo8hsnNQOW20AWEakR2LLyP7cWrgt7StyLkpiK+0dSicfLyIVk
sQ2/b7DQD+7JIaOwElsF0nht1wmvIiIHkuAesZVoZbeivHhps83UmUErV2e/I/UNc1VMivpzMJpS
3Z5MyhLU/xMC+wDgNy4bZWNF7vrGj5X/Q8txdlwDkhI/BfnRyZ2AlkJCcgJaEAdaas3o8jjuzTRV
09OUCXcggNG8AGws3L4MthhqxpJjq2pOh4GAG5fpfI4VKD7DjMYkGS7ozlsJeLNYOhqpTzQI3zlM
8Z6BqTUGcxYDRHUJEHmRzaNdJT9Ze2nnfphEU2EwyeQWpugzGUX3K5CdMFYONwqtu+WORrbN+jTq
GDDrnkNAmX1QXnAr7lLlMIhwuFyMd7QDpeU7W5e3NTp+b9gswg1rkHBT6dbFVrqCDT8jBZ7YskeW
hPr/OLJ47bgvupyYR+2PYcgv3TpQh4hUoWUGUyjwmGO2XgRCxy7ztC56KP2yJzegmeEBDNrlaTtw
YYk61tHDP9avPle+1+SxknAJMWBoS/w7p2hoBT628HnD/laiffRw+vIi1YzIw8jweVe+TqU18J4w
OEvcJqQGAzyQegwS/bTwsKfOF8MhK5isER4Dq0AA3vA/B5SucrBFPLEBcS1gGngO/Gi0fGZyGJiL
FPwAJh+sCy2G7HnNEtEYTQGcl0if8FBIgf3KNRDL8XniKTuwWcEG6s+0z589AzcAfHGKT+gpDq/5
z3ljo+bUH1tT7MBZLNpnDSbiP8RZW1ECTIX75sTjSTC/Id2UMFB9Yefaw/h1jyVavDGQ5tFb5D8D
Hb/NhNefxKXYoO8WB41c041/ufmec5k82Er0UQb+iXHynJ1hHzwoFnX9Ko2VxH2Jd5AniFnSxZ90
ZPqOzW+Xdf3cbjHw8Atvtof7IxA9/HyQiZj4DuqbEGcvqBENJ83w23thyZn7oV1l0aefyKM0b/jE
u99zjOengTzlwfdoKcwz3w9dZjg/LsJrJvMDttHFY5mf0EDW2Y910MoRtKt2EpyRdvrprQuudxed
RQRGSM22/W3PMLhkYEauxTvk4SN2igklOa0E/xHaV8dQwe7T2nY1HmRJBon/6TeUiDp9ckvE78bp
OEci2w4dBcEDrSgg07SkS9PyYcsbQ3F9Q/b71NcE+A6Pkm70FqQKOFwK58HMd4lOhXzoKaJUCNLe
IOPIt4TdUv28A2MRExffcxBv2H0BdEffX1IcT1t39OvSgAPnIWkMgaKkufKwC8rk8RFKhkMLqyK5
a5Kl6hts+ZMbV5bi2ocd+nmsfLGVbDBLBEESaYSk0GjhD8U5fNAw0LYkpbTIWHWZIKiu3xLk2WDQ
0F/ur9Jyi64LnDE/sz7GdSyIMQcZV469SeJAOgIRNpfztPz1/YPo+6ewUYjdKN1ysAHKShka6WEp
c0mMuuLokdl9ZkTeSuK52tXYQqQlyBFxr5xCs8+iqABofe4KJHbR5h3JvOg8/WAWO8Bi5tB3FH7w
Fu0AWKsng/HIbxVOUvA71+0kuiaqisUnsqKdjYu2BlR6OKgYtqFZatV5EGujuZOFTJdU86qIJ4fM
H0p3Z/5Y0GcxcF6TeS2n5U7lE42k/z6YReeCtDmRgqMbPtl0nFlfHQY1reeds9c8uZxMhLy7ZMew
joxaAYXWo5J5ufHKju661at0+dJwfvVa9DNXZ4RqBaRqned1b+1cVwubpk+U96UiAUFOIQUGQBUS
+AFIVBaJGcotzmQANdpeyDFi82K6nA/O3ggzVVRSF1hBGEjMwEl41xLYIaPpaW6RgkY6kTw+9kv/
G7KV8feUcYS+AxtdAWd89x1Lh2epKhBVa2cZAZTQtsZyQ0zH4t9csyv3AGUjb+Qkkvf4gbMZD0M0
lnxucOtpQvRdW3zR43NUkYKMsPFFQ5AGj9ry25yAuTp8SVsaKRoRLYRfA5gEcun60aodX3wZg3GT
XZ4Q9JTHcZ5qoRutKSkB77Q9YN++WiChxuAWiRbT8uVB8Kb8raeDFJILJBBK2FyyzEyW8ke2FnLT
MKG8Ssp9hNxcFj+H1eszR93wpMtnxzRgsAxxfCrYU8xabcL5TTi5mOAEFR21h0H8bLNQwpl2pA+Y
zH2znoRTX4ln2hguH7xz6VKzd+KwGYkruGkMLyIX0YnuZhMFx54q0a3sKU9zeRHD3UEfSXKcsSCB
TWUJRocDdqhPaTld0O0XFOiwqzMdbK5mQco6DOH1zsLE/0c716SAQzpKiSNxhuCzIIdkJ1UppALK
lVMNrCK/a8mhIK/hlqRUEqe4nsEstMxLjPhCQ5KFXEmH233PTcGJQwG5/PwPZ8PxrKldMpBYa8l4
oFIvA1mHeny1UmJBZOaYHR2Dbvka/FcQ99wcm7kSD9hC909vLRyy05lDyIeAjaY9zaEzB5eITBdw
WlXHHlTfHBCzQd2AwiBMe9IMzwcTaXZDAyujHXV2PSHsNuTYhEAHldHZa5u6XMnfB7/M7F7bKaec
brftDrbgtQ+xxk7EyLH/iikP4EsT+sGenYvdN9QgTJ9hMxsmBcSe8NaIyHuTZPm8mCQ6GqvVSAUh
4FYSOH5aO/MZnQqN6LywPkLHsZ8sXc8dpWDfkH3HFT7j+fI6XN0Cg0lGTJ3wxNc/YtgRx9oJ6PJ8
PLu6TB2IRRNoPMlXK9mTkD6dQnnM/Vkqpxw5qA8VV2lLRrtgEz68UQMTq9nvjfXaOXOLfc2hXJDU
+5OFrKvqlPsS5MybOwaoZ9S8Dc3FJQUy8z/ogCT0YohFfeHBR+IdhoBR1P58mvem8k8RSpZMvCG4
PfGN0PSOYh7PEZW6sWkdDLByOsOBqF7yHZkY9rnuqo44JNnKsAKrVD4Dp+68MiB8ROoIZmK9NoF/
6KaBGBL3bGVtlxoYVg8gY3JsDUwPQwPKWoYSooyi0b0Ok4s/17Tjb1UQv12QpZRdV142gkZv6Oe4
0EKtJK+IbxCCAfY6BBi/ql7aBq6GmFEBzqcf7Z9Y3lo1R1EXbE9d5Y2IAiEJnXRE/T3iB44ANI90
dgxJwlyaMWYoa1DB3J+2vmQQYZ1SjfTYmHq/k5WAYrP6TMe7oq/3BoEY+vyxQW9sBr8fjO9NzA7F
f2QRanF3eRMAoD6miKx5D/k/SZEjHLZZdgtkgEQ6AVTm3jGCtMA/ISqJuTpeHiUFzPLNaPLdcjG9
5hBdQ52WNRHlFmSDg5KdMCiwvac5yTQp1uAA0R0v+ELelug/p+lUXIYY+/DpnRxk5olV5mBGRGOH
aBNjjuOiYdT/Ysf/1dGSRjDCmKPShllMNKLaoGZILDaKrN3nG40FTB6uLLY0TOKNltA9n1BzYP5U
PGvMBoVugzqNOc8tlhAvRGm1ETgZGv6KZO5HG5SA+SDa23wYEkhc4uHMAbZ6q8k2Wic/nrxHRc3P
YBiFpBJbt6TCUJ7hOkY7p3rqT/ka0aYcac2okmC14d6ivyqD079vw4Ta7uHv4Fq0UYUtTW+yI1f4
r8H7qBkTtKapXMUH+2Dc5SszSr2gKX/uYgTD9C7eCuQLZ/RvGcn4X8U3MpNp2r+kfQbA2Jlwttin
AX6EIUnwWix2MgBh6Qk5lCfcCMNlzDITa1bggqb5XPrK8hIWwGK6bcZIaNZfLn0gV1AfpS8f6DPd
6/xRNxeLx7ShhL7on6wz9ILJP5l2w/Q3IFiYCiXEql2SftjU3zTUDlm07/bkUcGNq1gC+aQd3SBW
M9plEpT1zzCPMlqrrbunTJhg134Vr4Asu8hKA7+5bgyFuyfViyzOl5sXZ78mbdAoO+tB593i2jJS
iibXwZk2DIFSMiF8U9BJv9y/Q9I+VHS0P5vqII4Lzd5HBn75bRB8OSLLSrtWijy+RjB/SAOoXHN6
ga+l2jc7t4cE0LKMvtPNIvBEsm5CQatt12ivBTTVBH9aIEcOAVeAaAtObGwYKoMU3UMBZQm5ie0O
Zk+TtuCQcST8BFDWOCvqbTlBJ6pT4K9ok4I/v7LuaiJ2iGqTguzMzCV1Y29wEnRNBl7Yr4u3o9cr
niqt2C9blJ8cpUUKWEcBzLyfxHbLkNCJQSoT+sT+gsmiI4JYOOSqqD9b/p3AzzlZP+KX5fqA7aCT
952Uipac8DaJc9688/9p6GPugQFyJJ4mHti83fshOIPWbGDmit4znVdWxXZhhe3WWNQchq+cD5Uy
YAKtw6Ym5TipRdwsuzitr1Ol2mtOC66x2erZ2CAHxWGkyXn0SeMmKbUrVWfd6xCiCV3lRc7Gav5D
Y7Aym+5Y0p75OYg9laH9jSaop4zocmEJ4Z5HTUkvQc6GcXxxIgFY9p0SGYS/KGoEHhbhnuCsE6pL
Z0nBfrlMQ79VvNGAkywu+7O13bn1Hft55x8KlILTAP5LD0b7puhYqZXtPR777jcNEOQ+SsXc/ghb
NMD2fRRbGpMdzQyUBs/V9kdJe1wXmZ/vssEp9inOcU3rDqYNFphWjKXuyHoQVG+kezh98p+WXQg8
PirEbnujBPa3UtIkA9BTYEWVzk2NTbBr/zB6VoJ/iocniz31Preo/OvOexX4yCQbQon7TgeqEs7m
r90enQW0Dp3i86umlPxKR18fJLyccaEKvmfzq/J2Ud1c+lQCzFVO1fjU480wEVNjGB/MDllZWojW
zo2+j1MpDlJGLJNGyk/47pasEtm9/kqtTi7PkCuaDT7Zt+SZMKQM8gvBCEmVzVqGcGr38EHshDrq
eA5kDiRkI51c78wZEQRem9GDV0DrVqyh/uhn8B87FZMU/2Pyvg1W83bz+tMdbbDK/8eQXY3svIpZ
u/BwGpqHezM5nBNc8NzXO+xTeHV33DHOK6BqQU4I8Z8KX0C0NjIDyHiTmOroQQ/vu0oHlXO4tPH2
tcxo0UkZaHIGLN+SsMoibk4BG1G+xHmWlDkMi5mlY51Zy911QIPcu/uSaR//SxgUoAyE/FMS4b0m
kAymZalgPvUAYW7M88un6s4+TJsx0/vF0ix58UMJqbzu50B1Y3ZaqFFul2/fXPA25bGRqNmC7AwP
mTtxfOWJp1O1aNkqbRUFZTL+D+dsd6Kd2ZeW+HcWwrS9i/Ngz1EKkluSMS07aJQtqD9jGn7sXeVG
5tP9ZHQhNdvmN356xDgm9EyprNleSuLIM7jIBv/GytHtNXgqpRWalKnas1ozF+tJPTnW+G8cq1yV
gQjyZYvOLCO9whpzf4yO8aLEBZOdqzj/qX68z4fG6B22QGXP9V4WIsVD+xNRNk79U/6ny6BxQR/I
vy4ahSSdT3SmJVNbuXr0D6UK9Q1X4jJ7s/8XeMAlmhbhs8ScMvavhAwi+0/qcG67LnlZyaAfZakC
91ao0GJW+OvmI2a2TMQG+ek2uE0jtwLl/chUFG2IAOoF6o1M64XmwQsXival0TumzTvLGFj5v2+P
EsklASbzYcyYP07SixetF8ilNTXUmxBwBsAN1mVl3CF7Pyy/yG71UVMWN7SnYJu3Iaj+iASg7DGL
mqtDlSI3XpnzuY4lloJfcQNP85NnMGDUdgi0/YQl72jKj+gvHuzahriaRoDBsfG9fWSBqR0pDJfP
Rc1XGdDko85HYmrFUVKrDptwuwTuXXJDMpQeqeK5vkSbg3xB9D/fSZlNMfTx9SCUN/36Y/EsXAmu
dOGHT+Oh1sSRecLVL+CRsfyQcJzaY2tTGx011X4r+TtBg6SWEwkcdC/TvrgVTXbOqLN6O/nxuVDu
FwoYDBs0R4e1/ZFc4MIWuvKvEDkxzskDvT/KYCX39I8pmkLBE1eIp4Fip8+4vaMvrfzeJksz2w+Z
k6+vL/ypa5Ey7E4=
`protect end_protected

