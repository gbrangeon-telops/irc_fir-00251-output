

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gjKSpUobpdaEiN+EJKINegy9RfobWzPNNvSuynmxBaCaiXpZzE42DUdhJsa9nuNl5zrnRUR14CdT
xujtPqnMVQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VxmOSrOiNTkpjQCdEraeE2yE2mnMFQ7pRVDUX9VslB9rFCGD7dNvbneDVpuQoePUk+nSB0IAqnFe
/NakjC9Wt9azzGAltfbGlSpsCZYTQJMARswgnWL4Fmc2+3tN+okF6OFM1YLClj1yRXdxl+CDsxQ1
FBT8tPlhn++ZNTP2k9k=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aXqd6ynCn5cZfxJpxEun0CmjLX7cGy8EmIQDak6IkAJ5uWqWXRabnrZlR7iXAJjslJ8VJzSbOvYm
rNknXsQKfebDaT1iefkZ0I0Z762iOiWvIR0eap12f4JcJvz9RAzeBAaW4ZyAkczx3IYLwFNzh/0g
2pHrl6Pls+OFuVt68hp3jwzH7c003L035HPpddZ6HFBcZ3MJeQ/LoNxx+FWSqyEG8xTwd196QL6n
uNyNqC2ytbe6mU9D/s5w5KpomKyiSs16Q1gq8Rj3swuI/cDlyu2A84YTnDD1OVt7+ooOZIymcF7C
BaBzVPlYihS6ibZatAmcUNJ2pZYltRbTtDOOXw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S9smd62+t/cc6T+Az0vn0kXxFJK9ox1swzdVaJK3ag284vMfjrlnVswyLQNkD6M2BaUNuZuzevou
xaHfzJcTFt8YvMUaEn6TameCIs5/mTCxVsde0MlJlF2crCf3fZHzWj5ooeKnlSFJXuUK/R6CGS8a
2vO0yBw4ZENNd3h5OqE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cOFUj+LOfMo1PTF/10pikQPB0v1eZ+hPEU+cjnPIX80Jf3IXfuV5X+QqrEh3UZH/0+YwNN5uc8yz
3GcUBcrBnY3TVkMqnhGUk3sy243Fxp5BXFf4yGZm4BbuFXxSAKu5Q+k+UOvWrFZfWdNI4lYLdSEu
b+Pg0ebBc04YBsQL8j7TFN2y60Hw4npf4Ha1Oh0Q36x952OAGQt/kpvEYJz+iBAv7Wj4b3IJAFhe
Hz1SVdnrXpsS0DFFqDApZsueRszhz8yuOSjC5Se+b7SzsP1onkP7OL41tcS1dxgV6XpqQDe6m87o
cIvrt9MVp/aWXYppakvqJEuPRZUIN54B2pTOpA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6256)
`protect data_block
TkVMXuiwS5+/V5KSCIWINAZfej6TlblzHCR5hyoxPdtNmz6oTqQ0V8/parg0pENugq1wT0RTbHfV
fRn8ENj+6Pio2MxcxtFOpIjwzFc7SUx40EtJuRVYxvRO7Ru22+pFhjSXEsLPRAbDBv47K+JntoN5
ZZM4f2ic0X0FIE9QM6L7bKbS4Ackp22fEVIFIbw8TX+PTjZBeH1U0azWolQ8RN3iztZ5xeMZXait
mKcEbUrjI32KSSSd+RPOfefrT0YF15TKDJ5Hr0/b6sCezt7u9EyIxR2R8utcT9n2hLsczS3Zdym2
rQCegmKJMy6Lfg+a1I3QtmBe7kPGg10dMNVt/n9idDS/MFluEgB+/iTwkMW+PYSD3YDBc5LXFsMC
O43q38/xXbS0PNmzySwKy6zGbvbBwwyuj2PXnx+Hoblrp4YCJBVRTzNCR9pg09uy/CyqFP1WWrSE
s3l93o1LCxnlzm6iFAe2DduzZK+YBnKEUuicTigSbbo3tRhQ88FUfcSFUqsv1wWEURRjhX8WJnEA
JajPMhkt2lB4CM2rVUh0PtWkn71Yrxg86/MFsliO7wIW5ceuCJjpjiw/0cl+tEpJsp+Laxts8KhY
4dOOxYIB4MZ+nTfqqmtd3EQRqx+Z/M80RJuadOSQuE8VHFDdVAyLjg9iVSbkwcv0PAdFNRS6TY+U
rFhBzku2qKH/JUWTUSnB0/bn6mUqrWHoRSGVKVDfILO6KlSou/EnVX0ZFmPfGCoqoiYRySo1Admn
yScoN7CMhEOAjMtabynXa2wd3qif0kJuIR7HCZGpAusC6j2hUzrUYZlbs+h49VXlllfQZP68Zmv8
XiKTeFgBsCRUroWPJgAy73dBwoma93hS+yHhL5Ow7pPopfP76uFK5nijUzYV3LQTEBSY46QAemLz
KqRFsIsHWTP7xXqGDYbxZ5PzmtYlZhz19HxUsUBu5DEXUdXUvkkBIx6ZS6vpUSlvUyj7gbGOABho
EtHDLBHdxEEELvBLVJqKwYL4GTd2n1vPRAVcKBJUxK1E0VzTrFxzuJJGz3XQu5WtaMziY9lp99HU
uF6GjzGq4DIkMAVY3nzVRMrpST39nsmdmbViyz+8MU9hHibpmZnPHC+AYSSwRr6Oo1b+liQnzV94
C8iOTrf1390HuMfJe2WRgeVMcUgCvxnadUYjKlZVUT3JsNV2kjnUh4ON36nhUMt+5R75Cj+A5owk
j3+jgy9WVN3nqUCyLvKGyzl5UvJV6R9mVhgK80wOGF2y01RTNeMlPlfgISipTWWLmart28hQR4B7
BoNRYiOh+Q/Et+ywfXQWrBNwuJOfdXxLrT7Exg/uLpVN4NPlK39N6g82n21Wnu2BOJ/tdXT/OOnc
p3SDjYG4LBCjAkfHpoTDoynNW8K+UEuENdSmbn26h+Gygux78hUpExKs+qtIAwKfBN5/3jkkYoWw
k46dxyj0X4YJ7EAvy9uOIWVajyASHCxqGwP1u74Et1Laxf6ZWBpxCCvWFoDUxOtM3nQrOZ11fFRR
abDlleU9arCagbsHLZxHyrJ+3aWa6Twh2Z321d+FaZ0ZRJkh/hH07PjoD6YifnTcoZ8BB4bd9/ga
U6fgdAFdhOA8Zj+dbmDONxIlvmFlCBe/YQX0oSdAfngPJ5cAvjuRmgurpI3vGV6yg3JCu5eIAVdu
+5mIQBUuryrGWnouaEgQ0g91NLvTCZVBYe8Yc/jqY9k/1y5RLbEqQ+/CBKx61fQVCDvaZum/Prah
aXAvnFn7xW5o4QKLSGvkR1QspwOTjIMFVgMNlKkgMhJj1u96dtiEDI+U9QzYfRLpNYnv0zLuLX+7
KCAmvWmErDLXv1ngWmTo1feEjUN5yo+F1KtKAzUgXDZxxRnZ7mXmiIHfGf4JRZH03wgL7a2xxGpy
Ef56BpRQr+Zap1qydRCnTRdWVOhrmuZwTPdJBMPwlHiCKTTQnZoVpdIGJEGD4EP8z9e6Xuey9QrG
2XBy2e97rdfjfeRbgUS4eV0luDFNn5z9Ka6ZFjXjPqns5/ALegmnLb8wQ00ql8t9zvO4UjwB1uDa
b1Q2/8ptUsb+E7cA1WEfo4SNUo/LpjLqut/9oV/sC6dFQLE0ND9z6bTzXB226gjMc0OlwyR5PuZg
iz7Arghu/CsCGAfbEJbaWXmwVVLa/NrRL+wvacG121ock50O3gfhp7xvEqvzmCfHlnbyVxlz76t1
JP/hqC2Fc8FjPLW18i/ac1pPsQy3wd5u75ClNvfrc2JEaDPqxvmzTCE4tYugKW1tDwWIbqQY6+Uf
rZ6h2M4N9CT39t5Zz7J8J1pNeeO8uGke5+R+HYLsb+ff72hP7b1cnrPpMMPw2eIXrnj/wPkz8W0b
/QVxw5tGgks+xmePMbm3thQA+9PsGAqQICLkf3UhAL7/g42NXoFWwm8gW++rQNIuznnaHRgg30iF
lU8IWWY+S8kEAp4giZKPM4RoE0sJYUQgBqSUeVgx+EH4ArE0S24h1+Ob8kh2RLdDvOd9t0nDH+JP
sV6PvSGIOMEhZbymyONuSw0zs3I/djdZht5SNJRvD1gqaJ5GbALdZLBqEnF3DbMh4p/3S559hG6l
dNQba0rPRbmrpLlsxz2B57y1GrMGOijwMZAcL6wGF7UB+gQJTM0mkOYzkn2LtVxfp0WbU963MGHC
KgcoxZeLZO/PsMXQsv8vCFclVh+zzezkrgjJbnUjaRA786b6P9wXzTj6KMu8jNed9Q1MP5fWGEOz
hcxsj1OMDYWe+RhpfTxh+NAOZi/8N9mJ7PCZTq3rWRm0x0Zp1rOfqS4YM4/86YbeKkKlOMJkAiiF
kHsxav4ETzb1HYsN/Lj7DocXe2a8CPgdegXYjGwTjFwlG7PtcCiWOVDXp35axfXBSS7fOREQV+Oy
Aa0KU1AyNi2Gf5v6kjVLf72njZg5lZ3m1PZy1/3K+VK1jQV3tWQxvkMcgDo+E8uGzx9YXL0rJ5v9
7Iw2U4215HzyH9eogMzIKD4BfQRSkqU2RIpAZAEF9B4k+ImMpb3rro+hC1IEB1Pk5scg2XB0l8Hj
P1Fkk0Tvbwl/DmYhDeBLIZBZMeldTCCD5nXgYJGxOnhtaqxjxOaaOZILJR/PDHbQfCGlE0YzaYLU
3rbkbcRAMXSmhnlb19ARRK09h6iqefl/0pvwHjC/uM9Bi5mztBz+tMSv0IQ1rvZyRm9rUEGehMLf
M1AccwUkDewTgjcO9mrrklNP+1OzVpJyHyJnX0gMzx66mqnIxmEQKd0V+Cggx2W4EPlCCg7Nbui5
/8O4aXsxmnp7lj7TQpCvRJRypP96jtRD+CNcBZb7o7GgZ6PET3+6rkfXJmfq5w8/mIIKPEIKbsv3
IgjIvExmnv69A9YJTQ0vy7yRKjbf28OIK0mZ5IjKoaK+fsvZMa7ZhsomjjdrMlpw2sTEDKZzQ9OZ
khE/I5q2Rb7XWXXwJ8A2y8PP586L7LB8WhHCMAHKShJJvqC0Td0rXkyQcQCzjILRr3Rky+pXbgGT
EgBfPZnFW9NciZfMX9b/mhJlXIbWS27Pfl/CKqmWxlXEuFQ+fIn0hhAXH37iJ6IDlPQH3XPWBu1f
8TPJNtyZxgLPlRub7+Ljf6PFvoFjU9j9Uw/X5SQUigOu0ihBc9fUrZe9kgALP0EhYHRlwuL447qR
JdCIAzoaCMl+yP1u6cN1PT9gaRHsXtblSZvobwimq3oRKpPTvz3PHUkJzkEWfSP9VhhzFi70T436
BO4/thxU+pRU9XUHQhEvneBlnTX5tzvrifxBca/QGE/Il2UmkPmeqxasw3G1+794Lg92X44vUPcg
c6NgSRC1K9TUUIXs4VgcCSHRqlV0/1n55iiLS4tc7WRaS/4cVsyRmTeUfAIwhHJXpBq5I75Ujt2h
8LoYUNeup8Ce5GlTf89vOFLK+QOi64G76rN1Kf4KLBb6dDcbGjbvyeYWgNVD6nW9JYGNuhtUwsaA
cAeg2bqRYmCM+Cj3lUkm9G99tTunRLrVIOZF9Ojxhb+vAHkIixwji8dnW5+VlvxsGbkCXjwAW3Tb
rsWKLLG6wkUXJZEmeXpq5qIgNEtodPpk6vgUkvMMLpfla+C9oqumXvRxTu3NFfQsGWFQEh+vDaVW
I2C5VPCwHfTbaiHyGv5igPHtgpRsw62aD9IGk6lqvF2xf4KlgBFY+Pc3pDXxd8HeDPa+T7pJEMs9
1r7M2oOn2QRmX4l1cY0MzlCALdH82MiOlt//Gafjn5a8L/U7Rud7lptFstZflrHw5CAwiN94iAv3
cvoxXRsLcdy/b3ScW5NK3Yapy8grBM5ifOcuMvZRMfRb/nO0dVJw9FiSTTiemSZPW8ON04TNDf9O
y1blXU5/hPZWjyD4z9uluqJUyGEMESiHFiY03OmEGyR4+xj3LGPLzH08M3oco/juUayVn+OF/+2/
z71lfsxS06VdEaZihxDqlv7i7XxUhgqY0K0BkVQnhgcjeQUFLVTpY4sveUsipXN8DwNNoA56Ldrc
rPhKqrl9iJStVB1eL7GYu7cJqCXF2hWGtvwiqrnrhc+JH62Sm3/T1xvknNq0ljjqkYG+edXlITEE
Wneyq09UJD8f8/FOLoQzcV+au4erYlGy+I6FqHfwmgOr6Hgwn4FKM0ZLad5imybgROeu+HtAVpBK
jHYZJlDtLhcUAwR6iiUsUtPFY5SD7DRABouSiAiVL+lHjqetQdDq6S+6Hhnfyk11JC3dU/IKSp/9
jUi19L8MHqUPCXab1XL0HkTB6kuA/TC7CgMvwK4JHuPITkEY+Z5m6CtgtE0gFESCtnHOtvtsE1Dt
LexpbnhgUoMNTxgeCE9V/nh+v15dLspKBrDD2P4C7hRbc7OTxUjzRt8UxLAvI8V7CYQ2AKw6ph7x
5G8zKwfRd0e8Z5S9U4cURT2h/qALjCVjJOdMfBaHA0hEM+ca/oIX5nkaNjv5bcm34SBnOpqZGQn2
7IUnRHdzg+vhsh5z0z1HnMLjp0Qy+2w+AYS8g+bq+XZ6AIJJ8m1B2Enwwa4gHMdnmMGJH+WXejf1
87Gz+KhcLXwjJNMaSk8UIPwsYzRyu8KkI2yZsUWfeqLJYP03Z8Vpko4xI+lKIe5kke3QASf3Ltrn
vgGO7xk4kFIWzyeKD3xIx1KlnjgeiJz39eoKiq+q4vQNABKdzlDjIVfZqgBvBPLoxRLlrBNgXHeR
/LyPoRkcYQFkDuCewtIdNCwPctIY8wJbxnjzSG34MjKWWVw1ZfBVvAXwAA3DTirsVw8C4HEyZBFK
y71BYxfUXttrSHIbog/k40w7JuW4bIj+mHlgO3CINP4Hbrh/Vo0QrHaOdEVMAFKRb2ug9FNdAb8j
D+oPa564sHffmXpAxlsEfizK0+JNIOYOda0eFNKIVa0Ywa/ZfsYvh8FUk0PYRJAEudazzZDG8CPb
W5dP5SqcEj08fYVlixo33dJLty809HDxD+aV9DrDZTmagPWu2LhSSTa7cQUfXqXzAyoFnkQNzvoG
eK4cnACMTbaY1ApAa3S7+8qfQHKamctwNEzIan/MDDvZFwX4n64B8MPNm7OiCiUGOk2CNuKz7bOA
e4RJpUjhQ8h59YEeS+EyO9FpuZOekTta6GuCnLzHjJcVlmbdv9ny1YkgZp3DgEFDtpqV6CtlUclb
114c+zKOf7NkRHvA8RwYiVCKasYvTOrKnnKkB+bQslOYyGrsLU7+b9nV7MnEHwcnlNoAIrUQlDGC
1kTqEnh/6vsUtiNj4Vefku3R2v7o6oZku9hVOFplEdfNNpg75uJbWmywzP6AcFlY+aRmzWNXht2Q
WAZUoX0C86TL97xKiKBukCSPtJzS/LjL4SUn1tlMjXSSQ2E8/IbiBDn2uxD8/j19QWJIVyKossLa
438d8mamyHB/Lip4NwmVfpVDTb3qbMcc6INw7L+wUEiFLd2h4twKbBL3c2/4bTPkOEE57AtUaBwx
4rQ0FcZQ4iCYurWhdLEEJ0TpKDGpIHpsCKUsslF5i+Giw7HUcu2B1Z8Ibf3JQ4okAYAGvOD+bWRQ
MqC26MCJvkZ2u5IEIpOabAuJYTib7rBBOsxiFg8mRbXAOSj2J+cpZHrRbcqYt8En64jZTHZhGP2g
NYINdTwM+22v5MdblZSC5XR4gK/3PSsRf5GI8h+BrnoAxenz5rj0zl6Xoj3D4sQOd80ME6MYxsJF
jNoVRgv1NO3QUtNmcknGzUddHYUKT0ZpkCzSpsY5/OocF+6yV4yZVED2idPilzjbCplV5nUqwbO7
yFYr2kno6HcTkwWG9Ul7RTc0tIuAKfl2WIedWhz8Hn/3K4vaUzUoY9chJLvUBybW0CextCftP96u
lMc3FKUI7lR9xLRBGS87itnboVD3aFIUY0RBZbbqVz9vAA/mq9MhV28OXP23s4JuYbebaPCBaac6
NdUA5MDuGziLlcY2Vnl6LqD+y/34vc8t3o1bVTZJZQSpvzCOLncd2pWIpeQ10WfqZ8eCYfEVhWVy
vIHaYUIOR3JGwGbHj6wTZGRYtxhCgOqTa9p+ExKufE1N2RTVhg/paptmufoBH+aj9Ufk76BQ9RFW
Fwq002MVvmasjV+rF816h3kG4LoQMHBT46/NSCMxyxAGHe+J20tz9sOqwhhyKn4HSsIQ05Y1Q7vl
DC4kf+u0+Rj78DSV2RJBWdJK1YcwYRhavvKqFa2ZMdlCQ0/IhRCZA8W8JuNmZ1b2Yci92PmtED9y
QauVe0W0xIZNHqjx5ZvYJ9vwEzr32BQTYcY296vwu5l9JBAFuLWuMx3GS8Zf/NnK5iCeWd/wrn/Z
hqHy2oCW8hfJiTNZjDRSUCnIJdjLFIzGigntEJTcmBX7NHs4Es9ooY8wblZcmY3SZHyjosSMIypx
GknCaph0VxPfBhmg5o4RgT3T/YXr5J/MkMH/KH8OemB3zTqurCGOgH3IHJUVzZscpjTB9IdczOS2
4xONVLaR6DI+8RF/IPI27R1a+tjhGGxUDkcYRWxOiBsIL/iIymfntnHIWcbC9IGCGACK2oPzy9nD
JBjbFequQYby9K5tg7oKZHhcpCp22AXmMNpWTg/WXHn0cCco1BbnzxKGyecb21RD3R14NRQA53h6
AwP+uPjVlILtDdcgvBxOvm3ESv75giRmMnBI8mWweomeLszwwF8A2irpFlFHYj80aWcqGEqTQCOl
86xPLgnDXUfBL1FXBGeL+8EX09Ee6l6+iptxdDgn7MYqCpujjQe8CAB/Zo9i0hhhHg8HWEP34WN9
gkAbJ4wF+alz8Tg8jt5hgauEf9QllRDfUeWc9nf4EXy2xrRkqnPGa6vNAy+HVYnCKzbueZUbHTvA
8VZW8DIXzErh1w6NnzFq1ZzBPtn13YHpe7Bob9uINw9mzQFSVyw1lGCIo5Q5SlJpgzmpLGQKqSIJ
tMDR+2XNpK6/EBOWocC7EFE25YVekE49cUitq484SdYKT0zXq4KiZGeM6xWpiELGNqQlIOltNZqY
cCtQs/6hfKlYdrIOqJQ69USbXphP40xHn7yGvwvqsWt/59v1kpwBy6kZjPn3l3LPHyOeS86Lt2fr
q+DDA8bS5NVpM6TXJu1zdIjwyr2hmvnF7ydKnhjgueeGr0u/YAZ/ABKrNPTVW4YLRCoHfIUzo/ve
KCoYlZKNy8VvN+BDY5enDj/s5lJNJL9iaGL0sNE32dh7BcvIZFKXDJ1cCahHi/iSKk9i4ngF3g98
KJn0oH2tVWCXGjtgeW9X0OXE1pRX1BNwjDc+ABSeN8J0weHbY4ReAWeCyjB8jA4OR/wjiRsL9PhY
WNnzte8Ld3M/0U7wQUKGqfcpyX+ZMxyc6OUr/ui/WviiSEgXCwOReQ1iLXvfL/gEceWwtNMBJtj8
LXM29rWIGyTYiQRWphZ/wBdA6TS+88R3dThzyFXTsyNc0pGkxYoZ9jsjgvLMTOb26xNTD999WENa
DGKiOuSBMOIcWefsIcs86cHmy7mHCOrtvG/OkQBXWiKIAHcu6fX9F8u+VgmrMM+rlA0aFe3HHsyz
8eMj0dNBdAoHa8QehfCEf4hgHOVC6sXxeEciSMgGkZW0EReg17snL+zSPcgpDiZvKYVe8I4J+ie4
YMo2bZszw/22P9o1QdUsgAnw0up6ydkr0kS7oO8demOUESKv3IFf9VXqcu/qMIEX4iFdqn96yP54
HXeg0tRVs1Xwo/VkQ3zq2KkLUH0razpFvHWK8+rNWBldL2fxHyMF7vQf2ldrBbDCUTC85xd6Lae9
29pl+EFYKowZWDjD0QXCDVMVVZPsybDO8s/RtOeATDMdYp1ZgfaowX4UVo05ylDk0xf+ZZeNztr4
7UDYDkOS9smu84QdSPrfhwZLgyx2UjPb+p+bCmuXD0a5TGrp1W/2J6eqRA==
`protect end_protected

