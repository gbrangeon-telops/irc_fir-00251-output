

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gQ4CxdvWgnieRLRQ2AMwpJaA+X4QUP23A7mcpTzLH1nina2JWDwyro/SbR0koY81VxQ8tVNBYSg8
3s+EjSEjvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gPnHmBrjBHDleV2Jfu7AAgNyinLiMa4GswbueiHBD8y67DvELbF4ryETXsYzyyRC60JDgiQTY9xS
mNBL0n+tguqX8nripcl2WvUcK2rEIU4vEmrY5Xa0k52V9uCE29ruqODz0JXngqZvaosAn7R3hB73
7cI2IgLWPL6sayUHq1M=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bim7wErRMWV5FSeSCuJLdGVUUYEH+U9HzwEGlgElmMU1LE1rxBL3MWBw6E1Qg5kGmxPZcrNQKg7b
PLZUD5Dv3VyvXW/HR3jI7P5DnwdmPcuCjrrkZwCh4jjzor7rIj0AM8ubprUHwkpicj6rKGNYRGRi
+lmT6hjwlretXlYwE1YClKFDSDei0UBfS9a5tRfCcNpmoCaImXf0uTOJ8unbujREQZSIp1snYBqM
Q6qvNMpDqcLoVSU7OrgHQdnonXWYqY/ILDCjdL1o02B+xcnkuGf+oGCDs8KSCPuzYvirbLqI8N91
feufkvRKEcc9+CQ7U9kVuEQ2Z+MB8XwJtiWwVA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HhRynIQ+TRImN/1ISEgCruTQGOfZ7yQ0AeSPRr1UgeSXeBV4/j+sqUVwy6KpjxjyOB8/Up1pUaXk
C62p4kvtT61bX2llnNuuYjikfaIxGUWJ2S1a+GpileS7Ui7iwtZy8qreshTy7qb9L+4SycH2S0Vs
ofqZzZCA27OgdUdAA0M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RhnO7aE6HcfX9+ngWNOvpaRDGHOLotkXich9kwwYcDEBAwcff538vS/s9YC3iM7OnnDBzfIjK9PG
hZTnV6Wbh+heW3iD6MhhmPxC3a+3h3Xr7G6V/gV+8tP3qbjwLdyiI3Y3Tl9GXzeddtSNdvaD6764
1AS1CtRtG1cyGvfnXyGxmyDzJ91rqIOqSJbBOVjL0a+NolFyEU0BYVthKlZ39r7JI1kVtcM5XAND
LnFrRp5p6iEzVZDFdricPTs3V2FwNDnZSvZ0QADHlENUl1ofRaFRtXOEIahTDRwJJzBMRTba/K/s
3AtKBuzpWzTyvSqo+1PWwgrrClt60fAvHko0Yg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12608)
`protect data_block
Hx6lQiyT4Q2KXSxeMxtyzjCY+izU6u0vHCbcQhyGQFpwmko14NXEMDtJsnP3gFgvfsMKbR/V5Qw+
uZQ5U6Gi/5FRCPfdStLclQ0+I+mSAff644FlIXcJzX2xC5Gf9/vcBJigWJyw3IIsbExwDlcP1PRi
aT7H6m3+vnlY+4EXI1YFGkXMYOznJuV3JLE4mUedd5HPiZkoYtkI0FhfcyQbCdUk7wwELCXN/UcY
8OwWvVsXIkvImBay++wUCNGK0Vv2MiIRqdEjHELV5+lT4yJDDufejAJlq+bTZIuU4hr5wW//u/MK
z1Spl+M83WU2UUUbw14zKqmNo+3z47ybwrrHTgdWm5eevGc3JmIK6+xACotDLaDNoXtPCS+ZGRwH
12svpAs4EX7E7T/wZx02foLSdLutvvl7nxhAifkoFHdT0GlIPKJ4j7Fwei0tCWlF1f27stN34Lxf
wQOSGuM8RuBmYhpHcCY5fGWhX5yaHAYMPUNxISASlBlVUL6TZdZ0Avfamq//FPvvNqLlCIQLhPUt
Bc8GuOAgCh6LbKwxOhRQV636ih265Xgt/AGtZpCvoMZeBxF5gyKv1ttLTJSzAN+jKmNL/037h6XT
2EyhG+GbSSjNgGJnvDVuDCyRfo5D5x+Uxz7S+1Q7a31O/QVOGH8HV9BrHDz17ORcowliODquXuqp
gKK8NHSqXlPZ2CqL97AydoXkPc7RfMYn/GmOWEQHP0HGX3faqK6QwEqHVGiAtRV0SS74Lv6iADI9
WCdMZKEQEiNEqV8tduSNEgArLvqq9GkNRs7322eyq3th8eZo99yLmYw9Om8u9jT03qF4kyhcx/cV
vsUh0XbgqHAeH0OFULmWDtC24z3WyJ4g+2eIXXuO6sIpURImy+ZK44C/wPXA+CgYysenwvpfxWbn
uhOUU7YsAgSD17RdCoKgJJYOLDz+vtG8gZFV5Y8jSIHnscny9M0tHJT5VEAQZoEBb3Y5wI41xWK8
wiXBGsCPFkeEkWbyxe7AYF06m8xkMiti7AJaAK93scKoQG6aT5C64FDRKVki33PQSXnqf8KZ+M55
yarh0VlLm93VAyYxlSDUedRJ2cpvwDqNHZExYpP7qspZyKoOm2zuj/gvA9fWFeiJmbn0xL3BotbC
UpfBMb0BH5YrKxU425ihOKmGnflZKSP3FvqBIELa1fExDCTP9pvgf8a/E1rEUkd5kr7sMVi6L7bp
V/OzK43+81qx6bKEkIb8QD1CkF3VJn2HF1nUxpPuERC7Ud5nR29/oFBe1Y6Aa8UvDUPr85nnis/l
oNw+a0yn5Os6CHfz7B8vQOospVOjz1cT88rO5nNeGK5Sfcyu8J1jv7VH7gbm45kaVJr2ob2yIgP7
FIT6WC6SGYj9x6thUCUyylPX2t7yveUW2dnKnwJan2CZE9hWc3k3xwRyXiun4DUON6UhAhHVfpTB
bQVt4XUWiXP45AMq9wwyoXWqW2/qR9WqXacwDNNbmSWalD3zxA/xQW1EzYFaF7/0n6cgvIq1lOIH
lPqDJHFZQzwhBuksALfr6+SwMcS0Zb2OOnXMT+RHDtKuGWY72JahRv9Dzqvm3445eqEQ38QUZaij
ZRMBX5ufVYNPDyDs2bGP+w95syRTIGZJrJui5PRN/8Yv9o2PRMFC/V3T4RcMyp2y7JnaDO7xiqao
QoyaHm0U42ox9SuzcfsSl1k8oB1FeMV7hsf8CHjTYAaiXZNrKZLJPpMeMP3dlxteWgBmm8oFUiMd
kaQaencT6qCjHyqR+NNQtfzPVLhhM3GtrVUT0f0JOIFXCMEA/xxgKRHEOrAKAzJMPJhn3yJ2Jayh
F0NraRN8cPC9SYhXKRiSDAgS/RaFiC2/UNEU2FkhMOloPVTPaTstHIKRgTUgRjRKdyMM8XcpbXmi
cX/u1Km1Iu8HTqMf57AC/GZ7t9/FzEiQmxRXY1n985ktTbzO/nXOsU5AiAvZ3aOT7YGLn8cqzS5/
+oDU9OX4nu4p8FiLKBdJljLcC4DvITSryIfGthaTKNzhamqrj8rtRICi+CiXt04Ait2ErJa80aaJ
QyLHa9+7O9x4sB1gF+vsNaKeVjoZydn3tsk7lkeAGL03JNBx6BWe9j6Cpl05o2C3Kfwm3vBeKOOl
gD0NOmjIeH674fcKcdh5XVFhr9iOI9Vka3/fWgPrznLhdgBIrKFu/+eh4Mp8g7H8ydR4FQcfuFhZ
xxrk2Nq6GRApIHBy+6x6gI+71cRd6nkdgDv8PqSdJUy3n2ktX+dGhIN44+cuqdhRHEKeK8PGdvrZ
/UKxHnDhYgZJxcZzXmcwYjx5pGFHoDWw6XGOPhNW5zlRLfY2dvSjBWBYu+/pjzYla+PiCmf5HNFL
SXQW22S9YEXsm55/gwZM3Scuhuz0+NGVfC032pS2nvOVtiGn17wabYP37rh/B1i+pgHDEl7a22W3
ZQL8V0lcaq2RCDdSbmfMf1wMO2Xjfy57RGVlO4vhAfUTq7ayI2LrfN4rRvDjy2uCeQYreSqgDNkf
LUrop6pUMwHNTR+6WevFraITIIgvPTNA4HFd9D92JdnuQz/8mM8p+Un54UiCMpdCKwfEDrHplAR9
0ZXVZ8KhAbuKRnO+q0s1tTHVer4R2xoCB3TuFdpTHUOIzxn7sRBCSfDWKZvYehaVNFkrC7jH/8YH
18ol3007zon/BfN/mg62WSjSgIVrtqu3NQLztjTbsWUZSOySaMASEQ1pa2PSoXiMGuN3p7MTTy8W
8Ykf6kHSGfauQubnp6BQmBaSYgci3oohzvq/f2DYqwJmJFtn4GNlXwpQeRVpaam5egb8hNlb80Ao
gtKbY11Y1LpIqmud+hPIm+WDBElhS0zS4Wvh9a1zf0SKnLbLGu90TL8m33LY4vLcspfpojJw2H8K
5/6WZqFdKl8O4BnRyYpALnjaJFwifnlcomU1QjS0pXe2r9yT1nCqt0RJwx7kbUmm6d76cz2/MMy4
Z732MCa0ZlQkAFAaxQsmftYmuo1N2vfuo01O0bY3kX8JXjebwc0l/+cZovx4gypyiFlIqVufz/hi
IdGKM/5Y2beYHaRJ0Tof43tz7e/AwyGQVCTQ8VOQgE7mA4runWk3o7opsTszqdEGzM0i+V5h53so
lLaA8Dn0P+Rz0pQXikwhzWJfBM7fn8gZNiGUyVvqZWXSWxM5BWzlqzq4Gyag+BEwygXPQKRhhcR0
rYLl/Aj0rljA6OlELe4z1qhd9h1qZkJ1YOpRGdyl8GVAChdJBqjejPc/xi9Dxs8kqtIOT5hdr6G+
n0BE6SLEpc95s5n0M+Kp06eZxzRpTlJrw0b8pKDfa9/TdCHaQVufnnvztrFp6Q4J65CyAWrDv73C
jQ73FQMZIs/XS8d73EoYMrtU6JcEMnLvjP7rxhVLuvmt/rfes2Yse5LjJ+e9LXg6bRS9mNDwqoWr
vnp0Xdjj+XkHIAEkaqbg8oH25tAO2r5k5XhKzq2FWybewInJ37BjS8hOq05zV1XGFsMLsvDmo+2w
mi4R26Pd52CkT69C21KuzzTyIqIpQGYDmZ+MxJqUiwPCMqfWxPvmTB4gpbOWZG+HkUV9b4TtMQmm
kf46EtF4q5bZ8zS31Lld1jslHCY+/payevXFwXYlE8EPyUWM9Hz2ct7gJMRQAqpcQVD+n0U5SRmm
svCB7zRzXpSmMKufPls10ILvOZ1F7sa0ErBUcoJQgPJmUPMTYUZCaVDkcb7YFZdbD3ZzIZb7vD7I
Unk6Sxm69BXK6E4nBfp/6BwPQv9ePsxXYt5ZwjDoC6TrWYJ+b0iErjBzKVQSET31RNzAk8uknNkJ
gsLhcxdBBoJ/j4t/Pp9xU4QbP4dNyb+OlIAf2QnSQsiEHzFwbr/koEMzZBj/y7pqERJbNLKCHeFF
AOWOImeMqVCmjJ3slT4H8p6TbVeUUZi6HYAjb2oH0jNzJjlm1jyy9JsT15CxQ0zuVnyaub2Qno5c
2kSmmIg/k48arZxwE5sCVOqofWtm90mlJw3w8BfP+NdxWKqJ7TylxJgAwfqo4TyXUuf3muRVZYuY
BCxkJzVXYXSgHjIzzf9FnKde/h1qvjRfVgZNujv0jHRPoRX1boogi/ZYzMk4klyw85VlD16lYEv3
wlOsDLB7PHnabc1t16pUKISjkryxda7ymg12P3k4vsB17MKk3sPVZvwbkKDeel9+XOIBh9FeOBLC
Z/tE8um2ZEiW3wbyosHEkW2vOgovjT/uEOh0RiIUj54DXiJWkwKcKhdfbIsgVe+wHYytWxcFOnWA
xINDQaukXnrQETLtlZi7aN9yAfB6mkyGmclqck+AwdjZQecGYih4l8SAHl0UxDYh3RQCFHXfAMx3
76djReUphFjkLCbifXE4SHtq7qumazgFE/dV7dsTMLw7FrEvl0qTVM1K4ktjvERdi0S2n03AFYlv
fpEWukq+kJivxbaskTVw9BU3j5ZL6tyBGiPxJNciCxt4zNQ4i+IT5GSHgcuxOIGFJPYU/DfEkxlL
KCM2IjPbGXAXZWlrAi7Br9oD2r+nITti8l+uKL6jEnkvynhUQszm1lUrrRSB8LOPcmRj1hTD7EX0
LIK0NdtAx0BQdayKi/e4G6V1HLGphXP5/8PAjZ55YU40uQocXxyHws/LtSJmX1boSWykDvMH738I
pZRd8AQySucIjvHBNNiTbKWqP3Md7B//6nBWuam0+LPTR9mglXvUsiEubt/urnevwONYCBmTZyya
Xz+ZinVve/CoE2va+uluQc7fKlSAyfvOO90HfMSjYlg9FawPYZYNsK/yad9Mqg+wMtBV1nWGfqCS
JlAkUca6F++7WeUC4062vR1kWhBgx/I5l2bMj1fOEQukk0g0iUK+fSAQfvSiOXHxmnvYMwQ2ZrUs
t5WSsvjJPhRP2XMazCzuYqiXNpoQPbqJ7b4bJXuKb2kKjjqjcqOsJgCZxPAQ9NKzH076zmuhHWCd
/mhk8hI9HSrId0EVdjn/CIv2UnBS8fVo6eEloGebCp/O53ef3Phqcbztx+/vigg76BcEiVPkPGXM
TncOCwSHw5o+6FhAaE458IykPy1TMnhSeY2keUjvlMZfeiOAGb+Ae9NDdDlgF2VdmB+qR6Q16H5O
26apjWj5tBjcqlC0Lce/B4FvlRbAo7JeAtlBgzgOJ7aveGtdzdeUHWNsXy9xFdtDcOF+mZp8JUQO
GLr2BNiiNANMbMlrxL+gaEMXwQeqRqc8n3b3hKCSrwesXSvoPz2Sij/GVRmsg0cSpmPWMcf1QOUG
HFyg2wn5GPa0Q3U0b5d/1UEdTh6GINAIYWg0zxMMzZ5zfBY65kgOebf7PNRRZ4U1rQLTyImqFj/h
nVZ9LO9s6M+515jxrN3zioIyS2nSqDOTV3OxK0OcId/a4J3PE2QbwGCbYpGgPlgtpHmuOAQCbSBb
pcfAeZrYM29meGAKfU+xsF5AtijNjtibbYkD29Iv4mb+m1Kz7hn/a1GLvaDwrA+dD7sf0k1AU3zM
lQNeEoqSKujrJ7Wnqubh4uUrIhsXKlE22YvxonFoCXmAJ7xUUdywb4VE+Ad8h1XG2wktmWCNfxTg
u+Vt4z1F1FI5OauffHBJ3/Cq/20RyIf1BsI0bHuKCjqijF4M0W7jLKJZIHQP1oP1Udp4Slhe94+5
dTg8iJAqed1h2wsYt2yiDCdXxDUZJi+BVY2yWzpa9rn/cRFs+pzWPeBjwhKwjSMPGNqhw9zN86wr
1TGALJdVsvyVbzygkPN9pz7N8Ohn4rDARaQjA+lByDVEZ41vi5vQ5KkpOVVc64422uvWM/t9cgMh
mw6tBDYkrT0Dv9aizJzIEb7rfv//HHfyuNW69ls3fRWx+xwt0Ssbs4iYuQoeyjkacWXJTCdkr+ZF
px3IUt6pfz/ybaWwdwjWT6pLwSZN0k0kGv+HS59b8CqA7X+2P36k7NTJBb7KzW+MvlyF2VBC0dPa
npux690Ai39BHVotaZhdMZfwmLZZYrPxJbhGdAXbyItmBm5cvqKPu4ZyseQvVPUVgWX70mKchcmJ
xLI20PCf76GdWzhVrSlDnNYtad239UxAUjaoLuHdd6t0KItuJOVeLPCE2qu7+DVIU0/AL0+/61e3
8NnfgRrbw80KMdI5hrtrhQ8yw2SoZqa2wsGoPMkLE7cx74OVoFDw1kW+6Gf263Kkq7b1wLh5kbLB
mwAIl44oQbdiJ4zPGoyXhhEV5pQ+lEhSaaHJMu5DEis2y0DeN0vKUQu73GsYLr/l30nOfHtBRhw9
eWAXTBG0QepatIKHo9hRjPBrjRt9Csq3361d1iffZQQhtpQUCHKj2pKPTB5cV8wTTxEWgkHrnZvB
fQ7MtkPtDUIggQNqKj/KXxBibeBUjeavXmDRDluzG0IcgHhmIJZJE4YcbmtHX/bPybkGDImh2/4E
rMLWHElqETWLWXYO8zDZJH7rvbnYD/e1SSbNmlr5XI5N5ca6x6m48bF7zciJ7tzbjlHsktm2+cSW
PA1/WFEOo6NUOnaPkeWT/x7fIrk4FS5GtSa3pUd5UPuZ+8r+tMHJ8UF3Ei5uMH9t706f2T6wj7nT
Ipjo+okKRhM3SxCNH8Vo0PXDKpr6Vz9Xvlh9P2UPVpwjW2P8XFrIpJ9aQSsQVjqHaqSdYN+5NHIJ
WGopLK0Uoln0WXBDbS588tlWMYO6M0TGtDdjZthNNM03jBz6PxD2CJ0+jqh11WOd/jSzfPkXhnNp
M2EmUEGHt0xzPUVQghQqggDb7z/BGZqSMj0HAFSDrhUsTnDZ0zV0NnLgQXYA2xBBGKNFiWUqSeTu
tCx0Qx3Pcp9Oa8TFCko+OtWtmPT5RqLSYwnqSSaplfbd23T/6RxLqc/4fhsPQfn/X+FpLSWdJuYR
g7VUyB/ZNx6OmQYtkzUckoulb/Ios1IrYVjHiBt/ZJpO07YC6pDum+JgehBNd6RtLBC/JK3lpM3W
UvFzbmG26V4jhfBt/cBM6tiKJE8zSzpsAyo7gYuM5PY9bkyvllzPWpxY9Y9JIVXRnNatIHxKx3VE
K6b8A27gxsUfLCG0gdvyNmYIwEn0pQQLSbXIVOzIiY/Q1AglRSLx9sPQpz4G1WGBjTdYas5rbrL6
1xLIjly5nf8fNtMBJg2Rey0Wroq6LxExizNDtH2g5AsS1B75If/PAyk3xQEUQKFY1AMT6Fhap/JY
uY875AzY/xseOCl92DAGEPWiaLeNM2rmysuKCjc3KBD2Sf1opKBcHqOwrFKR8my9ybcXSOgwFWju
QeZvDKZLWL5WhzL2chzEZNQ5hrO7BV+pXeT+eiiyPFqLaObLI6dKdcSOuqybPJ5Yj4PbaLI5VVbB
ms0wC6UVtkCXprSiDOOJZ5zR3G/4V2c+Pn2rXwzVjx3W1iPaEFC0Is+q3UGtQ5yeFc6mNFXVM6SA
Be5EQbi0mdoFAQY7/p7LkGITytywk6mnkr5dtIubvyzpuBLLeOEaeRoBADGXFq4o2d6ASXcHrP6H
E6aMAacedB+YbK/+7Bc7XR/OECU+I8o+DK/xHz4TKWUP0DuFL7iXr7eRbAJVQyrrmy0jdEk2kkkE
XuNHA3eONLmADRP7lyBLM+nEbrFz7nxQ+KAMNsvrfgOexBlV5LeVbltK6TY5FKjgV1y4c+bACwzF
KHNSRmQILoAwHcCs39I63aziW3xqSbjX6+ffMFUfrzdI4MVnHY3VIAl76QnhDlXAh7HjhpvcECQc
jZoFX5YjyHlvSmFq/HfU4ZcTseZXo/k01WxF8eA39BF5VCTVFnOX6Yr6H5gdp02E4SWAfBHjXHUG
ZVo9XPXaqPivywWq6dt2vCVOlEy0dlv6hnXNDJWUE/BFGqw2jV32c8zcGOCoSNfbseujaNMYqAn9
/V9OBZK6QLz6BzYyCrghTusjmuKAWFJ9zy+2prNuVKb85jwKxW649myl8SLkIM1g0bsCMU4ZFHhI
/nw6lPmjXoq7CD6DTVmUaXW8WCq+UYqnfFbz5rOVvODRbdOKU+s6T2GiHXDQ3CHIFnYgZUoj6ndu
RD8/oHu3FOTbN8YfpxudD5XZT4jsRSr7sb+coWFzLH+e/mBPOF4ZhK7ohvCGzEwn+mFCYM7uSIQ6
DtAUkRPeeUNnqs0RnIbmHtkHYlZtegLMCVvTl4vtW+N1EfgRZMyWn88jbqTkwhTd4qlfpnN9yXgk
ifclvveBG7h3RnW4GRmK0xGSDL36oU5QlPJ99Uuv/gJvmqpLOnBPPkO+Tdrheo8wrPQpZuMBur7O
f0fMxolZutAkNcK2ha7oBoPT1vVtkwYU6e0xWpYHm4jVQ/OLCL+3U13NO35q3SjuwlE5wuf053fd
Txf97jwi10Jff2jjb7CmYTVasvC8WAMB6FbSuHXnfeP6nQ0KbMBU0ecrG3maBUk4acS2nC4j6W+K
M7TYy/L2ru1oO+IlU/WBl07YwCQcEKPZ2SZi6lm2ff1oDiaZLeItqPUmdw2gmFg0bs31UcD/qAJn
I6/KHt1ciwWkTDjDPd3WzJkfKGLZIyR1/kJDHI8E5emGvJXItrtvRH+DXmt4Yp0WzwgpCYV1LCC1
VlCliq4JEDeOHDm9mFkZLmv+KK7CmWBDtUGlfLSO/khCYeGSgBhEzo1ULotC3DQskZXu4NcJ6wkY
u7S1ThXCLcknf+VVZ8w7I0f49AvtolvffoxOa0MFhtW1IPXFGnnx81LOWyh128sv486IZcT5kHu/
/RlZCc3rNHxBywyUVMP282jBYIwfOEN6m6rbd8KO2GT+kqR/7B1ya3IdE7DjaAN3tk21pjfTGOed
fLTmrKuLgGg0cup79telC7IXlYP4ggIij14byk3/cK28SgsDO4tvI9iiPuV7peSXAgts+v+SY/w+
D724lKPuma3tghpLKOWfRnTjy5CuFvD4GYgjnu3+knypQU2xmNKRnW7k2N6Ncy0VW8hzoinysC85
fyubfd0pS0EBGq06KmuyC9St5YA6jdcBe9RbmYUFWruhdV11u+p0mx8JaO6Pd3opvvSgEpeKk8Tv
UDzCq4kZMEwabFS0L7TaIGPMsdjse0Ed6AHsmxkURQdPHGb6KlUB9vAi0WnCkKRd2PxwDf+aWvQV
mC5Pk+b7PH2kXr7JuIC8E2nzjJQBsq7TMqF3iBePcx0F4nX+YjZlou/Eq14bIdFntq58qs0tKAkM
RKJThVg+rwbVP+9uDyCH0jfgKWAFYBAJUet66wiNfmpellUgSBwUKTrUZa53O3ZLp4qjp5y2w3Kk
nDxRCgMKqNCo7P21gnq2bLJq6Q4awVXJ+H/mlxaWe2mdMXlGsXJogIY5RGtP5g7F1jrfLVgQAr5v
EQUZPxudIlZh3z29h6gvZZE3dGYF847H0A2PEhlb30txbZsE62jImFA5eV3R7HMvDGOyiWelKajy
oAzIkZQSiZBAVbkRy2GlsQMYQE/9U0Ur5Roa8AAULv6J30+ofLR/gH1B8HOuzq1U45n6wH5idxIu
4GgVqQXwNOcChfyPl6um+rBQqx3H9br9/jN7Nd5wLHP8nhsu1TvcvrwA8ZzhRcrtJnSMPScFayx6
/IDcZtnd66jRnf/sxKhOVnXEeNjumttzJowIwKvPTFfdFJ+MOtg4Ww4l+O3L4z/kN3JxgxIQ0t47
E4laoxiS0YqneM/gIHOhwr2dXa6RZ4+mQeqIl6cdx8w6mYKHrf71p9jJ8PZfvbl7lDx7Jwh74Xyy
kmXgA2tK9cIT3DKYn8LO4YMSvQQyePtFhcUt5Yfa8XLHfEehHHbSm6tlJR1/jZUegVk2UcH8WWgZ
RyxufVHRNrHK66m0WwqjlLQ1pAFDPY3BaRWdZ16XfJ+vpAC7huuxFF1iOfaumHSKE6qYb+jWMjoy
oa6Pw3lYUtT+48qt1JlDr+IGdMGw5TQeBO/f8FgI5ZBI4QYN5OmIrRbbSo0aOLDDQ0CGcEnPold/
rReWZFxlCp4v1j7Hjz54PGVKpyKlYDbOEhMIn8Gy5CtMGPYtR6mKNB6O0cq5QVJqidbsKi9SEFlU
DXk3F56U8MuWigUyNN3DcyTqTGd5odkeFjSId8gcXevj9bUMcvCuVo3PQODk/n28efdvlz4976je
qLNmOZ+4nLxVOQn/aIjdy1Hw7p0eFhYQAUQ86eQyEUIldgJW8nUMM38dS2c96RAoMnOe9WwKKDcp
Lhddu0WymmPsaEDse9FoFXrqKRN6cU+jWv3fkuYAAfJG87jUm5boEinGBn70/Ah/z3/pZnuy1vqF
paLiQWuDRjS3gcGer7LLhuzi+E4lTbCXRHmrzf5QTjFcXBg+Lx++HFTShTcXcsz8aJ7LRh5LOHzq
M6y0yChIiGQpHwlAf4P+KdJvNAU5BZ1u0nBiUm27sEH1HoKiRgiESIcVdTLSYB9k9R2mXrYf4CUC
e548aTzcncz1pf7AxXHEJSGJVgcTm3zxkrwb31qShATOdiALy6Z9QYi7pwBrXvcG83sC5/Zb7XFq
LcUU0FgWU2SaY0l6+tF9x7i1jQ2N2MN90u4QBPEAuZIEGF3CjUMiZVbsZmWSZTgbLfcRk1GWBKYU
VhhfQTsOP0ZgWHnYjvkFMYjfnH57atkz6Gb52an+kdI8AMBvXL/7fDwCX0oIxiDJza4F4mRSMleZ
rsiVghi3lQFkH+4O3WCmF6ob17hhesEG5vPFdtxDDpeC9sX6mYNAfNPePZJLZjZMdGAFIqTd9IkW
fKv9j9AFzAkYjL2KNnD8zAYiFnfqklrOYGL8c79rhf0Y29ruFlE6O6PWQ5CLLw87VTu0LdWHMETv
u/biHImUg4gXw3+/sUDhxg3srNfgYro05cJLJG5yibae75QBOSrajaCzewMETY8QRnUcC8HtT9rD
IDvC4hZViRahZJQj75+6xtu+99cQE9Qd0fbfGF5QmNKlnT+pLZv2fmuOsi1HpeIx+R4pSHyRLu3A
35CHyESHhuxmbIfCIxJVGw6jZfwAmvhXC4cmd+HV+Uv9dLCX6b6IuVT5LoY0whTSvcOLNu1zvh0x
pBXkqmf6l0OwKmssd136jqWl0gHXKqSOFIn6UKfJgkaVqpkPTuyo4WKzVGRD7VO5u6XCPcE8QyVl
jk9vshXldGKI6kib5pLEpgBQRbMAjp3ju/EyKjSaAjIY8DQRDlZKN/geEMeeBxYXf39p7CutfUVK
ADYjVqgdMzd7Freqv3tDqvotn85Cg5jb1qW+RssKS9ZmXo6IaSjsv7+rPxPh+CS44M43BYP3V+XP
Jwj7fvmR7Qadv0ibqoOgD9CT5gP7Fncjn7+XS4hMwtQ9BeCD/2GS61f4DB2Fx7IxzorMdoCzvCaP
mbbMIfSgCHWS7MLblOkZITdgaMbPmx4WLsTHDLNKe6muSonmUHI12Ci06vn1tpxjDf7mHsKVxQ9n
TM9s5IzqWzi0erIFIty4YHYTPleg9TNkFqM3A9UqpYAWi2HenEfUfqyaMCeXhDN17EP13DlM6Gcf
UrXgaHqkdid9UeoXItqFITcdbE+SMtTZB/zN1wyr8y1bDP5/rcAyBkPPaMrh0c7uMAH2h67iBClI
mAIYiP1DEUceh7YL2QVrimNmiQybS+nMJoam1tyDPWpiIMBUCQ89EM5tXQGqKx9BNfyxRfndWUhT
LEi09FdCiUof85UB6o91c2rj1+4bU2UQiMjggt3WzY2+5tkx+iKh9JOOZM7yhMUTqxTNq+aEUBsV
M2OanNOl9reIc22IhRXhhgI+vc0us/q4wDROy6P16nnBt6MuGmigf8aWMXQhmMiVUCV43VuezLlq
xGgYxfSlCakUjqLOp6KKjUfCGMqQIQ7OU5m81idW7eK7e5TiuB1HSwxrO72c1NizoYq6L4o0nCcd
wnt6jydCaWO0XowoCi5ieqw9VX/+94xnk3ZkdNRgzM23dlMr78n7UC2UF94D5x3AT31Zo3WTY2ED
0rWRG4CSBhLZZiXEL055q/VhkxhmjlbzR8wpPd0S1Eu8Qf2rsfWh+XfsKCGmIqHNAUs0+eK3JwsR
r1e/R7a3whNFR9tv/vFhE9yvXrRLQB4LLBkSJ9VnHseeC6hRL0X72TZQNOGAnm2WUj2edc5fI3kG
w9uu3fw1BBIybpxI+XG/oBt7U+5+PXRNi7ZH5KHBe/SxcptS5kZ97dMLCWDNBVjiMuVbrg0rMCv3
eruvw4PShD1N20CKA2LCH3Brf+80UDk+5KGaYLUgV7DMppSFyc72Hzm09KwTMaqfE3ljcMeW1aSk
B32NgfXzUBkVL/A9+iPjqBtfAkToTtQEluPDOEOLGpi3mcsBBemNbd/11FY9gAtWT454e+Ae9krZ
GySdA/zkDsVVYu5EMiejt7PrpZkX16ogeCKwSALghVe52oXfQjUB+wnBtZgttQn8/T9H/qi7d85j
IFjJGHd9LXSmcazlY2g+5SGaUZDsSn+zRTmJkVoNCNZYsBG4w8xAa0pgp/mC/WASv08Ud+guNLoD
EbFihyHUUSMiFWYobGxmVUEmWfJ96HhMjo9ADhjBEpFBP5xpQViupCrLJ2q1TKgfpKGWBiN8gIzy
stdCRNzJ4s0s2jqxZ0hiG4UgXjzp+53MjQH/kPH/FCK+qTz1pAysvYEw64hT4e9bOmoFmUXkgwOT
n8O/bfSXBfMdWH1Q62LfAVmyaLYNjy8M+xgdXQF7Yg7CvRtwf/csKGmBGJ7JpJGgXbO+HAgXzu7T
OpQ5oJX9bKtQOSg7tkWh2ykuNfY/NWJLyLJ3snvyc5rI40f6SDnA+xSM6RGujv62baHd6FfRjG4u
KV9606hDvFMLcgihFqZOGJ/DyrZDj1b54H7jO5cEQQGFMcqeyCNHvLK5Ot7MN9pYbR6lFZK77xji
dEuPlSK75umC70/wcSWR71jxELhZGIaaSShXCGjRu9hawfQZ83ZnLjHem0yqhxplU9PQ/fCvxE7m
4Fs+Dlz55wfhPsWuqo8d/IHuhecTvDUj4xBMe0MWveV/kcgw8tRG1SFRm5J7PqDOD+r9Xo+oAxO9
4/bw3G75MVymRXqmV4UUIhH47uMofIIx9qjwrLMt+rmJo0PsRjH6QG/lsCFvuj7RE8BmJalzTaPN
War2jgNNVGMpj5J+dq4lHIhaY6sk97dncxd8g0UiHnrON37fF8XR9yVgXFH2AOw64ZMsZ+OhdXqm
RioMK6PLzej8pYyse70ghzCV8Psb/1fZrV3UpnLTmsdbHeFPCAb+CnOrr/t/U+LrxIcJkOLcH3sU
oiM9Z5adD0aueS3PpfOD4q0/tb19PFF/G5AoVSgusviXW6C9fKa4nqliVHF+L00OdQAIcUkvTz9X
o8ozxGgaCbjBWbyBhVNC8AUG5+JsHwp0BbXeOPyVwzNO/MSWI/ha2ZM7xdOyDUHD700DoMia3JVe
A5ttIvulHZovylt+yf5CC8jXgBKf23cGRu/otFKSwumPu92J+HDzkuDMy118EwgM079kt7MdfNiN
t1nyb4OAKCEvNyKdfS8W2tTsMP6Wh1nc3bg3xJPuLz7ys9Hy1A20BT8tri5a+HQHdiBWnU+OvDSw
K5SYDAFyHY5Y2grooCnlGUiSTi2Ejgdxv1SYVbyMqfTLY2Y3O9Pi+K/S9eF703byBzFpqKL2enp/
8REECI3FqBOCZdoHwTEDxIN4vIEDJ2ppzd51Y1WLPecBpnahLBfoOXDeaFGX1u9EfeKvCIR9f7UU
ZFfAv6WpYeJZpsBDBYQhS5gJxtUWir/U4TUO4hB4Zb86OjRfrwIAasLUyC+pp9C2SrAMb6uokcYt
EaJRGoRtMMjqc0SUgptOANv5YcpbzYjI0CQZzhLZPO6LHy0R92g3JQJixoDmkyFbNgey0e2H2Yf1
CR1HAJxGkSBQzFHf2QdSWEhDT8u+nwD04U3KQk3r71zacpsKl7kOJGckveS2012oMi+mdVxTJMkl
qXSj0VuDsAwFz0a80gUgHigtCb5Yx4ZYiXG+QF/EVEAdInzNq4ty2yb6jHjp62zzaUWU8za6xSDy
eZjDdcGjxs58mKcttSHAlm5HLSiwcOQU2ZC990+4Lorf5f80WnMcqAlTB0Q1jNispRwNSPdvd99r
53H5YgrUenwqrjzWAf6mT4mGqKsrMGtWvQ98rrzpN95EAeHJoubcthPpkuKi6CznjFu0Ejh0Z2Ph
Dy7C0XgH9WdmNw3S+UmxcCWAfBXZgTEz0G0qbwXpMpigF/LSgPku5Ztm36G/4tgOeSUsJy4TUBy2
/1tYk/ARloisDhm8e2wsB+VkjSA91mR3v4mXdelfSxLOWvleSUaK6G7+RnaPBZlpOTSTFi40cpUN
P4/f3k6JtVeW6+XLSZiTyz/riQ8PfYRbbl53C30QENdGkf3pXqmLu5XN8wKBUMfg5Sy8wxuVkcc0
5LOXuc8QiDi2goLSbcw9r3rNS1LQgHjeJQp0XPsczkCarBQ86si1b5eGZubB8iFhDg6b7mTKigSP
d6lzCIDHlY3xeobvj0GxazIxWkCCozelaZgOteLNqD+jN8AhilB+H1YgjDRde0FJDViGJGSEqqy6
gCZmZQFFFHycigZaWugxXcNsQlhju13B/0UrFITEHp85Qum73lISGX2yqQFlVwEkq076o8xa0JoO
J8Sbe3V1iMKVfHU9Nh0dn81dyYjjwBD7rYRBIOqgwu54u4uYV10+fLAjC5ghLz9SdPtUohYjKyLo
GMtSjIoRl/j2Urv7NwzJPVA9PpOaumHyEwcKN+PjY3MGLnxD1emGybJTImpU43o0vKCwQosK5ggP
iKOeF59siwODe7zk/6zq/Z20B94NXj/x2/HRnCDJAcLEOKJcX/IP7rua3eEIb2i+dEEFk743wR+z
NzRpxK43URg4nFNpcacUbL7EBekmfcg/rKs727GSH5ox8BD3FkhX21OnO/Y0bGQkQkKsZRvtnQNI
ACZYZwMQSRSfdAVX5j0RyI2j+dxi+NtErT9XLaaW3/x39ztncGVmnyNghFVsuHr9RX0YvBUYRQgw
SybTZsQXVAmAnAS2tzff04m++TjEy2Y8tT1lHa3Ea0VpYLOuzm3YPT61CpVcu7B0szQeWaFO3aBR
T+vV1QbyybQ9DVNI6jyhy5KirS88lbxOyhcvheNEnibZOWDHoiHfRsR5L72/qMPhTyANKACQ+jeN
O04VTYCWqKqgEGfV83ib199eYgr9sZsxYcpSskVZrABY5ZYjUIWHdkASh9Rn1UC9THRqPX9knAIQ
qa4P+kbOmVOzG28LrSwfwYR8CsMEzTkem8/Z9z5KhwDUsJjfzigzLReh6VEAV05jsmTBWy/sfP7p
YWw+7D7tAIqlzCvgm7CCzRwLN17AiI4km4TBGU6YB3HUI2cphuZCjI1ZVZOuhHhNt9rtPpaK8UfU
z/9vIuh2ECUHbMl9N71tz3SVPwcOjbN/kYc8uABsXl3+iLf5bsRJHuRvqsGXVHOVxp4aPf3/uFxd
PPaiJXJS1axzjfcI9u199uHA3ewEwiRh1Vfti2NtFnOUiSvDuVmIJMsKykQ8VNBCH7WrGtGhdnw3
aFca02A6Acywwd3AmwaRizG85NSs8GMlw4lG0IN6UcRpmA7MgMxv1cPduA6+8GwoEfKOtaSNOkFE
BpSUrraA+67YJmlpEJshOGc6rfB4P9LX2YcKZ+ofknhhtQ2XSZnhu04smqpUkY1qEn5wOnCPSNyb
0UuyPgMS6szKivWbKYCpzIJ+NSdiAxPlMQcqJ3Mr5FnASNSLyNGC5/Bbnyva3uHK/+ITEpKE4aM5
9uDHXHnxShXRqRe22wkK/SuPI5cgCDPp28PRflWkloGC7y1EjJeWFZMa2gV8dF6oXkCIBdUTMee/
/mtc3B54iTRneZ7ZUgLCB568pCS6qnprIoL+H0TKuRwIy06PZDmK7r2XFXBQoRiR0NAxQcGHQRH0
GzQ3P8K4aOR4DWPgPk4AUM9fTNE3qgHDpXlPIBz6LLnEmBF3pMBYkVUB4zDkuwZFTwpEd8ZmC9mp
CrUcbBmYjVV7iPPN9x4Xv7wSWWXy/ncJ7MnHHmZ7RertxGz+lqPBLrMb8UdGvjfuLLWMVu2P/wph
j9z4yi4R4xSKSWnjaioyXnD/Y9HvmsbRcQef8diCaHsUZtNoudUkRJH1wKcxK3BEKmgDCswgDbUD
MjT4JP5fFP052w2AjDNr2cRDalgbYa0x3oWznqpCPMdcml4UylCkaBy8955RnpJvmdSL9gx62nUT
wfXEvz09eqWJblCrI8oiAhzzBKVub4rYCLJ4aJzsiKdY4pIFo1xO075zbvDBuVDY9rJ0y3/coD27
9sshR7mJ5ZeSj9cMh8djBboM2ITfCB7w3N96vHBJDXy56dWivCIW2u4IMNPrqR114kVIkA/OpEjT
qg1QkTz7P0NGBH7uuySYVR5WcBmATf6HgSllPTodeLjm8U8WTnlv1B4yU4/rNX97EP8x6LyiTyLy
Lg9vkd80iw73dv6hAtGCzKDiBYTGs8bPQgzssoPqeP29QZi+y5UJl3wk7a7rjTzjpW3TI8a2yXWW
4jRdH8j0zPqC2SMbJP+X0pOR2nv2GtQYcyD9XMkASOggRtujRQpayMGYIUD8ihbFj6RDx7CB8LIZ
6VWP8um+oJ1j/f7MdHxL+46LYPIJSR6JSwoWSRNTnXcWpn94yvjhYsLh/AmbIr8WwMPBwoHTPf+J
ihftIaNFuIvVhJDngTAw6YRBxEPz1A3IxfiahQoug8TRUAqStE+f/AJFNfpdxHrvLfWtzNY34LVt
ogg+sJ4I3zB1FL3RDk9koCjLVYGPKMmJqD4w4qlLCRaFgQSEO+PUvH3L1w69c5hp5M5H1ISIC0tB
UtZubf2W/auw4zYG9klHnkqMKQqZkfFUsQMumFk4lWuFDVZWrcxnCwz5/IaBEN32uoATIyQTXNYB
jqX8nfQOJy3GBrU=
`protect end_protected

