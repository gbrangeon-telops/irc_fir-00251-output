

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
e2VQd/JkHeEe4mr54dnWM16g2399v0mhU+1ZT8oWFJUJCdyMu4+q7oH8u3QZmAK8Rcnxp+2SrcpO
m9pYEpjU5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e4k3IaAaNAlNFkvmIoO4qJK1gZoF/VExyr/L2EnpV2zV6AVGzYp83eEX/q7O167vsBLgWYGwRFsP
yi4sfYl5lIuJf2EmeuOEauZwESJuKd6uc1klxaADn7CdEBB8W/rBSaqjDoVCuWxTpK1As0yCX9BZ
RkI2Kfe6mL0Xs6sQpTo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IbtPpkhRONJmgAFUIssZ5lSlLGn92JCOk3a/5TU0b+nZGM9b2fJWwwoGbY/OL/gG3eCzPWC2mZ4Q
yQHVXagA0da67WaW3vnZMDAL5frakXXSrA2s87T1FAjqJLmQF7Unh7546PBsqL3OQpKa5tE2Qt9p
EVAvDXDTdLcKhvmEciakrtXwSTthowcA9uRLxUPk8f0EUO4CTfkvluf6ycg5PO6pxfumZFj/0WGs
vgTtbHeVNSCwdx/DPIPQrx/2AfRxSZujtPeD86jE5AaqkaHPmVodviYONlhtWin/aHIYEIBELmjP
OfgBpo4y7pdG2K9gwF+I76hLDXYgXkS1E3SJtA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jYNHOo/XTSvo0oBfqkgIM6041mVNycidzkShFA7DjL3O3k+3PIOaz1gxN4XAJeVyBTFZGUu9UNpb
lLYIK0sXIcMhzqD/csYXqYD72yk+XSADEYXGdJxFpJfGamCnDtSyBZIo7PBWUINe2Do8h7OVRMiK
aS7bCOSSci8hvDiZE80=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZHkoK3izETxxNJyR8GdmtFOEPHd8+4rIb//gPmmS/L1BfMiycMWs4JZ0IF56rYeBFqrbQeNtD9Va
BKnGrhYVPTrxcjX5+asuKlu46CBX/iIHEmzrKpr/LAUFIgJgUQFePcXNFNPZEAJsYZmhuSrzc2sY
05sJlmShgR0KVQTbBUWl7mt1DY93aBIhdhmiaHpULcmSxpAU6go9uAbU3jUM00ZMhYA25YYv6AEb
gg84k1+xXW4rmxbK8BWXOVrPImvNZoYgt8qi2fdGpgMvgaoBCq3Rxxbaiti+CXpWZdQ5NbjWArUp
y47h8RokwLA8qG0K8OF44wzHSSkCcalfq4pG0w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26336)
`protect data_block
9GQtJruIPdnk3dtCQBDUpj46CgKR869rdFok9j0i4XezkcjUydLbBTrWEdUeSEF3rmWXYLghvBRO
aClqtdk95MyCJhYR+7bX0DhAASQwJPAaT+6MUo5H1d0H7EBFHjulPgezX8cix0U4jj9JgZvBeUnd
lJ7FpPw3V9LlIniDO9BHlsNyvtgVYXPHRbdpQJ6qQiIqg3QsQZJDZlzg1HqPOJdk5PBaGeS+nMIe
dvFICpub88aSmCtgTSh5LbGy0AxgmJS1vV9j5ioy3mtT+xY1YX0QfvcbFNpJkJiAa7/hNkdENZbg
Y3/jEgs0mVTnxtScbHmqYGVPwGyWADfSJUQgqfH+bu88fKV1TX7VUUzTwiEiZDgvhubWW1WdjMvM
kv9pYNiAm4xAoKF0wkOehntGC4CHggUHzQ0oeictOhZ8GLA/y/kKqPLJyMT0WLCD5N/MeNxSZuB0
uopLXyNHjqKLmBEWxCTVc84073urcZ2Jo4RU0UH2KqDjb3R4COmbfpuo/eli4pJGhoCpcoWmULFO
o5uP+sllxUm6HDVC+X0+3Pi1jlbJ/f4/qdcj+I79U0JJCR+Lb8Xroy41uWnAAZlvwGH2CjG0KZLX
AdFn0U8rQCGA7YWGMAlxXKvhUOHe8W5RwTzJNFaMwuh4uzolkL5wOWKqLdOjTlu/2TARk8Kdkk05
wy+cI7LQ2vWOLVznIYVNeKrnPlNC0fKpSi1MZeb5P9V1XHBjR4xxcke662YKqddgsG785C5eed1u
VKCze2SKft0u4+9+9R76u4gJyH6kqCk63sqva138jUxVHJVLw/DWahvgMnBstKloESMi5IC7ve6F
Bdig05PV7eABIkGyJJ4/v6/ATkYaXJz1LrzbMFIZInyKJrZMVzWWCEoFoRCMsDyLqn05X1xZMqOx
VvRhmIXaoWDBSuJFvzp6EA1XzzaEq0ivkRE2pnZB6XunISbl0t/fnQ/y6pADp4X9D8ZLfoEwoE9l
CA4D+fUtSEOg6Zh1XOUYQb3SlA6MYc+jLNbPIEkxY5W6+zXqB7hTG6MdNOaWlv0nFyaRP/vihg3i
3GxQJqt67Sj804e+NtM97HyMjtgmEgb3Q/j3STTUqO4VRicb7W5fxfo8yuJrF+VZHTtxLRA/ZmUB
/hiR4iWkSYNwGRTa5YcfRjUUoPrlBnmjLzCCAPlWEpTGo8Zndo5X7XoDXY5ohisg7jFTzKY+UcI6
Kv0Ikj6S0F0ja9VIzPuPBYRKLwBLWHskt3/WSqJc7ne9Be8VZoFug0PNzGvu2SIgme3AkWPzfHjb
4XgYGtRAaB1d3Mz2BdFw6U/BtwHxWu5pan8kP3tT2OtUXbrxW0p7l+A9tG2F/guCmyxPrncMt3+R
2n5AuJ5gqLSHugpgAWC7rW0Yab0+Yn1zfE4Xc7953HjQd+iSZT00HKmxZxai1ae2xRUYAc3QO8GN
LLk48H8Lq5Y1BM1T4yiADuYlXT/NKWFegQZ4fSlnyNI8PVa0/N/Y9IcX2J1+vA0gzlQ9Nu+CUQjS
3HhzAo25e9JqlteiI1/PBmWNxETOpi5WljE5V9IUteIruCYGScvoroETpJvEum17w5DeYRtdMIxy
vX4rDuH8YrCyvKR92QTGkqOEqr16csh1ePVBekl0coG3ifzcgIRqs3R5JFZh5923K1hkSMq6WeOl
qc6jRlws5GF1DJ3IFBSELbdD3iFdeJWTa655ktcuVT5PKnQaZnLqQ2d8hpOi6QrvATa078B2K2UD
fUHk3ctUx0maYyIIrlxOvidnV6uKZcWnZb/xWXoVj8r3Xz6cFQWjLM0hUti4bhS1M2lwODydOWjE
alyaj0JSI37HohGqUGgwrT21Ok3nrv1rn7evmciiQxBOKMtS7Ndi3rzCJYejCihqA4Y7+OSHoHz3
HQOFG0AlAiRhVtRNEtEpqHDetD1+1IUlcDna+fJbd9F2SDA2U+IMuYH8WoY5eHsM0JfNFYVCWhwh
7CS8uxAKKHoLwEwLKlEtaGGjEmMpwIrqd8oYhtObMmNrhhcfejopY/Ndv+2NOCmfWcdIRD9C93tn
b9AMLeAS49YMnTV19Ba7YuPYxKfJCDmQNGUCdXRnECMuVbF6FJgO06egfjLB0L9fl+3Zu+eSV5a1
625VqbgHlZx6vjDJv8pi0Q0y0WqFIJhRr4aZu9XzDfbg/10DQKXyusN1n24ORqgeAmTvOeouUxQY
m+nqjjPhau+oFW6xvYAhYcQm5piHKXbvavUtjW0nADgyUmS0/Rr01lP4J/pbxScyMnCYtWu6nYeU
tcOO0vKuCyWv6MZyfy1ix/EhxpXKwWAFeUGu3BJjbHhb5yOUFYGdMpsZHP6WcTU6ftQaegh48YDK
krPgDjjpPF6fluTEu7AAdYEK5O6gOQg2b8hvKG+thm2dsSbzJPvamxA8roIbx/+TYsx3rmCP+oQB
Cnj8va6tswJ90g+3vBT3bCBb20yLVxQOrqsRkpYYeXlwVQO37w3NWuiAlZAeuZkg03qraWPSX+xu
XUHjXz85887+TMglYYHzsu9c5vzd6aPOtpsZfZEhPahLgdnJP29JDskoOOgj8rNFv2fPmJqrio2p
hyiHJUQ9gKVRkjsBL4WvXSBdJTz3VVg//Q51UmxEA8YxN8YUGQW9stxUP11AVJ2LPwODz0pGbF/f
xDJUFL9OzZ3TCeEhzfjzcYMswKrKjb1CtoPDeSZbk73ZbPMr/aaJELNoi3iICT6LPWoiZ2YmqJbx
3JnWjVIGq0iX2WO0ktSoZDp9N2q3g46Nt+6ToSVf+Ynx3e1k/Z+Ldb/LWqgg5gQvokpkGYw4IwwX
wYQXxwdcdsFaW36p2Gkfq5O0ngmzq9tC5t8jO4mY3sKlhghrLRLUYgg5wphUU12UvzsrBBoG8Mdy
2GZAMyNPMkboqveWScm9n5RCOhhxsmLoCbjfqweallkFnXrCGVG2Pg6D3s5/1BgY53T3kZxJjcTQ
PaC6miqunmyYVGNw5cIgUXftoSxpvHgXmwZEx4h3YrGWTEZSqtgZ5beNysFOjIH3TONa51uYwJXZ
j06BdKZyVi6KHEUFnMk/LXqaPbQvHyc02IhXqJM+NjvGuW3LiU1+bIWc56N1LQRwcSHCESpoFd7t
xcaXcny+bR0Jobhz2qsxT94Pt8qbXHOvQGgKhMmv+gtNYiZ2w0WnBKV0stURZvaU+qri9NNYX4rs
SaKHSWWmOKE5kQ0EbOAVWQ32Qf8VcXa5ZetTjeoG6n+3Y3AmZ1BtFD6vhEPNsbMHTEQpT+eRH+7A
bGybLYdh/GDNelXGNQ08OU82JahuoG9C/dNnDFFq9Yjy3dSgK2qMrHdvjULu3vNh8icm7L4YITCJ
KvF2uNBtjSiB51m2o1GmDSgAlfocMKgDXgeILiVN1utMFReKUVZGNTGp8KakyXTK1mkFt7Yz9z3Z
GVbNsf5ZtlQd94z5Bm5g7e5EsRI2GrkF6/IJqB1v7g6QTM1W1Lt0sP72mQprnx56b2+j9AhmHygx
269k7m3Cu1sfkBb20z1WSZg+iJDkazXtg7gU2y3kT0YkQHcUkVNzLl6fduUAhl06uPcAr+zkBHtu
bMiAZ1wxGj2xjm708w28ACnpG2+ewUJBlgSW5LB6UqSpzHQ09F0LRYmhgfPQfuWKck1OH/Imj3q5
l0xAl6VWj8PSn57gY+MeWzEYKGYOHqvti24nnINyMFrzyAtvALw2YJLBXUocZwSFp9Ok8kONRKYi
Z9kEp7hmtBMMLdGabI7u4Duq1ZJ0BVLhdbzQLPicDeC53AwHpHqGGxN0uaWXQxKheclpmiCXkRcv
sOGdXG+Hpvfrrupf1//vx/Qldex/oMnZ4kiKBcHrjmOHtOeKdkkhUFVIr5/UyovgfYIN6w1o8Ha4
JBQavUeky/2gbKE9ati9mNjwGYOVV+Nc6xujoNUGLtlxV6gWWHd/xz+Zl+k/VbQIyEZY5tWHdAMd
RdI1cvZ6CHYNirxdFGFOBkQiq9hK9UyjRGkafldl/knObly5qgusXh7Q6xnNLvMRX5pVnG/hNN4n
XDWujJS0belD7OoVJWk5zNj8hP+5S4NL3qhHIyZRCzwsUfep+/1zJHpwtK7c/cGp1lxRL5nnTy9Z
Zoe1FB3SnazhIVeI3UF25+ODprEl8q5i1ScGCRU4AkTH7Poo8aFC4nE5oVd/FrKU6x5G3K37lmak
DkYGRQeWAPj7jesUpxYpHeHx0JKAok683aLr8gt1WUFvCHts882iXeWPN4eshm1dr//priyh2wto
BKUM53AZu215O9Cdt8ofi/BeIhOh6v2jW55MAzZW9efAA47lT52PBxNtg1MKpagij5yVe51gwlU/
DAXxB4uyzDMA2AjBdAkiGBnk0WGKQkHgdHwCxLJs3EtcJRdl7iTl9vPxDLr2cZ9DRVX+woey677B
96jtIV3Sy2L3SxzfunvtvEQX09kczGYQ/fFIL2OuSLkaxs6oGwhNb6OsAV8+uSdA9TgVGDTnMw77
9C2yhB9eT4lN9sVvBaFD6mcZ1cpNilhoz29Fv48G0fNq6DCXbZ4BpDiVfc9s+EG05o/yOgHq5g/O
2wk3MPgb9asm3e3wbU+bROB2BDyyKHsmdLYHjh+idNyRpOsG2fhclPFbBZvOOPG27uXd3+aJxYmb
GhMVzAFQbd4m0z/bLVbhZKqNh+A0sTUzzOuVSc4k96HoUUUB5obIUsqgz9vN8TOfKx2EmqeAEx+s
WsM7XLB27jLCLOHdeXpf022wte+WKcSUdy27yq6rDIDz9Hr9MVBngmZCdRewNLIhxkO5Igr76vn7
t83qJII/vgc9TVACHjGakuInfKKWDeN+IGB1X/IoR6418IkP/LKIeux8UAG3VOY0QVNu1FkWpxQo
cRUymPy4I4rLpSEFbrh2igeVeo3ghNmoSz775s53iXh44nKpOETc/KVWoPJQ/+vYreOa8S6LSIuh
KAqFUdKEdWmJeyKD2CUFgdXMLdQ+qRWO5kbI6XKW2r5NiBX38Pmhkq0+SkI4F5TIuHQ2Wmo6uKTd
Wg9sJ/fSWgtmRy4JSwMe+F1TlkuCQG/U7Lvc5cQ2n2ffN0x+pai8LOvtfm0hXSbH9/GgWvYztez+
R+9uMX8iLAPtna75/6S2xxLVQCxQNY5wqYXzzyJIRrkK5b3usaRd6NKSnD3GndYeLWLunqGDTjaR
YISy4vvZUhT/fjjbH6Afdv6grIXmRlUkqMSd3a32uCm9W5nQylp/3nBkizP6UshFiKQTvRUaBOZQ
hRrESjveoifSFAaMWFegj0enElUS3ZWguIQo0h3q4f1scceDt6ZXMOzZfW96QMNdvkGkPE0V20jq
NztzroTo+mwxQv0Fp3xBl1K6lRUg9tMTzyAzDPZMp80MN1pj4gDKA13EI53iMKdd8bRS74X2o8J1
e/3ceOmD33gZp4JMp5UTXSOciZ5+yPI8oVoM/zYUKUFPFBPPMo6QYEs1MbeBiwZYBeB3CBPiFHij
ZfvuNPwYLODrmBshf0jEFeiIn8a6a6u0rWiqEug0+M07uLOQDYp+r1iAIKYYksAbDsgJWPRysmjr
9mC8Xo4yqUaNtztjlVNIjRnLEw7xjHAFmP/hCq788ego7jZ4OataoRqoF9s4Hkz+XqjdOiqcimai
W8gec1/XuxTCKucgKqVh4/HfhDzxOKJakfbkEDwLnTPPgJsXKjcFCLYZEqZvwE3y14oj6JFheIJQ
A5st7oQtoUAG3/biGge07qrZXS440I9U1tLtXTzPnXmWQ1MqVQ13kjgBDNAExBuVuvlRCN3sQl/Y
wCR3mh2P6eekAIpyXujYFCesAe0Blx9HFVhVOKkCtbP3SQkFFzwFyKpC29vTTwl2zAAAo3Pz5pkO
MO/XzwsV5wxKmzmV+oor78WScCeBxTjQTMDtNtprrxNtWDZ1HZKrWyzUWkEx0REcHtWZKzNlhaV7
PRvb347nsmIQXW2z24Y+gUx3gDj8810oRylYimrW27yd+XtnuCvRP52OeGuBiz4AdAyv6umJ5mw2
Lr5meN6dyZV2I904plNp/eQcV9InV9TkfzN9Ftg0ggrxEQC9n5XbHgXGVOXGFM+8uz5DofW1AXao
8JUnFdoUax3dbM2AOTQdBPXWFDmgMiQ+NbZYRm8ewZFvA+j1Yg7lqPObhywk2a1+zQRnwxROrkt0
PzpqVJsjQbn9xfqoBEcYt7a/Uv5yKYGkAeZiULNZrin7tP9uuk41QNku5DFqTqPOAeTNwNGO57fp
Tt6dWigrB7xfSM0MyW5beWfnufggqko/rjhPFGltS62pm9TtNkx2pgD04sV2cPTMpfSZVuTW8ybX
N7ajYIfcuYLvNmxUeZLPZGMEVY4IXLU+sFUc1pDKzO80KQR1aNDeccWvU9ZHoMuYiAbXAu2pYPWM
9GDZhEct5z3EgRK6UDuwu7ZVtFh9RQtcawHZzgqHtMBl6HRb7WillWZDXKSEEqDtmrIK12W+Xt7A
PkC8BaT/NGbAuMws0cJVvQuvAibtut7XWKvrhZPX/QiSnjDNeVCh2QDcxH7tJZsMUTnNCuOoYGl0
jHhack+2qh/Y8dh14Mi2inQTpvlWdsLVrXxJFprE0DHCEAwxkiZE+vJuijm91zzBt0F90OqWl84r
MlGz0j1GxtAjxOw4LGmZaWCgb76CvSSpVxwYRk8dB/Zwh8SO88AHS2nI9OEw1b+zvONHm6QUXunW
i+7N1LZrbRcav0st4Be3AJ8Xhh1CNnvTV3nIoByNDE3LgUx8wOsWcta9CINJ6Msb9134VGOg89Tq
SMlljQDnIrIVRJjhzGz75aY5N2vQXvUbq3T/N6ljk8yjiaxIeBoUoa9vGGSduVLOWCYBOP0ZBCn0
HNXv9uutW7jVJqZZoovQeCEaHaMkPTnwBwaHredsU1f2Pg14y37c7OQKOUh+8O9qzulxNwLwpg+t
uz628CUQqzyEwTLx0QWXE8UAz/8Jwl12hLQu39prhQVxWb5cpeHWTIflzpVBohfa86dSzKZ9edkP
XqnVfKeGgtQ/o7MQSEwS8eAfG29TVfWe2aqp8xJOVQYZNikpAvWeq6DpMJ/fOrzNWbwS4f+vY2R1
nLsjH7PlH/jEQh+y0QkrCKbh75YaNpwZUwReJX1dTdWrONXnBGxh5X2YZA8dCudXGvSo8yNh/I8a
4hmtJkbw2oUSIqBiuKqQT1vsRnpdqZolFVpeXfw4dOE70duxDxXYkTkOommk8LcfVOefHZtjMDnG
cdHTKQgq4dBlP+nsx5rH5RvZN5w76t317E/1Nni5SZgy0CseSDSnNkCszno0DJBbl3X24CUqXfRi
HoNaK1TOpjZIUCwnX1tSRuTnWls9zLW6nljhjOoW9ceAfqy/216udkogmOy3pNRv4sDsrNW9Qddg
bPpq9PlgmgTjYjWvwnSNJYKm2jkPtjjWahooLSZmz5EYVCB0iDEMWG2yugNwyFwTS9KG/bbAdQZB
R/U5NrUoKRVKWMH+1iZA6gRn7E76iaLFZHjdgn9C+3TNY107kN34XuPfhMxda4iyJqMm0zBlgqxv
rKk8HKs6Xx2oa6hKLQGa8/PhV+mI+W/NI5ULDEYwjRGyObGDIG7rOmLUAfGkYNxSQJM+Uk29EfDL
MurbeaE/vFktyyu/xGLHTZIiGjHjK+ZHZMmqPgs4EvSzEvGwqAoET0ES1Kzte05L7Y3/el6NzKP8
jExJ8D7Iq4Bhmj/C8CGrQL0oxKwdXsmIRPrYdvG/XR07R7e6NzB16h/fIch1IPnVWi8O5LA8xqeB
0jF+7sb/ih/XFdF5jiV1Ev5kRcDE0x0iq81PONh0020MUdyciSQiJMIqNumK+3nymjmZkAsBi2WO
bddoPJWFW1mqeHtseoS4+zjk7ul6b5neH0iZPiawqPBH+VZAlZ0T3qJRIkDPVGNT7bb7kihPgM9o
GzV2HGKQZbKew7zuovJFF5KvG4ozPOegxeF+KoXIAhJLBhsMCpWjktIuwEXUWzDADmwwYvR1IvIt
a29SLhXRlDgmEAU8GnGVN7ZB0jnQuy8ifEKl3PrDHK0crkzgIaZud+o9mhw4eUVajXvJL2l4ian2
ec+3NY7RPp2NdR+PSYrWy8UIkxeZeT2/uqjYSJAmcSpgirY1SPmQi7o3Zl6dP2oQ+iDKPnCVtESy
y8aS12UDThtR8cxQfInZ3zBLgJsWrsdkkm4r1BaERANTDOWKA/IX/RzrZhXtiWcqC1mlsy7LkCab
XNXBPK/uDskrhuzR9U50PNg2bHmNVikD6pZuGeoAElN5FcjDfZHN4NoGSN6VL/bvY7DVTqvHhIxV
tFONzLDrkD1pC8vBMV7eei2y+BppNoaFac06r0uQYdJV2PR2jexVDw1ahWA7GdyH1BYHZB2mCp45
pPtx919QlzahDMuKvHU9rsQm1mW9uH+LO/kQwdqQLEtGQqKMtlegzuo8u5Kd0j6bcgZ8PLIR7sIr
Sv1RwDof2axRC8bNnJZCrJdzhP26QJHsgpwJEsEb5Ra5ZhDH6q2wnek9o9kpI0NASNsdSC8HyPY3
VnzOSyDVCk5h/ZFQyZTdHFUTKs7AFqDrLYD5/fMW10q//9P4/ap8LLdWYqpmnUhNmojXUu1ORurf
YNgwbK/CD6w0Gxq30Aaj7dgYlWNHAd00XGHGz67Rqe3ftDH6qVeAaEI030Lm3z9BWjN3eMZKksEC
SZBHzgEwEW6c2uXUzvTidy7swJYb6vF0OdJv7ujkiVAn9rjIabBo6EaB1Je7S+H0QiS2QPSTH/Oq
4aVEEm5LC2ObXgQ7qvxKBe/ci2PCpOXBPCzC2V5oladvTfkSLdFBUl0/ltl5vz5Daqx4aaIsp4MB
KROxXfwcryDtZRXn/HmWxsfg1IDUUw3HTRQIb2irwz4UsIlQ4uCBqOXaFf2mjdBE4O/rZWKB0Agu
5dQlV/v6DCoBcw9otGdR0uVpln5eLe2pG/oEXI+Len1t4y2r4h9w0SkBu+ASH3UknZm01PG9a8iM
/Erhrz5bOVoOgX3SIAw92JXsNwbIaU+UNQKcOon048iMNKzU/GODbXLh2VfbdAJ4NDk/d7RRMGtt
5xVZywVvEfIDq/WWcFhPKxel5xbzKUCcyCBYwHQIrZZMF7PItrBtvobgGqEK8RlavXTQ4dNdb+5R
43eXTFSxCXpkbe6PbS9TbBKf2BKMpev4kEM2MkcBUOb++SqTMo9RLRnnMUMfLjO0ARPwblGoMwtf
ETQvXhAZFcv1NjeVzuVpRUke5syyOLu6zRoMnorJ9+yYP16v0oy9MbN8awthO1jx6WsZaqclsdjj
Ib1N5gmAnUu+LBfKn2AvPoH+Dw3cXLXkJHT37m0e0yO+P9FqWbEkFv5QZvia5fY0Puvn35xrhSA0
uiXqMKGvqFzIktq3sVpOIGpm59oIJ528eLxC5FqaEfx/phK19o3BT+LoqBA+aYzx3qgZqKhYfOnx
0YIYetOfI9Y13LVm+bwHw0G3CWMO0nas+xeCJVZfDL/OIWdboEyX3CUNxJuC7WyEfE5iS7vnar+R
LiB0xCjN+GVEHta8YSZ85+c5RIvGhhBXthXbktbZefzvWkGLlHLcHw4mGbPpjuOOyK91rXI4iuVr
yNWO4hp2Zzwz50wt6Oy5VWXYpyCaNgy86SM1B6pgutMdKGgsIkKwlG2trCv+qCzOEm4Y3qDC96wx
RNEDEdiXZEwcktDeGD8meq8YPrHmnQylMJNT2OkY96P8WXMkxTxEJNSBlB1vXncdBJSRZzd3j2TZ
zWFHo3m3zRdwQ9hNHLT4fwSjMLe8kuynyTvkyPJ+aBfdGaH7ggG7mfJRWi9IISYyOQLEVRTPcfUh
+7JNthEDZdDCNBLkrADP91eW1KThqmENhJECDaLUrtkKjdKtDe6kf4dcMjRjjr01t1LwH5GI2TeE
sWfZB/xRxJN+eI2FAE54QYpBQQ6WsREfAtiFSSXIsewlvZVUOLB9G8KKjc6Gke3vLavaEXMv2rbp
YRYorwrqkU9UOL/H6AXmOqUteix3Le2exgnMBTBZc5ytbNMPqlJTPhzgLwQxuJxy6GprcjZXT71B
WQjhBcgsyiy1bPtD2CKdhQ+M5pUwnEd+ibh0xRVy3/joU4RIk2a7U7Rns3r/yGFqRev/mswVUpzg
rSi/MBaPM2GYAugcggA5TbDb5Tf0TR0scFlDkJpssz6XFbEa8qk3dDWQB98mkoqZD3d+kvnVrJNC
T0e9jKP3yKH96czwEaKza6Kazvb0WYa1oSk2q8PS21ZFtXgxcbpxQEuOHxUkuT6DvWNMZ2JENziN
FFbgi1+wfdCLNF51BrSlhUzjwcObX9Yxd1oSpgiCgbotGZF4mrV/qTb5Cwc6AsZCjAP5NnfMXzJe
x28dzdmaZQKYGGqikBzl70luATnd16/+VajcjgUlm1+tva5vsDcqxWpse5mQX3RpOnL+dGbznjpj
gnd4lp99brdqc1GstVquqa6BIOb50Fkugy84rKdugH4V2EfYyom7BCAtFUEGqEBW7daBSkLdH060
DOff7amebIZOaPFmqF1PG42Ie0/uPgmZN1Zz7Hehibqt/+zhZToFNEXlElVXO9q8wLE8S0h9I66k
i6R4eeJOIoqxas93GXwBtjwN6QqMB1VK2jFBL19YrDZe8xWGDx9w7BpotGJCUxHeFAxaaIz1RS5a
y8TSFPYgCNoFtBbH2GXkb7nvSzrsKFirNwP+35qqEkuxHWZtb89XOO2bBzwCd2hJUQjqjVdxHjde
tNphfDG4pJy4mLjO7JTGR8GsfDddty98OEXEO4mkV6+dAzKuUXWWQ+Q18K6876vjxuBBd9wyfRwK
mfm6goYs//J5RwPZ5J30Vj4oxjI8xFMm18ybATuO00LI7kJP9BgP330JCQAC2lpC7rbvIGbvUdo8
gruklMJVfS5BxuqJDPSTNq+2E0q9lda/sszhETXEc5YQz++5q3Id1io52FvuQM+Yrjod9HL/KqOB
KKsAgJLGZtM8jskx8mko+d+GzlCiCGVl0nYgRbBXOrfq4UO+yBzrvRhureKfzcqGi65IPp8M4o3S
FRI2mrpgezrR/gf5XouEjAdjMdazUJPaZFcxTolb/+Rn4b8u9BfB2IoU5vFe/mTsxg2t2p5m1MOc
4PvnnQBRdwfPjUY5ODWDM6NHyUEPzWxH3ZAdx4DpD/h9sPbjZ0JEzHLy3vylljwfLqIba9a6jP//
Ht1rrDFZ19j+hj/bNwhpJ6jCfbvlyOkjPz4wccmezgCh47T38ra5NfeYGmar+U255Ep2Gj21/LGT
t5CoTHCV+un3M6wgrEqK9vmiH4QSt1/UPXNuPpc7aVRSCivHb54LXUfke+HO3nQNF+oOKBKdHyvl
z1+zmV6rYeKph0hduLRjDQUtZyM19F5eyQwJDCk6dvs4hUMtoG3L2QSUKhpTQ4b8QOCaMuYqb94T
R3xB0pRu8fpPC35wGJeT7t0FtOpUxSqYXDmN08WmDTK2ffAAPMxxCxb9fEEWZr7It7ZystmSrVQX
pCzo4IBztdd6+uecAF3efMw/2pj7ejl8TMqCpb4Du2HA/FWvfo5HP9qOfA5C3p5YfSopH6ZMvBlQ
6Z/l5VfZpyUlLlIn8r25eaeHEemAn4pPyVXUOuQSXCznNZs2ZlqHEZnmCxycvp0wNj6DdT91HL0X
4nlVak/qq5IklfTV3pg5phCfCZ2vKpc0bR+pguwd50en0t98VmXaDG+WnQ5or4PSLtB4YvdoaA1H
zRpUTJQWSNTRtmzyQxX1Wig3BJpMfullR5uRylqCZiPaX2eILJJWbrp3KkFXCfGdFImHenFBg/FN
NmhH/K8LlIcmJ+n+AecJ92DDf75SDZ+4qZWBfs8bGFksXgd1+3YcOyCFVXJjULCtiBxK8/Efz5V2
qz3Ia7vbJO+TzKYYYkwrMVy92a8KmTqc7ee9aSQBJyldMwItosVLneII9o09TbyTu51A4wQuwmg5
PyL7VeKud/JGCLsDrCd+pNDW/2q9PwLWZHrtrxDjERybClOVwLNRvSgWvd+2WOfLrwF6I8NnoXOX
lKnOvoDtFwhjpQZ/G1GgMEGksmYWH8RlJjCzhi10BP+0qFH57fxRBTV/Kk10FWGcxT2ejbq2k6e9
qWdWO8cWoGyPoqGZ8zkkgW2NZHYvDsJDO1ZIrr0P16IAjJiFJd8ZQL1Khv+J8iw01NZK5PKSoOMa
c2Tw+tC36x5NEdX/Qp+az6Q+0SgjqvTjMbnkEaiSG6DMfCfyLXIs/HSa+XaOGoiHQ4R7vQJEoALF
EfWg4KbLbbHeohYSqLH8wntk0J/RWbaxuGwFsa3kx2Y4WyDGFszaRFt60ew66wp8DSKqFtaDrKe+
HF8pkX2MFT9kUbdXcTnkBSsnNp9skXwPagSm2wf3VBILhCv09c20njIOHoIRcaCAUUMEcCES0JG5
ByaCeXzqf+sTMB0QnFp7n0sR5ZobwHefl5pIdkHKpcdxQmbRN9vZHZfaVFbFpUq1CwZNkeekwrXW
ncTcxaBV/7JvC7rRYbcFxRe7uWJIvLXWoY5khXYVRA8LbopQsTY5MrGnjqeW0nx1g5wZLvVvzmlD
cM4pV+C1VMYhcNI/D2L1KHx3b9/WEAqY8g85wPELiOn+6XgXR6StsgFaCtY7VgKCHbxNum0F+lj4
Ids1Z43jm5Gf4irRJ3FixT8cTc18wU9FUeJpEW5ElyNQFidz9s0lSuvC/r0Z/MvnEBLAsLdITFMj
myScRO1zlUaI98OnPNtGqPRvAWI4lXaHGgup+flQFPy9MsdvmbPoOgFEJPYPUf9eKEGnqX5oP3eU
XyoWvwqtYOtBfoG6OZhIysGDe23iF100Gazpx/pZC0QeU93NtNdUjGs6UM2IYLvASOJI0flyFOH0
wusCto8oaZhYQh1Bduo4ehm9odkJgKDqENS3Sobmi3Htx83TGxtYTDyEZLNhFfEVGGX2ikkDJ9tN
EbrK+Y7H+QbsSkBr1tJti0ThI79VR9BimgR4q/CqpORYq1pNwDqSVr/kTSnrqqDWLS8XowgYOKY5
opryhAbRop5XhlzsJemuHDPpj04XxT8iADPLee1VrWMf6meXfz4OpZltpVRtT5c9Fo12oSsSC2eO
orJAVJf6j9qKQYSJhJuA+hw7WtHAqS1l2bh53aq+Todonae5ZAfEWaaJ0uU0uTQToy9N0wALitH3
QqLMvb1WK0zLnMZe8CdHxWDBzPcVsW/Z23ze9H1Ig0IGvrKr72hw+oQA+b993hMBCbZ4cqVVSs3u
FnmPtEN/fOpKl6J/HVYFAiwnFR+K2j3IeAnr++WBnCi/nyeuWEJ9Y9IT2AD/DSi+5uv+HC/JEd2M
o0UBcEckDMw2Qte3ccBCr5Jm45RZ702GsbB0dIrWh4vupVC6FTgkBcUur50IaGECTreN151Wa77k
4tfazhUQ17m51280yrWj+jOf8wV51nS62uBJomXtmc4rbUzWHEa7SP3wE7BjOPq52w5QyMLl5Bd5
iX1wTXQ44ABMpL0EODpRvY2hwZMI/BA5/hSiWt2cQZFZzlB97mFL1DqU6XAloFFCq8rvqMDhVIOy
OKLM91XsYfp0X1BIPgQ6cBZOv4e99dlwCF8a3sV39AH18tWyqaQ92Qn/sqyUZhB5FYT9YYM0tbP6
wMiMkTVQHiJjdw0BIpYE8o9cCjILBjMCrieSyLPF3Zj/IK0sL4qOvjssE2zgsGpwzYkfuQeFuK3R
0PhbPNlQtItOKyS4ikO4vZO5ufhojm4pro7I5CzRKO9qMr455Xubzk+BPWWnF9+WiYKv9MICLyvJ
ex99zOH7k/R4MU83mwy6yKbafXb1ZYvnyZIOGl0Sb3rpK2QFSY2nTm0LxvTEfdD4qs4RX9qsIko9
RClckdoEqPpuCKeNzyPn55IcGlgGYPhDjGypqtz4jF3HFkzKgyzbFTyZGHSCCzZRJCfGY56xJbdF
JMuAsS0tK73+FMcG3GlIGE0Qdxdaf6oFchlPQMrY7eyfmlyxU2U1jvv5dUIvNpxCBcx6E88XfgEo
eTmmQ07c0r1h7PH/mgQAMsbxYxAZRz9j2NbVkp+bNi04/BE92xGzRWds/pXsgWulAW5ZM0A43Wbi
vzJIKUNzph/w1WJS9lHhQ2oG2Hw3r3+CeP8f5UgZ6209Z3CkBQJTFb8kDSD6/kKwm3T4oHu8FuVX
5wdTsc9zzoPK3eGfEQs9hoolrFWrLHd7xPMpIzo8npROwbk7eCajYkXlnBiLd5yHubfDzoV5UkBf
QHetcTL8DdRjMVuJG0iPwic/gi/maOQBaM3Ytr6fjOTIKb2yXdDTfW+veTCFx8ZUh5RdusePLRiu
YiMRD/vNXxqX+/MwTaUhw+wjx/3+FXA5Db4tPrXAMth5+Y5KYHRz+IteDuiSOVVU3vLa8l3uDZYo
Edo/40U3FytQfRLckJLjDXEpz8nbaEh/OBfKE1CP/T64Z706Tkc/dhjtx5R/N6pLM81BLgPKK1MT
nbUfsruUNSEuuvFAKxFe+rC9XyO1JdzVrzPLWZM7sVHiLLDrGFC+k0+4PwbYdFnEDVT3lpDDhiwQ
d10U8fVZq/FsqiHw8fJTRVpla5agJtallbgywj8terZz0qvgbIq8COxTZBd/j0smVMgl0UOW+0rA
bknI5luvtO/390v44sVHF6QbsghqetwGP0klGTct3S3B4kDiK1k9+ZYoAysm3sWVvHv2FT5TVSOp
buEvMQ7VLRN+OvUDEJMnGSw1vLIk5fd7J6xFtR7ANwU8o58StbRCwZu6zN3HMSWLdpetMmVGlDo2
vwzDEMWXLzEoUZrxmuQc2qSvC0oRZ+QyXEk8htfpQ8Xf1ebvRPWczuwYppzBaCC4OpAtWS9BazQi
lyNx3aveUt6wfkHsKPWd3HpYX21X5T/me84a9o5cIc4sDWmvBMhH3WxDlK2wzpgrYnXwzFzlfuHY
oapF3qc7gYcAsJaYAuSRnMZE+4/41NJB3mwlMBw+vD6YGYg8VlIJ+LiOVdl/0sYDHih1MJ2AR3Tm
cOceZzvPVDECbnJ40Xd2m2eHb5YeJ4KtTInQeIdc/YvOwXKhmOnYit18dh2wFghTrOjAuugatHDg
Y6aSBYMmDk69LMbYZmaxaiLggL5DpdpgRdZDFFiURtrgoTsYOTkzHrlPzqkZgxmRhTW503n4Ugvx
UWxnIfWhf3W85EFFzWSjFfAN+mDChSpsng5idxJ6npd9ySn2Q8vMp4RFHuFNk6YuxxHmRXZ/DFUZ
8TAYmAt7eA8g4hDsou3zCPaL3SOiDRvvEe1BzBQW1KILmCIgOW4f1o6PxB3F2Gbs8l/oxO1HBB2/
rHKHtXP6wQIqZgRgp4uVGeAOmZenQ0yZdH50Mb4QT5j2R9aOxaLznQoiuuq/26N041d52WhIBVjw
v0Vbj+OXZjODtOY53mW2lePA5PdBYe/efsOmRfflt62xU8hujkrRRBSxbMwfWVn9Rqq1ncfujaej
hNex4BuaaFUQSJ4+g/I1gfNJk3nfQmydjrCOKJwd/30JuSOiNyyvvIo4TWmLpeoQz8RpC1tr78LV
kg6hCtTricSSIfU1vfFD7yPDMryUB5zcugShirbbgWHslOAxlL4u4e+MpqPYtNtI9ylHzgXFjV4h
X5a9r0hR7kgm0lwskXPeg2j7Om+Hy6td4oofhUp9Vu2919TgJ89oWQZ2NNgtefdlgeVLlQW9OS1U
j2KhNs3CQnLBfZ/s/IrrN+KdAOMWcOL7WvB1bFhVeATF/fzy1grJFKeMbk/kGnLEQM7HV+t9dole
+yB31/YiZN0YpSbHTYJVGvHE/eZiDj4aG5TmQSELsKBnJKFfGhNems8O4IK68yDDDhV2UqAWRlBW
qGQUYQUkYZQ1uhuMBjiw7KvghVc1QmwadaTGAyauqbm4a7JXmRpagl5j4szKVdYjB2uZf1HEt4iL
n/i71iPbYjPkSefMD/VwfVqfpbmPzxZsiEwq816E2FVKc4NiKW5TL96QYgOwuw/6UmpdMqAIqGLe
ySW9rA0qqI7JJtVZF5YhY1L7I7dK2JYv7UVOY3hKenH8P+LpbofoZbYbwVw9cBpyzbWFebGUyKTu
lvauNrGKHCpsylHGO2eMI71HeUOffYtKCafkbovnfoyf/0DBvFyIoc4Dpu37MoMsc3uHc7LOo/+m
j0qsRDMDW+irxOwKVjxkdnxgBxcEsjT3Ko6otmSEsHLyZ2fsRqA2exWD0r9lk6eaR51m1yLhu3Zw
2nJcEL6YYGQx+gGm24Fq87cDcWHdsG45tA+629BHPkzsR1kxAqWb/9lkLOQ0j/zQB9f/rlEXHTho
y3I0mB1/2eZ/erJIO8/lhiV5ollK0fcV4livnm/kx1Bmepnw2cFLcQk+KDlvWhNcxlQMHUpZH2Fx
Awc2M126WBvqkuMFcxyfjmIs/Wi2AGe18H3de8vOvrsWbBD890XoDkenfTnwWiQnErrhPnq6ajF1
9fNIXQm4ObPUUAzL/de1v/HxaUnT5ZPq0ci5M7t0m5B0EmKZDw6Z/lURMWmglNlJEj86yRq2YyUN
S5E4jawkPd2Mm8d/yPyW0UsebP70TJ5eUcD85j/VP3ypoCdNqaVpT0S4xy8tYoSXUuIuogt4qWGO
zGodl8X3RoDrQ6iuRST92/sNGDDT15LEKXbizEFINCFcngkrms11huqid/Ijd7Ixp0V6FOAbTNtU
dq7EsDkNZwQVacZZgIsvUl8vykZhHNwKTmohfu+XQ2wKYKVRBehuQTmSQbyWJ3jhDqCiHGg70gkG
TRkgdo1DozN7gvI86LaOO53u4Hf4TIVv6j9G0j7HVu6broc3crR3r8h9NQrS1hWQngcJ+nsbvAJA
xzMuMtKOMbFJvyrYR78L+D4myKMXGxhbSg2wa82O9YlqMnLSgyoCpjGXp9AKBi7RgR1HZA+ccH28
IZf4EQu2+IEMT7DTdCJdCyw24/kAWFpP13Cn/jiLMbcTshpuyRf2cf5Q1mvqKi4jq602YCFlzrsU
AnEevEnmGRh2I1GnJmAbXYyE8Pw2hC8FH5dz89IaQaZ95g84VSADVUD7HojZPIFNcWuCZTAdq5NP
P5jqGoF63BKH2g0XV6qKja51KI3lkVn2tWgJ+hiJDBZNTOKvzKQ9no0tkCj7i9e40IFKV0+TLsIo
BTWo/zSJASavQZTNgL5HQ6YtlMV/vtmun7oMDWwsUaj0ILmRiSvorG0iXA/BNMZRUnP1UAkcCpFV
mtQZSlk1gtGUcwsgiC32h43WQWMyV6uUWkgFtbDKPPZ9ao/SjXwSmtTZfgaTydkU5SBX16/VECPj
/dzofcFDHTN3WaHskf5s0iguhtuCIoQSXPg0rmFrMX0RbNVmoIQen1c88dVyXie0bvKLWhif1o3t
sVPofVyszctEtCEuakB4/ADy00vqyUPRBZN4ZX+9RWYzRNPpl4BovTNsksHojxvE3fAtR5TidcPw
im79OBlWfJzA51YC3R9QKQN2FSsHppVQC+5B1iQBCWtOxlBqPJon8mSkzIAr+FKtgaU+4GHqQ/cS
bfACmK/wDpRtVsO7yD7giW0OmR3In3APuoI2ifICueOHw2hj5PsEVj845zyCmLbRyVba0kOVqjFv
ZzWfeGRBczU7RQD8lOON7o+S/ZnKWPAXvqYaeJOsjgX9WiCLA4ivl3KkODiZ2xZvXiy+n2Z7jENT
20hmXRGS9KGZOE7wM4Zsj/9m9UjrRwYtaouK58TjSCLjxzaYGOO0KAbfHxHi4qJ9dSvncCyUZ3/y
pA58ruk/7KjEgptb53DLSqRh1GW6UnfMHWkw7W/Osi4InZA8/RP/5a1dvzpm2/n4Yhry+ma6hfRZ
Yx8vixCqZGkfMn8nGwIDC5VkiCQvtpBZq/bDdFEA5NI67dn20UssA+dt8W0G7duVxlH6YPTEh5xq
t8B191dIJZAQLq44vOBHPOcHvVI3o/Ks2NIwGbShmlTg1o2MkC4Kh0oGWkI5Wl63uZ6UyVOmowCK
N8Qr9ksBBUIx9ZlJ/IlXxljeVPzjFmztr1YdfAgmqGs+W04BbHewyBpIxOGaOxbslMHOtPx/6Y13
lNjTAGV5KweZ8pcaldHsgH7Yl5hiKbUJrGcXTfoaHh+FmimQCIT4WgEU5DTFbV0cMaPml2UKJH7T
nVKWY+GE6MSxNFZ2Jsdh7TQrL0JrquCm/8D5y0V5qmsKRKpTwOopB54/FcDW+AoaOP9K4EIrS+FX
53Xq/7V/NI45p+FnQmipwq8PzXADX6PQBOeIkPG8lnxeamMiB6O3PWLBfbjOIf1j3B2y/HgsJOeZ
I8yuixo791L83U5P49GalhAHWJPS6KSmPb5Ynbk0saEr0Ulsl0YhDZ5vhMkeQhgHPXYi7xGbdRNr
HPR54ljKmcOrgah9kLIacLMqYsv2Eo5DbEUEqyS4CjXtmBvXhQq8AtQCEdsoM080nOy5SVYw0JY/
4t7mo29pN0/gnOGg/cIKVI92LQBl0lJ+JRfInrcxVtrCGKXcbi2ZRAodVY/TUWMRQawwekE7WwAD
8TQDryDcW5uJ5EEEjOJ6LHOwuqWdh+BSZTp8Tg44wutWz0f4kPufOFnu3SPVxjF95KWysIq41ZTc
HwMeOzOJHOfu1V4k5E0cG8pWUlBvfTRCihdNBDsbZGn8FIv8HDKOH6/4k6e79akaDMChVo0wwwJb
3SU8vN0JuVLSE14tb6XOZi0ZrkkHKFM44NFo9A0OoKU7OJJqJek5anwVE7/hLMgA4HL2+MItx4/J
YUT/YrHzlJUx2A675ssA9XbIX6i/98lD2Qo7O6wr/jh62/JbZUmsHM2RGN19YRJoY6I92gVlqha/
cPeOvmXMBrsyPrrnq6yg5K42eLz0fIFCXe0PELHreRzZlibntR4Sc3TsAnRlrYcOkm4ffLsJzK5z
/9ylgm66Tu08/6FWk8uCSEHCu20PQe8N+1lCC6qOH4Bn1aKmhgpjla48+77Cauupy8p3Zk/maKMT
5WolxDGv7WfgnikFYIh/pRjersa6au7O0prf3j6eGnTyP5fzjXTauDU9PXUuiCGxiv7abwN5P6Ta
T0i7WB80e8FokjQgLGtRCOyamEt0dCsF9cL9Z1AvPqwX+ZZLzBPBh2oxer8l0QcwxN0S4CXDzs+E
8xEWLfY2GDok8sLofaM2lapcnT5x4ZpraVmd6RCaDCErNrDHrbL+bEa+2tbwGn9iJS0kHEnEZd3+
QbAZkGr1BhauFD9Fjtal//cHQMa4daMOrOcMXjLVF7lOeKE5X8CcL9ys/4VVIzQ4O2LqlecS5h/W
P1Z/LukmAUWX6vzMkpHT1NIbV9GiJArMbwJgUjxglGF/C+1QU+N0ZnQoVdNEYX7d9S9S9N+usv/t
D2q6ZW+oYPI7OQGnmUvTJQx24ypPiwYn9LTTtnU/8ZH8QU2P8IqmeSK3mszjZbAUkKT00Rwgcbog
9rvjDJUVYeJO93TGK7KxYRFOa7spTnwL9BdTuL9Z2Ll0W6T2cvT/olqS95UfGg9WB837pPZ7ackg
V4vCUnpzsvlYFR9lTaH8pm6+s9UVWW5ZVoWA+UYu2KyaR9ZnosL5fMFkUEP+EyjmlR2dXNWNSFuc
FW+Kog84FyO3wVeNj30fT9FfGKF0cauylpx5dhPpc/gA0rnBXADExhJOCRxtzKjVJaL9bLIiyiQB
J6igOSOq18nO/5o72IiOmAGGL9ZkrN2M18FUwj82PhFJwEDy8NNHi7PtybRe5xClEJsuCN3rE7pL
QdYsztNzVjsa+CvlipMRkO4Sl4x69OQ9poWv5O268tcBJayDeNWo/CyWzLVoDpiHoxfm5B2yZpDv
TwteGk30zkNYCJbwje7XDBVo8WdR8oBxiVUgX8cdvLnsD8dDstkOFgHh7FhZ3SxgDCIFYEhUOx+H
SNjzOKggJwTGpql826desdEXNidCmNGajweu9f89ybwtd6u7Q6Lh5kYdmNGyy2jpzrPDY+xJXIeT
vYZ315+fHndOwo6BCS1PPTt0wXAPhMoo7Z78Da7hYfu/pt+3SR7xGuDkUfd40wdmgjF9W2Gzkaal
mhZvDxRj0H1sXHoMu0X3Y+qhIQwo3zXxDcp/GWnfm8DGl+BOCeUWSZsRzGm6eHFZuWd/XqYkferW
LduI36lJVUh0iYhLArSghWPQJYkN/HI41qDpi3CD3fpyUnIMVJhwfVvnHOHEZL0V6v5/gv7fK5fq
E82AFSvfojX1vSeJXXIfs+gCyxXbtQirKY5lNEmJUnB6NmmFDMInWfNh07IFP1mQpjjo3WnbSGSZ
+GEIyK9xWgISFVykns2CpaVhMtGfU6MdEKAg3BaiRacR+VxOnTgYAZT7OPJy+SAC2ZlmYDT7OVsL
TW5RruPoX/Ea+kOkf2EU7ug/dKdUwTCoCg43FKZ+QEhcFCRY9WeAKb5uuA4mTVpKqJWvsP/XL3Sw
XVva3L3MDRkVRBvw/cGF+1Uf8gHXq0uo59/XL+/PA5WgYcis0vzgMjbHiDvdMhOM7KLg20ODQv8k
fmUnoKsbjBcbXQc3EjR1UJUm7W/XHEJbR+QpUqLOGZ3nOkFIh5kZVi32IFrf1AHUxgNLa9XmdLHQ
5UjnOPCzGgd6gTOhWuMM+9DZuG7LW+ELVA6x9jIz8ipXgQ6YdRxUX8HrhkG/CqtQVfQUHdUWsVNp
9KMvjDJZBz6PKwON3x7WyMJEvGPutSIsA9lT4lVCN2Da8ktpqD6o5BaTHTNnsJLhhXsmJ9XhNwXV
G4vfeB0TQuFYupQQNOkLzlHLsSxFsTh1U28XUPnQp3oeL0AcT3juPb6wWqcmwdbVVWnCpfauPIsb
frXXYpxNAPCS+QYiZjdQjpiY3AYw9I8P59bg/CeJTdNQBVn9LwdTO2kzbIUrlJtZ7RzlDzN5GLE1
5G+NtoBvl3JnYk9Bjciak/Etu+H2+MF0/q+mlSbj/Ws2O2G4SqnPcHQrK5srpvzBrnkmaN/KVmLD
qFB2K1RU0J9AMbDGq+EqTcuGYp3UqEVZzde1u9cgy7C9xQv0bEK6sgBbch9YGwToYkKYei3/weZR
KdqXo9lwXuDmh0W9bK2J6ytC++2a8Lg4MtFGGMUHdsxjdtvR+TGiSCCk0KNNt77RISTRcsL3WjE5
HFiT/P3yT99FY5hVtYISXUZ66VFSvI3TRoLbQT8a5qBFfpCFBimTew25r7PHLjT+5hDMs6XUb3Ex
Axy24zXUxiYwhqzlEn8yvG3fMPCnTCkBLZH1CD4uac0oY5M30j1Ti43ULIuO8Q1yOFd61SbwdC4q
9NuQksDBIDt7eXvxFBDqYBepFSJ3urDQEcPC/cBQ+Y9jLlJIKyGOIIIj20wORfabzDBmzmLGTX6j
SSMUiEmNx53a1F/UsgqJ5oX6xOhsGkgCL1HO3lNKBEVFnfIf1qZzngZ92UjA/twHFWoPWZQ8atc0
YcuC0KqlUsvX706NMR/7eZt1LfnOZti+M1kHDq4XKSYrQ0snkMnj9MrlDRQeC3MYYhpPcJmcmKpT
2A1eKkkyowvRJFdNbgFizV2FTnAWBh+h8gc2lJ0BWmvyB+JJwx/rzhxskxUvE8ME9bv2BEnJExLk
ro/yERQX2TLJpTQv4atvsrRYbh47186IJZk994jRIdUdJlqFiUPubmD3JQp1jV//ADb9CFWa6jWh
zTBZMXSU1W4COYvjqrORruLOJWwDFVz1IZwB9CCY0pix8fcFC/axFi0BEOOM/3p4tJbSymUQJr3i
NxM8qs2wt+jEfa9dWB+YJQTtoJX0DebSGouoWAs11BisDF013rPAS6IJAq9/ucRlUZNMU7Ye5RJk
LKc0YpEhfQ+CGi8GzJn78R6RZv93WlCT7O2db6HCP3zgA5E2BvoHkkYoN+BFGBqA0Z2q5Xt9WPdo
qKCi3frdQqXsUSgHRBHOTaarGXqeoHAMi79Oh4nDJcREW9Zb5n6WfGjyEHPxl4W6wo3yRQzB8YuB
kjldTH5hsmYfDZvUEWTqp5wKZqS7ahKnoFijcnjlYODybk54fDt/nvUATGNKiE5uZ2bj7yLJ5Swp
WWBA4Olrj0iEXVpxKcxMcf7iG4FCD2rgiTL9i86ai+yFCUD1l6jzoQIDwok2UQ9YnkCe/SApEz9X
obNHSyzbnnSI+b/M3cdHkXAB3e4MyS42BOzA/PnaKaaVNZLcTVsKPbA6613K20IA+BeLbrEk44aJ
W5X3QLkip6WevdWUAsVi5XyRFWCmaeKIPAQPPmyHMlS26lmhTXKuInoS3R88W0J3BuR3AIWa90mS
rY2nBjB6jOMBODn0SKg/+afnONkg4MQ6l1JdVsNp9iFlt5HS3uMGrhzG3gbM8uMJ2XzA6p55mq5c
YHh/mZwJzTAJPGITIVZUj9XdgS+WlNGuz7E3OZFxKnRg6EtNFD4TemkWOfyojPyQSB1R01DM2F8w
l5MUcDpi8tRFzUo7AXYSBRlmUZNZFfhjnZj9tqpLyPKTLDNmlc29EkHLT938qAYD4I8EioFhxbOA
HBcLT3PMkId570K/yU2Mk9RYMSE7F2ZZwOKDrvneyPcScAg6+S+TTx/FRLVnMaNSwa31vXZe02c6
i8ydrga/O+UXPJxLaYpl93laJm6ST2lOJgCE1JeZz+xBsAOzgOO02R3ssdXUGuPeD6VdkbY3upgr
mVyCJK1xU8tPNA0FvUxKNb1imiRh0q5oCzGOhQbRA3SGz4vgao12PR/LOJJyUrFWMsYrkm1qF1As
Ak/QYAcicDmcHPMZzxZ+iEGYf1sVYYPhCsUlSYuQg0untLWvlfO9S5Mtmb4pfBsqfRpv5EwV1mzH
zKSU1JJlWU4KOa5vDJxZcxge0ek/V7s6KEqbTi/sIwciNM6sZtYY3V34AGupL66xd0q6HPdo9S79
omp+PoslP8vhRT1uOY7YKYRYVPZzY8J/gKpy8ZKMoWTjKvxxjVlM7xE2WXgBO1tD2io87YAmNziO
NFelE0kdpq500wOMlsEvEiUF/gTsZ4LwFDzEgjfNfgHcOijqe8bI5Z8SajrXUCKWvpQvhExu3bVz
giPONparlv5rZ9tpjVhiLagEJPGBU69l9dlLP6VZeDQUp9YmW++ZVaoEwtHffVoeYHS8Fo5DMTq9
gVTumQul7IRHm/orICjwc5B9jlOePIbiZE8M18mn8YdV2U8Y5/0i7iDV5GY8gMqLCpl9JYC9gqbu
ATVBrRizEAGZLKeLMnx6BpzxodSEoTil2F9ocHN/4EZvG/7yTLtXq5GMqh9tR2TtZDZSts85OMFF
h178KUW2aT0XS2Ksf655u54F4mDkLS6A4dAH7SKfx5Vhp+QZkqJJolQdXE9HBumXOA02YUk0kzfw
b1/sCfQRAJmEx+Ylq0oviG48Ch7dTGHhzX3c2oKXGIiPfHYSB6vAeEOEV39s9Byiu9kszV7QCnQr
dvjtrFtHU0vpzhPlI3gUNHOHvNv0t4cyES21Pm/wEdXQZG594oL6AmnkkrKnzcNEMhrbEmVfrBUM
/L+EyBVgzk8UXM0h0/abFAS173Vk/b9ivKu92+UXH7fA688bR152Gv9JpnAC7UUiP5r67l52xQPQ
sRJrU6tK+1SU1W7LO9OSbSBfoH629puROtE794jmYszDK/O/yhPqV+fiJibWhW2whfnH9OTzGZWf
dsYLHENC1470jb9rolwA1Q2IQC9+rDNqw8zyL2lk+dVha2Lk0YgrB2ymGpYtr0pN7gJ4xoSE+O4r
E5/TkjO9+XQa2x4sjCmZx35Z8zTfRldWSRCxoxuFRd9s7e4eDqMNWkGDBG579YKDJIgyklA4Ohuv
wejAg3f/QziD7eItsZtArwgd5tdAium72C+9EKmN2hM1TtKR1cJN/Krog0555hciKWQDKoU9TenF
oQKCW3/eUSYzZ/OKFBK6LrNV8k0YVXRT4HPUaC9XyzmwTx8X6Rwno17dIM6F1y48ChaGTR3H7CKd
3nWPEcYO8pT6U6mvl2Z0zX9lrZm+dIPX8dCmu4gQRfF5ERXh5xqK9CtM0R0ZG0uQzv6zeTZUfh0n
jJkty0obKjOF6UyD2tNdW6HVRTTMrmrvaMOYY7m3s1NWHqAlzxpIz1biiR296g8Pe1Su0isyTW/z
x5hDEfG5mFwes4tfPiAkecgT5Qr+gnYOofBzZ8OBmBFatdTTd9rKk6qRQy8AjHQRHHgGeOnzjC8j
PFFViKVRTANmB+eWv+mcuOq01t8qw4dgnUxs+hqYWaS0cLDOZupqwcVIZ2urGZTw8uF9rPTbPPk/
jFlAwPo3QlIfHeT34ECJZ1I3Xi+Ad3GE890Su569+mc+BczJQuMUQN7W0k5YNwYfHQ6hrvqV0YeP
6Kn0NshdGMMzsR8tapuwGEPUmc90WEDoxHkh4/++EN6JlCPYMcgTaOznICYRorFzSe2EJ6Nk91bk
sDl+RgxCMoKrcF+uzE+W3HGw0Ba1Gk8t/yHadmhmwzqGa5U1tJcNHwHV9DqxwUhT4RRapl6WUyrf
3H6kPu32aP4GVi6tCZIeqvA5wRs7WzGmgd+rFZm2VxF1v4/Oupfkjv4mS7jCrrqvj3WzSdv/0sF1
3Xz2Qxn+UMEk9iebRqSp8frOrA308D7vV4YWXe6u+ZJX7kmwYvN63u8x3YE65E/c+VorFjHxAIr9
cLjFLkkc6cvIf+YLGi+smUknLEMHEHTQjTYuiP3VlQkS+zx08oTASNvV9+GwLIBT8yRinWaYverC
IaIQ7el/K6/c26BHI8poNMvtkkCUAi4emqsulA9ryqJ87lgKMJv/bIg1XNccy0d/Ax11rwI9w5cT
wb3Gjt2eOyuuNf9Ibs0uaCUNAvU3O1kSxvbQQYDtfZEDclcVqnC2Rww9fdFrFqV2/5JhNbommY5y
bbzmYljDNWdhyWynzOeKbZZL5gn75v5ssMuHo3J1HNqqAMlwgdXthzyj/uwaOU45IoaxfmKnQWq6
yuWtLmUsvfv3qvg67cs+dbuhyn9qYHENs5XycpqncW3+uNNkrvaOKGGWVZ9N+lDZ7+U7N0pszfHE
mUXwa4icb1UXrN5lKMsTssv9DGfygiV0oudpcEQYtW94h0JnoymRHy2/XIfBcTQE6JZDUto3cUTL
Y7p76yoOgsan1FhF9RE3tUay12INaSKrBHIQMcEL5SNpcRAC2QYW7NlSG3bOR22rhj9U2Jhh7bg5
tjldQxLTCz7/LPAqYRqIOkdsGiuErxokuqfwHj4n4LmFVzvKskhwhQ0UVr0WPkGRNAk/GCK6/rmD
0+9xXLcdAtTAkyvtpDmhxizgEP1XntkgFipG/3/y7RUXbeYvG4pM66U//7AUjvhy9rMZeIXysNR5
AZGRDnlBJ1008fyxNRPArPPp8zQAea/M6Jq678CSKGJUNILk73cBDBT2/W3zF9CdtYMLeriMjTgG
7fPS1NcBy9S0p/lp6h21vNCvchMfQG+tM7hPpeTfQVMOgf02WU797cXyEGtdjiEGz2JItICNciw7
T4czutnSTPcOvdhMv2xhhAppsmdZbpxwAP5iQoUEj2Kd1DBbEDbeg95I24QDCri9Ky9z0xzCuTn4
xQU7x5mpWIZR3JX4Z8hC0eg5iw0BmAkRo8KAAdSg7AfiLL2mHrew+dTMlulOJyqL5JTQ8gUFccPg
77V52fqyVG5VRyaKG2xq4NHRQpWbdxSjagrpX+bp5/nMmPnbFYNJT76ee82NgNlHYjpNaQiyZuBl
3mUzcqe3+mVuHNuk5vWhc0kTQMWJCtVPA8g6FyAqxdb8I85lw/hkDEgJg8r/sTai5ORKvQ9PR8yv
+BkiY8826/zUI0EoIL/UCisYb7A96FM45k71nYEZfQzf7rZbamyG9Wit6fD44zOdDMMwcXCVNjRf
ClV6F2v5aVH0AxdQfE0rY41DEPrAlFPoElT1XPRWeAhWeasd86wnh9c/6lwhEQRQ8c/gaKKBSJ1E
EQykGP0GPSVRl5Y/i6PJ3OTR/x/CuLT2CM5ZeTSg22RJuve7wesAV23+Lt3n+Es9PUWAqskieiTE
tOs4RNDXtO5aBGy73eXiZNKWntqkLJPviWqY3hg3hM3d976iGMnx9C9oxnU5MGlhn/B3w/ycM5qo
K8SxniON0TpOwxHL+hHSzqlXdBRrVTqMGn3t2Eq9l3OYpYeJDH+EnvP80YSIaw7fyt7r/eb/pAiX
KWlUas/kbD4s5vWGKxQtRLJR/2TpdrRHhkWaqU5oE44wOlXKUwPZDvK/e/TjSNTZZ887wZk+rjGF
ot3wHR9C0Or8KrWoA7nof3HGEFkT7Lkypg/Fc9KSMo8i73+nZCMIxpLz0A7Deql8WtoiBOMgTfbl
UvZ31ekP6kEyYl3Eeyf67S2yN8LqkLa7+QHakJvGEpA9pEovDQxY++wD69cbQNkpDYkiljlPwp2i
dOrMPuMj8TFBuPbZhZIuRLKHuxI9dH5XIFKXrBH1wpQa1N2P787ilGWRddWNYQ1NZNSrLPv04zXT
OBYURbjkY026VBQVkzU96NMqYUzan1oPxp4C7AGQQJMCNhSciOHHIb2eTuQqtHMU9KnZynOJ7aEc
D0mFrCK5E7ejxmrzdN1aym8nfkvyUTxPTOXdXlEskM0/Ee0NGhG61VVW0+gELtMov1EGpuJevGoI
Tgdg3wa2bRM4hcuh8X7/cERyvL/E3gubot3wN0j/CJQCBaIwkRtnp7uOj4HTdy8qRcJbqwboOsGi
/Dasu7RFDxq1MRd2Jv1soU9JPt8/RipflEPczesfZf5SUQWMXlWszE/nefWqZqw2eZNn6THBKWWU
+ZqUM3eiJ4a2DxFkT8XcC6W5eWtWcbcluYQY6HbmD5/pY5qhxWlprq5r2Z0z2r5K7u1wFuSxO2mC
tnV0GPI4oak4oHero0ZDr3TaV2iNpqtnCxuOs8ZUetlzITbhTh07Ic8TqI5enrzGg6CKYDoiYcoS
5mUXIm7K6EM6oJn/wjxD1To8+W5wiEFtOqA6HZfZapZfZoGhzbRx68vgApftFWPvt8WdG4uyTk9V
Sa8hMhZsn7u4zk2brbDv1epkMcaEJHMHFRPbUjVX+qFMstZI22BmgRORFPmvZ8C3B5HYMJECiZ0j
XNQbUEjkC+Zp5KyfK+Y5bGEZY54KexeP8jgbSIk71p+fj+x0OW6SwQ71XsWoUW7LR6NBoDsglIxK
P7mcFEo5C2VSYdIptzDmHq2AVAlYoGCMZ0OWQDp/B6JhrjwmpHfT8TzknEwTa/nOMUEmQP24lXIN
Z0OPrjjPLI0m6IZtH4oN4ZOb4rPzgPzXbNErFnb334JEWXsUwmfI78kDfD8nFxt0n5AGczmL46Fb
iFcFlozyTrdCLwn4LGABCOB750LYp2S1ZXD6iGCx5JJfAQprxqY/6IMcGcWUE2bE4Kh8W3u5heN8
6i423qoKyIW3NYAKE4jKp6YWuo2cjuiHY8WnsYQilZ9yAVnJSG8aPAG7zn9jZLpbQvwfbeH/c+hF
Qpl1wdUNS5sHyjFes3sOAMOAPgVovdFIQzRYBw7taWLZCkmfklYTfx0h9mzUq7Yb7zFeMq+sA29F
IggZHjGl2eH9wfOh6VeVBy1F2NflvzSHiBUrbAY1EE47L95p4rbq51vJoPcc2O9UNvbxVzPnyos3
gwDtq7B68j3W+Nx+XTV5Ov4WfiehmkV/nmbf28o164LxH1JUbVXeKIP8IFeDSDX9LIbBz/YQ7US9
poUD7U0C4Tc9UlAZcg5gMW1bIZfFZirkEg0LJ+0ooWejl1eU2fRiQzt4A5K02SXj7Ey4k7VXR0vM
O7Bp/GeYbhlnZLTVhsoRkzHauCfOH9n2VaF1NcC7+gTBdhsEDPLBRJU/XcCQphzxz45ZWb8gRgDm
rA7P06Y8T7BxDwbYzQgU4MG9kuqwyLzgzrDikjWNJdIrXvX2uwMNE5jlR3m8hRTv/SbX1q/aH2jC
1+qwoLouWxqkVnzyXaEWO1XhDjRJVuwvYkiYMjReUHlIG4YPi+E8NKoWUOUNJTQodtVSCciuBI2b
JJRJsFfMZMCTxe7m2UlZcZiyfbFB//EiValkL0yndeqcCp72EED+d90SGMxfR0uXO19IdiS4zm18
mZ7etSCk8ida+RChtEV7TRZg9bjb09A1FbWTy5CTETOUGfFmSdvCjgxx2swXnxHexlkAbGTkxgBz
KQpUxm5NTPqcKZtO//y7BuRQjI2JwbpW1tcsf1mezcCpVTXihfxoc2K8wMOCg6I7fmNENjxLcNsY
/ZUhWDNXb6/+LGThgU3oIcusv+4LW+RpfcCAIUoHlLqBWBTSfBU66WswWHJTq0T5R3RmKC+AxPGz
JbxzOSKWFY5fT0G6KhDeTY/o+KJ4RXMvZBRo6sxM7K42MiLayp+KKQ1L1MA05KO/n+fWfm2KpmuT
a3VQoPAcI2E/MspxStveTnki8KxPb2V1zWarvrTcYCkm24+4ESoizV3YLIVpLTUQOMxRdC54I6GR
kw+g1FLUXPzLtLE/EBJUd+LtBaw1a9xrzZjtmSe3nRrSRSyGLx/g2/0o7ERKfJh8tQPBEoMqZGwY
yOTFqt49KCWQXBWZoRnUtRZtnaOGzkdOnoRWzCW0uFusOeqp609UPSD3VTGXK9OS2doq92Cu9HFQ
vKVhgVgNyC9rMh3sJVUKRkBCTqpPA3Evrs4UI4sWeUgrVMHPLXiKxga4LeZYDk/HawHgTh9YmHRR
8og/+YnbKdWj4pJWs8s4d6cZYMkrDEnZPyyS/skJxqDo/xi5Yo3eFJd9cUEpxVbAMu8bfhObF/FD
jDJUqIOyRrnsuFtFK/BsuybYz9geGVd9cUR8iM0w9SclNKH5QuDgoRfCXpgke8a43jK4ERKIuqvG
MW0aKRqUDivW6tt6y4M7H/f4PP4YXCbGIvUt6oGVTWzDkhdCAtOkN6fYlMUEZsXG1jDgELLxGZuE
FT6qI5NY7NHiWE9EMAD9Olnc2+rvORWtGI9jOWe3fReEH6hxvRiX3BCLICbgGybpBhfvnm2q6FKO
tYjOfaF1sve4IWcn3I7R8WHY1wIDiJyERoGqH9O/zdF2kQ7uLvqWtnXMqLTjbehQe7O2n3EFETx3
Do1QaRHPE2Estz1QyvGAS02uWKyq+MxFldiIhSj89HIOyMsY1myJQwkUpaIvml68Nd7shiRM0yRb
hq4aQRWowrzrRMxM84t6tJ1RSzVlMGFSLpVSYpXEawzVSTzyueBfa8kJRmFt1/UzRYb9WuHZTUv1
T8BI2fq2veCtbZ9KKC7lWjDiSovm5QbaQhzufzd6jMyT1yZvLZHpcexMtOjkNBApQmpavOXDdM/u
7nteBKsbQetosl0N853/IhHueKYM84k2SjWsVMl9pRp/D8Kwx/8lNQTuAfVJ/HCjQbdwOkQppXds
Ck8x97eRI684tAEX1KGk+oO66pzD+51vED5fTDnZuLkAaVHTYBeUVzG70FAXxliwb6sHn8dILOxs
N7QmAzxLoTIRAJcSRNgjt8WUdYv+rHgyID7cmGwxmhVRX+ZYrm1TAA9yuSHUdmf8sUmK2NOBYyvv
xChCir0S4BYlER9APOMpjZFmtF3RWtJAGASGzg1T1rV7VqDYNwUf0F4WexXW8hL1aK05pSzsb5Wh
8BNliS3HOS4xG3NVcEwcPwHO/h0MKpv7gxzFsfRv63JHY/PW9t9yJ4xuTEj2Xw1pEc9NxJcdc5h8
+h2/ZClsXjA9j4M0GmUjcUsPkA+9eepdXA4CE/CvzW/bBJe+h+NImFPQjTSM8RYAcp4jeP64e2ta
KxS/bzDULWqwbLUsijijDz2nl8xtDPgaZWBkbDG5maJmAblaP7UhaYrHwsuTeRLWGIrIklk13DRM
JVrvMAdP0Y3l230WCZdG+iVj6LNV89KrmFD/zghkG/GrBhGNuL0412prNLpDYELhiI5Wdz6YcjnR
7yzH6NoJYtbEJ5Lx78Y4N8OX3gP0hr+t8FbDTegoknVepEZWfMDmS+ERxRF7uEOx/ZpvlLtTU9n0
WfIp95Xj03L7AA5xA/hbcd3lsbZcRYhfA4T0StW+5c/bIOVhWXR+lPPeW7/fOv3uWHNIUqz3tYtB
Nj5q43Wf2cTmDeP8LLRPSuDvxUo54A+Ig7z1675IfOYkOeHIpSv50HpNkdal3uGEiG8M9R8MjrP9
kBkOAPMPX/2an+NHuY+ILwVloIhab5y0Gh+h14ZPm6ibuglyTkhyPB5l8BRai/RPjyG54HDvt02l
fvc8CkZATl/XpmMUMFqcNnk3k6S4I2322B9GTY6Yyy9Lvr5tq8s33NId0KeaW2Y3+w9C7mAMuiOJ
tfIY5lOLYxhE3XUEtlILe00xfXRU7g0KKXa7PqKsa4DBuzCAmmfsK0TZyp5tXWmk5NYiTmbTNT53
sdqtmB8mqM2/OrxQxru3ISSPlloNFlHKfrYcLmRUnjq2G7L6oKB7BkfjQR65egWNfsU74WMGh69h
lXCMMgIXRhE2JNqjs3eP/oh7fdKAJwD8c4+0+g3j8WSO7qIXu3a8yWVZSrdd9Sd67HMs5f6B4WX2
RIPxzkKX7qwzeXkSVU5aEfgfvRB61jGDV0zqNi2eRVZzEaGDPexTgk3oIHeprlbpQaszpNy+uYuR
ICtCd/IrzHNfUjMW5evgYiS4lQ2UUSGnHpSpiGRcawPS5/pPXYVm7hQ4eZJRnmVTNf/fKx2yhMxE
YYaoi8CHwdMO9Km+iycKySR6zzS7df8GzT3/Vx0sa8wehbjOTYXPAW3xW1Ra3MLAnos/JjyidFux
ntUEGEldZ131ef5DgN55cuh+UekqWIiXvEBAa0lXINAp3Jttc/thEFvoLdqFnAox0xehgIGIAiNG
QAWDQS5G43g47JzO+ZoOMu0gCZ0KU/tk/alMh+kHPBHtfVRB2x1oKPuN672FiGgJ5aNAMgt4YiRh
h1hVe887vyoc5Xsgi6/DSfzjwRaeBMqiGkYvBiKncbp1GMO1tBzb8R7WiHmCn0PrX3uyPRXKydxt
+2hOrapp2PIDf2rV2/bJASTxTa5uF/dPi/7rQmlCRFk1s0Yfoyo3xZSrfLSTo2zeadWSP2G216Wa
5kVRRDsnThvaJ04kBehUZYKsmOUQctk4AKENeuJilaAY3bpfRTD0SK6mXeu0+s7PTc8LRRWaCr9J
iPgPlqxWpXuz+LsBNhYW3L3D3YNyG+ei8XiXOBRi6gUJHHumV++u72GI0sv0PcYaray3Vw+cdKea
+V8bRBxa3bZrF5VQR5kU8utjLJLEsxT0RnFNO6KLCGYpGYr8OzcqeAov8JA53vez2kcwfeIuFzyO
lBJg4HpSES4h4UthZBr9PpTJSzsGT06R0RDgtKr7vDv0tWS3LbYXtvh7U+MZzF6P433veQf0DTpt
bU7rL8L5DnWmS89SAZZSItI9SSLHUsEOVXim/Gatv91SPEaIEsIVePCkimy74FPEh1Zjctmf4woc
+p3NUP16E6wPTRfomLthSpOOdvDF8J8xFCzLraHCS73c0pMPHQrW2D7Elg6zjU8Ugj+1qBTF+Hr4
5jQYORKEYQqXvdeEsSPyMEzD1tf44IJ3OH+56wmNBCn7MzFD9g+Dolu5s8ncedf4HhR4JQIuEuPU
C8KwYJr2X2/Stbbwl47dI+LAH3mBQwEent1jLQtkiwBgVUjIPbl0okPAR2Fv2dYlmRdJt5p2Zu2o
rkS5kZaPDfUwtZqL4WgemVtVnH6bmQWnhtjGRMFM6bmzKZg/205CwonN9/prAo3jnJNnYxN8609D
FUiwz+6QZAnrLLJbpi3IjnCwPdfYuLFIOrg6DFRpJPE3BZMDmf6eZHzeBfypV1ffnQVwmN00740J
Y5G2s+lAko2PUNAnDHxZJaoWdOheoSD/cnaiYSqKdtDK9Xf0B3vBf2PUHhzeJVNFCqr0F7uZINv7
N8A0rIqluvr80n1gEFxak3m+gUWvc9PIV0Et7qteULOz4mB50OBnbfO4HcFk9sHDhEXxkTuAVtGw
dVwigYW2zSkx1Q8N7MNGX6I/oXzykALZUaZmoOxB13TmThEPDuVQYn37WQvqSxnvD7ZhBuIRvioZ
ejwiCDV4FjwEbijvyFr0s2zAfKjicBlUeczazsmbHr8c2BCB3juEhdQjjQcY6pKanwG+Vd1saxDc
URCq/4Zzmlv99+hLWCIw4Su1bqYsKc5lfD0WtwDQqP2Zw5JtVROEQQsJ+qQkJy3f3yob/6Y9/Zuy
pq5FtmdFBnViBxijinnp4e3LV9/neK6r2DvWt2KRW2F9V/uqYUB0FZ9DMRsy42KF8IAxQoYHxfKk
TTIQfzVq58y4rC9HHbGFc0ENeaLO0zpChcu/OoTRs4GSLIi4SGFpofRYG1Tv5Pnu1f5s8BHjpEeF
vjGkDlnb9tEwXA7PHCtpUh/fkn29jp6xq1wu5A4UFO+CjHHp3u9ISN/eEexyIn+IlV1DR0uwDsy/
pGKvrKqC8l+vPySnohII66yYhOoqU4ieYqhQRbnH1fLkoCJYGmNeEHMMYSfqpU7OrNuQu/0zTkSv
zOVqDvCREw+eoXVIPIpp59bdMYNENERZy3+ZXbQGzSqW5gPFcB6JP/EDFmGQYoa/6zAM5+Wl/9sT
csBWcKib6D8A/6zf1TIPnKOH8C0TGFIrWUbtRp7YiLIa+qofrIty6GInJ6ZJr4RMeMHXmcXKrx5o
IkJYoNiqYGU7yzoOkJHF53eoG4/+ecOQ8Ro0ZEQw/JjtGjOB5sHXouo54uEQffmSTc7lG2onxiDp
UxYZbf7CvHhUvOeH0mvkxCYB+5WQOm8divkFqL6N+HtSZBMionbQgItWe5zlN0RGqI9BwuuTUQVH
muoSU9jKPj+7tR3qGd5z0tzH+4DLkiUfCZ3lgTyypVWD/fsHuym4P+HdpCw50hc8fUdHuuM8GKDt
lDep2qwQsEvm7CuQPnnPCOFFh3TbbwVGmbbEn+yKn70Zvxs69iFm5fOnFX7kexNJz6FENeJIFvzz
c1wcWbRjUbaYBrxiCPmkX5BIQjFMmMWVNf7k5yMpYb6fUwwD75FwxIfUotlVmWPhBqFP0BRZuxBU
+I6n9eGmXwKxt7mSK5nx7dUv/fTUhldQ7HOZryMEq4O6x6n2NAIOn4raACGjgyRPQZfN3ddqdOFC
U6blKBijmj8XeXvKwqXMX7oKItJuLks8OhcCYNlegcVNEZeiSk+PAIO81fkS5X28l89lc5Gzfx5u
m4y4MDse0feyeuAI3Z4dZVN+Fvi/Op5L6KfK8CG/tFYfene4mc/kiKQD+9zVP1+Bsx/5/h1zVRyJ
myXACZAvY/F6T8vzd0iRwJPODfbygqVNw9gjt6MUegdlr7kP0yyHNmzWxhtE55EKxunKnETHxp4V
3E5LluHFSb77uhxcsHGYm56C1dtN3gXRO1hP9NSehj7SO7HOTxnlIF2huzt+AKMi+amcLplixNEW
KI79+INNib0BuZcC+nzpMLGz+HJ266wTk07i8L9lXHDyKJd86QbNXDVEjM1fCGq0SBzClpf3EFD3
w8M0SBo7qnQl2jN3qVAMU/KI2nXAoBacPsrDsmNovHr1Y4jDbcdAr3i8al+aGtRi3G4yoZcah6wT
htJ7ytKi2d4cJUAwJeavVKUWw19dlBSVMo5zN0NeXmTs9pMGYs9wHeNPgWgRSrybfLqlkHwko5s/
J/qBP0QSeiq4LXuct+Ic3T+aHJ/EV1zQ6cY2BxhPzgy+BiS5jI37prdlAmt1Zky29NKoFE96Q2lQ
D1AtVBrWrBFuga2p9eRUqu3gN/rEcaV7FH8lrNyu/XehT41fNd/U77fcKQGrgQkKJs1Plc67BFhf
M6EQ3LF9fWnPeWPNm7a+VPWTvL5QPBXUdozrLLV7jJoGOXtQRZ+wCt2zHz/Bkn7ncgqh/+fb4Rsc
wfDf5n9+KBu46q9KZOr2NQtjv13BgX/mhs0Xhp9Heui2SSZLMQ6AUT2Sy5MRGaHgjKxdAQzrtI+0
eFY2B490gjXScAaM2RuFECCSksu28wm+ABXu+4TZWaxQo7PFJlKLhZCjl+Enj53DNFoOhS3eghmG
hvxhOGSTRTmRpN2NbBUix3gNAW8H6Sf5/ZoRMlne11MeOpNSLeDqOE7W55axVoYxsVa6AUWdIK98
n1cUymonK6oBeNj6/N3h3G7hkU5mtZbBGVQWa8czsmH+IF+CXuIIPsNQnZdOE5DPssMsW+pU2q4f
3G2pU99miQ8A1kUwfiukcv33O97mSdL06rFL0VY+1m6amEoN1E0vQ4muZjOV397L0NoJ8o+9+r1Z
RBCRGqSfNL9CY0P+C32QNrFX0TdfeBIfpbLe5Z72xtNQEkgicnMm9kJ1ylpwPVNwq9Jhd+TiV27U
GCeBGnfVr9ktxnIm+Z8Q7VTUBH/1UkT9SrsipiILGjab6qd0jhZbGaqhA4p6Wng14LesTVmmHqpZ
6haxsWSB9iUxB6WbGRm0chr+Bc/XEBSFwz8u2WAwa1tyJ4iXYy4DsTOm7Ev6Gs3rhzTnglQNE7m8
d/0IYqfNTfZv2QRl3v5v0r238SGNXfOxwjYO2EfMwHeAB7Z6Gpw2RbONFB9N7YvEA5J9RKP+PuQN
n47GzPJ1lMMxBo0Aj7e1s5ycuT4GLAiMMy4Ie+/1iXH3fGyASbbM+S207LfeoFQLcGQFaqKVv7ax
I2Rcirz76GLvXQtF3zC6vU+ssdBHP6AasLy6g0i2y4hq8sWofMiHsuGV/n9jK2rbut+ug1oigSDY
CmXiwFjzGEdP1e3PtjQbZen54pDXLJAF/mUcuB0FCnytdclyn+I/0ghPdzCndf4rQhJSy6gCZQrV
mtZKnXrQFQyhBb8VOYeprIQ9V1MdC0U1itWF24rW1RuE4Mr/T4XQIWFKq9Se1qbDLu3NGfiDqyYX
K6+VYlPW28k7Ot0ezHC4oUib6BgS9Gk1cABnY920mfZM8hvde9KANnYV+Z+77KTOJ9W8gxONrzBJ
pbOt/Bo7KoSIJaiqn6kWi9Y7ZB0kuvdwKTxcK9ceHVTeiAlpNPhVj2j/a1IXSTvyk9RqLFlVK3tg
ImwxwLIK237EoELVNank4nlYgjz+oOdCrz/0k4YOueCdgOhmNVoP6y2SGydPeeqZJ9XA5zApw1sT
lOdbh75XsupNRRixz81Um8EPVM0MQlhbdZHCvIZGP0TBdnG7LmYi2zfEm04KXNtc4DEVLdg6MvIU
/Hms7hbKncBNYi6ee3y5ywIXJIZ9wsAeU/rsYj2Ww0a/g0vN4yEfW/tlLb2OzMT19giqXlK0Cl8D
Vvw=
`protect end_protected

