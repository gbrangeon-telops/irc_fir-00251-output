

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HUpwfbtoJu5ljZH1PD1nirfZUiqEH4rdOJmHG3byOsiHMKK3LegkCLnxPuPlk+MO+z4ctY9AQVS+
qDXnVNabAA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J5amwDwAOhmwY1AI7aPhS8ck8cUzk3ZbW/PSkoxcoFtS5AuFiIpCT9Eh2Lt0JzHUUKx72jQhC4xP
E8DYUPCIo40JuI++9z5fK4HwpQiCOB47OP9CCbDUXkdRdGgF4e6aIOfD40xCprloxnLZWVs0yawE
2eWpDksVPZ7exWV5yp8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kHeSBUaR4Gb9xyNR7/PmBoZ6gckk9p1h7+VOSSxhgJTOkeDKrcZOdIV1GDgFDrDQ7kzRgTiYYdNg
fXk4UhiKwBVyrTjV2sMzg3+WqoUQIK6Jy3j+rnKZ0FHbaJ/B0H/GfbBoAdHe7Ll2JvXvA2JrUnjB
cZCpVeHDgAOSHC+pzlRSIpPSacSQtQcR7XQ/3XaxnZYRC7uHkv276AbG3wIpLBG2zxIX3ZP+ackQ
pH7/JslwJLo+2yMp03WDL60KY4dKN4/3Cbuq0p9ZXqs2Y5D7OEUZNxyvOtt0dnCx89ZP9OSkU6+U
STforoN1MyOGgJ2YZ3QN/z5I0fk2RYpfEM9JsA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lu2s7AKqknRcUE5f3UmM0sxhb8YGklEChkrpjNpqeFmWrHZVTV653SjxOWSucZRxKRWERgvAD5Ge
f+lfXprxLknFOXVThhIZcoGHsP1dAaIYcRFINHuR+NXvmYc17FBsIljnkMKM4grLGNoBCK5BU3oj
+OpUaEAqYZcR3Ny7rME=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZNNygMQdh+aYmFNm+RRdz6IwBodkqsu7V9fE3BGXF5I2MBgRK6iGinaX8yLwnKR/gy2F4SnWUzqm
SM6Hy+mVD8IIS+xm7ukIVwLbM9+0zez0kJn+qWOW6DSjxPXqHRWy3fQI42FtwyVBs6pb7/W8Q9NM
y83XMjmhW9gbYNHIHq5e9D7ao/9WQ1Ytg4YhUY4H4cSzY2tHj3tbIsVO5Swzs3K1mz8KunAK9qzN
WNyQE7ctUOauX1bPhyKN8vZcKzkl7x8jPe9GO6BDBcCZS9DeY3P2LTqajNPbMa7b+rdlszJkVZWF
aXg8+G+Fp5cfd6qUK77FET8A+G+lv6qs6bNgOw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26160)
`protect data_block
ImqtntXWwDiZQUewAZk4ucR/htTX/1hdyhTUD36cpIKDKEcCfTdwHdF5tNP5ZnvQPqE6MJuIQNJI
dYK0eYn0h5tkURWINb4ZWinJY+yNYfx7yOem3Ak1eQsRebwLcjAJsIV+WdbPekdtdzsBE+xK31FJ
uZlI+eAmTy4925MiC0yg9sHRIgBJKlL1Qs0w8nDowYSkCc7u0BCdEMdTcXbiUkRQm1qZxJzZ4anE
K4nDWsa6jgHYpbGvTORLk9JdPZ2r25kWMf0kjccTvi3PRT/0DbMQK4Ffd4IWqiKtyXQuqGh9OCBZ
RCmFFZzeDBQ50FDXpsIMjT+abRYxKN6rw2C28JPDTxNuTVeHHC9cwWE/dZ7Xitfc+7ZRKTw4/O96
1ToRM9S6m7lxOvaiT0CTkODqk54V516lVihA5jomYktpQ1rh81QrirTWR4Rq1P9cFWgaZjdwAutT
Vy4a3FVFWBIPU9AcWc0c2ML/6/hvk/mK0EDPQt7+W3tO1G9wj9jKB+SG9o0oNHLjc+iMM8SUDlzV
j/4RTBGRmexAGXw7DYOvyWNM6B4i5W5+eGT7Z9dzJEUrEE0VlLVwOHjD8Ei8YYvpInRTKoWHGO/+
kEY9hHtG42Ae9VGPwZr8Zl2PQ+irlIRkL6AEYR6G4sFgFtsz6a5MfWFxrDXTb3k1v8GN0qud6hFq
PdHcN7vpMTo/DviuIo9GSTV/42DgBsV7x+wVtddyoPsTGd8mX4B2SuHCMyXIlf8+1mjQGjmljxyf
iG4bN7cHtRnwTvCxQSEayaGM0WuMdq++D2pB2o2KKa6Z5cIV9X5Wya7MPsp1HlkhMz/C755g+tqV
67SitIfUUZgdXLrpQ3pn5aQYExAOvyoVoS9Clr5qPNdOw1ZC4vJEcO30xpjjE+deo1w2C5B/nm+6
bQj9UbGhU5t8AAFrJ27V8cwx9iTh+Plm+zgj+yLk2yOFVRoeeuiJNmwu7vxW7IRYEIgor/zcLV6/
YfT6LMC2UzUjxXnclhUPoVTpJv0BL6Wsku0KBCR2/trEiRa7Uw08JjBsCdGFsoSUTP0eboaXSSGB
vgKzpf77vII1isAoZ6emWD3w8tX8Y6e+UNbunffKLZPHookYUJSGq4v6nsSF3w74JzpuG/JvWrNS
qgWkmPmKwjHgJKMxM85I4N5Yqwa1k7/g7/4bVsySNlkjtKVYgbv04Lgp1GrW6wCDoOjH0/mjkE11
2Og1hb+M2w/QTQcCvX9rdQvWUoTuT24dCrdmJa7iXqMMedBamYozcv1N7jfYWGUnOou6zW9y7EeN
TtXND55Cs4I0Ixs/36jWhCnGxK83wSGBBf5uB6MuwmxE96VD1cR7VLDD2oUeNw59HNC0uNXhuCMD
dn3UNw4W6zBq0g8c+jrGqFX+TQpTGuMC+RweiCydZeoBcUZWRcfIGfy4b/7ejUOICDzXCHPWnat5
FtT8Mnye57gCcvyjWt5HvJiNzFOL/yl9sx3FsVhoe4uzHHLEkbid4w/9iJzHmNjeZjqAne0g5GS/
akO0LmfFD03dXtJMU/u2nsj0eucqDyk3Nye45osZWh77rCYtUZIhbR3fFKKRNmrIMhdjbKzIK2T9
LGmMMAhMmX+GntzYBL3hLnBOcUFAFT6SPsuaFUFq9GDm5eR7ASkItneBcOPCrgNg31DJUi3TPQlA
G+lyVTfRDlZc3/+HFW7jLWi7g0U4z4ESdyFfaUn7xk0Z+8AqlUlevbo4qvLKouxrcqVPmNu99vaH
wH0eDSkzTYtor4HXFSHGIfIPqm4g0D8icAJPhak5h5v4ZnqhcnQm8cUPtdOBw+pngz1G9o/v8apt
fIWG2++C3AexsO4ekly9HvUG6SLiSeZP4HP9wrabGQJm9/xryxc1ZOmzHvbknIQkn4ZSXaGK53oz
nZCZ8++jmmKnenMKzCP/8kAGzD0lxCRyCXEHVyT4DYshluPy2ypa5YAri4RsFDxq+UXJWCfBVXvM
ol3hP+LzT7ye+Cc4Lc5fl9ZVoeX87TkTOVPSnu+iZY++ZwIHqgbCcc0gYSX9TYzlFk0T1VFPYOH9
S9UilZq0U8v/GmhMMJ1QbywUptPdwtQFtFr0YL5RH7CDju79ZQh9Xqu9SBWZoHd4IogDGPZvNCTv
AoK+OTdj+dVeQ/c1Gng7jBsi6+RDj+i6kVZlfF1B09Pryhw1zcUMQNbxdnJ980+ATX32crg65Pc8
l9Qh2riDyFWgavAslzXff7yBG7CAmsEw7kNE2YZ7yGyv5ZPES8VvQaTv/QzS0ANSlU7SE80hbZhE
cG+gJTnJYRDOHmAUFdjxz2EjNRNywCAbkGlgYGUlSsE4pktaav4S/KVXpWocOkiGDh34ik6+vWfK
ZG/eNh/ISMsjZeLa+n+bYfARg7YdpODCvvtiVbQTbQ+wLzuEQ10PrFG8+ccdne23F9mku0V5glpx
JZwFkYzHdpC3jZN9hvnhYy8RAmzfLKiCT8x6iInAOdJRBHj9jtSSk4zY7tVtYac0sTgX/RxH0LM7
gpLCbVxtHXGqzAodNhPDWhiDAiyDbhmR+BmBr99Fgq1/viEvmNnf07403k3jLinuCWtNcX2coMEH
+/hwAoFxS7zg93zUHYevMrwJwE/+0+SrLxJ0BJfjx08fh6cNVefUwHrsTwpBxp++hKVo1LUWQB0V
1GWpnNBMl/r3DpGFQPe62W8dmdDu5b/xu3Ma0fWyrqWthyBIH4OszW0F2QCc8XiOrOZdBmuJxu6G
pyX5LZa4z9uT67ZJphkiGG7s8BSuJYlMMBn2qITypm2mzoIlZl0uiBaWBNSnLndjdo5u2MqMxfqR
5WP35hYVaRC1KUKq8Wsf3nljZrKNlqD+2UFp6zHlA74tVDat87GduHbvQHS+Z7Tsi/UW4jPH+8eU
TSkWTmzm5HldstVoVpc6PgoO69si/RP0q1n5seSp/q/6uWWlNhmCOtLI53gmNfLTws6/jWi5nR42
03vC9dxOrOJFGwD8P0PMwUPs3vHX04YmsiJWKQiaPVQDIxlY+CZjxocvshvo6zVCIsn5FXtZNdD9
W2xIzxTc8wi5A8RL5pudlJCUcW3zT7MgCc/g3WKJ0VfdyoXD8U8Ycku08DvVAS2OxCgMRGweY05j
kFwkw5I+mlcl4is2XvktO5pJgyoQ4mQbNyx9azU20D0YplzbPP2D1DXk0/GWwqjpR73TN65lwlhu
fqyle1Rm37A3kbmwzdSWp0mGuVRRKWrW+S8/ViLd6aaxi0aY9lCVTfQWb0BECYdaTqSIiPHBdDmB
2hJkVNndJtuBf5reWFmeRAiL2itwlvybgUaGNkZBeLOl9GoCeDArvQl3R5LB1G9E8ChrcEDApuoP
UrVdi9Khsfq+x8MzHs9rxhcXaIA2LxDy8doj/8AEx5rnLWJZtrAytuFPVQRcqQz/Pmh3d/NNdGFb
y7PFVzNKl7mLsucZwcgdl+fMs0gKSbN8qS0vdHn44BVEV7/Io7qJKY3WNPHToUU/cjshX6XvTbDY
nCWfPBEx5e+FhAg4yFFskHcO/6hrIfjAlodIJJSHsnMCxSg3z5im1tHf3eoKZ9GK09OwdPBwFbDz
nTrRjlRdRRJZ+rIwRyjm6uWCwZ4ezUX3X/HfQDCceaKzqUH6OJmHhBa2eysW1QVtBxVBcpW9qkwP
A8tIJ5VZIUgLsrQlG5KhDx7+hym7R6koRj8DNSLjtHNM4eMI8e0Bbpq3dEbMinMKde5cnc9k5f2U
9YMt4Zo0K2ahUyV5DQO4OrkhnyPdW/Qw7QEoomZNDchJa2EONBX6e8LEukYI3N7+4MZLz1Ep4K+z
33fuiLoeQ5kGly7hzG2ivdc7ilWGfXKy9ulDDrRnyLTjsHwkcEw2lr2M3GAXQlAsfAuVkpbxZdoO
bLzX8L7OkwsDcSVXQXjGXtNOPytVSimNrxgocMPQA7DRVSEBiCu1m/XaXIBrCvouxHHzj9QHfzwp
c8xENZiHcc5TR4pi6vRy0axRyMLNysMQjKGUYpBM3TYfSNaR3+4LQ3BfZhzNkQ3BwocZsY2EbQMn
IkGPbMMCV6dXCxROZ4X/BrE90lj2ZCe+PpAB7YRU/7VtKS5qXsspvpKc/PI7ceGBtnU73sVPXebo
HNiZ6tTe5FA4VYhiUForfxydxK8PlZEmgyrlGQGKwaq0xGArkN7rgVSEjFeEbM8MQjZBETbUiBmE
8T48n6JqXZ6a0gmiT4nwi2CEmsKK7eIT6yGs/iQh20mXOa1Nya5VmWZpfojNZlrIk8mDbtsJvsa0
KoX3tkViwHQKQoDuJ5KTzz1UXGUl5OP4OPpYRhB6ZFAb27zglayi/SfhRQ3TuQCL8BdJQ8ElWHGJ
Lz8aMX/rmAi4Ogj9ZHnhdRy1rWSrsGxOwTbP9ujWkViBoxMSZC3TRigr2CUvY5obmqPUXnVDzatI
hGSAdQrqJV58XNMeTd6Z35FA2Qht8STrxb/UEyhPXuV+5Rxb/Zh8VGkySiD1QQ4b+IpA1aXX1MQV
xPgbyh+yWBI7YQmLQ7P/3f8gcSYqHiPC6YvfFeWYsqe1RvtJATFSNfMQTddLc1nqR1GQt7xN44VQ
AeGkdeaEnBzn/mhLY8zgkhLdOfHffCYt2CGQ5kfgVU1mAxplZILqSqyhLJ3zSnr9zcZKDxdSaoyo
Qp4HjSiajjPnB2/y0Da45b7+EzU2gmcpO4IYUqYnk2liXDrV8KgpL80AThP2Uy2iuGQHIFBb0+FY
yJhS/TR/zsw1jXSDiEmkFi3hT2wb/zx+fzrOk3flPkxi1MKLgFM22GWh6PpNLZr+Zk0s4TQZ1AdV
rXWz85Or5rhLHKaB5QBTMNz/HuUcusDnQGXzaRoLzD30RvfqenmtdEoTTV4IlpbeYUPjiskFE04u
fD9CN8HD8NIpSGPDectr62Np7ww6XSztiiGWTiHLWEdkqhKZz1HyqR8PSomr06fBVp5Wa8ZJ57fV
rojN9ybAsbI/dl1lHe/9qPSaj2XdBRDPebwSP2d01Zhwj+67rB34VzXNM4U4/UzqThZ3ztobh06F
SNI1Y6ET8iaSZMt89f8AszhP6ee4mTpAf2/pwTTfY5xtPjX6gb41UClrwMBDUA9Y2jrZWUpmZLIq
wg5VbKZPxGEwio2sTAVAEp+r5oIzNLwspVG4TXrcwsuiV8ubM/uxuca2QZw0uOQt9odpkKha3TZx
ZtOH1Pr7FXSmAaf+4pYWTiMIGy1Dwkb0vqIUygjALJG2U3trDne4ZZ6wzyyQxaJLFy85rGtKR8r0
Nbe7Sfm4ggSggSbb0B0wnnZrlYqrpnvhIGSFekDpP/7EURUuif+59jyiHr8hJBAoROXsJtdNUJ4K
gXPouclM6betTGyz8v/0ig49iSLtNeROwk+ZlIj8UcjNw6Z6Zz7iIzBzzxZm3S1tJ0OxhbEoY2bw
O/2bJNrKR7ys2c6J+1eIkQ7Eob0QK5OFPKr3y9kid1PhJobb9vBGamhXilPKmDDAnRSss+pXSUxO
J1H62PtrGuMG3nbU3dGKkBV9oLQQ9v56QolueSqd2kEB1SRWUrBeulR7F6uy5Tg/Yg8/QsOT/Ufq
EpuOsQWujNY8bzCWJw4bt3i2z5vEH2t4sf4pNF6+epbG+91iQDLHheMZzu+ZoZilUyRpYWgxIJnN
Pjxix8j8Osrmj94HdjX8KhwcEYlobHGxS/GdpT9G+fe8Rw9EyOye7/pXF3FUSLJ/h2wWQinp8EB2
tSauIO8Muy6xxWvSeb5xTaQEeeMsFDZZU+LNA8uF8JOu8QY7+vkIq5vhDlEbiVqQXpouc3O6I2h3
/bTQmsTHYkiaLxNOfaR+KBToa61KzAVcB/Lb6xCE12sTul5UIoExfPfyeJ5F9dqhQ2bCk7DWQtcM
GNfOEn2AS4nvggwKfOkWo3c1tCwELoW1LMzBI/gGJ2XRNXLIXo220uRjwU2z9ZW/JvcotEKL5y+e
GCXQKD/L5U88YmPhoUmC1gDa+VaBHIrV3T6la8XX5KMe86zM8Nf0ZADdMX7nNEUrP+pvBxtWFzyt
BBA/Gl2QWAVcKsEHuiZz+GZBylgEyhw43Ev0tjtr9x9NaMvU2YUuUYqbHzFvr2VNq6Ua51F1z9XS
9UoQOrnykDzBQMfzJrS8zaqEy1KMOg2CV7TTVHHkME5jPRCmUR2vAGarUuzILVZXDii7QK7+qLxd
x5KVbZYz79oda0Nj8Xhl5P7DIaomQcbnAm45KQRA9WqdidVBtTOAUHIAwA02dsikR6qU8LaJPfz6
idloNlZDQUYZWf1/HBsBCaojdT7zZiaDbtZrznEQN6jNfWXD+yLYhJORj7K0A9GWqBFPgS3RU63Z
p1m41IMAhle58OSj5y4nEij+cVA/61HiadUlJqc6uj07AHgQ4gPEOSepMiPNUEJ89JzcveNi0HRM
FGCNoNHPN6+aY12MCifrxDV/5GqcEXVvT3jDShf4Dlo8SYLRXF8LN1hmu9QOsSmeZPKCQHcc5uAk
6N54mNaj+S8dta7z4azwWV6w/oNu6y7Q9E7pM7kpG/or/gWPEdWehiUTx1pZ+gVqxfvw1groE2YU
SrwdIkFfcqeoRA7BAMRqEwL1TJ5QdeXZwV04p4ouVQ9tPRfQJq3yWaOC5CvRAparZXO58xWWMyja
RdsfKC5MEbmVdPLDR+TeBaBODha89MvOONIrZL/Co7U88L9a8X7VcU4vndkcJDsNhVwNSwMpqn97
PmErhVirLVZOdP1xF79BDekwiKPzVY1TqtteL04uyJtJVxERrQz237XywT2joJjJW7WqwCobyTnp
IeNl9z0P31jq9l2ajUt+XrCXcIy/ph/W8ao0oqoGL5BlDEKrgoSxhzJD2A8idloz9H5q1CAcR2js
/w6W+YrMBXp4bcv2v3JPZvW0xCEMeypFeyIk9Wwd0NijoonhLNXG47Z7MeijtPH19ta+TTxJb4GG
9JBRPe9AfnySgDPwH2aKmNeS3VAjnWtMNj1MUbYkk8Xk+caRbuZIiniRzYaaBODhVGN2UgBHOTh3
heItS7byW56FrR8Ap1f1WJY6f255RQma8CXA0tqdLndOIM7qobganhEgBzXWYeg0whGoS5arQN9y
Ttg9z4uUIyLr8frsiAjoTWe9NA8P4DnzjHWN7o9UXAldR3wXFu+w3UHmXKiRMW7amj1OAWQnJkRi
xVam38R/jftLrGG+KzytTOLvDLeNNYozWjUk0r3+nWP2yEB5Rt7iSGcxaWsTZhL9cdNfaosFKm0P
SvawPEffUSHO0p75EkI4qjDxDR+c9d+EP1c49PI/8WK+YOQI4ZVhzYqlFZOI2l1QRAZ80M/bv4pU
T5GD4YDuTPdOVcS4X9g1pu9CETq76D/nw7+NZ4AfUgDoSgKzG35j3Mg7rq9bxSZPd4QI9tMgMpr+
VKublgJ0R08xGyWv8naXwnHv9mMRONasq7YLUt+cY9qihci5VP71UVUkZSOi+OtArOLiVNhctuPI
JYGT1EQP4px6zj1gkmBj/ol8TxUsNFezL+mEzU/pmgDjUwSBq2TYhuMG8PZe9F4LOW5hKyeq3zzb
xPIsE9DBQbPeH5p7QQmuDtXFYlQMvfRD/jbTH00ti1AhxKmDOUbUHWgfPt9tfRsbBlPjeyhUcteX
maXiDlREZrhGi1PFM2jFcx0miPEisd4I4vcFsd3oPbxaa+3tlBfEworDV5ai+Ts9j6pb7+8/1wuI
sZlnvaKcpem6+cdEtM3o4P3+OKQg/pcIzAIKX8zfJURSIF6QZ9+FUkEZJLqiEvRU91JKkQMCAzLz
d2rzwxRG2nNz/YFT43lw0m0OMNwF4Y1rcWqEneQuhsDggN2P26KF3FX2HE5CWUZQh9I7n/CnNRO8
Ml1C/6OyjfmpLerk0Q5pC0uYaD47iv0GAvcg/SXQtU/XGJ2S2YqPWlL4hBMmnTU9DrnfERBxzXAW
MSctX5rS10Kiy+fu9jz03d/ExRB+hnC5gRCeMmM8ZFzdISDTmpAbwPivqoWzde/6JQRN86Iw8loX
gu4m8SreZWsSfkzNvT89H2ednk6acZLSFw/ZdoIBddcjJUveF0AzFG8qBTlL09DD0N8QVKycU/vP
sN9GSC1jkgJvBxhmKuEbeLDyRV+aL6aWvG1f20yp3iCmDvFQI5xbVVKGFqmOgiYzp2lXs8Vxa4xM
ckkSbfpYGPtrWABtAaKTXV1dUWzfQUwdVg0L5m+vwX/oiObDvdY31CwfTsZiypOat0Beq3AK7fGF
Qj5Z54obmccUdxXHxIhFqv3jK4ceGEcmvVaxf6sF4wfoDYshUNuketHKk2oi1bKiwZNxogyHERGM
8xNK2YA59CT8u8ONep4j3YKdorTzKp81abKIzyfcr+qEPmCCRhzfMe+X+m3s8KWONesStS2l71ay
BmhAW+RshhY0r/WQyKiNbrZ4/gWKOSjBXQWgOgJh2X/tTcdA7LYE18sJy62gHLbs+tW8s4FKXma9
SUv1/zoTXQ29r/KTq06KndvN/LdN11QQN6Qb77MhXRv098pHe7RIBjDrvpLG+3Bhe51aoKrHiwNY
nm9B6AUJFDrmWB9HtWXbElvRF1QUdV6jtf6uZ4PqJZGdVDqIK6t8l0Cz8VHR+iid5P4Nj7LogKdb
am1fbA2yJYHynAob4V8Yc/XLOO9Oyy8WQKPIXiNJnikKn2ulqu/mG4wejNAcR1w8gCcfCM5XAM5V
uGSWVqXasYmfsnGae/j9yOIBZ+p36VvQYOafNLiqP6pmWx5d3lHa4r/eZfvh4MuCmOirjkkTkEPU
kgMLUeJNVnOCx2NMkQrjW1J8j4xhR75F4L72fIiUP2ozZWFDJTfMrNhv3ZMXf3wenupLEnJjLEot
xxJIjfEAqIJSiZPPgyUfyZDrQKMWWmQVS4IlJaJ2ymTiogSd3LcsGeh0Tk2Ef/zGKedJkIK5Xp4A
n0HFL+HHXUb88yL7d7Q98sR7cEZ6kFFgL0LyOgm9VxvKx9+Cut0/VfqvovizYD13Z03DRXtRHbGJ
gk2kx9ItWTav8f4MgnwbN7A33l1MIVRjpr/JYQ5iBcuGTM5c6phZJBBVKIsB8c1lefQcI7cn6St/
hxvkkrq7Buo41bh33ie9dmyo5jo2dGx5Gb+HlQp8X1z2oeSeu6Y1df81LhzDVmyWDZ99XLGvGqCi
Kgm+Qt5XYGLMYkXjDCOVBk1os4Ln5QZE5a5yl8DFrmOfUYAxdZej86pGnpxOByKGvL1Keh3WRMyz
wpgVCm/XZgdfDyYIJBUxO/abkn4xecNfu7xOzaK7uVbP9DNiUEu4ddAOYLoic3aON0BTA5vDwlX0
bWT+ncfAq5lc0jGJmm4p9MroneNuXvxJtZ63oRfMV6ytUTi/joqD/AiA9ZpEZz8pqTki0svloX6o
mpKCHLVjbsP2NSzPSz1CPGLU1wett4P35HUMMFfz/C4qPjWLYH184u427SOypThej/Ga4fpA5XEN
YfuLjEtKjGdGFjVoUZ1vcCerhk8Dmv4LZZ2hLCHBGo2GGriPw25aefVGLU2e9HImUnFhZEwwQKbA
3nnCefE3kAnYDn0ep4r2Vn/B5/5RPIYVFWntNhYs3yvIhjYFa9+kYaIOzXQvTj4DcM69KDtiU4xf
qSHx3ucNpP5gQAO0oe1Wgkj62bh6toBEYGzh4yxMKePtEtYD8Htg+axhv4QszMXK8cB1hHM1dnmt
yZEzGFhzrpPqEps1qJnfwtAHsfv8g0omVyNnkW1I81i3L1KaaQPF4OeUu61/YP9ykDtTrTdO7k7R
cPXanQppNzwvcSEyKKbJyQHyIl/A6gPqzPaNOZL7XM77HF5eH/zQ4ujxJ9SxO3pN7UBmCOygtn7r
BLzSu4DIDe2WyyT9QWJGDxJw0G67xyDaz18v1w8wViHd6GwBZYMETaBBsn8FJlc70kI+QqEta6nP
1aHd3tcSCph594KpLul65U6WgLgpbyJ2KxR6DIU+MbWkds4c5GJomccUEkdPHLq9gx9waubtmWQZ
v1NvZ4AIQmqr4ESZa3Yb4jNY7H1127ltQTjOZ+VrKUZzowR2jkFL36dCHincGLczYyDem246Qglu
S/FqCq/R86vklfvzCSt6xC0QVysX/F8nRAAJi4L0fga6TE0iHh6JXCuzsBd9meCYXtULS6EC0WBj
aasnhak2PeDtvqtQ8+MnWZaHusmJENHjyZdXITER5Yu7l1fh7R7OlIAuvDdFQuw3sTT4Hb3lh1z3
OrLBMPLfA+okF7ozGl2Li2rOVqJ/loCrxhdnx3Ywg5+DlFvXh/VGLJbgWC1UzeQ3bTpYlCm6K/SL
jMrZTyMJK8o5Sbf10hjM/vPLAeUy6F5mqiCTXSq5SBfmzRFKG30jwgjHLfjFpv3ZdOmyCrc1ZgnQ
xKJHHVcjcBdPSgUtzHm/z4q9LGWeF6m5bXm3sOvBkMODekAInOFbzsLp1IviYMjqx3qn4AfWuvOx
bfCIrqfc08JdcYAObIhsFphrYaH5i/jaHTUJEivs16CAseCUJYVxWbcNrp2AQz92A0vUHfRwaLmX
Vx2IuvRWC1Ls9flZOAamuRHiPeAOcDsj8okhsJm/30e7LCvkifONwESZywZB7igU3DQVGdzalWVS
PyVsLo8q4rnDvC0JurMzYpLuoiT2pTap1RTQADGA/12DSjuyRV32+3Qmb4C3jKbsHsm3h/rkDCfw
x1GZCwFgvMG5FMUqv5Dmnpnp5kqUC51qvzRKGuKP4cDC6s9Nk49KKgNLobDEb612LWwg63HuZAiH
5wju/DxJ6/VIdh05l6WGCGRuyj+3APM0OFRL3LjJeM99bw1kRb2AccNM+FFTUrEYJeatWgDatm2D
mH4L7LRVD4HYZyUW07bo96aRSkN6DDDHSQxaiPvvMKauuP3mGRTwlsicJZEfjAOv+hneTaLKtnZm
wM19fhXCu4uR6SnXRFo2VzLS1gCnelM6cmFJjq5bL3o02DkAibDvYO7LPgFlU+b8knP0Z+dxaT0i
aWG96EPn/YrkRHuUzG3ekrtnLRwC1Iv2Xc3VHjBzVn5GHbNmsBCyx2ndJU3Waa1Y2z1Nz3HfiihV
l/MtSSWWqWqZWKP5+KbtBy+Nqikmkj8MBtWwDwAvVT1dJpR1VOzAv1ibC3mlOqwxrBz4PZmTwxvP
NGb5P1Nzf4FfNDtlawO1x9hYBfnvgr8h03jy3R1CIab9nrUwHHi5Yb02FYBB6d4MsNHY2VeGMody
u1pPRkkyjbbfUVEf+vkgHXztBlvhXVXdsrfDO42neoOux0xi/dzMKEgSBdDWPKz40sNUNVxkwyps
A4UvS3Uqs3peA49W1RpZVP4QVXyrO5kabbIWTeIwOevzyjnXOdTVM2QZrB72GL39jieU8x3OBhy1
TLLFF0HIR9uqMe825xqy7XtmQai2odLV9T9pHAMwe7sRBFYLsERunE20pWixqFgJ1R0sTYguAKb8
2zNc6qm7//puxrMuXGii7bILsJyMekFR/KBY3glZwUH1hr6DrTBENh6DeSdvgJSLDvJyqSak+N0B
36mWHLF/nqp3+saQGIdW6tpWdnMWIWKvpnnx3Hy+8fqDGVYYu8eW2U319vLx9FZ2dEVfsV+3R6zw
x6OSfpBLU7LXUjYhGukX+27VleAEKgcgJJkFIJRvn09KF6s01dEpFysFqSGo6K3akfxgWf6NcmfT
uR6ZBP+yuhcm4B8bIWUfzDn+mS91XifpOMib70QuHwGo0JKmEPo4b7AnmtKy171sL8sBsfvRemL8
MH55ag0i/EYrhoozkJPYL4bRG+swy4obIEewtw9juQDuLeYjWd4U1m5IrDvAg7bA22s8umyoggGW
I2a1QLrHWb21Fb0PPg4Lxfq/zgVsw7e/Ze5fZus7cBp1ojrTcVbFPfrU60qb10u453XrvMrjeUdS
iHWkw0h0BqqEaNNLxt+df7UqQhMz1KPKKGgyiAbEGioPv4hjFLaG+u3cJt4r2XkGUdu2fxiLbgO/
IWsXcXGoWcqWY0JzR0w5Q90CLTcS89CBOXTeqNvc4D6O2ZK8bNFABB+nNbYBN4ZR9b4N/dRTwh6k
UUSoesJQe4lJo74H5gI+KkVzJHReJP+uGcctVGupFvXiB05njRc+/jaNTuUBK7l2tcI40pM2yOGj
v/smf95h50fasf5U7msM5pm7KH7UamfLkS8brTcyBYFt2trP0BeZh3F+L6fKIgavyR0olYOVZD9+
FWIpzC/mFA7EDbse2OW1OVAwAPsJlKq0Jzor+AMOOZsEjr0/qXNI8683xNqPaEW6okgRES261Rmq
+vv6+XwRKWdKc7zX+peUPTT1W0Wd646tJNXSol/NTMOliV7OF4Js16VXQTkZ3LY1w+Uzy6g0tn+1
tH2LX2OO3p8HqNX31SB74lD7lFyU5E7qotPCaSi+oSK4KgtWPx6KinrubxV0KS4ymmgk7YAi4LUm
dtOpwHL99M9WEvp7dTAQs/M+8rNtZTbqPHZsAMEAqFZFzNK8cojSvayaFZ3imviJzmijjVsmDMhV
k1xzHxaL+YIRknNIGT01yfKKQbouyRodpaClH33g44bzAfC8gurbUlXQfxRh0Voo2fR0sqOdyY96
6Frjzh6+EIPXo72+fpA4GohJCix6m7edSaecfO3pzGiXR97ohoHnNGWxgN0UzovIS71FPlAnoiGj
amJIbl7NskoTWsI2jH7WnlIhzmn7/FRx3Ufp8mF1zZdQNA5sO5ypv0XDFhf4gZCIcFHycEnEFVmL
tLtVxVfQIDoCnZ4v732fJUz2B7KE5eCf0eOuHJURxflqyeQSfMNirVFQXgkk1E1HU85W+m8GbkWY
rtMUIaqKuUbmDC6obb2jJNOJGyIXOB+DQyc0RH1JDwEL6/4wHD5cI9YiOp2rgA9wWGzY/8luOv9z
oPsTYR9ahhsPXftYrRMjo5jGQhT5qk35fCIxw7HlCiuuw6ebFDDhRLkVsH3WDkua5cYMgsi3vM5J
AFNp+dYToHdAUM3Gu7X6oKghDeuLoIMNIV0shmGuuxCtEhgz0FOvxVv8vpvNTl/d+pbHoK7IY8is
7kj0raJpx9pXeUjCZYytFd+hk43qZDOAnhbCsxmN3hY4tHJrblqnoizKqLOUCOGy3+92IrRWr9O5
4fKgAzL8XqU3KLGVP7lW499CEx5eOPe2zWHimQLj4jmZMJ4KpYm+ZWz02e4FOcYqd7g2ITmRjzYL
Krzhn9Uh8iUnLW6K96dabI5EA4sa73wOYxB+vH6pZ8tgppPam81hOr2xVL4CsEHHZ4Z3jtdvyVtO
wEbNSZKJ6P1srhHUl1OTwqin0+fWMl0DUNrzYMbSIc2z07yoeGkeMzae9NgqO0Ff/Lr+QATra82X
goKdlW+ZEiHC2Chtz0b77zL4WPcLBLb4z9c5+2pMd4u+B1MdJ4ZeqwmDakC3e9VwnRByPKOdWYf1
NNUfetdlHs2xaY9DOH+/2pAzfgCTUEArTy60lOfiMXS21EX0ujuPvqFR/sa7mC+GHoZPkplvK2E2
7NZ8i5AvyAO1DOM9FCDkHpoH9nDKbotlkKiHQa5txmvuKzfRsCEGlx/g1REcP4WXX/mz/ZGL/jeK
6waWOzyPnSe31b46UOlp5RuglRYjoG/1gPzkX6vjRQ/VVNrk6MaBIlk0CG7OOiILNvLaZlfnNp5D
WlYRW1QGZ2/UQJI3dDAxCjddFYJ4O75vCAOwmHt61kl8B8TrT7UgoEb2mhYJM/xpcFptD8Uh6AHV
0oo4mgb2xhngw/fIOM9M/aFNLdgkgFm6rU92IqX5Zq5WK13m5kzUPDhqnsrLAMxjGNTL/JeEoMrC
Z6c/9+HCA1HTd85oViCexTWonUY+wofmE2znFk6atIYpvvjlYDAT7KjrqE/8GSTrVQs9ziAXyR9z
N/lSkjl0Sa++4/WUr5DjZQKVbsG5jewCRLKkPCSm3HiRoQgoEELItwuxBJLKipdBX/OVecUuNFnm
a1GUks1HsedTYEes3R8My+jmnnzs0HHpll5MZazhGvYWDo5BlOjq9/90nUSOrzkAqzL2XZ4wqPRQ
qqmTpYg9CmrcPo2evaYfvtgvz3bvjLG9U1MEyWBtRwWoaVq0m4051dDlPN6ewUSWvgnmGIsm7ImC
iDpCl6cEwxn7tEgS65L3QDktvpXKUFtYR316zdiR934vNdaJlTE4n9URfWxxEUFsvF4GwFxjmSBL
Kd/FxMSti26ayVhdDp4YmiwXVH0eoV9klLjQbnrPEUEqOajNcbCUAMexiO6Kt/f28zBvVrg1N+pW
jlojjZosEk8QDdcpMYwqX4WvmJDxPj2kalQl4C7b3Kx4KYuVkpy35pydliLzb8M0TBMMZx4fiw9z
QKvluBbr5HSU1gSPHPDtSkuNtTaCSg/516uudVq7PzcTw9D0RUTVgjGXNC48ZPGQx/XAoXX2e1QA
4ttgcKVyMgAuZ1gjNVYJXbAikNa4U0561qyJRqMMuJDdssz3HLfpJsVIDq46ag96KYMdvqwQXGpG
dC9O5x3zDz+g2aior2oeM9z+VHZIFRyMMLKyqMg2tMpZNN3Wz09jrLYfV+ISo4v4NN0gIwWwJcvh
2PGQuTJ9L8Y+CmAjY6Gk0ALlUCEx7xDkExGcbTqWX2XirvKVwAsN3w0m5U+Z1gyv46mWYro/QqoJ
LuvpBpJlMitWRSy7LskEmes344gAo/R0/LBBnCWOWj/9bC6D/oWIhYCKR93r+xSEvzVhGOuaUAja
ya21/9BRSfMNZdspC1Axls3rHPMgoyJHiLkCJZxTkgSgm1QL/5otCgceetwLc23RomUjQtq0D3lU
2Xm3tgCNfhicVVWZSbBcaIeAiAw/yfdeJrMlI3k0cw6YyE2JL9dJWEIGxzqbA1BTPOMtDdlun/yy
keIflYke8Nsj+N76YUwOra6XvdiSsGnCtmEv2V0D/+0asLRbqaaLjOkX1sZqKxljyP68ipiQzZOr
BoeII+QjLRpTRAW4IVSuH18GF3Oky0wKVYei0yH2/PEyxviIFDXgm03scKLjJrVrE6DMJ3TmwECF
AEKVVogI21qaeH1Mx+mIt+uE8F0frKiGNvvbFa//6PmBJ0XRi8SLOU1BzaOwz2g/dr9JI1g4s5AN
0z5XDUptXH3t5rq3V0evH0AQrn+U2ZglN57F3evems5H4VpCx5z+xnL86v/sNC2hBPWxPjQBWtMx
OP2tx7WLYg+zpwN4JOet4GyKsvcRZO5rIrwKznQ15D9/hbDd5/AifWgDhFleMOLo0FqGa94oXD0G
dDVFIjvaO6oVlnQVVfrdw4y7Qd+14h4jmJKJrptsIoFXYZS2yz+jQEl48lQfbRUoJR15dqr+rFIS
VWL4mgRXdn5c0JFVi6AAxuak1aTrhDUWvRHLcav4VXRkrALMisgnPhlKNUQQVrQpYxQRDkMqH2l+
3HyN41ee82cB/k17B6SRS12IB7eGmDMdA7NPaeLLbqXBUZ4jdAZYEMoAVLsbZx7iNF+DWQpy5c4t
O9QZ5JHloz3mpVRmX8NJ4cSrtoxkCOId3g3e17R1VoqsNWRVzIFoKC95fwM93qeEaFsM56d+INam
aUlvRVCNEgxs/fGJyjjs6tGRNYQAgQHVZyI7qdCoXXgtjZ+zl5AkNyrMknrhOPc6DFbc+hjuzBdN
k0sB3xlqS9w5ligC0QVtGUEtCEsFZhcE0fmbmXQ86cmNka8UzO/KZrBbDt1eSU5JmpWkyJSaASsO
yF4CpPOQ8oBqK5YtjmY9Ji8J55+4xtxVhrknJQs54PKk2yJVgCRy6yk+6DaTnc1g2tjqlFfGCRKn
Or2WpE2nAwgmjMfOlEQHd8/Oss8rwfuRkopk9KSChO3Ap+zLDTcWsLaCvSd+7bPxJDej+zcDW37u
6SfMm6a8Ag9j1eud7mV2sNSvjZCfBYdmgA+bD2Bh5yM85UikZH2m2JWnH3k7Jclf3i09z4FAMWvj
AdZI3qtwlBks7m0r2am8JUp/HUCp4OZR70w+ghTyxLEM4C2iHkSdxdXpGCRhi8pl+OlkTRuKSECv
5x+IcoGzw2b4E9zaThiHdoXLzrCUFvVlgZ9qIKZwUoha2pEO/sK2s3KKyt3sDDVr2VY8tGTPT8hV
nbgQ2Ev7kd38H7rXm/qrR1+3NfvshF6fSmItiJkf/cnM3JIQBes9aQrT3BFER4SDbeuUWvZT0oGI
XGjMRAII+BlRV7aTybinT/y1PzOuiLYjVi5jF76NUE1voKXdPAEps3cHv/ljCHzHp6617aSfKNdP
eS9ZGH+QN8XDfzv4MvKDBeYB5J61rWnWBMgfygWi1prpq5DocpuM0Lp4enE5ODmlxD1A/8hRLe1e
RWB0YXQPcLwfQtIK1d1RvFtKp8utQ7OoPM0k0NV/R0kpp8PoDL+9C0xXOMjYTHFAaBQhWsM8a9Qs
kG5BAQafAna1cJaVOxn4yMrImXPyKiQk8iVQ90XXvvCg5vVGbUaL29MiWiqKwTR/oUlXFW5jzwMM
lfjfUXCokXoLdfNsCPCfP70Dlp6ToCsxRpSfiJFTpKnLW2092jWcANb8PTzZT9L3SCy8KqgYSfYt
9jo1TKAGPSJgXioLKN4e+9jPc1Kdad3rdN51xuqREa38GkRKJ+JawdBUIhRBE1sljEGv6wqACcoC
CxJDWSd66rFAvce++DXAiQ+0jk4o/NboqPW+BUTNEzmlLWN9DdUklxNRknIanQRDo6aQpD8LygZI
SLi/xmNbSJrLukIjo4m+yX7aSl6GQANf0Ff6Ux21KBLeKpQfkgBeHo65Mvi4drhUtkSDOydQEnQQ
n2zA/GAzQ508sfXK0Qrrol1o+Wm8MGi6gemBBLE5Ro+AowMVcUjZkAmuLMB8vGaLo+Sw0g3uvhl0
Y8jK1gM+eyCi3Ppl1PWlw13BK32W4yWdYe5CrOX4ZShBH34l+h74/4LQRnRyJxsGWjiQ/PAgh8Wq
BQntWL/rN1rrUCqtnARqWADD/DdYsYEZRgcZJff9glL4L8nerHXpHA/CFA5lCUpoSuyw0PfT3Ib1
aWGnO1pzFuuR4vtTslMD8WO4g26gnKZUJeFZqc6B171Ah3S0tSdDk8uwLTc71MoIf8EhsrjqNBLZ
3+gziDSvbZP+xXRDQjm9iRsI87dVaaWdull3EKM7svimjt4dS9g3qfiCEWpmMFzMkuLY0triKQK+
WymNpvx4RvjOxk0lLwP2nbdQvskUssa2Q8voeS4QzNx1xpSIqo7TMJDEeW61A62gELNnk39Y7+qM
fWKOJX0XqfRGZBPwo0xJ+Q6lCplRzdVTpzMRz2BjM8L1lDCKGrBaDjiWf58YQjMpGSWb6prGiFR6
+cNA7+QMMVr15VpFDG188BXRv1ZcJXE41P//+Da3HDFgUjvmWoLouheHbOEGDG1fKR88gKKX7uD4
5xH51JCF27GQV6rs8XnXUdvMHxTfCIpdOEWd2cPNe5lJlCmRXRoIUvt/CikWsALNV6x3Ha0AzuIq
fPGQb6vuqEAbOma33g/YBRzOXstQeZYmJk758UPwQWLfIWZzjM7jXf3R3KjQSbqtDD0qstqnJCnk
iYiA2diF4oOxJ+gdMEI1InSMLKwfYsYatbMIvTPwKA6hbYhpGHLtBMDTXhyC/8T7GhexIMVFEaxw
dogB9F7FGwFMBkG/eV6Ogbvemqe6J2T5goNPS05cxzXUXKBqdbsbdjah5ydGJrNJl4UGbvBOpx8B
gBP/FWQlLaUtZsB+JorKgHijJ7GVm/QcY44nXrw9FAM1J3zFqcXCwd4rrHx3IlSdJuoGh5iilkSd
CuBIM6fHOgezLn8T7pPWfzSe1EczBkQK4buqNY0GjnVRQEuFS0Mn+4x79WGBj+TKbcPbCKJwEMa/
+3RrHVSl7z59PjFnlUvLJ0ZVUzBB1rpZ0ElvaE4NgdcoZv8eYFpxofp0o3uPBT3yLD0r/uQ1/8xg
rL45xcNKPAdagyEqiLRaG8RQdhLFzh1cr8gxIe+k7Vxs86DRdsJQjGYlutXBvxWjhIuGcYRLmaCr
t038m5tNT5p3ZZVYf5iS6dCUycF8zu6AQ13MRqFCO9B9DoXMdOYCrJJRk/x1QACU761GI0FgcXuI
N4Cd7RTcjcJ970zMMLWw+/yytXuHrcG10qw+wipk5u0Ec7onGLuLVED0pImi7DkzcD2UkKOQ/9Tt
1uj8f72jHwGvMA2rdeK+CuuIqPeXm6565PhocPCw7IjdO+CPovutVFEXqufGUXcIIJXIngsfOZ+n
8o6dFqnX9FYY63Bojf4JiGDr9OX26ySjIgY3spJ8ewlSkI5ImJJpD/b0nhs9nOPdTiFOU5RXU6yw
SP84pFZplP5aScGQgRmEQUOVE43AR1a/vlB5MoLskacBaN9wRZR95cTRpyvgmE1joQXu0HJFctGW
ynTuH6+DIsVpcT7bFJUnawMkcjaUjOy5Map9bdb475927UkYVY1lfQwa9WOFOY9Q9hST3BIM3lJH
uoRPJEpzEVMY8BEeOWw6kDzxrGr9mj+gYJhqvmHgwWCr1+PmWVylaRbCPd+6oqWVIInvYendsIal
Yn4yC1Lgl43z3hVnpDcWIc0GwpLhU1xjwT4fA0zv8l5m5hVsz0I/Hm4Hj6K+/MqrzEPgQagSbb4j
PzxEKFkXKu9C3r1/47qcmtOqmAEV+Sft9vf7UjEsTfL/KLQ3LreV1GbQNLnU6/a7u+eXZfVpbc+h
CmaBFPMM/CPP8AEODlgTF+2cT7vaksw/A9vxAP9nXPX5xnl+FGy3umAhINfwvouGelMDCbOOpQO/
MdB1EazL4Hi/uYkHnQtKEtjzxGpCfsKc1NtXTg9HkkWaHQVhvJom7oTJVEs+KkqSeD43OyLyZ6iS
xMRwaSRvuIrlHeSxEAAKRNrI11axATl2dnPnQO2jZtE8+vI1px97e+QorFpOa+8B5OkrjW71Y3Xf
T4ofGxlGMsxwuJ2AAn0z+UA3ZeUOfv5aKDT6aZdrHtP34irGsguJvLEvrL2GWiMhN77DQZqxLL+4
MBVn4xjQD4shx5jS13FXzU+FTdXrHqAkSnJ3C4y+ce1G1Ivlq82F7j6waFEuXVB0eO54gM0nbluY
lVQvUxtNRavFFk+nUDOC7TQQUZ9A8s93x3ojxKWD8l0MLBdedfdve//xxGtYzWiN34gbjwcYfGcq
B3KTNqTTZFVD1ym9WiHBuohim439gT4UqxeNhwtWNDS7Q/tpu8QViciL7uTlL3x16iC2t0602+I6
HhpnNP8C+KCOz1n/Y7hqX9O3oI6/aOps/psiky9ypdOzAMkNKphy2xjrHtRbOawQtxbd5XzYsEYK
9Rm4j+ThXcfCRmpP0OGBrs9kb4ESvr6KuVcd39pWb5Yr0rN2Mo4QOJ697QjyKzWOref0Aqx6/nZD
Ozasp8Ho039yPWDnaKNDVOep+wlZ8R3ndDWQnhQqS4IwGvtwAdYDwdiGWZf1oWaC2p02pmC6EB6L
qDf1RMZWTmGArsCJpf5YCyxU6kQyY7SuSFjJv8LtQXeuKcBJaMlGzWmc62e8aGLRnpAQL1H5Aw8a
GHfh+tXuyci0Awe6RWPxNuyKl3i7OgTXKpbDzUyTdEhrGDK3HF32zPO1DVLWgVNk8Q+pd5WOuHWH
/23M8y5/9d/1nh1fs4mNMUofMOhZOdFjznEgylvh4O9JXZVxHXWlGjNCI1qdRbbHGZ4BjFmqVnN4
juvxUKh7K/Iie2+VZWbzWs3r6GdIe1+Co9B5XCvWmc1B9sDI3bcmucGVofcn+6NPk5wLNyrQWo/I
h+oV+NwdFH5oMH/Gb7hp0R8v2+l7+aQKnPj2ZcPH8mLKY3vOI70xJFOyudfhuGjBFiuBR2/pg2Pg
D1+a4ouyrtRboNL+Ls2SxmaPKBV9ZNkjrbYmCnr6WnxD23KlyPxJadew5XCeD0OjkCf5mwhy2JOH
psxrnWyw5CTeHdLEfFwhIQcfBBNxQypcFbABDNcO0eMkzPQFsjnk2g2OacOAMA/wtftK5YXOVzHH
mjXgxqa1cDaezXIYbbLVXr5S4uLJapy6GElyT/Fg3+gTQyo8r89HIe9Od4/OiEpWFX+jq/fYAnSV
G8Cx6f5npoLQFXhyQE4LsskaDvc8vGUuOrVZR8Dfl1uRUAGLBHB9wc+RpV9xRJizahJ1zHPtaE0d
cdV9UL1Bx6wqbve7tbSS4dTshY+ouK6oxzmUqH1s0IfJ9B/GpU0S5wwRN/t9g+0+XYcekrPzTSdy
Quz9fgesO7UGRnY1JLXAswEehcs8VdY1AL/943SFdBtsziaevZlRLM4R17tz41QYkO0hg5gFT+TV
aDZRcT0pr41bwFaF2IS/VJH/gjWBkkev0diYiglEYQ9dvbXsx/B9CZpVaBtxH7YfvqnpIQAXTdCY
6magpfbmRVNpK8AP8Cm+1hqXvYlu+TgAwqdlIFCOFrDAZ0kPcWDLJGlFhsA18DrwNZ+p2K7Waf+8
G4p5TaL3j+fxKEla9Rh5Gu8hxUpIA7VM6qfB1X3wUOlPxVSwfnTOUrwaLRk/p8AVcx2dqXPDWv2G
+3Qad6qrcKcUXU6wm75Em/5CLhO0xQJEkU3zhJMIzBzP6rjd002WvDFbZk4y5hOSZmCX9+pzzJ6E
b2UzxiHgV/dtYsh9SFyQoWODmULvmX4DYXwZ5jG4GDPV7LAWnj3g19G1nm+ewwRjDThNNDmnThfJ
bNN01qb5WVXuYjkg7LxZGA+Y6J+r8Su/80Apgv6iEgoOO3oTanJnRwOtcoZJxiyzWM7hw2fwquF5
iww4R5ZAzi0QL3DM112xBTJiUR4xcRTd++hXM9gLz9qY78J4XXC0f++4Znsm2lZlP81xoRKta1E9
7+m7DQBSeIVrNtVXCggzuzRKrW3nSwJz22RW1cPxrhOF6AtePcZyfQgv34ixmIsHf1DD5kRGA8bu
yT1EHzj9F9QeWgMPbvb8ofLh18wv8L5JjWXmfiM3wfV/j2gRsGkhmBbBmNsGucSmQlh+GcgEoN4R
UWw7lA38bvTrB7+PDxsSRNDgaTO3lzDQyxBWDV8RsfjRuGmoe0+b9ioSO0J2bP/GR36DGdHyuFMv
/WhCE289XmN5uZo3Ix9ZUs7hdf3yBhpb9Y7zpmNrVB0H5OwVuWWw4BBqEnRqfD96TnkLwnU4fts1
z6ZrZLMye1jFm1YWU26qHxZXZNG5u/dgIcOpA0JHxI5X3wE7URcFfxjHb4ff/RukWL0MwTKWiFYK
jNphcfbDuKUp9mqzqFDqnCHUy8WhESF7U7iOVxJo88gVFDYJwJ7/kKAOoI1kSfoQd+7ADT1NP7Dm
O6bXUIZonmFQ9UnoHweTLbwjivHo3oJ7BxsaaKXUxp+dRdVlWTE3qJc8oW47cnDy6JblJGG4XCaU
LKmaULhnFhklyf3vrgQtcBLhoBZ/Rw6nk8oklXedokdeyrxMXKcWOr4Xd9kp6YYBCEyS59EF7+e4
TBwbFXWp+pb8J3obYHb6onSWN2J8V51BK6i3YNh5CoViPy5G1TGgSyGK5rDJaFKO1439dNn4IcJu
potO1jn3N0+eB8YBjegN7o/vJLr/JRxu7oCyy5KLbHC5ccjh2w2p+OxwiEuhNfBBRxMFNZnVVYdX
9pDxwqSS4O5Gc8lPghXwsZLoeY8jpxoQ9EjOJFJULOebVcmZD3cxliKiREJJkXrilXgnSTL/lx2g
LL0YQ92SBy5XK9iPGzD53jxTKZy70XlO4fBQho3ZiDT4chpgxOi+WYCDbngUc8ODV6YVlsX8K6bp
pgARVCa9qhvSwUcnLbXlC6/mMTebuYzDPKMX+YilYO5n1fSyxUHVzdd62cpnexEU70ABId7C40UG
bmJh4NTCkF5sqBP1nuage/2JQLYwkJZ+YjA0fA8cJexfRIhE4uspkE1r6+J62xR0JcLytFuVekxh
zw/fDZyUfqibqPEDKtwJOi5IwZukFsiPvSv8UkJt7g2z7hdgef9dPou0OakhvrrlFNcCEq6UT9PX
f4nsxFCRenmEYAzD82MvsmV39Satz8IkI1ABoJmvmqaMTvxawxfLSlaxgUvhqJrfkwEKRGmuGMqD
rLLDrvnXkU6o4tMH7ZZFnzYU9eFYhcNgcRxhH6TWaflz+FgqhAV7oyH3bqGn4Twoh8RBvlD/tVj9
E9mowM4F6epVy0ArY8VqAQGppwIBP7lQmOPHujUEFkM+dblKd5pSEUJNS8NkTNFWWHDStOYnb0oi
+SKD/HkbeYI98f2dy0cmIL3E+bi41deB8h/y51tAUpGcQqo+8bDjKXUP4w3T4hV/fG65pAbuwN2V
fKhO1nRDiNe4IXeDcyu8sTGdvoqfazkldf+FRynUcITvvW+t90z7wEKLQBDPb6TKky7B8ZGdO+vW
tHWNrtEfg2Rg51xnnNvEW6q4bmJG8s0+KBEENcirQaDConParYSazDKZTgzwMLI+4A0j+NyBK1SL
5K8+5rtfVMI5JCj4IrdDtKRc4F0zY35d/6nDg28ehYzHfWm1K5HZ79FgdZ8l38kT/ZuLQJOzqV9X
tg6paYijrSHTXMgoFPk1GDBBdyOq6BbnF5VWr6CFLplBlPDg3FvOao4oTM45d1Qt73eoBy+qvXHv
gKNjpUHOo5TQ98jgfMKiXQ2ze6ZHawRR8pS5gvEKToykjW4aKrSNZywSeEmbQNWmzlpo6LGWeDQO
VXkbDe6/BE08nigp/FVr5K7L1qGGnWieWWXl8LB85k6pZjCXlzTNAlkSKDyaLVsHJpk/Ma7W4sAC
A5LazEC7iebJwg3Fdx3LAAwGARsNaeLug1NziAkYGe+JTZueLmJVolvNu0VkIlx3olKLx/8jlEqT
T1Uzv/EfaG585JrqYXHfT7HhtTCItzmGWVOVtvTqgTTRrLeBlsoLcTFUFfUnc0m4gz1xQyXoD4fl
1HNdjW4exP7+WKhiQyKnsNRMDOFF/WGR13pzvoA5iqtJljSUEIcLSSB5B06r5cRL2K60Y2Cf9lZz
JNNduxEpb7Ag79RGAqVcHbFUvblblET4PP2Oa+n5Qq0m1phcoYnbn7a3Ao6ocbN7LYjKt+FLCIt+
5ebhn0YZay58YnXiXngZ6iY6CMhH6GpMVdIaqdOMsL9AuQejj921FkIErVW/f3uYI7g01mON8kwv
37IvGnKr/g1d1E+m+bwJLudQQIWMaYFqTnh5+cWnxyqp1+OVqrY0awZm8G3PWaCWpL5XEjDhgGbr
HewP3toVsVMgnico0MjcKfYUrFym1JhtFN2D2AkNbkuEKmuIFg/dkbSiNsV5aMEyHmMcLxKwTb5u
UXV9B4wpg/d8DLNEOk1oKYnGO4rSX0Am6lPA2/VHr/cmxXlQyGsJZEJXubesdEnqx5B817NWgWx7
zfr+kbzLfUAdpD5h9V9iJ+pJ0LyYeHfWkKSKYSQ5jw5+6sr3CBi4LyGoTe7fkIc1eaTN6ESoKzCc
jjOQL1TfPn76nC97ZGtGYvWB93/qeyzfbdw16PvE/+8pB1dCTwak8jW3+BRXaY3b1jXIYJmNdYlR
jLWFcHUORppiTcH8kwXh9bmRkct+HzLHiIb2uSM+mlqAnnE8JWIuIlQcjN5LpQKyLGSt7Gc2UdJd
sOnHnwEx4c/eDbHRD4vHGuoxcdfDUR2ndggzEgPrM1hMS+s/lmmoJPcmRDyUnGY0L6nMewCFou7H
e57brEGaUqed2WHnBY5vsZJSGs5gdxIjtJBxp6zmKV7BtvPcPwQzd3/kmPX1A0A1E0qihCclbkhw
g+Veq2vLkLRpef45Y2Sr3DjI1bwI7UatKsJKNOu+/t2xSqSvQIBOlVlu2JQRBz8uYqNKCmmes7nS
dYgua8oTwVAdHMXwbco04oGmFbMjHHDXGNnc6vx9GrmolAecB2e4ctgHxfh7WJ+HSq9GfzsQKmJ3
8vPhtsWLpg0+/Gh2x1ut9swZe7vdWWHlWdEdwFPjkoDiEWKJF2Rh5QoeWq/NIxjtdAHZWibFx+xz
mFhKYgvW+r3f+KDwOBkfRVSUOqDTvKWmzFOpb2mtEfbb9viyX+Qj1wI/p7yHqvICHtMOb+D4e+Wn
iNc7pi1xSfMBTo4rTkRd3X94IKTuI+aDWfIZVMZBPsFI2Un8dT1x5ChWmCrk0VF8xg7yW739DLRZ
VNNkLaI+BKnqvSRLs5Y72SKIV7mXerjang3E2arXVeaddlk9ea8SsU+mL0VcUHylFX4iBzZp+oVo
urwpyCHZLwLuxLKVz8THJNzOVBaw95Qt3YleX44xR9vui6LLrIqSssNQFcFNEIHnpgAftS/pKZIS
A/pj4KJhi/nnyBUJSPKVWaS+tkDG+slOkkI0yTja0vb8ph4sgoxrIV1FEQVivxboQxpgWB7j+sLp
mfuzN+Ad0M3EYBpEInef/BwVqFpFy1D+xGwYEAUeTY0DhROB+rgL48zJpqygv3A+Tq7hOoN628bi
uceL024yPeEF3CVQz7QuE15JaDCWrR55BVwMtmayU7YlQNUJ7lDml1TC40DB55Fmq08PfkiDwfhi
O5PEdVfpv3VbfUxQpzRHELRJQ4N+Dyqnqi3K9vZK0sN0itcaD+Nva9KQZ0EKou/U2sVVaR0LWBZD
MZNIiyn4GPDI60SWEcssG+Pe7NKhYkX3YHCHnkT+5KXotFQbpanZX5jizZwTUQ+XA0oQ8qbZJf5a
F+H3bDwIdBIZHZTrKN+2ZrKt13J5kfcZv+7OM4zB+VH1f693SY3sYlBj3A257eJmMMl2XweuYZHC
lGzRfAwQlpXDt9fJtcMEazo9eNUqmpE4urzjE8gn8InHOjJ7HJa6vVK29J4t5N3Gfzmxg0rLFIyn
C5tQVxl1NzalkvRJKJ01ZqNBLvDIIHf5qevXPK/QIYQHKDMaZCP4UWXb6bz/lj4dMihaTBE/rpgK
2hlEcjVhrE2lmyrD7At5PUuHuz4f9TjZd14E/eHdbZB2VmF+Xof3Eqr4wXDnlQAyPctr1Ouvtxqs
IXrVohjBwjQ0maXC5Sg2dUDpeatCid9bHW3hjgfzXBOM9AkdL7tocTx8440rYmVANvhzBbj4VQlA
ImVficpwMyiNHIlAxCaj053rplf3PaF/wcl/hWonfGz8ztEH2Q/8KkDfK3cXgod7JwvkqI5XqI09
E8okJocgCe2Y+6Fz2SFnyp82IAScOLNKigzsdp5QD3pxI1BjK5W2lPM8cG+BTir+kD7jKlVFagMf
znwZvKXcJusC1P0gVKNjf4MrwH2C8WIhav1x6ptMZNxO8jnanI2928L+UlkMJcL4JfrwDIcl+su1
DoYshF6vbEikiq49ZPASkaVIhptMEN+uLtfsti1hN6IJEmzXevjnavR11/vVFPIa9/H+1GPJWuaI
2gzDz8GzzZJnhyyHY57fQLJD4dl1xBAZ6X1f5MMT6/mRn1x2tHHalufP07yNkBENWMJB7aYcUD9P
M/aS6XZBS7CG/+VpzaVdxTT2VGPWhcoq00iHPziv15ajPgOsLR6fFiaqottBGzlDFvRx1Jq31DGE
ZzKiuzO38LFFW8siZOXqzzpKS7oe2smzDDlBRe/jve25zGYW82vXowrrrPellOfuNCppghhQjCbF
0NNpn3opCPapK6gTvYajEf4PW9+qDSK+DPPxKZxciYS36EYO+eEGpJwrV9yVHqiOFhCzsS7xGhVY
QzaGSydNFiNgFqFrjcBb0pKeulp4nfDfDeRDJ9wRL/DRkYvf0YHAEb9Bm0qiiGqcqvUJmxOObzBr
9oQjgl3/M/kxaqwnje9arVgfcNlNMjt4qlrNyzur5yMOxgvi30qAfHWnw8S3P+3lurSt6oq9n6rL
YU8g4ku2x03X5poxlfv7PciBqGKNwpolem4e2RrXhQs03lLlL5gXWjzJ4Q8Lqn0b/lCquUJsiFYR
YfFA3H6GLW3DYJQ+nOWNNekwBx0m4bwTZGe1D/RIiT/cghkm3eSx/ewV7va4+qbqlYzc/F83ZFwJ
KqcKt4mDhenyCUDcvsfJlmSnEiW8ePSiRajTBGmhbag8EERNcRXdPEZHwY94R9wboJnyBgeX7vrC
PM6Y+HnFNT0DdomFZZ8L1FDQrkeQLsJQPB7v690aOFXoJnqxnZq32+NrbEXeu+SMYxbJn6LkwDHE
x/DWTSWCNFgLp2qhUyfCPwgpWAAaoFy4Jo95Zo07ZUObRiodO5fmFwJH5gmKE5VOR33LHDlYlKUv
1zD9I9NiXFPOWlDWmlWmnhAVlRQBTM97Mw8ca7a4u3ntO02/MjHvSC6I6sTUaNgd1WQOZE/gMrco
EN59IZMZweo0NubdlgmendGrebRa19rcuJwuubywwmnzhjQfrVL9mqmzPmSIVq3QderMnheoXaq4
qHvbSOtOvt+YXfOanxBY3Y46fVYigDkTBajJZRpAY0TkPebVgXHGwvSo2AX5rsXvm31a3lLt9xck
YUIS33J0mC5IITjXtfBSiN3lZ26sFU9eJihoqfypD/DiiQhn0Noq0SRcbGZV+Z5s4HMVlxnlTQML
FqvQ/qX3qgJFvBvzPYWMhQlk5akmpDJK90sikUlTKW1c/4slYUpa4E2Xgypynq+iEeSniizcEhMg
nsDFjVcKiaR3/vOBl97a91Ku1jJQ5B6OsR9vLJuGS1X/veYb2D6oSKeG+Tggdf2GYL+db068tz1/
3gvhynsudpfavf1PTA4o8EH7eJwTCVWSCrlBJjpLItnvzvaEunvUZPt459SgjLA3gA2ObjcK2rB/
Jeldjz9Ef3+nxU7Y2Y5j+UFabSt1WjyChtJL2CrDi6DQPks1e9xXPw1k4qdRO4BG06GsCfTnbAzu
SKjLFKakEg/lIpy9xFLJBWEoARrA323I2xeDc/E2HZwn34IVa3YI0cSZTwB6gzkU4Bp3eEWvJdBp
mQ4U/5fJ3VL2ull2OmdPE1KbPAs2ez+lBpmg0io70jo4wMvpXT3u3KOEDn9a1LOonqcpCQEy+UYk
I/+HICLSx8MrADd1zNOLPrGY375TywSeZu6DOYFQmIV5WdwlDN7SgUUbCEhiFehRbc9E9YcFZA09
zZk79x2lYq1D4rstGJ6j/CJHLaz/WzzI6n6rdm81sFZGL7R8sGLDB3DT+fkIyVk5xKapcuciBSax
NflTYu8L1l4dKrrP0PwWVPpVmdO3ZMWiNszh+74mOuL6nICEOCVBuu+nK8v4jaBOUSGlzyKoo56o
8GOYJMt02yln4DrnRWynNLozYqtAoeu+L0ricPlGrf8RKqAD1HKRdk+th5STb7iTFVtJI4FD/8fI
M7SYu0oD6+hNXA0pPLqavzEJO5wUpLaBBz7UftdoXvAO0GyuqR/jem5E5ROvJizcm34uce/KzoDP
O4A0uww6dOybLzr7mXBONpyYgWdyohjvmh5taRqbjmuOIKmGnipijDdyMITDgj2UqDET4h5MeMQh
zlx8B7XvS+eAFTSztPsqkKzpJSn2pDucFKDYe6ppbS+O7RY6mfnCSMAE2QNbZHHB1Yu/2PHlqCQ+
HrXY8GGELUgFkXQ5gRStxgThehF57vhu+xbLandysgFWIC9yR9IWwKS/zyxpknpJQAn9eDyJO8X2
iArMPXvzRmz/mdYfslsImrSbRxP36MCQeQzHKinSIGbZsimzfu2U+7SHfBTuOZsiKpUwU30rk6Bf
931C7LXhWaAaaJxYhT7N7Vrjj8wK6rOPXTNdwtGQKWUv5MV4Ixv7+fVQ5gdyVed/tBKjHCSO4zTh
ePYecjawgevpD468TOZD646di23oZPMIV0923o+KS4fbeEvsJfcJaV6BUCRymhl2vkNV03mFB25O
3hRIicfPm43TKZV7EtIva5ga1+rXhzFXZEyXsMsQFkggejtoiZksU7CW71vfFJ0SzofozYdoXtYG
f5pKh5yueKdMmyzDIviG/EbbiGxm+UncGACio/ctgGXfozxeNLhwpCLXs68dAJcXnHmBqLDx/Gn+
wTKP0Ht29YuHWnXQzHDvrx28BEkg3iNE5QK0Cf0W1YeHohbvgPzvYmMKtJiytrTuMI2zM7VEc6LV
C5/vMd7HbYuZcxIB1prvtMDgJ5rHUVdEywJ/Cf6peAT9cnb4/sZf5hCTkGMBffa7T0GcL3CdwGUv
l3S/S8RIQlmomKiWWCm20RoVkiu3649KP/OIDTB0hK+aJkXorSnS0LLL5hjbwKobVh30XbA6990Q
6gdm9Wvn4gVhtr6cfUPh7U4pq6B9Wy9mn3vy4lD5IjZR97jtVVqE+kMc3EdxJQ7MDRs3b6r2LysM
1WtXuFnnXCpp0NSlPqV+Td6rfc+9NkVJJF30s0WqEVAMqMw3n6Q0PwwjQcxDRwQckuNwoAsAd1aa
4hZi3nJUTPoObMlAsr3Jjrg54w7u3+gS7lqmuX6sX3AfMO6441+Qz6GYKEtOa5iU+ZL+66XBLmjO
t1OCumbmRbr3P72rU6gu9eRbtVLfx4L067ycBG+nKPXOg+HDnffrYUAgy4RSIC1FNfTSXBgQoVE6
ZSRlrN8YLQkD2MMI10F4AqAehEHMj56fydl+54ENVY6lovn6GIoZ6SAqyVXvvV8bLL/lROFEvqxZ
jHUgIo2zjx3c/d5Uw75SYpptE/nGvA9QWVKFCFJo4FZxjER+PVZZU/OvJf2TSnkK9eyPje/0BOSt
u1od0oeROpVHl7EhtXxBGNidPeNamyiEcL6llwxVZs56OESfdj4e/QD2hCelaiCtzV8ALTA6G3c0
xmDSvb3WRDTjwTgekt+66A+dl111V+fnEc4sKjGrGXYzsLUCDP2sSsibgeFYCO4xkwqdGjAWR1Ok
VPm5npekf7HMk3n7sUzFRT9DCWCUD4UStgmvQRpsBb/scbRfsImlSohwgLWrGo0yj6oYfTKYKgaA
4QsgELEmqpveYRqE4+0RDs10T2YpkFNSHZ6T/mJIC80TSgkJygD/6wSM8dunMXVBajqchQZnis8q
xRAlGq9f3QoG8ol6h67DROdsFbRMn3Vr4o/t7kJCGzJQlkFasOWjUB51Vh+cfjmRt/2CAXaMk9gW
35DeU83zOVO5DRzhJxkhn1WJ9wbsRLDhXOfmY6/lK1fLtO5YaEk4A2Q3aGk/w+pP148UH0ugEyW5
p2pIpsO+1D4mxfTO+0T2Zol9Qfw75Dc2gNJDf/fR5bQPmS7U/ybzmfVpwY/ZFfjlu00PIvSJdV71
GsTmb4v4blQ9I1fmTloKsBylggMjDxRrFCndNJrrnpuKALhaKEXBWHuBPCtyLRXbh+7td1a+P1NU
zFVxAkJMEsYKBc85EYlsja2Vd0Sk8Ns+wTZ49f7DPP8//8P+D6atqw/r45udxmMQoJ+Z6eIICj5B
4ZnNv8wUg+TBlV1Ld1GPAVo9a4nqd/2ZCcn3Pa1s1gL/ZCc+1idGqgrLGS2hLndcpOQfYdQmCM4P
XXoGLVKpIUgIC1IJAETh8Oiygd1tz1wvNs5fvxhphFEF8I1hLgGe8HOrHyZ75op3hmdzyxmyDX7h
4c+8ElrvS9ZFc454oA3RUuDvqDYpiBmwDPddXZzfcVoeiWhxcYwB9JICHNpEG3s0+c3VV5ZNP/5x
DHvMAwfr7S5fjFkrR1ut0q0ajkPxefPokcmLknwUWiKEJRFtbKYbQ0lSciKIuQPtsdn8vHWZVhiC
QNizVZ3nfQBDb0ua5PQKqxHqKotfugntx1HrJQiCAcza4cFfGf2rmvIdLWj2kEDghnDUtSeQzZwL
fN/ZHad5F2ZhUw3JqPeayu15rHkRQz33Mg1xIu596kZJnfWrJHajel6cg940sts9kpYTkjFu7/t5
DOqcdotb0f6VcOdXmirmvZwnaJJxANiYS/CL7B/owjnbb/neiv9R91u1SwpQFz4LUrJWmkwAvjrN
nVjRJoIAVTuNzies5LfWgqQ6tV49FZfk7cuOWabmNjMYAYTIFzG5WZMJQ1f+ASsxtFPvZNpQA4oz
olMQwrDKuwVj1ew/JW2f+Si1yFwN5ohQhT90PpyDm8/jZ85oi0wcYmKwTOk9/aUryVOMYbukLtHF
dlouKQia5bkRrSj5EngYY3YQvWSZ3jp6gFnvu4l3c4zI1qvuQ1WDnW+dgxqO1CYcu0n9AjFgmfoM
Sb1kjlGjcfs2qP4lDvcgsah21Gx1PuKUeRAB7cH3lRQGjk7uXf7j04lb/0PKOy8JLBDy0CUs6whj
wxqIMGAYWYrcnS36+U/rPFavgzg3lHZL/uYrrNR57iHg93di52HqDPuQbiWT7L3W2aezpce8iQRI
zHUoSZdogX0+/Se4OIovhZodiWg0yliEO2nAW5lL/9ex6syOQjDXpeQg+uwp7fMW8HnaXa95/YAP
dwRGGD3tc6YEL/UEQsaRqEEZ+8JVzQFX2pPBuJAeom1sTfAG6nDsdyu3BcvXbq3e7R9tttshC8ul
1UShNxbcXajjJrx/riRbweXfNwpK4IP12fNp3KUJddZJKXgobVaEpBHbFx1KHKzWaQoX4sG5PEIy
Xd5CZZWSjI75hjUNj47UT3nzYk/7lMstvtkyoEzsxbqfD9iMQXlE9+Q7PFhpL0SJ0JKRwxAMq21N
CydR7Bb38FVQhMMy4BcImYKHLeLTzZWamcFHPUpo5slG+B/cv5zSNSpogAJkkTlRQDrgKI3h4qSd
6Z6AorElbHMMPr2UjA0AyrJOr9OcPrE1FQnWEw3bKt6qHzejtvRY4nWKoiWOKokGheCQzvnCmMlI
luG/TwlJQJTorCfH6xQ46l3NahDw4IuPxBrmduNivSY552gnXw9ud4aLJsENjcookhsBs3meJ/0c
yz8r48LrizxKuymLzUqxXPaUDUfXb+Ia0BC92isreaUvYHAKKEBgr+ptfwhZUeJIVQ9La1N7U+mE
QhBaHoWTIHKNPvmZUNIT0fL8QlHqTiozhw4TOcnZQC12PZDUC/iqw9l46comW4JkxsmxI5qEgqjL
qA5M8oTNkPCeex/gIw2BEOoNViTyTO5srwp/jhfcuetnlMewiM8vaWsOBUhxkIV6EnFQQTjUSOyw
tFKtupfhjQwRK6g6meBzRqqFXJmeoQLMHV02jOM5bEQ3j+kqN/CMNUUOJ03b7vYq3RNuuERs9F9g
I5pQPSYQkDJIDKU7ImPKAt1IbzBm329fRFGMMYTL8tqK8odAzI3YY8lGns5wSPy7V2dQHKdItRBp
36C3weKIezWyH6P0t0aBkT6/UlKkTCJAQviMyLVNeCJJ8oo0K7ckeiJg2dVWRONAr7cTNMwx7IXH
pSFcQJeOnx5zurQELcept8Y+FNDV3VtLAOxdVlN6bwNesH6+iLCewyc2W26kWfdTSw7vfj6msNWd
DlgC3sC6mdBgqF0YX7bkMl6CftiicJI9HFO5lss0vb39zBJU8RXj+Y6zR9Et4Up53lHJUxAuBsBU
jgbMc0MplhFxcGmRM5z4Hf30hbObq66Omjp45u0zL/SE6U5hYagDJnVJn1IGfIyNx0p+OmR6PoGo
qBgEp/b1+cVABg5ifYeEi/9NXmWo6OBvpNuQ8DaPErHc+4aAdVy449GGgG3ILscxpUZAWUwPsOSp
973CZnA6+AKYImGnzAoBIX4HYso2bli3kiaHs4ARepDMwL/ZvP3K4nbbOMyHVvd/0O4tw8AUZ4Xw
bZcQft/nHX+ZZEiTWJVlc4jnXH9a9z0nE3rtUhbL2VdVBCWG/xkXm3G9Dir0mb0RRdFtfpg7C83K
il2GnE7UgMJfHdwBC9cdOSAkBKQP6ro9a2ocIr86XEBn9iesoyeMLQj8gPo/D3896FhQH2OZX5Cv
McGHTh4jRBWaQryoRla/MjDGdkl0eJWB9CxJ8Ik5haiif3BhfvBY3y8Knh0JSZ0kSBWTIf73pfvD
L1dRFXyeDvVL5ukV/dyZxQG23RmzE7jdN/uDl5HWwnlvwoA63DqKdrHvrSWflLwL8kN9K+yZtwJm
h/exSj3hQlTk6RqW1ev7lf6ON43mGCWCNBOFfgKGjDCJgMpAixxz1RYGNpgMqhD/MoI0oQrlAZfm
tgoAj21eof8LahEERgjamo5kfWCEyS9dD7d8GY0xG4s6SDdnmsIR0DecLmUnWofmOjSeyHsNgdgB
q0ZX3HT2xcKZXASqy2TPu1U3iSoPxmNuoZYS/53whG568YieXo+RqN2+I/hbFBgjv3IAAfVBefN4
N8vi4Ydk8XH/BGs1T7izt/drsWneSCBcunfJP8BCzhOWXday1GfvS5SxJRXX45Iksr5yIgoToiAm
2xU8iGQfagfkqeP2XZxmMSU4TgyqXCRe5+bdWPXC0vWwkt6iQmjVNf3f5GQjiOisjcwLtutp8MVm
fLN0ybiwDIEmd1Z6pYOEgEkGTFxR3PjWmqe7YowgvvR+J0eQkdW2NgY4S0bLJu2E1zkH7/+mLWcY
FJPZ2ueNNcQRcfCTnLnb6KA/moKR6o69zubWS+uE/rOdorpXyHhl8Gnub5KyqNDkkMkIgFKpUlxa
yvwH+lqq7V05GUS+q4LokdB5PzjbUA1izTYzZwlgjz6ZENCAhJ6dZCrTxULgFDe0BxtqIrx0iXAG
lZZOY5/01l4G3RPTlXfcRWtXZJGpT5dSiWdQQH3Ujn2tTzm9992mwSTcXEVeOOz46SqR/DJZv1LT
Y22rlefJGVfgL6/w73wk7/uZ+rLzCgXCkyYWYQCEfd9HxgLh9jDGuTnOea29vUOmlWhAwyQIXTvr
BBP/ooAdpJK1LsnxS9avzN2CyJXW6aan8mKsuUjBBnKbMM++SPg0D5MHrjdHzyIdEnm4Pw4Eo5iP
pak0zP40n5bR59O9c/7lxOiCuOdWM+B54NhB+AUiaJ/xPIKCuqORiZbUxvwaXuHgysxCerhuSyEg
FB8T6eGKopOEAsylWSQRlHPZ5s0Iq2nuiGb/kxkL8nEzGYpcj70Zaa4zJnCcigRNSK5gob8ApfNx
wpdQQZIksLqJUSsGeHLjE4MHWb9X1KiDPxI5p14HWWztWkR991B22mxhjJTpTf022aLQvSGoetCZ
XFBt5vJByWdY4ROaV6F2ji8QUjl1OLuUbm/DtPMquacCAec206DrsZaBSP4ALB5ZkucFf0mOZGkj
GDA4RJYWOOcOfOxshirFP+lFTgOjsj7WLVVOI3JQeTWF10d8ouPj2S/FIj9IFVfinNXBqgjUxSfZ
2EmNoNTim7MQbW7nzyNAnZAeUWQO1uZYJFyd238KCjCIJb7FA0RlInA4Lqn0Hn+DQfOJFdvwLA2y
RLuvuC9B8dM2nctJFHgRz9sANmvscEIt+wtLyG6wfk5NnGZOTkZR0tbz9HY05oTaf0p0dIdHEsw3
ME3396XX3gE7JMBZW6WZIEnhBu+pah0nAjWUdZ1fJxwq5QzvDmpcQqmseDl02yHgC6kTRZj+kfbt
+ymK2AsP541WFCwnVZKPn6XFsdsFt7HvtUhH+Zy1i3x9zuGvhO0/PF4p3OdPiMxaDIzeo5pV+mXp
9uPhJnqnVl9oOef8VrkcNjfQTUPa4MfJWRfWeh4qLhBl3AIdUoGLEFGKMSVG/5WOGTM/Q5SCTwAU
sMfEVY0QR8ER/HN9bTMqimIxuLsVTIcqZrCaZWyVfcV95RCx4yMQxwmAP0UNCOXLVIo0/7/kuTvN
QTlWtAbEkzcTMPkfzHpCOT32TfpSoMNECaLXGRKcuLgkubIcskXicfWDkXIZxKiR2+20/Xbqm1z3
87fPzWbjVIYtVbT97sAS1eG6v5gstkbKpE7fuNcYqvYM2qDCO+2x1RgHqiAd7fOnPeNd5yO/y3EW
PflCotorE2ynEnESFqBwBwrGCqNAR6E+evxzBkPXXFosZukb4ri4VFvnZJfvdobZ4lPCFpHIPz+n
C1b3UjIPDqPgdWdhGJyatrxdJQdrL0iY3pDE7UdM9cy1SMnIZ9B8+SN/AQuXHDxUcJyT6tUD3rL/
erZce+2nRyuxrFe3hrZLeZQuFlAmZBPVp0KdCaae1UhfBSW3gLSa3Tky2JNCI+OjVi7sOpVRk2a5
xghRX8BRI8ITY6l/uoNCifGV+EqqQeHWwx+lFoAZ4flAaI1rA5Ksw8J5K2VzzxkP6ZEqheAmj4uE
m1yYctlyiydNcuqXEywcI/ivEn4AcOMJtJPAD2VyrTQQLqDvd/FLqJZCPvSo1tR9OqkU/FqX0dqy
M1OkjUkz9gZxcKOCFV8fz4iHRMSqJFVqXtpoWEeWxs2nVqlxFHUs7IY5nB8ltBzgaVgAd+iueSfi
GI7lxdvOu7F7zm5VuEZi5tLaJkECeznzIxhjkIIhCK5H9PzSNunR8UFJ1/Besmlu9MI4ZI/B+Dq8
KjWHE/+Kl7DmCx4Geas01NgYaq8L9QqFkKSI7cFYySKMaB9Wu7QqN9LuCnE14WEoGBVJj3GMLfcX
uDuPhYRqhL9HH8W+tTgag9MkJPdSriOdd2LmlsXhuNuZVQ0XpdzEDXZ3VQHT2Zd8/EHmgz8HY+3I
2mk5rWiqrW0MdzfYITjEPYDjoe1gzpTUvGKDuH0je1J6AWeerwFvm1RQnj/02kulXdjl8ptEWF30
tMxFBniABvlWp4y3kwXYgFT442/dITvrvS00Bw/7BsTWdTUIWOL3g313xfuFAMllHBiSSFKUOUKw
/Mq96YiX9OwOtYlcR89lYJBi8dG2uAp23kPbJ5js/36w/2/i/B8G0Yjm6UCqELHoeATH01Xo8/SK
ieienYKQL+IeAG13jcLfkh+qPdZHTwy8EDj+63XbZ1TIZk+H73SpZ9qcWKIxkkJTiFXSJwiNJsTg
qjFEYzuhfXSAqF3xnd4ojjnDmnHrqZ7kI9IMPR8UWjPsMnZIn5pfkMdE+Bk5mHZgqBt6HEDiSlRy
kiV8V7A8WQPCzr1aAAZ6S2QWCNesCRkfNLOKhR4IwZWowL8b7B3ixSEr9okixRbK6ZKuiYX8v2tb
uNurfXmZo+53R1sHGAFo9jl31fKHR7X8TfZkZQCYmF7bPltAgy548cbiAmkrcEYPPrq+viCAMslZ
oKuTncLmQx+51TeZfjFrotg8k0CGd0jFTqZs1yYD1XjMUHusVvWas31U7nftHGtf4xg8Y3L7
`protect end_protected

