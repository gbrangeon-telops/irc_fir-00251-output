

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JoMCOWeb5WJCBfHoFXpAeueDDgvCDiGp3AckCc481MQYfkwqbKzf91lDJ35VGRkR+lnFDdba8hVh
ebdPAvk8sQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bZP6jV/nU5x88OLSeX17wUzGVM/1H7fFl1OvjJVlfPM0WRyEzOpDDBDAUuNgnxFvzLOKKYEuQdGX
W9Azus4jUwU+zlgsaiCb1S5W3YMjUJKtbRQ/PvNNulBlTlfZaMHLAox9gfCqP4OK4hzymuRCwSK9
PA7SK6I+FbKAacX9y/g=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
38Ya3DupjVbpSJ4i6CmxC3OEuL9qNwdAvGt4GnhSmvDhP9C+krqPc261IqfCwYzwzxzaeMibTDWx
/h5fHzYF2I5fsXilkoEoRxiVUecJo1YSbQfTJW8OEBtN5aYD4EfWNZxg7GXemsfNXYAT3IQ9OGaZ
Z3OnlMzYiNTbG4DNtpaaHWOF6C1ZcpZaMxg6JA0ZIcSPls5SVALLcDt5FUbDAqBNYpV4JoWo+qsc
FnhESB/fKp4TYpfMu8ZebNdGwLZE/v7NBBWsur4E5vgpE96o2V2PrhB/yUkeOaYd/sqFfOVAPPYH
mOxmomWznEckwZ7yWdfaca/+EES9Dh2xe5bnww==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D5raxCdsBjNBeucgp+JNk0QydQuZbfT0hk9FPoXi6WfKMKGXanrHw+M0M2EvNOZMUencxzfv6CtL
nCmVqYCrBCTP3KURzHM5DqNYzQyp0kj6XGMA+Q1QHtCCtnTEsuFMkRdychCBXeOcnfn0sPqhPAb+
dDkLPxvSvOkSf8WjYwI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KE84+0MQOal9OYCn+WiAXywM19zQ4xYNV40iodnIlowR+vSp+kbADs/ClNTsY+01AbPMnO8ZTgZN
CGRjsRjKcpFcdHcCbRqcEDPJE7OK/v9PEqPDH9NFgGw1pSJUkP9IpUNC9/uKTepjTRYkaMQQIcwb
MA905J1RyQ1JTo8+T7ZjypavwIpWqfh9+/OtTNQBqe8xPN3IUu4u+7M4P7P5w0QOtT0XGFUOVu4C
5WyMVCFrGwdZoGJ0XcMR+keGC+lH3zgKGf7XDuZwC5nPj50Jr/CWT4G590JXwyjmGrh+LuEInmJ7
dRdHoyo/UrKvxi9s4oal4X1UmgumWAW7Jj7wfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
WoUSqohl2pRrU0zYISOEgS3fjCl6/1MuPsOWkfrW9IFHSBiaW/ILUNrqMgFH5IbNUI89QtTfH3Tz
g2P/OC8csKMuFvO5xiQS1aggRY7ashXHm7JNisgAK2iI1CRW7KJA1FbcxnZBAdq5y9cpHTya5tPv
OdYwNg/KYZVz9Vy9EXaKvCl+Bj1KkBqtsI3usRMwIUy60RESStnUe76XvV3Ct3gBAxpExNUA5QgH
nBXrEwjc9rLVVISzr5v+lPXze1yKza4F72Jbg6ZeLxQJSOhtZOOkb6v1WBx4iWEMuprm0HgIZT/n
p1YuWFJ+hpF68ShGI5pUU6mEy/OUW2Tis79Q1yV+JrfxGDWffbgrtbJxH8a2EpgNkqOgryLF41Xv
+/PSDg/t6WInmZ5ReUQtz+V9jY0XArHW1+U0/f5j+byluSg02YRJfyYBNGxXmWSfMyIUO0f49f4M
m1VwRGYfgQfc9AIMREkZk4TSsYJazLPCyBVXJBQugsbYLmENNxrQUWugCJjoge/1j+3MToZ0Wp84
kKIiVF+EL3BAeueORChxtvOiz9Z8WxLvwePIKjcOrGQdg4z6keHQt8K87+FQB2ObTYFw9eJbefSK
DfXgRWDO3PJfQLOdR0aD6ywdFdGIw2p6D051RteAwHYrYz7eCTRYPBz7eQUKu1eEh6ttCUMLzOZz
zv/MktC/dPOYj2+dThxoawypAAw2ZDjFD/5ZaFKrVNvOYuF3X93bzSosou5CPQsO4o8g8Z0lGVMY
RW6/RnqvHlaA4q2WpktuLTbsnBZ3/qcD29z+rPNHDWR5veZOpfj4IyCHwu1p6vZLgur4w6y8CSp1
y2EAu/QhEmSbEKRyBJwinnOZT1neayuXHiPGCjMHzSW7tnyVdUVh5Anmcf/RkDTrgbWse46mUzyo
+a6RfCuSvEgHFtxkeN2Bxmy3gnrekLXEAHwcx1YmCmxSXNT+QX/bJ7mQgFci7tbukwi0yVICBSFV
Swae+KZD9iia6m955QseEURW2XHFtCvyhPCRmmC/NyKmfA0XwSVlJUVLI6rQ/7VUwX7YH7rYsXbd
BichUGBdlnwLggMxkCEz/LqrByIAkziIYliMioAFUoNUs7IXM7sgqvdyQEBuMlCy6YfjyhCzC7xL
WwUBD3WSsu5b3khbt/oYcw7flHRynHrob4qLub19iX7Em4m306MBbaXgDkkylzdsAYxkw7VG4z/Q
Y4pvar1aiLGLdH/SJbunY7S0qgjNipSANEK8U0mASwSzyZTp+MX8oOqca1A9Mls8y7pMrAEUTrsF
n3IRT64Njamcm0ebbYHgvkRmkUGVY3R3irOk+UEoUXQYKdRaLPXERPS4DXg5rxRg0YLY7VcBaelk
54TDGIfPtp88mJVxgfsIiC3X6fiWvmRJ31FO7KlA4a3RID8daqunwri6fPJ2NDcCu1yBzE7GIFO0
beLRD7AVCQTjx5D1hQmR4QF0RBGlvLRDQ09cAaShGWdkZbLABlASZIRWapNhPIckiI0Ei2WBzOg2
MKnaTlTZl67K29rmU5vRd21heisyaEa+G6JQQn4vOtjOoqiJ96pVY8uRH5w6rqStJubmVlDbp6vS
mpS2+emb8xI6vijteGetXTkMeWU2H+InSJVS+46yXwEK2+ov40rplpdCD8AmCWRMdwyAswfHx721
cYLAXrtcNbdURfndOHe6wgdUeMlcOWnXL84fhBi4TrrnUSNdK1AJhGCfoWMuH+scfZ3dn2PsBGVy
zvGIcju5FjFdJ+nF5Fjdo7jpmEVht3kB23mKnqeYsjovQC7hDeGnV+TIPXCcOTal/YBz4+vHFHHA
f3HqG8GBqQY4bizYVpPPJLKFfoY/e+6vxGWTb8a+My+idGw2WprP/EqBykwWm1/pobzaoT+OEMDC
2VRLj8tXslasCxjxk2sHfTVnGerMxmlkJw/kUvHNA4Kg7RUsuYHPqjSoerKgfWVQFE0PmRto/dQ5
2ztYgrtUyfceAaAU4ZrB3MwKU3WC7aLYJWCtcbzPkdRptJagH/1i979QgvjCp3iHMqgFv+WVMZzr
u0OWm8K4oiRdECs2A5aEryX6ZwI+OocbWASMDB/ROPHOVXFYbu0QosOHPrNF3T5D+9Nxgufh9D+W
dLmSzOs83+ggUkE9zvQCZ2fQ5cEp8lX4tsTY05qpU2Op/m7OzOIoDMXHkk2Bhaezv5cPV62g2U4q
5wVkRVP4bLfKCUuC6Fuv5NSIoSSdk8566rSSePChlMaHcohTmGpNOXRSbvRwsdhF6ZiM6Q0o+eM0
UvWbGWPcIVLEoNnlzfWb6s9LNXsC8t8exOj/GiH7jPgsBeUYdls2nf53YqKFgjqaJVQTwsPUFEt7
fUvhEE0fVGXsfmbPqEdpSr3huI+EXeukY1HFn7FHkY3vVWYzXzB/Kf1tYoWfcsBwyQQPQO3SmZmr
BWuSPP7hD0AcRQuhGb2hVGU4pd2F01IRmUc8wmnZLrqRo0jH9fLHdyg5c+njOPbfqsRLE68Z6VGs
tcjx5YLQNshfZ88MCqcqLyEHQbFlW69e/UAa4+ReALHQCZ7BDxtLS1w9JnmvUbnHxBy6gMlYRkr/
BhYD3gmm26MrB39+2wJeSTKxridgZ7ByFJ+R4g9gto1mDf8PK3IPrlRNdIqY8RyT4aTEcwXNY/Xi
Xm5uNbU1vI7/4OXtECR6A9sbog2g49OlLpwS1gjczb5YKRWOBst/5/C6UkWJq2ADozluUn/azydi
KKnd35L9WKxLUcRpA/uKO8xZmnJotvxX+OyIH+Kx9o9l0ex+qcV8w0UgiZlpN2xQN04HCieEn/dD
bKxOBYnASS4xL52ez+RSpklT1q6EhJJ44q2azTWo64iXTHIKcTAFJ8/JWChiz7ItANhtedUJoBG8
TID3rCVATNgE+ScqjamKTY1nl76cJRaTJhNyLGDurkJf/s2kiTS+R+Pgxs5ie+/XHwM6byVVk+Lh
c8/ZDhWPoKddUR5iyS2dkiRs7zwyaxwTIRtqCEe9L+lfYQNDytcYoBEae++6UpzdDu+c9dnSDUS6
A6uQTaHqd8UMM84GH7HZOgUWyfyzkLmI9llNvFQ1PlYTHfmWdAZzG/rr80ZKrSOM+6YEJ/FkvZ4c
RdoKDXhvbpSq45SMlh4yMI+VVXVF1bkxUpfred2J+UGR0chT2vYb9/NierefaWZCVSIzLcp/IEvg
IVly0q+Js0Z1vk6cS/Kn8RGbvawC9iq7NJck9gWl+nMee8sQlyZt819eQrNLCcBQc5VfAFziVaFj
6EFsVaPSMDu/56Xh8eZP6/NLN3CUk9n8nTLsYDDn4lOIPvUQ9hQsmm09pEnwvqXa0LzKdoZOpdyP
dZ4+l8QZP7wqtUWF0RSgBHAZ0NvPqqGpytrYPMPzsFzpLkTwZqngE8jSdYbQSr+Kfa7aPgd9XFvq
RMPGTWRkZF/WexMSA1ZSBLrnglmAS+E7mk+U73kMbIA7fWr+orVgcTYS20+uyNFlG+WlRdtFupVU
gEPiorTEcnT9QTxaZHe7t13zBOPL+kQxWF3AtvdGgcizDbPYWPCchXz9e5i5o4RdJIwZ2ZwWHqsU
e97Wig0ejqFeXFOuxomR10AjbYTETtTH+/mEUnBSQWp3cXMs01MpPvEzGJe46nZPZ9iLXyIt3OEW
MwZ9XdZGBll4AI4ijrrviuAdCAOuKvszK2LN+Z6j0wm9J8UoccSxuHbblh6zfwTzwzdp/ghEeCB8
GeKgimKEYRBa9ab8BdwX1l1iMqhocpk1wQT91yOdZEItkFPQi2lsIpYOe6DhfirvTaPLspGCwbWv
c9Lb6p70+RpkCfXUOJhYOFV5VnCQ68jzM4tFOLV5/Ee8W0Yd/GEzConBPi2i21kZADR05UNO1k8z
uWPnWcc8CNxrXKdvlU85thjIt61RHZOwRi320MlGmjHB5BxF/KYy34ucGZ4FulGY0LkQqDzt5B1p
sDFYkrVAES0GpPFqXYkJ11wDFrX50KBsyxhgQW5hp0E1RVfA6bb2EQU/D4A4lpcHhXxZVj6VOlkz
5Xu0yh8Cmq5olMaq9E1ooI4osaKgxdNChgHnU+Pvs0qa7qR22j2uohJZBVlLIItbPnI7rp9s/Fvx
i1osqRbeaIZiEAqRGcr0EuWJGCf9hn+6hR8LFcyucg4iWxQEOUmMAhd6t22Vjk/r4lfKYztjzhlu
0tomAW/JPabhRKASyumiAv7/6j9UlMTxoKse+/QgvuII21Z8QugzC1S9QmhmFbcnNtz7VkKOI0EU
5CJZ6suFBSypLN8/kPzxeMHYJkWmJJmbKc0+0ecLkKCUIwBfkj+C8Us/sWrHLRXXg7XsGd6srOsy
igc5dT+4g2KmBu3g8jgpGCU2s8OO+nGdwesFpfsrrjf9Go2pq44fcRcGSRHHerSdQzpp7fTa1ZQL
MTVfeJJJt5HCE7V3ogC8txoaArGErapAtOw9dAiw9wverX/Go1QynSc8NVpwwtDI0FDL8Hw/7sGk
82yK01qaAWjEoTQ9r7pnW0v4HE58Lnxu5d9LXE1/JMfPp8twGmo9i8LmNISgVfjD/tIWXsnXS8G0
k+iNixt8hZw6YXYRiqv7JF3LAT8YUwUMEoOhGXp00dEPl390yaYdM70xmjqV4KTmES0pcjg0EL55
WRgeuwgXJv36/x/g0V/Cm91J4A1fcCOO51Wfs9YIY2bSb1Wc17tu5bOi1LcP/iigbKOU4/ri4hJr
ne/5N6iOEoYAAck29c3z0xIUFSxwZPL8LsK6K3ZHshSy+i4i7QPmfIYe/Vd0bqynkv8s9mnpKUMj
OsZT/GIp6DE/l/jB4mSL2U5hWeVWo4rC5XGYO888N79oaaltyUON/4GgxteMpfnRIxKIZoUZqi3Z
wBh7+G8SLXDmGfYW156p5waRpoB0VNgZfaUf29RlswMKTknaAbWc78NnMnsi6GTvGW2j61eXmx5F
yhmbf/Hl8rYvZGRz3SVDbd6FBiDL7ZmVJ0uoGOG6Ur52fEyGyyEd8axWjNHuFSElovSzYnd+2yf1
7TH6VZhM+5mbzNDO3+e2O5ot59J9ZxabZnZg1fCLGq7F9AAkTNPa12/qg5/CEnnD4jML6e5jR2WY
lmWbhXr6wLf9J85ZZyqM3R7e47hxvPyiKU4IBNrqY4XtFdbuNYKlkZotNqZonBAZ3kjRe8b5qMt+
KoRuGcSdPcqKEngAlgV5PhGbY2FgbJ3DHywNuCg49+FTiGYmecEKk1PcEn5H40t6gUuMkwD5ZL04
h5b4M/kQ0oD9iiV+L4Ob7vUCSTm92s0Ks78G4cXZECMGOFTVTlO70kHDFS+LJ75uAiy4cNciJ8N9
BWra3AxfezZfw3TX3ep5u28vkkpSwse7y57SO0pTV0PTaUbMXl45FA5bY1Adw21B6SyF3uNaFmQG
Hcw8sAxy2nbOZHg0R34hCD9M5Kl8VDXBBnSpXj0HPOo1W8CrEZwEMdGTzxDP2s+VpYHZ/Veo0jex
sGWAFziGaql5AyuSTEs2z6DiF8JL6P4VcKSVaCNa7hYi5wsdI/b0Tjv6kLiPT2jvjYhofz3fyILg
Hgz59MMlr3tiPxQQm33js0MCrdbJ7EtY6Jx/NuJ32m9nNj9+nGmz+Qjnm8Rafo2kvLARQGBKU5Yf
eP3SZIhVYg/fBmh9ydFpNNi+QNE0BXym4F6D5Ytez/IHjCKDfDKsoXoR9xFQBgbaMzcoKbPOHjY7
BqD3qWTcB2jKzsRkTiVBbUX/Bj9713lcneeIZQYZdzV3DrnZbg+p2oDlSQ/sqUv2rXYf3BqsAk94
AZeWR0FeHGqYdusQYvfglLVbpqWly61H2z/P0s69BAAsH8oiCk4qoAuWy3TJUSa/1hDnL1zytcQ/
H4N2RuzwTQ9GwuzzJIHrzNxAQua9g2RIzYC0TFjfW+gdSKmWuvgMKC7nPfE5CpNMcG7CA61gGpd8
x++1w9TVmq1eJmYbv6WsebrpV0DkYr/R4UqXn0fxWjatzWxdl3aj5+gQU5UEtYe4ANvhOoWCHuJK
4weU3244F5O1lCvqEeP09rEjPNYli3Wup70Jmqudgk2EnZ66RqOno9EZ3Btcyr97PTnIaixEbbq3
hk7NPT+lBtfeGID4Bi2RN3sIePEuBDbjLrYZSkei9ZPMU2KGk4BBcDp3EnhVgJA1kTN+HGd3dIBn
sbo5Kiz4C25L29A7WJCSKeQj59wEOgaco2Eg0ljP1X999kOE6W/ab8BwrD3+g/BbobfCe80qiDbp
iGRKX2e1E+kt2h+6Y8iRHKYfpKRLK844wLNe0gP00JDjykkUVBuCJUDB3w88yJtpWZ/uisMN0BVf
43egco5hUAfCHZhPVEu0acEbTLZyG0gov06KrrOmCAulmg8jjZ8wKsRn5QDmwjtbsDV/CHy1jg4v
AW0ES7ScqJu5tcnt2YVU+dspGKvdLVV+wWf/dXeXvEXVzf1ay4u+EdWN6ZIDqP6/ZzU1sYzmqHM3
qgLpCU0bV03QSO9PQlQR8VK404uwexp7lL6eXtyLIJAciBYJzs1TzQH6YN5/k2BSxlT1ZzTLRGmd
GgXkT4H4NjHwaAB+dwzA1+1A2sGpsQFh+IlDFAdEQ4EetpPNa8qEJqB0msYaulUZenL+7dc6CydE
TDBBrDXWPhGQwQJGzRt25vh9AYwW8+ZImrN9Oqo/te2MDiS1qEV4fAFQSDeD1bTr6ugUFx3WR+Jb
BB6GzWika2RmyGSPsXrETrHbtnlE4DaaJ+tBwf7FcIlF6Ch2nDPqvCmsDHhbH2Yi8AZ71D9lc+jB
pllYEscsF0N0GIVhJ31+jJhhJJsyfgh8EjYC6rKEm3WpUL5H0N1lMMvhifJxwyyhZYWkZinWF6Rn
/zUdqFivqxIXRSvXDxJr8raKv94vQZe13HFHsYcjT49UBi4IFF7Iyqb6v2w4C5k23qUwXOYAjtI5
Q233OhdlVKo27IT4cqvFECQbhdbPxGRodYYyEh1VstL/ONRtjL7i8mGMGfz5gbWe3Y/H2W9lIsxv
R+7QYTYUvpv2Giz8oS2haycUQMQXwEpuvXtuj5sdlwf2gr3vgLt8PYJAz/0+Rap2ZoNxgYlEQWE4
STzC9et9DKNNX6WT4aoN26zN+VTULVFk2SYbW9ynHl0nytbkV86cULbGdCBxa/UOKZmB9Myumvik
aMRX91ur92Yk+W+KT2qrYNJNEBnnfJKy5cYCqpM86dEQBj7vXFkSuNzU/1Bu4yEHATS3DtVNlebF
uvq0YiLvBpc1B9aSqk5gcvkX2gkA9vD8IL8ioLmhD1kw0iSkSqs+so4xyM0XhNydFgf7Eyb7ZY1N
heBSuj4FkYfDTgXJQlV8X0cwy4GuJUbTWFZvURir5dCTn+xhHD84Us8mMCbUzNS+25VJGjHZHe/6
ymZhNADt0S68dnmhz/NRM52vS7+kexqW/hBbr5aN2rjU5ICw/WbGiWwfcE9Jig4dDJYs2IUWRYGr
nrR8XFe8Fq9U7zBcf9gCdgfv06uKYUBgzngd2YyzFaTRZPwjXnJ9V0apYlZ9OUfdVZgrco56J13V
PbSy8782ptjGCNQ2o53NYEwYR8jCeJt1W5Vymza2ZGpp96qeI1851yg6VuT1YrUJEEp6W3HDL79O
vdF7JpXD/Kobnr4HBtniwijRR6kz0hiejD8PAyUxI0bI+XShhufFUHIqVzZ4+WNVJzFm/zGkQfd6
d6Tog2AJYDH5MDaJZdQ0hxgSNVmkyddSwzhhK36mZoCj2UMrsMeRYMMQn7AQfe+gppk0Y74lIgjn
+nqt9SlOOnZtsg==
`protect end_protected

