

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
US2mB3ZU2xYMwSgf2KG3QONmAU5qxOR5gFmXyP3MzegSXblZ76jq0dw3DGi2XivflSREvQG+tGNr
93kJJN9RHg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cVCcDe3dO8A3aQlcacvtDrMlOeMM3iFulWP1GnL0AstVpxpdCCRRxU3UHiCxbevv+1Dnaf6o7WxT
G4MiJBrZR0NZpyZrN6elCTa1aex/x1et3mJ/kXtaSnXZDYRGWgFlsFwFLktb6kdkyrjtbx1rPCM3
CfbtCvTObEIGzIf/FJI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ybpmXaWiA2h4ouUhToF83n5FZ6mSwY7i2SbAGhh214jlEV4EAw60pDdsC9S1DXRUJs2H5ijqRHjq
O6r3TnjNUgOULu96coukm/eTQWKkKJe9Aqdi1COsXCRXpY/qPst8iFpcYgvP7x9BLqj2FuOVCOp1
vBc1X163t+3g+Wnu5wdB02cYtsPg85Aym4KDvpdGC2+lcbTElJIi+JurCHNEVSPxn/s/byKj9Aee
BWqSso/XFdRP+TM7huy2D0efcTINLjUE/2qeG1Z2VdFBpyOvUXxDlOhNEr+qAiw/pCiqNyrHCapM
TfSbH498t2P5uuhd9n2zpj2CUOFq13OvODvHsg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o4nr3qLm7Rem+yVuZpGX2Dwzye61TgXXpiZsrYTQhxAIOttLQ5qy48oMqssSkd1Afuq4E1AgeeLD
pr9heGHoD5AjWxk13hv9r2YUI3BND7NaVLyrx7mIkF/pxjMjFTBF3rI5FZuYgxY00aftrEFjG/AI
XeOeb4w/KZQIUde+tJY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dHlANyrutuNgAtytsZMPMatpxiEBkM3u/gDZ64fIbSRqU16FBJ0WguNKCot1/TeXAq8CSJHQCt8x
3wxDlxfMsEEJdw5OF5Pn172rV07Ce6wZ30zB83ou1uUKjnNgy6pYqTworLe5Tj4SYl9VY0bcZ0g/
rN0niMih/6g+8XwbbPNRS7in3icwjpeqxdXwsRyEX3dbCrKVz4LXcfmP+ybNfKunFSp+imrzoFLt
cLJF8o/HdEoH/59p1whEdIyNin1+Ra+5d2hGnILLEgUP28LNS8Xr0dqjxGFNrkIDmtSmsmF2E1fl
JbLYu0fIIENjFn9nAJCzGQU523347ABwMPcyhA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5328)
`protect data_block
0jmFEyNUBXIKVLvveRXwAggcUvhkwn0G8kqGRKZFpQjQOt4zXvKFYKd2RhJpTZW1loUUVYdJzmgg
0C2UhopTnXArJkenbXs3vkTTeqn4mUVbI3GGEzcF5Cr8Pu/j6Z8W7R0DQP6F4u0CcmYSePEf98B1
Yy6mZKMKziB5mVniB9cc+fiKGc7rF8vNqR+p90+Dv59Lls2DI0PdrdPOk+Q27kBIvASFLXPB4yh4
s6/s5xzLHnKCaMLFwmLrtJKGseSGniIBi2x9cZZuICNuYSsiX+lKeuhrZMjnY+st+M4jgEW9fzQR
B0PTgX9fgrWamOIk0X9D3UbOlPotjKFf390QuFJOdFb11UteyUxuweYDmEVSISiu/TJDWfFdJ03L
OqM0bIQXaJLm7140sYZVtD+TXEih7Rve9XTtDcL57SE9K+TRL9T6rtL2ghcWep5bTfHXYmDcnvJD
3TdUiabbweyD6CBj3CPPX8+MouxuAuRTR9RVU7Wy/eER6JbrWnmz6lEBrVdoioI1BiEqIXP7L4jb
NpVkcaaw0V/BfMSaAlPMegaXO/xPd6Ajsex9PWRNEvcDwU8ApSEULpgAIn1NZ76mOJpQKwfmWrAg
Vbzlud75T56z56Vh/lotQK6/ESnDxzOEa5n14XVSJH4yIpEW6feEhc3JcZnI8tWfBfRYJtMpOEjK
ayJyDXF7Dhkb9+zSU7jrQ2fGlS273hU3xiX/qu7qYu7TejNzJZS8d0EWhqUGtIat3yzh1MZEoydg
EKsH3T4+A3aTC0/ULrfWnL+9WipqWS4ELkjjfuRu4kt2lJkiO1KWbVan7CneaROOeOtnXrPM+t/F
RWMs6wN3MN+tUWeh1WISCOLjE3o3KHKO/pyhLA5CRP0yYKoXrrpvT/pgriMWgfxCgHdhGoSWqPi4
/a5fhGWJKnujj1KySu1fBSJP2ydnKu7Md9y6NqhP+wYC5uiwNk3GJwiMwic4KWpecHRyBXIW3LC6
pgnAX97bavoKyIIABKo3F1kdsfv6ZQXIRvwlspvSqBZbBi9ZF6S6hood7o3LanHcLf+xuY1czRXh
0RBt7Kab+5OAYecKooSbdkrQ1VFiAI9Xa/l85eXw8cPEO6rDK7mfedeWu/O574RYiA4gf+YqiIYR
zk8D0AECsyL0w9IYe7oL0L57i0z7UR3kGGFKVkNMbHaND88Pn98fjYa7/B/vQgHWY6m28goBp+uF
dwZOlFiZrs8Wc/3wCaLeuJJALdWyZpRnkbCdySU8yq+KVbxHsrbZGCKkycYs1Hxi9//X85igVJhP
BdAquQNW3X5XSzjV0iB9iVvt6pdgodrsVsvs3fQsXSwZVkqd0p45kevqam33x9neUbNUNkC4pXMq
KMHauyZWSh0qXnzAXiPDAeoWbypzxKPR0smyCjG/t3/Twgnw1MQ9Cw7iwarT1TkwmRnLKiNehXrB
m+w8LhMgTAV97beDDPP+2jvD4ba2aV0R44eVYtxuRkyJHLa8vYmyR2mfxPj5/8Wlk7zw5Tfr2hTl
KXFAAv7eQXtDGDF+PIE+UhbbvVAK9oe/UmROb+eWTmERFMmVC+L9YXFPbNoVyQaLwwxUO/DC8m0I
9v4D12LSZqEW+2K4/lBfIsmRc78i5MFEuy8cltmMXnaCAxhHqioXkXixwxl7/AyxDR7ePvURt2Xk
Od1c+37YjTTpTmojNAM6+5kfyR1WpY6FPdlrNSVP4vyHKG/dZXaEpSVIMPLqRLsw8+8dsEulsRHg
Ze0o9QsdVRhGStHWwXx13K5zlrXWheJ96Zf4wF7MUlZLN1z6/MDFMHdbHeZ+kekRv1SDuHRx1IWo
WtjCfpDaE8B9cidDi27jSP7DYh2Eyjb1H5kfQw+Nz5hZFESwr4nEXo9IFBpurFBDq32ptz58iXjc
AheXFQcxyOO1qYrtJpoHaBJp9Imke58CZTKOo7e0z04JfObt1/jkcsGVmImKre+NHFep6SsGZDeJ
y3glfGasRpJDn4deYGkZ3X+hKg0GhyQB1E9dFNZ8yXgJFpF01JBMDLMXkcmFU3pQA/ZAw+Rq99hf
blJeVBbSb9gmT+SQ0Pa8UyTJewMI/3IiIF+xlALMNp/iVwR6JLbi+p9doCQQvviwaYr7oyD43ygK
UyF+AUpv6QyIz4lUqZG4mXS7tB7LkCJ4V9haIhP3un55H6W3gHJZnyKiKWzF+7PSCw7Shewd+h+t
kA5zQbENXgQlOpOx0iFmHpBqkV+9JoCKcZjCJZSeGUlAwDnGFkY3q9xw2wTSADiLviHhWfBkBTcu
oGv0owEMk4oYPy8B+teg93GAQMEfrMVqEp0JBsBNwrr+5gD2RGbWK0sno8huHOd4KHWnpmiZ6UD4
bhZVJ4OEnnjnLpJ4unPw5QbbrjeY7VIFIrkQpT09eRr+qi0qrHZs1GJcoN08x1YoZ2bY/19fxeXV
7PappYUj760iqF+fwjB+d/1m1We9gq+VR0urswIXFLeDJTHIBgBuNPGgEQTYbMVceviwHsEYuqEE
6IwflkdttT2ljYEU14hlWiRev1TuNxIF6t4gx0Pcc8oMHr1CmZCO6IFNNgnihwb59z+o0Ab0DJl3
y+qGxogILWCqWyu5R3Z9m/bMibGRyVI8uR21QF7littiVI4qXlUKnLeWHYIG+7a5dc7vsMc5DtqW
EiRtHcuPNUrXSRrzh/oYv0caeGykAF/NsxzziL3fpCP4diX4YyEcutzCbRK8b/FP7YyoJobblQKu
MmK6EPD1Vd+2j43Qlr+FoSS2Vguz05VzreWzgLCzrZOqGxgRTSbGB5Wel84BMZFTxqCCAcoVZFCr
0OZOO6ZXYUdWUinLxB0X4I8YVdp3GqBf/CboZUZY/NgEycP/GnRCe3TAFczQIRzAFd85q3jElcb1
S/GRa/mkOCJoNAQAR7nFKBJFOL+7gHOU3idnI3jw0h+6B4qhxbloKBS+F+Mpkeuxp/Scsgy41GmN
q1x4OFoiuxoT/QmC0JLuBTjBbFHkRgPa1YaFHqAWR2xWzxlNMcGDvTXSEoj9bQP5Rxoq/upVLPjW
zKbwRXcAGLkOw/gr/ogVTRqH0Kba++MItJOB6l2NZ7YXP+R17UDpsHcfHF6RE6rqRIl/J43bQGCx
KPmLWjuTgt1/90jSY67T+qDkGxvSvILP7LbXZk4+/zCX7Oa+yf6sjxMzDSJwyayqoNKFTYqHLfvU
Fk5jmA8+UvnNOFx/IJnCTAD8UuR/mNYUiy84SC/nthKewF3pojMh2fzP6TMJzluAXmKSgs8wB5vr
vcmXUjni/njWj6uYu63Iz4MJGjm47ow50z21zctS9/SuucbpnwJCDTLUXWKmpfYyl1GLdIVapVSL
pPX0E5feZKnFFy/7BBuifxYIEXQqupil64L/1UhKYtTu3XZgZI/G8cypO3+8r5PiI0JTVYGUKeLa
k8RqZfKYvyr72zL34n6zxB+YEKUpE2irYN17ShEiYf4XsYCycx1R89km7+E7Gtabfm/IA5bgk52L
mOZRgGQI52izUwOSdMDweJaW3YoK/NRPjkk7Yqmwp6IhSfiJTDyz3FQH45Zsr6OqolNd9yclvWCG
JTyub9r6R6/KS+zpLmvLo6tHlQI/w6YZy+w0RYL5iU5fPL7aC6E2y7dSmx5Mwe1wFXIKoPi0jx2m
erwEJmME+KU2r2K4/iK/IPgTmj26/UPigg139kPpsBQQWFWMGq5Psjol/JgXwlecgwOegEzfO3qM
dxCUHa+EMzErNomSH+UWVJQvx5RZFw6gxK10vVo1APlzEz/wOuZh33kAmUfFICOg8IeZ1gPHB1zZ
/Pb4LvENmz2yw8VzNYQhZf5mspB8gtiwrQoxRO8eDBNl8aPnQWWcqNCh8Wx8x+2cnqkgD0dWhLng
HbUR93dl5972fdn9PsFpl+o/g3D+cG1kjuh5kbStO81Ra8UdVM5LbxEciDcuiYSZNSlTogvu+dQ6
qDx1vDnL8/NqpZdA6P+ZlSPtJiPDVGSAhUa8X9HhJj5uIKe3d4w9PJewgav5LxdaTH8m+HOjWx8W
m6zEq7NAHm8e3ifoYsjRxrjoNkSvs0wuAXt0Yu8/+X3aQJCEn6qUkePcvxPISkxN8RoEFkk5aQVr
hAfEUAsQHKftjPBmXhmdl7C68lwaaiDDLEIYvrltjsnKdQeG/pD+Xduo05Fox6l7zxG3band30Ll
BkWbWkriwldkXD7VrSfcQZ0R2hpIAJ9QELl1wxdlk+vppOa+TvC+kA3N4Iufnb1uKQGOACl5QEl6
UGLBHQ86FeW1mFB658x5JVMXB03Mkv07H1oPfiFlX0BlSSTrzashfQTuknS1zjzrYRyKrBd0p4za
uYQXLMLudgGkSyd+h98rYFSsGcNKKWAaC+jDthwDd2ViiUoL25+WacNTo6K0XbVgxX9yNggdPjyH
b5/irhQ0gZx0WJj0wdBDw/oJ/m9Tzsfd5GU4qEhPY8zdaS9SZZlhRbRhhFuvN/pKpFlHgO6mAxkm
S8gSv57Jh+F5wqjnFsUNlmn+FqvjxYGh/HagXreeOwLfBoN2V/t4e/bN/A7dYBW+UXAGuiR2MOLP
raCX7NjRU1iL3m/rJK3yRf+iitqISYk2Fy+cJ+77ql5GbPCxfV/7lcry3Mux5YCpMXp/ySPVVVlb
1cLKS9N6KdmbY//aYihHLIIApjy/xHCXDvGlmqu9ShVw5zqQ9Jdmu2O/webOKznHBxVwopJZbs7T
rKZU4cJIP6f4Yh3TazAuWZihqnTJMPtyc8qLEzNb99TWdJgan6YrP4dWfUwew6YYIX/f+kOhXlyt
D2hkPrH18leuwG6TUVw7l3l399FcxqaJI2RDVCszsUhc4vxZQj5iO/J1papI/VmmzU5KGiL12Erh
1mlw7SOrhwbyYYIyqarQUwYqyXnCRMmv6ioB+I+dHJ+P6I2DYHbUcArriucXWIHV6L+Ni/PnmmH2
Ydmo2bufMmaK5Ry8WzIoqfMlEbMevTnmhFLMN8/EyXTHOJ8nFVROrRK9gWfQ6B2332JYexqiX3O/
DFzW9v5O8zd87A2Gpigu17mu/cTf83lFddae87ufGjgAEy72mOOUUXKG7JKXzH1/elAlOKAzX5qQ
VplfCchIWmrCQH8JQQ1hkqmsxgztcg7whtw+aQlE+6GxrQnYA7Y4WDV5jnpnIh8SCux+F9XOxDTD
4MgJldnw/T3PO/1miSYxz94+hAIkRfiw6MNB8sOBtBzXjs16i+15elgDEaNNNI0Hk2+3R0egTO1L
QU+rZgB8LlOlivrHkmb4xEd+6zctcTq0fn6/I65UE4vkjWwcxDGt2sxYWIM7LKGd7sMGKhyFQ0RI
55bf6Y1ei+MU/iQJ0uziVaNs2MXL1IoooeySGZXEVwRt33qgtNtIM4PxLpyyuZ4+7SEuP0jK9qqu
7jtJ4IQ2tJ4g5bAv7YmTXZlUkpvD+zqZWHqkPSJrf+GGhofSEh8ycglBWfr+HkPmdgD95GdeIHis
X6h7W3nHEZc5D1eFe8KEBwASLh8hSBEsOhXtlT9E1tE0oBJ0Ml5zV3bjXMDzpnxchxcX0jdGr/Al
7aYH3l4v0Dzx0Gn+FMsgvOvDefeWlg5RgFz78YPGvWt5uMIb16rxjO605jaT69v2/gCMS8e/dJWF
impglALCV9FSkTaEsj0T+VlCrayfQ1Xl+hCLSL3sXT1fDKXfMHi2tc7EiDa49ZBGb52r6AAXxbxh
N5ufsyjSJdcskuSZeO4ndxzFbnNHIJx5rOVUekfqmwobK6uGudtaSHfrErEr0x4p0Gy28CmoeVNs
KJswMbdXxXJ1OQXdb15wLyl6CIRbQOz9w9fuZa78G3NFGVzDOonFuUZjtzrH+EseT7cELWjiYK0I
QK95D5wMXn+cpkGGT1KCHodVwZ3eJbBSEosLhjpBKT9KTt57rapflrmg4NapiyzuLktaLd2fnkQf
H4iLmsUwQDj7s+sguxp9sBcNHqnJo3GHuzW+CWxp0XMihc/3tPAPv+o56OedBz0xYsD6d1myd0ee
YMrONmR/reQYQnEachxcLke54rB1Xc1ajiJfkLmiMbEmSE9hlSXmb5CqGlpFrl+gIMtwW9ZlYFZL
FawNpgFZJgknZNn2xqCoWBvA78YE89rbxRldeFSSIA5dDWsNJo8DlpLPVbqj3RkpuW+kDMXpFGdP
CtO5Xz3IxVFiTiKfGNcrVM7KsMU6cVJo887Cm9rGYr5HguZRelKOonJBlUsQzEk90/wh3GgJQPwS
WG2ARBYfPuZT+pCQWlq/+I4bp/bcZjKSptTZbR8ANmVQZwbj9zWFRsjHm42URTkdi2kl0gQ5YGad
BVuMDvQxPDZ7MOcYEdwH+QhcRjfIoJ2i1XwWC+DijdeSZP066mrkDP2BkhRvLleoSZSWSm+vbEJa
/TKJHvV8b9QCVuq8xS6QsUzLlb+M7X7LDiHsSvoOkw+3OIiKB3v6HkQ4qcexN5li6yA1HN66bClk
FgPPhx5SvodBdp9ORIRoUmpDnBMLJXv1RyB31gjndqpep0IfCCmgoM+7AQMxlmCewsHpg67OOD5w
+KB8hJBPmA5bk9Z83BYfu4627bGuJGsFscGB4te4P24oYfaPZ3kBU4raEXhLqgT1yN+r2VhF7kQJ
QMKaEJL5uHDHwVQq0xOQO+fSucHCO58LDnvYyyMFcddOsO81RpiAt/qQ1kIEtizP3hYv+WX2nnC1
89XnYHELXK+rlHm1Tk3unEs/RwpKwVku2Cit5EdDOj5zn+LjP8nbaRnLp1A7viDgCADzROr9KQXb
gtBQ3wvdUoFp88tXh8aF9n2lZM9cLX2YK7tUey1eI+id/e1od2n2IaKbiWErzod2fUSpRkeMeMoJ
apBuktkJz0ERb7pUadqlrmcDa4NNDrGsUnm+UH2/SWCu7VvFw3v1RTMes9EWS7mCRhcAMwrKKcbr
X6GyZw6JwHIf9C8GD8n6YYRQRTXWXQdzBcnF6cfVm5yYOdAV+4YpSLYMOIooAp8WJgUqlpDtj25R
nzo3ZH2uh/7s4aoUN5jiuhD7DI+mRxB/Rmd3jTN/MMXXkzttQzjKIPXigPttXZCncZG2rUr+llkS
8xSehFhzHxhQ6HbbOoaZTTTl7l6vfqfX8XL0
`protect end_protected

