

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2013"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SPpb0sHtYr+7D0Z/NdHkBGKHFj6bPnAk4zCT9Qd9jSi/NZdzqHWXjKwgFh3NrYG/AQMVJcT4R9KU
T1kWm6bsuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PM0w38wqoKZTqxD5ZMv+He7u+x4mAKOhS9vNWqYsLtlMu2ni98hkp4Js0D7iFCQdcFCu3Jaj2Vqe
E0m1H+UGB6We+zPa+TnTKUC9+mxtEW7xpi8i+GVKfIfe89n3euEibIBIS0WLtZypuPRjuzr2TWw/
TpBFYS1oUTQ1qwWguI8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2013_09", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OIEbVz6QJBHT228fhImFLc7Q94gbSg/QOSgeKpAp1zRCxot1azeNL0EHN3pwZU9Qs6kuTNEAn7+w
agqdilWN9rl3uQlRBfW5KbIj2khza90rK/4UYrbcPGQyMxF8l/LBS9RaSzH8pqlJgQ4YfgwGNaq6
EHHkNL7CBEprP8VBO3A9geAIYBWstNirz3P/01jzH8PT87csZHkt/KV+1ancvBdl8zy3Pi5RrOtK
WdR5qLkbXJ6m4DjaubrW8HdK/fqusuCVkVGxmajuQw899iRpx5AiTEwKYKOor3msJGxdK7STL4ZT
S1m+Ec1GdsxDwYBgiKT0A3c1/unIYBS6y17V2A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y9qoE+tEhAFEsAZgxeFxNUflksEoY80RYly6rjz4X/QwncMYkOdY5w8AxmW4IYZfWprQfyfkxMrN
8JuXogLHC84iIPhEFIhJ/+RivFHW4gCUIf9NTOGEkQza7hd31B0/7LZttbZHcfTR5stmYGMhB9xi
VCriwe4C9iR9zFvOJxk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eCcOM7HngIZB2JCDRQ//SPPOptJbtDQ6WJM03A6xR3t8OhM7+MFavTdB4aR11UrppwUsYiZCHTBc
4AdaSSNbTEcILhRaZMNZ85hgqiNgFb3YTJu8ZIWifM+Ad5U1zkzbH1xsVssRl/Sl+cf+TCDh9Psd
UOpjIzWfsyGgyfaSSbczC/DMklBqFcyspqzOP0YGdgI4It3e5xnwDvYeewRqIZggj0RyjkJH8PxJ
o1XlyTZFQZIIFN0x8sDbcPdsUekU3pOCvI9JK89jigNzKmLJRotLEgZQt0B8gMiz/gm5u0+k01OA
f/7Xo9TSexSaZ5evmswsNTBQhg4v8j39bgkh9Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7744)
`protect data_block
UDIi0UOGNjwzFlPmuAd8Xdy8fTyU9TDP1mnZfLDQxdoAdI7Wcs9fFvj5LsUpAIRjteag22tQSlRC
jm3USX+QX3kodrG+/D3AiAy7kYQciWm5DXn9oBTe0roPbC4A6lf4FQ5BrO4Py1rKYumbkG4ydy0R
0I5jv6GzDpZLafLCESbUGeCmzfFQZEgGfml8Ygb9Z2TxElBGhiZlIbvHQK0GjFI/iRYTPbkVFLT0
Q/CPOuAOoLQ/7Xox04TeAsXdDgpe08GCgMcmAZom5YksFgSTmDKa/pKaAb1chvAGSNaFKFNTcF75
BXp0+QCVO8NHydXXWr8w+3SnF7thGSWW4wqL9wxAmVJrP5OO7L+J0JEu6Yz4c/WaSzPQnIlBITZI
Iwn6O6W3oqn5/B57Wd+eGycOQTDP33xqD4q5Ti6PFN4qY8t6xxFb1jolu8tvcMsAOYpLaBgepuMJ
yCxFd41oPcX65u/ATbZ64wlLwEzBFPI2D+B/U1mtpHPeRkQ9lVGyHP+TB3zn4KBFMD/2sXYrxkFI
JpdNTrfHzMfisqbr4kqmSUgeUHZ6f5PTsWddLsn8lN9DmHPsi2qbvwQfjwal+xMf9yc90/EXDE8k
nIOoB2MM7Bi1rdMDV7fVilB35ShKWkPJ/YI6AjnI25bWdTxrwpcOBhDGejr67Rx7f2CHnNQXEa3r
VbaLa1bqTfTjOuuaREi6RmiokGW498hy5NOBekChkR5uSbD2jpxxsbQy+LHPWEdlz78j84N+zpAX
rB43DpcKmVDrULB3q8nm/FpCgO3K0kVC+VQurVXkYcfyDom1fWXhjcecfWo+WYPxqRx3ZR0mI0RU
idT+LSokiPThq5YeEY4zhaL6hh5l/PYyg3HtKWVbWozLwLT1jXZJFsqhkOaipo7VQLejtgbnN3Sg
jdOPLLjyueURc44yfnz9GfBOg+BctO7MlYH5jiZx90rBa7MbgCDbQguZJj4EgIaYJbyHGYlTXwJg
MO3mBrVnkbYI2nTZGqiyWCUk3k4Czsnw6Hyvkp/T5cN6c43qUCTJztYLTVN69y/nzCsrJ+VUqg5r
U9T+YQyjHOsGrAx2kFhgTYS9RSy0jP3iUQBLB5UXd5P3K1h2OuUyH0AfToRi4FWOaP6e7jxRgqms
2cQ05qZYQrFgTWLjKRmBw6ih65tPPv3uibF5a8Lcob52C6PUEVny7Zz+gPicFL5fNBWK3bEaJmRz
vGV9LAXSomwyeVmDjngXn/LSyB1g9DzGvhjFUsJ8/hZK1/61fB3gnX0PRqdyS0XlWbPBS2JmeLhV
6UOthHBdIunW13B2UyV8GVxIoIaoE/Ld/L7R6LR/S9XaAI3A2rwnyCPFkZgZ75FIShfcszJuAEQ3
AlV9Uaq8Q2n83ZFwGxGjqitWkRdBaLkRXB9qkVpqQAMLxGTiHY0D5gPBmsIlgLCpzGZfR1UIJ0GP
ouGnsvCYXLLJ8/imgBEYjrBgqygQYl2oed2cK872PyzNOZkS8qGz4/p5mATA7jq72ZzjLTVOlTae
vgviVnTXY77qfWTPzkxIR1RvkOIZyUpUbQIT8QPq0h+aGvsq/yOFAl78wyQSgbNdFTxn+uK3iaMh
ovSelQ3s9AlgG4ilIxAGQQW1s3868LNVywH4B7KYnBD3yqSUrdipHTtTG9n3LNHsm6CDLumL1r72
s/krQEQH+7/g06rikkQT3d0Z00zaHHffzgFgCn/JV8yXUZ/wBoNpPhDujO9IfatFiRZbPfgoOozu
RyZODFthtJfpRHYv10vx790TQW16suQhBtpiixRkp9cd9iTkf+q0Yjlac0UFCRBTuKKN6lIWEb5P
OMRe/ukTeEcJfknqEA8sfjrlCZYXuiS3U8sj/0mVFXj3BxfU+xJy/lE/I1DlZdHygKSgHaNRNB9q
Tynp1dzfk1jhYkTettsMkBBoqB052N+NRJbAVb0/DswaxwT93CXT5A6qWDceEIC98pA5SMijHM2U
FXCN236hfLv8/iXZ22An5+t50U9ryX3LfgjVyzInl3/A7Yg0vjlahjsFJSXZdP0VIyidF0qimRJo
6p6sA7Dh2UhBtJDokVMagh322JUO9kvzetwBqNXoyGH8zAJEY6CiPF7AxmrlB4Q9kW/lJAGo2p0c
cZSnbESw128pGnyBUcDVPbevrtaa3dMNpBi1AKAWU38cwVLhoVYE71k4xvUraQprjAjd82M3inYS
FtZvXW+iqM8Y2rH8BsEnYVoZTQnxptatLqAhvyjNmQ1tkv3izaYaPYw1eLXuG8VZm92nP3F1xyo2
uaTIBqYD6y1/p1yAIQ7Ykz0vgfYLoa/4SZrEdI2lSCWjvm+6K5HBF383dhRISCNOiMPVtF5p98/5
hDAO76FISzT2HNrTrH5dT/dCufrzEnY5/1rRgUurBGvYNgkwvrRYeG6OZnq1B1I9XXeforpRsgMn
pSouO+zo5HFrs8ybRbVqJp2glAgIwMEDki8Ztmn9zCzdtix6lkWss6E0+kAc0f8W3FnnxJ4pWzTL
//Z93fwfco0xhjtDyhmRhPOgafeZu+sGacIjPYnvIqUvXqPPK/PRwxKnd/MlVIbsdGu9nc+XtDoa
0UlXs9Pi0E3exA6/TKAUPsL89S8xrQM5MWyLGJv6hy84G6+38W4rvnkYJtHs2WpVb8q3FodozuW6
a+mzzbFtSHkErTXEgRAyUp+8KbYjPT0qkAxesXGo3r70sYO7EHAgEYKytkZB4Ou9gqM8qrJ5eISV
mMoGWoh/mEf3ApQSGtVEL3fLavDFYfeEo8AmTzG5rGKZyffrDqsTcKMqGpJAbQ6sMjXcDhCSQF0K
1/u+m6l4/RbDsBMTd4wWPVE5E4/2NXQJqSChv+B7DTXO8TaMG8cTFWCpgtynJo7b5Iv2Pf147OoE
O7iuc/8yK9LtQS3xPwEQ1OCD5YciMc2+CArXORcDvA0G/fjWQJkv0Qd729uLDwmXlVkVAbJZaBzn
BDahE84tlzXXERl1lA0Bb7DcCAl+Rj7lTwEUeeHOBntjg4uPhjIbRjSH2ki600Xh5WRyxWty1f2T
6yiTzPJW9jmt5nClRtAW6tPN1EnFEv6wi66Y4yhvaWPEMmxDcbwbGw31umJITGzE9pg4WbeJvPYz
eQ0dGfFyr+OVmb8w4kdSHbmZ+Xm14xSDFmBE5uCEr42+M/L7I533Ed4MAm878ow0Mt6+lncFUCMg
3TmQoC2HjpP20FqAga7/fNRUDXhDvrXe64uqR52By8RRdGXRDd22oo+LJudNz7T104x3nYVZyGcv
yxWeMAXJD+YAGm3qPi8ctHkG8UcyZ1kiPLplxXoI58FFFK8Na8/ZXwi5b4ovX4fkK/9XKq9Pg1uf
h8josRV0Wq4+U7FxFm/nFay4Zosg0cbpvIDNcW91SAN/Pgds+Uaie1IcBnpN4bxqM7Dsf2liHzEB
a7vMyaC88U73sBCnjRf0OuinHR5cutu+d9YTIOb9z3nZE6+dsZE8+RWjWTcwCD7FeSjjNC6/ZRIH
pxzLWZx8qUmBI+xboBT1P0l9SWX5eV+YEriHguQOxJJ+wuFtiGrHIEtJzQEyBT83Mkzopm/AkeDr
VUSCUnLNGsXOFmE8qV4eslTWwFtTubolhnqF3s/tRENRkqTrH8iYmqpV53fztCNMiMkyzUIQVRGG
KEq9KdnZJnFguoUhhKPhBQvzaFZyQkELqFeK/6YfulvH96zZA7lArSCbQasv3XgRuS5or1HricVt
/Tt/TWSc+zLZm5vXq1kFkKz3Zj8OW0zLPbX7g6FJGW+WoOp70lxaI33HSlt/P1hm+kuPd71sXnVt
O0NLEn5ltwJKKezIvaD2Jfd9v24r3pgXbQUEqPuf6sU4JrOAvioRyMHRsK/f51RXybPNpzwm8sec
FCg4oBDWL1Q3qL8ZShBWj3oiZmwoOvt3TtFcg8QcTFHFD2KjUhma2B5z95EpcYlA5r4NnKWN7CW3
BtoRN4Uj/ttJPRtRD0+p1+IiuFX3MT5IRbgHQUAMoWR0YfMdtHf6WfBLs5cklLTWUzZ/LFC+MP3j
SIYbhYCE/Y3DRFWVa+A+2hNAuUEq/rkfg62MTMPXOGvicC+AaUc2m5Zpgrf45L7p+I4lL1zXuJFS
EkJpzVznt/V9iCUO3n8hsCiae1KLtQniHFT9I6YhDj0W0WVnvYJHhchAkljuImA1gZU/TLf3Kudj
Irqim5JcrXu8i4KAciPK3sGur6+tDywWHz7sFbV75aFNRqME7w1G5Kt2L6zi+u2iEfh33hYs3guj
2fB2+xwculT1ffcV5nVsvhIZaeLa8gqeKOBm/cHpOOu27g3idDC9XQ+2Z3Wky8ME9GMTiRQfpUaJ
By4Zm/3AmPbozNyJCIoIxQ+lpxWR59XqC8Q2BbxELi563bq2AbdJmQbqi+cLP/rzt08W59Baz/v+
+2uYEsa70w+UAAlS7NMI0BxXXgiNHOlAge2JqZHII/rkclQXzHtZ0cCQK3NAsIVkx+IEazgY2GP/
i4ABQayy8MTTECWSh45y0TJFQmInQj2xi6tc9vhIUOgFtFffJQQ//Jj6UxoMPHCELtX1NeNYUJFM
xEsyfJBk+FeEKe04IiYAZZHIH7d5qoGk/Sci6ExEh4U37xDp5XyvJZZZMHW2pURT/xubG+WEmoUz
s/shY2RxIWCgZWY0UoyfSEotK7xiAYGYl3e6XkDJDKRrHh7aCofjHjtGomDPoZwk+NvzikoA1UdD
MyLUgT7v2f7/JLk7CtzR4ueW0VYOdpmrsXocWhMHgf2ByxhghJ54mvWzYgpFwKf9g6hmyWhSXKvn
84VMYKMoGK8mVQF/o9o1G883OdAbw4y1EN5FEKofBlOIbZsCz+zBct2qK3SbmBw0WM3Lw/8+5K1R
8LlCf1Jr7KymePvGRx/DURwtYRvlrFij9BAp9E1m0A4StJkKhtY9JB+eiz1kgEfWLT3gixFjvaMi
6w9/r6K41tucfXE+k0mf1vw8ruuH28vl9hqAVO73cOWyqxrJGJijsm3bsURTA52H4AT7sX1gjj9H
PdE54Ml7sIklIN3DDJ51J6qUm4CVcBUqDSIRMAkoCmKpcmWc1L3FjRJ7GHJI2XawvD7i5c25CKD0
BReAQMOae4lGc4byxsTuepdg5+LHOXTHmslheXeKzLNn3aUaiP+uh0Gj6QzEkRg/Cj2kvWaXDogz
3mLPcMmfFinXWxebUvXq6TzBt+LZ8dDyl5+2PFvbes2ZlZXiEcAWiVtZ+9/Zt8EVt3C1tmpilTw2
nCUYaxdB7tBonnsnfVjjxLJKUDkxkW8wzx3BkJ027I/iTBuR8d3oSRB3Lzr3Km/FL6oeWepEQKy8
AFJ+RNAvt3nrra2cOkrwReA1qNZbOtJbcNM8ebVx7HBl4t4FUYELs4qZfo21Wq/pxmcg6MVQ42vZ
Y9xdef/9LK7Vl96jVR+76nJOnmU9hScM68si6fpUZ8+1usJ6UgfUuTM3UYH8JNuFvFafyokXOY9W
oCj4EgGqHT12f4vWfFl/+llpIHARZ5AIEYbKrBe6REp5zo2Q1UXmMNbCsC9thEBMNGMXcBHvQHzV
3pyaec5J5JLc3bnsK2nCDFKlGR4sSDgjZ/R2/sfFsU3OB1c7R56Wbw9/WIMRjyHUWV0TXz6oErR6
KO0wtPt7LFrDuEPGpl4hWJoLvGOjw++FtG3Ec8dL13f4vq4JIe2IGSRtVzA/2qIQ5jJ9k3X0sjrv
Zq+B6Y6oCGw/aqE9vpt6sPEWLy6f7Xge83NgXAkXyYXC1LPKhhcl0fuE63QCo2nIblM3GzoXQ/6u
ZuoL9lT9mO4TTDzkSTvqZ6JPwbUeeJfX6sgCOPFxmUgXukZifnZyVtIpJIRmffRO7tPaz7G3UvF1
GHAhH4oR2D5nKNQc77+Sts7clixN+906rNjYlEyQRzhypOy1BllD2xamnr4xrkSf8kTlA7M47JnX
V8pa9AKJ526jUx01eWzu5/LPYmaX9RdtyCBT20kiyGLsPvxFqW6hvFbJ9961A/OM8lagYaW6/wDI
6QGXgYvjzOQhXMHvhX0aTGm2YGd2BEMj2+Om6l6hsf8hHv7HGH1uMQZtkmAdDeCBiPnCz+05QBtQ
NE5rRiWaRrJgMklcUkAdhsAr9eT7WUhD29I30slYEO9xwqDzRIshjvkxAQPxecoLTxY+CgUAy3qe
SH+vPFj21rH6/tLOhG3ME4fHqrRbjYCdfDr7+OiR8NFKtgUV9tUKpQ9GobAo7ho7Uo7PBUzhb3mP
n9Knhzp5XThtQyf5e6PHA9HYmIA/zunCP5w6wOFBcTTsxn6EVnJELhxvWk/HUc91XffjLb+L95pp
g8IijtLOt2KxRvjw6V3BDkfwZS4szYC8UsG/xNRLR15EhGesG8EGSMIT0TAGdz/LlD5EdiQ/tCqL
cDiuBK41sMf8US3pbd0THoFZOWeWpaCxfjMz7428DOJcKpub+i1O61oi4eoEJlpecSZ+NezmX9r0
WTolhsl2k0d+2I/1khEWdbqBeTYJQzTvAiBkPRyMaBWVaFcacw2Zj6XRdue8NI59WUhC8f+qcENt
WUfHH1Nv5f6Tkcdfi3OgQXd8TmgzL4arhLdRxVpYeJ4BfSDZE7yIcl2zE/wrIXEwCtX1hHjoFZmZ
C4Qgnm1T8w1M8W7+c0DiLaxlVJdOiOarP566uKvxqwmod3gpqZpC6f4OkqJuqX/G1sCiyLFlZT1C
frHlWfzMj19MPwHizbUccz2f5ozfzjt0iydLDYt8SN/g0rx4wUarJYutdEnBLwqG8fc6e7YHZ9N8
QfPAX8YEiMI4qDsoY7MEmv6A9pt2j0AP1M7qRXDudeWrwO5n9605AWFv3YvPdGQrcMk9c8YwRqwc
sExqmn9GTIQ70ji1q8IeNLO/0+Ie31czmgF0ySA+y8/7r8hYZLCu8KnfEeBgcqef5dHxuiEw80yz
wqdPf6UEtKXpYW2JCeedbRyTQ7gaPzdRlLGcK7yXnY+iXYUKPE4Mw52dl7SmrE8wKEqWD66xMBnO
W9zbh246zb5M3jYd+/vb0DCIOHK3QmrBu9WH+vlqYlA0dFcYi6uag/6N6f4zRck7/lmFoIthO2S4
2kjouvJIcReOAriw9OYSHQfwyrlBrftWP+WgH63PQJCQGur+fX9EssJOwF6K9K1tsCk1rHJbOvDo
bnd4IiLB89LAjNjRpFT955DyKDBOD/5GhtzZP1mOmrxQ5AW5M714hFssEQyYGc+jQ1xAzu2jpKec
3hDOgFsM025kNPYBC92pozBroOvGSILPfTGstIHc6W4eRBIORqR8yXJGR7AlO559RHZaYWHqO0P/
A8CVjx7cyLvVdPCduEGl0bwZlv0KWQlKkXO3A1j9abVahYKJ45aN7rcq9rzxbr3iG2L14/MzGjbv
VmVDHsrSq0KKTI5aAH1ZLCBcnu18XZV8EyTv1wAWACiHvGPEFqC72Yqr7PLmnHQSlRXl4Wb/idsZ
c6o2T7oElVr8DRH19PuUkOnFk/BijH+tqQ7+1yBkDWhsT2fjgvMJi54lwaUGDDnplNY6ysTd6Zt3
IHptTUCoDNiVqYrpIRNMJaX/TkAVJmXgFOi3W+FHfREyzvY/o9vQCUsW5RkLBLMf7Eh8hq2XJ/y2
802EAKl5GPGo6xcfom/fk8Dp3pDUnu4GszyTHWD4rIIOiS5qr7Xz/dMRoOFS9fCQ3ruKjq0VWNfG
yl5IwdyCzSkBOquPJSRDUt6QbjNZpx2x+cmKqRfw5yhwkKMfrVpoPL9ze8ioG0NP+Sh+v+kA5O+H
WqIDLrvPMHENgELH8qWmEoQ6LmMlRjQOSZDYXAsRUS8l0NDS2TK+XLb3f4cCfFE16eWdOU/cyqT8
f/9mXMcwAFcuoUo86d4LweDimNLJT1Qv0E25mZv1zmiw46ZuoRPSiv8e4+k+Va1rwn+gDRA8eLkr
TG3cfWnKVTga0mGtxyo7LM+qrr3dJ6ISFJzNIP9AhWbBWdK9RAVH/dqr+fbwg3KyTzgV7EaAmhMl
BxZbf7ab9L1OtJPYQ13XvsOcpgYTrkHFh4pWJikbkMxLR3ml9kIZ0I+6y5HVw9dez/oYxQ783qu/
odm6wVeIh9fBOCwsEMOEYAp733GGR9QCCljhbD6FKomD6AKXQcZsyjtBZFWxUPAk57UAge9crPpZ
l8qvP6xJFP9JVMc/Ync0bug+iObM3tAk2ZHA0m3pozN+rJqwBIK4sCO884Axput2TvtVHWvLqlU2
diQjmxICO18WIyby3qNXukrDw71zqzQd99RgvZ5BA/x7sqXbObFmro/Gg35UgbMiJKTBG8teQbGw
fCtDfR/PkhWMg0502cQM7FcVCxhZn/D7ANeh30FrU9ZirLi35vPG+RWWuVANxdFvjkFqw0OIkYHZ
/Z8Q1xRRtu7l5L2faP4E3syRa+Pdd2Nlp4WJZ58gp6swn6TZq3KjR4+fShyAkM8CxbfzIa/uqJZU
iHdSfdU4j9Hy+XopYwDfjYLV4bbWq4mdoHXViWAD29lptrLTB1kRbnGCd4Bmtn/8FAImRmFlM3vA
eSV3isqBH+9yVJOUeiyIpLjEka8oPoOw0h9P7G6jvZXLIaMgjEhklhMV+xsO+pQuKTXZJpi1FjHs
SrD/BUjTKepwLX9dtLl7cnJQ0UeiuIaJ1qQXSPr6OqJP1pkMqcnoiPlV/Gr8XZ16ODIPXGriB6cF
KzBLo+E5Orm96Fzt546vsHrzdSZTHNHUkIr/sm/k4IquBLfLRdU7NDx9uJ32E0hhcYwVh13Plmer
tKULafwANp/44lfHhEfv24L92sPICjiVIRF3NpBkgcXeK60fnq8GJhBu7l9gJIPWBvYbemqtqGAF
JivJFwBbOXe9ZE1+OkXJH8b1ZUAseRHdTkMeRcIEFz5bVbxouWgSb8IBL5plPBtCiAW6tdi6SaTY
7cABiaYzZM74D56Y0FhczM507p9H6DfGn6zPzTAqD8QJ946uf7O3q6g13pzeJrJu2o2JY9bLd5Q+
nMODoSUwkfGUr+UtWfdazpPShhjZJfdQAivAgFw0YCwLHZhRdkGrB04xfTFDy6gi1Vm6irIpP8ks
TvLLHbYKr5zTH+e/DV4K5hLFN2FpmZXLpDdYg+qY+YDAQ+wF/IQCabcspL2QxjPBv06csQXnSN8W
bBHUZo8U4a9zV5yWdoRTGH086GytqB0juPN08gsaZjazK+jwJit62YJusxfh/SkrH8khHa9WVq73
t018KtWGKDjUnQidzwvxrQSuZnRPeHXxUm0Om45qPtzYeVictR3+KwX9t+r4+reoTUcL1UqB5aaR
Zss6PErR6m4TnQGKwDqso619O1zngoW6H48IDWOJdDrwVmshFYPQMkn1O6Gl1Kub/bMYg4fPFW+u
yCZkf79nFsqEVLC895V3gp9CdsmXEtg0/cWOsQqZQFfsygg0DLdzRgxUCiq+QfTiSs3JNEkMoQTw
skBlwFM76ZIqv/YzMCtjbbj7v8/r8CKfKZGoWSnNfj3H6lu3HuoTMmOJs+NEnllR+W6TDPO6qle1
HH9zVpMp6udFw49KtAcGiIllgZdMhRtGiVQ5yQEd0V76jpq9RsdnZfwsAqK1fzjV+vt+9PfJcl6+
ViWOWKTpIivcaaCwRlfBCIGCcFQVxBsacGpQo8M7AnmWt21uLFUrA9VQw1Cl0Vd0EKbYDb/ZVltn
Me9rc1RPgt64Qf5R+q42kr82nWw7aeC0S3hQYK4KFhDNfSEOX29KkrSYHDN+v0fBDGar5QzcjAiY
uCwGp25a5bcJLs30ctF9FvwJCLGgjw4Aiuhdst4PlcUIguIiD9nXqHgBeui78S9RcY6iY7UHuaXM
aE1VYv8e+wXLX+91HCxdc7NLJgkKvkGb7fCmTbLfaWR2doK/Ma1I2F8Kd4dAM7Rtiq5zYMckl0vE
PkaxzSCXzbq+2BaqyRkBkaF7uKCiH0aaQf/pTRt5DMSlDMBwSxryqqPDPeFPivlviajWlHBCalQ+
OEIOmYO3JyeIsNYBCW51OrNSVM18BxAryGpzvOiMf3Z2bbLBQz7/5QWZRPs9bgnnewCK8SpiAUrE
qqgfdXwNrRpQt9B6mZghYU7TXg/jJun9ex3tujhjE0EnfU6oA/O6/xI26tdj8+Yk/SW2c0CvtW0M
jEwEuSn1t9seP2YlnE4qApwnd+2yjhZnmyP9PND7YCoGzEjWkYoCWSJ2FvMOG/uL1rPEPwd/lz4x
NSJ9kuNw/Tkf74boUBhBTmpn0coNw/nL2KpI2jWW2SUIT3X2LuF+/ZmaxL60ze2rqfWyDTOEopKw
ZJTvMBFAmVbJrK/ML0pt/iA5WWoFDLyebdRS+tXiKwLM0jdUhyXfoEnNT+s9iUxhqA==
`protect end_protected

